library verilog;
use verilog.vl_types.all;
entity xor_boh_tb is
end xor_boh_tb;
