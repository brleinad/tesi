module enc_lut(s,enc_s);
`include "constants.v"

input [NBIT:0] s;
output reg [NBIT:0] enc_s;
always @(*)
begin
    case(s)
	0 : enc_s = 0;
	1 : enc_s = 256;
	2 : enc_s = 128;
	3 : enc_s = 384;
	4 : enc_s = 64;
	5 : enc_s = 320;
	6 : enc_s = 288;
	7 : enc_s = 448;
	8 : enc_s = 32;
	9 : enc_s = 272;
	10 : enc_s = 264;
	11 : enc_s = 416;
	12 : enc_s = 260;
	13 : enc_s = 400;
	14 : enc_s = 392;
	15 : enc_s = 480;
	16 : enc_s = 8;
	17 : enc_s = 258;
	18 : enc_s = 257;
	19 : enc_s = 388;
	20 : enc_s = 192;
	21 : enc_s = 386;
	22 : enc_s = 385;
	23 : enc_s = 464;
	24 : enc_s = 160;
	25 : enc_s = 352;
	26 : enc_s = 336;
	27 : enc_s = 456;
	28 : enc_s = 328;
	29 : enc_s = 452;
	30 : enc_s = 450;
	31 : enc_s = 496;
	32 : enc_s = 16;
	33 : enc_s = 144;
	34 : enc_s = 136;
	35 : enc_s = 324;
	36 : enc_s = 132;
	37 : enc_s = 322;
	38 : enc_s = 321;
	39 : enc_s = 449;
	40 : enc_s = 130;
	41 : enc_s = 304;
	42 : enc_s = 296;
	43 : enc_s = 432;
	44 : enc_s = 292;
	45 : enc_s = 424;
	46 : enc_s = 420;
	47 : enc_s = 488;
	48 : enc_s = 129;
	49 : enc_s = 290;
	50 : enc_s = 289;
	51 : enc_s = 418;
	52 : enc_s = 280;
	53 : enc_s = 417;
	54 : enc_s = 408;
	55 : enc_s = 484;
	56 : enc_s = 276;
	57 : enc_s = 404;
	58 : enc_s = 402;
	59 : enc_s = 482;
	60 : enc_s = 401;
	61 : enc_s = 481;
	62 : enc_s = 472;
	63 : enc_s = 504;
	64 : enc_s = 4;
	65 : enc_s = 96;
	66 : enc_s = 80;
	67 : enc_s = 274;
	68 : enc_s = 72;
	69 : enc_s = 273;
	70 : enc_s = 268;
	71 : enc_s = 396;
	72 : enc_s = 68;
	73 : enc_s = 266;
	74 : enc_s = 265;
	75 : enc_s = 394;
	76 : enc_s = 262;
	77 : enc_s = 393;
	78 : enc_s = 390;
	79 : enc_s = 468;
	80 : enc_s = 66;
	81 : enc_s = 261;
	82 : enc_s = 259;
	83 : enc_s = 389;
	84 : enc_s = 224;
	85 : enc_s = 387;
	86 : enc_s = 368;
	87 : enc_s = 466;
	88 : enc_s = 208;
	89 : enc_s = 360;
	90 : enc_s = 356;
	91 : enc_s = 465;
	92 : enc_s = 354;
	93 : enc_s = 460;
	94 : enc_s = 458;
	95 : enc_s = 500;
	96 : enc_s = 65;
	97 : enc_s = 200;
	98 : enc_s = 196;
	99 : enc_s = 353;
	100 : enc_s = 194;
	101 : enc_s = 344;
	102 : enc_s = 340;
	103 : enc_s = 457;
	104 : enc_s = 193;
	105 : enc_s = 338;
	106 : enc_s = 337;
	107 : enc_s = 454;
	108 : enc_s = 332;
	109 : enc_s = 453;
	110 : enc_s = 451;
	111 : enc_s = 498;
	112 : enc_s = 176;
	113 : enc_s = 330;
	114 : enc_s = 329;
	115 : enc_s = 440;
	116 : enc_s = 326;
	117 : enc_s = 436;
	118 : enc_s = 434;
	119 : enc_s = 497;
	120 : enc_s = 325;
	121 : enc_s = 433;
	122 : enc_s = 428;
	123 : enc_s = 492;
	124 : enc_s = 426;
	125 : enc_s = 490;
	126 : enc_s = 489;
	127 : enc_s = 508;
	128 : enc_s = 2;
	129 : enc_s = 48;
	130 : enc_s = 40;
	131 : enc_s = 168;
	132 : enc_s = 36;
	133 : enc_s = 164;
	134 : enc_s = 162;
	135 : enc_s = 323;
	136 : enc_s = 34;
	137 : enc_s = 161;
	138 : enc_s = 152;
	139 : enc_s = 312;
	140 : enc_s = 148;
	141 : enc_s = 308;
	142 : enc_s = 306;
	143 : enc_s = 425;
	144 : enc_s = 33;
	145 : enc_s = 146;
	146 : enc_s = 145;
	147 : enc_s = 305;
	148 : enc_s = 140;
	149 : enc_s = 300;
	150 : enc_s = 298;
	151 : enc_s = 422;
	152 : enc_s = 138;
	153 : enc_s = 297;
	154 : enc_s = 294;
	155 : enc_s = 421;
	156 : enc_s = 293;
	157 : enc_s = 419;
	158 : enc_s = 412;
	159 : enc_s = 486;
	160 : enc_s = 24;
	161 : enc_s = 137;
	162 : enc_s = 134;
	163 : enc_s = 291;
	164 : enc_s = 133;
	165 : enc_s = 284;
	166 : enc_s = 282;
	167 : enc_s = 410;
	168 : enc_s = 131;
	169 : enc_s = 281;
	170 : enc_s = 278;
	171 : enc_s = 409;
	172 : enc_s = 277;
	173 : enc_s = 406;
	174 : enc_s = 405;
	175 : enc_s = 485;
	176 : enc_s = 112;
	177 : enc_s = 275;
	178 : enc_s = 270;
	179 : enc_s = 403;
	180 : enc_s = 269;
	181 : enc_s = 398;
	182 : enc_s = 397;
	183 : enc_s = 483;
	184 : enc_s = 267;
	185 : enc_s = 395;
	186 : enc_s = 391;
	187 : enc_s = 476;
	188 : enc_s = 376;
	189 : enc_s = 474;
	190 : enc_s = 473;
	191 : enc_s = 506;
	192 : enc_s = 20;
	193 : enc_s = 104;
	194 : enc_s = 100;
	195 : enc_s = 263;
	196 : enc_s = 98;
	197 : enc_s = 240;
	198 : enc_s = 232;
	199 : enc_s = 372;
	200 : enc_s = 97;
	201 : enc_s = 228;
	202 : enc_s = 226;
	203 : enc_s = 370;
	204 : enc_s = 225;
	205 : enc_s = 369;
	206 : enc_s = 364;
	207 : enc_s = 470;
	208 : enc_s = 88;
	209 : enc_s = 216;
	210 : enc_s = 212;
	211 : enc_s = 362;
	212 : enc_s = 210;
	213 : enc_s = 361;
	214 : enc_s = 358;
	215 : enc_s = 469;
	216 : enc_s = 209;
	217 : enc_s = 357;
	218 : enc_s = 355;
	219 : enc_s = 467;
	220 : enc_s = 348;
	221 : enc_s = 462;
	222 : enc_s = 461;
	223 : enc_s = 505;
	224 : enc_s = 84;
	225 : enc_s = 204;
	226 : enc_s = 202;
	227 : enc_s = 346;
	228 : enc_s = 201;
	229 : enc_s = 345;
	230 : enc_s = 342;
	231 : enc_s = 459;
	232 : enc_s = 198;
	233 : enc_s = 341;
	234 : enc_s = 339;
	235 : enc_s = 455;
	236 : enc_s = 334;
	237 : enc_s = 444;
	238 : enc_s = 442;
	239 : enc_s = 502;
	240 : enc_s = 197;
	241 : enc_s = 333;
	242 : enc_s = 331;
	243 : enc_s = 441;
	244 : enc_s = 327;
	245 : enc_s = 438;
	246 : enc_s = 437;
	247 : enc_s = 501;
	248 : enc_s = 316;
	249 : enc_s = 435;
	250 : enc_s = 430;
	251 : enc_s = 499;
	252 : enc_s = 429;
	253 : enc_s = 494;
	254 : enc_s = 493;
	255 : enc_s = 510;
	256 : enc_s = 1;
	257 : enc_s = 18;
	258 : enc_s = 17;
	259 : enc_s = 82;
	260 : enc_s = 12;
	261 : enc_s = 81;
	262 : enc_s = 76;
	263 : enc_s = 195;
	264 : enc_s = 10;
	265 : enc_s = 74;
	266 : enc_s = 73;
	267 : enc_s = 184;
	268 : enc_s = 70;
	269 : enc_s = 180;
	270 : enc_s = 178;
	271 : enc_s = 314;
	272 : enc_s = 9;
	273 : enc_s = 69;
	274 : enc_s = 67;
	275 : enc_s = 177;
	276 : enc_s = 56;
	277 : enc_s = 172;
	278 : enc_s = 170;
	279 : enc_s = 313;
	280 : enc_s = 52;
	281 : enc_s = 169;
	282 : enc_s = 166;
	283 : enc_s = 310;
	284 : enc_s = 165;
	285 : enc_s = 309;
	286 : enc_s = 307;
	287 : enc_s = 427;
	288 : enc_s = 6;
	289 : enc_s = 50;
	290 : enc_s = 49;
	291 : enc_s = 163;
	292 : enc_s = 44;
	293 : enc_s = 156;
	294 : enc_s = 154;
	295 : enc_s = 302;
	296 : enc_s = 42;
	297 : enc_s = 153;
	298 : enc_s = 150;
	299 : enc_s = 301;
	300 : enc_s = 149;
	301 : enc_s = 299;
	302 : enc_s = 295;
	303 : enc_s = 423;
	304 : enc_s = 41;
	305 : enc_s = 147;
	306 : enc_s = 142;
	307 : enc_s = 286;
	308 : enc_s = 141;
	309 : enc_s = 285;
	310 : enc_s = 283;
	311 : enc_s = 414;
	312 : enc_s = 139;
	313 : enc_s = 279;
	314 : enc_s = 271;
	315 : enc_s = 413;
	316 : enc_s = 248;
	317 : enc_s = 411;
	318 : enc_s = 407;
	319 : enc_s = 491;
	320 : enc_s = 5;
	321 : enc_s = 38;
	322 : enc_s = 37;
	323 : enc_s = 135;
	324 : enc_s = 35;
	325 : enc_s = 120;
	326 : enc_s = 116;
	327 : enc_s = 244;
	328 : enc_s = 28;
	329 : enc_s = 114;
	330 : enc_s = 113;
	331 : enc_s = 242;
	332 : enc_s = 108;
	333 : enc_s = 241;
	334 : enc_s = 236;
	335 : enc_s = 399;
	336 : enc_s = 26;
	337 : enc_s = 106;
	338 : enc_s = 105;
	339 : enc_s = 234;
	340 : enc_s = 102;
	341 : enc_s = 233;
	342 : enc_s = 230;
	343 : enc_s = 380;
	344 : enc_s = 101;
	345 : enc_s = 229;
	346 : enc_s = 227;
	347 : enc_s = 378;
	348 : enc_s = 220;
	349 : enc_s = 377;
	350 : enc_s = 374;
	351 : enc_s = 487;
	352 : enc_s = 25;
	353 : enc_s = 99;
	354 : enc_s = 92;
	355 : enc_s = 218;
	356 : enc_s = 90;
	357 : enc_s = 217;
	358 : enc_s = 214;
	359 : enc_s = 373;
	360 : enc_s = 89;
	361 : enc_s = 213;
	362 : enc_s = 211;
	363 : enc_s = 371;
	364 : enc_s = 206;
	365 : enc_s = 366;
	366 : enc_s = 365;
	367 : enc_s = 478;
	368 : enc_s = 86;
	369 : enc_s = 205;
	370 : enc_s = 203;
	371 : enc_s = 363;
	372 : enc_s = 199;
	373 : enc_s = 359;
	374 : enc_s = 350;
	375 : enc_s = 477;
	376 : enc_s = 188;
	377 : enc_s = 349;
	378 : enc_s = 347;
	379 : enc_s = 475;
	380 : enc_s = 343;
	381 : enc_s = 471;
	382 : enc_s = 463;
	383 : enc_s = 509;
	384 : enc_s = 3;
	385 : enc_s = 22;
	386 : enc_s = 21;
	387 : enc_s = 85;
	388 : enc_s = 19;
	389 : enc_s = 83;
	390 : enc_s = 78;
	391 : enc_s = 186;
	392 : enc_s = 14;
	393 : enc_s = 77;
	394 : enc_s = 75;
	395 : enc_s = 185;
	396 : enc_s = 71;
	397 : enc_s = 182;
	398 : enc_s = 181;
	399 : enc_s = 335;
	400 : enc_s = 13;
	401 : enc_s = 60;
	402 : enc_s = 58;
	403 : enc_s = 179;
	404 : enc_s = 57;
	405 : enc_s = 174;
	406 : enc_s = 173;
	407 : enc_s = 318;
	408 : enc_s = 54;
	409 : enc_s = 171;
	410 : enc_s = 167;
	411 : enc_s = 317;
	412 : enc_s = 158;
	413 : enc_s = 315;
	414 : enc_s = 311;
	415 : enc_s = 446;
	416 : enc_s = 11;
	417 : enc_s = 53;
	418 : enc_s = 51;
	419 : enc_s = 157;
	420 : enc_s = 46;
	421 : enc_s = 155;
	422 : enc_s = 151;
	423 : enc_s = 303;
	424 : enc_s = 45;
	425 : enc_s = 143;
	426 : enc_s = 124;
	427 : enc_s = 287;
	428 : enc_s = 122;
	429 : enc_s = 252;
	430 : enc_s = 250;
	431 : enc_s = 445;
	432 : enc_s = 43;
	433 : enc_s = 121;
	434 : enc_s = 118;
	435 : enc_s = 249;
	436 : enc_s = 117;
	437 : enc_s = 246;
	438 : enc_s = 245;
	439 : enc_s = 443;
	440 : enc_s = 115;
	441 : enc_s = 243;
	442 : enc_s = 238;
	443 : enc_s = 439;
	444 : enc_s = 237;
	445 : enc_s = 431;
	446 : enc_s = 415;
	447 : enc_s = 507;
	448 : enc_s = 7;
	449 : enc_s = 39;
	450 : enc_s = 30;
	451 : enc_s = 110;
	452 : enc_s = 29;
	453 : enc_s = 109;
	454 : enc_s = 107;
	455 : enc_s = 235;
	456 : enc_s = 27;
	457 : enc_s = 103;
	458 : enc_s = 94;
	459 : enc_s = 231;
	460 : enc_s = 93;
	461 : enc_s = 222;
	462 : enc_s = 221;
	463 : enc_s = 382;
	464 : enc_s = 23;
	465 : enc_s = 91;
	466 : enc_s = 87;
	467 : enc_s = 219;
	468 : enc_s = 79;
	469 : enc_s = 215;
	470 : enc_s = 207;
	471 : enc_s = 381;
	472 : enc_s = 62;
	473 : enc_s = 190;
	474 : enc_s = 189;
	475 : enc_s = 379;
	476 : enc_s = 187;
	477 : enc_s = 375;
	478 : enc_s = 367;
	479 : enc_s = 503;
	480 : enc_s = 15;
	481 : enc_s = 61;
	482 : enc_s = 59;
	483 : enc_s = 183;
	484 : enc_s = 55;
	485 : enc_s = 175;
	486 : enc_s = 159;
	487 : enc_s = 351;
	488 : enc_s = 47;
	489 : enc_s = 126;
	490 : enc_s = 125;
	491 : enc_s = 319;
	492 : enc_s = 123;
	493 : enc_s = 254;
	494 : enc_s = 253;
	495 : enc_s = 479;
	496 : enc_s = 31;
	497 : enc_s = 119;
	498 : enc_s = 111;
	499 : enc_s = 251;
	500 : enc_s = 95;
	501 : enc_s = 247;
	502 : enc_s = 239;
	503 : enc_s = 495;
	504 : enc_s = 63;
	505 : enc_s = 223;
	506 : enc_s = 191;
	507 : enc_s = 447;
	508 : enc_s = 127;
	509 : enc_s = 383;
	510 : enc_s = 255;
	default : enc_s = 0;
    endcase
end
endmodule
