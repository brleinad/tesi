
module gen_linear_part ( a, b, n, s );
  input [9:0] a;
  input [9:0] b;
  input [2034:0] n;
  output [9:0] s;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724;

  XOR4D0 U1 ( .A1(b[9]), .A2(a[9]), .A3(n1), .A4(n2), .Z(s[9]) );
  XOR4D0 U2 ( .A1(n[2028]), .A2(n3), .A3(n[2030]), .A4(n[2029]), .Z(n2) );
  XOR4D0 U3 ( .A1(n[2023]), .A2(n[2022]), .A3(n4), .A4(n5), .Z(n3) );
  XOR3D0 U4 ( .A1(n6), .A2(n7), .A3(n[2021]), .Z(n5) );
  XOR4D0 U5 ( .A1(n[2014]), .A2(n8), .A3(n[2016]), .A4(n[2015]), .Z(n7) );
  XOR4D0 U6 ( .A1(n[2009]), .A2(n[2008]), .A3(n9), .A4(n10), .Z(n8) );
  XOR3D0 U7 ( .A1(n11), .A2(n12), .A3(n[2007]), .Z(n10) );
  XOR4D0 U8 ( .A1(n[2000]), .A2(n13), .A3(n[2002]), .A4(n[2001]), .Z(n12) );
  XOR4D0 U9 ( .A1(n[1995]), .A2(n[1994]), .A3(n14), .A4(n15), .Z(n13) );
  XOR3D0 U10 ( .A1(n16), .A2(n17), .A3(n[1993]), .Z(n15) );
  XOR4D0 U11 ( .A1(n[1986]), .A2(n18), .A3(n[1988]), .A4(n[1987]), .Z(n17) );
  XOR4D0 U12 ( .A1(n[1981]), .A2(n[1980]), .A3(n19), .A4(n20), .Z(n18) );
  XOR3D0 U13 ( .A1(n21), .A2(n22), .A3(n[1979]), .Z(n20) );
  XOR4D0 U14 ( .A1(n[1972]), .A2(n23), .A3(n[1974]), .A4(n[1973]), .Z(n22) );
  XOR4D0 U15 ( .A1(n[1967]), .A2(n[1966]), .A3(n24), .A4(n25), .Z(n23) );
  XOR3D0 U16 ( .A1(n26), .A2(n27), .A3(n[1965]), .Z(n25) );
  XOR4D0 U17 ( .A1(n[1958]), .A2(n28), .A3(n[1960]), .A4(n[1959]), .Z(n27) );
  XOR4D0 U18 ( .A1(n[1953]), .A2(n[1952]), .A3(n29), .A4(n30), .Z(n28) );
  XOR3D0 U19 ( .A1(n31), .A2(n32), .A3(n[1951]), .Z(n30) );
  XOR4D0 U20 ( .A1(n[1944]), .A2(n33), .A3(n[1946]), .A4(n[1945]), .Z(n32) );
  XOR4D0 U21 ( .A1(n[1939]), .A2(n[1938]), .A3(n34), .A4(n35), .Z(n33) );
  XOR3D0 U22 ( .A1(n36), .A2(n37), .A3(n[1937]), .Z(n35) );
  XOR4D0 U23 ( .A1(n[1930]), .A2(n38), .A3(n[1932]), .A4(n[1931]), .Z(n37) );
  XOR4D0 U24 ( .A1(n[1925]), .A2(n[1924]), .A3(n39), .A4(n40), .Z(n38) );
  XOR3D0 U25 ( .A1(n41), .A2(n42), .A3(n[1923]), .Z(n40) );
  XOR4D0 U26 ( .A1(n[1916]), .A2(n43), .A3(n[1918]), .A4(n[1917]), .Z(n42) );
  XOR4D0 U27 ( .A1(n[1911]), .A2(n[1910]), .A3(n44), .A4(n45), .Z(n43) );
  XOR3D0 U28 ( .A1(n46), .A2(n47), .A3(n[1909]), .Z(n45) );
  XOR4D0 U29 ( .A1(n[1902]), .A2(n48), .A3(n[1904]), .A4(n[1903]), .Z(n47) );
  XOR4D0 U30 ( .A1(n[1897]), .A2(n[1896]), .A3(n49), .A4(n50), .Z(n48) );
  XOR3D0 U31 ( .A1(n51), .A2(n52), .A3(n[1895]), .Z(n50) );
  XOR4D0 U32 ( .A1(n[1888]), .A2(n53), .A3(n[1890]), .A4(n[1889]), .Z(n52) );
  XOR4D0 U33 ( .A1(n[1883]), .A2(n[1882]), .A3(n54), .A4(n55), .Z(n53) );
  XOR3D0 U34 ( .A1(n56), .A2(n57), .A3(n[1881]), .Z(n55) );
  XOR4D0 U35 ( .A1(n[1874]), .A2(n58), .A3(n[1876]), .A4(n[1875]), .Z(n57) );
  XOR4D0 U36 ( .A1(n[1869]), .A2(n[1868]), .A3(n59), .A4(n60), .Z(n58) );
  XOR3D0 U37 ( .A1(n61), .A2(n62), .A3(n[1867]), .Z(n60) );
  XOR4D0 U38 ( .A1(n[1860]), .A2(n63), .A3(n[1862]), .A4(n[1861]), .Z(n62) );
  XOR4D0 U39 ( .A1(n[1855]), .A2(n[1854]), .A3(n64), .A4(n65), .Z(n63) );
  XOR3D0 U40 ( .A1(n66), .A2(n67), .A3(n[1853]), .Z(n65) );
  XOR4D0 U41 ( .A1(n[1846]), .A2(n68), .A3(n[1848]), .A4(n[1847]), .Z(n67) );
  XOR4D0 U42 ( .A1(n[1841]), .A2(n[1840]), .A3(n69), .A4(n70), .Z(n68) );
  XOR3D0 U43 ( .A1(n71), .A2(n72), .A3(n[1839]), .Z(n70) );
  XOR4D0 U44 ( .A1(n[1832]), .A2(n73), .A3(n[1834]), .A4(n[1833]), .Z(n72) );
  XOR4D0 U45 ( .A1(n[1827]), .A2(n[1826]), .A3(n74), .A4(n75), .Z(n73) );
  XOR3D0 U46 ( .A1(n76), .A2(n77), .A3(n[1825]), .Z(n75) );
  XOR4D0 U47 ( .A1(n[1818]), .A2(n78), .A3(n[1820]), .A4(n[1819]), .Z(n77) );
  XOR4D0 U48 ( .A1(n[1813]), .A2(n[1812]), .A3(n79), .A4(n80), .Z(n78) );
  XOR3D0 U49 ( .A1(n81), .A2(n82), .A3(n[1811]), .Z(n80) );
  XOR4D0 U50 ( .A1(n[1804]), .A2(n83), .A3(n[1806]), .A4(n[1805]), .Z(n82) );
  XOR4D0 U51 ( .A1(n[1799]), .A2(n[1798]), .A3(n84), .A4(n85), .Z(n83) );
  XOR3D0 U52 ( .A1(n86), .A2(n87), .A3(n[1797]), .Z(n85) );
  XOR4D0 U53 ( .A1(n[1790]), .A2(n88), .A3(n[1792]), .A4(n[1791]), .Z(n87) );
  XOR4D0 U54 ( .A1(n[1785]), .A2(n[1784]), .A3(n89), .A4(n90), .Z(n88) );
  XOR3D0 U55 ( .A1(n91), .A2(n92), .A3(n[1783]), .Z(n90) );
  XOR4D0 U56 ( .A1(n[1776]), .A2(n93), .A3(n[1778]), .A4(n[1777]), .Z(n92) );
  XOR4D0 U57 ( .A1(n[1771]), .A2(n[1770]), .A3(n94), .A4(n95), .Z(n93) );
  XOR3D0 U58 ( .A1(n96), .A2(n97), .A3(n[1769]), .Z(n95) );
  XOR4D0 U59 ( .A1(n[1762]), .A2(n98), .A3(n[1764]), .A4(n[1763]), .Z(n97) );
  XOR4D0 U60 ( .A1(n[1757]), .A2(n[1756]), .A3(n99), .A4(n100), .Z(n98) );
  XOR3D0 U61 ( .A1(n101), .A2(n102), .A3(n[1755]), .Z(n100) );
  XOR4D0 U62 ( .A1(n[1748]), .A2(n103), .A3(n[1750]), .A4(n[1749]), .Z(n102)
         );
  XOR4D0 U63 ( .A1(n[1743]), .A2(n[1742]), .A3(n104), .A4(n105), .Z(n103) );
  XOR3D0 U64 ( .A1(n106), .A2(n107), .A3(n[1741]), .Z(n105) );
  XOR4D0 U65 ( .A1(n[1734]), .A2(n108), .A3(n[1736]), .A4(n[1735]), .Z(n107)
         );
  XOR4D0 U66 ( .A1(n[1729]), .A2(n[1728]), .A3(n109), .A4(n110), .Z(n108) );
  XOR3D0 U67 ( .A1(n111), .A2(n112), .A3(n[1727]), .Z(n110) );
  XOR4D0 U68 ( .A1(n[1720]), .A2(n113), .A3(n[1722]), .A4(n[1721]), .Z(n112)
         );
  XOR4D0 U69 ( .A1(n[1715]), .A2(n[1714]), .A3(n114), .A4(n115), .Z(n113) );
  XOR3D0 U70 ( .A1(n116), .A2(n117), .A3(n[1713]), .Z(n115) );
  XOR4D0 U71 ( .A1(n[1706]), .A2(n118), .A3(n[1708]), .A4(n[1707]), .Z(n117)
         );
  XOR4D0 U72 ( .A1(n[1701]), .A2(n[1700]), .A3(n119), .A4(n120), .Z(n118) );
  XOR3D0 U73 ( .A1(n121), .A2(n122), .A3(n[1699]), .Z(n120) );
  XOR4D0 U74 ( .A1(n[1692]), .A2(n123), .A3(n[1694]), .A4(n[1693]), .Z(n122)
         );
  XOR4D0 U75 ( .A1(n[1687]), .A2(n[1686]), .A3(n124), .A4(n125), .Z(n123) );
  XOR3D0 U76 ( .A1(n126), .A2(n127), .A3(n[1685]), .Z(n125) );
  XOR4D0 U77 ( .A1(n[1678]), .A2(n128), .A3(n[1680]), .A4(n[1679]), .Z(n127)
         );
  XOR4D0 U78 ( .A1(n[1673]), .A2(n[1672]), .A3(n129), .A4(n130), .Z(n128) );
  XOR3D0 U79 ( .A1(n131), .A2(n132), .A3(n[1671]), .Z(n130) );
  XOR4D0 U80 ( .A1(n[1664]), .A2(n133), .A3(n[1666]), .A4(n[1665]), .Z(n132)
         );
  XOR4D0 U81 ( .A1(n[1659]), .A2(n[1658]), .A3(n134), .A4(n135), .Z(n133) );
  XOR3D0 U82 ( .A1(n136), .A2(n137), .A3(n[1657]), .Z(n135) );
  XOR4D0 U83 ( .A1(n[1650]), .A2(n138), .A3(n[1652]), .A4(n[1651]), .Z(n137)
         );
  XOR4D0 U84 ( .A1(n[1645]), .A2(n[1644]), .A3(n139), .A4(n140), .Z(n138) );
  XOR3D0 U85 ( .A1(n141), .A2(n142), .A3(n[1643]), .Z(n140) );
  XOR4D0 U86 ( .A1(n[1636]), .A2(n143), .A3(n[1638]), .A4(n[1637]), .Z(n142)
         );
  XOR4D0 U87 ( .A1(n[1631]), .A2(n[1630]), .A3(n144), .A4(n145), .Z(n143) );
  XOR3D0 U88 ( .A1(n146), .A2(n147), .A3(n[1629]), .Z(n145) );
  XOR4D0 U89 ( .A1(n[1622]), .A2(n148), .A3(n[1624]), .A4(n[1623]), .Z(n147)
         );
  XOR4D0 U90 ( .A1(n[1617]), .A2(n[1616]), .A3(n149), .A4(n150), .Z(n148) );
  XOR3D0 U91 ( .A1(n151), .A2(n152), .A3(n[1615]), .Z(n150) );
  XOR4D0 U92 ( .A1(n[1608]), .A2(n153), .A3(n[1610]), .A4(n[1609]), .Z(n152)
         );
  XOR4D0 U93 ( .A1(n[1603]), .A2(n[1602]), .A3(n154), .A4(n155), .Z(n153) );
  XOR3D0 U94 ( .A1(n156), .A2(n157), .A3(n[1601]), .Z(n155) );
  XOR4D0 U95 ( .A1(n[1594]), .A2(n158), .A3(n[1596]), .A4(n[1595]), .Z(n157)
         );
  XOR4D0 U96 ( .A1(n[1589]), .A2(n[1588]), .A3(n159), .A4(n160), .Z(n158) );
  XOR3D0 U97 ( .A1(n161), .A2(n162), .A3(n[1587]), .Z(n160) );
  XOR4D0 U98 ( .A1(n[1580]), .A2(n163), .A3(n[1582]), .A4(n[1581]), .Z(n162)
         );
  XOR4D0 U99 ( .A1(n[1575]), .A2(n[1574]), .A3(n164), .A4(n165), .Z(n163) );
  XOR3D0 U100 ( .A1(n166), .A2(n167), .A3(n[1573]), .Z(n165) );
  XOR4D0 U101 ( .A1(n[1566]), .A2(n168), .A3(n[1568]), .A4(n[1567]), .Z(n167)
         );
  XOR4D0 U102 ( .A1(n[1561]), .A2(n[1560]), .A3(n169), .A4(n170), .Z(n168) );
  XOR3D0 U103 ( .A1(n171), .A2(n172), .A3(n[1559]), .Z(n170) );
  XOR4D0 U104 ( .A1(n[1552]), .A2(n173), .A3(n[1554]), .A4(n[1553]), .Z(n172)
         );
  XOR4D0 U105 ( .A1(n[1547]), .A2(n[1546]), .A3(n174), .A4(n175), .Z(n173) );
  XOR3D0 U106 ( .A1(n176), .A2(n177), .A3(n[1545]), .Z(n175) );
  XOR4D0 U107 ( .A1(n[1538]), .A2(n178), .A3(n[1540]), .A4(n[1539]), .Z(n177)
         );
  XOR4D0 U108 ( .A1(n[1533]), .A2(n[1532]), .A3(n179), .A4(n180), .Z(n178) );
  XOR3D0 U109 ( .A1(n181), .A2(n182), .A3(n[1531]), .Z(n180) );
  XOR4D0 U110 ( .A1(n[1524]), .A2(n183), .A3(n[1526]), .A4(n[1525]), .Z(n182)
         );
  XOR4D0 U111 ( .A1(n[1519]), .A2(n[1518]), .A3(n184), .A4(n185), .Z(n183) );
  XOR3D0 U112 ( .A1(n186), .A2(n187), .A3(n[1517]), .Z(n185) );
  XOR4D0 U113 ( .A1(n[1510]), .A2(n188), .A3(n[1512]), .A4(n[1511]), .Z(n187)
         );
  XOR4D0 U114 ( .A1(n[1505]), .A2(n[1504]), .A3(n189), .A4(n190), .Z(n188) );
  XOR3D0 U115 ( .A1(n191), .A2(n192), .A3(n[1503]), .Z(n190) );
  XOR4D0 U116 ( .A1(n[1496]), .A2(n193), .A3(n[1498]), .A4(n[1497]), .Z(n192)
         );
  XOR4D0 U117 ( .A1(n[1491]), .A2(n[1490]), .A3(n194), .A4(n195), .Z(n193) );
  XOR3D0 U118 ( .A1(n196), .A2(n197), .A3(n[1489]), .Z(n195) );
  XOR4D0 U119 ( .A1(n[1482]), .A2(n198), .A3(n[1484]), .A4(n[1483]), .Z(n197)
         );
  XOR4D0 U120 ( .A1(n[1477]), .A2(n[1476]), .A3(n199), .A4(n200), .Z(n198) );
  XOR3D0 U121 ( .A1(n201), .A2(n202), .A3(n[1475]), .Z(n200) );
  XOR4D0 U122 ( .A1(n[1468]), .A2(n203), .A3(n[1470]), .A4(n[1469]), .Z(n202)
         );
  XOR4D0 U123 ( .A1(n[1463]), .A2(n[1462]), .A3(n204), .A4(n205), .Z(n203) );
  XOR3D0 U124 ( .A1(n206), .A2(n207), .A3(n[1461]), .Z(n205) );
  XOR4D0 U125 ( .A1(n[1454]), .A2(n208), .A3(n[1456]), .A4(n[1455]), .Z(n207)
         );
  XOR4D0 U126 ( .A1(n[1449]), .A2(n[1448]), .A3(n209), .A4(n210), .Z(n208) );
  XOR3D0 U127 ( .A1(n211), .A2(n212), .A3(n[1447]), .Z(n210) );
  XOR4D0 U128 ( .A1(n[1440]), .A2(n213), .A3(n[1442]), .A4(n[1441]), .Z(n212)
         );
  XOR4D0 U129 ( .A1(n[1435]), .A2(n[1434]), .A3(n214), .A4(n215), .Z(n213) );
  XOR3D0 U130 ( .A1(n216), .A2(n217), .A3(n[1433]), .Z(n215) );
  XOR4D0 U131 ( .A1(n[1426]), .A2(n218), .A3(n[1428]), .A4(n[1427]), .Z(n217)
         );
  XOR4D0 U132 ( .A1(n[1421]), .A2(n[1420]), .A3(n219), .A4(n220), .Z(n218) );
  XOR3D0 U133 ( .A1(n221), .A2(n222), .A3(n[1419]), .Z(n220) );
  XOR4D0 U134 ( .A1(n[1412]), .A2(n223), .A3(n[1414]), .A4(n[1413]), .Z(n222)
         );
  XOR4D0 U135 ( .A1(n[1407]), .A2(n[1406]), .A3(n224), .A4(n225), .Z(n223) );
  XOR3D0 U136 ( .A1(n226), .A2(n227), .A3(n[1405]), .Z(n225) );
  XOR4D0 U137 ( .A1(n[1398]), .A2(n228), .A3(n[1400]), .A4(n[1399]), .Z(n227)
         );
  XOR4D0 U138 ( .A1(n[1393]), .A2(n[1392]), .A3(n229), .A4(n230), .Z(n228) );
  XOR3D0 U139 ( .A1(n231), .A2(n232), .A3(n[1391]), .Z(n230) );
  XOR4D0 U140 ( .A1(n[1384]), .A2(n233), .A3(n[1386]), .A4(n[1385]), .Z(n232)
         );
  XOR4D0 U141 ( .A1(n[1379]), .A2(n[1378]), .A3(n234), .A4(n235), .Z(n233) );
  XOR3D0 U142 ( .A1(n236), .A2(n237), .A3(n[1377]), .Z(n235) );
  XOR4D0 U143 ( .A1(n[1370]), .A2(n238), .A3(n[1372]), .A4(n[1371]), .Z(n237)
         );
  XOR4D0 U144 ( .A1(n[1365]), .A2(n[1364]), .A3(n239), .A4(n240), .Z(n238) );
  XOR3D0 U145 ( .A1(n241), .A2(n242), .A3(n[1363]), .Z(n240) );
  XOR4D0 U146 ( .A1(n[1356]), .A2(n243), .A3(n[1358]), .A4(n[1357]), .Z(n242)
         );
  XOR4D0 U147 ( .A1(n[1351]), .A2(n[1350]), .A3(n244), .A4(n245), .Z(n243) );
  XOR3D0 U148 ( .A1(n246), .A2(n247), .A3(n[1349]), .Z(n245) );
  XOR4D0 U149 ( .A1(n[1342]), .A2(n248), .A3(n[1344]), .A4(n[1343]), .Z(n247)
         );
  XOR4D0 U150 ( .A1(n[1337]), .A2(n[1336]), .A3(n249), .A4(n250), .Z(n248) );
  XOR3D0 U151 ( .A1(n251), .A2(n252), .A3(n[1335]), .Z(n250) );
  XOR4D0 U152 ( .A1(n[1328]), .A2(n253), .A3(n[1330]), .A4(n[1329]), .Z(n252)
         );
  XOR4D0 U153 ( .A1(n[1323]), .A2(n[1322]), .A3(n254), .A4(n255), .Z(n253) );
  XOR3D0 U154 ( .A1(n256), .A2(n257), .A3(n[1321]), .Z(n255) );
  XOR4D0 U155 ( .A1(n[1314]), .A2(n258), .A3(n[1316]), .A4(n[1315]), .Z(n257)
         );
  XOR4D0 U156 ( .A1(n[1309]), .A2(n[1308]), .A3(n259), .A4(n260), .Z(n258) );
  XOR3D0 U157 ( .A1(n261), .A2(n262), .A3(n[1307]), .Z(n260) );
  XOR4D0 U158 ( .A1(n[1300]), .A2(n263), .A3(n[1302]), .A4(n[1301]), .Z(n262)
         );
  XOR4D0 U159 ( .A1(n[1295]), .A2(n[1294]), .A3(n264), .A4(n265), .Z(n263) );
  XOR3D0 U160 ( .A1(n266), .A2(n267), .A3(n[1293]), .Z(n265) );
  XOR4D0 U161 ( .A1(n[1286]), .A2(n268), .A3(n[1288]), .A4(n[1287]), .Z(n267)
         );
  XOR4D0 U162 ( .A1(n[1281]), .A2(n[1280]), .A3(n269), .A4(n270), .Z(n268) );
  XOR3D0 U163 ( .A1(n271), .A2(n272), .A3(n[1279]), .Z(n270) );
  XOR4D0 U164 ( .A1(n[1272]), .A2(n273), .A3(n[1274]), .A4(n[1273]), .Z(n272)
         );
  XOR4D0 U165 ( .A1(n[1267]), .A2(n[1266]), .A3(n274), .A4(n275), .Z(n273) );
  XOR3D0 U166 ( .A1(n276), .A2(n277), .A3(n[1265]), .Z(n275) );
  XOR4D0 U167 ( .A1(n[1258]), .A2(n278), .A3(n[1260]), .A4(n[1259]), .Z(n277)
         );
  XOR4D0 U168 ( .A1(n[1253]), .A2(n[1252]), .A3(n279), .A4(n280), .Z(n278) );
  XOR3D0 U169 ( .A1(n281), .A2(n282), .A3(n[1251]), .Z(n280) );
  XOR4D0 U170 ( .A1(n[1244]), .A2(n283), .A3(n[1246]), .A4(n[1245]), .Z(n282)
         );
  XOR4D0 U171 ( .A1(n[1239]), .A2(n[1238]), .A3(n284), .A4(n285), .Z(n283) );
  XOR3D0 U172 ( .A1(n286), .A2(n287), .A3(n[1237]), .Z(n285) );
  XOR4D0 U173 ( .A1(n[1230]), .A2(n288), .A3(n[1232]), .A4(n[1231]), .Z(n287)
         );
  XOR4D0 U174 ( .A1(n[1225]), .A2(n[1224]), .A3(n289), .A4(n290), .Z(n288) );
  XOR3D0 U175 ( .A1(n291), .A2(n292), .A3(n[1223]), .Z(n290) );
  XOR4D0 U176 ( .A1(n[1216]), .A2(n293), .A3(n[1218]), .A4(n[1217]), .Z(n292)
         );
  XOR4D0 U177 ( .A1(n[1211]), .A2(n[1210]), .A3(n294), .A4(n295), .Z(n293) );
  XOR3D0 U178 ( .A1(n296), .A2(n297), .A3(n[1209]), .Z(n295) );
  XOR4D0 U179 ( .A1(n[1202]), .A2(n298), .A3(n[1204]), .A4(n[1203]), .Z(n297)
         );
  XOR4D0 U180 ( .A1(n[1197]), .A2(n[1196]), .A3(n299), .A4(n300), .Z(n298) );
  XOR3D0 U181 ( .A1(n301), .A2(n302), .A3(n[1195]), .Z(n300) );
  XOR4D0 U182 ( .A1(n[1188]), .A2(n303), .A3(n[1190]), .A4(n[1189]), .Z(n302)
         );
  XOR4D0 U183 ( .A1(n[1183]), .A2(n[1182]), .A3(n304), .A4(n305), .Z(n303) );
  XOR3D0 U184 ( .A1(n306), .A2(n307), .A3(n[1181]), .Z(n305) );
  XOR4D0 U185 ( .A1(n[1174]), .A2(n308), .A3(n[1176]), .A4(n[1175]), .Z(n307)
         );
  XOR4D0 U186 ( .A1(n[1169]), .A2(n[1168]), .A3(n309), .A4(n310), .Z(n308) );
  XOR3D0 U187 ( .A1(n311), .A2(n312), .A3(n[1167]), .Z(n310) );
  XOR4D0 U188 ( .A1(n[1160]), .A2(n313), .A3(n[1162]), .A4(n[1161]), .Z(n312)
         );
  XOR4D0 U189 ( .A1(n[1155]), .A2(n[1154]), .A3(n314), .A4(n315), .Z(n313) );
  XOR3D0 U190 ( .A1(n316), .A2(n317), .A3(n[1153]), .Z(n315) );
  XOR4D0 U191 ( .A1(n[1146]), .A2(n318), .A3(n[1148]), .A4(n[1147]), .Z(n317)
         );
  XOR4D0 U192 ( .A1(n[1141]), .A2(n[1140]), .A3(n319), .A4(n320), .Z(n318) );
  XOR3D0 U193 ( .A1(n321), .A2(n322), .A3(n[1139]), .Z(n320) );
  XOR4D0 U194 ( .A1(n[1132]), .A2(n323), .A3(n[1134]), .A4(n[1133]), .Z(n322)
         );
  XOR4D0 U195 ( .A1(n[1127]), .A2(n[1126]), .A3(n324), .A4(n325), .Z(n323) );
  XOR3D0 U196 ( .A1(n326), .A2(n327), .A3(n[1125]), .Z(n325) );
  XOR4D0 U197 ( .A1(n[1118]), .A2(n328), .A3(n[1120]), .A4(n[1119]), .Z(n327)
         );
  XOR4D0 U198 ( .A1(n[1113]), .A2(n[1112]), .A3(n329), .A4(n330), .Z(n328) );
  XOR3D0 U199 ( .A1(n331), .A2(n332), .A3(n[1111]), .Z(n330) );
  XOR4D0 U200 ( .A1(n[1104]), .A2(n333), .A3(n[1106]), .A4(n[1105]), .Z(n332)
         );
  XOR4D0 U201 ( .A1(n[1099]), .A2(n[1098]), .A3(n334), .A4(n335), .Z(n333) );
  XOR3D0 U202 ( .A1(n336), .A2(n337), .A3(n[1097]), .Z(n335) );
  XOR4D0 U203 ( .A1(n[1090]), .A2(n338), .A3(n[1092]), .A4(n[1091]), .Z(n337)
         );
  XOR4D0 U204 ( .A1(n[1085]), .A2(n[1084]), .A3(n339), .A4(n340), .Z(n338) );
  XOR3D0 U205 ( .A1(n341), .A2(n342), .A3(n[1083]), .Z(n340) );
  XOR4D0 U206 ( .A1(n[1076]), .A2(n343), .A3(n[1078]), .A4(n[1077]), .Z(n342)
         );
  XOR4D0 U207 ( .A1(n[1071]), .A2(n[1070]), .A3(n344), .A4(n345), .Z(n343) );
  XOR3D0 U208 ( .A1(n346), .A2(n347), .A3(n[1069]), .Z(n345) );
  XOR4D0 U209 ( .A1(n[1062]), .A2(n348), .A3(n[1064]), .A4(n[1063]), .Z(n347)
         );
  XOR4D0 U210 ( .A1(n[1057]), .A2(n[1056]), .A3(n349), .A4(n350), .Z(n348) );
  XOR3D0 U211 ( .A1(n351), .A2(n352), .A3(n[1055]), .Z(n350) );
  XOR4D0 U212 ( .A1(n[1048]), .A2(n353), .A3(n[1050]), .A4(n[1049]), .Z(n352)
         );
  XOR4D0 U213 ( .A1(n[1043]), .A2(n[1042]), .A3(n354), .A4(n355), .Z(n353) );
  XOR3D0 U214 ( .A1(n356), .A2(n357), .A3(n[1041]), .Z(n355) );
  XOR4D0 U215 ( .A1(n[1034]), .A2(n358), .A3(n[1036]), .A4(n[1035]), .Z(n357)
         );
  XOR4D0 U216 ( .A1(n[1029]), .A2(n[1028]), .A3(n359), .A4(n360), .Z(n358) );
  XOR3D0 U217 ( .A1(n361), .A2(n362), .A3(n[1027]), .Z(n360) );
  XOR3D0 U218 ( .A1(n[1022]), .A2(n[1021]), .A3(n363), .Z(n362) );
  XOR3D0 U219 ( .A1(n364), .A2(n365), .A3(n[1020]), .Z(n363) );
  XOR4D0 U220 ( .A1(n[1013]), .A2(n[1012]), .A3(n[1015]), .A4(n[1014]), .Z(
        n365) );
  XOR4D0 U221 ( .A1(n[1017]), .A2(n[1016]), .A3(n[1019]), .A4(n[1018]), .Z(
        n364) );
  XOR4D0 U222 ( .A1(n[1024]), .A2(n[1023]), .A3(n[1026]), .A4(n[1025]), .Z(
        n361) );
  XOR4D0 U223 ( .A1(n[1031]), .A2(n[1030]), .A3(n[1033]), .A4(n[1032]), .Z(
        n359) );
  XOR4D0 U224 ( .A1(n[1038]), .A2(n[1037]), .A3(n[1040]), .A4(n[1039]), .Z(
        n356) );
  XOR4D0 U225 ( .A1(n[1045]), .A2(n[1044]), .A3(n[1047]), .A4(n[1046]), .Z(
        n354) );
  XOR4D0 U226 ( .A1(n[1052]), .A2(n[1051]), .A3(n[1054]), .A4(n[1053]), .Z(
        n351) );
  XOR4D0 U227 ( .A1(n[1059]), .A2(n[1058]), .A3(n[1061]), .A4(n[1060]), .Z(
        n349) );
  XOR4D0 U228 ( .A1(n[1066]), .A2(n[1065]), .A3(n[1068]), .A4(n[1067]), .Z(
        n346) );
  XOR4D0 U229 ( .A1(n[1073]), .A2(n[1072]), .A3(n[1075]), .A4(n[1074]), .Z(
        n344) );
  XOR4D0 U230 ( .A1(n[1080]), .A2(n[1079]), .A3(n[1082]), .A4(n[1081]), .Z(
        n341) );
  XOR4D0 U231 ( .A1(n[1087]), .A2(n[1086]), .A3(n[1089]), .A4(n[1088]), .Z(
        n339) );
  XOR4D0 U232 ( .A1(n[1094]), .A2(n[1093]), .A3(n[1096]), .A4(n[1095]), .Z(
        n336) );
  XOR4D0 U233 ( .A1(n[1101]), .A2(n[1100]), .A3(n[1103]), .A4(n[1102]), .Z(
        n334) );
  XOR4D0 U234 ( .A1(n[1108]), .A2(n[1107]), .A3(n[1110]), .A4(n[1109]), .Z(
        n331) );
  XOR4D0 U235 ( .A1(n[1115]), .A2(n[1114]), .A3(n[1117]), .A4(n[1116]), .Z(
        n329) );
  XOR4D0 U236 ( .A1(n[1122]), .A2(n[1121]), .A3(n[1124]), .A4(n[1123]), .Z(
        n326) );
  XOR4D0 U237 ( .A1(n[1129]), .A2(n[1128]), .A3(n[1131]), .A4(n[1130]), .Z(
        n324) );
  XOR4D0 U238 ( .A1(n[1136]), .A2(n[1135]), .A3(n[1138]), .A4(n[1137]), .Z(
        n321) );
  XOR4D0 U239 ( .A1(n[1143]), .A2(n[1142]), .A3(n[1145]), .A4(n[1144]), .Z(
        n319) );
  XOR4D0 U240 ( .A1(n[1150]), .A2(n[1149]), .A3(n[1152]), .A4(n[1151]), .Z(
        n316) );
  XOR4D0 U241 ( .A1(n[1157]), .A2(n[1156]), .A3(n[1159]), .A4(n[1158]), .Z(
        n314) );
  XOR4D0 U242 ( .A1(n[1164]), .A2(n[1163]), .A3(n[1166]), .A4(n[1165]), .Z(
        n311) );
  XOR4D0 U243 ( .A1(n[1171]), .A2(n[1170]), .A3(n[1173]), .A4(n[1172]), .Z(
        n309) );
  XOR4D0 U244 ( .A1(n[1178]), .A2(n[1177]), .A3(n[1180]), .A4(n[1179]), .Z(
        n306) );
  XOR4D0 U245 ( .A1(n[1185]), .A2(n[1184]), .A3(n[1187]), .A4(n[1186]), .Z(
        n304) );
  XOR4D0 U246 ( .A1(n[1192]), .A2(n[1191]), .A3(n[1194]), .A4(n[1193]), .Z(
        n301) );
  XOR4D0 U247 ( .A1(n[1199]), .A2(n[1198]), .A3(n[1201]), .A4(n[1200]), .Z(
        n299) );
  XOR4D0 U248 ( .A1(n[1206]), .A2(n[1205]), .A3(n[1208]), .A4(n[1207]), .Z(
        n296) );
  XOR4D0 U249 ( .A1(n[1213]), .A2(n[1212]), .A3(n[1215]), .A4(n[1214]), .Z(
        n294) );
  XOR4D0 U250 ( .A1(n[1220]), .A2(n[1219]), .A3(n[1222]), .A4(n[1221]), .Z(
        n291) );
  XOR4D0 U251 ( .A1(n[1227]), .A2(n[1226]), .A3(n[1229]), .A4(n[1228]), .Z(
        n289) );
  XOR4D0 U252 ( .A1(n[1234]), .A2(n[1233]), .A3(n[1236]), .A4(n[1235]), .Z(
        n286) );
  XOR4D0 U253 ( .A1(n[1241]), .A2(n[1240]), .A3(n[1243]), .A4(n[1242]), .Z(
        n284) );
  XOR4D0 U254 ( .A1(n[1248]), .A2(n[1247]), .A3(n[1250]), .A4(n[1249]), .Z(
        n281) );
  XOR4D0 U255 ( .A1(n[1255]), .A2(n[1254]), .A3(n[1257]), .A4(n[1256]), .Z(
        n279) );
  XOR4D0 U256 ( .A1(n[1262]), .A2(n[1261]), .A3(n[1264]), .A4(n[1263]), .Z(
        n276) );
  XOR4D0 U257 ( .A1(n[1269]), .A2(n[1268]), .A3(n[1271]), .A4(n[1270]), .Z(
        n274) );
  XOR4D0 U258 ( .A1(n[1276]), .A2(n[1275]), .A3(n[1278]), .A4(n[1277]), .Z(
        n271) );
  XOR4D0 U259 ( .A1(n[1283]), .A2(n[1282]), .A3(n[1285]), .A4(n[1284]), .Z(
        n269) );
  XOR4D0 U260 ( .A1(n[1290]), .A2(n[1289]), .A3(n[1292]), .A4(n[1291]), .Z(
        n266) );
  XOR4D0 U261 ( .A1(n[1297]), .A2(n[1296]), .A3(n[1299]), .A4(n[1298]), .Z(
        n264) );
  XOR4D0 U262 ( .A1(n[1304]), .A2(n[1303]), .A3(n[1306]), .A4(n[1305]), .Z(
        n261) );
  XOR4D0 U263 ( .A1(n[1311]), .A2(n[1310]), .A3(n[1313]), .A4(n[1312]), .Z(
        n259) );
  XOR4D0 U264 ( .A1(n[1318]), .A2(n[1317]), .A3(n[1320]), .A4(n[1319]), .Z(
        n256) );
  XOR4D0 U265 ( .A1(n[1325]), .A2(n[1324]), .A3(n[1327]), .A4(n[1326]), .Z(
        n254) );
  XOR4D0 U266 ( .A1(n[1332]), .A2(n[1331]), .A3(n[1334]), .A4(n[1333]), .Z(
        n251) );
  XOR4D0 U267 ( .A1(n[1339]), .A2(n[1338]), .A3(n[1341]), .A4(n[1340]), .Z(
        n249) );
  XOR4D0 U268 ( .A1(n[1346]), .A2(n[1345]), .A3(n[1348]), .A4(n[1347]), .Z(
        n246) );
  XOR4D0 U269 ( .A1(n[1353]), .A2(n[1352]), .A3(n[1355]), .A4(n[1354]), .Z(
        n244) );
  XOR4D0 U270 ( .A1(n[1360]), .A2(n[1359]), .A3(n[1362]), .A4(n[1361]), .Z(
        n241) );
  XOR4D0 U271 ( .A1(n[1367]), .A2(n[1366]), .A3(n[1369]), .A4(n[1368]), .Z(
        n239) );
  XOR4D0 U272 ( .A1(n[1374]), .A2(n[1373]), .A3(n[1376]), .A4(n[1375]), .Z(
        n236) );
  XOR4D0 U273 ( .A1(n[1381]), .A2(n[1380]), .A3(n[1383]), .A4(n[1382]), .Z(
        n234) );
  XOR4D0 U274 ( .A1(n[1388]), .A2(n[1387]), .A3(n[1390]), .A4(n[1389]), .Z(
        n231) );
  XOR4D0 U275 ( .A1(n[1395]), .A2(n[1394]), .A3(n[1397]), .A4(n[1396]), .Z(
        n229) );
  XOR4D0 U276 ( .A1(n[1402]), .A2(n[1401]), .A3(n[1404]), .A4(n[1403]), .Z(
        n226) );
  XOR4D0 U277 ( .A1(n[1409]), .A2(n[1408]), .A3(n[1411]), .A4(n[1410]), .Z(
        n224) );
  XOR4D0 U278 ( .A1(n[1416]), .A2(n[1415]), .A3(n[1418]), .A4(n[1417]), .Z(
        n221) );
  XOR4D0 U279 ( .A1(n[1423]), .A2(n[1422]), .A3(n[1425]), .A4(n[1424]), .Z(
        n219) );
  XOR4D0 U280 ( .A1(n[1430]), .A2(n[1429]), .A3(n[1432]), .A4(n[1431]), .Z(
        n216) );
  XOR4D0 U281 ( .A1(n[1437]), .A2(n[1436]), .A3(n[1439]), .A4(n[1438]), .Z(
        n214) );
  XOR4D0 U282 ( .A1(n[1444]), .A2(n[1443]), .A3(n[1446]), .A4(n[1445]), .Z(
        n211) );
  XOR4D0 U283 ( .A1(n[1451]), .A2(n[1450]), .A3(n[1453]), .A4(n[1452]), .Z(
        n209) );
  XOR4D0 U284 ( .A1(n[1458]), .A2(n[1457]), .A3(n[1460]), .A4(n[1459]), .Z(
        n206) );
  XOR4D0 U285 ( .A1(n[1465]), .A2(n[1464]), .A3(n[1467]), .A4(n[1466]), .Z(
        n204) );
  XOR4D0 U286 ( .A1(n[1472]), .A2(n[1471]), .A3(n[1474]), .A4(n[1473]), .Z(
        n201) );
  XOR4D0 U287 ( .A1(n[1479]), .A2(n[1478]), .A3(n[1481]), .A4(n[1480]), .Z(
        n199) );
  XOR4D0 U288 ( .A1(n[1486]), .A2(n[1485]), .A3(n[1488]), .A4(n[1487]), .Z(
        n196) );
  XOR4D0 U289 ( .A1(n[1493]), .A2(n[1492]), .A3(n[1495]), .A4(n[1494]), .Z(
        n194) );
  XOR4D0 U290 ( .A1(n[1500]), .A2(n[1499]), .A3(n[1502]), .A4(n[1501]), .Z(
        n191) );
  XOR4D0 U291 ( .A1(n[1507]), .A2(n[1506]), .A3(n[1509]), .A4(n[1508]), .Z(
        n189) );
  XOR4D0 U292 ( .A1(n[1514]), .A2(n[1513]), .A3(n[1516]), .A4(n[1515]), .Z(
        n186) );
  XOR4D0 U293 ( .A1(n[1521]), .A2(n[1520]), .A3(n[1523]), .A4(n[1522]), .Z(
        n184) );
  XOR4D0 U294 ( .A1(n[1528]), .A2(n[1527]), .A3(n[1530]), .A4(n[1529]), .Z(
        n181) );
  XOR4D0 U295 ( .A1(n[1535]), .A2(n[1534]), .A3(n[1537]), .A4(n[1536]), .Z(
        n179) );
  XOR4D0 U296 ( .A1(n[1542]), .A2(n[1541]), .A3(n[1544]), .A4(n[1543]), .Z(
        n176) );
  XOR4D0 U297 ( .A1(n[1549]), .A2(n[1548]), .A3(n[1551]), .A4(n[1550]), .Z(
        n174) );
  XOR4D0 U298 ( .A1(n[1556]), .A2(n[1555]), .A3(n[1558]), .A4(n[1557]), .Z(
        n171) );
  XOR4D0 U299 ( .A1(n[1563]), .A2(n[1562]), .A3(n[1565]), .A4(n[1564]), .Z(
        n169) );
  XOR4D0 U300 ( .A1(n[1570]), .A2(n[1569]), .A3(n[1572]), .A4(n[1571]), .Z(
        n166) );
  XOR4D0 U301 ( .A1(n[1577]), .A2(n[1576]), .A3(n[1579]), .A4(n[1578]), .Z(
        n164) );
  XOR4D0 U302 ( .A1(n[1584]), .A2(n[1583]), .A3(n[1586]), .A4(n[1585]), .Z(
        n161) );
  XOR4D0 U303 ( .A1(n[1591]), .A2(n[1590]), .A3(n[1593]), .A4(n[1592]), .Z(
        n159) );
  XOR4D0 U304 ( .A1(n[1598]), .A2(n[1597]), .A3(n[1600]), .A4(n[1599]), .Z(
        n156) );
  XOR4D0 U305 ( .A1(n[1605]), .A2(n[1604]), .A3(n[1607]), .A4(n[1606]), .Z(
        n154) );
  XOR4D0 U306 ( .A1(n[1612]), .A2(n[1611]), .A3(n[1614]), .A4(n[1613]), .Z(
        n151) );
  XOR4D0 U307 ( .A1(n[1619]), .A2(n[1618]), .A3(n[1621]), .A4(n[1620]), .Z(
        n149) );
  XOR4D0 U308 ( .A1(n[1626]), .A2(n[1625]), .A3(n[1628]), .A4(n[1627]), .Z(
        n146) );
  XOR4D0 U309 ( .A1(n[1633]), .A2(n[1632]), .A3(n[1635]), .A4(n[1634]), .Z(
        n144) );
  XOR4D0 U310 ( .A1(n[1640]), .A2(n[1639]), .A3(n[1642]), .A4(n[1641]), .Z(
        n141) );
  XOR4D0 U311 ( .A1(n[1647]), .A2(n[1646]), .A3(n[1649]), .A4(n[1648]), .Z(
        n139) );
  XOR4D0 U312 ( .A1(n[1654]), .A2(n[1653]), .A3(n[1656]), .A4(n[1655]), .Z(
        n136) );
  XOR4D0 U313 ( .A1(n[1661]), .A2(n[1660]), .A3(n[1663]), .A4(n[1662]), .Z(
        n134) );
  XOR4D0 U314 ( .A1(n[1668]), .A2(n[1667]), .A3(n[1670]), .A4(n[1669]), .Z(
        n131) );
  XOR4D0 U315 ( .A1(n[1675]), .A2(n[1674]), .A3(n[1677]), .A4(n[1676]), .Z(
        n129) );
  XOR4D0 U316 ( .A1(n[1682]), .A2(n[1681]), .A3(n[1684]), .A4(n[1683]), .Z(
        n126) );
  XOR4D0 U317 ( .A1(n[1689]), .A2(n[1688]), .A3(n[1691]), .A4(n[1690]), .Z(
        n124) );
  XOR4D0 U318 ( .A1(n[1696]), .A2(n[1695]), .A3(n[1698]), .A4(n[1697]), .Z(
        n121) );
  XOR4D0 U319 ( .A1(n[1703]), .A2(n[1702]), .A3(n[1705]), .A4(n[1704]), .Z(
        n119) );
  XOR4D0 U320 ( .A1(n[1710]), .A2(n[1709]), .A3(n[1712]), .A4(n[1711]), .Z(
        n116) );
  XOR4D0 U321 ( .A1(n[1717]), .A2(n[1716]), .A3(n[1719]), .A4(n[1718]), .Z(
        n114) );
  XOR4D0 U322 ( .A1(n[1724]), .A2(n[1723]), .A3(n[1726]), .A4(n[1725]), .Z(
        n111) );
  XOR4D0 U323 ( .A1(n[1731]), .A2(n[1730]), .A3(n[1733]), .A4(n[1732]), .Z(
        n109) );
  XOR4D0 U324 ( .A1(n[1738]), .A2(n[1737]), .A3(n[1740]), .A4(n[1739]), .Z(
        n106) );
  XOR4D0 U325 ( .A1(n[1745]), .A2(n[1744]), .A3(n[1747]), .A4(n[1746]), .Z(
        n104) );
  XOR4D0 U326 ( .A1(n[1752]), .A2(n[1751]), .A3(n[1754]), .A4(n[1753]), .Z(
        n101) );
  XOR4D0 U327 ( .A1(n[1759]), .A2(n[1758]), .A3(n[1761]), .A4(n[1760]), .Z(n99) );
  XOR4D0 U328 ( .A1(n[1766]), .A2(n[1765]), .A3(n[1768]), .A4(n[1767]), .Z(n96) );
  XOR4D0 U329 ( .A1(n[1773]), .A2(n[1772]), .A3(n[1775]), .A4(n[1774]), .Z(n94) );
  XOR4D0 U330 ( .A1(n[1780]), .A2(n[1779]), .A3(n[1782]), .A4(n[1781]), .Z(n91) );
  XOR4D0 U331 ( .A1(n[1787]), .A2(n[1786]), .A3(n[1789]), .A4(n[1788]), .Z(n89) );
  XOR4D0 U332 ( .A1(n[1794]), .A2(n[1793]), .A3(n[1796]), .A4(n[1795]), .Z(n86) );
  XOR4D0 U333 ( .A1(n[1801]), .A2(n[1800]), .A3(n[1803]), .A4(n[1802]), .Z(n84) );
  XOR4D0 U334 ( .A1(n[1808]), .A2(n[1807]), .A3(n[1810]), .A4(n[1809]), .Z(n81) );
  XOR4D0 U335 ( .A1(n[1815]), .A2(n[1814]), .A3(n[1817]), .A4(n[1816]), .Z(n79) );
  XOR4D0 U336 ( .A1(n[1822]), .A2(n[1821]), .A3(n[1824]), .A4(n[1823]), .Z(n76) );
  XOR4D0 U337 ( .A1(n[1829]), .A2(n[1828]), .A3(n[1831]), .A4(n[1830]), .Z(n74) );
  XOR4D0 U338 ( .A1(n[1836]), .A2(n[1835]), .A3(n[1838]), .A4(n[1837]), .Z(n71) );
  XOR4D0 U339 ( .A1(n[1843]), .A2(n[1842]), .A3(n[1845]), .A4(n[1844]), .Z(n69) );
  XOR4D0 U340 ( .A1(n[1850]), .A2(n[1849]), .A3(n[1852]), .A4(n[1851]), .Z(n66) );
  XOR4D0 U341 ( .A1(n[1857]), .A2(n[1856]), .A3(n[1859]), .A4(n[1858]), .Z(n64) );
  XOR4D0 U342 ( .A1(n[1864]), .A2(n[1863]), .A3(n[1866]), .A4(n[1865]), .Z(n61) );
  XOR4D0 U343 ( .A1(n[1871]), .A2(n[1870]), .A3(n[1873]), .A4(n[1872]), .Z(n59) );
  XOR4D0 U344 ( .A1(n[1878]), .A2(n[1877]), .A3(n[1880]), .A4(n[1879]), .Z(n56) );
  XOR4D0 U345 ( .A1(n[1885]), .A2(n[1884]), .A3(n[1887]), .A4(n[1886]), .Z(n54) );
  XOR4D0 U346 ( .A1(n[1892]), .A2(n[1891]), .A3(n[1894]), .A4(n[1893]), .Z(n51) );
  XOR4D0 U347 ( .A1(n[1899]), .A2(n[1898]), .A3(n[1901]), .A4(n[1900]), .Z(n49) );
  XOR4D0 U348 ( .A1(n[1906]), .A2(n[1905]), .A3(n[1908]), .A4(n[1907]), .Z(n46) );
  XOR4D0 U349 ( .A1(n[1913]), .A2(n[1912]), .A3(n[1915]), .A4(n[1914]), .Z(n44) );
  XOR4D0 U350 ( .A1(n[1920]), .A2(n[1919]), .A3(n[1922]), .A4(n[1921]), .Z(n41) );
  XOR4D0 U351 ( .A1(n[1927]), .A2(n[1926]), .A3(n[1929]), .A4(n[1928]), .Z(n39) );
  XOR4D0 U352 ( .A1(n[1934]), .A2(n[1933]), .A3(n[1936]), .A4(n[1935]), .Z(n36) );
  XOR4D0 U353 ( .A1(n[1941]), .A2(n[1940]), .A3(n[1943]), .A4(n[1942]), .Z(n34) );
  XOR4D0 U354 ( .A1(n[1948]), .A2(n[1947]), .A3(n[1950]), .A4(n[1949]), .Z(n31) );
  XOR4D0 U355 ( .A1(n[1955]), .A2(n[1954]), .A3(n[1957]), .A4(n[1956]), .Z(n29) );
  XOR4D0 U356 ( .A1(n[1962]), .A2(n[1961]), .A3(n[1964]), .A4(n[1963]), .Z(n26) );
  XOR4D0 U357 ( .A1(n[1969]), .A2(n[1968]), .A3(n[1971]), .A4(n[1970]), .Z(n24) );
  XOR4D0 U358 ( .A1(n[1976]), .A2(n[1975]), .A3(n[1978]), .A4(n[1977]), .Z(n21) );
  XOR4D0 U359 ( .A1(n[1983]), .A2(n[1982]), .A3(n[1985]), .A4(n[1984]), .Z(n19) );
  XOR4D0 U360 ( .A1(n[1990]), .A2(n[1989]), .A3(n[1992]), .A4(n[1991]), .Z(n16) );
  XOR4D0 U361 ( .A1(n[1997]), .A2(n[1996]), .A3(n[1999]), .A4(n[1998]), .Z(n14) );
  XOR4D0 U362 ( .A1(n[2004]), .A2(n[2003]), .A3(n[2006]), .A4(n[2005]), .Z(n11) );
  XOR4D0 U363 ( .A1(n[2011]), .A2(n[2010]), .A3(n[2013]), .A4(n[2012]), .Z(n9)
         );
  XOR4D0 U364 ( .A1(n[2018]), .A2(n[2017]), .A3(n[2020]), .A4(n[2019]), .Z(n6)
         );
  XOR4D0 U365 ( .A1(n[2025]), .A2(n[2024]), .A3(n[2027]), .A4(n[2026]), .Z(n4)
         );
  XOR4D0 U366 ( .A1(n[2032]), .A2(n[2031]), .A3(n[2034]), .A4(n[2033]), .Z(n1)
         );
  XOR3D0 U367 ( .A1(n366), .A2(n367), .A3(n[1011]), .Z(s[8]) );
  XOR4D0 U368 ( .A1(a[8]), .A2(n368), .A3(n[1006]), .A4(b[8]), .Z(n367) );
  XOR4D0 U369 ( .A1(n[1002]), .A2(n[1001]), .A3(n369), .A4(n370), .Z(n368) );
  XOR3D0 U370 ( .A1(n371), .A2(n372), .A3(n[1000]), .Z(n370) );
  XOR4D0 U371 ( .A1(n[992]), .A2(n373), .A3(n[994]), .A4(n[993]), .Z(n372) );
  XOR4D0 U372 ( .A1(n[987]), .A2(n[986]), .A3(n374), .A4(n375), .Z(n373) );
  XOR3D0 U373 ( .A1(n376), .A2(n377), .A3(n[985]), .Z(n375) );
  XOR4D0 U374 ( .A1(n[978]), .A2(n378), .A3(n[980]), .A4(n[979]), .Z(n377) );
  XOR4D0 U375 ( .A1(n[973]), .A2(n[972]), .A3(n379), .A4(n380), .Z(n378) );
  XOR3D0 U376 ( .A1(n381), .A2(n382), .A3(n[971]), .Z(n380) );
  XOR4D0 U377 ( .A1(n[964]), .A2(n383), .A3(n[966]), .A4(n[965]), .Z(n382) );
  XOR4D0 U378 ( .A1(n[959]), .A2(n[958]), .A3(n384), .A4(n385), .Z(n383) );
  XOR3D0 U379 ( .A1(n386), .A2(n387), .A3(n[957]), .Z(n385) );
  XOR4D0 U380 ( .A1(n[950]), .A2(n388), .A3(n[952]), .A4(n[951]), .Z(n387) );
  XOR4D0 U381 ( .A1(n[945]), .A2(n[944]), .A3(n389), .A4(n390), .Z(n388) );
  XOR3D0 U382 ( .A1(n391), .A2(n392), .A3(n[943]), .Z(n390) );
  XOR4D0 U383 ( .A1(n[936]), .A2(n393), .A3(n[938]), .A4(n[937]), .Z(n392) );
  XOR4D0 U384 ( .A1(n[931]), .A2(n[930]), .A3(n394), .A4(n395), .Z(n393) );
  XOR3D0 U385 ( .A1(n396), .A2(n397), .A3(n[929]), .Z(n395) );
  XOR4D0 U386 ( .A1(n[922]), .A2(n398), .A3(n[924]), .A4(n[923]), .Z(n397) );
  XOR4D0 U387 ( .A1(n[917]), .A2(n[916]), .A3(n399), .A4(n400), .Z(n398) );
  XOR3D0 U388 ( .A1(n401), .A2(n402), .A3(n[915]), .Z(n400) );
  XOR4D0 U389 ( .A1(n[908]), .A2(n403), .A3(n[910]), .A4(n[909]), .Z(n402) );
  XOR4D0 U390 ( .A1(n[903]), .A2(n[902]), .A3(n404), .A4(n405), .Z(n403) );
  XOR3D0 U391 ( .A1(n406), .A2(n407), .A3(n[901]), .Z(n405) );
  XOR4D0 U392 ( .A1(n[894]), .A2(n408), .A3(n[896]), .A4(n[895]), .Z(n407) );
  XOR4D0 U393 ( .A1(n[889]), .A2(n[888]), .A3(n409), .A4(n410), .Z(n408) );
  XOR3D0 U394 ( .A1(n411), .A2(n412), .A3(n[887]), .Z(n410) );
  XOR4D0 U395 ( .A1(n[880]), .A2(n413), .A3(n[882]), .A4(n[881]), .Z(n412) );
  XOR4D0 U396 ( .A1(n[875]), .A2(n[874]), .A3(n414), .A4(n415), .Z(n413) );
  XOR3D0 U397 ( .A1(n416), .A2(n417), .A3(n[873]), .Z(n415) );
  XOR4D0 U398 ( .A1(n[866]), .A2(n418), .A3(n[868]), .A4(n[867]), .Z(n417) );
  XOR4D0 U399 ( .A1(n[861]), .A2(n[860]), .A3(n419), .A4(n420), .Z(n418) );
  XOR3D0 U400 ( .A1(n421), .A2(n422), .A3(n[859]), .Z(n420) );
  XOR4D0 U401 ( .A1(n[852]), .A2(n423), .A3(n[854]), .A4(n[853]), .Z(n422) );
  XOR4D0 U402 ( .A1(n[847]), .A2(n[846]), .A3(n424), .A4(n425), .Z(n423) );
  XOR3D0 U403 ( .A1(n426), .A2(n427), .A3(n[845]), .Z(n425) );
  XOR4D0 U404 ( .A1(n[838]), .A2(n428), .A3(n[840]), .A4(n[839]), .Z(n427) );
  XOR4D0 U405 ( .A1(n[833]), .A2(n[832]), .A3(n429), .A4(n430), .Z(n428) );
  XOR3D0 U406 ( .A1(n431), .A2(n432), .A3(n[831]), .Z(n430) );
  XOR4D0 U407 ( .A1(n[824]), .A2(n433), .A3(n[826]), .A4(n[825]), .Z(n432) );
  XOR4D0 U408 ( .A1(n[819]), .A2(n[818]), .A3(n434), .A4(n435), .Z(n433) );
  XOR3D0 U409 ( .A1(n436), .A2(n437), .A3(n[817]), .Z(n435) );
  XOR4D0 U410 ( .A1(n[810]), .A2(n438), .A3(n[812]), .A4(n[811]), .Z(n437) );
  XOR4D0 U411 ( .A1(n[805]), .A2(n[804]), .A3(n439), .A4(n440), .Z(n438) );
  XOR3D0 U412 ( .A1(n441), .A2(n442), .A3(n[803]), .Z(n440) );
  XOR4D0 U413 ( .A1(n[796]), .A2(n443), .A3(n[798]), .A4(n[797]), .Z(n442) );
  XOR4D0 U414 ( .A1(n[791]), .A2(n[790]), .A3(n444), .A4(n445), .Z(n443) );
  XOR3D0 U415 ( .A1(n446), .A2(n447), .A3(n[789]), .Z(n445) );
  XOR4D0 U416 ( .A1(n[782]), .A2(n448), .A3(n[784]), .A4(n[783]), .Z(n447) );
  XOR4D0 U417 ( .A1(n[777]), .A2(n[776]), .A3(n449), .A4(n450), .Z(n448) );
  XOR3D0 U418 ( .A1(n451), .A2(n452), .A3(n[775]), .Z(n450) );
  XOR4D0 U419 ( .A1(n[768]), .A2(n453), .A3(n[770]), .A4(n[769]), .Z(n452) );
  XOR4D0 U420 ( .A1(n[763]), .A2(n[762]), .A3(n454), .A4(n455), .Z(n453) );
  XOR3D0 U421 ( .A1(n456), .A2(n457), .A3(n[761]), .Z(n455) );
  XOR4D0 U422 ( .A1(n[754]), .A2(n458), .A3(n[756]), .A4(n[755]), .Z(n457) );
  XOR4D0 U423 ( .A1(n[749]), .A2(n[748]), .A3(n459), .A4(n460), .Z(n458) );
  XOR3D0 U424 ( .A1(n461), .A2(n462), .A3(n[747]), .Z(n460) );
  XOR4D0 U425 ( .A1(n[740]), .A2(n463), .A3(n[742]), .A4(n[741]), .Z(n462) );
  XOR4D0 U426 ( .A1(n[735]), .A2(n[734]), .A3(n464), .A4(n465), .Z(n463) );
  XOR3D0 U427 ( .A1(n466), .A2(n467), .A3(n[733]), .Z(n465) );
  XOR4D0 U428 ( .A1(n[726]), .A2(n468), .A3(n[728]), .A4(n[727]), .Z(n467) );
  XOR4D0 U429 ( .A1(n[721]), .A2(n[720]), .A3(n469), .A4(n470), .Z(n468) );
  XOR3D0 U430 ( .A1(n471), .A2(n472), .A3(n[719]), .Z(n470) );
  XOR4D0 U431 ( .A1(n[712]), .A2(n473), .A3(n[714]), .A4(n[713]), .Z(n472) );
  XOR4D0 U432 ( .A1(n[707]), .A2(n[706]), .A3(n474), .A4(n475), .Z(n473) );
  XOR3D0 U433 ( .A1(n476), .A2(n477), .A3(n[705]), .Z(n475) );
  XOR4D0 U434 ( .A1(n[698]), .A2(n478), .A3(n[700]), .A4(n[699]), .Z(n477) );
  XOR4D0 U435 ( .A1(n[693]), .A2(n[692]), .A3(n479), .A4(n480), .Z(n478) );
  XOR3D0 U436 ( .A1(n481), .A2(n482), .A3(n[691]), .Z(n480) );
  XOR4D0 U437 ( .A1(n[684]), .A2(n483), .A3(n[686]), .A4(n[685]), .Z(n482) );
  XOR4D0 U438 ( .A1(n[679]), .A2(n[678]), .A3(n484), .A4(n485), .Z(n483) );
  XOR3D0 U439 ( .A1(n486), .A2(n487), .A3(n[677]), .Z(n485) );
  XOR4D0 U440 ( .A1(n[670]), .A2(n488), .A3(n[672]), .A4(n[671]), .Z(n487) );
  XOR4D0 U441 ( .A1(n[665]), .A2(n[664]), .A3(n489), .A4(n490), .Z(n488) );
  XOR3D0 U442 ( .A1(n491), .A2(n492), .A3(n[663]), .Z(n490) );
  XOR4D0 U443 ( .A1(n[656]), .A2(n493), .A3(n[658]), .A4(n[657]), .Z(n492) );
  XOR4D0 U444 ( .A1(n[651]), .A2(n[650]), .A3(n494), .A4(n495), .Z(n493) );
  XOR3D0 U445 ( .A1(n496), .A2(n497), .A3(n[649]), .Z(n495) );
  XOR4D0 U446 ( .A1(n[642]), .A2(n498), .A3(n[644]), .A4(n[643]), .Z(n497) );
  XOR4D0 U447 ( .A1(n[637]), .A2(n[636]), .A3(n499), .A4(n500), .Z(n498) );
  XOR3D0 U448 ( .A1(n501), .A2(n502), .A3(n[635]), .Z(n500) );
  XOR4D0 U449 ( .A1(n[628]), .A2(n503), .A3(n[630]), .A4(n[629]), .Z(n502) );
  XOR4D0 U450 ( .A1(n[623]), .A2(n[622]), .A3(n504), .A4(n505), .Z(n503) );
  XOR3D0 U451 ( .A1(n506), .A2(n507), .A3(n[621]), .Z(n505) );
  XOR4D0 U452 ( .A1(n[614]), .A2(n508), .A3(n[616]), .A4(n[615]), .Z(n507) );
  XOR4D0 U453 ( .A1(n[609]), .A2(n[608]), .A3(n509), .A4(n510), .Z(n508) );
  XOR3D0 U454 ( .A1(n511), .A2(n512), .A3(n[607]), .Z(n510) );
  XOR4D0 U455 ( .A1(n[600]), .A2(n513), .A3(n[602]), .A4(n[601]), .Z(n512) );
  XOR4D0 U456 ( .A1(n[595]), .A2(n[594]), .A3(n514), .A4(n515), .Z(n513) );
  XOR3D0 U457 ( .A1(n516), .A2(n517), .A3(n[593]), .Z(n515) );
  XOR4D0 U458 ( .A1(n[586]), .A2(n518), .A3(n[588]), .A4(n[587]), .Z(n517) );
  XOR4D0 U459 ( .A1(n[581]), .A2(n[580]), .A3(n519), .A4(n520), .Z(n518) );
  XOR3D0 U460 ( .A1(n521), .A2(n522), .A3(n[579]), .Z(n520) );
  XOR4D0 U461 ( .A1(n[572]), .A2(n523), .A3(n[574]), .A4(n[573]), .Z(n522) );
  XOR4D0 U462 ( .A1(n[567]), .A2(n[566]), .A3(n524), .A4(n525), .Z(n523) );
  XOR3D0 U463 ( .A1(n526), .A2(n527), .A3(n[565]), .Z(n525) );
  XOR4D0 U464 ( .A1(n[558]), .A2(n528), .A3(n[560]), .A4(n[559]), .Z(n527) );
  XOR4D0 U465 ( .A1(n[553]), .A2(n[552]), .A3(n529), .A4(n530), .Z(n528) );
  XOR3D0 U466 ( .A1(n531), .A2(n532), .A3(n[551]), .Z(n530) );
  XOR4D0 U467 ( .A1(n[544]), .A2(n533), .A3(n[546]), .A4(n[545]), .Z(n532) );
  XOR4D0 U468 ( .A1(n[539]), .A2(n[538]), .A3(n534), .A4(n535), .Z(n533) );
  XOR3D0 U469 ( .A1(n536), .A2(n537), .A3(n[537]), .Z(n535) );
  XOR4D0 U470 ( .A1(n[530]), .A2(n538), .A3(n[532]), .A4(n[531]), .Z(n537) );
  XOR4D0 U471 ( .A1(n[525]), .A2(n[524]), .A3(n539), .A4(n540), .Z(n538) );
  XOR3D0 U472 ( .A1(n541), .A2(n542), .A3(n[523]), .Z(n540) );
  XOR4D0 U473 ( .A1(n[516]), .A2(n543), .A3(n[518]), .A4(n[517]), .Z(n542) );
  XOR4D0 U474 ( .A1(n[511]), .A2(n[510]), .A3(n544), .A4(n545), .Z(n543) );
  XOR3D0 U475 ( .A1(n546), .A2(n547), .A3(n[509]), .Z(n545) );
  XOR4D0 U476 ( .A1(n[502]), .A2(n[501]), .A3(n[504]), .A4(n[503]), .Z(n547)
         );
  XOR4D0 U477 ( .A1(n[506]), .A2(n[505]), .A3(n[508]), .A4(n[507]), .Z(n546)
         );
  XOR4D0 U478 ( .A1(n[513]), .A2(n[512]), .A3(n[515]), .A4(n[514]), .Z(n544)
         );
  XOR4D0 U479 ( .A1(n[520]), .A2(n[519]), .A3(n[522]), .A4(n[521]), .Z(n541)
         );
  XOR4D0 U480 ( .A1(n[527]), .A2(n[526]), .A3(n[529]), .A4(n[528]), .Z(n539)
         );
  XOR4D0 U481 ( .A1(n[534]), .A2(n[533]), .A3(n[536]), .A4(n[535]), .Z(n536)
         );
  XOR4D0 U482 ( .A1(n[541]), .A2(n[540]), .A3(n[543]), .A4(n[542]), .Z(n534)
         );
  XOR4D0 U483 ( .A1(n[548]), .A2(n[547]), .A3(n[550]), .A4(n[549]), .Z(n531)
         );
  XOR4D0 U484 ( .A1(n[555]), .A2(n[554]), .A3(n[557]), .A4(n[556]), .Z(n529)
         );
  XOR4D0 U485 ( .A1(n[562]), .A2(n[561]), .A3(n[564]), .A4(n[563]), .Z(n526)
         );
  XOR4D0 U486 ( .A1(n[569]), .A2(n[568]), .A3(n[571]), .A4(n[570]), .Z(n524)
         );
  XOR4D0 U487 ( .A1(n[576]), .A2(n[575]), .A3(n[578]), .A4(n[577]), .Z(n521)
         );
  XOR4D0 U488 ( .A1(n[583]), .A2(n[582]), .A3(n[585]), .A4(n[584]), .Z(n519)
         );
  XOR4D0 U489 ( .A1(n[590]), .A2(n[589]), .A3(n[592]), .A4(n[591]), .Z(n516)
         );
  XOR4D0 U490 ( .A1(n[597]), .A2(n[596]), .A3(n[599]), .A4(n[598]), .Z(n514)
         );
  XOR4D0 U491 ( .A1(n[604]), .A2(n[603]), .A3(n[606]), .A4(n[605]), .Z(n511)
         );
  XOR4D0 U492 ( .A1(n[611]), .A2(n[610]), .A3(n[613]), .A4(n[612]), .Z(n509)
         );
  XOR4D0 U493 ( .A1(n[618]), .A2(n[617]), .A3(n[620]), .A4(n[619]), .Z(n506)
         );
  XOR4D0 U494 ( .A1(n[625]), .A2(n[624]), .A3(n[627]), .A4(n[626]), .Z(n504)
         );
  XOR4D0 U495 ( .A1(n[632]), .A2(n[631]), .A3(n[634]), .A4(n[633]), .Z(n501)
         );
  XOR4D0 U496 ( .A1(n[639]), .A2(n[638]), .A3(n[641]), .A4(n[640]), .Z(n499)
         );
  XOR4D0 U497 ( .A1(n[646]), .A2(n[645]), .A3(n[648]), .A4(n[647]), .Z(n496)
         );
  XOR4D0 U498 ( .A1(n[653]), .A2(n[652]), .A3(n[655]), .A4(n[654]), .Z(n494)
         );
  XOR4D0 U499 ( .A1(n[660]), .A2(n[659]), .A3(n[662]), .A4(n[661]), .Z(n491)
         );
  XOR4D0 U500 ( .A1(n[667]), .A2(n[666]), .A3(n[669]), .A4(n[668]), .Z(n489)
         );
  XOR4D0 U501 ( .A1(n[674]), .A2(n[673]), .A3(n[676]), .A4(n[675]), .Z(n486)
         );
  XOR4D0 U502 ( .A1(n[681]), .A2(n[680]), .A3(n[683]), .A4(n[682]), .Z(n484)
         );
  XOR4D0 U503 ( .A1(n[688]), .A2(n[687]), .A3(n[690]), .A4(n[689]), .Z(n481)
         );
  XOR4D0 U504 ( .A1(n[695]), .A2(n[694]), .A3(n[697]), .A4(n[696]), .Z(n479)
         );
  XOR4D0 U505 ( .A1(n[702]), .A2(n[701]), .A3(n[704]), .A4(n[703]), .Z(n476)
         );
  XOR4D0 U506 ( .A1(n[709]), .A2(n[708]), .A3(n[711]), .A4(n[710]), .Z(n474)
         );
  XOR4D0 U507 ( .A1(n[716]), .A2(n[715]), .A3(n[718]), .A4(n[717]), .Z(n471)
         );
  XOR4D0 U508 ( .A1(n[723]), .A2(n[722]), .A3(n[725]), .A4(n[724]), .Z(n469)
         );
  XOR4D0 U509 ( .A1(n[730]), .A2(n[729]), .A3(n[732]), .A4(n[731]), .Z(n466)
         );
  XOR4D0 U510 ( .A1(n[737]), .A2(n[736]), .A3(n[739]), .A4(n[738]), .Z(n464)
         );
  XOR4D0 U511 ( .A1(n[744]), .A2(n[743]), .A3(n[746]), .A4(n[745]), .Z(n461)
         );
  XOR4D0 U512 ( .A1(n[751]), .A2(n[750]), .A3(n[753]), .A4(n[752]), .Z(n459)
         );
  XOR4D0 U513 ( .A1(n[758]), .A2(n[757]), .A3(n[760]), .A4(n[759]), .Z(n456)
         );
  XOR4D0 U514 ( .A1(n[765]), .A2(n[764]), .A3(n[767]), .A4(n[766]), .Z(n454)
         );
  XOR4D0 U515 ( .A1(n[772]), .A2(n[771]), .A3(n[774]), .A4(n[773]), .Z(n451)
         );
  XOR4D0 U516 ( .A1(n[779]), .A2(n[778]), .A3(n[781]), .A4(n[780]), .Z(n449)
         );
  XOR4D0 U517 ( .A1(n[786]), .A2(n[785]), .A3(n[788]), .A4(n[787]), .Z(n446)
         );
  XOR4D0 U518 ( .A1(n[793]), .A2(n[792]), .A3(n[795]), .A4(n[794]), .Z(n444)
         );
  XOR4D0 U519 ( .A1(n[800]), .A2(n[799]), .A3(n[802]), .A4(n[801]), .Z(n441)
         );
  XOR4D0 U520 ( .A1(n[807]), .A2(n[806]), .A3(n[809]), .A4(n[808]), .Z(n439)
         );
  XOR4D0 U521 ( .A1(n[814]), .A2(n[813]), .A3(n[816]), .A4(n[815]), .Z(n436)
         );
  XOR4D0 U522 ( .A1(n[821]), .A2(n[820]), .A3(n[823]), .A4(n[822]), .Z(n434)
         );
  XOR4D0 U523 ( .A1(n[828]), .A2(n[827]), .A3(n[830]), .A4(n[829]), .Z(n431)
         );
  XOR4D0 U524 ( .A1(n[835]), .A2(n[834]), .A3(n[837]), .A4(n[836]), .Z(n429)
         );
  XOR4D0 U525 ( .A1(n[842]), .A2(n[841]), .A3(n[844]), .A4(n[843]), .Z(n426)
         );
  XOR4D0 U526 ( .A1(n[849]), .A2(n[848]), .A3(n[851]), .A4(n[850]), .Z(n424)
         );
  XOR4D0 U527 ( .A1(n[856]), .A2(n[855]), .A3(n[858]), .A4(n[857]), .Z(n421)
         );
  XOR4D0 U528 ( .A1(n[863]), .A2(n[862]), .A3(n[865]), .A4(n[864]), .Z(n419)
         );
  XOR4D0 U529 ( .A1(n[870]), .A2(n[869]), .A3(n[872]), .A4(n[871]), .Z(n416)
         );
  XOR4D0 U530 ( .A1(n[877]), .A2(n[876]), .A3(n[879]), .A4(n[878]), .Z(n414)
         );
  XOR4D0 U531 ( .A1(n[884]), .A2(n[883]), .A3(n[886]), .A4(n[885]), .Z(n411)
         );
  XOR4D0 U532 ( .A1(n[891]), .A2(n[890]), .A3(n[893]), .A4(n[892]), .Z(n409)
         );
  XOR4D0 U533 ( .A1(n[898]), .A2(n[897]), .A3(n[900]), .A4(n[899]), .Z(n406)
         );
  XOR4D0 U534 ( .A1(n[905]), .A2(n[904]), .A3(n[907]), .A4(n[906]), .Z(n404)
         );
  XOR4D0 U535 ( .A1(n[912]), .A2(n[911]), .A3(n[914]), .A4(n[913]), .Z(n401)
         );
  XOR4D0 U536 ( .A1(n[919]), .A2(n[918]), .A3(n[921]), .A4(n[920]), .Z(n399)
         );
  XOR4D0 U537 ( .A1(n[926]), .A2(n[925]), .A3(n[928]), .A4(n[927]), .Z(n396)
         );
  XOR4D0 U538 ( .A1(n[933]), .A2(n[932]), .A3(n[935]), .A4(n[934]), .Z(n394)
         );
  XOR4D0 U539 ( .A1(n[940]), .A2(n[939]), .A3(n[942]), .A4(n[941]), .Z(n391)
         );
  XOR4D0 U540 ( .A1(n[947]), .A2(n[946]), .A3(n[949]), .A4(n[948]), .Z(n389)
         );
  XOR4D0 U541 ( .A1(n[954]), .A2(n[953]), .A3(n[956]), .A4(n[955]), .Z(n386)
         );
  XOR4D0 U542 ( .A1(n[961]), .A2(n[960]), .A3(n[963]), .A4(n[962]), .Z(n384)
         );
  XOR4D0 U543 ( .A1(n[968]), .A2(n[967]), .A3(n[970]), .A4(n[969]), .Z(n381)
         );
  XOR4D0 U544 ( .A1(n[975]), .A2(n[974]), .A3(n[977]), .A4(n[976]), .Z(n379)
         );
  XOR4D0 U545 ( .A1(n[982]), .A2(n[981]), .A3(n[984]), .A4(n[983]), .Z(n376)
         );
  XOR4D0 U546 ( .A1(n[989]), .A2(n[988]), .A3(n[991]), .A4(n[990]), .Z(n374)
         );
  XOR4D0 U547 ( .A1(n[996]), .A2(n[995]), .A3(n[998]), .A4(n[997]), .Z(n371)
         );
  XOR4D0 U548 ( .A1(n[1004]), .A2(n[1003]), .A3(n[999]), .A4(n[1005]), .Z(n369) );
  XOR4D0 U549 ( .A1(n[1008]), .A2(n[1007]), .A3(n[1010]), .A4(n[1009]), .Z(
        n366) );
  XOR4D0 U550 ( .A1(n548), .A2(n549), .A3(n550), .A4(n[495]), .Z(s[7]) );
  XOR3D0 U551 ( .A1(n[498]), .A2(n[497]), .A3(n[496]), .Z(n550) );
  XOR4D0 U552 ( .A1(a[7]), .A2(n551), .A3(n[492]), .A4(b[7]), .Z(n549) );
  XOR4D0 U553 ( .A1(n[487]), .A2(n[486]), .A3(n552), .A4(n553), .Z(n551) );
  XOR3D0 U554 ( .A1(n554), .A2(n555), .A3(n[485]), .Z(n553) );
  XOR4D0 U555 ( .A1(n[478]), .A2(n556), .A3(n[480]), .A4(n[479]), .Z(n555) );
  XOR4D0 U556 ( .A1(n[473]), .A2(n[472]), .A3(n557), .A4(n558), .Z(n556) );
  XOR3D0 U557 ( .A1(n559), .A2(n560), .A3(n[471]), .Z(n558) );
  XOR4D0 U558 ( .A1(n[464]), .A2(n561), .A3(n[466]), .A4(n[465]), .Z(n560) );
  XOR4D0 U559 ( .A1(n[459]), .A2(n[458]), .A3(n562), .A4(n563), .Z(n561) );
  XOR3D0 U560 ( .A1(n564), .A2(n565), .A3(n[457]), .Z(n563) );
  XOR4D0 U561 ( .A1(n[450]), .A2(n566), .A3(n[452]), .A4(n[451]), .Z(n565) );
  XOR4D0 U562 ( .A1(n[445]), .A2(n[444]), .A3(n567), .A4(n568), .Z(n566) );
  XOR3D0 U563 ( .A1(n569), .A2(n570), .A3(n[443]), .Z(n568) );
  XOR4D0 U564 ( .A1(n[436]), .A2(n571), .A3(n[438]), .A4(n[437]), .Z(n570) );
  XOR4D0 U565 ( .A1(n[431]), .A2(n[430]), .A3(n572), .A4(n573), .Z(n571) );
  XOR3D0 U566 ( .A1(n574), .A2(n575), .A3(n[429]), .Z(n573) );
  XOR4D0 U567 ( .A1(n[422]), .A2(n576), .A3(n[424]), .A4(n[423]), .Z(n575) );
  XOR4D0 U568 ( .A1(n[417]), .A2(n[416]), .A3(n577), .A4(n578), .Z(n576) );
  XOR3D0 U569 ( .A1(n579), .A2(n580), .A3(n[415]), .Z(n578) );
  XOR4D0 U570 ( .A1(n[408]), .A2(n581), .A3(n[410]), .A4(n[409]), .Z(n580) );
  XOR4D0 U571 ( .A1(n[403]), .A2(n[402]), .A3(n582), .A4(n583), .Z(n581) );
  XOR3D0 U572 ( .A1(n584), .A2(n585), .A3(n[401]), .Z(n583) );
  XOR4D0 U573 ( .A1(n[394]), .A2(n586), .A3(n[396]), .A4(n[395]), .Z(n585) );
  XOR4D0 U574 ( .A1(n[389]), .A2(n[388]), .A3(n587), .A4(n588), .Z(n586) );
  XOR3D0 U575 ( .A1(n589), .A2(n590), .A3(n[387]), .Z(n588) );
  XOR4D0 U576 ( .A1(n[380]), .A2(n591), .A3(n[382]), .A4(n[381]), .Z(n590) );
  XOR4D0 U577 ( .A1(n[375]), .A2(n[374]), .A3(n592), .A4(n593), .Z(n591) );
  XOR3D0 U578 ( .A1(n594), .A2(n595), .A3(n[373]), .Z(n593) );
  XOR4D0 U579 ( .A1(n[366]), .A2(n596), .A3(n[368]), .A4(n[367]), .Z(n595) );
  XOR4D0 U580 ( .A1(n[361]), .A2(n[360]), .A3(n597), .A4(n598), .Z(n596) );
  XOR3D0 U581 ( .A1(n599), .A2(n600), .A3(n[359]), .Z(n598) );
  XOR4D0 U582 ( .A1(n[352]), .A2(n601), .A3(n[354]), .A4(n[353]), .Z(n600) );
  XOR4D0 U583 ( .A1(n[347]), .A2(n[346]), .A3(n602), .A4(n603), .Z(n601) );
  XOR3D0 U584 ( .A1(n604), .A2(n605), .A3(n[345]), .Z(n603) );
  XOR4D0 U585 ( .A1(n[338]), .A2(n606), .A3(n[340]), .A4(n[339]), .Z(n605) );
  XOR4D0 U586 ( .A1(n[333]), .A2(n[332]), .A3(n607), .A4(n608), .Z(n606) );
  XOR3D0 U587 ( .A1(n609), .A2(n610), .A3(n[331]), .Z(n608) );
  XOR4D0 U588 ( .A1(n[324]), .A2(n611), .A3(n[326]), .A4(n[325]), .Z(n610) );
  XOR4D0 U589 ( .A1(n[319]), .A2(n[318]), .A3(n612), .A4(n613), .Z(n611) );
  XOR3D0 U590 ( .A1(n614), .A2(n615), .A3(n[317]), .Z(n613) );
  XOR4D0 U591 ( .A1(n[310]), .A2(n616), .A3(n[312]), .A4(n[311]), .Z(n615) );
  XOR4D0 U592 ( .A1(n[305]), .A2(n[304]), .A3(n617), .A4(n618), .Z(n616) );
  XOR3D0 U593 ( .A1(n619), .A2(n620), .A3(n[303]), .Z(n618) );
  XOR4D0 U594 ( .A1(n[296]), .A2(n621), .A3(n[298]), .A4(n[297]), .Z(n620) );
  XOR4D0 U595 ( .A1(n[291]), .A2(n[290]), .A3(n622), .A4(n623), .Z(n621) );
  XOR3D0 U596 ( .A1(n624), .A2(n625), .A3(n[289]), .Z(n623) );
  XOR4D0 U597 ( .A1(n[282]), .A2(n626), .A3(n[284]), .A4(n[283]), .Z(n625) );
  XOR4D0 U598 ( .A1(n[277]), .A2(n[276]), .A3(n627), .A4(n628), .Z(n626) );
  XOR3D0 U599 ( .A1(n629), .A2(n630), .A3(n[275]), .Z(n628) );
  XOR4D0 U600 ( .A1(n[268]), .A2(n631), .A3(n[270]), .A4(n[269]), .Z(n630) );
  XOR4D0 U601 ( .A1(n[263]), .A2(n[262]), .A3(n632), .A4(n633), .Z(n631) );
  XOR3D0 U602 ( .A1(n634), .A2(n635), .A3(n[261]), .Z(n633) );
  XOR3D0 U603 ( .A1(n[256]), .A2(n[255]), .A3(n636), .Z(n635) );
  XOR3D0 U604 ( .A1(n637), .A2(n638), .A3(n[254]), .Z(n636) );
  XOR4D0 U605 ( .A1(n[247]), .A2(n[246]), .A3(n[249]), .A4(n[248]), .Z(n638)
         );
  XOR4D0 U606 ( .A1(n[251]), .A2(n[250]), .A3(n[253]), .A4(n[252]), .Z(n637)
         );
  XOR4D0 U607 ( .A1(n[258]), .A2(n[257]), .A3(n[260]), .A4(n[259]), .Z(n634)
         );
  XOR4D0 U608 ( .A1(n[265]), .A2(n[264]), .A3(n[267]), .A4(n[266]), .Z(n632)
         );
  XOR4D0 U609 ( .A1(n[272]), .A2(n[271]), .A3(n[274]), .A4(n[273]), .Z(n629)
         );
  XOR4D0 U610 ( .A1(n[279]), .A2(n[278]), .A3(n[281]), .A4(n[280]), .Z(n627)
         );
  XOR4D0 U611 ( .A1(n[286]), .A2(n[285]), .A3(n[288]), .A4(n[287]), .Z(n624)
         );
  XOR4D0 U612 ( .A1(n[293]), .A2(n[292]), .A3(n[295]), .A4(n[294]), .Z(n622)
         );
  XOR4D0 U613 ( .A1(n[300]), .A2(n[299]), .A3(n[302]), .A4(n[301]), .Z(n619)
         );
  XOR4D0 U614 ( .A1(n[307]), .A2(n[306]), .A3(n[309]), .A4(n[308]), .Z(n617)
         );
  XOR4D0 U615 ( .A1(n[314]), .A2(n[313]), .A3(n[316]), .A4(n[315]), .Z(n614)
         );
  XOR4D0 U616 ( .A1(n[321]), .A2(n[320]), .A3(n[323]), .A4(n[322]), .Z(n612)
         );
  XOR4D0 U617 ( .A1(n[328]), .A2(n[327]), .A3(n[330]), .A4(n[329]), .Z(n609)
         );
  XOR4D0 U618 ( .A1(n[335]), .A2(n[334]), .A3(n[337]), .A4(n[336]), .Z(n607)
         );
  XOR4D0 U619 ( .A1(n[342]), .A2(n[341]), .A3(n[344]), .A4(n[343]), .Z(n604)
         );
  XOR4D0 U620 ( .A1(n[349]), .A2(n[348]), .A3(n[351]), .A4(n[350]), .Z(n602)
         );
  XOR4D0 U621 ( .A1(n[356]), .A2(n[355]), .A3(n[358]), .A4(n[357]), .Z(n599)
         );
  XOR4D0 U622 ( .A1(n[363]), .A2(n[362]), .A3(n[365]), .A4(n[364]), .Z(n597)
         );
  XOR4D0 U623 ( .A1(n[370]), .A2(n[369]), .A3(n[372]), .A4(n[371]), .Z(n594)
         );
  XOR4D0 U624 ( .A1(n[377]), .A2(n[376]), .A3(n[379]), .A4(n[378]), .Z(n592)
         );
  XOR4D0 U625 ( .A1(n[384]), .A2(n[383]), .A3(n[386]), .A4(n[385]), .Z(n589)
         );
  XOR4D0 U626 ( .A1(n[391]), .A2(n[390]), .A3(n[393]), .A4(n[392]), .Z(n587)
         );
  XOR4D0 U627 ( .A1(n[398]), .A2(n[397]), .A3(n[400]), .A4(n[399]), .Z(n584)
         );
  XOR4D0 U628 ( .A1(n[405]), .A2(n[404]), .A3(n[407]), .A4(n[406]), .Z(n582)
         );
  XOR4D0 U629 ( .A1(n[412]), .A2(n[411]), .A3(n[414]), .A4(n[413]), .Z(n579)
         );
  XOR4D0 U630 ( .A1(n[419]), .A2(n[418]), .A3(n[421]), .A4(n[420]), .Z(n577)
         );
  XOR4D0 U631 ( .A1(n[426]), .A2(n[425]), .A3(n[428]), .A4(n[427]), .Z(n574)
         );
  XOR4D0 U632 ( .A1(n[433]), .A2(n[432]), .A3(n[435]), .A4(n[434]), .Z(n572)
         );
  XOR4D0 U633 ( .A1(n[440]), .A2(n[439]), .A3(n[442]), .A4(n[441]), .Z(n569)
         );
  XOR4D0 U634 ( .A1(n[447]), .A2(n[446]), .A3(n[449]), .A4(n[448]), .Z(n567)
         );
  XOR4D0 U635 ( .A1(n[454]), .A2(n[453]), .A3(n[456]), .A4(n[455]), .Z(n564)
         );
  XOR4D0 U636 ( .A1(n[461]), .A2(n[460]), .A3(n[463]), .A4(n[462]), .Z(n562)
         );
  XOR4D0 U637 ( .A1(n[468]), .A2(n[467]), .A3(n[470]), .A4(n[469]), .Z(n559)
         );
  XOR4D0 U638 ( .A1(n[475]), .A2(n[474]), .A3(n[477]), .A4(n[476]), .Z(n557)
         );
  XOR4D0 U639 ( .A1(n[482]), .A2(n[481]), .A3(n[484]), .A4(n[483]), .Z(n554)
         );
  XOR4D0 U640 ( .A1(n[489]), .A2(n[488]), .A3(n[491]), .A4(n[490]), .Z(n552)
         );
  XOR4D0 U641 ( .A1(n[494]), .A2(n[493]), .A3(n[500]), .A4(n[499]), .Z(n548)
         );
  XOR4D0 U642 ( .A1(b[6]), .A2(a[6]), .A3(n639), .A4(n640), .Z(s[6]) );
  XOR4D0 U643 ( .A1(n[239]), .A2(n641), .A3(n[241]), .A4(n[240]), .Z(n640) );
  XOR4D0 U644 ( .A1(n[234]), .A2(n[233]), .A3(n642), .A4(n643), .Z(n641) );
  XOR3D0 U645 ( .A1(n644), .A2(n645), .A3(n[232]), .Z(n643) );
  XOR4D0 U646 ( .A1(n[225]), .A2(n646), .A3(n[227]), .A4(n[226]), .Z(n645) );
  XOR4D0 U647 ( .A1(n[220]), .A2(n[219]), .A3(n647), .A4(n648), .Z(n646) );
  XOR3D0 U648 ( .A1(n649), .A2(n650), .A3(n[218]), .Z(n648) );
  XOR4D0 U649 ( .A1(n[211]), .A2(n651), .A3(n[213]), .A4(n[212]), .Z(n650) );
  XOR4D0 U650 ( .A1(n[206]), .A2(n[205]), .A3(n652), .A4(n653), .Z(n651) );
  XOR3D0 U651 ( .A1(n654), .A2(n655), .A3(n[204]), .Z(n653) );
  XOR4D0 U652 ( .A1(n[197]), .A2(n656), .A3(n[199]), .A4(n[198]), .Z(n655) );
  XOR4D0 U653 ( .A1(n[192]), .A2(n[191]), .A3(n657), .A4(n658), .Z(n656) );
  XOR3D0 U654 ( .A1(n659), .A2(n660), .A3(n[190]), .Z(n658) );
  XOR4D0 U655 ( .A1(n[183]), .A2(n661), .A3(n[185]), .A4(n[184]), .Z(n660) );
  XOR4D0 U656 ( .A1(n[178]), .A2(n[177]), .A3(n662), .A4(n663), .Z(n661) );
  XOR3D0 U657 ( .A1(n664), .A2(n665), .A3(n[176]), .Z(n663) );
  XOR4D0 U658 ( .A1(n[169]), .A2(n666), .A3(n[171]), .A4(n[170]), .Z(n665) );
  XOR4D0 U659 ( .A1(n[164]), .A2(n[163]), .A3(n667), .A4(n668), .Z(n666) );
  XOR3D0 U660 ( .A1(n669), .A2(n670), .A3(n[162]), .Z(n668) );
  XOR4D0 U661 ( .A1(n[155]), .A2(n671), .A3(n[157]), .A4(n[156]), .Z(n670) );
  XOR4D0 U662 ( .A1(n[150]), .A2(n[149]), .A3(n672), .A4(n673), .Z(n671) );
  XOR3D0 U663 ( .A1(n674), .A2(n675), .A3(n[148]), .Z(n673) );
  XOR4D0 U664 ( .A1(n[141]), .A2(n676), .A3(n[143]), .A4(n[142]), .Z(n675) );
  XOR4D0 U665 ( .A1(n[136]), .A2(n[135]), .A3(n677), .A4(n678), .Z(n676) );
  XOR3D0 U666 ( .A1(n679), .A2(n680), .A3(n[134]), .Z(n678) );
  XOR3D0 U667 ( .A1(n[129]), .A2(n[128]), .A3(n681), .Z(n680) );
  XOR3D0 U668 ( .A1(n682), .A2(n683), .A3(n[127]), .Z(n681) );
  XOR4D0 U669 ( .A1(n[120]), .A2(n[119]), .A3(n[122]), .A4(n[121]), .Z(n683)
         );
  XOR4D0 U670 ( .A1(n[124]), .A2(n[123]), .A3(n[126]), .A4(n[125]), .Z(n682)
         );
  XOR4D0 U671 ( .A1(n[131]), .A2(n[130]), .A3(n[133]), .A4(n[132]), .Z(n679)
         );
  XOR4D0 U672 ( .A1(n[138]), .A2(n[137]), .A3(n[140]), .A4(n[139]), .Z(n677)
         );
  XOR4D0 U673 ( .A1(n[145]), .A2(n[144]), .A3(n[147]), .A4(n[146]), .Z(n674)
         );
  XOR4D0 U674 ( .A1(n[152]), .A2(n[151]), .A3(n[154]), .A4(n[153]), .Z(n672)
         );
  XOR4D0 U675 ( .A1(n[159]), .A2(n[158]), .A3(n[161]), .A4(n[160]), .Z(n669)
         );
  XOR4D0 U676 ( .A1(n[166]), .A2(n[165]), .A3(n[168]), .A4(n[167]), .Z(n667)
         );
  XOR4D0 U677 ( .A1(n[173]), .A2(n[172]), .A3(n[175]), .A4(n[174]), .Z(n664)
         );
  XOR4D0 U678 ( .A1(n[180]), .A2(n[179]), .A3(n[182]), .A4(n[181]), .Z(n662)
         );
  XOR4D0 U679 ( .A1(n[187]), .A2(n[186]), .A3(n[189]), .A4(n[188]), .Z(n659)
         );
  XOR4D0 U680 ( .A1(n[194]), .A2(n[193]), .A3(n[196]), .A4(n[195]), .Z(n657)
         );
  XOR4D0 U681 ( .A1(n[201]), .A2(n[200]), .A3(n[203]), .A4(n[202]), .Z(n654)
         );
  XOR4D0 U682 ( .A1(n[208]), .A2(n[207]), .A3(n[210]), .A4(n[209]), .Z(n652)
         );
  XOR4D0 U683 ( .A1(n[215]), .A2(n[214]), .A3(n[217]), .A4(n[216]), .Z(n649)
         );
  XOR4D0 U684 ( .A1(n[222]), .A2(n[221]), .A3(n[224]), .A4(n[223]), .Z(n647)
         );
  XOR4D0 U685 ( .A1(n[229]), .A2(n[228]), .A3(n[231]), .A4(n[230]), .Z(n644)
         );
  XOR4D0 U686 ( .A1(n[236]), .A2(n[235]), .A3(n[238]), .A4(n[237]), .Z(n642)
         );
  XOR4D0 U687 ( .A1(n[243]), .A2(n[242]), .A3(n[245]), .A4(n[244]), .Z(n639)
         );
  XOR3D0 U688 ( .A1(n684), .A2(n685), .A3(n[118]), .Z(s[5]) );
  XOR4D0 U689 ( .A1(a[5]), .A2(n686), .A3(n[113]), .A4(b[5]), .Z(n685) );
  XOR4D0 U690 ( .A1(n[108]), .A2(n[107]), .A3(n687), .A4(n688), .Z(n686) );
  XOR3D0 U691 ( .A1(n689), .A2(n690), .A3(n[106]), .Z(n688) );
  XOR4D0 U692 ( .A1(n[100]), .A2(n691), .A3(n[102]), .A4(n[101]), .Z(n690) );
  XOR4D0 U693 ( .A1(n[94]), .A2(n[93]), .A3(n692), .A4(n693), .Z(n691) );
  XOR3D0 U694 ( .A1(n694), .A2(n695), .A3(n[92]), .Z(n693) );
  XOR4D0 U695 ( .A1(n[85]), .A2(n696), .A3(n[87]), .A4(n[86]), .Z(n695) );
  XOR4D0 U696 ( .A1(n[80]), .A2(n[79]), .A3(n697), .A4(n698), .Z(n696) );
  XOR3D0 U697 ( .A1(n699), .A2(n700), .A3(n[78]), .Z(n698) );
  XOR4D0 U698 ( .A1(n[71]), .A2(n701), .A3(n[73]), .A4(n[72]), .Z(n700) );
  XOR4D0 U699 ( .A1(n[66]), .A2(n[65]), .A3(n702), .A4(n703), .Z(n701) );
  XOR3D0 U700 ( .A1(n704), .A2(n705), .A3(n[64]), .Z(n703) );
  XOR4D0 U701 ( .A1(n[57]), .A2(n[56]), .A3(n[59]), .A4(n[58]), .Z(n705) );
  XOR4D0 U702 ( .A1(n[61]), .A2(n[60]), .A3(n[63]), .A4(n[62]), .Z(n704) );
  XOR4D0 U703 ( .A1(n[68]), .A2(n[67]), .A3(n[70]), .A4(n[69]), .Z(n702) );
  XOR4D0 U704 ( .A1(n[75]), .A2(n[74]), .A3(n[77]), .A4(n[76]), .Z(n699) );
  XOR4D0 U705 ( .A1(n[82]), .A2(n[81]), .A3(n[84]), .A4(n[83]), .Z(n697) );
  XOR4D0 U706 ( .A1(n[89]), .A2(n[88]), .A3(n[91]), .A4(n[90]), .Z(n694) );
  XOR4D0 U707 ( .A1(n[96]), .A2(n[95]), .A3(n[98]), .A4(n[97]), .Z(n692) );
  XOR4D0 U708 ( .A1(n[104]), .A2(n[103]), .A3(n[99]), .A4(n[105]), .Z(n689) );
  XOR4D0 U709 ( .A1(n[110]), .A2(n[109]), .A3(n[112]), .A4(n[111]), .Z(n687)
         );
  XOR4D0 U710 ( .A1(n[115]), .A2(n[114]), .A3(n[117]), .A4(n[116]), .Z(n684)
         );
  XOR4D0 U711 ( .A1(n706), .A2(n707), .A3(n708), .A4(n[50]), .Z(s[4]) );
  XOR3D0 U712 ( .A1(n[53]), .A2(n[52]), .A3(n[51]), .Z(n708) );
  XOR4D0 U713 ( .A1(a[4]), .A2(n709), .A3(n[47]), .A4(b[4]), .Z(n707) );
  XOR4D0 U714 ( .A1(n[42]), .A2(n[41]), .A3(n710), .A4(n711), .Z(n709) );
  XOR3D0 U715 ( .A1(n712), .A2(n713), .A3(n[40]), .Z(n711) );
  XOR3D0 U716 ( .A1(n[35]), .A2(n[34]), .A3(n714), .Z(n713) );
  XOR3D0 U717 ( .A1(n715), .A2(n716), .A3(n[33]), .Z(n714) );
  XOR4D0 U718 ( .A1(n[26]), .A2(n[25]), .A3(n[28]), .A4(n[27]), .Z(n716) );
  XOR4D0 U719 ( .A1(n[30]), .A2(n[29]), .A3(n[32]), .A4(n[31]), .Z(n715) );
  XOR4D0 U720 ( .A1(n[37]), .A2(n[36]), .A3(n[39]), .A4(n[38]), .Z(n712) );
  XOR4D0 U721 ( .A1(n[44]), .A2(n[43]), .A3(n[46]), .A4(n[45]), .Z(n710) );
  XOR4D0 U722 ( .A1(n[49]), .A2(n[48]), .A3(n[55]), .A4(n[54]), .Z(n706) );
  XOR4D0 U723 ( .A1(b[3]), .A2(a[3]), .A3(n717), .A4(n718), .Z(s[3]) );
  XOR3D0 U724 ( .A1(n[20]), .A2(n[19]), .A3(n719), .Z(n718) );
  XOR3D0 U725 ( .A1(n720), .A2(n721), .A3(n[18]), .Z(n719) );
  XOR4D0 U726 ( .A1(n[11]), .A2(n[10]), .A3(n[13]), .A4(n[12]), .Z(n721) );
  XOR4D0 U727 ( .A1(n[15]), .A2(n[14]), .A3(n[17]), .A4(n[16]), .Z(n720) );
  XOR4D0 U728 ( .A1(n[22]), .A2(n[21]), .A3(n[24]), .A4(n[23]), .Z(n717) );
  XOR3D0 U729 ( .A1(n722), .A2(n723), .A3(n[9]), .Z(s[2]) );
  XOR4D0 U730 ( .A1(b[2]), .A2(a[2]), .A3(n[4]), .A4(n[3]), .Z(n723) );
  XOR4D0 U731 ( .A1(n[6]), .A2(n[5]), .A3(n[8]), .A4(n[7]), .Z(n722) );
  XOR3D0 U732 ( .A1(b[1]), .A2(a[1]), .A3(n724), .Z(s[1]) );
  XOR3D0 U733 ( .A1(n[2]), .A2(n[1]), .A3(n[0]), .Z(n724) );
  XOR2D0 U734 ( .A1(b[0]), .A2(a[0]), .Z(s[0]) );
endmodule


module gen_nonlinear_part ( a, b, n );
  input [9:0] a;
  input [9:0] b;
  output [2034:0] n;


  INVD0 U2 ( .I(1'b1), .ZN(n[1]) );
  INVD0 U4 ( .I(1'b1), .ZN(n[2]) );
  INVD0 U6 ( .I(1'b1), .ZN(n[5]) );
  INVD0 U8 ( .I(1'b1), .ZN(n[6]) );
  INVD0 U10 ( .I(1'b1), .ZN(n[8]) );
  INVD0 U12 ( .I(1'b1), .ZN(n[9]) );
  INVD0 U14 ( .I(1'b1), .ZN(n[13]) );
  INVD0 U16 ( .I(1'b1), .ZN(n[14]) );
  INVD0 U18 ( .I(1'b1), .ZN(n[16]) );
  INVD0 U20 ( .I(1'b1), .ZN(n[17]) );
  INVD0 U22 ( .I(1'b1), .ZN(n[20]) );
  INVD0 U24 ( .I(1'b1), .ZN(n[21]) );
  INVD0 U26 ( .I(1'b1), .ZN(n[23]) );
  INVD0 U28 ( .I(1'b1), .ZN(n[24]) );
  INVD0 U30 ( .I(1'b1), .ZN(n[29]) );
  INVD0 U32 ( .I(1'b1), .ZN(n[30]) );
  INVD0 U34 ( .I(1'b1), .ZN(n[32]) );
  INVD0 U36 ( .I(1'b1), .ZN(n[33]) );
  INVD0 U38 ( .I(1'b1), .ZN(n[36]) );
  INVD0 U40 ( .I(1'b1), .ZN(n[37]) );
  INVD0 U42 ( .I(1'b1), .ZN(n[39]) );
  INVD0 U44 ( .I(1'b1), .ZN(n[40]) );
  INVD0 U46 ( .I(1'b1), .ZN(n[44]) );
  INVD0 U48 ( .I(1'b1), .ZN(n[45]) );
  INVD0 U50 ( .I(1'b1), .ZN(n[47]) );
  INVD0 U52 ( .I(1'b1), .ZN(n[48]) );
  INVD0 U54 ( .I(1'b1), .ZN(n[51]) );
  INVD0 U56 ( .I(1'b1), .ZN(n[52]) );
  INVD0 U58 ( .I(1'b1), .ZN(n[54]) );
  INVD0 U60 ( .I(1'b1), .ZN(n[55]) );
  INVD0 U62 ( .I(1'b1), .ZN(n[61]) );
  INVD0 U64 ( .I(1'b1), .ZN(n[62]) );
  INVD0 U66 ( .I(1'b1), .ZN(n[64]) );
  INVD0 U68 ( .I(1'b1), .ZN(n[65]) );
  INVD0 U70 ( .I(1'b1), .ZN(n[68]) );
  INVD0 U72 ( .I(1'b1), .ZN(n[69]) );
  INVD0 U74 ( .I(1'b1), .ZN(n[71]) );
  INVD0 U76 ( .I(1'b1), .ZN(n[72]) );
  INVD0 U78 ( .I(1'b1), .ZN(n[76]) );
  INVD0 U80 ( .I(1'b1), .ZN(n[77]) );
  INVD0 U82 ( .I(1'b1), .ZN(n[79]) );
  INVD0 U84 ( .I(1'b1), .ZN(n[80]) );
  INVD0 U86 ( .I(1'b1), .ZN(n[83]) );
  INVD0 U88 ( .I(1'b1), .ZN(n[84]) );
  INVD0 U90 ( .I(1'b1), .ZN(n[86]) );
  INVD0 U92 ( .I(1'b1), .ZN(n[87]) );
  INVD0 U94 ( .I(1'b1), .ZN(n[92]) );
  INVD0 U96 ( .I(1'b1), .ZN(n[93]) );
  INVD0 U98 ( .I(1'b1), .ZN(n[95]) );
  INVD0 U100 ( .I(1'b1), .ZN(n[96]) );
  INVD0 U102 ( .I(1'b1), .ZN(n[99]) );
  INVD0 U104 ( .I(1'b1), .ZN(n[100]) );
  INVD0 U106 ( .I(1'b1), .ZN(n[102]) );
  INVD0 U108 ( .I(1'b1), .ZN(n[103]) );
  INVD0 U110 ( .I(1'b1), .ZN(n[107]) );
  INVD0 U112 ( .I(1'b1), .ZN(n[108]) );
  INVD0 U114 ( .I(1'b1), .ZN(n[110]) );
  INVD0 U116 ( .I(1'b1), .ZN(n[111]) );
  INVD0 U118 ( .I(1'b1), .ZN(n[114]) );
  INVD0 U120 ( .I(1'b1), .ZN(n[115]) );
  INVD0 U122 ( .I(1'b1), .ZN(n[117]) );
  INVD0 U124 ( .I(1'b1), .ZN(n[118]) );
  INVD0 U126 ( .I(1'b1), .ZN(n[125]) );
  INVD0 U128 ( .I(1'b1), .ZN(n[126]) );
  INVD0 U130 ( .I(1'b1), .ZN(n[128]) );
  INVD0 U132 ( .I(1'b1), .ZN(n[129]) );
  INVD0 U134 ( .I(1'b1), .ZN(n[132]) );
  INVD0 U136 ( .I(1'b1), .ZN(n[133]) );
  INVD0 U138 ( .I(1'b1), .ZN(n[135]) );
  INVD0 U140 ( .I(1'b1), .ZN(n[136]) );
  INVD0 U142 ( .I(1'b1), .ZN(n[140]) );
  INVD0 U144 ( .I(1'b1), .ZN(n[141]) );
  INVD0 U146 ( .I(1'b1), .ZN(n[143]) );
  INVD0 U148 ( .I(1'b1), .ZN(n[144]) );
  INVD0 U150 ( .I(1'b1), .ZN(n[147]) );
  INVD0 U152 ( .I(1'b1), .ZN(n[148]) );
  INVD0 U154 ( .I(1'b1), .ZN(n[150]) );
  INVD0 U156 ( .I(1'b1), .ZN(n[151]) );
  INVD0 U158 ( .I(1'b1), .ZN(n[156]) );
  INVD0 U160 ( .I(1'b1), .ZN(n[157]) );
  INVD0 U162 ( .I(1'b1), .ZN(n[159]) );
  INVD0 U164 ( .I(1'b1), .ZN(n[160]) );
  INVD0 U166 ( .I(1'b1), .ZN(n[163]) );
  INVD0 U168 ( .I(1'b1), .ZN(n[164]) );
  INVD0 U170 ( .I(1'b1), .ZN(n[166]) );
  INVD0 U172 ( .I(1'b1), .ZN(n[167]) );
  INVD0 U174 ( .I(1'b1), .ZN(n[171]) );
  INVD0 U176 ( .I(1'b1), .ZN(n[172]) );
  INVD0 U178 ( .I(1'b1), .ZN(n[174]) );
  INVD0 U180 ( .I(1'b1), .ZN(n[175]) );
  INVD0 U182 ( .I(1'b1), .ZN(n[178]) );
  INVD0 U184 ( .I(1'b1), .ZN(n[179]) );
  INVD0 U186 ( .I(1'b1), .ZN(n[181]) );
  INVD0 U188 ( .I(1'b1), .ZN(n[182]) );
  INVD0 U190 ( .I(1'b1), .ZN(n[188]) );
  INVD0 U192 ( .I(1'b1), .ZN(n[189]) );
  INVD0 U194 ( .I(1'b1), .ZN(n[191]) );
  INVD0 U196 ( .I(1'b1), .ZN(n[192]) );
  INVD0 U198 ( .I(1'b1), .ZN(n[195]) );
  INVD0 U200 ( .I(1'b1), .ZN(n[196]) );
  INVD0 U202 ( .I(1'b1), .ZN(n[198]) );
  INVD0 U204 ( .I(1'b1), .ZN(n[199]) );
  INVD0 U206 ( .I(1'b1), .ZN(n[203]) );
  INVD0 U208 ( .I(1'b1), .ZN(n[204]) );
  INVD0 U210 ( .I(1'b1), .ZN(n[206]) );
  INVD0 U212 ( .I(1'b1), .ZN(n[207]) );
  INVD0 U214 ( .I(1'b1), .ZN(n[210]) );
  INVD0 U216 ( .I(1'b1), .ZN(n[211]) );
  INVD0 U218 ( .I(1'b1), .ZN(n[213]) );
  INVD0 U220 ( .I(1'b1), .ZN(n[214]) );
  INVD0 U222 ( .I(1'b1), .ZN(n[219]) );
  INVD0 U224 ( .I(1'b1), .ZN(n[220]) );
  INVD0 U226 ( .I(1'b1), .ZN(n[222]) );
  INVD0 U228 ( .I(1'b1), .ZN(n[223]) );
  INVD0 U230 ( .I(1'b1), .ZN(n[226]) );
  INVD0 U232 ( .I(1'b1), .ZN(n[227]) );
  INVD0 U234 ( .I(1'b1), .ZN(n[229]) );
  INVD0 U236 ( .I(1'b1), .ZN(n[230]) );
  INVD0 U238 ( .I(1'b1), .ZN(n[234]) );
  INVD0 U240 ( .I(1'b1), .ZN(n[235]) );
  INVD0 U242 ( .I(1'b1), .ZN(n[237]) );
  INVD0 U244 ( .I(1'b1), .ZN(n[238]) );
  INVD0 U246 ( .I(1'b1), .ZN(n[241]) );
  INVD0 U248 ( .I(1'b1), .ZN(n[242]) );
  INVD0 U250 ( .I(1'b1), .ZN(n[244]) );
  INVD0 U252 ( .I(1'b1), .ZN(n[245]) );
  INVD0 U254 ( .I(1'b1), .ZN(n[253]) );
  INVD0 U256 ( .I(1'b1), .ZN(n[254]) );
  INVD0 U258 ( .I(1'b1), .ZN(n[256]) );
  INVD0 U260 ( .I(1'b1), .ZN(n[257]) );
  INVD0 U262 ( .I(1'b1), .ZN(n[260]) );
  INVD0 U264 ( .I(1'b1), .ZN(n[261]) );
  INVD0 U266 ( .I(1'b1), .ZN(n[263]) );
  INVD0 U268 ( .I(1'b1), .ZN(n[264]) );
  INVD0 U270 ( .I(1'b1), .ZN(n[268]) );
  INVD0 U272 ( .I(1'b1), .ZN(n[269]) );
  INVD0 U274 ( .I(1'b1), .ZN(n[271]) );
  INVD0 U276 ( .I(1'b1), .ZN(n[272]) );
  INVD0 U278 ( .I(1'b1), .ZN(n[275]) );
  INVD0 U280 ( .I(1'b1), .ZN(n[276]) );
  INVD0 U282 ( .I(1'b1), .ZN(n[278]) );
  INVD0 U284 ( .I(1'b1), .ZN(n[279]) );
  INVD0 U286 ( .I(1'b1), .ZN(n[284]) );
  INVD0 U288 ( .I(1'b1), .ZN(n[285]) );
  INVD0 U290 ( .I(1'b1), .ZN(n[287]) );
  INVD0 U292 ( .I(1'b1), .ZN(n[288]) );
  INVD0 U294 ( .I(1'b1), .ZN(n[291]) );
  INVD0 U296 ( .I(1'b1), .ZN(n[292]) );
  INVD0 U298 ( .I(1'b1), .ZN(n[294]) );
  INVD0 U300 ( .I(1'b1), .ZN(n[295]) );
  INVD0 U302 ( .I(1'b1), .ZN(n[299]) );
  INVD0 U304 ( .I(1'b1), .ZN(n[300]) );
  INVD0 U306 ( .I(1'b1), .ZN(n[302]) );
  INVD0 U308 ( .I(1'b1), .ZN(n[303]) );
  INVD0 U310 ( .I(1'b1), .ZN(n[306]) );
  INVD0 U312 ( .I(1'b1), .ZN(n[307]) );
  INVD0 U314 ( .I(1'b1), .ZN(n[309]) );
  INVD0 U316 ( .I(1'b1), .ZN(n[310]) );
  INVD0 U318 ( .I(1'b1), .ZN(n[316]) );
  INVD0 U320 ( .I(1'b1), .ZN(n[317]) );
  INVD0 U322 ( .I(1'b1), .ZN(n[319]) );
  INVD0 U324 ( .I(1'b1), .ZN(n[320]) );
  INVD0 U326 ( .I(1'b1), .ZN(n[323]) );
  INVD0 U328 ( .I(1'b1), .ZN(n[324]) );
  INVD0 U330 ( .I(1'b1), .ZN(n[326]) );
  INVD0 U332 ( .I(1'b1), .ZN(n[327]) );
  INVD0 U334 ( .I(1'b1), .ZN(n[331]) );
  INVD0 U336 ( .I(1'b1), .ZN(n[332]) );
  INVD0 U338 ( .I(1'b1), .ZN(n[334]) );
  INVD0 U340 ( .I(1'b1), .ZN(n[335]) );
  INVD0 U342 ( .I(1'b1), .ZN(n[338]) );
  INVD0 U344 ( .I(1'b1), .ZN(n[339]) );
  INVD0 U346 ( .I(1'b1), .ZN(n[341]) );
  INVD0 U348 ( .I(1'b1), .ZN(n[342]) );
  INVD0 U350 ( .I(1'b1), .ZN(n[347]) );
  INVD0 U352 ( .I(1'b1), .ZN(n[348]) );
  INVD0 U354 ( .I(1'b1), .ZN(n[350]) );
  INVD0 U356 ( .I(1'b1), .ZN(n[351]) );
  INVD0 U358 ( .I(1'b1), .ZN(n[354]) );
  INVD0 U360 ( .I(1'b1), .ZN(n[355]) );
  INVD0 U362 ( .I(1'b1), .ZN(n[357]) );
  INVD0 U364 ( .I(1'b1), .ZN(n[358]) );
  INVD0 U366 ( .I(1'b1), .ZN(n[362]) );
  INVD0 U368 ( .I(1'b1), .ZN(n[363]) );
  INVD0 U370 ( .I(1'b1), .ZN(n[365]) );
  INVD0 U372 ( .I(1'b1), .ZN(n[366]) );
  INVD0 U374 ( .I(1'b1), .ZN(n[369]) );
  INVD0 U376 ( .I(1'b1), .ZN(n[370]) );
  INVD0 U378 ( .I(1'b1), .ZN(n[372]) );
  INVD0 U380 ( .I(1'b1), .ZN(n[373]) );
  INVD0 U382 ( .I(1'b1), .ZN(n[380]) );
  INVD0 U384 ( .I(1'b1), .ZN(n[381]) );
  INVD0 U386 ( .I(1'b1), .ZN(n[383]) );
  INVD0 U388 ( .I(1'b1), .ZN(n[384]) );
  INVD0 U390 ( .I(1'b1), .ZN(n[387]) );
  INVD0 U392 ( .I(1'b1), .ZN(n[388]) );
  INVD0 U394 ( .I(1'b1), .ZN(n[390]) );
  INVD0 U396 ( .I(1'b1), .ZN(n[391]) );
  INVD0 U398 ( .I(1'b1), .ZN(n[395]) );
  INVD0 U400 ( .I(1'b1), .ZN(n[396]) );
  INVD0 U402 ( .I(1'b1), .ZN(n[398]) );
  INVD0 U404 ( .I(1'b1), .ZN(n[399]) );
  INVD0 U406 ( .I(1'b1), .ZN(n[402]) );
  INVD0 U408 ( .I(1'b1), .ZN(n[403]) );
  INVD0 U410 ( .I(1'b1), .ZN(n[405]) );
  INVD0 U412 ( .I(1'b1), .ZN(n[406]) );
  INVD0 U414 ( .I(1'b1), .ZN(n[411]) );
  INVD0 U416 ( .I(1'b1), .ZN(n[412]) );
  INVD0 U418 ( .I(1'b1), .ZN(n[414]) );
  INVD0 U420 ( .I(1'b1), .ZN(n[415]) );
  INVD0 U422 ( .I(1'b1), .ZN(n[418]) );
  INVD0 U424 ( .I(1'b1), .ZN(n[419]) );
  INVD0 U426 ( .I(1'b1), .ZN(n[421]) );
  INVD0 U428 ( .I(1'b1), .ZN(n[422]) );
  INVD0 U430 ( .I(1'b1), .ZN(n[426]) );
  INVD0 U432 ( .I(1'b1), .ZN(n[427]) );
  INVD0 U434 ( .I(1'b1), .ZN(n[429]) );
  INVD0 U436 ( .I(1'b1), .ZN(n[430]) );
  INVD0 U438 ( .I(1'b1), .ZN(n[433]) );
  INVD0 U440 ( .I(1'b1), .ZN(n[434]) );
  INVD0 U442 ( .I(1'b1), .ZN(n[436]) );
  INVD0 U444 ( .I(1'b1), .ZN(n[437]) );
  INVD0 U446 ( .I(1'b1), .ZN(n[443]) );
  INVD0 U448 ( .I(1'b1), .ZN(n[444]) );
  INVD0 U450 ( .I(1'b1), .ZN(n[446]) );
  INVD0 U452 ( .I(1'b1), .ZN(n[447]) );
  INVD0 U454 ( .I(1'b1), .ZN(n[450]) );
  INVD0 U456 ( .I(1'b1), .ZN(n[451]) );
  INVD0 U458 ( .I(1'b1), .ZN(n[453]) );
  INVD0 U460 ( .I(1'b1), .ZN(n[454]) );
  INVD0 U462 ( .I(1'b1), .ZN(n[458]) );
  INVD0 U464 ( .I(1'b1), .ZN(n[459]) );
  INVD0 U466 ( .I(1'b1), .ZN(n[461]) );
  INVD0 U468 ( .I(1'b1), .ZN(n[462]) );
  INVD0 U470 ( .I(1'b1), .ZN(n[465]) );
  INVD0 U472 ( .I(1'b1), .ZN(n[466]) );
  INVD0 U474 ( .I(1'b1), .ZN(n[468]) );
  INVD0 U476 ( .I(1'b1), .ZN(n[469]) );
  INVD0 U478 ( .I(1'b1), .ZN(n[474]) );
  INVD0 U480 ( .I(1'b1), .ZN(n[475]) );
  INVD0 U482 ( .I(1'b1), .ZN(n[477]) );
  INVD0 U484 ( .I(1'b1), .ZN(n[478]) );
  INVD0 U486 ( .I(1'b1), .ZN(n[481]) );
  INVD0 U488 ( .I(1'b1), .ZN(n[482]) );
  INVD0 U490 ( .I(1'b1), .ZN(n[484]) );
  INVD0 U492 ( .I(1'b1), .ZN(n[485]) );
  INVD0 U494 ( .I(1'b1), .ZN(n[489]) );
  INVD0 U496 ( .I(1'b1), .ZN(n[490]) );
  INVD0 U498 ( .I(1'b1), .ZN(n[492]) );
  INVD0 U500 ( .I(1'b1), .ZN(n[493]) );
  INVD0 U502 ( .I(1'b1), .ZN(n[496]) );
  INVD0 U504 ( .I(1'b1), .ZN(n[497]) );
  INVD0 U506 ( .I(1'b1), .ZN(n[499]) );
  INVD0 U508 ( .I(1'b1), .ZN(n[500]) );
  INVD0 U510 ( .I(1'b1), .ZN(n[509]) );
  INVD0 U512 ( .I(1'b1), .ZN(n[510]) );
  INVD0 U514 ( .I(1'b1), .ZN(n[512]) );
  INVD0 U516 ( .I(1'b1), .ZN(n[513]) );
  INVD0 U518 ( .I(1'b1), .ZN(n[516]) );
  INVD0 U520 ( .I(1'b1), .ZN(n[517]) );
  INVD0 U522 ( .I(1'b1), .ZN(n[519]) );
  INVD0 U524 ( .I(1'b1), .ZN(n[520]) );
  INVD0 U526 ( .I(1'b1), .ZN(n[524]) );
  INVD0 U528 ( .I(1'b1), .ZN(n[525]) );
  INVD0 U530 ( .I(1'b1), .ZN(n[527]) );
  INVD0 U532 ( .I(1'b1), .ZN(n[528]) );
  INVD0 U534 ( .I(1'b1), .ZN(n[531]) );
  INVD0 U536 ( .I(1'b1), .ZN(n[532]) );
  INVD0 U538 ( .I(1'b1), .ZN(n[534]) );
  INVD0 U540 ( .I(1'b1), .ZN(n[535]) );
  INVD0 U542 ( .I(1'b1), .ZN(n[540]) );
  INVD0 U544 ( .I(1'b1), .ZN(n[541]) );
  INVD0 U546 ( .I(1'b1), .ZN(n[543]) );
  INVD0 U548 ( .I(1'b1), .ZN(n[544]) );
  INVD0 U550 ( .I(1'b1), .ZN(n[547]) );
  INVD0 U552 ( .I(1'b1), .ZN(n[548]) );
  INVD0 U554 ( .I(1'b1), .ZN(n[550]) );
  INVD0 U556 ( .I(1'b1), .ZN(n[551]) );
  INVD0 U558 ( .I(1'b1), .ZN(n[555]) );
  INVD0 U560 ( .I(1'b1), .ZN(n[556]) );
  INVD0 U562 ( .I(1'b1), .ZN(n[558]) );
  INVD0 U564 ( .I(1'b1), .ZN(n[559]) );
  INVD0 U566 ( .I(1'b1), .ZN(n[562]) );
  INVD0 U568 ( .I(1'b1), .ZN(n[563]) );
  INVD0 U570 ( .I(1'b1), .ZN(n[565]) );
  INVD0 U572 ( .I(1'b1), .ZN(n[566]) );
  INVD0 U574 ( .I(1'b1), .ZN(n[572]) );
  INVD0 U576 ( .I(1'b1), .ZN(n[573]) );
  INVD0 U578 ( .I(1'b1), .ZN(n[575]) );
  INVD0 U580 ( .I(1'b1), .ZN(n[576]) );
  INVD0 U582 ( .I(1'b1), .ZN(n[579]) );
  INVD0 U584 ( .I(1'b1), .ZN(n[580]) );
  INVD0 U586 ( .I(1'b1), .ZN(n[582]) );
  INVD0 U588 ( .I(1'b1), .ZN(n[583]) );
  INVD0 U590 ( .I(1'b1), .ZN(n[587]) );
  INVD0 U592 ( .I(1'b1), .ZN(n[588]) );
  INVD0 U594 ( .I(1'b1), .ZN(n[590]) );
  INVD0 U596 ( .I(1'b1), .ZN(n[591]) );
  INVD0 U598 ( .I(1'b1), .ZN(n[594]) );
  INVD0 U600 ( .I(1'b1), .ZN(n[595]) );
  INVD0 U602 ( .I(1'b1), .ZN(n[597]) );
  INVD0 U604 ( .I(1'b1), .ZN(n[598]) );
  INVD0 U606 ( .I(1'b1), .ZN(n[603]) );
  INVD0 U608 ( .I(1'b1), .ZN(n[604]) );
  INVD0 U610 ( .I(1'b1), .ZN(n[606]) );
  INVD0 U612 ( .I(1'b1), .ZN(n[607]) );
  INVD0 U614 ( .I(1'b1), .ZN(n[610]) );
  INVD0 U616 ( .I(1'b1), .ZN(n[611]) );
  INVD0 U618 ( .I(1'b1), .ZN(n[613]) );
  INVD0 U620 ( .I(1'b1), .ZN(n[614]) );
  INVD0 U622 ( .I(1'b1), .ZN(n[618]) );
  INVD0 U624 ( .I(1'b1), .ZN(n[619]) );
  INVD0 U626 ( .I(1'b1), .ZN(n[621]) );
  INVD0 U628 ( .I(1'b1), .ZN(n[622]) );
  INVD0 U630 ( .I(1'b1), .ZN(n[625]) );
  INVD0 U632 ( .I(1'b1), .ZN(n[626]) );
  INVD0 U634 ( .I(1'b1), .ZN(n[628]) );
  INVD0 U636 ( .I(1'b1), .ZN(n[629]) );
  INVD0 U638 ( .I(1'b1), .ZN(n[636]) );
  INVD0 U640 ( .I(1'b1), .ZN(n[637]) );
  INVD0 U642 ( .I(1'b1), .ZN(n[639]) );
  INVD0 U644 ( .I(1'b1), .ZN(n[640]) );
  INVD0 U646 ( .I(1'b1), .ZN(n[643]) );
  INVD0 U648 ( .I(1'b1), .ZN(n[644]) );
  INVD0 U650 ( .I(1'b1), .ZN(n[646]) );
  INVD0 U652 ( .I(1'b1), .ZN(n[647]) );
  INVD0 U654 ( .I(1'b1), .ZN(n[651]) );
  INVD0 U656 ( .I(1'b1), .ZN(n[652]) );
  INVD0 U658 ( .I(1'b1), .ZN(n[654]) );
  INVD0 U660 ( .I(1'b1), .ZN(n[655]) );
  INVD0 U662 ( .I(1'b1), .ZN(n[658]) );
  INVD0 U664 ( .I(1'b1), .ZN(n[659]) );
  INVD0 U666 ( .I(1'b1), .ZN(n[661]) );
  INVD0 U668 ( .I(1'b1), .ZN(n[662]) );
  INVD0 U670 ( .I(1'b1), .ZN(n[667]) );
  INVD0 U672 ( .I(1'b1), .ZN(n[668]) );
  INVD0 U674 ( .I(1'b1), .ZN(n[670]) );
  INVD0 U676 ( .I(1'b1), .ZN(n[671]) );
  INVD0 U678 ( .I(1'b1), .ZN(n[674]) );
  INVD0 U680 ( .I(1'b1), .ZN(n[675]) );
  INVD0 U682 ( .I(1'b1), .ZN(n[677]) );
  INVD0 U684 ( .I(1'b1), .ZN(n[678]) );
  INVD0 U686 ( .I(1'b1), .ZN(n[682]) );
  INVD0 U688 ( .I(1'b1), .ZN(n[683]) );
  INVD0 U690 ( .I(1'b1), .ZN(n[685]) );
  INVD0 U692 ( .I(1'b1), .ZN(n[686]) );
  INVD0 U694 ( .I(1'b1), .ZN(n[689]) );
  INVD0 U696 ( .I(1'b1), .ZN(n[690]) );
  INVD0 U698 ( .I(1'b1), .ZN(n[692]) );
  INVD0 U700 ( .I(1'b1), .ZN(n[693]) );
  INVD0 U702 ( .I(1'b1), .ZN(n[699]) );
  INVD0 U704 ( .I(1'b1), .ZN(n[700]) );
  INVD0 U706 ( .I(1'b1), .ZN(n[702]) );
  INVD0 U708 ( .I(1'b1), .ZN(n[703]) );
  INVD0 U710 ( .I(1'b1), .ZN(n[706]) );
  INVD0 U712 ( .I(1'b1), .ZN(n[707]) );
  INVD0 U714 ( .I(1'b1), .ZN(n[709]) );
  INVD0 U716 ( .I(1'b1), .ZN(n[710]) );
  INVD0 U718 ( .I(1'b1), .ZN(n[714]) );
  INVD0 U720 ( .I(1'b1), .ZN(n[715]) );
  INVD0 U722 ( .I(1'b1), .ZN(n[717]) );
  INVD0 U724 ( .I(1'b1), .ZN(n[718]) );
  INVD0 U726 ( .I(1'b1), .ZN(n[721]) );
  INVD0 U728 ( .I(1'b1), .ZN(n[722]) );
  INVD0 U730 ( .I(1'b1), .ZN(n[724]) );
  INVD0 U732 ( .I(1'b1), .ZN(n[725]) );
  INVD0 U734 ( .I(1'b1), .ZN(n[730]) );
  INVD0 U736 ( .I(1'b1), .ZN(n[731]) );
  INVD0 U738 ( .I(1'b1), .ZN(n[733]) );
  INVD0 U740 ( .I(1'b1), .ZN(n[734]) );
  INVD0 U742 ( .I(1'b1), .ZN(n[737]) );
  INVD0 U744 ( .I(1'b1), .ZN(n[738]) );
  INVD0 U746 ( .I(1'b1), .ZN(n[740]) );
  INVD0 U748 ( .I(1'b1), .ZN(n[741]) );
  INVD0 U750 ( .I(1'b1), .ZN(n[745]) );
  INVD0 U752 ( .I(1'b1), .ZN(n[746]) );
  INVD0 U754 ( .I(1'b1), .ZN(n[748]) );
  INVD0 U756 ( .I(1'b1), .ZN(n[749]) );
  INVD0 U758 ( .I(1'b1), .ZN(n[752]) );
  INVD0 U760 ( .I(1'b1), .ZN(n[753]) );
  INVD0 U762 ( .I(1'b1), .ZN(n[755]) );
  INVD0 U764 ( .I(1'b1), .ZN(n[756]) );
  INVD0 U766 ( .I(1'b1), .ZN(n[764]) );
  INVD0 U768 ( .I(1'b1), .ZN(n[765]) );
  INVD0 U770 ( .I(1'b1), .ZN(n[767]) );
  INVD0 U772 ( .I(1'b1), .ZN(n[768]) );
  INVD0 U774 ( .I(1'b1), .ZN(n[771]) );
  INVD0 U776 ( .I(1'b1), .ZN(n[772]) );
  INVD0 U778 ( .I(1'b1), .ZN(n[774]) );
  INVD0 U780 ( .I(1'b1), .ZN(n[775]) );
  INVD0 U782 ( .I(1'b1), .ZN(n[779]) );
  INVD0 U784 ( .I(1'b1), .ZN(n[780]) );
  INVD0 U786 ( .I(1'b1), .ZN(n[782]) );
  INVD0 U788 ( .I(1'b1), .ZN(n[783]) );
  INVD0 U790 ( .I(1'b1), .ZN(n[786]) );
  INVD0 U792 ( .I(1'b1), .ZN(n[787]) );
  INVD0 U794 ( .I(1'b1), .ZN(n[789]) );
  INVD0 U796 ( .I(1'b1), .ZN(n[790]) );
  INVD0 U798 ( .I(1'b1), .ZN(n[795]) );
  INVD0 U800 ( .I(1'b1), .ZN(n[796]) );
  INVD0 U802 ( .I(1'b1), .ZN(n[798]) );
  INVD0 U804 ( .I(1'b1), .ZN(n[799]) );
  INVD0 U806 ( .I(1'b1), .ZN(n[802]) );
  INVD0 U808 ( .I(1'b1), .ZN(n[803]) );
  INVD0 U810 ( .I(1'b1), .ZN(n[805]) );
  INVD0 U812 ( .I(1'b1), .ZN(n[806]) );
  INVD0 U814 ( .I(1'b1), .ZN(n[810]) );
  INVD0 U816 ( .I(1'b1), .ZN(n[811]) );
  INVD0 U818 ( .I(1'b1), .ZN(n[813]) );
  INVD0 U820 ( .I(1'b1), .ZN(n[814]) );
  INVD0 U822 ( .I(1'b1), .ZN(n[817]) );
  INVD0 U824 ( .I(1'b1), .ZN(n[818]) );
  INVD0 U826 ( .I(1'b1), .ZN(n[820]) );
  INVD0 U828 ( .I(1'b1), .ZN(n[821]) );
  INVD0 U830 ( .I(1'b1), .ZN(n[827]) );
  INVD0 U832 ( .I(1'b1), .ZN(n[828]) );
  INVD0 U834 ( .I(1'b1), .ZN(n[830]) );
  INVD0 U836 ( .I(1'b1), .ZN(n[831]) );
  INVD0 U838 ( .I(1'b1), .ZN(n[834]) );
  INVD0 U840 ( .I(1'b1), .ZN(n[835]) );
  INVD0 U842 ( .I(1'b1), .ZN(n[837]) );
  INVD0 U844 ( .I(1'b1), .ZN(n[838]) );
  INVD0 U846 ( .I(1'b1), .ZN(n[842]) );
  INVD0 U848 ( .I(1'b1), .ZN(n[843]) );
  INVD0 U850 ( .I(1'b1), .ZN(n[845]) );
  INVD0 U852 ( .I(1'b1), .ZN(n[846]) );
  INVD0 U854 ( .I(1'b1), .ZN(n[849]) );
  INVD0 U856 ( .I(1'b1), .ZN(n[850]) );
  INVD0 U858 ( .I(1'b1), .ZN(n[852]) );
  INVD0 U860 ( .I(1'b1), .ZN(n[853]) );
  INVD0 U862 ( .I(1'b1), .ZN(n[858]) );
  INVD0 U864 ( .I(1'b1), .ZN(n[859]) );
  INVD0 U866 ( .I(1'b1), .ZN(n[861]) );
  INVD0 U868 ( .I(1'b1), .ZN(n[862]) );
  INVD0 U870 ( .I(1'b1), .ZN(n[865]) );
  INVD0 U872 ( .I(1'b1), .ZN(n[866]) );
  INVD0 U874 ( .I(1'b1), .ZN(n[868]) );
  INVD0 U876 ( .I(1'b1), .ZN(n[869]) );
  INVD0 U878 ( .I(1'b1), .ZN(n[873]) );
  INVD0 U880 ( .I(1'b1), .ZN(n[874]) );
  INVD0 U882 ( .I(1'b1), .ZN(n[876]) );
  INVD0 U884 ( .I(1'b1), .ZN(n[877]) );
  INVD0 U886 ( .I(1'b1), .ZN(n[880]) );
  INVD0 U888 ( .I(1'b1), .ZN(n[881]) );
  INVD0 U890 ( .I(1'b1), .ZN(n[883]) );
  INVD0 U892 ( .I(1'b1), .ZN(n[884]) );
  INVD0 U894 ( .I(1'b1), .ZN(n[891]) );
  INVD0 U896 ( .I(1'b1), .ZN(n[892]) );
  INVD0 U898 ( .I(1'b1), .ZN(n[894]) );
  INVD0 U900 ( .I(1'b1), .ZN(n[895]) );
  INVD0 U902 ( .I(1'b1), .ZN(n[898]) );
  INVD0 U904 ( .I(1'b1), .ZN(n[899]) );
  INVD0 U906 ( .I(1'b1), .ZN(n[901]) );
  INVD0 U908 ( .I(1'b1), .ZN(n[902]) );
  INVD0 U910 ( .I(1'b1), .ZN(n[906]) );
  INVD0 U912 ( .I(1'b1), .ZN(n[907]) );
  INVD0 U914 ( .I(1'b1), .ZN(n[909]) );
  INVD0 U916 ( .I(1'b1), .ZN(n[910]) );
  INVD0 U918 ( .I(1'b1), .ZN(n[913]) );
  INVD0 U920 ( .I(1'b1), .ZN(n[914]) );
  INVD0 U922 ( .I(1'b1), .ZN(n[916]) );
  INVD0 U924 ( .I(1'b1), .ZN(n[917]) );
  INVD0 U926 ( .I(1'b1), .ZN(n[922]) );
  INVD0 U928 ( .I(1'b1), .ZN(n[923]) );
  INVD0 U930 ( .I(1'b1), .ZN(n[925]) );
  INVD0 U932 ( .I(1'b1), .ZN(n[926]) );
  INVD0 U934 ( .I(1'b1), .ZN(n[929]) );
  INVD0 U936 ( .I(1'b1), .ZN(n[930]) );
  INVD0 U938 ( .I(1'b1), .ZN(n[932]) );
  INVD0 U940 ( .I(1'b1), .ZN(n[933]) );
  INVD0 U942 ( .I(1'b1), .ZN(n[937]) );
  INVD0 U944 ( .I(1'b1), .ZN(n[938]) );
  INVD0 U946 ( .I(1'b1), .ZN(n[940]) );
  INVD0 U948 ( .I(1'b1), .ZN(n[941]) );
  INVD0 U950 ( .I(1'b1), .ZN(n[944]) );
  INVD0 U952 ( .I(1'b1), .ZN(n[945]) );
  INVD0 U954 ( .I(1'b1), .ZN(n[947]) );
  INVD0 U956 ( .I(1'b1), .ZN(n[948]) );
  INVD0 U958 ( .I(1'b1), .ZN(n[954]) );
  INVD0 U960 ( .I(1'b1), .ZN(n[955]) );
  INVD0 U962 ( .I(1'b1), .ZN(n[957]) );
  INVD0 U964 ( .I(1'b1), .ZN(n[958]) );
  INVD0 U966 ( .I(1'b1), .ZN(n[961]) );
  INVD0 U968 ( .I(1'b1), .ZN(n[962]) );
  INVD0 U970 ( .I(1'b1), .ZN(n[964]) );
  INVD0 U972 ( .I(1'b1), .ZN(n[965]) );
  INVD0 U974 ( .I(1'b1), .ZN(n[969]) );
  INVD0 U976 ( .I(1'b1), .ZN(n[970]) );
  INVD0 U978 ( .I(1'b1), .ZN(n[972]) );
  INVD0 U980 ( .I(1'b1), .ZN(n[973]) );
  INVD0 U982 ( .I(1'b1), .ZN(n[976]) );
  INVD0 U984 ( .I(1'b1), .ZN(n[977]) );
  INVD0 U986 ( .I(1'b1), .ZN(n[979]) );
  INVD0 U988 ( .I(1'b1), .ZN(n[980]) );
  INVD0 U990 ( .I(1'b1), .ZN(n[985]) );
  INVD0 U992 ( .I(1'b1), .ZN(n[986]) );
  INVD0 U994 ( .I(1'b1), .ZN(n[988]) );
  INVD0 U996 ( .I(1'b1), .ZN(n[989]) );
  INVD0 U998 ( .I(1'b1), .ZN(n[992]) );
  INVD0 U1000 ( .I(1'b1), .ZN(n[993]) );
  INVD0 U1002 ( .I(1'b1), .ZN(n[995]) );
  INVD0 U1004 ( .I(1'b1), .ZN(n[996]) );
  INVD0 U1006 ( .I(1'b1), .ZN(n[1000]) );
  INVD0 U1008 ( .I(1'b1), .ZN(n[1001]) );
  INVD0 U1010 ( .I(1'b1), .ZN(n[1003]) );
  INVD0 U1012 ( .I(1'b1), .ZN(n[1004]) );
  INVD0 U1014 ( .I(1'b1), .ZN(n[1007]) );
  INVD0 U1017 ( .I(1'b1), .ZN(n[1008]) );
  INVD0 U1019 ( .I(1'b1), .ZN(n[1010]) );
  INVD0 U1021 ( .I(1'b1), .ZN(n[1011]) );
  INVD0 U1023 ( .I(1'b1), .ZN(n[1021]) );
  INVD0 U1025 ( .I(1'b1), .ZN(n[1022]) );
  INVD0 U1027 ( .I(1'b1), .ZN(n[1024]) );
  INVD0 U1029 ( .I(1'b1), .ZN(n[1025]) );
  INVD0 U1031 ( .I(1'b1), .ZN(n[1028]) );
  INVD0 U1033 ( .I(1'b1), .ZN(n[1029]) );
  INVD0 U1035 ( .I(1'b1), .ZN(n[1031]) );
  INVD0 U1037 ( .I(1'b1), .ZN(n[1032]) );
  INVD0 U1039 ( .I(1'b1), .ZN(n[1036]) );
  INVD0 U1041 ( .I(1'b1), .ZN(n[1037]) );
  INVD0 U1043 ( .I(1'b1), .ZN(n[1039]) );
  INVD0 U1045 ( .I(1'b1), .ZN(n[1040]) );
  INVD0 U1047 ( .I(1'b1), .ZN(n[1043]) );
  INVD0 U1049 ( .I(1'b1), .ZN(n[1044]) );
  INVD0 U1051 ( .I(1'b1), .ZN(n[1046]) );
  INVD0 U1053 ( .I(1'b1), .ZN(n[1047]) );
  INVD0 U1055 ( .I(1'b1), .ZN(n[1052]) );
  INVD0 U1057 ( .I(1'b1), .ZN(n[1053]) );
  INVD0 U1059 ( .I(1'b1), .ZN(n[1055]) );
  INVD0 U1061 ( .I(1'b1), .ZN(n[1056]) );
  INVD0 U1063 ( .I(1'b1), .ZN(n[1059]) );
  INVD0 U1065 ( .I(1'b1), .ZN(n[1060]) );
  INVD0 U1067 ( .I(1'b1), .ZN(n[1062]) );
  INVD0 U1069 ( .I(1'b1), .ZN(n[1063]) );
  INVD0 U1071 ( .I(1'b1), .ZN(n[1067]) );
  INVD0 U1073 ( .I(1'b1), .ZN(n[1068]) );
  INVD0 U1075 ( .I(1'b1), .ZN(n[1070]) );
  INVD0 U1077 ( .I(1'b1), .ZN(n[1071]) );
  INVD0 U1079 ( .I(1'b1), .ZN(n[1074]) );
  INVD0 U1081 ( .I(1'b1), .ZN(n[1075]) );
  INVD0 U1083 ( .I(1'b1), .ZN(n[1077]) );
  INVD0 U1085 ( .I(1'b1), .ZN(n[1078]) );
  INVD0 U1087 ( .I(1'b1), .ZN(n[1084]) );
  INVD0 U1089 ( .I(1'b1), .ZN(n[1085]) );
  INVD0 U1091 ( .I(1'b1), .ZN(n[1087]) );
  INVD0 U1093 ( .I(1'b1), .ZN(n[1088]) );
  INVD0 U1095 ( .I(1'b1), .ZN(n[1091]) );
  INVD0 U1097 ( .I(1'b1), .ZN(n[1092]) );
  INVD0 U1099 ( .I(1'b1), .ZN(n[1094]) );
  INVD0 U1101 ( .I(1'b1), .ZN(n[1095]) );
  INVD0 U1103 ( .I(1'b1), .ZN(n[1099]) );
  INVD0 U1105 ( .I(1'b1), .ZN(n[1100]) );
  INVD0 U1107 ( .I(1'b1), .ZN(n[1102]) );
  INVD0 U1109 ( .I(1'b1), .ZN(n[1103]) );
  INVD0 U1111 ( .I(1'b1), .ZN(n[1106]) );
  INVD0 U1113 ( .I(1'b1), .ZN(n[1107]) );
  INVD0 U1115 ( .I(1'b1), .ZN(n[1109]) );
  INVD0 U1117 ( .I(1'b1), .ZN(n[1110]) );
  INVD0 U1119 ( .I(1'b1), .ZN(n[1115]) );
  INVD0 U1121 ( .I(1'b1), .ZN(n[1116]) );
  INVD0 U1123 ( .I(1'b1), .ZN(n[1118]) );
  INVD0 U1125 ( .I(1'b1), .ZN(n[1119]) );
  INVD0 U1127 ( .I(1'b1), .ZN(n[1122]) );
  INVD0 U1129 ( .I(1'b1), .ZN(n[1123]) );
  INVD0 U1131 ( .I(1'b1), .ZN(n[1125]) );
  INVD0 U1133 ( .I(1'b1), .ZN(n[1126]) );
  INVD0 U1135 ( .I(1'b1), .ZN(n[1130]) );
  INVD0 U1137 ( .I(1'b1), .ZN(n[1131]) );
  INVD0 U1139 ( .I(1'b1), .ZN(n[1133]) );
  INVD0 U1141 ( .I(1'b1), .ZN(n[1134]) );
  INVD0 U1143 ( .I(1'b1), .ZN(n[1137]) );
  INVD0 U1145 ( .I(1'b1), .ZN(n[1138]) );
  INVD0 U1147 ( .I(1'b1), .ZN(n[1140]) );
  INVD0 U1149 ( .I(1'b1), .ZN(n[1141]) );
  INVD0 U1151 ( .I(1'b1), .ZN(n[1148]) );
  INVD0 U1153 ( .I(1'b1), .ZN(n[1149]) );
  INVD0 U1155 ( .I(1'b1), .ZN(n[1151]) );
  INVD0 U1157 ( .I(1'b1), .ZN(n[1152]) );
  INVD0 U1159 ( .I(1'b1), .ZN(n[1155]) );
  INVD0 U1161 ( .I(1'b1), .ZN(n[1156]) );
  INVD0 U1163 ( .I(1'b1), .ZN(n[1158]) );
  INVD0 U1165 ( .I(1'b1), .ZN(n[1159]) );
  INVD0 U1167 ( .I(1'b1), .ZN(n[1163]) );
  INVD0 U1169 ( .I(1'b1), .ZN(n[1164]) );
  INVD0 U1171 ( .I(1'b1), .ZN(n[1166]) );
  INVD0 U1173 ( .I(1'b1), .ZN(n[1167]) );
  INVD0 U1175 ( .I(1'b1), .ZN(n[1170]) );
  INVD0 U1177 ( .I(1'b1), .ZN(n[1171]) );
  INVD0 U1179 ( .I(1'b1), .ZN(n[1173]) );
  INVD0 U1181 ( .I(1'b1), .ZN(n[1174]) );
  INVD0 U1183 ( .I(1'b1), .ZN(n[1179]) );
  INVD0 U1185 ( .I(1'b1), .ZN(n[1180]) );
  INVD0 U1187 ( .I(1'b1), .ZN(n[1182]) );
  INVD0 U1189 ( .I(1'b1), .ZN(n[1183]) );
  INVD0 U1191 ( .I(1'b1), .ZN(n[1186]) );
  INVD0 U1193 ( .I(1'b1), .ZN(n[1187]) );
  INVD0 U1195 ( .I(1'b1), .ZN(n[1189]) );
  INVD0 U1197 ( .I(1'b1), .ZN(n[1190]) );
  INVD0 U1199 ( .I(1'b1), .ZN(n[1194]) );
  INVD0 U1201 ( .I(1'b1), .ZN(n[1195]) );
  INVD0 U1203 ( .I(1'b1), .ZN(n[1197]) );
  INVD0 U1205 ( .I(1'b1), .ZN(n[1198]) );
  INVD0 U1207 ( .I(1'b1), .ZN(n[1201]) );
  INVD0 U1209 ( .I(1'b1), .ZN(n[1202]) );
  INVD0 U1211 ( .I(1'b1), .ZN(n[1204]) );
  INVD0 U1213 ( .I(1'b1), .ZN(n[1205]) );
  INVD0 U1215 ( .I(1'b1), .ZN(n[1211]) );
  INVD0 U1217 ( .I(1'b1), .ZN(n[1212]) );
  INVD0 U1219 ( .I(1'b1), .ZN(n[1214]) );
  INVD0 U1221 ( .I(1'b1), .ZN(n[1215]) );
  INVD0 U1223 ( .I(1'b1), .ZN(n[1218]) );
  INVD0 U1225 ( .I(1'b1), .ZN(n[1219]) );
  INVD0 U1227 ( .I(1'b1), .ZN(n[1221]) );
  INVD0 U1229 ( .I(1'b1), .ZN(n[1222]) );
  INVD0 U1231 ( .I(1'b1), .ZN(n[1226]) );
  INVD0 U1233 ( .I(1'b1), .ZN(n[1227]) );
  INVD0 U1235 ( .I(1'b1), .ZN(n[1229]) );
  INVD0 U1237 ( .I(1'b1), .ZN(n[1230]) );
  INVD0 U1239 ( .I(1'b1), .ZN(n[1233]) );
  INVD0 U1241 ( .I(1'b1), .ZN(n[1234]) );
  INVD0 U1243 ( .I(1'b1), .ZN(n[1236]) );
  INVD0 U1245 ( .I(1'b1), .ZN(n[1237]) );
  INVD0 U1247 ( .I(1'b1), .ZN(n[1242]) );
  INVD0 U1249 ( .I(1'b1), .ZN(n[1243]) );
  INVD0 U1251 ( .I(1'b1), .ZN(n[1245]) );
  INVD0 U1253 ( .I(1'b1), .ZN(n[1246]) );
  INVD0 U1255 ( .I(1'b1), .ZN(n[1249]) );
  INVD0 U1257 ( .I(1'b1), .ZN(n[1250]) );
  INVD0 U1259 ( .I(1'b1), .ZN(n[1252]) );
  INVD0 U1261 ( .I(1'b1), .ZN(n[1253]) );
  INVD0 U1263 ( .I(1'b1), .ZN(n[1257]) );
  INVD0 U1265 ( .I(1'b1), .ZN(n[1258]) );
  INVD0 U1267 ( .I(1'b1), .ZN(n[1260]) );
  INVD0 U1269 ( .I(1'b1), .ZN(n[1261]) );
  INVD0 U1271 ( .I(1'b1), .ZN(n[1264]) );
  INVD0 U1273 ( .I(1'b1), .ZN(n[1265]) );
  INVD0 U1275 ( .I(1'b1), .ZN(n[1267]) );
  INVD0 U1277 ( .I(1'b1), .ZN(n[1268]) );
  INVD0 U1279 ( .I(1'b1), .ZN(n[1276]) );
  INVD0 U1281 ( .I(1'b1), .ZN(n[1277]) );
  INVD0 U1283 ( .I(1'b1), .ZN(n[1279]) );
  INVD0 U1285 ( .I(1'b1), .ZN(n[1280]) );
  INVD0 U1287 ( .I(1'b1), .ZN(n[1283]) );
  INVD0 U1289 ( .I(1'b1), .ZN(n[1284]) );
  INVD0 U1291 ( .I(1'b1), .ZN(n[1286]) );
  INVD0 U1293 ( .I(1'b1), .ZN(n[1287]) );
  INVD0 U1295 ( .I(1'b1), .ZN(n[1291]) );
  INVD0 U1297 ( .I(1'b1), .ZN(n[1292]) );
  INVD0 U1299 ( .I(1'b1), .ZN(n[1294]) );
  INVD0 U1301 ( .I(1'b1), .ZN(n[1295]) );
  INVD0 U1303 ( .I(1'b1), .ZN(n[1298]) );
  INVD0 U1305 ( .I(1'b1), .ZN(n[1299]) );
  INVD0 U1307 ( .I(1'b1), .ZN(n[1301]) );
  INVD0 U1309 ( .I(1'b1), .ZN(n[1302]) );
  INVD0 U1311 ( .I(1'b1), .ZN(n[1307]) );
  INVD0 U1313 ( .I(1'b1), .ZN(n[1308]) );
  INVD0 U1315 ( .I(1'b1), .ZN(n[1310]) );
  INVD0 U1317 ( .I(1'b1), .ZN(n[1311]) );
  INVD0 U1319 ( .I(1'b1), .ZN(n[1314]) );
  INVD0 U1321 ( .I(1'b1), .ZN(n[1315]) );
  INVD0 U1323 ( .I(1'b1), .ZN(n[1317]) );
  INVD0 U1325 ( .I(1'b1), .ZN(n[1318]) );
  INVD0 U1327 ( .I(1'b1), .ZN(n[1322]) );
  INVD0 U1329 ( .I(1'b1), .ZN(n[1323]) );
  INVD0 U1331 ( .I(1'b1), .ZN(n[1325]) );
  INVD0 U1333 ( .I(1'b1), .ZN(n[1326]) );
  INVD0 U1335 ( .I(1'b1), .ZN(n[1329]) );
  INVD0 U1337 ( .I(1'b1), .ZN(n[1330]) );
  INVD0 U1339 ( .I(1'b1), .ZN(n[1332]) );
  INVD0 U1341 ( .I(1'b1), .ZN(n[1333]) );
  INVD0 U1343 ( .I(1'b1), .ZN(n[1339]) );
  INVD0 U1345 ( .I(1'b1), .ZN(n[1340]) );
  INVD0 U1347 ( .I(1'b1), .ZN(n[1342]) );
  INVD0 U1349 ( .I(1'b1), .ZN(n[1343]) );
  INVD0 U1351 ( .I(1'b1), .ZN(n[1346]) );
  INVD0 U1353 ( .I(1'b1), .ZN(n[1347]) );
  INVD0 U1355 ( .I(1'b1), .ZN(n[1349]) );
  INVD0 U1357 ( .I(1'b1), .ZN(n[1350]) );
  INVD0 U1359 ( .I(1'b1), .ZN(n[1354]) );
  INVD0 U1361 ( .I(1'b1), .ZN(n[1355]) );
  INVD0 U1363 ( .I(1'b1), .ZN(n[1357]) );
  INVD0 U1365 ( .I(1'b1), .ZN(n[1358]) );
  INVD0 U1367 ( .I(1'b1), .ZN(n[1361]) );
  INVD0 U1369 ( .I(1'b1), .ZN(n[1362]) );
  INVD0 U1371 ( .I(1'b1), .ZN(n[1364]) );
  INVD0 U1373 ( .I(1'b1), .ZN(n[1365]) );
  INVD0 U1375 ( .I(1'b1), .ZN(n[1370]) );
  INVD0 U1377 ( .I(1'b1), .ZN(n[1371]) );
  INVD0 U1379 ( .I(1'b1), .ZN(n[1373]) );
  INVD0 U1381 ( .I(1'b1), .ZN(n[1374]) );
  INVD0 U1383 ( .I(1'b1), .ZN(n[1377]) );
  INVD0 U1385 ( .I(1'b1), .ZN(n[1378]) );
  INVD0 U1387 ( .I(1'b1), .ZN(n[1380]) );
  INVD0 U1389 ( .I(1'b1), .ZN(n[1381]) );
  INVD0 U1391 ( .I(1'b1), .ZN(n[1385]) );
  INVD0 U1393 ( .I(1'b1), .ZN(n[1386]) );
  INVD0 U1395 ( .I(1'b1), .ZN(n[1388]) );
  INVD0 U1397 ( .I(1'b1), .ZN(n[1389]) );
  INVD0 U1399 ( .I(1'b1), .ZN(n[1392]) );
  INVD0 U1401 ( .I(1'b1), .ZN(n[1393]) );
  INVD0 U1403 ( .I(1'b1), .ZN(n[1395]) );
  INVD0 U1405 ( .I(1'b1), .ZN(n[1396]) );
  INVD0 U1407 ( .I(1'b1), .ZN(n[1403]) );
  INVD0 U1409 ( .I(1'b1), .ZN(n[1404]) );
  INVD0 U1411 ( .I(1'b1), .ZN(n[1406]) );
  INVD0 U1413 ( .I(1'b1), .ZN(n[1407]) );
  INVD0 U1415 ( .I(1'b1), .ZN(n[1410]) );
  INVD0 U1417 ( .I(1'b1), .ZN(n[1411]) );
  INVD0 U1419 ( .I(1'b1), .ZN(n[1413]) );
  INVD0 U1421 ( .I(1'b1), .ZN(n[1414]) );
  INVD0 U1423 ( .I(1'b1), .ZN(n[1418]) );
  INVD0 U1425 ( .I(1'b1), .ZN(n[1419]) );
  INVD0 U1427 ( .I(1'b1), .ZN(n[1421]) );
  INVD0 U1429 ( .I(1'b1), .ZN(n[1422]) );
  INVD0 U1431 ( .I(1'b1), .ZN(n[1425]) );
  INVD0 U1433 ( .I(1'b1), .ZN(n[1426]) );
  INVD0 U1435 ( .I(1'b1), .ZN(n[1428]) );
  INVD0 U1437 ( .I(1'b1), .ZN(n[1429]) );
  INVD0 U1439 ( .I(1'b1), .ZN(n[1434]) );
  INVD0 U1441 ( .I(1'b1), .ZN(n[1435]) );
  INVD0 U1443 ( .I(1'b1), .ZN(n[1437]) );
  INVD0 U1445 ( .I(1'b1), .ZN(n[1438]) );
  INVD0 U1447 ( .I(1'b1), .ZN(n[1441]) );
  INVD0 U1449 ( .I(1'b1), .ZN(n[1442]) );
  INVD0 U1451 ( .I(1'b1), .ZN(n[1444]) );
  INVD0 U1453 ( .I(1'b1), .ZN(n[1445]) );
  INVD0 U1455 ( .I(1'b1), .ZN(n[1449]) );
  INVD0 U1457 ( .I(1'b1), .ZN(n[1450]) );
  INVD0 U1459 ( .I(1'b1), .ZN(n[1452]) );
  INVD0 U1461 ( .I(1'b1), .ZN(n[1453]) );
  INVD0 U1463 ( .I(1'b1), .ZN(n[1456]) );
  INVD0 U1465 ( .I(1'b1), .ZN(n[1457]) );
  INVD0 U1467 ( .I(1'b1), .ZN(n[1459]) );
  INVD0 U1469 ( .I(1'b1), .ZN(n[1460]) );
  INVD0 U1471 ( .I(1'b1), .ZN(n[1466]) );
  INVD0 U1473 ( .I(1'b1), .ZN(n[1467]) );
  INVD0 U1475 ( .I(1'b1), .ZN(n[1469]) );
  INVD0 U1477 ( .I(1'b1), .ZN(n[1470]) );
  INVD0 U1479 ( .I(1'b1), .ZN(n[1473]) );
  INVD0 U1481 ( .I(1'b1), .ZN(n[1474]) );
  INVD0 U1483 ( .I(1'b1), .ZN(n[1476]) );
  INVD0 U1485 ( .I(1'b1), .ZN(n[1477]) );
  INVD0 U1487 ( .I(1'b1), .ZN(n[1481]) );
  INVD0 U1489 ( .I(1'b1), .ZN(n[1482]) );
  INVD0 U1491 ( .I(1'b1), .ZN(n[1484]) );
  INVD0 U1493 ( .I(1'b1), .ZN(n[1485]) );
  INVD0 U1495 ( .I(1'b1), .ZN(n[1488]) );
  INVD0 U1497 ( .I(1'b1), .ZN(n[1489]) );
  INVD0 U1499 ( .I(1'b1), .ZN(n[1491]) );
  INVD0 U1501 ( .I(1'b1), .ZN(n[1492]) );
  INVD0 U1503 ( .I(1'b1), .ZN(n[1497]) );
  INVD0 U1505 ( .I(1'b1), .ZN(n[1498]) );
  INVD0 U1507 ( .I(1'b1), .ZN(n[1500]) );
  INVD0 U1509 ( .I(1'b1), .ZN(n[1501]) );
  INVD0 U1511 ( .I(1'b1), .ZN(n[1504]) );
  INVD0 U1513 ( .I(1'b1), .ZN(n[1505]) );
  INVD0 U1515 ( .I(1'b1), .ZN(n[1507]) );
  INVD0 U1517 ( .I(1'b1), .ZN(n[1508]) );
  INVD0 U1519 ( .I(1'b1), .ZN(n[1512]) );
  INVD0 U1521 ( .I(1'b1), .ZN(n[1513]) );
  INVD0 U1523 ( .I(1'b1), .ZN(n[1515]) );
  INVD0 U1525 ( .I(1'b1), .ZN(n[1516]) );
  INVD0 U1527 ( .I(1'b1), .ZN(n[1519]) );
  INVD0 U1529 ( .I(1'b1), .ZN(n[1520]) );
  INVD0 U1531 ( .I(1'b1), .ZN(n[1522]) );
  INVD0 U1533 ( .I(1'b1), .ZN(n[1523]) );
  INVD0 U1535 ( .I(1'b1), .ZN(n[1532]) );
  INVD0 U1537 ( .I(1'b1), .ZN(n[1533]) );
  INVD0 U1539 ( .I(1'b1), .ZN(n[1535]) );
  INVD0 U1541 ( .I(1'b1), .ZN(n[1536]) );
  INVD0 U1543 ( .I(1'b1), .ZN(n[1539]) );
  INVD0 U1545 ( .I(1'b1), .ZN(n[1540]) );
  INVD0 U1547 ( .I(1'b1), .ZN(n[1542]) );
  INVD0 U1549 ( .I(1'b1), .ZN(n[1543]) );
  INVD0 U1551 ( .I(1'b1), .ZN(n[1547]) );
  INVD0 U1553 ( .I(1'b1), .ZN(n[1548]) );
  INVD0 U1555 ( .I(1'b1), .ZN(n[1550]) );
  INVD0 U1557 ( .I(1'b1), .ZN(n[1551]) );
  INVD0 U1559 ( .I(1'b1), .ZN(n[1554]) );
  INVD0 U1561 ( .I(1'b1), .ZN(n[1555]) );
  INVD0 U1563 ( .I(1'b1), .ZN(n[1557]) );
  INVD0 U1565 ( .I(1'b1), .ZN(n[1558]) );
  INVD0 U1567 ( .I(1'b1), .ZN(n[1563]) );
  INVD0 U1569 ( .I(1'b1), .ZN(n[1564]) );
  INVD0 U1571 ( .I(1'b1), .ZN(n[1566]) );
  INVD0 U1573 ( .I(1'b1), .ZN(n[1567]) );
  INVD0 U1575 ( .I(1'b1), .ZN(n[1570]) );
  INVD0 U1577 ( .I(1'b1), .ZN(n[1571]) );
  INVD0 U1579 ( .I(1'b1), .ZN(n[1573]) );
  INVD0 U1581 ( .I(1'b1), .ZN(n[1574]) );
  INVD0 U1583 ( .I(1'b1), .ZN(n[1578]) );
  INVD0 U1585 ( .I(1'b1), .ZN(n[1579]) );
  INVD0 U1587 ( .I(1'b1), .ZN(n[1581]) );
  INVD0 U1589 ( .I(1'b1), .ZN(n[1582]) );
  INVD0 U1591 ( .I(1'b1), .ZN(n[1585]) );
  INVD0 U1593 ( .I(1'b1), .ZN(n[1586]) );
  INVD0 U1595 ( .I(1'b1), .ZN(n[1588]) );
  INVD0 U1597 ( .I(1'b1), .ZN(n[1589]) );
  INVD0 U1599 ( .I(1'b1), .ZN(n[1595]) );
  INVD0 U1601 ( .I(1'b1), .ZN(n[1596]) );
  INVD0 U1603 ( .I(1'b1), .ZN(n[1598]) );
  INVD0 U1605 ( .I(1'b1), .ZN(n[1599]) );
  INVD0 U1607 ( .I(1'b1), .ZN(n[1602]) );
  INVD0 U1609 ( .I(1'b1), .ZN(n[1603]) );
  INVD0 U1611 ( .I(1'b1), .ZN(n[1605]) );
  INVD0 U1613 ( .I(1'b1), .ZN(n[1606]) );
  INVD0 U1615 ( .I(1'b1), .ZN(n[1610]) );
  INVD0 U1617 ( .I(1'b1), .ZN(n[1611]) );
  INVD0 U1619 ( .I(1'b1), .ZN(n[1613]) );
  INVD0 U1621 ( .I(1'b1), .ZN(n[1614]) );
  INVD0 U1623 ( .I(1'b1), .ZN(n[1617]) );
  INVD0 U1625 ( .I(1'b1), .ZN(n[1618]) );
  INVD0 U1627 ( .I(1'b1), .ZN(n[1620]) );
  INVD0 U1629 ( .I(1'b1), .ZN(n[1621]) );
  INVD0 U1631 ( .I(1'b1), .ZN(n[1626]) );
  INVD0 U1633 ( .I(1'b1), .ZN(n[1627]) );
  INVD0 U1635 ( .I(1'b1), .ZN(n[1629]) );
  INVD0 U1637 ( .I(1'b1), .ZN(n[1630]) );
  INVD0 U1639 ( .I(1'b1), .ZN(n[1633]) );
  INVD0 U1641 ( .I(1'b1), .ZN(n[1634]) );
  INVD0 U1643 ( .I(1'b1), .ZN(n[1636]) );
  INVD0 U1645 ( .I(1'b1), .ZN(n[1637]) );
  INVD0 U1647 ( .I(1'b1), .ZN(n[1641]) );
  INVD0 U1649 ( .I(1'b1), .ZN(n[1642]) );
  INVD0 U1651 ( .I(1'b1), .ZN(n[1644]) );
  INVD0 U1653 ( .I(1'b1), .ZN(n[1645]) );
  INVD0 U1655 ( .I(1'b1), .ZN(n[1648]) );
  INVD0 U1657 ( .I(1'b1), .ZN(n[1649]) );
  INVD0 U1659 ( .I(1'b1), .ZN(n[1651]) );
  INVD0 U1661 ( .I(1'b1), .ZN(n[1652]) );
  INVD0 U1663 ( .I(1'b1), .ZN(n[1659]) );
  INVD0 U1665 ( .I(1'b1), .ZN(n[1660]) );
  INVD0 U1667 ( .I(1'b1), .ZN(n[1662]) );
  INVD0 U1669 ( .I(1'b1), .ZN(n[1663]) );
  INVD0 U1671 ( .I(1'b1), .ZN(n[1666]) );
  INVD0 U1673 ( .I(1'b1), .ZN(n[1667]) );
  INVD0 U1675 ( .I(1'b1), .ZN(n[1669]) );
  INVD0 U1677 ( .I(1'b1), .ZN(n[1670]) );
  INVD0 U1679 ( .I(1'b1), .ZN(n[1674]) );
  INVD0 U1681 ( .I(1'b1), .ZN(n[1675]) );
  INVD0 U1683 ( .I(1'b1), .ZN(n[1677]) );
  INVD0 U1685 ( .I(1'b1), .ZN(n[1678]) );
  INVD0 U1687 ( .I(1'b1), .ZN(n[1681]) );
  INVD0 U1689 ( .I(1'b1), .ZN(n[1682]) );
  INVD0 U1691 ( .I(1'b1), .ZN(n[1684]) );
  INVD0 U1693 ( .I(1'b1), .ZN(n[1685]) );
  INVD0 U1695 ( .I(1'b1), .ZN(n[1690]) );
  INVD0 U1697 ( .I(1'b1), .ZN(n[1691]) );
  INVD0 U1699 ( .I(1'b1), .ZN(n[1693]) );
  INVD0 U1701 ( .I(1'b1), .ZN(n[1694]) );
  INVD0 U1703 ( .I(1'b1), .ZN(n[1697]) );
  INVD0 U1705 ( .I(1'b1), .ZN(n[1698]) );
  INVD0 U1707 ( .I(1'b1), .ZN(n[1700]) );
  INVD0 U1709 ( .I(1'b1), .ZN(n[1701]) );
  INVD0 U1711 ( .I(1'b1), .ZN(n[1705]) );
  INVD0 U1713 ( .I(1'b1), .ZN(n[1706]) );
  INVD0 U1715 ( .I(1'b1), .ZN(n[1708]) );
  INVD0 U1717 ( .I(1'b1), .ZN(n[1709]) );
  INVD0 U1719 ( .I(1'b1), .ZN(n[1712]) );
  INVD0 U1721 ( .I(1'b1), .ZN(n[1713]) );
  INVD0 U1723 ( .I(1'b1), .ZN(n[1715]) );
  INVD0 U1725 ( .I(1'b1), .ZN(n[1716]) );
  INVD0 U1727 ( .I(1'b1), .ZN(n[1722]) );
  INVD0 U1729 ( .I(1'b1), .ZN(n[1723]) );
  INVD0 U1731 ( .I(1'b1), .ZN(n[1725]) );
  INVD0 U1733 ( .I(1'b1), .ZN(n[1726]) );
  INVD0 U1735 ( .I(1'b1), .ZN(n[1729]) );
  INVD0 U1737 ( .I(1'b1), .ZN(n[1730]) );
  INVD0 U1739 ( .I(1'b1), .ZN(n[1732]) );
  INVD0 U1741 ( .I(1'b1), .ZN(n[1733]) );
  INVD0 U1743 ( .I(1'b1), .ZN(n[1737]) );
  INVD0 U1745 ( .I(1'b1), .ZN(n[1738]) );
  INVD0 U1747 ( .I(1'b1), .ZN(n[1740]) );
  INVD0 U1749 ( .I(1'b1), .ZN(n[1741]) );
  INVD0 U1751 ( .I(1'b1), .ZN(n[1744]) );
  INVD0 U1753 ( .I(1'b1), .ZN(n[1745]) );
  INVD0 U1755 ( .I(1'b1), .ZN(n[1747]) );
  INVD0 U1757 ( .I(1'b1), .ZN(n[1748]) );
  INVD0 U1759 ( .I(1'b1), .ZN(n[1753]) );
  INVD0 U1761 ( .I(1'b1), .ZN(n[1754]) );
  INVD0 U1763 ( .I(1'b1), .ZN(n[1756]) );
  INVD0 U1765 ( .I(1'b1), .ZN(n[1757]) );
  INVD0 U1767 ( .I(1'b1), .ZN(n[1760]) );
  INVD0 U1769 ( .I(1'b1), .ZN(n[1761]) );
  INVD0 U1771 ( .I(1'b1), .ZN(n[1763]) );
  INVD0 U1773 ( .I(1'b1), .ZN(n[1764]) );
  INVD0 U1775 ( .I(1'b1), .ZN(n[1768]) );
  INVD0 U1777 ( .I(1'b1), .ZN(n[1769]) );
  INVD0 U1779 ( .I(1'b1), .ZN(n[1771]) );
  INVD0 U1781 ( .I(1'b1), .ZN(n[1772]) );
  INVD0 U1783 ( .I(1'b1), .ZN(n[1775]) );
  INVD0 U1785 ( .I(1'b1), .ZN(n[1776]) );
  INVD0 U1787 ( .I(1'b1), .ZN(n[1778]) );
  INVD0 U1789 ( .I(1'b1), .ZN(n[1779]) );
  INVD0 U1791 ( .I(1'b1), .ZN(n[1787]) );
  INVD0 U1793 ( .I(1'b1), .ZN(n[1788]) );
  INVD0 U1795 ( .I(1'b1), .ZN(n[1790]) );
  INVD0 U1797 ( .I(1'b1), .ZN(n[1791]) );
  INVD0 U1799 ( .I(1'b1), .ZN(n[1794]) );
  INVD0 U1801 ( .I(1'b1), .ZN(n[1795]) );
  INVD0 U1803 ( .I(1'b1), .ZN(n[1797]) );
  INVD0 U1805 ( .I(1'b1), .ZN(n[1798]) );
  INVD0 U1807 ( .I(1'b1), .ZN(n[1802]) );
  INVD0 U1809 ( .I(1'b1), .ZN(n[1803]) );
  INVD0 U1811 ( .I(1'b1), .ZN(n[1805]) );
  INVD0 U1813 ( .I(1'b1), .ZN(n[1806]) );
  INVD0 U1815 ( .I(1'b1), .ZN(n[1809]) );
  INVD0 U1817 ( .I(1'b1), .ZN(n[1810]) );
  INVD0 U1819 ( .I(1'b1), .ZN(n[1812]) );
  INVD0 U1821 ( .I(1'b1), .ZN(n[1813]) );
  INVD0 U1823 ( .I(1'b1), .ZN(n[1818]) );
  INVD0 U1825 ( .I(1'b1), .ZN(n[1819]) );
  INVD0 U1827 ( .I(1'b1), .ZN(n[1821]) );
  INVD0 U1829 ( .I(1'b1), .ZN(n[1822]) );
  INVD0 U1831 ( .I(1'b1), .ZN(n[1825]) );
  INVD0 U1833 ( .I(1'b1), .ZN(n[1826]) );
  INVD0 U1835 ( .I(1'b1), .ZN(n[1828]) );
  INVD0 U1837 ( .I(1'b1), .ZN(n[1829]) );
  INVD0 U1839 ( .I(1'b1), .ZN(n[1833]) );
  INVD0 U1841 ( .I(1'b1), .ZN(n[1834]) );
  INVD0 U1843 ( .I(1'b1), .ZN(n[1836]) );
  INVD0 U1845 ( .I(1'b1), .ZN(n[1837]) );
  INVD0 U1847 ( .I(1'b1), .ZN(n[1840]) );
  INVD0 U1849 ( .I(1'b1), .ZN(n[1841]) );
  INVD0 U1851 ( .I(1'b1), .ZN(n[1843]) );
  INVD0 U1853 ( .I(1'b1), .ZN(n[1844]) );
  INVD0 U1855 ( .I(1'b1), .ZN(n[1850]) );
  INVD0 U1857 ( .I(1'b1), .ZN(n[1851]) );
  INVD0 U1859 ( .I(1'b1), .ZN(n[1853]) );
  INVD0 U1861 ( .I(1'b1), .ZN(n[1854]) );
  INVD0 U1863 ( .I(1'b1), .ZN(n[1857]) );
  INVD0 U1865 ( .I(1'b1), .ZN(n[1858]) );
  INVD0 U1867 ( .I(1'b1), .ZN(n[1860]) );
  INVD0 U1869 ( .I(1'b1), .ZN(n[1861]) );
  INVD0 U1871 ( .I(1'b1), .ZN(n[1865]) );
  INVD0 U1873 ( .I(1'b1), .ZN(n[1866]) );
  INVD0 U1875 ( .I(1'b1), .ZN(n[1868]) );
  INVD0 U1877 ( .I(1'b1), .ZN(n[1869]) );
  INVD0 U1879 ( .I(1'b1), .ZN(n[1872]) );
  INVD0 U1881 ( .I(1'b1), .ZN(n[1873]) );
  INVD0 U1883 ( .I(1'b1), .ZN(n[1875]) );
  INVD0 U1885 ( .I(1'b1), .ZN(n[1876]) );
  INVD0 U1887 ( .I(1'b1), .ZN(n[1881]) );
  INVD0 U1889 ( .I(1'b1), .ZN(n[1882]) );
  INVD0 U1891 ( .I(1'b1), .ZN(n[1884]) );
  INVD0 U1893 ( .I(1'b1), .ZN(n[1885]) );
  INVD0 U1895 ( .I(1'b1), .ZN(n[1888]) );
  INVD0 U1897 ( .I(1'b1), .ZN(n[1889]) );
  INVD0 U1899 ( .I(1'b1), .ZN(n[1891]) );
  INVD0 U1901 ( .I(1'b1), .ZN(n[1892]) );
  INVD0 U1903 ( .I(1'b1), .ZN(n[1896]) );
  INVD0 U1905 ( .I(1'b1), .ZN(n[1897]) );
  INVD0 U1907 ( .I(1'b1), .ZN(n[1899]) );
  INVD0 U1909 ( .I(1'b1), .ZN(n[1900]) );
  INVD0 U1911 ( .I(1'b1), .ZN(n[1903]) );
  INVD0 U1913 ( .I(1'b1), .ZN(n[1904]) );
  INVD0 U1915 ( .I(1'b1), .ZN(n[1906]) );
  INVD0 U1917 ( .I(1'b1), .ZN(n[1907]) );
  INVD0 U1919 ( .I(1'b1), .ZN(n[1914]) );
  INVD0 U1921 ( .I(1'b1), .ZN(n[1915]) );
  INVD0 U1923 ( .I(1'b1), .ZN(n[1917]) );
  INVD0 U1925 ( .I(1'b1), .ZN(n[1918]) );
  INVD0 U1927 ( .I(1'b1), .ZN(n[1921]) );
  INVD0 U1929 ( .I(1'b1), .ZN(n[1922]) );
  INVD0 U1931 ( .I(1'b1), .ZN(n[1924]) );
  INVD0 U1933 ( .I(1'b1), .ZN(n[1925]) );
  INVD0 U1935 ( .I(1'b1), .ZN(n[1929]) );
  INVD0 U1937 ( .I(1'b1), .ZN(n[1930]) );
  INVD0 U1939 ( .I(1'b1), .ZN(n[1932]) );
  INVD0 U1941 ( .I(1'b1), .ZN(n[1933]) );
  INVD0 U1943 ( .I(1'b1), .ZN(n[1936]) );
  INVD0 U1945 ( .I(1'b1), .ZN(n[1937]) );
  INVD0 U1947 ( .I(1'b1), .ZN(n[1939]) );
  INVD0 U1949 ( .I(1'b1), .ZN(n[1940]) );
  INVD0 U1951 ( .I(1'b1), .ZN(n[1945]) );
  INVD0 U1953 ( .I(1'b1), .ZN(n[1946]) );
  INVD0 U1955 ( .I(1'b1), .ZN(n[1948]) );
  INVD0 U1957 ( .I(1'b1), .ZN(n[1949]) );
  INVD0 U1959 ( .I(1'b1), .ZN(n[1952]) );
  INVD0 U1961 ( .I(1'b1), .ZN(n[1953]) );
  INVD0 U1963 ( .I(1'b1), .ZN(n[1955]) );
  INVD0 U1965 ( .I(1'b1), .ZN(n[1956]) );
  INVD0 U1967 ( .I(1'b1), .ZN(n[1960]) );
  INVD0 U1969 ( .I(1'b1), .ZN(n[1961]) );
  INVD0 U1971 ( .I(1'b1), .ZN(n[1963]) );
  INVD0 U1973 ( .I(1'b1), .ZN(n[1964]) );
  INVD0 U1975 ( .I(1'b1), .ZN(n[1967]) );
  INVD0 U1977 ( .I(1'b1), .ZN(n[1968]) );
  INVD0 U1979 ( .I(1'b1), .ZN(n[1970]) );
  INVD0 U1981 ( .I(1'b1), .ZN(n[1971]) );
  INVD0 U1983 ( .I(1'b1), .ZN(n[1977]) );
  INVD0 U1985 ( .I(1'b1), .ZN(n[1978]) );
  INVD0 U1987 ( .I(1'b1), .ZN(n[1980]) );
  INVD0 U1989 ( .I(1'b1), .ZN(n[1981]) );
  INVD0 U1991 ( .I(1'b1), .ZN(n[1984]) );
  INVD0 U1993 ( .I(1'b1), .ZN(n[1985]) );
  INVD0 U1995 ( .I(1'b1), .ZN(n[1987]) );
  INVD0 U1997 ( .I(1'b1), .ZN(n[1988]) );
  INVD0 U1999 ( .I(1'b1), .ZN(n[1992]) );
  INVD0 U2001 ( .I(1'b1), .ZN(n[1993]) );
  INVD0 U2003 ( .I(1'b1), .ZN(n[1995]) );
  INVD0 U2005 ( .I(1'b1), .ZN(n[1996]) );
  INVD0 U2007 ( .I(1'b1), .ZN(n[1999]) );
  INVD0 U2009 ( .I(1'b1), .ZN(n[2000]) );
  INVD0 U2011 ( .I(1'b1), .ZN(n[2002]) );
  INVD0 U2013 ( .I(1'b1), .ZN(n[2003]) );
  INVD0 U2015 ( .I(1'b1), .ZN(n[2008]) );
  INVD0 U2017 ( .I(1'b1), .ZN(n[2009]) );
  INVD0 U2019 ( .I(1'b1), .ZN(n[2011]) );
  INVD0 U2021 ( .I(1'b1), .ZN(n[2012]) );
  INVD0 U2023 ( .I(1'b1), .ZN(n[2015]) );
  INVD0 U2025 ( .I(1'b1), .ZN(n[2016]) );
  INVD0 U2027 ( .I(1'b1), .ZN(n[2018]) );
  INVD0 U2029 ( .I(1'b1), .ZN(n[2019]) );
  INVD0 U2031 ( .I(1'b1), .ZN(n[2023]) );
  INVD0 U2033 ( .I(1'b1), .ZN(n[2024]) );
  INVD0 U2035 ( .I(1'b1), .ZN(n[2026]) );
  INVD0 U2037 ( .I(1'b1), .ZN(n[2027]) );
  INVD0 U2039 ( .I(1'b1), .ZN(n[2030]) );
  INVD0 U2041 ( .I(1'b1), .ZN(n[2031]) );
  INVD0 U2043 ( .I(1'b1), .ZN(n[2033]) );
  INVD0 U2045 ( .I(1'b1), .ZN(n[2034]) );
  AN2D0 U2047 ( .A1(b[8]), .A2(n[1009]), .Z(n[2032]) );
  AN2D0 U2048 ( .A1(n[1006]), .A2(b[8]), .Z(n[2029]) );
  AN2D0 U2049 ( .A1(n[1005]), .A2(b[8]), .Z(n[2028]) );
  AN2D0 U2050 ( .A1(n[1002]), .A2(b[8]), .Z(n[2025]) );
  AN2D0 U2051 ( .A1(n[999]), .A2(b[8]), .Z(n[2022]) );
  AN2D0 U2052 ( .A1(n[998]), .A2(b[8]), .Z(n[2021]) );
  AN2D0 U2053 ( .A1(n[997]), .A2(b[8]), .Z(n[2020]) );
  AN2D0 U2054 ( .A1(n[994]), .A2(b[8]), .Z(n[2017]) );
  AN2D0 U2055 ( .A1(n[991]), .A2(b[8]), .Z(n[2014]) );
  AN2D0 U2056 ( .A1(n[990]), .A2(b[8]), .Z(n[2013]) );
  AN2D0 U2057 ( .A1(n[987]), .A2(b[8]), .Z(n[2010]) );
  AN2D0 U2058 ( .A1(n[984]), .A2(b[8]), .Z(n[2007]) );
  AN2D0 U2059 ( .A1(n[983]), .A2(b[8]), .Z(n[2006]) );
  AN2D0 U2060 ( .A1(n[982]), .A2(b[8]), .Z(n[2005]) );
  AN2D0 U2061 ( .A1(n[981]), .A2(b[8]), .Z(n[2004]) );
  AN2D0 U2062 ( .A1(n[978]), .A2(b[8]), .Z(n[2001]) );
  AN2D0 U2063 ( .A1(n[975]), .A2(b[8]), .Z(n[1998]) );
  AN2D0 U2064 ( .A1(n[974]), .A2(b[8]), .Z(n[1997]) );
  AN2D0 U2065 ( .A1(n[971]), .A2(b[8]), .Z(n[1994]) );
  AN2D0 U2066 ( .A1(n[968]), .A2(b[8]), .Z(n[1991]) );
  AN2D0 U2067 ( .A1(n[967]), .A2(b[8]), .Z(n[1990]) );
  AN2D0 U2068 ( .A1(n[966]), .A2(b[8]), .Z(n[1989]) );
  AN2D0 U2069 ( .A1(n[963]), .A2(b[8]), .Z(n[1986]) );
  AN2D0 U2070 ( .A1(n[960]), .A2(b[8]), .Z(n[1983]) );
  AN2D0 U2071 ( .A1(n[959]), .A2(b[8]), .Z(n[1982]) );
  AN2D0 U2072 ( .A1(n[956]), .A2(b[8]), .Z(n[1979]) );
  AN2D0 U2073 ( .A1(n[953]), .A2(b[8]), .Z(n[1976]) );
  AN2D0 U2074 ( .A1(n[952]), .A2(b[8]), .Z(n[1975]) );
  AN2D0 U2075 ( .A1(n[951]), .A2(b[8]), .Z(n[1974]) );
  AN2D0 U2076 ( .A1(n[950]), .A2(b[8]), .Z(n[1973]) );
  AN2D0 U2077 ( .A1(n[949]), .A2(b[8]), .Z(n[1972]) );
  AN2D0 U2078 ( .A1(n[946]), .A2(b[8]), .Z(n[1969]) );
  AN2D0 U2079 ( .A1(n[943]), .A2(b[8]), .Z(n[1966]) );
  AN2D0 U2080 ( .A1(n[942]), .A2(b[8]), .Z(n[1965]) );
  AN2D0 U2081 ( .A1(n[939]), .A2(b[8]), .Z(n[1962]) );
  AN2D0 U2082 ( .A1(n[936]), .A2(b[8]), .Z(n[1959]) );
  AN2D0 U2083 ( .A1(n[935]), .A2(b[8]), .Z(n[1958]) );
  AN2D0 U2084 ( .A1(n[934]), .A2(b[8]), .Z(n[1957]) );
  AN2D0 U2085 ( .A1(n[931]), .A2(b[8]), .Z(n[1954]) );
  AN2D0 U2086 ( .A1(n[928]), .A2(b[8]), .Z(n[1951]) );
  AN2D0 U2087 ( .A1(n[927]), .A2(b[8]), .Z(n[1950]) );
  AN2D0 U2088 ( .A1(n[924]), .A2(b[8]), .Z(n[1947]) );
  AN2D0 U2089 ( .A1(n[921]), .A2(b[8]), .Z(n[1944]) );
  AN2D0 U2090 ( .A1(n[920]), .A2(b[8]), .Z(n[1943]) );
  AN2D0 U2091 ( .A1(n[919]), .A2(b[8]), .Z(n[1942]) );
  AN2D0 U2092 ( .A1(n[918]), .A2(b[8]), .Z(n[1941]) );
  AN2D0 U2093 ( .A1(n[915]), .A2(b[8]), .Z(n[1938]) );
  AN2D0 U2094 ( .A1(n[912]), .A2(b[8]), .Z(n[1935]) );
  AN2D0 U2095 ( .A1(n[911]), .A2(b[8]), .Z(n[1934]) );
  AN2D0 U2096 ( .A1(n[908]), .A2(b[8]), .Z(n[1931]) );
  AN2D0 U2097 ( .A1(n[905]), .A2(b[8]), .Z(n[1928]) );
  AN2D0 U2098 ( .A1(n[904]), .A2(b[8]), .Z(n[1927]) );
  AN2D0 U2099 ( .A1(n[903]), .A2(b[8]), .Z(n[1926]) );
  AN2D0 U2100 ( .A1(n[900]), .A2(b[8]), .Z(n[1923]) );
  AN2D0 U2101 ( .A1(n[897]), .A2(b[8]), .Z(n[1920]) );
  AN2D0 U2102 ( .A1(n[896]), .A2(b[8]), .Z(n[1919]) );
  AN2D0 U2103 ( .A1(n[893]), .A2(b[8]), .Z(n[1916]) );
  AN2D0 U2104 ( .A1(n[890]), .A2(b[8]), .Z(n[1913]) );
  AN2D0 U2105 ( .A1(n[889]), .A2(b[8]), .Z(n[1912]) );
  AN2D0 U2106 ( .A1(n[888]), .A2(b[8]), .Z(n[1911]) );
  AN2D0 U2107 ( .A1(n[887]), .A2(b[8]), .Z(n[1910]) );
  AN2D0 U2108 ( .A1(n[886]), .A2(b[8]), .Z(n[1909]) );
  AN2D0 U2109 ( .A1(n[885]), .A2(b[8]), .Z(n[1908]) );
  AN2D0 U2110 ( .A1(n[882]), .A2(b[8]), .Z(n[1905]) );
  AN2D0 U2111 ( .A1(n[879]), .A2(b[8]), .Z(n[1902]) );
  AN2D0 U2112 ( .A1(n[878]), .A2(b[8]), .Z(n[1901]) );
  AN2D0 U2113 ( .A1(n[875]), .A2(b[8]), .Z(n[1898]) );
  AN2D0 U2114 ( .A1(n[872]), .A2(b[8]), .Z(n[1895]) );
  AN2D0 U2115 ( .A1(n[871]), .A2(b[8]), .Z(n[1894]) );
  AN2D0 U2116 ( .A1(n[870]), .A2(b[8]), .Z(n[1893]) );
  AN2D0 U2117 ( .A1(n[867]), .A2(b[8]), .Z(n[1890]) );
  AN2D0 U2118 ( .A1(n[864]), .A2(b[8]), .Z(n[1887]) );
  AN2D0 U2119 ( .A1(n[863]), .A2(b[8]), .Z(n[1886]) );
  AN2D0 U2120 ( .A1(n[860]), .A2(b[8]), .Z(n[1883]) );
  AN2D0 U2121 ( .A1(n[857]), .A2(b[8]), .Z(n[1880]) );
  AN2D0 U2122 ( .A1(n[856]), .A2(b[8]), .Z(n[1879]) );
  AN2D0 U2123 ( .A1(n[855]), .A2(b[8]), .Z(n[1878]) );
  AN2D0 U2124 ( .A1(n[854]), .A2(b[8]), .Z(n[1877]) );
  AN2D0 U2125 ( .A1(n[851]), .A2(b[8]), .Z(n[1874]) );
  AN2D0 U2126 ( .A1(n[848]), .A2(b[8]), .Z(n[1871]) );
  AN2D0 U2127 ( .A1(n[847]), .A2(b[8]), .Z(n[1870]) );
  AN2D0 U2128 ( .A1(n[844]), .A2(b[8]), .Z(n[1867]) );
  AN2D0 U2129 ( .A1(n[841]), .A2(b[8]), .Z(n[1864]) );
  AN2D0 U2130 ( .A1(n[840]), .A2(b[8]), .Z(n[1863]) );
  AN2D0 U2131 ( .A1(n[839]), .A2(b[8]), .Z(n[1862]) );
  AN2D0 U2132 ( .A1(n[836]), .A2(b[8]), .Z(n[1859]) );
  AN2D0 U2133 ( .A1(n[833]), .A2(b[8]), .Z(n[1856]) );
  AN2D0 U2134 ( .A1(n[832]), .A2(b[8]), .Z(n[1855]) );
  AN2D0 U2135 ( .A1(n[829]), .A2(b[8]), .Z(n[1852]) );
  AN2D0 U2136 ( .A1(n[826]), .A2(b[8]), .Z(n[1849]) );
  AN2D0 U2137 ( .A1(n[825]), .A2(b[8]), .Z(n[1848]) );
  AN2D0 U2138 ( .A1(n[824]), .A2(b[8]), .Z(n[1847]) );
  AN2D0 U2139 ( .A1(n[823]), .A2(b[8]), .Z(n[1846]) );
  AN2D0 U2140 ( .A1(n[822]), .A2(b[8]), .Z(n[1845]) );
  AN2D0 U2141 ( .A1(n[819]), .A2(b[8]), .Z(n[1842]) );
  AN2D0 U2142 ( .A1(n[816]), .A2(b[8]), .Z(n[1839]) );
  AN2D0 U2143 ( .A1(n[815]), .A2(b[8]), .Z(n[1838]) );
  AN2D0 U2144 ( .A1(n[812]), .A2(b[8]), .Z(n[1835]) );
  AN2D0 U2145 ( .A1(n[809]), .A2(b[8]), .Z(n[1832]) );
  AN2D0 U2146 ( .A1(n[808]), .A2(b[8]), .Z(n[1831]) );
  AN2D0 U2147 ( .A1(n[807]), .A2(b[8]), .Z(n[1830]) );
  AN2D0 U2148 ( .A1(n[804]), .A2(b[8]), .Z(n[1827]) );
  AN2D0 U2149 ( .A1(n[801]), .A2(b[8]), .Z(n[1824]) );
  AN2D0 U2150 ( .A1(n[800]), .A2(b[8]), .Z(n[1823]) );
  AN2D0 U2151 ( .A1(n[797]), .A2(b[8]), .Z(n[1820]) );
  AN2D0 U2152 ( .A1(n[794]), .A2(b[8]), .Z(n[1817]) );
  AN2D0 U2153 ( .A1(n[793]), .A2(b[8]), .Z(n[1816]) );
  AN2D0 U2154 ( .A1(n[792]), .A2(b[8]), .Z(n[1815]) );
  AN2D0 U2155 ( .A1(n[791]), .A2(b[8]), .Z(n[1814]) );
  AN2D0 U2156 ( .A1(n[788]), .A2(b[8]), .Z(n[1811]) );
  AN2D0 U2157 ( .A1(n[785]), .A2(b[8]), .Z(n[1808]) );
  AN2D0 U2158 ( .A1(n[784]), .A2(b[8]), .Z(n[1807]) );
  AN2D0 U2159 ( .A1(n[781]), .A2(b[8]), .Z(n[1804]) );
  AN2D0 U2160 ( .A1(n[778]), .A2(b[8]), .Z(n[1801]) );
  AN2D0 U2161 ( .A1(n[777]), .A2(b[8]), .Z(n[1800]) );
  AN2D0 U2162 ( .A1(n[776]), .A2(b[8]), .Z(n[1799]) );
  AN2D0 U2163 ( .A1(n[773]), .A2(b[8]), .Z(n[1796]) );
  AN2D0 U2164 ( .A1(n[770]), .A2(b[8]), .Z(n[1793]) );
  AN2D0 U2165 ( .A1(n[769]), .A2(b[8]), .Z(n[1792]) );
  AN2D0 U2166 ( .A1(n[766]), .A2(b[8]), .Z(n[1789]) );
  AN2D0 U2167 ( .A1(n[763]), .A2(b[8]), .Z(n[1786]) );
  AN2D0 U2168 ( .A1(n[762]), .A2(b[8]), .Z(n[1785]) );
  AN2D0 U2169 ( .A1(n[761]), .A2(b[8]), .Z(n[1784]) );
  AN2D0 U2170 ( .A1(n[760]), .A2(b[8]), .Z(n[1783]) );
  AN2D0 U2171 ( .A1(n[759]), .A2(b[8]), .Z(n[1782]) );
  AN2D0 U2172 ( .A1(n[758]), .A2(b[8]), .Z(n[1781]) );
  AN2D0 U2173 ( .A1(n[757]), .A2(b[8]), .Z(n[1780]) );
  AN2D0 U2174 ( .A1(n[754]), .A2(b[8]), .Z(n[1777]) );
  AN2D0 U2175 ( .A1(n[751]), .A2(b[8]), .Z(n[1774]) );
  AN2D0 U2176 ( .A1(n[750]), .A2(b[8]), .Z(n[1773]) );
  AN2D0 U2177 ( .A1(n[747]), .A2(b[8]), .Z(n[1770]) );
  AN2D0 U2178 ( .A1(n[744]), .A2(b[8]), .Z(n[1767]) );
  AN2D0 U2179 ( .A1(n[743]), .A2(b[8]), .Z(n[1766]) );
  AN2D0 U2180 ( .A1(n[742]), .A2(b[8]), .Z(n[1765]) );
  AN2D0 U2181 ( .A1(n[739]), .A2(b[8]), .Z(n[1762]) );
  AN2D0 U2182 ( .A1(n[736]), .A2(b[8]), .Z(n[1759]) );
  AN2D0 U2183 ( .A1(n[735]), .A2(b[8]), .Z(n[1758]) );
  AN2D0 U2184 ( .A1(n[732]), .A2(b[8]), .Z(n[1755]) );
  AN2D0 U2185 ( .A1(n[729]), .A2(b[8]), .Z(n[1752]) );
  AN2D0 U2186 ( .A1(n[728]), .A2(b[8]), .Z(n[1751]) );
  AN2D0 U2187 ( .A1(n[727]), .A2(b[8]), .Z(n[1750]) );
  AN2D0 U2188 ( .A1(n[726]), .A2(b[8]), .Z(n[1749]) );
  AN2D0 U2189 ( .A1(n[723]), .A2(b[8]), .Z(n[1746]) );
  AN2D0 U2190 ( .A1(n[720]), .A2(b[8]), .Z(n[1743]) );
  AN2D0 U2191 ( .A1(n[719]), .A2(b[8]), .Z(n[1742]) );
  AN2D0 U2192 ( .A1(n[716]), .A2(b[8]), .Z(n[1739]) );
  AN2D0 U2193 ( .A1(n[713]), .A2(b[8]), .Z(n[1736]) );
  AN2D0 U2194 ( .A1(n[712]), .A2(b[8]), .Z(n[1735]) );
  AN2D0 U2195 ( .A1(n[711]), .A2(b[8]), .Z(n[1734]) );
  AN2D0 U2196 ( .A1(n[708]), .A2(b[8]), .Z(n[1731]) );
  AN2D0 U2197 ( .A1(n[705]), .A2(b[8]), .Z(n[1728]) );
  AN2D0 U2198 ( .A1(n[704]), .A2(b[8]), .Z(n[1727]) );
  AN2D0 U2199 ( .A1(n[701]), .A2(b[8]), .Z(n[1724]) );
  AN2D0 U2200 ( .A1(n[698]), .A2(b[8]), .Z(n[1721]) );
  AN2D0 U2201 ( .A1(n[697]), .A2(b[8]), .Z(n[1720]) );
  AN2D0 U2202 ( .A1(n[696]), .A2(b[8]), .Z(n[1719]) );
  AN2D0 U2203 ( .A1(n[695]), .A2(b[8]), .Z(n[1718]) );
  AN2D0 U2204 ( .A1(n[694]), .A2(b[8]), .Z(n[1717]) );
  AN2D0 U2205 ( .A1(n[691]), .A2(b[8]), .Z(n[1714]) );
  AN2D0 U2206 ( .A1(n[688]), .A2(b[8]), .Z(n[1711]) );
  AN2D0 U2207 ( .A1(n[687]), .A2(b[8]), .Z(n[1710]) );
  AN2D0 U2208 ( .A1(n[684]), .A2(b[8]), .Z(n[1707]) );
  AN2D0 U2209 ( .A1(n[681]), .A2(b[8]), .Z(n[1704]) );
  AN2D0 U2210 ( .A1(n[680]), .A2(b[8]), .Z(n[1703]) );
  AN2D0 U2211 ( .A1(n[679]), .A2(b[8]), .Z(n[1702]) );
  AN2D0 U2212 ( .A1(n[676]), .A2(b[8]), .Z(n[1699]) );
  AN2D0 U2213 ( .A1(n[673]), .A2(b[8]), .Z(n[1696]) );
  AN2D0 U2214 ( .A1(n[672]), .A2(b[8]), .Z(n[1695]) );
  AN2D0 U2215 ( .A1(n[669]), .A2(b[8]), .Z(n[1692]) );
  AN2D0 U2216 ( .A1(n[666]), .A2(b[8]), .Z(n[1689]) );
  AN2D0 U2217 ( .A1(n[665]), .A2(b[8]), .Z(n[1688]) );
  AN2D0 U2218 ( .A1(n[664]), .A2(b[8]), .Z(n[1687]) );
  AN2D0 U2219 ( .A1(n[663]), .A2(b[8]), .Z(n[1686]) );
  AN2D0 U2220 ( .A1(n[660]), .A2(b[8]), .Z(n[1683]) );
  AN2D0 U2221 ( .A1(n[657]), .A2(b[8]), .Z(n[1680]) );
  AN2D0 U2222 ( .A1(n[656]), .A2(b[8]), .Z(n[1679]) );
  AN2D0 U2223 ( .A1(n[653]), .A2(b[8]), .Z(n[1676]) );
  AN2D0 U2224 ( .A1(n[650]), .A2(b[8]), .Z(n[1673]) );
  AN2D0 U2225 ( .A1(n[649]), .A2(b[8]), .Z(n[1672]) );
  AN2D0 U2226 ( .A1(n[648]), .A2(b[8]), .Z(n[1671]) );
  AN2D0 U2227 ( .A1(n[645]), .A2(b[8]), .Z(n[1668]) );
  AN2D0 U2228 ( .A1(n[642]), .A2(b[8]), .Z(n[1665]) );
  AN2D0 U2229 ( .A1(n[641]), .A2(b[8]), .Z(n[1664]) );
  AN2D0 U2230 ( .A1(n[638]), .A2(b[8]), .Z(n[1661]) );
  AN2D0 U2231 ( .A1(n[635]), .A2(b[8]), .Z(n[1658]) );
  AN2D0 U2232 ( .A1(n[634]), .A2(b[8]), .Z(n[1657]) );
  AN2D0 U2233 ( .A1(n[633]), .A2(b[8]), .Z(n[1656]) );
  AN2D0 U2234 ( .A1(n[632]), .A2(b[8]), .Z(n[1655]) );
  AN2D0 U2235 ( .A1(n[631]), .A2(b[8]), .Z(n[1654]) );
  AN2D0 U2236 ( .A1(n[630]), .A2(b[8]), .Z(n[1653]) );
  AN2D0 U2237 ( .A1(n[627]), .A2(b[8]), .Z(n[1650]) );
  AN2D0 U2238 ( .A1(n[624]), .A2(b[8]), .Z(n[1647]) );
  AN2D0 U2239 ( .A1(n[623]), .A2(b[8]), .Z(n[1646]) );
  AN2D0 U2240 ( .A1(n[620]), .A2(b[8]), .Z(n[1643]) );
  AN2D0 U2241 ( .A1(n[617]), .A2(b[8]), .Z(n[1640]) );
  AN2D0 U2242 ( .A1(n[616]), .A2(b[8]), .Z(n[1639]) );
  AN2D0 U2243 ( .A1(n[615]), .A2(b[8]), .Z(n[1638]) );
  AN2D0 U2244 ( .A1(n[612]), .A2(b[8]), .Z(n[1635]) );
  AN2D0 U2245 ( .A1(n[609]), .A2(b[8]), .Z(n[1632]) );
  AN2D0 U2246 ( .A1(n[608]), .A2(b[8]), .Z(n[1631]) );
  AN2D0 U2247 ( .A1(n[605]), .A2(b[8]), .Z(n[1628]) );
  AN2D0 U2248 ( .A1(n[602]), .A2(b[8]), .Z(n[1625]) );
  AN2D0 U2249 ( .A1(n[601]), .A2(b[8]), .Z(n[1624]) );
  AN2D0 U2250 ( .A1(n[600]), .A2(b[8]), .Z(n[1623]) );
  AN2D0 U2251 ( .A1(n[599]), .A2(b[8]), .Z(n[1622]) );
  AN2D0 U2252 ( .A1(n[596]), .A2(b[8]), .Z(n[1619]) );
  AN2D0 U2253 ( .A1(n[593]), .A2(b[8]), .Z(n[1616]) );
  AN2D0 U2254 ( .A1(n[592]), .A2(b[8]), .Z(n[1615]) );
  AN2D0 U2255 ( .A1(n[589]), .A2(b[8]), .Z(n[1612]) );
  AN2D0 U2256 ( .A1(n[586]), .A2(b[8]), .Z(n[1609]) );
  AN2D0 U2257 ( .A1(n[585]), .A2(b[8]), .Z(n[1608]) );
  AN2D0 U2258 ( .A1(n[584]), .A2(b[8]), .Z(n[1607]) );
  AN2D0 U2259 ( .A1(n[581]), .A2(b[8]), .Z(n[1604]) );
  AN2D0 U2260 ( .A1(n[578]), .A2(b[8]), .Z(n[1601]) );
  AN2D0 U2261 ( .A1(n[577]), .A2(b[8]), .Z(n[1600]) );
  AN2D0 U2262 ( .A1(n[574]), .A2(b[8]), .Z(n[1597]) );
  AN2D0 U2263 ( .A1(n[571]), .A2(b[8]), .Z(n[1594]) );
  AN2D0 U2264 ( .A1(n[570]), .A2(b[8]), .Z(n[1593]) );
  AN2D0 U2265 ( .A1(n[569]), .A2(b[8]), .Z(n[1592]) );
  AN2D0 U2266 ( .A1(n[568]), .A2(b[8]), .Z(n[1591]) );
  AN2D0 U2267 ( .A1(n[567]), .A2(b[8]), .Z(n[1590]) );
  AN2D0 U2268 ( .A1(n[564]), .A2(b[8]), .Z(n[1587]) );
  AN2D0 U2269 ( .A1(n[561]), .A2(b[8]), .Z(n[1584]) );
  AN2D0 U2270 ( .A1(n[560]), .A2(b[8]), .Z(n[1583]) );
  AN2D0 U2271 ( .A1(n[557]), .A2(b[8]), .Z(n[1580]) );
  AN2D0 U2272 ( .A1(n[554]), .A2(b[8]), .Z(n[1577]) );
  AN2D0 U2273 ( .A1(n[553]), .A2(b[8]), .Z(n[1576]) );
  AN2D0 U2274 ( .A1(n[552]), .A2(b[8]), .Z(n[1575]) );
  AN2D0 U2275 ( .A1(n[549]), .A2(b[8]), .Z(n[1572]) );
  AN2D0 U2276 ( .A1(n[546]), .A2(b[8]), .Z(n[1569]) );
  AN2D0 U2277 ( .A1(n[545]), .A2(b[8]), .Z(n[1568]) );
  AN2D0 U2278 ( .A1(n[542]), .A2(b[8]), .Z(n[1565]) );
  AN2D0 U2279 ( .A1(n[539]), .A2(b[8]), .Z(n[1562]) );
  AN2D0 U2280 ( .A1(n[538]), .A2(b[8]), .Z(n[1561]) );
  AN2D0 U2281 ( .A1(n[537]), .A2(b[8]), .Z(n[1560]) );
  AN2D0 U2282 ( .A1(n[536]), .A2(b[8]), .Z(n[1559]) );
  AN2D0 U2283 ( .A1(n[533]), .A2(b[8]), .Z(n[1556]) );
  AN2D0 U2284 ( .A1(n[530]), .A2(b[8]), .Z(n[1553]) );
  AN2D0 U2285 ( .A1(n[529]), .A2(b[8]), .Z(n[1552]) );
  AN2D0 U2286 ( .A1(n[526]), .A2(b[8]), .Z(n[1549]) );
  AN2D0 U2287 ( .A1(n[523]), .A2(b[8]), .Z(n[1546]) );
  AN2D0 U2288 ( .A1(n[522]), .A2(b[8]), .Z(n[1545]) );
  AN2D0 U2289 ( .A1(n[521]), .A2(b[8]), .Z(n[1544]) );
  AN2D0 U2290 ( .A1(n[518]), .A2(b[8]), .Z(n[1541]) );
  AN2D0 U2291 ( .A1(n[515]), .A2(b[8]), .Z(n[1538]) );
  AN2D0 U2292 ( .A1(n[514]), .A2(b[8]), .Z(n[1537]) );
  AN2D0 U2293 ( .A1(n[511]), .A2(b[8]), .Z(n[1534]) );
  AN2D0 U2294 ( .A1(n[508]), .A2(b[8]), .Z(n[1531]) );
  AN2D0 U2295 ( .A1(n[507]), .A2(b[8]), .Z(n[1530]) );
  AN2D0 U2296 ( .A1(n[506]), .A2(b[8]), .Z(n[1529]) );
  AN2D0 U2297 ( .A1(n[505]), .A2(b[8]), .Z(n[1528]) );
  AN2D0 U2298 ( .A1(n[504]), .A2(b[8]), .Z(n[1527]) );
  AN2D0 U2299 ( .A1(n[503]), .A2(b[8]), .Z(n[1526]) );
  AN2D0 U2300 ( .A1(n[502]), .A2(b[8]), .Z(n[1525]) );
  AN2D0 U2301 ( .A1(n[501]), .A2(b[8]), .Z(n[1524]) );
  AN2D0 U2302 ( .A1(a[8]), .A2(n[1009]), .Z(n[1521]) );
  AN2D0 U2303 ( .A1(a[8]), .A2(n[1006]), .Z(n[1518]) );
  AN2D0 U2304 ( .A1(a[8]), .A2(n[1005]), .Z(n[1517]) );
  AN2D0 U2305 ( .A1(a[8]), .A2(n[1002]), .Z(n[1514]) );
  AN2D0 U2306 ( .A1(a[8]), .A2(n[999]), .Z(n[1511]) );
  AN2D0 U2307 ( .A1(n[488]), .A2(b[7]), .Z(n[999]) );
  AN2D0 U2308 ( .A1(a[8]), .A2(n[998]), .Z(n[1510]) );
  AN2D0 U2309 ( .A1(b[7]), .A2(n[487]), .Z(n[998]) );
  AN2D0 U2310 ( .A1(a[8]), .A2(n[997]), .Z(n[1509]) );
  AN2D0 U2311 ( .A1(b[7]), .A2(n[486]), .Z(n[997]) );
  AN2D0 U2312 ( .A1(a[8]), .A2(n[994]), .Z(n[1506]) );
  AN2D0 U2313 ( .A1(b[7]), .A2(n[483]), .Z(n[994]) );
  AN2D0 U2314 ( .A1(a[8]), .A2(n[991]), .Z(n[1503]) );
  AN2D0 U2315 ( .A1(b[7]), .A2(n[480]), .Z(n[991]) );
  AN2D0 U2316 ( .A1(a[8]), .A2(n[990]), .Z(n[1502]) );
  AN2D0 U2317 ( .A1(b[7]), .A2(n[479]), .Z(n[990]) );
  AN2D0 U2318 ( .A1(a[8]), .A2(n[987]), .Z(n[1499]) );
  AN2D0 U2319 ( .A1(b[7]), .A2(n[476]), .Z(n[987]) );
  AN2D0 U2320 ( .A1(a[8]), .A2(n[984]), .Z(n[1496]) );
  AN2D0 U2321 ( .A1(b[7]), .A2(n[473]), .Z(n[984]) );
  AN2D0 U2322 ( .A1(a[8]), .A2(n[983]), .Z(n[1495]) );
  AN2D0 U2323 ( .A1(b[7]), .A2(n[472]), .Z(n[983]) );
  AN2D0 U2324 ( .A1(a[8]), .A2(n[982]), .Z(n[1494]) );
  AN2D0 U2325 ( .A1(b[7]), .A2(n[471]), .Z(n[982]) );
  AN2D0 U2326 ( .A1(a[8]), .A2(n[981]), .Z(n[1493]) );
  AN2D0 U2327 ( .A1(b[7]), .A2(n[470]), .Z(n[981]) );
  AN2D0 U2328 ( .A1(a[8]), .A2(n[978]), .Z(n[1490]) );
  AN2D0 U2329 ( .A1(b[7]), .A2(n[467]), .Z(n[978]) );
  AN2D0 U2330 ( .A1(a[8]), .A2(n[975]), .Z(n[1487]) );
  AN2D0 U2331 ( .A1(b[7]), .A2(n[464]), .Z(n[975]) );
  AN2D0 U2332 ( .A1(a[8]), .A2(n[974]), .Z(n[1486]) );
  AN2D0 U2333 ( .A1(b[7]), .A2(n[463]), .Z(n[974]) );
  AN2D0 U2334 ( .A1(a[8]), .A2(n[971]), .Z(n[1483]) );
  AN2D0 U2335 ( .A1(b[7]), .A2(n[460]), .Z(n[971]) );
  AN2D0 U2336 ( .A1(a[8]), .A2(n[968]), .Z(n[1480]) );
  AN2D0 U2337 ( .A1(b[7]), .A2(n[457]), .Z(n[968]) );
  AN2D0 U2338 ( .A1(a[8]), .A2(n[967]), .Z(n[1479]) );
  AN2D0 U2339 ( .A1(b[7]), .A2(n[456]), .Z(n[967]) );
  AN2D0 U2340 ( .A1(a[8]), .A2(n[966]), .Z(n[1478]) );
  AN2D0 U2341 ( .A1(b[7]), .A2(n[455]), .Z(n[966]) );
  AN2D0 U2342 ( .A1(a[8]), .A2(n[963]), .Z(n[1475]) );
  AN2D0 U2343 ( .A1(b[7]), .A2(n[452]), .Z(n[963]) );
  AN2D0 U2344 ( .A1(a[8]), .A2(n[960]), .Z(n[1472]) );
  AN2D0 U2345 ( .A1(b[7]), .A2(n[449]), .Z(n[960]) );
  AN2D0 U2346 ( .A1(a[8]), .A2(n[959]), .Z(n[1471]) );
  AN2D0 U2347 ( .A1(b[7]), .A2(n[448]), .Z(n[959]) );
  AN2D0 U2348 ( .A1(a[8]), .A2(n[956]), .Z(n[1468]) );
  AN2D0 U2349 ( .A1(b[7]), .A2(n[445]), .Z(n[956]) );
  AN2D0 U2350 ( .A1(a[8]), .A2(n[953]), .Z(n[1465]) );
  AN2D0 U2351 ( .A1(b[7]), .A2(n[442]), .Z(n[953]) );
  AN2D0 U2352 ( .A1(a[8]), .A2(n[952]), .Z(n[1464]) );
  AN2D0 U2353 ( .A1(b[7]), .A2(n[441]), .Z(n[952]) );
  AN2D0 U2354 ( .A1(a[8]), .A2(n[951]), .Z(n[1463]) );
  AN2D0 U2355 ( .A1(b[7]), .A2(n[440]), .Z(n[951]) );
  AN2D0 U2356 ( .A1(a[8]), .A2(n[950]), .Z(n[1462]) );
  AN2D0 U2357 ( .A1(b[7]), .A2(n[439]), .Z(n[950]) );
  AN2D0 U2358 ( .A1(a[8]), .A2(n[949]), .Z(n[1461]) );
  AN2D0 U2359 ( .A1(b[7]), .A2(n[438]), .Z(n[949]) );
  AN2D0 U2360 ( .A1(a[8]), .A2(n[946]), .Z(n[1458]) );
  AN2D0 U2361 ( .A1(b[7]), .A2(n[435]), .Z(n[946]) );
  AN2D0 U2362 ( .A1(a[8]), .A2(n[943]), .Z(n[1455]) );
  AN2D0 U2363 ( .A1(b[7]), .A2(n[432]), .Z(n[943]) );
  AN2D0 U2364 ( .A1(a[8]), .A2(n[942]), .Z(n[1454]) );
  AN2D0 U2365 ( .A1(b[7]), .A2(n[431]), .Z(n[942]) );
  AN2D0 U2366 ( .A1(a[8]), .A2(n[939]), .Z(n[1451]) );
  AN2D0 U2367 ( .A1(b[7]), .A2(n[428]), .Z(n[939]) );
  AN2D0 U2368 ( .A1(a[8]), .A2(n[936]), .Z(n[1448]) );
  AN2D0 U2369 ( .A1(b[7]), .A2(n[425]), .Z(n[936]) );
  AN2D0 U2370 ( .A1(a[8]), .A2(n[935]), .Z(n[1447]) );
  AN2D0 U2371 ( .A1(b[7]), .A2(n[424]), .Z(n[935]) );
  AN2D0 U2372 ( .A1(a[8]), .A2(n[934]), .Z(n[1446]) );
  AN2D0 U2373 ( .A1(b[7]), .A2(n[423]), .Z(n[934]) );
  AN2D0 U2374 ( .A1(a[8]), .A2(n[931]), .Z(n[1443]) );
  AN2D0 U2375 ( .A1(b[7]), .A2(n[420]), .Z(n[931]) );
  AN2D0 U2376 ( .A1(a[8]), .A2(n[928]), .Z(n[1440]) );
  AN2D0 U2377 ( .A1(b[7]), .A2(n[417]), .Z(n[928]) );
  AN2D0 U2378 ( .A1(a[8]), .A2(n[927]), .Z(n[1439]) );
  AN2D0 U2379 ( .A1(b[7]), .A2(n[416]), .Z(n[927]) );
  AN2D0 U2380 ( .A1(a[8]), .A2(n[924]), .Z(n[1436]) );
  AN2D0 U2381 ( .A1(b[7]), .A2(n[413]), .Z(n[924]) );
  AN2D0 U2382 ( .A1(a[8]), .A2(n[921]), .Z(n[1433]) );
  AN2D0 U2383 ( .A1(b[7]), .A2(n[410]), .Z(n[921]) );
  AN2D0 U2384 ( .A1(a[8]), .A2(n[920]), .Z(n[1432]) );
  AN2D0 U2385 ( .A1(b[7]), .A2(n[409]), .Z(n[920]) );
  AN2D0 U2386 ( .A1(a[8]), .A2(n[919]), .Z(n[1431]) );
  AN2D0 U2387 ( .A1(b[7]), .A2(n[408]), .Z(n[919]) );
  AN2D0 U2388 ( .A1(a[8]), .A2(n[918]), .Z(n[1430]) );
  AN2D0 U2389 ( .A1(b[7]), .A2(n[407]), .Z(n[918]) );
  AN2D0 U2390 ( .A1(a[8]), .A2(n[915]), .Z(n[1427]) );
  AN2D0 U2391 ( .A1(b[7]), .A2(n[404]), .Z(n[915]) );
  AN2D0 U2392 ( .A1(a[8]), .A2(n[912]), .Z(n[1424]) );
  AN2D0 U2393 ( .A1(b[7]), .A2(n[401]), .Z(n[912]) );
  AN2D0 U2394 ( .A1(a[8]), .A2(n[911]), .Z(n[1423]) );
  AN2D0 U2395 ( .A1(b[7]), .A2(n[400]), .Z(n[911]) );
  AN2D0 U2396 ( .A1(a[8]), .A2(n[908]), .Z(n[1420]) );
  AN2D0 U2397 ( .A1(b[7]), .A2(n[397]), .Z(n[908]) );
  AN2D0 U2398 ( .A1(a[8]), .A2(n[905]), .Z(n[1417]) );
  AN2D0 U2399 ( .A1(b[7]), .A2(n[394]), .Z(n[905]) );
  AN2D0 U2400 ( .A1(a[8]), .A2(n[904]), .Z(n[1416]) );
  AN2D0 U2401 ( .A1(b[7]), .A2(n[393]), .Z(n[904]) );
  AN2D0 U2402 ( .A1(a[8]), .A2(n[903]), .Z(n[1415]) );
  AN2D0 U2403 ( .A1(b[7]), .A2(n[392]), .Z(n[903]) );
  AN2D0 U2404 ( .A1(a[8]), .A2(n[900]), .Z(n[1412]) );
  AN2D0 U2405 ( .A1(b[7]), .A2(n[389]), .Z(n[900]) );
  AN2D0 U2406 ( .A1(a[8]), .A2(n[897]), .Z(n[1409]) );
  AN2D0 U2407 ( .A1(b[7]), .A2(n[386]), .Z(n[897]) );
  AN2D0 U2408 ( .A1(a[8]), .A2(n[896]), .Z(n[1408]) );
  AN2D0 U2409 ( .A1(b[7]), .A2(n[385]), .Z(n[896]) );
  AN2D0 U2410 ( .A1(a[8]), .A2(n[893]), .Z(n[1405]) );
  AN2D0 U2411 ( .A1(b[7]), .A2(n[382]), .Z(n[893]) );
  AN2D0 U2412 ( .A1(a[8]), .A2(n[890]), .Z(n[1402]) );
  AN2D0 U2413 ( .A1(b[7]), .A2(n[379]), .Z(n[890]) );
  AN2D0 U2414 ( .A1(a[8]), .A2(n[889]), .Z(n[1401]) );
  AN2D0 U2415 ( .A1(b[7]), .A2(n[378]), .Z(n[889]) );
  AN2D0 U2416 ( .A1(a[8]), .A2(n[888]), .Z(n[1400]) );
  AN2D0 U2417 ( .A1(b[7]), .A2(n[377]), .Z(n[888]) );
  AN2D0 U2418 ( .A1(a[8]), .A2(n[887]), .Z(n[1399]) );
  AN2D0 U2419 ( .A1(b[7]), .A2(n[376]), .Z(n[887]) );
  AN2D0 U2420 ( .A1(a[8]), .A2(n[886]), .Z(n[1398]) );
  AN2D0 U2421 ( .A1(b[7]), .A2(n[375]), .Z(n[886]) );
  AN2D0 U2422 ( .A1(a[8]), .A2(n[885]), .Z(n[1397]) );
  AN2D0 U2423 ( .A1(b[7]), .A2(n[374]), .Z(n[885]) );
  AN2D0 U2424 ( .A1(a[8]), .A2(n[882]), .Z(n[1394]) );
  AN2D0 U2425 ( .A1(b[7]), .A2(n[371]), .Z(n[882]) );
  AN2D0 U2426 ( .A1(a[8]), .A2(n[879]), .Z(n[1391]) );
  AN2D0 U2427 ( .A1(b[7]), .A2(n[368]), .Z(n[879]) );
  AN2D0 U2428 ( .A1(a[8]), .A2(n[878]), .Z(n[1390]) );
  AN2D0 U2429 ( .A1(b[7]), .A2(n[367]), .Z(n[878]) );
  AN2D0 U2430 ( .A1(a[8]), .A2(n[875]), .Z(n[1387]) );
  AN2D0 U2431 ( .A1(b[7]), .A2(n[364]), .Z(n[875]) );
  AN2D0 U2432 ( .A1(a[8]), .A2(n[872]), .Z(n[1384]) );
  AN2D0 U2433 ( .A1(b[7]), .A2(n[361]), .Z(n[872]) );
  AN2D0 U2434 ( .A1(a[8]), .A2(n[871]), .Z(n[1383]) );
  AN2D0 U2435 ( .A1(b[7]), .A2(n[360]), .Z(n[871]) );
  AN2D0 U2436 ( .A1(a[8]), .A2(n[870]), .Z(n[1382]) );
  AN2D0 U2437 ( .A1(b[7]), .A2(n[359]), .Z(n[870]) );
  AN2D0 U2438 ( .A1(a[8]), .A2(n[867]), .Z(n[1379]) );
  AN2D0 U2439 ( .A1(b[7]), .A2(n[356]), .Z(n[867]) );
  AN2D0 U2440 ( .A1(a[8]), .A2(n[864]), .Z(n[1376]) );
  AN2D0 U2441 ( .A1(b[7]), .A2(n[353]), .Z(n[864]) );
  AN2D0 U2442 ( .A1(a[8]), .A2(n[863]), .Z(n[1375]) );
  AN2D0 U2443 ( .A1(b[7]), .A2(n[352]), .Z(n[863]) );
  AN2D0 U2444 ( .A1(a[8]), .A2(n[860]), .Z(n[1372]) );
  AN2D0 U2445 ( .A1(b[7]), .A2(n[349]), .Z(n[860]) );
  AN2D0 U2446 ( .A1(a[8]), .A2(n[857]), .Z(n[1369]) );
  AN2D0 U2447 ( .A1(b[7]), .A2(n[346]), .Z(n[857]) );
  AN2D0 U2448 ( .A1(a[8]), .A2(n[856]), .Z(n[1368]) );
  AN2D0 U2449 ( .A1(b[7]), .A2(n[345]), .Z(n[856]) );
  AN2D0 U2450 ( .A1(a[8]), .A2(n[855]), .Z(n[1367]) );
  AN2D0 U2451 ( .A1(b[7]), .A2(n[344]), .Z(n[855]) );
  AN2D0 U2452 ( .A1(a[8]), .A2(n[854]), .Z(n[1366]) );
  AN2D0 U2453 ( .A1(b[7]), .A2(n[343]), .Z(n[854]) );
  AN2D0 U2454 ( .A1(a[8]), .A2(n[851]), .Z(n[1363]) );
  AN2D0 U2455 ( .A1(b[7]), .A2(n[340]), .Z(n[851]) );
  AN2D0 U2456 ( .A1(a[8]), .A2(n[848]), .Z(n[1360]) );
  AN2D0 U2457 ( .A1(b[7]), .A2(n[337]), .Z(n[848]) );
  AN2D0 U2458 ( .A1(a[8]), .A2(n[847]), .Z(n[1359]) );
  AN2D0 U2459 ( .A1(b[7]), .A2(n[336]), .Z(n[847]) );
  AN2D0 U2460 ( .A1(a[8]), .A2(n[844]), .Z(n[1356]) );
  AN2D0 U2461 ( .A1(b[7]), .A2(n[333]), .Z(n[844]) );
  AN2D0 U2462 ( .A1(a[8]), .A2(n[841]), .Z(n[1353]) );
  AN2D0 U2463 ( .A1(b[7]), .A2(n[330]), .Z(n[841]) );
  AN2D0 U2464 ( .A1(a[8]), .A2(n[840]), .Z(n[1352]) );
  AN2D0 U2465 ( .A1(b[7]), .A2(n[329]), .Z(n[840]) );
  AN2D0 U2466 ( .A1(a[8]), .A2(n[839]), .Z(n[1351]) );
  AN2D0 U2467 ( .A1(b[7]), .A2(n[328]), .Z(n[839]) );
  AN2D0 U2468 ( .A1(a[8]), .A2(n[836]), .Z(n[1348]) );
  AN2D0 U2469 ( .A1(b[7]), .A2(n[325]), .Z(n[836]) );
  AN2D0 U2470 ( .A1(a[8]), .A2(n[833]), .Z(n[1345]) );
  AN2D0 U2471 ( .A1(b[7]), .A2(n[322]), .Z(n[833]) );
  AN2D0 U2472 ( .A1(a[8]), .A2(n[832]), .Z(n[1344]) );
  AN2D0 U2473 ( .A1(b[7]), .A2(n[321]), .Z(n[832]) );
  AN2D0 U2474 ( .A1(a[8]), .A2(n[829]), .Z(n[1341]) );
  AN2D0 U2475 ( .A1(b[7]), .A2(n[318]), .Z(n[829]) );
  AN2D0 U2476 ( .A1(a[8]), .A2(n[826]), .Z(n[1338]) );
  AN2D0 U2477 ( .A1(b[7]), .A2(n[315]), .Z(n[826]) );
  AN2D0 U2478 ( .A1(a[8]), .A2(n[825]), .Z(n[1337]) );
  AN2D0 U2479 ( .A1(b[7]), .A2(n[314]), .Z(n[825]) );
  AN2D0 U2480 ( .A1(a[8]), .A2(n[824]), .Z(n[1336]) );
  AN2D0 U2481 ( .A1(b[7]), .A2(n[313]), .Z(n[824]) );
  AN2D0 U2482 ( .A1(a[8]), .A2(n[823]), .Z(n[1335]) );
  AN2D0 U2483 ( .A1(b[7]), .A2(n[312]), .Z(n[823]) );
  AN2D0 U2484 ( .A1(a[8]), .A2(n[822]), .Z(n[1334]) );
  AN2D0 U2485 ( .A1(b[7]), .A2(n[311]), .Z(n[822]) );
  AN2D0 U2486 ( .A1(a[8]), .A2(n[819]), .Z(n[1331]) );
  AN2D0 U2487 ( .A1(b[7]), .A2(n[308]), .Z(n[819]) );
  AN2D0 U2488 ( .A1(a[8]), .A2(n[816]), .Z(n[1328]) );
  AN2D0 U2489 ( .A1(b[7]), .A2(n[305]), .Z(n[816]) );
  AN2D0 U2490 ( .A1(a[8]), .A2(n[815]), .Z(n[1327]) );
  AN2D0 U2491 ( .A1(b[7]), .A2(n[304]), .Z(n[815]) );
  AN2D0 U2492 ( .A1(a[8]), .A2(n[812]), .Z(n[1324]) );
  AN2D0 U2493 ( .A1(b[7]), .A2(n[301]), .Z(n[812]) );
  AN2D0 U2494 ( .A1(a[8]), .A2(n[809]), .Z(n[1321]) );
  AN2D0 U2495 ( .A1(b[7]), .A2(n[298]), .Z(n[809]) );
  AN2D0 U2496 ( .A1(a[8]), .A2(n[808]), .Z(n[1320]) );
  AN2D0 U2497 ( .A1(b[7]), .A2(n[297]), .Z(n[808]) );
  AN2D0 U2498 ( .A1(a[8]), .A2(n[807]), .Z(n[1319]) );
  AN2D0 U2499 ( .A1(b[7]), .A2(n[296]), .Z(n[807]) );
  AN2D0 U2500 ( .A1(a[8]), .A2(n[804]), .Z(n[1316]) );
  AN2D0 U2501 ( .A1(b[7]), .A2(n[293]), .Z(n[804]) );
  AN2D0 U2502 ( .A1(a[8]), .A2(n[801]), .Z(n[1313]) );
  AN2D0 U2503 ( .A1(b[7]), .A2(n[290]), .Z(n[801]) );
  AN2D0 U2504 ( .A1(a[8]), .A2(n[800]), .Z(n[1312]) );
  AN2D0 U2505 ( .A1(b[7]), .A2(n[289]), .Z(n[800]) );
  AN2D0 U2506 ( .A1(a[8]), .A2(n[797]), .Z(n[1309]) );
  AN2D0 U2507 ( .A1(b[7]), .A2(n[286]), .Z(n[797]) );
  AN2D0 U2508 ( .A1(a[8]), .A2(n[794]), .Z(n[1306]) );
  AN2D0 U2509 ( .A1(b[7]), .A2(n[283]), .Z(n[794]) );
  AN2D0 U2510 ( .A1(a[8]), .A2(n[793]), .Z(n[1305]) );
  AN2D0 U2511 ( .A1(b[7]), .A2(n[282]), .Z(n[793]) );
  AN2D0 U2512 ( .A1(a[8]), .A2(n[792]), .Z(n[1304]) );
  AN2D0 U2513 ( .A1(b[7]), .A2(n[281]), .Z(n[792]) );
  AN2D0 U2514 ( .A1(a[8]), .A2(n[791]), .Z(n[1303]) );
  AN2D0 U2515 ( .A1(b[7]), .A2(n[280]), .Z(n[791]) );
  AN2D0 U2516 ( .A1(a[8]), .A2(n[788]), .Z(n[1300]) );
  AN2D0 U2517 ( .A1(b[7]), .A2(n[277]), .Z(n[788]) );
  AN2D0 U2518 ( .A1(a[8]), .A2(n[785]), .Z(n[1297]) );
  AN2D0 U2519 ( .A1(b[7]), .A2(n[274]), .Z(n[785]) );
  AN2D0 U2520 ( .A1(a[8]), .A2(n[784]), .Z(n[1296]) );
  AN2D0 U2521 ( .A1(b[7]), .A2(n[273]), .Z(n[784]) );
  AN2D0 U2522 ( .A1(a[8]), .A2(n[781]), .Z(n[1293]) );
  AN2D0 U2523 ( .A1(b[7]), .A2(n[270]), .Z(n[781]) );
  AN2D0 U2524 ( .A1(a[8]), .A2(n[778]), .Z(n[1290]) );
  AN2D0 U2525 ( .A1(b[7]), .A2(n[267]), .Z(n[778]) );
  AN2D0 U2526 ( .A1(a[8]), .A2(n[777]), .Z(n[1289]) );
  AN2D0 U2527 ( .A1(b[7]), .A2(n[266]), .Z(n[777]) );
  AN2D0 U2528 ( .A1(a[8]), .A2(n[776]), .Z(n[1288]) );
  AN2D0 U2529 ( .A1(b[7]), .A2(n[265]), .Z(n[776]) );
  AN2D0 U2530 ( .A1(a[8]), .A2(n[773]), .Z(n[1285]) );
  AN2D0 U2531 ( .A1(b[7]), .A2(n[262]), .Z(n[773]) );
  AN2D0 U2532 ( .A1(a[8]), .A2(n[770]), .Z(n[1282]) );
  AN2D0 U2533 ( .A1(b[7]), .A2(n[259]), .Z(n[770]) );
  AN2D0 U2534 ( .A1(a[8]), .A2(n[769]), .Z(n[1281]) );
  AN2D0 U2535 ( .A1(b[7]), .A2(n[258]), .Z(n[769]) );
  AN2D0 U2536 ( .A1(a[8]), .A2(n[766]), .Z(n[1278]) );
  AN2D0 U2537 ( .A1(b[7]), .A2(n[255]), .Z(n[766]) );
  AN2D0 U2538 ( .A1(a[8]), .A2(n[763]), .Z(n[1275]) );
  AN2D0 U2539 ( .A1(b[7]), .A2(n[252]), .Z(n[763]) );
  AN2D0 U2540 ( .A1(a[8]), .A2(n[762]), .Z(n[1274]) );
  AN2D0 U2541 ( .A1(b[7]), .A2(n[251]), .Z(n[762]) );
  AN2D0 U2542 ( .A1(a[8]), .A2(n[761]), .Z(n[1273]) );
  AN2D0 U2543 ( .A1(b[7]), .A2(n[250]), .Z(n[761]) );
  AN2D0 U2544 ( .A1(a[8]), .A2(n[760]), .Z(n[1272]) );
  AN2D0 U2545 ( .A1(b[7]), .A2(n[249]), .Z(n[760]) );
  AN2D0 U2546 ( .A1(a[8]), .A2(n[759]), .Z(n[1271]) );
  AN2D0 U2547 ( .A1(b[7]), .A2(n[248]), .Z(n[759]) );
  AN2D0 U2548 ( .A1(a[8]), .A2(n[758]), .Z(n[1270]) );
  AN2D0 U2549 ( .A1(b[7]), .A2(n[247]), .Z(n[758]) );
  AN2D0 U2550 ( .A1(a[8]), .A2(n[757]), .Z(n[1269]) );
  AN2D0 U2551 ( .A1(b[7]), .A2(n[246]), .Z(n[757]) );
  AN2D0 U2552 ( .A1(a[8]), .A2(n[754]), .Z(n[1266]) );
  AN2D0 U2553 ( .A1(n[498]), .A2(a[7]), .Z(n[754]) );
  AN2D0 U2554 ( .A1(a[8]), .A2(n[751]), .Z(n[1263]) );
  AN2D0 U2555 ( .A1(a[7]), .A2(n[495]), .Z(n[751]) );
  AN2D0 U2556 ( .A1(a[8]), .A2(n[750]), .Z(n[1262]) );
  AN2D0 U2557 ( .A1(a[7]), .A2(n[494]), .Z(n[750]) );
  AN2D0 U2558 ( .A1(a[8]), .A2(n[747]), .Z(n[1259]) );
  AN2D0 U2559 ( .A1(a[7]), .A2(n[491]), .Z(n[747]) );
  AN2D0 U2560 ( .A1(a[8]), .A2(n[744]), .Z(n[1256]) );
  AN2D0 U2561 ( .A1(n[488]), .A2(a[7]), .Z(n[744]) );
  AN2D0 U2562 ( .A1(n[233]), .A2(b[6]), .Z(n[488]) );
  AN2D0 U2563 ( .A1(a[8]), .A2(n[743]), .Z(n[1255]) );
  AN2D0 U2564 ( .A1(n[487]), .A2(a[7]), .Z(n[743]) );
  AN2D0 U2565 ( .A1(b[6]), .A2(n[232]), .Z(n[487]) );
  AN2D0 U2566 ( .A1(a[8]), .A2(n[742]), .Z(n[1254]) );
  AN2D0 U2567 ( .A1(n[486]), .A2(a[7]), .Z(n[742]) );
  AN2D0 U2568 ( .A1(b[6]), .A2(n[231]), .Z(n[486]) );
  AN2D0 U2569 ( .A1(a[8]), .A2(n[739]), .Z(n[1251]) );
  AN2D0 U2570 ( .A1(n[483]), .A2(a[7]), .Z(n[739]) );
  AN2D0 U2571 ( .A1(b[6]), .A2(n[228]), .Z(n[483]) );
  AN2D0 U2572 ( .A1(a[8]), .A2(n[736]), .Z(n[1248]) );
  AN2D0 U2573 ( .A1(n[480]), .A2(a[7]), .Z(n[736]) );
  AN2D0 U2574 ( .A1(b[6]), .A2(n[225]), .Z(n[480]) );
  AN2D0 U2575 ( .A1(a[8]), .A2(n[735]), .Z(n[1247]) );
  AN2D0 U2576 ( .A1(n[479]), .A2(a[7]), .Z(n[735]) );
  AN2D0 U2577 ( .A1(b[6]), .A2(n[224]), .Z(n[479]) );
  AN2D0 U2578 ( .A1(a[8]), .A2(n[732]), .Z(n[1244]) );
  AN2D0 U2579 ( .A1(n[476]), .A2(a[7]), .Z(n[732]) );
  AN2D0 U2580 ( .A1(b[6]), .A2(n[221]), .Z(n[476]) );
  AN2D0 U2581 ( .A1(a[8]), .A2(n[729]), .Z(n[1241]) );
  AN2D0 U2582 ( .A1(n[473]), .A2(a[7]), .Z(n[729]) );
  AN2D0 U2583 ( .A1(b[6]), .A2(n[218]), .Z(n[473]) );
  AN2D0 U2584 ( .A1(a[8]), .A2(n[728]), .Z(n[1240]) );
  AN2D0 U2585 ( .A1(n[472]), .A2(a[7]), .Z(n[728]) );
  AN2D0 U2586 ( .A1(b[6]), .A2(n[217]), .Z(n[472]) );
  AN2D0 U2587 ( .A1(a[8]), .A2(n[727]), .Z(n[1239]) );
  AN2D0 U2588 ( .A1(n[471]), .A2(a[7]), .Z(n[727]) );
  AN2D0 U2589 ( .A1(b[6]), .A2(n[216]), .Z(n[471]) );
  AN2D0 U2590 ( .A1(a[8]), .A2(n[726]), .Z(n[1238]) );
  AN2D0 U2591 ( .A1(n[470]), .A2(a[7]), .Z(n[726]) );
  AN2D0 U2592 ( .A1(b[6]), .A2(n[215]), .Z(n[470]) );
  AN2D0 U2593 ( .A1(a[8]), .A2(n[723]), .Z(n[1235]) );
  AN2D0 U2594 ( .A1(n[467]), .A2(a[7]), .Z(n[723]) );
  AN2D0 U2595 ( .A1(b[6]), .A2(n[212]), .Z(n[467]) );
  AN2D0 U2596 ( .A1(a[8]), .A2(n[720]), .Z(n[1232]) );
  AN2D0 U2597 ( .A1(n[464]), .A2(a[7]), .Z(n[720]) );
  AN2D0 U2598 ( .A1(b[6]), .A2(n[209]), .Z(n[464]) );
  AN2D0 U2599 ( .A1(a[8]), .A2(n[719]), .Z(n[1231]) );
  AN2D0 U2600 ( .A1(n[463]), .A2(a[7]), .Z(n[719]) );
  AN2D0 U2601 ( .A1(b[6]), .A2(n[208]), .Z(n[463]) );
  AN2D0 U2602 ( .A1(a[8]), .A2(n[716]), .Z(n[1228]) );
  AN2D0 U2603 ( .A1(n[460]), .A2(a[7]), .Z(n[716]) );
  AN2D0 U2604 ( .A1(b[6]), .A2(n[205]), .Z(n[460]) );
  AN2D0 U2605 ( .A1(a[8]), .A2(n[713]), .Z(n[1225]) );
  AN2D0 U2606 ( .A1(n[457]), .A2(a[7]), .Z(n[713]) );
  AN2D0 U2607 ( .A1(b[6]), .A2(n[202]), .Z(n[457]) );
  AN2D0 U2608 ( .A1(a[8]), .A2(n[712]), .Z(n[1224]) );
  AN2D0 U2609 ( .A1(n[456]), .A2(a[7]), .Z(n[712]) );
  AN2D0 U2610 ( .A1(b[6]), .A2(n[201]), .Z(n[456]) );
  AN2D0 U2611 ( .A1(a[8]), .A2(n[711]), .Z(n[1223]) );
  AN2D0 U2612 ( .A1(n[455]), .A2(a[7]), .Z(n[711]) );
  AN2D0 U2613 ( .A1(b[6]), .A2(n[200]), .Z(n[455]) );
  AN2D0 U2614 ( .A1(a[8]), .A2(n[708]), .Z(n[1220]) );
  AN2D0 U2615 ( .A1(n[452]), .A2(a[7]), .Z(n[708]) );
  AN2D0 U2616 ( .A1(b[6]), .A2(n[197]), .Z(n[452]) );
  AN2D0 U2617 ( .A1(a[8]), .A2(n[705]), .Z(n[1217]) );
  AN2D0 U2618 ( .A1(n[449]), .A2(a[7]), .Z(n[705]) );
  AN2D0 U2619 ( .A1(b[6]), .A2(n[194]), .Z(n[449]) );
  AN2D0 U2620 ( .A1(a[8]), .A2(n[704]), .Z(n[1216]) );
  AN2D0 U2621 ( .A1(n[448]), .A2(a[7]), .Z(n[704]) );
  AN2D0 U2622 ( .A1(b[6]), .A2(n[193]), .Z(n[448]) );
  AN2D0 U2623 ( .A1(a[8]), .A2(n[701]), .Z(n[1213]) );
  AN2D0 U2624 ( .A1(n[445]), .A2(a[7]), .Z(n[701]) );
  AN2D0 U2625 ( .A1(b[6]), .A2(n[190]), .Z(n[445]) );
  AN2D0 U2626 ( .A1(a[8]), .A2(n[698]), .Z(n[1210]) );
  AN2D0 U2627 ( .A1(n[442]), .A2(a[7]), .Z(n[698]) );
  AN2D0 U2628 ( .A1(b[6]), .A2(n[187]), .Z(n[442]) );
  AN2D0 U2629 ( .A1(a[8]), .A2(n[697]), .Z(n[1209]) );
  AN2D0 U2630 ( .A1(n[441]), .A2(a[7]), .Z(n[697]) );
  AN2D0 U2631 ( .A1(b[6]), .A2(n[186]), .Z(n[441]) );
  AN2D0 U2632 ( .A1(a[8]), .A2(n[696]), .Z(n[1208]) );
  AN2D0 U2633 ( .A1(n[440]), .A2(a[7]), .Z(n[696]) );
  AN2D0 U2634 ( .A1(b[6]), .A2(n[185]), .Z(n[440]) );
  AN2D0 U2635 ( .A1(a[8]), .A2(n[695]), .Z(n[1207]) );
  AN2D0 U2636 ( .A1(n[439]), .A2(a[7]), .Z(n[695]) );
  AN2D0 U2637 ( .A1(b[6]), .A2(n[184]), .Z(n[439]) );
  AN2D0 U2638 ( .A1(a[8]), .A2(n[694]), .Z(n[1206]) );
  AN2D0 U2639 ( .A1(n[438]), .A2(a[7]), .Z(n[694]) );
  AN2D0 U2640 ( .A1(b[6]), .A2(n[183]), .Z(n[438]) );
  AN2D0 U2641 ( .A1(a[8]), .A2(n[691]), .Z(n[1203]) );
  AN2D0 U2642 ( .A1(n[435]), .A2(a[7]), .Z(n[691]) );
  AN2D0 U2643 ( .A1(b[6]), .A2(n[180]), .Z(n[435]) );
  AN2D0 U2644 ( .A1(a[8]), .A2(n[688]), .Z(n[1200]) );
  AN2D0 U2645 ( .A1(n[432]), .A2(a[7]), .Z(n[688]) );
  AN2D0 U2646 ( .A1(b[6]), .A2(n[177]), .Z(n[432]) );
  AN2D0 U2647 ( .A1(a[8]), .A2(n[687]), .Z(n[1199]) );
  AN2D0 U2648 ( .A1(n[431]), .A2(a[7]), .Z(n[687]) );
  AN2D0 U2649 ( .A1(b[6]), .A2(n[176]), .Z(n[431]) );
  AN2D0 U2650 ( .A1(a[8]), .A2(n[684]), .Z(n[1196]) );
  AN2D0 U2651 ( .A1(n[428]), .A2(a[7]), .Z(n[684]) );
  AN2D0 U2652 ( .A1(b[6]), .A2(n[173]), .Z(n[428]) );
  AN2D0 U2653 ( .A1(a[8]), .A2(n[681]), .Z(n[1193]) );
  AN2D0 U2654 ( .A1(n[425]), .A2(a[7]), .Z(n[681]) );
  AN2D0 U2655 ( .A1(b[6]), .A2(n[170]), .Z(n[425]) );
  AN2D0 U2656 ( .A1(a[8]), .A2(n[680]), .Z(n[1192]) );
  AN2D0 U2657 ( .A1(n[424]), .A2(a[7]), .Z(n[680]) );
  AN2D0 U2658 ( .A1(b[6]), .A2(n[169]), .Z(n[424]) );
  AN2D0 U2659 ( .A1(a[8]), .A2(n[679]), .Z(n[1191]) );
  AN2D0 U2660 ( .A1(n[423]), .A2(a[7]), .Z(n[679]) );
  AN2D0 U2661 ( .A1(b[6]), .A2(n[168]), .Z(n[423]) );
  AN2D0 U2662 ( .A1(a[8]), .A2(n[676]), .Z(n[1188]) );
  AN2D0 U2663 ( .A1(n[420]), .A2(a[7]), .Z(n[676]) );
  AN2D0 U2664 ( .A1(b[6]), .A2(n[165]), .Z(n[420]) );
  AN2D0 U2665 ( .A1(a[8]), .A2(n[673]), .Z(n[1185]) );
  AN2D0 U2666 ( .A1(n[417]), .A2(a[7]), .Z(n[673]) );
  AN2D0 U2667 ( .A1(b[6]), .A2(n[162]), .Z(n[417]) );
  AN2D0 U2668 ( .A1(a[8]), .A2(n[672]), .Z(n[1184]) );
  AN2D0 U2669 ( .A1(n[416]), .A2(a[7]), .Z(n[672]) );
  AN2D0 U2670 ( .A1(b[6]), .A2(n[161]), .Z(n[416]) );
  AN2D0 U2671 ( .A1(a[8]), .A2(n[669]), .Z(n[1181]) );
  AN2D0 U2672 ( .A1(n[413]), .A2(a[7]), .Z(n[669]) );
  AN2D0 U2673 ( .A1(b[6]), .A2(n[158]), .Z(n[413]) );
  AN2D0 U2674 ( .A1(a[8]), .A2(n[666]), .Z(n[1178]) );
  AN2D0 U2675 ( .A1(n[410]), .A2(a[7]), .Z(n[666]) );
  AN2D0 U2676 ( .A1(b[6]), .A2(n[155]), .Z(n[410]) );
  AN2D0 U2677 ( .A1(a[8]), .A2(n[665]), .Z(n[1177]) );
  AN2D0 U2678 ( .A1(n[409]), .A2(a[7]), .Z(n[665]) );
  AN2D0 U2679 ( .A1(b[6]), .A2(n[154]), .Z(n[409]) );
  AN2D0 U2680 ( .A1(a[8]), .A2(n[664]), .Z(n[1176]) );
  AN2D0 U2681 ( .A1(n[408]), .A2(a[7]), .Z(n[664]) );
  AN2D0 U2682 ( .A1(b[6]), .A2(n[153]), .Z(n[408]) );
  AN2D0 U2683 ( .A1(a[8]), .A2(n[663]), .Z(n[1175]) );
  AN2D0 U2684 ( .A1(n[407]), .A2(a[7]), .Z(n[663]) );
  AN2D0 U2685 ( .A1(b[6]), .A2(n[152]), .Z(n[407]) );
  AN2D0 U2686 ( .A1(a[8]), .A2(n[660]), .Z(n[1172]) );
  AN2D0 U2687 ( .A1(n[404]), .A2(a[7]), .Z(n[660]) );
  AN2D0 U2688 ( .A1(b[6]), .A2(n[149]), .Z(n[404]) );
  AN2D0 U2689 ( .A1(a[8]), .A2(n[657]), .Z(n[1169]) );
  AN2D0 U2690 ( .A1(n[401]), .A2(a[7]), .Z(n[657]) );
  AN2D0 U2691 ( .A1(b[6]), .A2(n[146]), .Z(n[401]) );
  AN2D0 U2692 ( .A1(a[8]), .A2(n[656]), .Z(n[1168]) );
  AN2D0 U2693 ( .A1(n[400]), .A2(a[7]), .Z(n[656]) );
  AN2D0 U2694 ( .A1(b[6]), .A2(n[145]), .Z(n[400]) );
  AN2D0 U2695 ( .A1(a[8]), .A2(n[653]), .Z(n[1165]) );
  AN2D0 U2696 ( .A1(n[397]), .A2(a[7]), .Z(n[653]) );
  AN2D0 U2697 ( .A1(b[6]), .A2(n[142]), .Z(n[397]) );
  AN2D0 U2698 ( .A1(a[8]), .A2(n[650]), .Z(n[1162]) );
  AN2D0 U2699 ( .A1(n[394]), .A2(a[7]), .Z(n[650]) );
  AN2D0 U2700 ( .A1(b[6]), .A2(n[139]), .Z(n[394]) );
  AN2D0 U2701 ( .A1(a[8]), .A2(n[649]), .Z(n[1161]) );
  AN2D0 U2702 ( .A1(n[393]), .A2(a[7]), .Z(n[649]) );
  AN2D0 U2703 ( .A1(b[6]), .A2(n[138]), .Z(n[393]) );
  AN2D0 U2704 ( .A1(a[8]), .A2(n[648]), .Z(n[1160]) );
  AN2D0 U2705 ( .A1(n[392]), .A2(a[7]), .Z(n[648]) );
  AN2D0 U2706 ( .A1(b[6]), .A2(n[137]), .Z(n[392]) );
  AN2D0 U2707 ( .A1(a[8]), .A2(n[645]), .Z(n[1157]) );
  AN2D0 U2708 ( .A1(n[389]), .A2(a[7]), .Z(n[645]) );
  AN2D0 U2709 ( .A1(b[6]), .A2(n[134]), .Z(n[389]) );
  AN2D0 U2710 ( .A1(a[8]), .A2(n[642]), .Z(n[1154]) );
  AN2D0 U2711 ( .A1(n[386]), .A2(a[7]), .Z(n[642]) );
  AN2D0 U2712 ( .A1(b[6]), .A2(n[131]), .Z(n[386]) );
  AN2D0 U2713 ( .A1(a[8]), .A2(n[641]), .Z(n[1153]) );
  AN2D0 U2714 ( .A1(n[385]), .A2(a[7]), .Z(n[641]) );
  AN2D0 U2715 ( .A1(b[6]), .A2(n[130]), .Z(n[385]) );
  AN2D0 U2716 ( .A1(a[8]), .A2(n[638]), .Z(n[1150]) );
  AN2D0 U2717 ( .A1(n[382]), .A2(a[7]), .Z(n[638]) );
  AN2D0 U2718 ( .A1(b[6]), .A2(n[127]), .Z(n[382]) );
  AN2D0 U2719 ( .A1(a[8]), .A2(n[635]), .Z(n[1147]) );
  AN2D0 U2720 ( .A1(n[379]), .A2(a[7]), .Z(n[635]) );
  AN2D0 U2721 ( .A1(b[6]), .A2(n[124]), .Z(n[379]) );
  AN2D0 U2722 ( .A1(a[8]), .A2(n[634]), .Z(n[1146]) );
  AN2D0 U2723 ( .A1(n[378]), .A2(a[7]), .Z(n[634]) );
  AN2D0 U2724 ( .A1(b[6]), .A2(n[123]), .Z(n[378]) );
  AN2D0 U2725 ( .A1(a[8]), .A2(n[633]), .Z(n[1145]) );
  AN2D0 U2726 ( .A1(n[377]), .A2(a[7]), .Z(n[633]) );
  AN2D0 U2727 ( .A1(b[6]), .A2(n[122]), .Z(n[377]) );
  AN2D0 U2728 ( .A1(a[8]), .A2(n[632]), .Z(n[1144]) );
  AN2D0 U2729 ( .A1(n[376]), .A2(a[7]), .Z(n[632]) );
  AN2D0 U2730 ( .A1(b[6]), .A2(n[121]), .Z(n[376]) );
  AN2D0 U2731 ( .A1(a[8]), .A2(n[631]), .Z(n[1143]) );
  AN2D0 U2732 ( .A1(n[375]), .A2(a[7]), .Z(n[631]) );
  AN2D0 U2733 ( .A1(b[6]), .A2(n[120]), .Z(n[375]) );
  AN2D0 U2734 ( .A1(a[8]), .A2(n[630]), .Z(n[1142]) );
  AN2D0 U2735 ( .A1(n[374]), .A2(a[7]), .Z(n[630]) );
  AN2D0 U2736 ( .A1(b[6]), .A2(n[119]), .Z(n[374]) );
  AN2D0 U2737 ( .A1(a[8]), .A2(n[627]), .Z(n[1139]) );
  AN2D0 U2738 ( .A1(n[371]), .A2(a[7]), .Z(n[627]) );
  AN2D0 U2739 ( .A1(n[243]), .A2(a[6]), .Z(n[371]) );
  AN2D0 U2740 ( .A1(a[8]), .A2(n[624]), .Z(n[1136]) );
  AN2D0 U2741 ( .A1(n[368]), .A2(a[7]), .Z(n[624]) );
  AN2D0 U2742 ( .A1(a[6]), .A2(n[240]), .Z(n[368]) );
  AN2D0 U2743 ( .A1(a[8]), .A2(n[623]), .Z(n[1135]) );
  AN2D0 U2744 ( .A1(n[367]), .A2(a[7]), .Z(n[623]) );
  AN2D0 U2745 ( .A1(a[6]), .A2(n[239]), .Z(n[367]) );
  AN2D0 U2746 ( .A1(a[8]), .A2(n[620]), .Z(n[1132]) );
  AN2D0 U2747 ( .A1(n[364]), .A2(a[7]), .Z(n[620]) );
  AN2D0 U2748 ( .A1(a[6]), .A2(n[236]), .Z(n[364]) );
  AN2D0 U2749 ( .A1(a[8]), .A2(n[617]), .Z(n[1129]) );
  AN2D0 U2750 ( .A1(n[361]), .A2(a[7]), .Z(n[617]) );
  AN2D0 U2751 ( .A1(n[233]), .A2(a[6]), .Z(n[361]) );
  AN2D0 U2752 ( .A1(n[106]), .A2(b[5]), .Z(n[233]) );
  AN2D0 U2753 ( .A1(a[8]), .A2(n[616]), .Z(n[1128]) );
  AN2D0 U2754 ( .A1(n[360]), .A2(a[7]), .Z(n[616]) );
  AN2D0 U2755 ( .A1(n[232]), .A2(a[6]), .Z(n[360]) );
  AN2D0 U2756 ( .A1(b[5]), .A2(n[105]), .Z(n[232]) );
  AN2D0 U2757 ( .A1(a[8]), .A2(n[615]), .Z(n[1127]) );
  AN2D0 U2758 ( .A1(n[359]), .A2(a[7]), .Z(n[615]) );
  AN2D0 U2759 ( .A1(n[231]), .A2(a[6]), .Z(n[359]) );
  AN2D0 U2760 ( .A1(b[5]), .A2(n[104]), .Z(n[231]) );
  AN2D0 U2761 ( .A1(a[8]), .A2(n[612]), .Z(n[1124]) );
  AN2D0 U2762 ( .A1(n[356]), .A2(a[7]), .Z(n[612]) );
  AN2D0 U2763 ( .A1(n[228]), .A2(a[6]), .Z(n[356]) );
  AN2D0 U2764 ( .A1(b[5]), .A2(n[101]), .Z(n[228]) );
  AN2D0 U2765 ( .A1(a[8]), .A2(n[609]), .Z(n[1121]) );
  AN2D0 U2766 ( .A1(n[353]), .A2(a[7]), .Z(n[609]) );
  AN2D0 U2767 ( .A1(n[225]), .A2(a[6]), .Z(n[353]) );
  AN2D0 U2768 ( .A1(b[5]), .A2(n[98]), .Z(n[225]) );
  AN2D0 U2769 ( .A1(a[8]), .A2(n[608]), .Z(n[1120]) );
  AN2D0 U2770 ( .A1(n[352]), .A2(a[7]), .Z(n[608]) );
  AN2D0 U2771 ( .A1(n[224]), .A2(a[6]), .Z(n[352]) );
  AN2D0 U2772 ( .A1(b[5]), .A2(n[97]), .Z(n[224]) );
  AN2D0 U2773 ( .A1(a[8]), .A2(n[605]), .Z(n[1117]) );
  AN2D0 U2774 ( .A1(n[349]), .A2(a[7]), .Z(n[605]) );
  AN2D0 U2775 ( .A1(n[221]), .A2(a[6]), .Z(n[349]) );
  AN2D0 U2776 ( .A1(b[5]), .A2(n[94]), .Z(n[221]) );
  AN2D0 U2777 ( .A1(a[8]), .A2(n[602]), .Z(n[1114]) );
  AN2D0 U2778 ( .A1(n[346]), .A2(a[7]), .Z(n[602]) );
  AN2D0 U2779 ( .A1(n[218]), .A2(a[6]), .Z(n[346]) );
  AN2D0 U2780 ( .A1(b[5]), .A2(n[91]), .Z(n[218]) );
  AN2D0 U2781 ( .A1(a[8]), .A2(n[601]), .Z(n[1113]) );
  AN2D0 U2782 ( .A1(n[345]), .A2(a[7]), .Z(n[601]) );
  AN2D0 U2783 ( .A1(n[217]), .A2(a[6]), .Z(n[345]) );
  AN2D0 U2784 ( .A1(b[5]), .A2(n[90]), .Z(n[217]) );
  AN2D0 U2785 ( .A1(a[8]), .A2(n[600]), .Z(n[1112]) );
  AN2D0 U2786 ( .A1(n[344]), .A2(a[7]), .Z(n[600]) );
  AN2D0 U2787 ( .A1(n[216]), .A2(a[6]), .Z(n[344]) );
  AN2D0 U2788 ( .A1(b[5]), .A2(n[89]), .Z(n[216]) );
  AN2D0 U2789 ( .A1(a[8]), .A2(n[599]), .Z(n[1111]) );
  AN2D0 U2790 ( .A1(n[343]), .A2(a[7]), .Z(n[599]) );
  AN2D0 U2791 ( .A1(n[215]), .A2(a[6]), .Z(n[343]) );
  AN2D0 U2792 ( .A1(b[5]), .A2(n[88]), .Z(n[215]) );
  AN2D0 U2793 ( .A1(a[8]), .A2(n[596]), .Z(n[1108]) );
  AN2D0 U2794 ( .A1(n[340]), .A2(a[7]), .Z(n[596]) );
  AN2D0 U2795 ( .A1(n[212]), .A2(a[6]), .Z(n[340]) );
  AN2D0 U2796 ( .A1(b[5]), .A2(n[85]), .Z(n[212]) );
  AN2D0 U2797 ( .A1(a[8]), .A2(n[593]), .Z(n[1105]) );
  AN2D0 U2798 ( .A1(n[337]), .A2(a[7]), .Z(n[593]) );
  AN2D0 U2799 ( .A1(n[209]), .A2(a[6]), .Z(n[337]) );
  AN2D0 U2800 ( .A1(b[5]), .A2(n[82]), .Z(n[209]) );
  AN2D0 U2801 ( .A1(a[8]), .A2(n[592]), .Z(n[1104]) );
  AN2D0 U2802 ( .A1(n[336]), .A2(a[7]), .Z(n[592]) );
  AN2D0 U2803 ( .A1(n[208]), .A2(a[6]), .Z(n[336]) );
  AN2D0 U2804 ( .A1(b[5]), .A2(n[81]), .Z(n[208]) );
  AN2D0 U2805 ( .A1(a[8]), .A2(n[589]), .Z(n[1101]) );
  AN2D0 U2806 ( .A1(n[333]), .A2(a[7]), .Z(n[589]) );
  AN2D0 U2807 ( .A1(n[205]), .A2(a[6]), .Z(n[333]) );
  AN2D0 U2808 ( .A1(b[5]), .A2(n[78]), .Z(n[205]) );
  AN2D0 U2809 ( .A1(a[8]), .A2(n[586]), .Z(n[1098]) );
  AN2D0 U2810 ( .A1(n[330]), .A2(a[7]), .Z(n[586]) );
  AN2D0 U2811 ( .A1(n[202]), .A2(a[6]), .Z(n[330]) );
  AN2D0 U2812 ( .A1(b[5]), .A2(n[75]), .Z(n[202]) );
  AN2D0 U2813 ( .A1(a[8]), .A2(n[585]), .Z(n[1097]) );
  AN2D0 U2814 ( .A1(n[329]), .A2(a[7]), .Z(n[585]) );
  AN2D0 U2815 ( .A1(n[201]), .A2(a[6]), .Z(n[329]) );
  AN2D0 U2816 ( .A1(b[5]), .A2(n[74]), .Z(n[201]) );
  AN2D0 U2817 ( .A1(a[8]), .A2(n[584]), .Z(n[1096]) );
  AN2D0 U2818 ( .A1(n[328]), .A2(a[7]), .Z(n[584]) );
  AN2D0 U2819 ( .A1(n[200]), .A2(a[6]), .Z(n[328]) );
  AN2D0 U2820 ( .A1(b[5]), .A2(n[73]), .Z(n[200]) );
  AN2D0 U2821 ( .A1(a[8]), .A2(n[581]), .Z(n[1093]) );
  AN2D0 U2822 ( .A1(n[325]), .A2(a[7]), .Z(n[581]) );
  AN2D0 U2823 ( .A1(n[197]), .A2(a[6]), .Z(n[325]) );
  AN2D0 U2824 ( .A1(b[5]), .A2(n[70]), .Z(n[197]) );
  AN2D0 U2825 ( .A1(a[8]), .A2(n[578]), .Z(n[1090]) );
  AN2D0 U2826 ( .A1(n[322]), .A2(a[7]), .Z(n[578]) );
  AN2D0 U2827 ( .A1(n[194]), .A2(a[6]), .Z(n[322]) );
  AN2D0 U2828 ( .A1(b[5]), .A2(n[67]), .Z(n[194]) );
  AN2D0 U2829 ( .A1(a[8]), .A2(n[577]), .Z(n[1089]) );
  AN2D0 U2830 ( .A1(n[321]), .A2(a[7]), .Z(n[577]) );
  AN2D0 U2831 ( .A1(n[193]), .A2(a[6]), .Z(n[321]) );
  AN2D0 U2832 ( .A1(b[5]), .A2(n[66]), .Z(n[193]) );
  AN2D0 U2833 ( .A1(a[8]), .A2(n[574]), .Z(n[1086]) );
  AN2D0 U2834 ( .A1(n[318]), .A2(a[7]), .Z(n[574]) );
  AN2D0 U2835 ( .A1(n[190]), .A2(a[6]), .Z(n[318]) );
  AN2D0 U2836 ( .A1(b[5]), .A2(n[63]), .Z(n[190]) );
  AN2D0 U2837 ( .A1(a[8]), .A2(n[571]), .Z(n[1083]) );
  AN2D0 U2838 ( .A1(n[315]), .A2(a[7]), .Z(n[571]) );
  AN2D0 U2839 ( .A1(n[187]), .A2(a[6]), .Z(n[315]) );
  AN2D0 U2840 ( .A1(b[5]), .A2(n[60]), .Z(n[187]) );
  AN2D0 U2841 ( .A1(a[8]), .A2(n[570]), .Z(n[1082]) );
  AN2D0 U2842 ( .A1(n[314]), .A2(a[7]), .Z(n[570]) );
  AN2D0 U2843 ( .A1(n[186]), .A2(a[6]), .Z(n[314]) );
  AN2D0 U2844 ( .A1(b[5]), .A2(n[59]), .Z(n[186]) );
  AN2D0 U2845 ( .A1(a[8]), .A2(n[569]), .Z(n[1081]) );
  AN2D0 U2846 ( .A1(n[313]), .A2(a[7]), .Z(n[569]) );
  AN2D0 U2847 ( .A1(n[185]), .A2(a[6]), .Z(n[313]) );
  AN2D0 U2848 ( .A1(b[5]), .A2(n[58]), .Z(n[185]) );
  AN2D0 U2849 ( .A1(a[8]), .A2(n[568]), .Z(n[1080]) );
  AN2D0 U2850 ( .A1(n[312]), .A2(a[7]), .Z(n[568]) );
  AN2D0 U2851 ( .A1(n[184]), .A2(a[6]), .Z(n[312]) );
  AN2D0 U2852 ( .A1(b[5]), .A2(n[57]), .Z(n[184]) );
  AN2D0 U2853 ( .A1(a[8]), .A2(n[567]), .Z(n[1079]) );
  AN2D0 U2854 ( .A1(n[311]), .A2(a[7]), .Z(n[567]) );
  AN2D0 U2855 ( .A1(n[183]), .A2(a[6]), .Z(n[311]) );
  AN2D0 U2856 ( .A1(b[5]), .A2(n[56]), .Z(n[183]) );
  AN2D0 U2857 ( .A1(a[8]), .A2(n[564]), .Z(n[1076]) );
  AN2D0 U2858 ( .A1(n[308]), .A2(a[7]), .Z(n[564]) );
  AN2D0 U2859 ( .A1(n[180]), .A2(a[6]), .Z(n[308]) );
  AN2D0 U2860 ( .A1(n[116]), .A2(a[5]), .Z(n[180]) );
  AN2D0 U2861 ( .A1(a[8]), .A2(n[561]), .Z(n[1073]) );
  AN2D0 U2862 ( .A1(n[305]), .A2(a[7]), .Z(n[561]) );
  AN2D0 U2863 ( .A1(n[177]), .A2(a[6]), .Z(n[305]) );
  AN2D0 U2864 ( .A1(a[5]), .A2(n[113]), .Z(n[177]) );
  AN2D0 U2865 ( .A1(a[8]), .A2(n[560]), .Z(n[1072]) );
  AN2D0 U2866 ( .A1(n[304]), .A2(a[7]), .Z(n[560]) );
  AN2D0 U2867 ( .A1(n[176]), .A2(a[6]), .Z(n[304]) );
  AN2D0 U2868 ( .A1(a[5]), .A2(n[112]), .Z(n[176]) );
  AN2D0 U2869 ( .A1(a[8]), .A2(n[557]), .Z(n[1069]) );
  AN2D0 U2870 ( .A1(n[301]), .A2(a[7]), .Z(n[557]) );
  AN2D0 U2871 ( .A1(n[173]), .A2(a[6]), .Z(n[301]) );
  AN2D0 U2872 ( .A1(a[5]), .A2(n[109]), .Z(n[173]) );
  AN2D0 U2873 ( .A1(a[8]), .A2(n[554]), .Z(n[1066]) );
  AN2D0 U2874 ( .A1(n[298]), .A2(a[7]), .Z(n[554]) );
  AN2D0 U2875 ( .A1(n[170]), .A2(a[6]), .Z(n[298]) );
  AN2D0 U2876 ( .A1(n[106]), .A2(a[5]), .Z(n[170]) );
  AN2D0 U2877 ( .A1(n[43]), .A2(b[4]), .Z(n[106]) );
  AN2D0 U2878 ( .A1(a[8]), .A2(n[553]), .Z(n[1065]) );
  AN2D0 U2879 ( .A1(n[297]), .A2(a[7]), .Z(n[553]) );
  AN2D0 U2880 ( .A1(n[169]), .A2(a[6]), .Z(n[297]) );
  AN2D0 U2881 ( .A1(n[105]), .A2(a[5]), .Z(n[169]) );
  AN2D0 U2882 ( .A1(a[8]), .A2(n[552]), .Z(n[1064]) );
  AN2D0 U2883 ( .A1(n[296]), .A2(a[7]), .Z(n[552]) );
  AN2D0 U2884 ( .A1(n[168]), .A2(a[6]), .Z(n[296]) );
  AN2D0 U2885 ( .A1(n[104]), .A2(a[5]), .Z(n[168]) );
  AN2D0 U2886 ( .A1(a[8]), .A2(n[549]), .Z(n[1061]) );
  AN2D0 U2887 ( .A1(n[293]), .A2(a[7]), .Z(n[549]) );
  AN2D0 U2888 ( .A1(n[165]), .A2(a[6]), .Z(n[293]) );
  AN2D0 U2889 ( .A1(n[101]), .A2(a[5]), .Z(n[165]) );
  AN2D0 U2890 ( .A1(b[4]), .A2(n[42]), .Z(n[105]) );
  AN2D0 U2891 ( .A1(a[8]), .A2(n[546]), .Z(n[1058]) );
  AN2D0 U2892 ( .A1(n[290]), .A2(a[7]), .Z(n[546]) );
  AN2D0 U2893 ( .A1(n[162]), .A2(a[6]), .Z(n[290]) );
  AN2D0 U2894 ( .A1(n[98]), .A2(a[5]), .Z(n[162]) );
  AN2D0 U2895 ( .A1(b[4]), .A2(n[35]), .Z(n[98]) );
  AN2D0 U2896 ( .A1(a[8]), .A2(n[545]), .Z(n[1057]) );
  AN2D0 U2897 ( .A1(n[289]), .A2(a[7]), .Z(n[545]) );
  AN2D0 U2898 ( .A1(n[161]), .A2(a[6]), .Z(n[289]) );
  AN2D0 U2899 ( .A1(n[97]), .A2(a[5]), .Z(n[161]) );
  AN2D0 U2900 ( .A1(b[4]), .A2(n[34]), .Z(n[97]) );
  AN2D0 U2901 ( .A1(a[8]), .A2(n[542]), .Z(n[1054]) );
  AN2D0 U2902 ( .A1(n[286]), .A2(a[7]), .Z(n[542]) );
  AN2D0 U2903 ( .A1(n[158]), .A2(a[6]), .Z(n[286]) );
  AN2D0 U2904 ( .A1(n[94]), .A2(a[5]), .Z(n[158]) );
  AN2D0 U2905 ( .A1(b[4]), .A2(n[31]), .Z(n[94]) );
  AN2D0 U2906 ( .A1(a[8]), .A2(n[539]), .Z(n[1051]) );
  AN2D0 U2907 ( .A1(n[283]), .A2(a[7]), .Z(n[539]) );
  AN2D0 U2908 ( .A1(n[155]), .A2(a[6]), .Z(n[283]) );
  AN2D0 U2909 ( .A1(n[91]), .A2(a[5]), .Z(n[155]) );
  AN2D0 U2910 ( .A1(b[4]), .A2(n[28]), .Z(n[91]) );
  AN2D0 U2911 ( .A1(a[8]), .A2(n[538]), .Z(n[1050]) );
  AN2D0 U2912 ( .A1(n[282]), .A2(a[7]), .Z(n[538]) );
  AN2D0 U2913 ( .A1(n[154]), .A2(a[6]), .Z(n[282]) );
  AN2D0 U2914 ( .A1(n[90]), .A2(a[5]), .Z(n[154]) );
  AN2D0 U2915 ( .A1(b[4]), .A2(n[27]), .Z(n[90]) );
  AN2D0 U2916 ( .A1(b[4]), .A2(n[41]), .Z(n[104]) );
  AN2D0 U2917 ( .A1(a[8]), .A2(n[537]), .Z(n[1049]) );
  AN2D0 U2918 ( .A1(n[281]), .A2(a[7]), .Z(n[537]) );
  AN2D0 U2919 ( .A1(n[153]), .A2(a[6]), .Z(n[281]) );
  AN2D0 U2920 ( .A1(n[89]), .A2(a[5]), .Z(n[153]) );
  AN2D0 U2921 ( .A1(b[4]), .A2(n[26]), .Z(n[89]) );
  AN2D0 U2922 ( .A1(a[8]), .A2(n[536]), .Z(n[1048]) );
  AN2D0 U2923 ( .A1(n[280]), .A2(a[7]), .Z(n[536]) );
  AN2D0 U2924 ( .A1(n[152]), .A2(a[6]), .Z(n[280]) );
  AN2D0 U2925 ( .A1(n[88]), .A2(a[5]), .Z(n[152]) );
  AN2D0 U2926 ( .A1(b[4]), .A2(n[25]), .Z(n[88]) );
  AN2D0 U2927 ( .A1(a[8]), .A2(n[533]), .Z(n[1045]) );
  AN2D0 U2928 ( .A1(n[277]), .A2(a[7]), .Z(n[533]) );
  AN2D0 U2929 ( .A1(n[149]), .A2(a[6]), .Z(n[277]) );
  AN2D0 U2930 ( .A1(n[85]), .A2(a[5]), .Z(n[149]) );
  AN2D0 U2931 ( .A1(n[53]), .A2(a[4]), .Z(n[85]) );
  AN2D0 U2932 ( .A1(a[8]), .A2(n[530]), .Z(n[1042]) );
  AN2D0 U2933 ( .A1(n[274]), .A2(a[7]), .Z(n[530]) );
  AN2D0 U2934 ( .A1(n[146]), .A2(a[6]), .Z(n[274]) );
  AN2D0 U2935 ( .A1(n[82]), .A2(a[5]), .Z(n[146]) );
  AN2D0 U2936 ( .A1(a[4]), .A2(n[50]), .Z(n[82]) );
  AN2D0 U2937 ( .A1(a[8]), .A2(n[529]), .Z(n[1041]) );
  AN2D0 U2938 ( .A1(n[273]), .A2(a[7]), .Z(n[529]) );
  AN2D0 U2939 ( .A1(n[145]), .A2(a[6]), .Z(n[273]) );
  AN2D0 U2940 ( .A1(n[81]), .A2(a[5]), .Z(n[145]) );
  AN2D0 U2941 ( .A1(a[4]), .A2(n[49]), .Z(n[81]) );
  AN2D0 U2942 ( .A1(a[8]), .A2(n[526]), .Z(n[1038]) );
  AN2D0 U2943 ( .A1(n[270]), .A2(a[7]), .Z(n[526]) );
  AN2D0 U2944 ( .A1(n[142]), .A2(a[6]), .Z(n[270]) );
  AN2D0 U2945 ( .A1(n[78]), .A2(a[5]), .Z(n[142]) );
  AN2D0 U2946 ( .A1(a[4]), .A2(n[46]), .Z(n[78]) );
  AN2D0 U2947 ( .A1(a[8]), .A2(n[523]), .Z(n[1035]) );
  AN2D0 U2948 ( .A1(n[267]), .A2(a[7]), .Z(n[523]) );
  AN2D0 U2949 ( .A1(n[139]), .A2(a[6]), .Z(n[267]) );
  AN2D0 U2950 ( .A1(n[75]), .A2(a[5]), .Z(n[139]) );
  AN2D0 U2951 ( .A1(n[43]), .A2(a[4]), .Z(n[75]) );
  AN2D0 U2952 ( .A1(n[12]), .A2(b[3]), .Z(n[43]) );
  AN2D0 U2953 ( .A1(a[8]), .A2(n[522]), .Z(n[1034]) );
  AN2D0 U2954 ( .A1(n[266]), .A2(a[7]), .Z(n[522]) );
  AN2D0 U2955 ( .A1(n[138]), .A2(a[6]), .Z(n[266]) );
  AN2D0 U2956 ( .A1(n[74]), .A2(a[5]), .Z(n[138]) );
  AN2D0 U2957 ( .A1(n[42]), .A2(a[4]), .Z(n[74]) );
  AN2D0 U2958 ( .A1(b[3]), .A2(n[11]), .Z(n[42]) );
  AN2D0 U2959 ( .A1(a[8]), .A2(n[521]), .Z(n[1033]) );
  AN2D0 U2960 ( .A1(n[265]), .A2(a[7]), .Z(n[521]) );
  AN2D0 U2961 ( .A1(n[137]), .A2(a[6]), .Z(n[265]) );
  AN2D0 U2962 ( .A1(n[73]), .A2(a[5]), .Z(n[137]) );
  AN2D0 U2963 ( .A1(n[41]), .A2(a[4]), .Z(n[73]) );
  AN2D0 U2964 ( .A1(b[3]), .A2(n[10]), .Z(n[41]) );
  AN2D0 U2965 ( .A1(a[8]), .A2(n[518]), .Z(n[1030]) );
  AN2D0 U2966 ( .A1(n[262]), .A2(a[7]), .Z(n[518]) );
  AN2D0 U2967 ( .A1(n[134]), .A2(a[6]), .Z(n[262]) );
  AN2D0 U2968 ( .A1(n[70]), .A2(a[5]), .Z(n[134]) );
  AN2D0 U2969 ( .A1(n[38]), .A2(a[4]), .Z(n[70]) );
  AN2D0 U2970 ( .A1(a[8]), .A2(n[515]), .Z(n[1027]) );
  AN2D0 U2971 ( .A1(n[259]), .A2(a[7]), .Z(n[515]) );
  AN2D0 U2972 ( .A1(n[131]), .A2(a[6]), .Z(n[259]) );
  AN2D0 U2973 ( .A1(n[67]), .A2(a[5]), .Z(n[131]) );
  AN2D0 U2974 ( .A1(n[35]), .A2(a[4]), .Z(n[67]) );
  AN2D0 U2975 ( .A1(a[3]), .A2(n[19]), .Z(n[35]) );
  AN2D0 U2976 ( .A1(a[8]), .A2(n[514]), .Z(n[1026]) );
  AN2D0 U2977 ( .A1(n[258]), .A2(a[7]), .Z(n[514]) );
  AN2D0 U2978 ( .A1(n[130]), .A2(a[6]), .Z(n[258]) );
  AN2D0 U2979 ( .A1(n[66]), .A2(a[5]), .Z(n[130]) );
  AN2D0 U2980 ( .A1(n[34]), .A2(a[4]), .Z(n[66]) );
  AN2D0 U2981 ( .A1(a[3]), .A2(n[18]), .Z(n[34]) );
  AN2D0 U2982 ( .A1(a[8]), .A2(n[511]), .Z(n[1023]) );
  AN2D0 U2983 ( .A1(n[255]), .A2(a[7]), .Z(n[511]) );
  AN2D0 U2984 ( .A1(n[127]), .A2(a[6]), .Z(n[255]) );
  AN2D0 U2985 ( .A1(n[63]), .A2(a[5]), .Z(n[127]) );
  AN2D0 U2986 ( .A1(n[31]), .A2(a[4]), .Z(n[63]) );
  AN2D0 U2987 ( .A1(a[3]), .A2(n[15]), .Z(n[31]) );
  AN2D0 U2988 ( .A1(a[8]), .A2(n[508]), .Z(n[1020]) );
  AN2D0 U2989 ( .A1(n[252]), .A2(a[7]), .Z(n[508]) );
  AN2D0 U2990 ( .A1(n[124]), .A2(a[6]), .Z(n[252]) );
  AN2D0 U2991 ( .A1(n[60]), .A2(a[5]), .Z(n[124]) );
  AN2D0 U2992 ( .A1(n[28]), .A2(a[4]), .Z(n[60]) );
  AN2D0 U2993 ( .A1(n[12]), .A2(a[3]), .Z(n[28]) );
  AN2D0 U2994 ( .A1(n[4]), .A2(a[2]), .Z(n[12]) );
  AN2D0 U2995 ( .A1(b[4]), .A2(n[38]), .Z(n[101]) );
  AN2D0 U2996 ( .A1(n[22]), .A2(a[3]), .Z(n[38]) );
  AN2D0 U2997 ( .A1(a[8]), .A2(n[507]), .Z(n[1019]) );
  AN2D0 U2998 ( .A1(n[251]), .A2(a[7]), .Z(n[507]) );
  AN2D0 U2999 ( .A1(n[123]), .A2(a[6]), .Z(n[251]) );
  AN2D0 U3000 ( .A1(n[59]), .A2(a[5]), .Z(n[123]) );
  AN2D0 U3001 ( .A1(n[27]), .A2(a[4]), .Z(n[59]) );
  AN2D0 U3002 ( .A1(n[11]), .A2(a[3]), .Z(n[27]) );
  AN2D0 U3003 ( .A1(a[2]), .A2(n[3]), .Z(n[11]) );
  AN2D0 U3004 ( .A1(a[8]), .A2(n[506]), .Z(n[1018]) );
  AN2D0 U3005 ( .A1(n[250]), .A2(a[7]), .Z(n[506]) );
  AN2D0 U3006 ( .A1(n[122]), .A2(a[6]), .Z(n[250]) );
  AN2D0 U3007 ( .A1(n[58]), .A2(a[5]), .Z(n[122]) );
  AN2D0 U3008 ( .A1(n[26]), .A2(a[4]), .Z(n[58]) );
  AN2D0 U3009 ( .A1(n[10]), .A2(a[3]), .Z(n[26]) );
  AN2D0 U3010 ( .A1(a[2]), .A2(b[2]), .Z(n[10]) );
  AN2D0 U3011 ( .A1(a[8]), .A2(n[505]), .Z(n[1017]) );
  AN2D0 U3012 ( .A1(n[249]), .A2(a[7]), .Z(n[505]) );
  AN2D0 U3013 ( .A1(n[121]), .A2(a[6]), .Z(n[249]) );
  AN2D0 U3014 ( .A1(n[57]), .A2(a[5]), .Z(n[121]) );
  AN2D0 U3015 ( .A1(n[25]), .A2(a[4]), .Z(n[57]) );
  AN2D0 U3016 ( .A1(b[3]), .A2(a[3]), .Z(n[25]) );
  AN2D0 U3017 ( .A1(a[8]), .A2(n[504]), .Z(n[1016]) );
  AN2D0 U3018 ( .A1(n[248]), .A2(a[7]), .Z(n[504]) );
  AN2D0 U3019 ( .A1(n[120]), .A2(a[6]), .Z(n[248]) );
  AN2D0 U3020 ( .A1(n[56]), .A2(a[5]), .Z(n[120]) );
  AN2D0 U3021 ( .A1(b[4]), .A2(a[4]), .Z(n[56]) );
  AN2D0 U3022 ( .A1(a[8]), .A2(n[503]), .Z(n[1015]) );
  AN2D0 U3023 ( .A1(n[247]), .A2(a[7]), .Z(n[503]) );
  AN2D0 U3024 ( .A1(n[119]), .A2(a[6]), .Z(n[247]) );
  AN2D0 U3025 ( .A1(b[5]), .A2(a[5]), .Z(n[119]) );
  AN2D0 U3026 ( .A1(a[8]), .A2(n[502]), .Z(n[1014]) );
  AN2D0 U3027 ( .A1(n[246]), .A2(a[7]), .Z(n[502]) );
  AN2D0 U3028 ( .A1(b[6]), .A2(a[6]), .Z(n[246]) );
  AN2D0 U3029 ( .A1(a[8]), .A2(n[501]), .Z(n[1013]) );
  AN2D0 U3030 ( .A1(b[7]), .A2(a[7]), .Z(n[501]) );
  AN2D0 U3031 ( .A1(a[8]), .A2(b[8]), .Z(n[1012]) );
  AN2D0 U3032 ( .A1(b[7]), .A2(n[498]), .Z(n[1009]) );
  AN2D0 U3033 ( .A1(b[6]), .A2(n[243]), .Z(n[498]) );
  AN2D0 U3034 ( .A1(b[5]), .A2(n[116]), .Z(n[243]) );
  AN2D0 U3035 ( .A1(b[4]), .A2(n[53]), .Z(n[116]) );
  AN2D0 U3036 ( .A1(b[3]), .A2(n[22]), .Z(n[53]) );
  AN2D0 U3037 ( .A1(b[2]), .A2(n[7]), .Z(n[22]) );
  AN2D0 U3038 ( .A1(b[7]), .A2(n[495]), .Z(n[1006]) );
  AN2D0 U3039 ( .A1(b[6]), .A2(n[240]), .Z(n[495]) );
  AN2D0 U3040 ( .A1(b[5]), .A2(n[113]), .Z(n[240]) );
  AN2D0 U3041 ( .A1(b[4]), .A2(n[50]), .Z(n[113]) );
  AN2D0 U3042 ( .A1(b[3]), .A2(n[19]), .Z(n[50]) );
  AN2D0 U3043 ( .A1(n[4]), .A2(b[2]), .Z(n[19]) );
  AN2D0 U3044 ( .A1(n[0]), .A2(a[1]), .Z(n[4]) );
  AN2D0 U3045 ( .A1(b[7]), .A2(n[494]), .Z(n[1005]) );
  AN2D0 U3046 ( .A1(b[6]), .A2(n[239]), .Z(n[494]) );
  AN2D0 U3047 ( .A1(b[5]), .A2(n[112]), .Z(n[239]) );
  AN2D0 U3048 ( .A1(b[4]), .A2(n[49]), .Z(n[112]) );
  AN2D0 U3049 ( .A1(b[3]), .A2(n[18]), .Z(n[49]) );
  AN2D0 U3050 ( .A1(n[3]), .A2(b[2]), .Z(n[18]) );
  AN2D0 U3051 ( .A1(a[1]), .A2(b[1]), .Z(n[3]) );
  AN2D0 U3052 ( .A1(b[7]), .A2(n[491]), .Z(n[1002]) );
  AN2D0 U3053 ( .A1(b[6]), .A2(n[236]), .Z(n[491]) );
  AN2D0 U3054 ( .A1(b[5]), .A2(n[109]), .Z(n[236]) );
  AN2D0 U3055 ( .A1(b[4]), .A2(n[46]), .Z(n[109]) );
  AN2D0 U3056 ( .A1(b[3]), .A2(n[15]), .Z(n[46]) );
  AN2D0 U3057 ( .A1(a[2]), .A2(n[7]), .Z(n[15]) );
  AN2D0 U3058 ( .A1(n[0]), .A2(b[1]), .Z(n[7]) );
  AN2D0 U3059 ( .A1(b[0]), .A2(a[0]), .Z(n[0]) );
endmodule


module gen_cla_decomposed ( a, b, s );
  input [9:0] a;
  input [9:0] b;
  output [9:0] s;

  wire   [2034:0] n;

  gen_nonlinear_part NLIN ( .a(a), .b(b), .n(n) );
  gen_linear_part LIN ( .a(a), .b(b), .n({1'b0, 1'b0, n[2032], 1'b0, 1'b0, 
        n[2029:2028], 1'b0, 1'b0, n[2025], 1'b0, 1'b0, n[2022:2020], 1'b0, 
        1'b0, n[2017], 1'b0, 1'b0, n[2014:2013], 1'b0, 1'b0, n[2010], 1'b0, 
        1'b0, n[2007:2004], 1'b0, 1'b0, n[2001], 1'b0, 1'b0, n[1998:1997], 
        1'b0, 1'b0, n[1994], 1'b0, 1'b0, n[1991:1989], 1'b0, 1'b0, n[1986], 
        1'b0, 1'b0, n[1983:1982], 1'b0, 1'b0, n[1979], 1'b0, 1'b0, 
        n[1976:1972], 1'b0, 1'b0, n[1969], 1'b0, 1'b0, n[1966:1965], 1'b0, 
        1'b0, n[1962], 1'b0, 1'b0, n[1959:1957], 1'b0, 1'b0, n[1954], 1'b0, 
        1'b0, n[1951:1950], 1'b0, 1'b0, n[1947], 1'b0, 1'b0, n[1944:1941], 
        1'b0, 1'b0, n[1938], 1'b0, 1'b0, n[1935:1934], 1'b0, 1'b0, n[1931], 
        1'b0, 1'b0, n[1928:1926], 1'b0, 1'b0, n[1923], 1'b0, 1'b0, 
        n[1920:1919], 1'b0, 1'b0, n[1916], 1'b0, 1'b0, n[1913:1908], 1'b0, 
        1'b0, n[1905], 1'b0, 1'b0, n[1902:1901], 1'b0, 1'b0, n[1898], 1'b0, 
        1'b0, n[1895:1893], 1'b0, 1'b0, n[1890], 1'b0, 1'b0, n[1887:1886], 
        1'b0, 1'b0, n[1883], 1'b0, 1'b0, n[1880:1877], 1'b0, 1'b0, n[1874], 
        1'b0, 1'b0, n[1871:1870], 1'b0, 1'b0, n[1867], 1'b0, 1'b0, 
        n[1864:1862], 1'b0, 1'b0, n[1859], 1'b0, 1'b0, n[1856:1855], 1'b0, 
        1'b0, n[1852], 1'b0, 1'b0, n[1849:1845], 1'b0, 1'b0, n[1842], 1'b0, 
        1'b0, n[1839:1838], 1'b0, 1'b0, n[1835], 1'b0, 1'b0, n[1832:1830], 
        1'b0, 1'b0, n[1827], 1'b0, 1'b0, n[1824:1823], 1'b0, 1'b0, n[1820], 
        1'b0, 1'b0, n[1817:1814], 1'b0, 1'b0, n[1811], 1'b0, 1'b0, 
        n[1808:1807], 1'b0, 1'b0, n[1804], 1'b0, 1'b0, n[1801:1799], 1'b0, 
        1'b0, n[1796], 1'b0, 1'b0, n[1793:1792], 1'b0, 1'b0, n[1789], 1'b0, 
        1'b0, n[1786:1780], 1'b0, 1'b0, n[1777], 1'b0, 1'b0, n[1774:1773], 
        1'b0, 1'b0, n[1770], 1'b0, 1'b0, n[1767:1765], 1'b0, 1'b0, n[1762], 
        1'b0, 1'b0, n[1759:1758], 1'b0, 1'b0, n[1755], 1'b0, 1'b0, 
        n[1752:1749], 1'b0, 1'b0, n[1746], 1'b0, 1'b0, n[1743:1742], 1'b0, 
        1'b0, n[1739], 1'b0, 1'b0, n[1736:1734], 1'b0, 1'b0, n[1731], 1'b0, 
        1'b0, n[1728:1727], 1'b0, 1'b0, n[1724], 1'b0, 1'b0, n[1721:1717], 
        1'b0, 1'b0, n[1714], 1'b0, 1'b0, n[1711:1710], 1'b0, 1'b0, n[1707], 
        1'b0, 1'b0, n[1704:1702], 1'b0, 1'b0, n[1699], 1'b0, 1'b0, 
        n[1696:1695], 1'b0, 1'b0, n[1692], 1'b0, 1'b0, n[1689:1686], 1'b0, 
        1'b0, n[1683], 1'b0, 1'b0, n[1680:1679], 1'b0, 1'b0, n[1676], 1'b0, 
        1'b0, n[1673:1671], 1'b0, 1'b0, n[1668], 1'b0, 1'b0, n[1665:1664], 
        1'b0, 1'b0, n[1661], 1'b0, 1'b0, n[1658:1653], 1'b0, 1'b0, n[1650], 
        1'b0, 1'b0, n[1647:1646], 1'b0, 1'b0, n[1643], 1'b0, 1'b0, 
        n[1640:1638], 1'b0, 1'b0, n[1635], 1'b0, 1'b0, n[1632:1631], 1'b0, 
        1'b0, n[1628], 1'b0, 1'b0, n[1625:1622], 1'b0, 1'b0, n[1619], 1'b0, 
        1'b0, n[1616:1615], 1'b0, 1'b0, n[1612], 1'b0, 1'b0, n[1609:1607], 
        1'b0, 1'b0, n[1604], 1'b0, 1'b0, n[1601:1600], 1'b0, 1'b0, n[1597], 
        1'b0, 1'b0, n[1594:1590], 1'b0, 1'b0, n[1587], 1'b0, 1'b0, 
        n[1584:1583], 1'b0, 1'b0, n[1580], 1'b0, 1'b0, n[1577:1575], 1'b0, 
        1'b0, n[1572], 1'b0, 1'b0, n[1569:1568], 1'b0, 1'b0, n[1565], 1'b0, 
        1'b0, n[1562:1559], 1'b0, 1'b0, n[1556], 1'b0, 1'b0, n[1553:1552], 
        1'b0, 1'b0, n[1549], 1'b0, 1'b0, n[1546:1544], 1'b0, 1'b0, n[1541], 
        1'b0, 1'b0, n[1538:1537], 1'b0, 1'b0, n[1534], 1'b0, 1'b0, 
        n[1531:1524], 1'b0, 1'b0, n[1521], 1'b0, 1'b0, n[1518:1517], 1'b0, 
        1'b0, n[1514], 1'b0, 1'b0, n[1511:1509], 1'b0, 1'b0, n[1506], 1'b0, 
        1'b0, n[1503:1502], 1'b0, 1'b0, n[1499], 1'b0, 1'b0, n[1496:1493], 
        1'b0, 1'b0, n[1490], 1'b0, 1'b0, n[1487:1486], 1'b0, 1'b0, n[1483], 
        1'b0, 1'b0, n[1480:1478], 1'b0, 1'b0, n[1475], 1'b0, 1'b0, 
        n[1472:1471], 1'b0, 1'b0, n[1468], 1'b0, 1'b0, n[1465:1461], 1'b0, 
        1'b0, n[1458], 1'b0, 1'b0, n[1455:1454], 1'b0, 1'b0, n[1451], 1'b0, 
        1'b0, n[1448:1446], 1'b0, 1'b0, n[1443], 1'b0, 1'b0, n[1440:1439], 
        1'b0, 1'b0, n[1436], 1'b0, 1'b0, n[1433:1430], 1'b0, 1'b0, n[1427], 
        1'b0, 1'b0, n[1424:1423], 1'b0, 1'b0, n[1420], 1'b0, 1'b0, 
        n[1417:1415], 1'b0, 1'b0, n[1412], 1'b0, 1'b0, n[1409:1408], 1'b0, 
        1'b0, n[1405], 1'b0, 1'b0, n[1402:1397], 1'b0, 1'b0, n[1394], 1'b0, 
        1'b0, n[1391:1390], 1'b0, 1'b0, n[1387], 1'b0, 1'b0, n[1384:1382], 
        1'b0, 1'b0, n[1379], 1'b0, 1'b0, n[1376:1375], 1'b0, 1'b0, n[1372], 
        1'b0, 1'b0, n[1369:1366], 1'b0, 1'b0, n[1363], 1'b0, 1'b0, 
        n[1360:1359], 1'b0, 1'b0, n[1356], 1'b0, 1'b0, n[1353:1351], 1'b0, 
        1'b0, n[1348], 1'b0, 1'b0, n[1345:1344], 1'b0, 1'b0, n[1341], 1'b0, 
        1'b0, n[1338:1334], 1'b0, 1'b0, n[1331], 1'b0, 1'b0, n[1328:1327], 
        1'b0, 1'b0, n[1324], 1'b0, 1'b0, n[1321:1319], 1'b0, 1'b0, n[1316], 
        1'b0, 1'b0, n[1313:1312], 1'b0, 1'b0, n[1309], 1'b0, 1'b0, 
        n[1306:1303], 1'b0, 1'b0, n[1300], 1'b0, 1'b0, n[1297:1296], 1'b0, 
        1'b0, n[1293], 1'b0, 1'b0, n[1290:1288], 1'b0, 1'b0, n[1285], 1'b0, 
        1'b0, n[1282:1281], 1'b0, 1'b0, n[1278], 1'b0, 1'b0, n[1275:1269], 
        1'b0, 1'b0, n[1266], 1'b0, 1'b0, n[1263:1262], 1'b0, 1'b0, n[1259], 
        1'b0, 1'b0, n[1256:1254], 1'b0, 1'b0, n[1251], 1'b0, 1'b0, 
        n[1248:1247], 1'b0, 1'b0, n[1244], 1'b0, 1'b0, n[1241:1238], 1'b0, 
        1'b0, n[1235], 1'b0, 1'b0, n[1232:1231], 1'b0, 1'b0, n[1228], 1'b0, 
        1'b0, n[1225:1223], 1'b0, 1'b0, n[1220], 1'b0, 1'b0, n[1217:1216], 
        1'b0, 1'b0, n[1213], 1'b0, 1'b0, n[1210:1206], 1'b0, 1'b0, n[1203], 
        1'b0, 1'b0, n[1200:1199], 1'b0, 1'b0, n[1196], 1'b0, 1'b0, 
        n[1193:1191], 1'b0, 1'b0, n[1188], 1'b0, 1'b0, n[1185:1184], 1'b0, 
        1'b0, n[1181], 1'b0, 1'b0, n[1178:1175], 1'b0, 1'b0, n[1172], 1'b0, 
        1'b0, n[1169:1168], 1'b0, 1'b0, n[1165], 1'b0, 1'b0, n[1162:1160], 
        1'b0, 1'b0, n[1157], 1'b0, 1'b0, n[1154:1153], 1'b0, 1'b0, n[1150], 
        1'b0, 1'b0, n[1147:1142], 1'b0, 1'b0, n[1139], 1'b0, 1'b0, 
        n[1136:1135], 1'b0, 1'b0, n[1132], 1'b0, 1'b0, n[1129:1127], 1'b0, 
        1'b0, n[1124], 1'b0, 1'b0, n[1121:1120], 1'b0, 1'b0, n[1117], 1'b0, 
        1'b0, n[1114:1111], 1'b0, 1'b0, n[1108], 1'b0, 1'b0, n[1105:1104], 
        1'b0, 1'b0, n[1101], 1'b0, 1'b0, n[1098:1096], 1'b0, 1'b0, n[1093], 
        1'b0, 1'b0, n[1090:1089], 1'b0, 1'b0, n[1086], 1'b0, 1'b0, 
        n[1083:1079], 1'b0, 1'b0, n[1076], 1'b0, 1'b0, n[1073:1072], 1'b0, 
        1'b0, n[1069], 1'b0, 1'b0, n[1066:1064], 1'b0, 1'b0, n[1061], 1'b0, 
        1'b0, n[1058:1057], 1'b0, 1'b0, n[1054], 1'b0, 1'b0, n[1051:1048], 
        1'b0, 1'b0, n[1045], 1'b0, 1'b0, n[1042:1041], 1'b0, 1'b0, n[1038], 
        1'b0, 1'b0, n[1035:1033], 1'b0, 1'b0, n[1030], 1'b0, 1'b0, 
        n[1027:1026], 1'b0, 1'b0, n[1023], 1'b0, 1'b0, n[1020:1012], 1'b0, 
        1'b0, n[1009], 1'b0, 1'b0, n[1006:1005], 1'b0, 1'b0, n[1002], 1'b0, 
        1'b0, n[999:997], 1'b0, 1'b0, n[994], 1'b0, 1'b0, n[991:990], 1'b0, 
        1'b0, n[987], 1'b0, 1'b0, n[984:981], 1'b0, 1'b0, n[978], 1'b0, 1'b0, 
        n[975:974], 1'b0, 1'b0, n[971], 1'b0, 1'b0, n[968:966], 1'b0, 1'b0, 
        n[963], 1'b0, 1'b0, n[960:959], 1'b0, 1'b0, n[956], 1'b0, 1'b0, 
        n[953:949], 1'b0, 1'b0, n[946], 1'b0, 1'b0, n[943:942], 1'b0, 1'b0, 
        n[939], 1'b0, 1'b0, n[936:934], 1'b0, 1'b0, n[931], 1'b0, 1'b0, 
        n[928:927], 1'b0, 1'b0, n[924], 1'b0, 1'b0, n[921:918], 1'b0, 1'b0, 
        n[915], 1'b0, 1'b0, n[912:911], 1'b0, 1'b0, n[908], 1'b0, 1'b0, 
        n[905:903], 1'b0, 1'b0, n[900], 1'b0, 1'b0, n[897:896], 1'b0, 1'b0, 
        n[893], 1'b0, 1'b0, n[890:885], 1'b0, 1'b0, n[882], 1'b0, 1'b0, 
        n[879:878], 1'b0, 1'b0, n[875], 1'b0, 1'b0, n[872:870], 1'b0, 1'b0, 
        n[867], 1'b0, 1'b0, n[864:863], 1'b0, 1'b0, n[860], 1'b0, 1'b0, 
        n[857:854], 1'b0, 1'b0, n[851], 1'b0, 1'b0, n[848:847], 1'b0, 1'b0, 
        n[844], 1'b0, 1'b0, n[841:839], 1'b0, 1'b0, n[836], 1'b0, 1'b0, 
        n[833:832], 1'b0, 1'b0, n[829], 1'b0, 1'b0, n[826:822], 1'b0, 1'b0, 
        n[819], 1'b0, 1'b0, n[816:815], 1'b0, 1'b0, n[812], 1'b0, 1'b0, 
        n[809:807], 1'b0, 1'b0, n[804], 1'b0, 1'b0, n[801:800], 1'b0, 1'b0, 
        n[797], 1'b0, 1'b0, n[794:791], 1'b0, 1'b0, n[788], 1'b0, 1'b0, 
        n[785:784], 1'b0, 1'b0, n[781], 1'b0, 1'b0, n[778:776], 1'b0, 1'b0, 
        n[773], 1'b0, 1'b0, n[770:769], 1'b0, 1'b0, n[766], 1'b0, 1'b0, 
        n[763:757], 1'b0, 1'b0, n[754], 1'b0, 1'b0, n[751:750], 1'b0, 1'b0, 
        n[747], 1'b0, 1'b0, n[744:742], 1'b0, 1'b0, n[739], 1'b0, 1'b0, 
        n[736:735], 1'b0, 1'b0, n[732], 1'b0, 1'b0, n[729:726], 1'b0, 1'b0, 
        n[723], 1'b0, 1'b0, n[720:719], 1'b0, 1'b0, n[716], 1'b0, 1'b0, 
        n[713:711], 1'b0, 1'b0, n[708], 1'b0, 1'b0, n[705:704], 1'b0, 1'b0, 
        n[701], 1'b0, 1'b0, n[698:694], 1'b0, 1'b0, n[691], 1'b0, 1'b0, 
        n[688:687], 1'b0, 1'b0, n[684], 1'b0, 1'b0, n[681:679], 1'b0, 1'b0, 
        n[676], 1'b0, 1'b0, n[673:672], 1'b0, 1'b0, n[669], 1'b0, 1'b0, 
        n[666:663], 1'b0, 1'b0, n[660], 1'b0, 1'b0, n[657:656], 1'b0, 1'b0, 
        n[653], 1'b0, 1'b0, n[650:648], 1'b0, 1'b0, n[645], 1'b0, 1'b0, 
        n[642:641], 1'b0, 1'b0, n[638], 1'b0, 1'b0, n[635:630], 1'b0, 1'b0, 
        n[627], 1'b0, 1'b0, n[624:623], 1'b0, 1'b0, n[620], 1'b0, 1'b0, 
        n[617:615], 1'b0, 1'b0, n[612], 1'b0, 1'b0, n[609:608], 1'b0, 1'b0, 
        n[605], 1'b0, 1'b0, n[602:599], 1'b0, 1'b0, n[596], 1'b0, 1'b0, 
        n[593:592], 1'b0, 1'b0, n[589], 1'b0, 1'b0, n[586:584], 1'b0, 1'b0, 
        n[581], 1'b0, 1'b0, n[578:577], 1'b0, 1'b0, n[574], 1'b0, 1'b0, 
        n[571:567], 1'b0, 1'b0, n[564], 1'b0, 1'b0, n[561:560], 1'b0, 1'b0, 
        n[557], 1'b0, 1'b0, n[554:552], 1'b0, 1'b0, n[549], 1'b0, 1'b0, 
        n[546:545], 1'b0, 1'b0, n[542], 1'b0, 1'b0, n[539:536], 1'b0, 1'b0, 
        n[533], 1'b0, 1'b0, n[530:529], 1'b0, 1'b0, n[526], 1'b0, 1'b0, 
        n[523:521], 1'b0, 1'b0, n[518], 1'b0, 1'b0, n[515:514], 1'b0, 1'b0, 
        n[511], 1'b0, 1'b0, n[508:501], 1'b0, 1'b0, n[498], 1'b0, 1'b0, 
        n[495:494], 1'b0, 1'b0, n[491], 1'b0, 1'b0, n[488:486], 1'b0, 1'b0, 
        n[483], 1'b0, 1'b0, n[480:479], 1'b0, 1'b0, n[476], 1'b0, 1'b0, 
        n[473:470], 1'b0, 1'b0, n[467], 1'b0, 1'b0, n[464:463], 1'b0, 1'b0, 
        n[460], 1'b0, 1'b0, n[457:455], 1'b0, 1'b0, n[452], 1'b0, 1'b0, 
        n[449:448], 1'b0, 1'b0, n[445], 1'b0, 1'b0, n[442:438], 1'b0, 1'b0, 
        n[435], 1'b0, 1'b0, n[432:431], 1'b0, 1'b0, n[428], 1'b0, 1'b0, 
        n[425:423], 1'b0, 1'b0, n[420], 1'b0, 1'b0, n[417:416], 1'b0, 1'b0, 
        n[413], 1'b0, 1'b0, n[410:407], 1'b0, 1'b0, n[404], 1'b0, 1'b0, 
        n[401:400], 1'b0, 1'b0, n[397], 1'b0, 1'b0, n[394:392], 1'b0, 1'b0, 
        n[389], 1'b0, 1'b0, n[386:385], 1'b0, 1'b0, n[382], 1'b0, 1'b0, 
        n[379:374], 1'b0, 1'b0, n[371], 1'b0, 1'b0, n[368:367], 1'b0, 1'b0, 
        n[364], 1'b0, 1'b0, n[361:359], 1'b0, 1'b0, n[356], 1'b0, 1'b0, 
        n[353:352], 1'b0, 1'b0, n[349], 1'b0, 1'b0, n[346:343], 1'b0, 1'b0, 
        n[340], 1'b0, 1'b0, n[337:336], 1'b0, 1'b0, n[333], 1'b0, 1'b0, 
        n[330:328], 1'b0, 1'b0, n[325], 1'b0, 1'b0, n[322:321], 1'b0, 1'b0, 
        n[318], 1'b0, 1'b0, n[315:311], 1'b0, 1'b0, n[308], 1'b0, 1'b0, 
        n[305:304], 1'b0, 1'b0, n[301], 1'b0, 1'b0, n[298:296], 1'b0, 1'b0, 
        n[293], 1'b0, 1'b0, n[290:289], 1'b0, 1'b0, n[286], 1'b0, 1'b0, 
        n[283:280], 1'b0, 1'b0, n[277], 1'b0, 1'b0, n[274:273], 1'b0, 1'b0, 
        n[270], 1'b0, 1'b0, n[267:265], 1'b0, 1'b0, n[262], 1'b0, 1'b0, 
        n[259:258], 1'b0, 1'b0, n[255], 1'b0, 1'b0, n[252:246], 1'b0, 1'b0, 
        n[243], 1'b0, 1'b0, n[240:239], 1'b0, 1'b0, n[236], 1'b0, 1'b0, 
        n[233:231], 1'b0, 1'b0, n[228], 1'b0, 1'b0, n[225:224], 1'b0, 1'b0, 
        n[221], 1'b0, 1'b0, n[218:215], 1'b0, 1'b0, n[212], 1'b0, 1'b0, 
        n[209:208], 1'b0, 1'b0, n[205], 1'b0, 1'b0, n[202:200], 1'b0, 1'b0, 
        n[197], 1'b0, 1'b0, n[194:193], 1'b0, 1'b0, n[190], 1'b0, 1'b0, 
        n[187:183], 1'b0, 1'b0, n[180], 1'b0, 1'b0, n[177:176], 1'b0, 1'b0, 
        n[173], 1'b0, 1'b0, n[170:168], 1'b0, 1'b0, n[165], 1'b0, 1'b0, 
        n[162:161], 1'b0, 1'b0, n[158], 1'b0, 1'b0, n[155:152], 1'b0, 1'b0, 
        n[149], 1'b0, 1'b0, n[146:145], 1'b0, 1'b0, n[142], 1'b0, 1'b0, 
        n[139:137], 1'b0, 1'b0, n[134], 1'b0, 1'b0, n[131:130], 1'b0, 1'b0, 
        n[127], 1'b0, 1'b0, n[124:119], 1'b0, 1'b0, n[116], 1'b0, 1'b0, 
        n[113:112], 1'b0, 1'b0, n[109], 1'b0, 1'b0, n[106:104], 1'b0, 1'b0, 
        n[101], 1'b0, 1'b0, n[98:97], 1'b0, 1'b0, n[94], 1'b0, 1'b0, n[91:88], 
        1'b0, 1'b0, n[85], 1'b0, 1'b0, n[82:81], 1'b0, 1'b0, n[78], 1'b0, 1'b0, 
        n[75:73], 1'b0, 1'b0, n[70], 1'b0, 1'b0, n[67:66], 1'b0, 1'b0, n[63], 
        1'b0, 1'b0, n[60:56], 1'b0, 1'b0, n[53], 1'b0, 1'b0, n[50:49], 1'b0, 
        1'b0, n[46], 1'b0, 1'b0, n[43:41], 1'b0, 1'b0, n[38], 1'b0, 1'b0, 
        n[35:34], 1'b0, 1'b0, n[31], 1'b0, 1'b0, n[28:25], 1'b0, 1'b0, n[22], 
        1'b0, 1'b0, n[19:18], 1'b0, 1'b0, n[15], 1'b0, 1'b0, n[12:10], 1'b0, 
        1'b0, n[7], 1'b0, 1'b0, n[4:3], 1'b0, 1'b0, n[0]}), .s(s) );
endmodule

