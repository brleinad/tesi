
module cla_adder ( a, b, s, cin, cout );
  input [255:0] a;
  input [255:0] b;
  output [255:0] s;
  input cin;
  output cout;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242,
         N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253,
         N254;
  wire   [254:0] g;
  wire   [255:0] p;
  wire   [255:1] c;

  XOR2D0 C2306 ( .A1(p[0]), .A2(cin), .Z(s[0]) );
  XOR2D0 C2305 ( .A1(p[1]), .A2(c[1]), .Z(s[1]) );
  XOR2D0 C2304 ( .A1(p[2]), .A2(c[2]), .Z(s[2]) );
  XOR2D0 C2303 ( .A1(p[3]), .A2(c[3]), .Z(s[3]) );
  XOR2D0 C2302 ( .A1(p[4]), .A2(c[4]), .Z(s[4]) );
  XOR2D0 C2301 ( .A1(p[5]), .A2(c[5]), .Z(s[5]) );
  XOR2D0 C2300 ( .A1(p[6]), .A2(c[6]), .Z(s[6]) );
  XOR2D0 C2299 ( .A1(p[7]), .A2(c[7]), .Z(s[7]) );
  XOR2D0 C2298 ( .A1(p[8]), .A2(c[8]), .Z(s[8]) );
  XOR2D0 C2297 ( .A1(p[9]), .A2(c[9]), .Z(s[9]) );
  XOR2D0 C2296 ( .A1(p[10]), .A2(c[10]), .Z(s[10]) );
  XOR2D0 C2295 ( .A1(p[11]), .A2(c[11]), .Z(s[11]) );
  XOR2D0 C2294 ( .A1(p[12]), .A2(c[12]), .Z(s[12]) );
  XOR2D0 C2293 ( .A1(p[13]), .A2(c[13]), .Z(s[13]) );
  XOR2D0 C2292 ( .A1(p[14]), .A2(c[14]), .Z(s[14]) );
  XOR2D0 C2291 ( .A1(p[15]), .A2(c[15]), .Z(s[15]) );
  XOR2D0 C2290 ( .A1(p[16]), .A2(c[16]), .Z(s[16]) );
  XOR2D0 C2289 ( .A1(p[17]), .A2(c[17]), .Z(s[17]) );
  XOR2D0 C2288 ( .A1(p[18]), .A2(c[18]), .Z(s[18]) );
  XOR2D0 C2287 ( .A1(p[19]), .A2(c[19]), .Z(s[19]) );
  XOR2D0 C2286 ( .A1(p[20]), .A2(c[20]), .Z(s[20]) );
  XOR2D0 C2285 ( .A1(p[21]), .A2(c[21]), .Z(s[21]) );
  XOR2D0 C2284 ( .A1(p[22]), .A2(c[22]), .Z(s[22]) );
  XOR2D0 C2283 ( .A1(p[23]), .A2(c[23]), .Z(s[23]) );
  XOR2D0 C2282 ( .A1(p[24]), .A2(c[24]), .Z(s[24]) );
  XOR2D0 C2281 ( .A1(p[25]), .A2(c[25]), .Z(s[25]) );
  XOR2D0 C2280 ( .A1(p[26]), .A2(c[26]), .Z(s[26]) );
  XOR2D0 C2279 ( .A1(p[27]), .A2(c[27]), .Z(s[27]) );
  XOR2D0 C2278 ( .A1(p[28]), .A2(c[28]), .Z(s[28]) );
  XOR2D0 C2277 ( .A1(p[29]), .A2(c[29]), .Z(s[29]) );
  XOR2D0 C2276 ( .A1(p[30]), .A2(c[30]), .Z(s[30]) );
  XOR2D0 C2275 ( .A1(p[31]), .A2(c[31]), .Z(s[31]) );
  XOR2D0 C2274 ( .A1(p[32]), .A2(c[32]), .Z(s[32]) );
  XOR2D0 C2273 ( .A1(p[33]), .A2(c[33]), .Z(s[33]) );
  XOR2D0 C2272 ( .A1(p[34]), .A2(c[34]), .Z(s[34]) );
  XOR2D0 C2271 ( .A1(p[35]), .A2(c[35]), .Z(s[35]) );
  XOR2D0 C2270 ( .A1(p[36]), .A2(c[36]), .Z(s[36]) );
  XOR2D0 C2269 ( .A1(p[37]), .A2(c[37]), .Z(s[37]) );
  XOR2D0 C2268 ( .A1(p[38]), .A2(c[38]), .Z(s[38]) );
  XOR2D0 C2267 ( .A1(p[39]), .A2(c[39]), .Z(s[39]) );
  XOR2D0 C2266 ( .A1(p[40]), .A2(c[40]), .Z(s[40]) );
  XOR2D0 C2265 ( .A1(p[41]), .A2(c[41]), .Z(s[41]) );
  XOR2D0 C2264 ( .A1(p[42]), .A2(c[42]), .Z(s[42]) );
  XOR2D0 C2263 ( .A1(p[43]), .A2(c[43]), .Z(s[43]) );
  XOR2D0 C2262 ( .A1(p[44]), .A2(c[44]), .Z(s[44]) );
  XOR2D0 C2261 ( .A1(p[45]), .A2(c[45]), .Z(s[45]) );
  XOR2D0 C2260 ( .A1(p[46]), .A2(c[46]), .Z(s[46]) );
  XOR2D0 C2259 ( .A1(p[47]), .A2(c[47]), .Z(s[47]) );
  XOR2D0 C2258 ( .A1(p[48]), .A2(c[48]), .Z(s[48]) );
  XOR2D0 C2257 ( .A1(p[49]), .A2(c[49]), .Z(s[49]) );
  XOR2D0 C2256 ( .A1(p[50]), .A2(c[50]), .Z(s[50]) );
  XOR2D0 C2255 ( .A1(p[51]), .A2(c[51]), .Z(s[51]) );
  XOR2D0 C2254 ( .A1(p[52]), .A2(c[52]), .Z(s[52]) );
  XOR2D0 C2253 ( .A1(p[53]), .A2(c[53]), .Z(s[53]) );
  XOR2D0 C2252 ( .A1(p[54]), .A2(c[54]), .Z(s[54]) );
  XOR2D0 C2251 ( .A1(p[55]), .A2(c[55]), .Z(s[55]) );
  XOR2D0 C2250 ( .A1(p[56]), .A2(c[56]), .Z(s[56]) );
  XOR2D0 C2249 ( .A1(p[57]), .A2(c[57]), .Z(s[57]) );
  XOR2D0 C2248 ( .A1(p[58]), .A2(c[58]), .Z(s[58]) );
  XOR2D0 C2247 ( .A1(p[59]), .A2(c[59]), .Z(s[59]) );
  XOR2D0 C2246 ( .A1(p[60]), .A2(c[60]), .Z(s[60]) );
  XOR2D0 C2245 ( .A1(p[61]), .A2(c[61]), .Z(s[61]) );
  XOR2D0 C2244 ( .A1(p[62]), .A2(c[62]), .Z(s[62]) );
  XOR2D0 C2243 ( .A1(p[63]), .A2(c[63]), .Z(s[63]) );
  XOR2D0 C2242 ( .A1(p[64]), .A2(c[64]), .Z(s[64]) );
  XOR2D0 C2241 ( .A1(p[65]), .A2(c[65]), .Z(s[65]) );
  XOR2D0 C2240 ( .A1(p[66]), .A2(c[66]), .Z(s[66]) );
  XOR2D0 C2239 ( .A1(p[67]), .A2(c[67]), .Z(s[67]) );
  XOR2D0 C2238 ( .A1(p[68]), .A2(c[68]), .Z(s[68]) );
  XOR2D0 C2237 ( .A1(p[69]), .A2(c[69]), .Z(s[69]) );
  XOR2D0 C2236 ( .A1(p[70]), .A2(c[70]), .Z(s[70]) );
  XOR2D0 C2235 ( .A1(p[71]), .A2(c[71]), .Z(s[71]) );
  XOR2D0 C2234 ( .A1(p[72]), .A2(c[72]), .Z(s[72]) );
  XOR2D0 C2233 ( .A1(p[73]), .A2(c[73]), .Z(s[73]) );
  XOR2D0 C2232 ( .A1(p[74]), .A2(c[74]), .Z(s[74]) );
  XOR2D0 C2231 ( .A1(p[75]), .A2(c[75]), .Z(s[75]) );
  XOR2D0 C2230 ( .A1(p[76]), .A2(c[76]), .Z(s[76]) );
  XOR2D0 C2229 ( .A1(p[77]), .A2(c[77]), .Z(s[77]) );
  XOR2D0 C2228 ( .A1(p[78]), .A2(c[78]), .Z(s[78]) );
  XOR2D0 C2227 ( .A1(p[79]), .A2(c[79]), .Z(s[79]) );
  XOR2D0 C2226 ( .A1(p[80]), .A2(c[80]), .Z(s[80]) );
  XOR2D0 C2225 ( .A1(p[81]), .A2(c[81]), .Z(s[81]) );
  XOR2D0 C2224 ( .A1(p[82]), .A2(c[82]), .Z(s[82]) );
  XOR2D0 C2223 ( .A1(p[83]), .A2(c[83]), .Z(s[83]) );
  XOR2D0 C2222 ( .A1(p[84]), .A2(c[84]), .Z(s[84]) );
  XOR2D0 C2221 ( .A1(p[85]), .A2(c[85]), .Z(s[85]) );
  XOR2D0 C2220 ( .A1(p[86]), .A2(c[86]), .Z(s[86]) );
  XOR2D0 C2219 ( .A1(p[87]), .A2(c[87]), .Z(s[87]) );
  XOR2D0 C2218 ( .A1(p[88]), .A2(c[88]), .Z(s[88]) );
  XOR2D0 C2217 ( .A1(p[89]), .A2(c[89]), .Z(s[89]) );
  XOR2D0 C2216 ( .A1(p[90]), .A2(c[90]), .Z(s[90]) );
  XOR2D0 C2215 ( .A1(p[91]), .A2(c[91]), .Z(s[91]) );
  XOR2D0 C2214 ( .A1(p[92]), .A2(c[92]), .Z(s[92]) );
  XOR2D0 C2213 ( .A1(p[93]), .A2(c[93]), .Z(s[93]) );
  XOR2D0 C2212 ( .A1(p[94]), .A2(c[94]), .Z(s[94]) );
  XOR2D0 C2211 ( .A1(p[95]), .A2(c[95]), .Z(s[95]) );
  XOR2D0 C2210 ( .A1(p[96]), .A2(c[96]), .Z(s[96]) );
  XOR2D0 C2209 ( .A1(p[97]), .A2(c[97]), .Z(s[97]) );
  XOR2D0 C2208 ( .A1(p[98]), .A2(c[98]), .Z(s[98]) );
  XOR2D0 C2207 ( .A1(p[99]), .A2(c[99]), .Z(s[99]) );
  XOR2D0 C2206 ( .A1(p[100]), .A2(c[100]), .Z(s[100]) );
  XOR2D0 C2205 ( .A1(p[101]), .A2(c[101]), .Z(s[101]) );
  XOR2D0 C2204 ( .A1(p[102]), .A2(c[102]), .Z(s[102]) );
  XOR2D0 C2203 ( .A1(p[103]), .A2(c[103]), .Z(s[103]) );
  XOR2D0 C2202 ( .A1(p[104]), .A2(c[104]), .Z(s[104]) );
  XOR2D0 C2201 ( .A1(p[105]), .A2(c[105]), .Z(s[105]) );
  XOR2D0 C2200 ( .A1(p[106]), .A2(c[106]), .Z(s[106]) );
  XOR2D0 C2199 ( .A1(p[107]), .A2(c[107]), .Z(s[107]) );
  XOR2D0 C2198 ( .A1(p[108]), .A2(c[108]), .Z(s[108]) );
  XOR2D0 C2197 ( .A1(p[109]), .A2(c[109]), .Z(s[109]) );
  XOR2D0 C2196 ( .A1(p[110]), .A2(c[110]), .Z(s[110]) );
  XOR2D0 C2195 ( .A1(p[111]), .A2(c[111]), .Z(s[111]) );
  XOR2D0 C2194 ( .A1(p[112]), .A2(c[112]), .Z(s[112]) );
  XOR2D0 C2193 ( .A1(p[113]), .A2(c[113]), .Z(s[113]) );
  XOR2D0 C2192 ( .A1(p[114]), .A2(c[114]), .Z(s[114]) );
  XOR2D0 C2191 ( .A1(p[115]), .A2(c[115]), .Z(s[115]) );
  XOR2D0 C2190 ( .A1(p[116]), .A2(c[116]), .Z(s[116]) );
  XOR2D0 C2189 ( .A1(p[117]), .A2(c[117]), .Z(s[117]) );
  XOR2D0 C2188 ( .A1(p[118]), .A2(c[118]), .Z(s[118]) );
  XOR2D0 C2187 ( .A1(p[119]), .A2(c[119]), .Z(s[119]) );
  XOR2D0 C2186 ( .A1(p[120]), .A2(c[120]), .Z(s[120]) );
  XOR2D0 C2185 ( .A1(p[121]), .A2(c[121]), .Z(s[121]) );
  XOR2D0 C2184 ( .A1(p[122]), .A2(c[122]), .Z(s[122]) );
  XOR2D0 C2183 ( .A1(p[123]), .A2(c[123]), .Z(s[123]) );
  XOR2D0 C2182 ( .A1(p[124]), .A2(c[124]), .Z(s[124]) );
  XOR2D0 C2181 ( .A1(p[125]), .A2(c[125]), .Z(s[125]) );
  XOR2D0 C2180 ( .A1(p[126]), .A2(c[126]), .Z(s[126]) );
  XOR2D0 C2179 ( .A1(p[127]), .A2(c[127]), .Z(s[127]) );
  XOR2D0 C2178 ( .A1(p[128]), .A2(c[128]), .Z(s[128]) );
  XOR2D0 C2177 ( .A1(p[129]), .A2(c[129]), .Z(s[129]) );
  XOR2D0 C2176 ( .A1(p[130]), .A2(c[130]), .Z(s[130]) );
  XOR2D0 C2175 ( .A1(p[131]), .A2(c[131]), .Z(s[131]) );
  XOR2D0 C2174 ( .A1(p[132]), .A2(c[132]), .Z(s[132]) );
  XOR2D0 C2173 ( .A1(p[133]), .A2(c[133]), .Z(s[133]) );
  XOR2D0 C2172 ( .A1(p[134]), .A2(c[134]), .Z(s[134]) );
  XOR2D0 C2171 ( .A1(p[135]), .A2(c[135]), .Z(s[135]) );
  XOR2D0 C2170 ( .A1(p[136]), .A2(c[136]), .Z(s[136]) );
  XOR2D0 C2169 ( .A1(p[137]), .A2(c[137]), .Z(s[137]) );
  XOR2D0 C2168 ( .A1(p[138]), .A2(c[138]), .Z(s[138]) );
  XOR2D0 C2167 ( .A1(p[139]), .A2(c[139]), .Z(s[139]) );
  XOR2D0 C2166 ( .A1(p[140]), .A2(c[140]), .Z(s[140]) );
  XOR2D0 C2165 ( .A1(p[141]), .A2(c[141]), .Z(s[141]) );
  XOR2D0 C2164 ( .A1(p[142]), .A2(c[142]), .Z(s[142]) );
  XOR2D0 C2163 ( .A1(p[143]), .A2(c[143]), .Z(s[143]) );
  XOR2D0 C2162 ( .A1(p[144]), .A2(c[144]), .Z(s[144]) );
  XOR2D0 C2161 ( .A1(p[145]), .A2(c[145]), .Z(s[145]) );
  XOR2D0 C2160 ( .A1(p[146]), .A2(c[146]), .Z(s[146]) );
  XOR2D0 C2159 ( .A1(p[147]), .A2(c[147]), .Z(s[147]) );
  XOR2D0 C2158 ( .A1(p[148]), .A2(c[148]), .Z(s[148]) );
  XOR2D0 C2157 ( .A1(p[149]), .A2(c[149]), .Z(s[149]) );
  XOR2D0 C2156 ( .A1(p[150]), .A2(c[150]), .Z(s[150]) );
  XOR2D0 C2155 ( .A1(p[151]), .A2(c[151]), .Z(s[151]) );
  XOR2D0 C2154 ( .A1(p[152]), .A2(c[152]), .Z(s[152]) );
  XOR2D0 C2153 ( .A1(p[153]), .A2(c[153]), .Z(s[153]) );
  XOR2D0 C2152 ( .A1(p[154]), .A2(c[154]), .Z(s[154]) );
  XOR2D0 C2151 ( .A1(p[155]), .A2(c[155]), .Z(s[155]) );
  XOR2D0 C2150 ( .A1(p[156]), .A2(c[156]), .Z(s[156]) );
  XOR2D0 C2149 ( .A1(p[157]), .A2(c[157]), .Z(s[157]) );
  XOR2D0 C2148 ( .A1(p[158]), .A2(c[158]), .Z(s[158]) );
  XOR2D0 C2147 ( .A1(p[159]), .A2(c[159]), .Z(s[159]) );
  XOR2D0 C2146 ( .A1(p[160]), .A2(c[160]), .Z(s[160]) );
  XOR2D0 C2145 ( .A1(p[161]), .A2(c[161]), .Z(s[161]) );
  XOR2D0 C2144 ( .A1(p[162]), .A2(c[162]), .Z(s[162]) );
  XOR2D0 C2143 ( .A1(p[163]), .A2(c[163]), .Z(s[163]) );
  XOR2D0 C2142 ( .A1(p[164]), .A2(c[164]), .Z(s[164]) );
  XOR2D0 C2141 ( .A1(p[165]), .A2(c[165]), .Z(s[165]) );
  XOR2D0 C2140 ( .A1(p[166]), .A2(c[166]), .Z(s[166]) );
  XOR2D0 C2139 ( .A1(p[167]), .A2(c[167]), .Z(s[167]) );
  XOR2D0 C2138 ( .A1(p[168]), .A2(c[168]), .Z(s[168]) );
  XOR2D0 C2137 ( .A1(p[169]), .A2(c[169]), .Z(s[169]) );
  XOR2D0 C2136 ( .A1(p[170]), .A2(c[170]), .Z(s[170]) );
  XOR2D0 C2135 ( .A1(p[171]), .A2(c[171]), .Z(s[171]) );
  XOR2D0 C2134 ( .A1(p[172]), .A2(c[172]), .Z(s[172]) );
  XOR2D0 C2133 ( .A1(p[173]), .A2(c[173]), .Z(s[173]) );
  XOR2D0 C2132 ( .A1(p[174]), .A2(c[174]), .Z(s[174]) );
  XOR2D0 C2131 ( .A1(p[175]), .A2(c[175]), .Z(s[175]) );
  XOR2D0 C2130 ( .A1(p[176]), .A2(c[176]), .Z(s[176]) );
  XOR2D0 C2129 ( .A1(p[177]), .A2(c[177]), .Z(s[177]) );
  XOR2D0 C2128 ( .A1(p[178]), .A2(c[178]), .Z(s[178]) );
  XOR2D0 C2127 ( .A1(p[179]), .A2(c[179]), .Z(s[179]) );
  XOR2D0 C2126 ( .A1(p[180]), .A2(c[180]), .Z(s[180]) );
  XOR2D0 C2125 ( .A1(p[181]), .A2(c[181]), .Z(s[181]) );
  XOR2D0 C2124 ( .A1(p[182]), .A2(c[182]), .Z(s[182]) );
  XOR2D0 C2123 ( .A1(p[183]), .A2(c[183]), .Z(s[183]) );
  XOR2D0 C2122 ( .A1(p[184]), .A2(c[184]), .Z(s[184]) );
  XOR2D0 C2121 ( .A1(p[185]), .A2(c[185]), .Z(s[185]) );
  XOR2D0 C2120 ( .A1(p[186]), .A2(c[186]), .Z(s[186]) );
  XOR2D0 C2119 ( .A1(p[187]), .A2(c[187]), .Z(s[187]) );
  XOR2D0 C2118 ( .A1(p[188]), .A2(c[188]), .Z(s[188]) );
  XOR2D0 C2117 ( .A1(p[189]), .A2(c[189]), .Z(s[189]) );
  XOR2D0 C2116 ( .A1(p[190]), .A2(c[190]), .Z(s[190]) );
  XOR2D0 C2115 ( .A1(p[191]), .A2(c[191]), .Z(s[191]) );
  XOR2D0 C2114 ( .A1(p[192]), .A2(c[192]), .Z(s[192]) );
  XOR2D0 C2113 ( .A1(p[193]), .A2(c[193]), .Z(s[193]) );
  XOR2D0 C2112 ( .A1(p[194]), .A2(c[194]), .Z(s[194]) );
  XOR2D0 C2111 ( .A1(p[195]), .A2(c[195]), .Z(s[195]) );
  XOR2D0 C2110 ( .A1(p[196]), .A2(c[196]), .Z(s[196]) );
  XOR2D0 C2109 ( .A1(p[197]), .A2(c[197]), .Z(s[197]) );
  XOR2D0 C2108 ( .A1(p[198]), .A2(c[198]), .Z(s[198]) );
  XOR2D0 C2107 ( .A1(p[199]), .A2(c[199]), .Z(s[199]) );
  XOR2D0 C2106 ( .A1(p[200]), .A2(c[200]), .Z(s[200]) );
  XOR2D0 C2105 ( .A1(p[201]), .A2(c[201]), .Z(s[201]) );
  XOR2D0 C2104 ( .A1(p[202]), .A2(c[202]), .Z(s[202]) );
  XOR2D0 C2103 ( .A1(p[203]), .A2(c[203]), .Z(s[203]) );
  XOR2D0 C2102 ( .A1(p[204]), .A2(c[204]), .Z(s[204]) );
  XOR2D0 C2101 ( .A1(p[205]), .A2(c[205]), .Z(s[205]) );
  XOR2D0 C2100 ( .A1(p[206]), .A2(c[206]), .Z(s[206]) );
  XOR2D0 C2099 ( .A1(p[207]), .A2(c[207]), .Z(s[207]) );
  XOR2D0 C2098 ( .A1(p[208]), .A2(c[208]), .Z(s[208]) );
  XOR2D0 C2097 ( .A1(p[209]), .A2(c[209]), .Z(s[209]) );
  XOR2D0 C2096 ( .A1(p[210]), .A2(c[210]), .Z(s[210]) );
  XOR2D0 C2095 ( .A1(p[211]), .A2(c[211]), .Z(s[211]) );
  XOR2D0 C2094 ( .A1(p[212]), .A2(c[212]), .Z(s[212]) );
  XOR2D0 C2093 ( .A1(p[213]), .A2(c[213]), .Z(s[213]) );
  XOR2D0 C2092 ( .A1(p[214]), .A2(c[214]), .Z(s[214]) );
  XOR2D0 C2091 ( .A1(p[215]), .A2(c[215]), .Z(s[215]) );
  XOR2D0 C2090 ( .A1(p[216]), .A2(c[216]), .Z(s[216]) );
  XOR2D0 C2089 ( .A1(p[217]), .A2(c[217]), .Z(s[217]) );
  XOR2D0 C2088 ( .A1(p[218]), .A2(c[218]), .Z(s[218]) );
  XOR2D0 C2087 ( .A1(p[219]), .A2(c[219]), .Z(s[219]) );
  XOR2D0 C2086 ( .A1(p[220]), .A2(c[220]), .Z(s[220]) );
  XOR2D0 C2085 ( .A1(p[221]), .A2(c[221]), .Z(s[221]) );
  XOR2D0 C2084 ( .A1(p[222]), .A2(c[222]), .Z(s[222]) );
  XOR2D0 C2083 ( .A1(p[223]), .A2(c[223]), .Z(s[223]) );
  XOR2D0 C2082 ( .A1(p[224]), .A2(c[224]), .Z(s[224]) );
  XOR2D0 C2081 ( .A1(p[225]), .A2(c[225]), .Z(s[225]) );
  XOR2D0 C2080 ( .A1(p[226]), .A2(c[226]), .Z(s[226]) );
  XOR2D0 C2079 ( .A1(p[227]), .A2(c[227]), .Z(s[227]) );
  XOR2D0 C2078 ( .A1(p[228]), .A2(c[228]), .Z(s[228]) );
  XOR2D0 C2077 ( .A1(p[229]), .A2(c[229]), .Z(s[229]) );
  XOR2D0 C2076 ( .A1(p[230]), .A2(c[230]), .Z(s[230]) );
  XOR2D0 C2075 ( .A1(p[231]), .A2(c[231]), .Z(s[231]) );
  XOR2D0 C2074 ( .A1(p[232]), .A2(c[232]), .Z(s[232]) );
  XOR2D0 C2073 ( .A1(p[233]), .A2(c[233]), .Z(s[233]) );
  XOR2D0 C2072 ( .A1(p[234]), .A2(c[234]), .Z(s[234]) );
  XOR2D0 C2071 ( .A1(p[235]), .A2(c[235]), .Z(s[235]) );
  XOR2D0 C2070 ( .A1(p[236]), .A2(c[236]), .Z(s[236]) );
  XOR2D0 C2069 ( .A1(p[237]), .A2(c[237]), .Z(s[237]) );
  XOR2D0 C2068 ( .A1(p[238]), .A2(c[238]), .Z(s[238]) );
  XOR2D0 C2067 ( .A1(p[239]), .A2(c[239]), .Z(s[239]) );
  XOR2D0 C2066 ( .A1(p[240]), .A2(c[240]), .Z(s[240]) );
  XOR2D0 C2065 ( .A1(p[241]), .A2(c[241]), .Z(s[241]) );
  XOR2D0 C2064 ( .A1(p[242]), .A2(c[242]), .Z(s[242]) );
  XOR2D0 C2063 ( .A1(p[243]), .A2(c[243]), .Z(s[243]) );
  XOR2D0 C2062 ( .A1(p[244]), .A2(c[244]), .Z(s[244]) );
  XOR2D0 C2061 ( .A1(p[245]), .A2(c[245]), .Z(s[245]) );
  XOR2D0 C2060 ( .A1(p[246]), .A2(c[246]), .Z(s[246]) );
  XOR2D0 C2059 ( .A1(p[247]), .A2(c[247]), .Z(s[247]) );
  XOR2D0 C2058 ( .A1(p[248]), .A2(c[248]), .Z(s[248]) );
  XOR2D0 C2057 ( .A1(p[249]), .A2(c[249]), .Z(s[249]) );
  XOR2D0 C2056 ( .A1(p[250]), .A2(c[250]), .Z(s[250]) );
  XOR2D0 C2055 ( .A1(p[251]), .A2(c[251]), .Z(s[251]) );
  XOR2D0 C2054 ( .A1(p[252]), .A2(c[252]), .Z(s[252]) );
  XOR2D0 C2053 ( .A1(p[253]), .A2(c[253]), .Z(s[253]) );
  XOR2D0 C2052 ( .A1(p[254]), .A2(c[254]), .Z(s[254]) );
  XOR2D0 C2051 ( .A1(p[255]), .A2(c[255]), .Z(s[255]) );
  AN2D0 C2050 ( .A1(p[254]), .A2(c[254]), .Z(N254) );
  OR2D0 C2049 ( .A1(g[254]), .A2(N254), .Z(c[255]) );
  AN2D0 C2048 ( .A1(p[253]), .A2(c[253]), .Z(N253) );
  OR2D0 C2047 ( .A1(g[253]), .A2(N253), .Z(c[254]) );
  AN2D0 C2046 ( .A1(p[252]), .A2(c[252]), .Z(N252) );
  OR2D0 C2045 ( .A1(g[252]), .A2(N252), .Z(c[253]) );
  AN2D0 C2044 ( .A1(p[251]), .A2(c[251]), .Z(N251) );
  OR2D0 C2043 ( .A1(g[251]), .A2(N251), .Z(c[252]) );
  AN2D0 C2042 ( .A1(p[250]), .A2(c[250]), .Z(N250) );
  OR2D0 C2041 ( .A1(g[250]), .A2(N250), .Z(c[251]) );
  AN2D0 C2040 ( .A1(p[249]), .A2(c[249]), .Z(N249) );
  OR2D0 C2039 ( .A1(g[249]), .A2(N249), .Z(c[250]) );
  AN2D0 C2038 ( .A1(p[248]), .A2(c[248]), .Z(N248) );
  OR2D0 C2037 ( .A1(g[248]), .A2(N248), .Z(c[249]) );
  AN2D0 C2036 ( .A1(p[247]), .A2(c[247]), .Z(N247) );
  OR2D0 C2035 ( .A1(g[247]), .A2(N247), .Z(c[248]) );
  AN2D0 C2034 ( .A1(p[246]), .A2(c[246]), .Z(N246) );
  OR2D0 C2033 ( .A1(g[246]), .A2(N246), .Z(c[247]) );
  AN2D0 C2032 ( .A1(p[245]), .A2(c[245]), .Z(N245) );
  OR2D0 C2031 ( .A1(g[245]), .A2(N245), .Z(c[246]) );
  AN2D0 C2030 ( .A1(p[244]), .A2(c[244]), .Z(N244) );
  OR2D0 C2029 ( .A1(g[244]), .A2(N244), .Z(c[245]) );
  AN2D0 C2028 ( .A1(p[243]), .A2(c[243]), .Z(N243) );
  OR2D0 C2027 ( .A1(g[243]), .A2(N243), .Z(c[244]) );
  AN2D0 C2026 ( .A1(p[242]), .A2(c[242]), .Z(N242) );
  OR2D0 C2025 ( .A1(g[242]), .A2(N242), .Z(c[243]) );
  AN2D0 C2024 ( .A1(p[241]), .A2(c[241]), .Z(N241) );
  OR2D0 C2023 ( .A1(g[241]), .A2(N241), .Z(c[242]) );
  AN2D0 C2022 ( .A1(p[240]), .A2(c[240]), .Z(N240) );
  OR2D0 C2021 ( .A1(g[240]), .A2(N240), .Z(c[241]) );
  AN2D0 C2020 ( .A1(p[239]), .A2(c[239]), .Z(N239) );
  OR2D0 C2019 ( .A1(g[239]), .A2(N239), .Z(c[240]) );
  AN2D0 C2018 ( .A1(p[238]), .A2(c[238]), .Z(N238) );
  OR2D0 C2017 ( .A1(g[238]), .A2(N238), .Z(c[239]) );
  AN2D0 C2016 ( .A1(p[237]), .A2(c[237]), .Z(N237) );
  OR2D0 C2015 ( .A1(g[237]), .A2(N237), .Z(c[238]) );
  AN2D0 C2014 ( .A1(p[236]), .A2(c[236]), .Z(N236) );
  OR2D0 C2013 ( .A1(g[236]), .A2(N236), .Z(c[237]) );
  AN2D0 C2012 ( .A1(p[235]), .A2(c[235]), .Z(N235) );
  OR2D0 C2011 ( .A1(g[235]), .A2(N235), .Z(c[236]) );
  AN2D0 C2010 ( .A1(p[234]), .A2(c[234]), .Z(N234) );
  OR2D0 C2009 ( .A1(g[234]), .A2(N234), .Z(c[235]) );
  AN2D0 C2008 ( .A1(p[233]), .A2(c[233]), .Z(N233) );
  OR2D0 C2007 ( .A1(g[233]), .A2(N233), .Z(c[234]) );
  AN2D0 C2006 ( .A1(p[232]), .A2(c[232]), .Z(N232) );
  OR2D0 C2005 ( .A1(g[232]), .A2(N232), .Z(c[233]) );
  AN2D0 C2004 ( .A1(p[231]), .A2(c[231]), .Z(N231) );
  OR2D0 C2003 ( .A1(g[231]), .A2(N231), .Z(c[232]) );
  AN2D0 C2002 ( .A1(p[230]), .A2(c[230]), .Z(N230) );
  OR2D0 C2001 ( .A1(g[230]), .A2(N230), .Z(c[231]) );
  AN2D0 C2000 ( .A1(p[229]), .A2(c[229]), .Z(N229) );
  OR2D0 C1999 ( .A1(g[229]), .A2(N229), .Z(c[230]) );
  AN2D0 C1998 ( .A1(p[228]), .A2(c[228]), .Z(N228) );
  OR2D0 C1997 ( .A1(g[228]), .A2(N228), .Z(c[229]) );
  AN2D0 C1996 ( .A1(p[227]), .A2(c[227]), .Z(N227) );
  OR2D0 C1995 ( .A1(g[227]), .A2(N227), .Z(c[228]) );
  AN2D0 C1994 ( .A1(p[226]), .A2(c[226]), .Z(N226) );
  OR2D0 C1993 ( .A1(g[226]), .A2(N226), .Z(c[227]) );
  AN2D0 C1992 ( .A1(p[225]), .A2(c[225]), .Z(N225) );
  OR2D0 C1991 ( .A1(g[225]), .A2(N225), .Z(c[226]) );
  AN2D0 C1990 ( .A1(p[224]), .A2(c[224]), .Z(N224) );
  OR2D0 C1989 ( .A1(g[224]), .A2(N224), .Z(c[225]) );
  AN2D0 C1988 ( .A1(p[223]), .A2(c[223]), .Z(N223) );
  OR2D0 C1987 ( .A1(g[223]), .A2(N223), .Z(c[224]) );
  AN2D0 C1986 ( .A1(p[222]), .A2(c[222]), .Z(N222) );
  OR2D0 C1985 ( .A1(g[222]), .A2(N222), .Z(c[223]) );
  AN2D0 C1984 ( .A1(p[221]), .A2(c[221]), .Z(N221) );
  OR2D0 C1983 ( .A1(g[221]), .A2(N221), .Z(c[222]) );
  AN2D0 C1982 ( .A1(p[220]), .A2(c[220]), .Z(N220) );
  OR2D0 C1981 ( .A1(g[220]), .A2(N220), .Z(c[221]) );
  AN2D0 C1980 ( .A1(p[219]), .A2(c[219]), .Z(N219) );
  OR2D0 C1979 ( .A1(g[219]), .A2(N219), .Z(c[220]) );
  AN2D0 C1978 ( .A1(p[218]), .A2(c[218]), .Z(N218) );
  OR2D0 C1977 ( .A1(g[218]), .A2(N218), .Z(c[219]) );
  AN2D0 C1976 ( .A1(p[217]), .A2(c[217]), .Z(N217) );
  OR2D0 C1975 ( .A1(g[217]), .A2(N217), .Z(c[218]) );
  AN2D0 C1974 ( .A1(p[216]), .A2(c[216]), .Z(N216) );
  OR2D0 C1973 ( .A1(g[216]), .A2(N216), .Z(c[217]) );
  AN2D0 C1972 ( .A1(p[215]), .A2(c[215]), .Z(N215) );
  OR2D0 C1971 ( .A1(g[215]), .A2(N215), .Z(c[216]) );
  AN2D0 C1970 ( .A1(p[214]), .A2(c[214]), .Z(N214) );
  OR2D0 C1969 ( .A1(g[214]), .A2(N214), .Z(c[215]) );
  AN2D0 C1968 ( .A1(p[213]), .A2(c[213]), .Z(N213) );
  OR2D0 C1967 ( .A1(g[213]), .A2(N213), .Z(c[214]) );
  AN2D0 C1966 ( .A1(p[212]), .A2(c[212]), .Z(N212) );
  OR2D0 C1965 ( .A1(g[212]), .A2(N212), .Z(c[213]) );
  AN2D0 C1964 ( .A1(p[211]), .A2(c[211]), .Z(N211) );
  OR2D0 C1963 ( .A1(g[211]), .A2(N211), .Z(c[212]) );
  AN2D0 C1962 ( .A1(p[210]), .A2(c[210]), .Z(N210) );
  OR2D0 C1961 ( .A1(g[210]), .A2(N210), .Z(c[211]) );
  AN2D0 C1960 ( .A1(p[209]), .A2(c[209]), .Z(N209) );
  OR2D0 C1959 ( .A1(g[209]), .A2(N209), .Z(c[210]) );
  AN2D0 C1958 ( .A1(p[208]), .A2(c[208]), .Z(N208) );
  OR2D0 C1957 ( .A1(g[208]), .A2(N208), .Z(c[209]) );
  AN2D0 C1956 ( .A1(p[207]), .A2(c[207]), .Z(N207) );
  OR2D0 C1955 ( .A1(g[207]), .A2(N207), .Z(c[208]) );
  AN2D0 C1954 ( .A1(p[206]), .A2(c[206]), .Z(N206) );
  OR2D0 C1953 ( .A1(g[206]), .A2(N206), .Z(c[207]) );
  AN2D0 C1952 ( .A1(p[205]), .A2(c[205]), .Z(N205) );
  OR2D0 C1951 ( .A1(g[205]), .A2(N205), .Z(c[206]) );
  AN2D0 C1950 ( .A1(p[204]), .A2(c[204]), .Z(N204) );
  OR2D0 C1949 ( .A1(g[204]), .A2(N204), .Z(c[205]) );
  AN2D0 C1948 ( .A1(p[203]), .A2(c[203]), .Z(N203) );
  OR2D0 C1947 ( .A1(g[203]), .A2(N203), .Z(c[204]) );
  AN2D0 C1946 ( .A1(p[202]), .A2(c[202]), .Z(N202) );
  OR2D0 C1945 ( .A1(g[202]), .A2(N202), .Z(c[203]) );
  AN2D0 C1944 ( .A1(p[201]), .A2(c[201]), .Z(N201) );
  OR2D0 C1943 ( .A1(g[201]), .A2(N201), .Z(c[202]) );
  AN2D0 C1942 ( .A1(p[200]), .A2(c[200]), .Z(N200) );
  OR2D0 C1941 ( .A1(g[200]), .A2(N200), .Z(c[201]) );
  AN2D0 C1940 ( .A1(p[199]), .A2(c[199]), .Z(N199) );
  OR2D0 C1939 ( .A1(g[199]), .A2(N199), .Z(c[200]) );
  AN2D0 C1938 ( .A1(p[198]), .A2(c[198]), .Z(N198) );
  OR2D0 C1937 ( .A1(g[198]), .A2(N198), .Z(c[199]) );
  AN2D0 C1936 ( .A1(p[197]), .A2(c[197]), .Z(N197) );
  OR2D0 C1935 ( .A1(g[197]), .A2(N197), .Z(c[198]) );
  AN2D0 C1934 ( .A1(p[196]), .A2(c[196]), .Z(N196) );
  OR2D0 C1933 ( .A1(g[196]), .A2(N196), .Z(c[197]) );
  AN2D0 C1932 ( .A1(p[195]), .A2(c[195]), .Z(N195) );
  OR2D0 C1931 ( .A1(g[195]), .A2(N195), .Z(c[196]) );
  AN2D0 C1930 ( .A1(p[194]), .A2(c[194]), .Z(N194) );
  OR2D0 C1929 ( .A1(g[194]), .A2(N194), .Z(c[195]) );
  AN2D0 C1928 ( .A1(p[193]), .A2(c[193]), .Z(N193) );
  OR2D0 C1927 ( .A1(g[193]), .A2(N193), .Z(c[194]) );
  AN2D0 C1926 ( .A1(p[192]), .A2(c[192]), .Z(N192) );
  OR2D0 C1925 ( .A1(g[192]), .A2(N192), .Z(c[193]) );
  AN2D0 C1924 ( .A1(p[191]), .A2(c[191]), .Z(N191) );
  OR2D0 C1923 ( .A1(g[191]), .A2(N191), .Z(c[192]) );
  AN2D0 C1922 ( .A1(p[190]), .A2(c[190]), .Z(N190) );
  OR2D0 C1921 ( .A1(g[190]), .A2(N190), .Z(c[191]) );
  AN2D0 C1920 ( .A1(p[189]), .A2(c[189]), .Z(N189) );
  OR2D0 C1919 ( .A1(g[189]), .A2(N189), .Z(c[190]) );
  AN2D0 C1918 ( .A1(p[188]), .A2(c[188]), .Z(N188) );
  OR2D0 C1917 ( .A1(g[188]), .A2(N188), .Z(c[189]) );
  AN2D0 C1916 ( .A1(p[187]), .A2(c[187]), .Z(N187) );
  OR2D0 C1915 ( .A1(g[187]), .A2(N187), .Z(c[188]) );
  AN2D0 C1914 ( .A1(p[186]), .A2(c[186]), .Z(N186) );
  OR2D0 C1913 ( .A1(g[186]), .A2(N186), .Z(c[187]) );
  AN2D0 C1912 ( .A1(p[185]), .A2(c[185]), .Z(N185) );
  OR2D0 C1911 ( .A1(g[185]), .A2(N185), .Z(c[186]) );
  AN2D0 C1910 ( .A1(p[184]), .A2(c[184]), .Z(N184) );
  OR2D0 C1909 ( .A1(g[184]), .A2(N184), .Z(c[185]) );
  AN2D0 C1908 ( .A1(p[183]), .A2(c[183]), .Z(N183) );
  OR2D0 C1907 ( .A1(g[183]), .A2(N183), .Z(c[184]) );
  AN2D0 C1906 ( .A1(p[182]), .A2(c[182]), .Z(N182) );
  OR2D0 C1905 ( .A1(g[182]), .A2(N182), .Z(c[183]) );
  AN2D0 C1904 ( .A1(p[181]), .A2(c[181]), .Z(N181) );
  OR2D0 C1903 ( .A1(g[181]), .A2(N181), .Z(c[182]) );
  AN2D0 C1902 ( .A1(p[180]), .A2(c[180]), .Z(N180) );
  OR2D0 C1901 ( .A1(g[180]), .A2(N180), .Z(c[181]) );
  AN2D0 C1900 ( .A1(p[179]), .A2(c[179]), .Z(N179) );
  OR2D0 C1899 ( .A1(g[179]), .A2(N179), .Z(c[180]) );
  AN2D0 C1898 ( .A1(p[178]), .A2(c[178]), .Z(N178) );
  OR2D0 C1897 ( .A1(g[178]), .A2(N178), .Z(c[179]) );
  AN2D0 C1896 ( .A1(p[177]), .A2(c[177]), .Z(N177) );
  OR2D0 C1895 ( .A1(g[177]), .A2(N177), .Z(c[178]) );
  AN2D0 C1894 ( .A1(p[176]), .A2(c[176]), .Z(N176) );
  OR2D0 C1893 ( .A1(g[176]), .A2(N176), .Z(c[177]) );
  AN2D0 C1892 ( .A1(p[175]), .A2(c[175]), .Z(N175) );
  OR2D0 C1891 ( .A1(g[175]), .A2(N175), .Z(c[176]) );
  AN2D0 C1890 ( .A1(p[174]), .A2(c[174]), .Z(N174) );
  OR2D0 C1889 ( .A1(g[174]), .A2(N174), .Z(c[175]) );
  AN2D0 C1888 ( .A1(p[173]), .A2(c[173]), .Z(N173) );
  OR2D0 C1887 ( .A1(g[173]), .A2(N173), .Z(c[174]) );
  AN2D0 C1886 ( .A1(p[172]), .A2(c[172]), .Z(N172) );
  OR2D0 C1885 ( .A1(g[172]), .A2(N172), .Z(c[173]) );
  AN2D0 C1884 ( .A1(p[171]), .A2(c[171]), .Z(N171) );
  OR2D0 C1883 ( .A1(g[171]), .A2(N171), .Z(c[172]) );
  AN2D0 C1882 ( .A1(p[170]), .A2(c[170]), .Z(N170) );
  OR2D0 C1881 ( .A1(g[170]), .A2(N170), .Z(c[171]) );
  AN2D0 C1880 ( .A1(p[169]), .A2(c[169]), .Z(N169) );
  OR2D0 C1879 ( .A1(g[169]), .A2(N169), .Z(c[170]) );
  AN2D0 C1878 ( .A1(p[168]), .A2(c[168]), .Z(N168) );
  OR2D0 C1877 ( .A1(g[168]), .A2(N168), .Z(c[169]) );
  AN2D0 C1876 ( .A1(p[167]), .A2(c[167]), .Z(N167) );
  OR2D0 C1875 ( .A1(g[167]), .A2(N167), .Z(c[168]) );
  AN2D0 C1874 ( .A1(p[166]), .A2(c[166]), .Z(N166) );
  OR2D0 C1873 ( .A1(g[166]), .A2(N166), .Z(c[167]) );
  AN2D0 C1872 ( .A1(p[165]), .A2(c[165]), .Z(N165) );
  OR2D0 C1871 ( .A1(g[165]), .A2(N165), .Z(c[166]) );
  AN2D0 C1870 ( .A1(p[164]), .A2(c[164]), .Z(N164) );
  OR2D0 C1869 ( .A1(g[164]), .A2(N164), .Z(c[165]) );
  AN2D0 C1868 ( .A1(p[163]), .A2(c[163]), .Z(N163) );
  OR2D0 C1867 ( .A1(g[163]), .A2(N163), .Z(c[164]) );
  AN2D0 C1866 ( .A1(p[162]), .A2(c[162]), .Z(N162) );
  OR2D0 C1865 ( .A1(g[162]), .A2(N162), .Z(c[163]) );
  AN2D0 C1864 ( .A1(p[161]), .A2(c[161]), .Z(N161) );
  OR2D0 C1863 ( .A1(g[161]), .A2(N161), .Z(c[162]) );
  AN2D0 C1862 ( .A1(p[160]), .A2(c[160]), .Z(N160) );
  OR2D0 C1861 ( .A1(g[160]), .A2(N160), .Z(c[161]) );
  AN2D0 C1860 ( .A1(p[159]), .A2(c[159]), .Z(N159) );
  OR2D0 C1859 ( .A1(g[159]), .A2(N159), .Z(c[160]) );
  AN2D0 C1858 ( .A1(p[158]), .A2(c[158]), .Z(N158) );
  OR2D0 C1857 ( .A1(g[158]), .A2(N158), .Z(c[159]) );
  AN2D0 C1856 ( .A1(p[157]), .A2(c[157]), .Z(N157) );
  OR2D0 C1855 ( .A1(g[157]), .A2(N157), .Z(c[158]) );
  AN2D0 C1854 ( .A1(p[156]), .A2(c[156]), .Z(N156) );
  OR2D0 C1853 ( .A1(g[156]), .A2(N156), .Z(c[157]) );
  AN2D0 C1852 ( .A1(p[155]), .A2(c[155]), .Z(N155) );
  OR2D0 C1851 ( .A1(g[155]), .A2(N155), .Z(c[156]) );
  AN2D0 C1850 ( .A1(p[154]), .A2(c[154]), .Z(N154) );
  OR2D0 C1849 ( .A1(g[154]), .A2(N154), .Z(c[155]) );
  AN2D0 C1848 ( .A1(p[153]), .A2(c[153]), .Z(N153) );
  OR2D0 C1847 ( .A1(g[153]), .A2(N153), .Z(c[154]) );
  AN2D0 C1846 ( .A1(p[152]), .A2(c[152]), .Z(N152) );
  OR2D0 C1845 ( .A1(g[152]), .A2(N152), .Z(c[153]) );
  AN2D0 C1844 ( .A1(p[151]), .A2(c[151]), .Z(N151) );
  OR2D0 C1843 ( .A1(g[151]), .A2(N151), .Z(c[152]) );
  AN2D0 C1842 ( .A1(p[150]), .A2(c[150]), .Z(N150) );
  OR2D0 C1841 ( .A1(g[150]), .A2(N150), .Z(c[151]) );
  AN2D0 C1840 ( .A1(p[149]), .A2(c[149]), .Z(N149) );
  OR2D0 C1839 ( .A1(g[149]), .A2(N149), .Z(c[150]) );
  AN2D0 C1838 ( .A1(p[148]), .A2(c[148]), .Z(N148) );
  OR2D0 C1837 ( .A1(g[148]), .A2(N148), .Z(c[149]) );
  AN2D0 C1836 ( .A1(p[147]), .A2(c[147]), .Z(N147) );
  OR2D0 C1835 ( .A1(g[147]), .A2(N147), .Z(c[148]) );
  AN2D0 C1834 ( .A1(p[146]), .A2(c[146]), .Z(N146) );
  OR2D0 C1833 ( .A1(g[146]), .A2(N146), .Z(c[147]) );
  AN2D0 C1832 ( .A1(p[145]), .A2(c[145]), .Z(N145) );
  OR2D0 C1831 ( .A1(g[145]), .A2(N145), .Z(c[146]) );
  AN2D0 C1830 ( .A1(p[144]), .A2(c[144]), .Z(N144) );
  OR2D0 C1829 ( .A1(g[144]), .A2(N144), .Z(c[145]) );
  AN2D0 C1828 ( .A1(p[143]), .A2(c[143]), .Z(N143) );
  OR2D0 C1827 ( .A1(g[143]), .A2(N143), .Z(c[144]) );
  AN2D0 C1826 ( .A1(p[142]), .A2(c[142]), .Z(N142) );
  OR2D0 C1825 ( .A1(g[142]), .A2(N142), .Z(c[143]) );
  AN2D0 C1824 ( .A1(p[141]), .A2(c[141]), .Z(N141) );
  OR2D0 C1823 ( .A1(g[141]), .A2(N141), .Z(c[142]) );
  AN2D0 C1822 ( .A1(p[140]), .A2(c[140]), .Z(N140) );
  OR2D0 C1821 ( .A1(g[140]), .A2(N140), .Z(c[141]) );
  AN2D0 C1820 ( .A1(p[139]), .A2(c[139]), .Z(N139) );
  OR2D0 C1819 ( .A1(g[139]), .A2(N139), .Z(c[140]) );
  AN2D0 C1818 ( .A1(p[138]), .A2(c[138]), .Z(N138) );
  OR2D0 C1817 ( .A1(g[138]), .A2(N138), .Z(c[139]) );
  AN2D0 C1816 ( .A1(p[137]), .A2(c[137]), .Z(N137) );
  OR2D0 C1815 ( .A1(g[137]), .A2(N137), .Z(c[138]) );
  AN2D0 C1814 ( .A1(p[136]), .A2(c[136]), .Z(N136) );
  OR2D0 C1813 ( .A1(g[136]), .A2(N136), .Z(c[137]) );
  AN2D0 C1812 ( .A1(p[135]), .A2(c[135]), .Z(N135) );
  OR2D0 C1811 ( .A1(g[135]), .A2(N135), .Z(c[136]) );
  AN2D0 C1810 ( .A1(p[134]), .A2(c[134]), .Z(N134) );
  OR2D0 C1809 ( .A1(g[134]), .A2(N134), .Z(c[135]) );
  AN2D0 C1808 ( .A1(p[133]), .A2(c[133]), .Z(N133) );
  OR2D0 C1807 ( .A1(g[133]), .A2(N133), .Z(c[134]) );
  AN2D0 C1806 ( .A1(p[132]), .A2(c[132]), .Z(N132) );
  OR2D0 C1805 ( .A1(g[132]), .A2(N132), .Z(c[133]) );
  AN2D0 C1804 ( .A1(p[131]), .A2(c[131]), .Z(N131) );
  OR2D0 C1803 ( .A1(g[131]), .A2(N131), .Z(c[132]) );
  AN2D0 C1802 ( .A1(p[130]), .A2(c[130]), .Z(N130) );
  OR2D0 C1801 ( .A1(g[130]), .A2(N130), .Z(c[131]) );
  AN2D0 C1800 ( .A1(p[129]), .A2(c[129]), .Z(N129) );
  OR2D0 C1799 ( .A1(g[129]), .A2(N129), .Z(c[130]) );
  AN2D0 C1798 ( .A1(p[128]), .A2(c[128]), .Z(N128) );
  OR2D0 C1797 ( .A1(g[128]), .A2(N128), .Z(c[129]) );
  AN2D0 C1796 ( .A1(p[127]), .A2(c[127]), .Z(N127) );
  OR2D0 C1795 ( .A1(g[127]), .A2(N127), .Z(c[128]) );
  AN2D0 C1794 ( .A1(p[126]), .A2(c[126]), .Z(N126) );
  OR2D0 C1793 ( .A1(g[126]), .A2(N126), .Z(c[127]) );
  AN2D0 C1792 ( .A1(p[125]), .A2(c[125]), .Z(N125) );
  OR2D0 C1791 ( .A1(g[125]), .A2(N125), .Z(c[126]) );
  AN2D0 C1790 ( .A1(p[124]), .A2(c[124]), .Z(N124) );
  OR2D0 C1789 ( .A1(g[124]), .A2(N124), .Z(c[125]) );
  AN2D0 C1788 ( .A1(p[123]), .A2(c[123]), .Z(N123) );
  OR2D0 C1787 ( .A1(g[123]), .A2(N123), .Z(c[124]) );
  AN2D0 C1786 ( .A1(p[122]), .A2(c[122]), .Z(N122) );
  OR2D0 C1785 ( .A1(g[122]), .A2(N122), .Z(c[123]) );
  AN2D0 C1784 ( .A1(p[121]), .A2(c[121]), .Z(N121) );
  OR2D0 C1783 ( .A1(g[121]), .A2(N121), .Z(c[122]) );
  AN2D0 C1782 ( .A1(p[120]), .A2(c[120]), .Z(N120) );
  OR2D0 C1781 ( .A1(g[120]), .A2(N120), .Z(c[121]) );
  AN2D0 C1780 ( .A1(p[119]), .A2(c[119]), .Z(N119) );
  OR2D0 C1779 ( .A1(g[119]), .A2(N119), .Z(c[120]) );
  AN2D0 C1778 ( .A1(p[118]), .A2(c[118]), .Z(N118) );
  OR2D0 C1777 ( .A1(g[118]), .A2(N118), .Z(c[119]) );
  AN2D0 C1776 ( .A1(p[117]), .A2(c[117]), .Z(N117) );
  OR2D0 C1775 ( .A1(g[117]), .A2(N117), .Z(c[118]) );
  AN2D0 C1774 ( .A1(p[116]), .A2(c[116]), .Z(N116) );
  OR2D0 C1773 ( .A1(g[116]), .A2(N116), .Z(c[117]) );
  AN2D0 C1772 ( .A1(p[115]), .A2(c[115]), .Z(N115) );
  OR2D0 C1771 ( .A1(g[115]), .A2(N115), .Z(c[116]) );
  AN2D0 C1770 ( .A1(p[114]), .A2(c[114]), .Z(N114) );
  OR2D0 C1769 ( .A1(g[114]), .A2(N114), .Z(c[115]) );
  AN2D0 C1768 ( .A1(p[113]), .A2(c[113]), .Z(N113) );
  OR2D0 C1767 ( .A1(g[113]), .A2(N113), .Z(c[114]) );
  AN2D0 C1766 ( .A1(p[112]), .A2(c[112]), .Z(N112) );
  OR2D0 C1765 ( .A1(g[112]), .A2(N112), .Z(c[113]) );
  AN2D0 C1764 ( .A1(p[111]), .A2(c[111]), .Z(N111) );
  OR2D0 C1763 ( .A1(g[111]), .A2(N111), .Z(c[112]) );
  AN2D0 C1762 ( .A1(p[110]), .A2(c[110]), .Z(N110) );
  OR2D0 C1761 ( .A1(g[110]), .A2(N110), .Z(c[111]) );
  AN2D0 C1760 ( .A1(p[109]), .A2(c[109]), .Z(N109) );
  OR2D0 C1759 ( .A1(g[109]), .A2(N109), .Z(c[110]) );
  AN2D0 C1758 ( .A1(p[108]), .A2(c[108]), .Z(N108) );
  OR2D0 C1757 ( .A1(g[108]), .A2(N108), .Z(c[109]) );
  AN2D0 C1756 ( .A1(p[107]), .A2(c[107]), .Z(N107) );
  OR2D0 C1755 ( .A1(g[107]), .A2(N107), .Z(c[108]) );
  AN2D0 C1754 ( .A1(p[106]), .A2(c[106]), .Z(N106) );
  OR2D0 C1753 ( .A1(g[106]), .A2(N106), .Z(c[107]) );
  AN2D0 C1752 ( .A1(p[105]), .A2(c[105]), .Z(N105) );
  OR2D0 C1751 ( .A1(g[105]), .A2(N105), .Z(c[106]) );
  AN2D0 C1750 ( .A1(p[104]), .A2(c[104]), .Z(N104) );
  OR2D0 C1749 ( .A1(g[104]), .A2(N104), .Z(c[105]) );
  AN2D0 C1748 ( .A1(p[103]), .A2(c[103]), .Z(N103) );
  OR2D0 C1747 ( .A1(g[103]), .A2(N103), .Z(c[104]) );
  AN2D0 C1746 ( .A1(p[102]), .A2(c[102]), .Z(N102) );
  OR2D0 C1745 ( .A1(g[102]), .A2(N102), .Z(c[103]) );
  AN2D0 C1744 ( .A1(p[101]), .A2(c[101]), .Z(N101) );
  OR2D0 C1743 ( .A1(g[101]), .A2(N101), .Z(c[102]) );
  AN2D0 C1742 ( .A1(p[100]), .A2(c[100]), .Z(N100) );
  OR2D0 C1741 ( .A1(g[100]), .A2(N100), .Z(c[101]) );
  AN2D0 C1740 ( .A1(p[99]), .A2(c[99]), .Z(N99) );
  OR2D0 C1739 ( .A1(g[99]), .A2(N99), .Z(c[100]) );
  AN2D0 C1738 ( .A1(p[98]), .A2(c[98]), .Z(N98) );
  OR2D0 C1737 ( .A1(g[98]), .A2(N98), .Z(c[99]) );
  AN2D0 C1736 ( .A1(p[97]), .A2(c[97]), .Z(N97) );
  OR2D0 C1735 ( .A1(g[97]), .A2(N97), .Z(c[98]) );
  AN2D0 C1734 ( .A1(p[96]), .A2(c[96]), .Z(N96) );
  OR2D0 C1733 ( .A1(g[96]), .A2(N96), .Z(c[97]) );
  AN2D0 C1732 ( .A1(p[95]), .A2(c[95]), .Z(N95) );
  OR2D0 C1731 ( .A1(g[95]), .A2(N95), .Z(c[96]) );
  AN2D0 C1730 ( .A1(p[94]), .A2(c[94]), .Z(N94) );
  OR2D0 C1729 ( .A1(g[94]), .A2(N94), .Z(c[95]) );
  AN2D0 C1728 ( .A1(p[93]), .A2(c[93]), .Z(N93) );
  OR2D0 C1727 ( .A1(g[93]), .A2(N93), .Z(c[94]) );
  AN2D0 C1726 ( .A1(p[92]), .A2(c[92]), .Z(N92) );
  OR2D0 C1725 ( .A1(g[92]), .A2(N92), .Z(c[93]) );
  AN2D0 C1724 ( .A1(p[91]), .A2(c[91]), .Z(N91) );
  OR2D0 C1723 ( .A1(g[91]), .A2(N91), .Z(c[92]) );
  AN2D0 C1722 ( .A1(p[90]), .A2(c[90]), .Z(N90) );
  OR2D0 C1721 ( .A1(g[90]), .A2(N90), .Z(c[91]) );
  AN2D0 C1720 ( .A1(p[89]), .A2(c[89]), .Z(N89) );
  OR2D0 C1719 ( .A1(g[89]), .A2(N89), .Z(c[90]) );
  AN2D0 C1718 ( .A1(p[88]), .A2(c[88]), .Z(N88) );
  OR2D0 C1717 ( .A1(g[88]), .A2(N88), .Z(c[89]) );
  AN2D0 C1716 ( .A1(p[87]), .A2(c[87]), .Z(N87) );
  OR2D0 C1715 ( .A1(g[87]), .A2(N87), .Z(c[88]) );
  AN2D0 C1714 ( .A1(p[86]), .A2(c[86]), .Z(N86) );
  OR2D0 C1713 ( .A1(g[86]), .A2(N86), .Z(c[87]) );
  AN2D0 C1712 ( .A1(p[85]), .A2(c[85]), .Z(N85) );
  OR2D0 C1711 ( .A1(g[85]), .A2(N85), .Z(c[86]) );
  AN2D0 C1710 ( .A1(p[84]), .A2(c[84]), .Z(N84) );
  OR2D0 C1709 ( .A1(g[84]), .A2(N84), .Z(c[85]) );
  AN2D0 C1708 ( .A1(p[83]), .A2(c[83]), .Z(N83) );
  OR2D0 C1707 ( .A1(g[83]), .A2(N83), .Z(c[84]) );
  AN2D0 C1706 ( .A1(p[82]), .A2(c[82]), .Z(N82) );
  OR2D0 C1705 ( .A1(g[82]), .A2(N82), .Z(c[83]) );
  AN2D0 C1704 ( .A1(p[81]), .A2(c[81]), .Z(N81) );
  OR2D0 C1703 ( .A1(g[81]), .A2(N81), .Z(c[82]) );
  AN2D0 C1702 ( .A1(p[80]), .A2(c[80]), .Z(N80) );
  OR2D0 C1701 ( .A1(g[80]), .A2(N80), .Z(c[81]) );
  AN2D0 C1700 ( .A1(p[79]), .A2(c[79]), .Z(N79) );
  OR2D0 C1699 ( .A1(g[79]), .A2(N79), .Z(c[80]) );
  AN2D0 C1698 ( .A1(p[78]), .A2(c[78]), .Z(N78) );
  OR2D0 C1697 ( .A1(g[78]), .A2(N78), .Z(c[79]) );
  AN2D0 C1696 ( .A1(p[77]), .A2(c[77]), .Z(N77) );
  OR2D0 C1695 ( .A1(g[77]), .A2(N77), .Z(c[78]) );
  AN2D0 C1694 ( .A1(p[76]), .A2(c[76]), .Z(N76) );
  OR2D0 C1693 ( .A1(g[76]), .A2(N76), .Z(c[77]) );
  AN2D0 C1692 ( .A1(p[75]), .A2(c[75]), .Z(N75) );
  OR2D0 C1691 ( .A1(g[75]), .A2(N75), .Z(c[76]) );
  AN2D0 C1690 ( .A1(p[74]), .A2(c[74]), .Z(N74) );
  OR2D0 C1689 ( .A1(g[74]), .A2(N74), .Z(c[75]) );
  AN2D0 C1688 ( .A1(p[73]), .A2(c[73]), .Z(N73) );
  OR2D0 C1687 ( .A1(g[73]), .A2(N73), .Z(c[74]) );
  AN2D0 C1686 ( .A1(p[72]), .A2(c[72]), .Z(N72) );
  OR2D0 C1685 ( .A1(g[72]), .A2(N72), .Z(c[73]) );
  AN2D0 C1684 ( .A1(p[71]), .A2(c[71]), .Z(N71) );
  OR2D0 C1683 ( .A1(g[71]), .A2(N71), .Z(c[72]) );
  AN2D0 C1682 ( .A1(p[70]), .A2(c[70]), .Z(N70) );
  OR2D0 C1681 ( .A1(g[70]), .A2(N70), .Z(c[71]) );
  AN2D0 C1680 ( .A1(p[69]), .A2(c[69]), .Z(N69) );
  OR2D0 C1679 ( .A1(g[69]), .A2(N69), .Z(c[70]) );
  AN2D0 C1678 ( .A1(p[68]), .A2(c[68]), .Z(N68) );
  OR2D0 C1677 ( .A1(g[68]), .A2(N68), .Z(c[69]) );
  AN2D0 C1676 ( .A1(p[67]), .A2(c[67]), .Z(N67) );
  OR2D0 C1675 ( .A1(g[67]), .A2(N67), .Z(c[68]) );
  AN2D0 C1674 ( .A1(p[66]), .A2(c[66]), .Z(N66) );
  OR2D0 C1673 ( .A1(g[66]), .A2(N66), .Z(c[67]) );
  AN2D0 C1672 ( .A1(p[65]), .A2(c[65]), .Z(N65) );
  OR2D0 C1671 ( .A1(g[65]), .A2(N65), .Z(c[66]) );
  AN2D0 C1670 ( .A1(p[64]), .A2(c[64]), .Z(N64) );
  OR2D0 C1669 ( .A1(g[64]), .A2(N64), .Z(c[65]) );
  AN2D0 C1668 ( .A1(p[63]), .A2(c[63]), .Z(N63) );
  OR2D0 C1667 ( .A1(g[63]), .A2(N63), .Z(c[64]) );
  AN2D0 C1666 ( .A1(p[62]), .A2(c[62]), .Z(N62) );
  OR2D0 C1665 ( .A1(g[62]), .A2(N62), .Z(c[63]) );
  AN2D0 C1664 ( .A1(p[61]), .A2(c[61]), .Z(N61) );
  OR2D0 C1663 ( .A1(g[61]), .A2(N61), .Z(c[62]) );
  AN2D0 C1662 ( .A1(p[60]), .A2(c[60]), .Z(N60) );
  OR2D0 C1661 ( .A1(g[60]), .A2(N60), .Z(c[61]) );
  AN2D0 C1660 ( .A1(p[59]), .A2(c[59]), .Z(N59) );
  OR2D0 C1659 ( .A1(g[59]), .A2(N59), .Z(c[60]) );
  AN2D0 C1658 ( .A1(p[58]), .A2(c[58]), .Z(N58) );
  OR2D0 C1657 ( .A1(g[58]), .A2(N58), .Z(c[59]) );
  AN2D0 C1656 ( .A1(p[57]), .A2(c[57]), .Z(N57) );
  OR2D0 C1655 ( .A1(g[57]), .A2(N57), .Z(c[58]) );
  AN2D0 C1654 ( .A1(p[56]), .A2(c[56]), .Z(N56) );
  OR2D0 C1653 ( .A1(g[56]), .A2(N56), .Z(c[57]) );
  AN2D0 C1652 ( .A1(p[55]), .A2(c[55]), .Z(N55) );
  OR2D0 C1651 ( .A1(g[55]), .A2(N55), .Z(c[56]) );
  AN2D0 C1650 ( .A1(p[54]), .A2(c[54]), .Z(N54) );
  OR2D0 C1649 ( .A1(g[54]), .A2(N54), .Z(c[55]) );
  AN2D0 C1648 ( .A1(p[53]), .A2(c[53]), .Z(N53) );
  OR2D0 C1647 ( .A1(g[53]), .A2(N53), .Z(c[54]) );
  AN2D0 C1646 ( .A1(p[52]), .A2(c[52]), .Z(N52) );
  OR2D0 C1645 ( .A1(g[52]), .A2(N52), .Z(c[53]) );
  AN2D0 C1644 ( .A1(p[51]), .A2(c[51]), .Z(N51) );
  OR2D0 C1643 ( .A1(g[51]), .A2(N51), .Z(c[52]) );
  AN2D0 C1642 ( .A1(p[50]), .A2(c[50]), .Z(N50) );
  OR2D0 C1641 ( .A1(g[50]), .A2(N50), .Z(c[51]) );
  AN2D0 C1640 ( .A1(p[49]), .A2(c[49]), .Z(N49) );
  OR2D0 C1639 ( .A1(g[49]), .A2(N49), .Z(c[50]) );
  AN2D0 C1638 ( .A1(p[48]), .A2(c[48]), .Z(N48) );
  OR2D0 C1637 ( .A1(g[48]), .A2(N48), .Z(c[49]) );
  AN2D0 C1636 ( .A1(p[47]), .A2(c[47]), .Z(N47) );
  OR2D0 C1635 ( .A1(g[47]), .A2(N47), .Z(c[48]) );
  AN2D0 C1634 ( .A1(p[46]), .A2(c[46]), .Z(N46) );
  OR2D0 C1633 ( .A1(g[46]), .A2(N46), .Z(c[47]) );
  AN2D0 C1632 ( .A1(p[45]), .A2(c[45]), .Z(N45) );
  OR2D0 C1631 ( .A1(g[45]), .A2(N45), .Z(c[46]) );
  AN2D0 C1630 ( .A1(p[44]), .A2(c[44]), .Z(N44) );
  OR2D0 C1629 ( .A1(g[44]), .A2(N44), .Z(c[45]) );
  AN2D0 C1628 ( .A1(p[43]), .A2(c[43]), .Z(N43) );
  OR2D0 C1627 ( .A1(g[43]), .A2(N43), .Z(c[44]) );
  AN2D0 C1626 ( .A1(p[42]), .A2(c[42]), .Z(N42) );
  OR2D0 C1625 ( .A1(g[42]), .A2(N42), .Z(c[43]) );
  AN2D0 C1624 ( .A1(p[41]), .A2(c[41]), .Z(N41) );
  OR2D0 C1623 ( .A1(g[41]), .A2(N41), .Z(c[42]) );
  AN2D0 C1622 ( .A1(p[40]), .A2(c[40]), .Z(N40) );
  OR2D0 C1621 ( .A1(g[40]), .A2(N40), .Z(c[41]) );
  AN2D0 C1620 ( .A1(p[39]), .A2(c[39]), .Z(N39) );
  OR2D0 C1619 ( .A1(g[39]), .A2(N39), .Z(c[40]) );
  AN2D0 C1618 ( .A1(p[38]), .A2(c[38]), .Z(N38) );
  OR2D0 C1617 ( .A1(g[38]), .A2(N38), .Z(c[39]) );
  AN2D0 C1616 ( .A1(p[37]), .A2(c[37]), .Z(N37) );
  OR2D0 C1615 ( .A1(g[37]), .A2(N37), .Z(c[38]) );
  AN2D0 C1614 ( .A1(p[36]), .A2(c[36]), .Z(N36) );
  OR2D0 C1613 ( .A1(g[36]), .A2(N36), .Z(c[37]) );
  AN2D0 C1612 ( .A1(p[35]), .A2(c[35]), .Z(N35) );
  OR2D0 C1611 ( .A1(g[35]), .A2(N35), .Z(c[36]) );
  AN2D0 C1610 ( .A1(p[34]), .A2(c[34]), .Z(N34) );
  OR2D0 C1609 ( .A1(g[34]), .A2(N34), .Z(c[35]) );
  AN2D0 C1608 ( .A1(p[33]), .A2(c[33]), .Z(N33) );
  OR2D0 C1607 ( .A1(g[33]), .A2(N33), .Z(c[34]) );
  AN2D0 C1606 ( .A1(p[32]), .A2(c[32]), .Z(N32) );
  OR2D0 C1605 ( .A1(g[32]), .A2(N32), .Z(c[33]) );
  AN2D0 C1604 ( .A1(p[31]), .A2(c[31]), .Z(N31) );
  OR2D0 C1603 ( .A1(g[31]), .A2(N31), .Z(c[32]) );
  AN2D0 C1602 ( .A1(p[30]), .A2(c[30]), .Z(N30) );
  OR2D0 C1601 ( .A1(g[30]), .A2(N30), .Z(c[31]) );
  AN2D0 C1600 ( .A1(p[29]), .A2(c[29]), .Z(N29) );
  OR2D0 C1599 ( .A1(g[29]), .A2(N29), .Z(c[30]) );
  AN2D0 C1598 ( .A1(p[28]), .A2(c[28]), .Z(N28) );
  OR2D0 C1597 ( .A1(g[28]), .A2(N28), .Z(c[29]) );
  AN2D0 C1596 ( .A1(p[27]), .A2(c[27]), .Z(N27) );
  OR2D0 C1595 ( .A1(g[27]), .A2(N27), .Z(c[28]) );
  AN2D0 C1594 ( .A1(p[26]), .A2(c[26]), .Z(N26) );
  OR2D0 C1593 ( .A1(g[26]), .A2(N26), .Z(c[27]) );
  AN2D0 C1592 ( .A1(p[25]), .A2(c[25]), .Z(N25) );
  OR2D0 C1591 ( .A1(g[25]), .A2(N25), .Z(c[26]) );
  AN2D0 C1590 ( .A1(p[24]), .A2(c[24]), .Z(N24) );
  OR2D0 C1589 ( .A1(g[24]), .A2(N24), .Z(c[25]) );
  AN2D0 C1588 ( .A1(p[23]), .A2(c[23]), .Z(N23) );
  OR2D0 C1587 ( .A1(g[23]), .A2(N23), .Z(c[24]) );
  AN2D0 C1586 ( .A1(p[22]), .A2(c[22]), .Z(N22) );
  OR2D0 C1585 ( .A1(g[22]), .A2(N22), .Z(c[23]) );
  AN2D0 C1584 ( .A1(p[21]), .A2(c[21]), .Z(N21) );
  OR2D0 C1583 ( .A1(g[21]), .A2(N21), .Z(c[22]) );
  AN2D0 C1582 ( .A1(p[20]), .A2(c[20]), .Z(N20) );
  OR2D0 C1581 ( .A1(g[20]), .A2(N20), .Z(c[21]) );
  AN2D0 C1580 ( .A1(p[19]), .A2(c[19]), .Z(N19) );
  OR2D0 C1579 ( .A1(g[19]), .A2(N19), .Z(c[20]) );
  AN2D0 C1578 ( .A1(p[18]), .A2(c[18]), .Z(N18) );
  OR2D0 C1577 ( .A1(g[18]), .A2(N18), .Z(c[19]) );
  AN2D0 C1576 ( .A1(p[17]), .A2(c[17]), .Z(N17) );
  OR2D0 C1575 ( .A1(g[17]), .A2(N17), .Z(c[18]) );
  AN2D0 C1574 ( .A1(p[16]), .A2(c[16]), .Z(N16) );
  OR2D0 C1573 ( .A1(g[16]), .A2(N16), .Z(c[17]) );
  AN2D0 C1572 ( .A1(p[15]), .A2(c[15]), .Z(N15) );
  OR2D0 C1571 ( .A1(g[15]), .A2(N15), .Z(c[16]) );
  AN2D0 C1570 ( .A1(p[14]), .A2(c[14]), .Z(N14) );
  OR2D0 C1569 ( .A1(g[14]), .A2(N14), .Z(c[15]) );
  AN2D0 C1568 ( .A1(p[13]), .A2(c[13]), .Z(N13) );
  OR2D0 C1567 ( .A1(g[13]), .A2(N13), .Z(c[14]) );
  AN2D0 C1566 ( .A1(p[12]), .A2(c[12]), .Z(N12) );
  OR2D0 C1565 ( .A1(g[12]), .A2(N12), .Z(c[13]) );
  AN2D0 C1564 ( .A1(p[11]), .A2(c[11]), .Z(N11) );
  OR2D0 C1563 ( .A1(g[11]), .A2(N11), .Z(c[12]) );
  AN2D0 C1562 ( .A1(p[10]), .A2(c[10]), .Z(N10) );
  OR2D0 C1561 ( .A1(g[10]), .A2(N10), .Z(c[11]) );
  AN2D0 C1560 ( .A1(p[9]), .A2(c[9]), .Z(N9) );
  OR2D0 C1559 ( .A1(g[9]), .A2(N9), .Z(c[10]) );
  AN2D0 C1558 ( .A1(p[8]), .A2(c[8]), .Z(N8) );
  OR2D0 C1557 ( .A1(g[8]), .A2(N8), .Z(c[9]) );
  AN2D0 C1556 ( .A1(p[7]), .A2(c[7]), .Z(N7) );
  OR2D0 C1555 ( .A1(g[7]), .A2(N7), .Z(c[8]) );
  AN2D0 C1554 ( .A1(p[6]), .A2(c[6]), .Z(N6) );
  OR2D0 C1553 ( .A1(g[6]), .A2(N6), .Z(c[7]) );
  AN2D0 C1552 ( .A1(p[5]), .A2(c[5]), .Z(N5) );
  OR2D0 C1551 ( .A1(g[5]), .A2(N5), .Z(c[6]) );
  AN2D0 C1550 ( .A1(p[4]), .A2(c[4]), .Z(N4) );
  OR2D0 C1549 ( .A1(g[4]), .A2(N4), .Z(c[5]) );
  AN2D0 C1548 ( .A1(p[3]), .A2(c[3]), .Z(N3) );
  OR2D0 C1547 ( .A1(g[3]), .A2(N3), .Z(c[4]) );
  AN2D0 C1546 ( .A1(p[2]), .A2(c[2]), .Z(N2) );
  OR2D0 C1545 ( .A1(g[2]), .A2(N2), .Z(c[3]) );
  AN2D0 C1544 ( .A1(p[1]), .A2(c[1]), .Z(N1) );
  OR2D0 C1543 ( .A1(g[1]), .A2(N1), .Z(c[2]) );
  AN2D0 C1542 ( .A1(p[0]), .A2(cin), .Z(N0) );
  OR2D0 C1541 ( .A1(g[0]), .A2(N0), .Z(c[1]) );
  XOR2D0 C1540 ( .A1(a[0]), .A2(b[0]), .Z(p[0]) );
  XOR2D0 C1539 ( .A1(a[1]), .A2(b[1]), .Z(p[1]) );
  XOR2D0 C1538 ( .A1(a[2]), .A2(b[2]), .Z(p[2]) );
  XOR2D0 C1537 ( .A1(a[3]), .A2(b[3]), .Z(p[3]) );
  XOR2D0 C1536 ( .A1(a[4]), .A2(b[4]), .Z(p[4]) );
  XOR2D0 C1535 ( .A1(a[5]), .A2(b[5]), .Z(p[5]) );
  XOR2D0 C1534 ( .A1(a[6]), .A2(b[6]), .Z(p[6]) );
  XOR2D0 C1533 ( .A1(a[7]), .A2(b[7]), .Z(p[7]) );
  XOR2D0 C1532 ( .A1(a[8]), .A2(b[8]), .Z(p[8]) );
  XOR2D0 C1531 ( .A1(a[9]), .A2(b[9]), .Z(p[9]) );
  XOR2D0 C1530 ( .A1(a[10]), .A2(b[10]), .Z(p[10]) );
  XOR2D0 C1529 ( .A1(a[11]), .A2(b[11]), .Z(p[11]) );
  XOR2D0 C1528 ( .A1(a[12]), .A2(b[12]), .Z(p[12]) );
  XOR2D0 C1527 ( .A1(a[13]), .A2(b[13]), .Z(p[13]) );
  XOR2D0 C1526 ( .A1(a[14]), .A2(b[14]), .Z(p[14]) );
  XOR2D0 C1525 ( .A1(a[15]), .A2(b[15]), .Z(p[15]) );
  XOR2D0 C1524 ( .A1(a[16]), .A2(b[16]), .Z(p[16]) );
  XOR2D0 C1523 ( .A1(a[17]), .A2(b[17]), .Z(p[17]) );
  XOR2D0 C1522 ( .A1(a[18]), .A2(b[18]), .Z(p[18]) );
  XOR2D0 C1521 ( .A1(a[19]), .A2(b[19]), .Z(p[19]) );
  XOR2D0 C1520 ( .A1(a[20]), .A2(b[20]), .Z(p[20]) );
  XOR2D0 C1519 ( .A1(a[21]), .A2(b[21]), .Z(p[21]) );
  XOR2D0 C1518 ( .A1(a[22]), .A2(b[22]), .Z(p[22]) );
  XOR2D0 C1517 ( .A1(a[23]), .A2(b[23]), .Z(p[23]) );
  XOR2D0 C1516 ( .A1(a[24]), .A2(b[24]), .Z(p[24]) );
  XOR2D0 C1515 ( .A1(a[25]), .A2(b[25]), .Z(p[25]) );
  XOR2D0 C1514 ( .A1(a[26]), .A2(b[26]), .Z(p[26]) );
  XOR2D0 C1513 ( .A1(a[27]), .A2(b[27]), .Z(p[27]) );
  XOR2D0 C1512 ( .A1(a[28]), .A2(b[28]), .Z(p[28]) );
  XOR2D0 C1511 ( .A1(a[29]), .A2(b[29]), .Z(p[29]) );
  XOR2D0 C1510 ( .A1(a[30]), .A2(b[30]), .Z(p[30]) );
  XOR2D0 C1509 ( .A1(a[31]), .A2(b[31]), .Z(p[31]) );
  XOR2D0 C1508 ( .A1(a[32]), .A2(b[32]), .Z(p[32]) );
  XOR2D0 C1507 ( .A1(a[33]), .A2(b[33]), .Z(p[33]) );
  XOR2D0 C1506 ( .A1(a[34]), .A2(b[34]), .Z(p[34]) );
  XOR2D0 C1505 ( .A1(a[35]), .A2(b[35]), .Z(p[35]) );
  XOR2D0 C1504 ( .A1(a[36]), .A2(b[36]), .Z(p[36]) );
  XOR2D0 C1503 ( .A1(a[37]), .A2(b[37]), .Z(p[37]) );
  XOR2D0 C1502 ( .A1(a[38]), .A2(b[38]), .Z(p[38]) );
  XOR2D0 C1501 ( .A1(a[39]), .A2(b[39]), .Z(p[39]) );
  XOR2D0 C1500 ( .A1(a[40]), .A2(b[40]), .Z(p[40]) );
  XOR2D0 C1499 ( .A1(a[41]), .A2(b[41]), .Z(p[41]) );
  XOR2D0 C1498 ( .A1(a[42]), .A2(b[42]), .Z(p[42]) );
  XOR2D0 C1497 ( .A1(a[43]), .A2(b[43]), .Z(p[43]) );
  XOR2D0 C1496 ( .A1(a[44]), .A2(b[44]), .Z(p[44]) );
  XOR2D0 C1495 ( .A1(a[45]), .A2(b[45]), .Z(p[45]) );
  XOR2D0 C1494 ( .A1(a[46]), .A2(b[46]), .Z(p[46]) );
  XOR2D0 C1493 ( .A1(a[47]), .A2(b[47]), .Z(p[47]) );
  XOR2D0 C1492 ( .A1(a[48]), .A2(b[48]), .Z(p[48]) );
  XOR2D0 C1491 ( .A1(a[49]), .A2(b[49]), .Z(p[49]) );
  XOR2D0 C1490 ( .A1(a[50]), .A2(b[50]), .Z(p[50]) );
  XOR2D0 C1489 ( .A1(a[51]), .A2(b[51]), .Z(p[51]) );
  XOR2D0 C1488 ( .A1(a[52]), .A2(b[52]), .Z(p[52]) );
  XOR2D0 C1487 ( .A1(a[53]), .A2(b[53]), .Z(p[53]) );
  XOR2D0 C1486 ( .A1(a[54]), .A2(b[54]), .Z(p[54]) );
  XOR2D0 C1485 ( .A1(a[55]), .A2(b[55]), .Z(p[55]) );
  XOR2D0 C1484 ( .A1(a[56]), .A2(b[56]), .Z(p[56]) );
  XOR2D0 C1483 ( .A1(a[57]), .A2(b[57]), .Z(p[57]) );
  XOR2D0 C1482 ( .A1(a[58]), .A2(b[58]), .Z(p[58]) );
  XOR2D0 C1481 ( .A1(a[59]), .A2(b[59]), .Z(p[59]) );
  XOR2D0 C1480 ( .A1(a[60]), .A2(b[60]), .Z(p[60]) );
  XOR2D0 C1479 ( .A1(a[61]), .A2(b[61]), .Z(p[61]) );
  XOR2D0 C1478 ( .A1(a[62]), .A2(b[62]), .Z(p[62]) );
  XOR2D0 C1477 ( .A1(a[63]), .A2(b[63]), .Z(p[63]) );
  XOR2D0 C1476 ( .A1(a[64]), .A2(b[64]), .Z(p[64]) );
  XOR2D0 C1475 ( .A1(a[65]), .A2(b[65]), .Z(p[65]) );
  XOR2D0 C1474 ( .A1(a[66]), .A2(b[66]), .Z(p[66]) );
  XOR2D0 C1473 ( .A1(a[67]), .A2(b[67]), .Z(p[67]) );
  XOR2D0 C1472 ( .A1(a[68]), .A2(b[68]), .Z(p[68]) );
  XOR2D0 C1471 ( .A1(a[69]), .A2(b[69]), .Z(p[69]) );
  XOR2D0 C1470 ( .A1(a[70]), .A2(b[70]), .Z(p[70]) );
  XOR2D0 C1469 ( .A1(a[71]), .A2(b[71]), .Z(p[71]) );
  XOR2D0 C1468 ( .A1(a[72]), .A2(b[72]), .Z(p[72]) );
  XOR2D0 C1467 ( .A1(a[73]), .A2(b[73]), .Z(p[73]) );
  XOR2D0 C1466 ( .A1(a[74]), .A2(b[74]), .Z(p[74]) );
  XOR2D0 C1465 ( .A1(a[75]), .A2(b[75]), .Z(p[75]) );
  XOR2D0 C1464 ( .A1(a[76]), .A2(b[76]), .Z(p[76]) );
  XOR2D0 C1463 ( .A1(a[77]), .A2(b[77]), .Z(p[77]) );
  XOR2D0 C1462 ( .A1(a[78]), .A2(b[78]), .Z(p[78]) );
  XOR2D0 C1461 ( .A1(a[79]), .A2(b[79]), .Z(p[79]) );
  XOR2D0 C1460 ( .A1(a[80]), .A2(b[80]), .Z(p[80]) );
  XOR2D0 C1459 ( .A1(a[81]), .A2(b[81]), .Z(p[81]) );
  XOR2D0 C1458 ( .A1(a[82]), .A2(b[82]), .Z(p[82]) );
  XOR2D0 C1457 ( .A1(a[83]), .A2(b[83]), .Z(p[83]) );
  XOR2D0 C1456 ( .A1(a[84]), .A2(b[84]), .Z(p[84]) );
  XOR2D0 C1455 ( .A1(a[85]), .A2(b[85]), .Z(p[85]) );
  XOR2D0 C1454 ( .A1(a[86]), .A2(b[86]), .Z(p[86]) );
  XOR2D0 C1453 ( .A1(a[87]), .A2(b[87]), .Z(p[87]) );
  XOR2D0 C1452 ( .A1(a[88]), .A2(b[88]), .Z(p[88]) );
  XOR2D0 C1451 ( .A1(a[89]), .A2(b[89]), .Z(p[89]) );
  XOR2D0 C1450 ( .A1(a[90]), .A2(b[90]), .Z(p[90]) );
  XOR2D0 C1449 ( .A1(a[91]), .A2(b[91]), .Z(p[91]) );
  XOR2D0 C1448 ( .A1(a[92]), .A2(b[92]), .Z(p[92]) );
  XOR2D0 C1447 ( .A1(a[93]), .A2(b[93]), .Z(p[93]) );
  XOR2D0 C1446 ( .A1(a[94]), .A2(b[94]), .Z(p[94]) );
  XOR2D0 C1445 ( .A1(a[95]), .A2(b[95]), .Z(p[95]) );
  XOR2D0 C1444 ( .A1(a[96]), .A2(b[96]), .Z(p[96]) );
  XOR2D0 C1443 ( .A1(a[97]), .A2(b[97]), .Z(p[97]) );
  XOR2D0 C1442 ( .A1(a[98]), .A2(b[98]), .Z(p[98]) );
  XOR2D0 C1441 ( .A1(a[99]), .A2(b[99]), .Z(p[99]) );
  XOR2D0 C1440 ( .A1(a[100]), .A2(b[100]), .Z(p[100]) );
  XOR2D0 C1439 ( .A1(a[101]), .A2(b[101]), .Z(p[101]) );
  XOR2D0 C1438 ( .A1(a[102]), .A2(b[102]), .Z(p[102]) );
  XOR2D0 C1437 ( .A1(a[103]), .A2(b[103]), .Z(p[103]) );
  XOR2D0 C1436 ( .A1(a[104]), .A2(b[104]), .Z(p[104]) );
  XOR2D0 C1435 ( .A1(a[105]), .A2(b[105]), .Z(p[105]) );
  XOR2D0 C1434 ( .A1(a[106]), .A2(b[106]), .Z(p[106]) );
  XOR2D0 C1433 ( .A1(a[107]), .A2(b[107]), .Z(p[107]) );
  XOR2D0 C1432 ( .A1(a[108]), .A2(b[108]), .Z(p[108]) );
  XOR2D0 C1431 ( .A1(a[109]), .A2(b[109]), .Z(p[109]) );
  XOR2D0 C1430 ( .A1(a[110]), .A2(b[110]), .Z(p[110]) );
  XOR2D0 C1429 ( .A1(a[111]), .A2(b[111]), .Z(p[111]) );
  XOR2D0 C1428 ( .A1(a[112]), .A2(b[112]), .Z(p[112]) );
  XOR2D0 C1427 ( .A1(a[113]), .A2(b[113]), .Z(p[113]) );
  XOR2D0 C1426 ( .A1(a[114]), .A2(b[114]), .Z(p[114]) );
  XOR2D0 C1425 ( .A1(a[115]), .A2(b[115]), .Z(p[115]) );
  XOR2D0 C1424 ( .A1(a[116]), .A2(b[116]), .Z(p[116]) );
  XOR2D0 C1423 ( .A1(a[117]), .A2(b[117]), .Z(p[117]) );
  XOR2D0 C1422 ( .A1(a[118]), .A2(b[118]), .Z(p[118]) );
  XOR2D0 C1421 ( .A1(a[119]), .A2(b[119]), .Z(p[119]) );
  XOR2D0 C1420 ( .A1(a[120]), .A2(b[120]), .Z(p[120]) );
  XOR2D0 C1419 ( .A1(a[121]), .A2(b[121]), .Z(p[121]) );
  XOR2D0 C1418 ( .A1(a[122]), .A2(b[122]), .Z(p[122]) );
  XOR2D0 C1417 ( .A1(a[123]), .A2(b[123]), .Z(p[123]) );
  XOR2D0 C1416 ( .A1(a[124]), .A2(b[124]), .Z(p[124]) );
  XOR2D0 C1415 ( .A1(a[125]), .A2(b[125]), .Z(p[125]) );
  XOR2D0 C1414 ( .A1(a[126]), .A2(b[126]), .Z(p[126]) );
  XOR2D0 C1413 ( .A1(a[127]), .A2(b[127]), .Z(p[127]) );
  XOR2D0 C1412 ( .A1(a[128]), .A2(b[128]), .Z(p[128]) );
  XOR2D0 C1411 ( .A1(a[129]), .A2(b[129]), .Z(p[129]) );
  XOR2D0 C1410 ( .A1(a[130]), .A2(b[130]), .Z(p[130]) );
  XOR2D0 C1409 ( .A1(a[131]), .A2(b[131]), .Z(p[131]) );
  XOR2D0 C1408 ( .A1(a[132]), .A2(b[132]), .Z(p[132]) );
  XOR2D0 C1407 ( .A1(a[133]), .A2(b[133]), .Z(p[133]) );
  XOR2D0 C1406 ( .A1(a[134]), .A2(b[134]), .Z(p[134]) );
  XOR2D0 C1405 ( .A1(a[135]), .A2(b[135]), .Z(p[135]) );
  XOR2D0 C1404 ( .A1(a[136]), .A2(b[136]), .Z(p[136]) );
  XOR2D0 C1403 ( .A1(a[137]), .A2(b[137]), .Z(p[137]) );
  XOR2D0 C1402 ( .A1(a[138]), .A2(b[138]), .Z(p[138]) );
  XOR2D0 C1401 ( .A1(a[139]), .A2(b[139]), .Z(p[139]) );
  XOR2D0 C1400 ( .A1(a[140]), .A2(b[140]), .Z(p[140]) );
  XOR2D0 C1399 ( .A1(a[141]), .A2(b[141]), .Z(p[141]) );
  XOR2D0 C1398 ( .A1(a[142]), .A2(b[142]), .Z(p[142]) );
  XOR2D0 C1397 ( .A1(a[143]), .A2(b[143]), .Z(p[143]) );
  XOR2D0 C1396 ( .A1(a[144]), .A2(b[144]), .Z(p[144]) );
  XOR2D0 C1395 ( .A1(a[145]), .A2(b[145]), .Z(p[145]) );
  XOR2D0 C1394 ( .A1(a[146]), .A2(b[146]), .Z(p[146]) );
  XOR2D0 C1393 ( .A1(a[147]), .A2(b[147]), .Z(p[147]) );
  XOR2D0 C1392 ( .A1(a[148]), .A2(b[148]), .Z(p[148]) );
  XOR2D0 C1391 ( .A1(a[149]), .A2(b[149]), .Z(p[149]) );
  XOR2D0 C1390 ( .A1(a[150]), .A2(b[150]), .Z(p[150]) );
  XOR2D0 C1389 ( .A1(a[151]), .A2(b[151]), .Z(p[151]) );
  XOR2D0 C1388 ( .A1(a[152]), .A2(b[152]), .Z(p[152]) );
  XOR2D0 C1387 ( .A1(a[153]), .A2(b[153]), .Z(p[153]) );
  XOR2D0 C1386 ( .A1(a[154]), .A2(b[154]), .Z(p[154]) );
  XOR2D0 C1385 ( .A1(a[155]), .A2(b[155]), .Z(p[155]) );
  XOR2D0 C1384 ( .A1(a[156]), .A2(b[156]), .Z(p[156]) );
  XOR2D0 C1383 ( .A1(a[157]), .A2(b[157]), .Z(p[157]) );
  XOR2D0 C1382 ( .A1(a[158]), .A2(b[158]), .Z(p[158]) );
  XOR2D0 C1381 ( .A1(a[159]), .A2(b[159]), .Z(p[159]) );
  XOR2D0 C1380 ( .A1(a[160]), .A2(b[160]), .Z(p[160]) );
  XOR2D0 C1379 ( .A1(a[161]), .A2(b[161]), .Z(p[161]) );
  XOR2D0 C1378 ( .A1(a[162]), .A2(b[162]), .Z(p[162]) );
  XOR2D0 C1377 ( .A1(a[163]), .A2(b[163]), .Z(p[163]) );
  XOR2D0 C1376 ( .A1(a[164]), .A2(b[164]), .Z(p[164]) );
  XOR2D0 C1375 ( .A1(a[165]), .A2(b[165]), .Z(p[165]) );
  XOR2D0 C1374 ( .A1(a[166]), .A2(b[166]), .Z(p[166]) );
  XOR2D0 C1373 ( .A1(a[167]), .A2(b[167]), .Z(p[167]) );
  XOR2D0 C1372 ( .A1(a[168]), .A2(b[168]), .Z(p[168]) );
  XOR2D0 C1371 ( .A1(a[169]), .A2(b[169]), .Z(p[169]) );
  XOR2D0 C1370 ( .A1(a[170]), .A2(b[170]), .Z(p[170]) );
  XOR2D0 C1369 ( .A1(a[171]), .A2(b[171]), .Z(p[171]) );
  XOR2D0 C1368 ( .A1(a[172]), .A2(b[172]), .Z(p[172]) );
  XOR2D0 C1367 ( .A1(a[173]), .A2(b[173]), .Z(p[173]) );
  XOR2D0 C1366 ( .A1(a[174]), .A2(b[174]), .Z(p[174]) );
  XOR2D0 C1365 ( .A1(a[175]), .A2(b[175]), .Z(p[175]) );
  XOR2D0 C1364 ( .A1(a[176]), .A2(b[176]), .Z(p[176]) );
  XOR2D0 C1363 ( .A1(a[177]), .A2(b[177]), .Z(p[177]) );
  XOR2D0 C1362 ( .A1(a[178]), .A2(b[178]), .Z(p[178]) );
  XOR2D0 C1361 ( .A1(a[179]), .A2(b[179]), .Z(p[179]) );
  XOR2D0 C1360 ( .A1(a[180]), .A2(b[180]), .Z(p[180]) );
  XOR2D0 C1359 ( .A1(a[181]), .A2(b[181]), .Z(p[181]) );
  XOR2D0 C1358 ( .A1(a[182]), .A2(b[182]), .Z(p[182]) );
  XOR2D0 C1357 ( .A1(a[183]), .A2(b[183]), .Z(p[183]) );
  XOR2D0 C1356 ( .A1(a[184]), .A2(b[184]), .Z(p[184]) );
  XOR2D0 C1355 ( .A1(a[185]), .A2(b[185]), .Z(p[185]) );
  XOR2D0 C1354 ( .A1(a[186]), .A2(b[186]), .Z(p[186]) );
  XOR2D0 C1353 ( .A1(a[187]), .A2(b[187]), .Z(p[187]) );
  XOR2D0 C1352 ( .A1(a[188]), .A2(b[188]), .Z(p[188]) );
  XOR2D0 C1351 ( .A1(a[189]), .A2(b[189]), .Z(p[189]) );
  XOR2D0 C1350 ( .A1(a[190]), .A2(b[190]), .Z(p[190]) );
  XOR2D0 C1349 ( .A1(a[191]), .A2(b[191]), .Z(p[191]) );
  XOR2D0 C1348 ( .A1(a[192]), .A2(b[192]), .Z(p[192]) );
  XOR2D0 C1347 ( .A1(a[193]), .A2(b[193]), .Z(p[193]) );
  XOR2D0 C1346 ( .A1(a[194]), .A2(b[194]), .Z(p[194]) );
  XOR2D0 C1345 ( .A1(a[195]), .A2(b[195]), .Z(p[195]) );
  XOR2D0 C1344 ( .A1(a[196]), .A2(b[196]), .Z(p[196]) );
  XOR2D0 C1343 ( .A1(a[197]), .A2(b[197]), .Z(p[197]) );
  XOR2D0 C1342 ( .A1(a[198]), .A2(b[198]), .Z(p[198]) );
  XOR2D0 C1341 ( .A1(a[199]), .A2(b[199]), .Z(p[199]) );
  XOR2D0 C1340 ( .A1(a[200]), .A2(b[200]), .Z(p[200]) );
  XOR2D0 C1339 ( .A1(a[201]), .A2(b[201]), .Z(p[201]) );
  XOR2D0 C1338 ( .A1(a[202]), .A2(b[202]), .Z(p[202]) );
  XOR2D0 C1337 ( .A1(a[203]), .A2(b[203]), .Z(p[203]) );
  XOR2D0 C1336 ( .A1(a[204]), .A2(b[204]), .Z(p[204]) );
  XOR2D0 C1335 ( .A1(a[205]), .A2(b[205]), .Z(p[205]) );
  XOR2D0 C1334 ( .A1(a[206]), .A2(b[206]), .Z(p[206]) );
  XOR2D0 C1333 ( .A1(a[207]), .A2(b[207]), .Z(p[207]) );
  XOR2D0 C1332 ( .A1(a[208]), .A2(b[208]), .Z(p[208]) );
  XOR2D0 C1331 ( .A1(a[209]), .A2(b[209]), .Z(p[209]) );
  XOR2D0 C1330 ( .A1(a[210]), .A2(b[210]), .Z(p[210]) );
  XOR2D0 C1329 ( .A1(a[211]), .A2(b[211]), .Z(p[211]) );
  XOR2D0 C1328 ( .A1(a[212]), .A2(b[212]), .Z(p[212]) );
  XOR2D0 C1327 ( .A1(a[213]), .A2(b[213]), .Z(p[213]) );
  XOR2D0 C1326 ( .A1(a[214]), .A2(b[214]), .Z(p[214]) );
  XOR2D0 C1325 ( .A1(a[215]), .A2(b[215]), .Z(p[215]) );
  XOR2D0 C1324 ( .A1(a[216]), .A2(b[216]), .Z(p[216]) );
  XOR2D0 C1323 ( .A1(a[217]), .A2(b[217]), .Z(p[217]) );
  XOR2D0 C1322 ( .A1(a[218]), .A2(b[218]), .Z(p[218]) );
  XOR2D0 C1321 ( .A1(a[219]), .A2(b[219]), .Z(p[219]) );
  XOR2D0 C1320 ( .A1(a[220]), .A2(b[220]), .Z(p[220]) );
  XOR2D0 C1319 ( .A1(a[221]), .A2(b[221]), .Z(p[221]) );
  XOR2D0 C1318 ( .A1(a[222]), .A2(b[222]), .Z(p[222]) );
  XOR2D0 C1317 ( .A1(a[223]), .A2(b[223]), .Z(p[223]) );
  XOR2D0 C1316 ( .A1(a[224]), .A2(b[224]), .Z(p[224]) );
  XOR2D0 C1315 ( .A1(a[225]), .A2(b[225]), .Z(p[225]) );
  XOR2D0 C1314 ( .A1(a[226]), .A2(b[226]), .Z(p[226]) );
  XOR2D0 C1313 ( .A1(a[227]), .A2(b[227]), .Z(p[227]) );
  XOR2D0 C1312 ( .A1(a[228]), .A2(b[228]), .Z(p[228]) );
  XOR2D0 C1311 ( .A1(a[229]), .A2(b[229]), .Z(p[229]) );
  XOR2D0 C1310 ( .A1(a[230]), .A2(b[230]), .Z(p[230]) );
  XOR2D0 C1309 ( .A1(a[231]), .A2(b[231]), .Z(p[231]) );
  XOR2D0 C1308 ( .A1(a[232]), .A2(b[232]), .Z(p[232]) );
  XOR2D0 C1307 ( .A1(a[233]), .A2(b[233]), .Z(p[233]) );
  XOR2D0 C1306 ( .A1(a[234]), .A2(b[234]), .Z(p[234]) );
  XOR2D0 C1305 ( .A1(a[235]), .A2(b[235]), .Z(p[235]) );
  XOR2D0 C1304 ( .A1(a[236]), .A2(b[236]), .Z(p[236]) );
  XOR2D0 C1303 ( .A1(a[237]), .A2(b[237]), .Z(p[237]) );
  XOR2D0 C1302 ( .A1(a[238]), .A2(b[238]), .Z(p[238]) );
  XOR2D0 C1301 ( .A1(a[239]), .A2(b[239]), .Z(p[239]) );
  XOR2D0 C1300 ( .A1(a[240]), .A2(b[240]), .Z(p[240]) );
  XOR2D0 C1299 ( .A1(a[241]), .A2(b[241]), .Z(p[241]) );
  XOR2D0 C1298 ( .A1(a[242]), .A2(b[242]), .Z(p[242]) );
  XOR2D0 C1297 ( .A1(a[243]), .A2(b[243]), .Z(p[243]) );
  XOR2D0 C1296 ( .A1(a[244]), .A2(b[244]), .Z(p[244]) );
  XOR2D0 C1295 ( .A1(a[245]), .A2(b[245]), .Z(p[245]) );
  XOR2D0 C1294 ( .A1(a[246]), .A2(b[246]), .Z(p[246]) );
  XOR2D0 C1293 ( .A1(a[247]), .A2(b[247]), .Z(p[247]) );
  XOR2D0 C1292 ( .A1(a[248]), .A2(b[248]), .Z(p[248]) );
  XOR2D0 C1291 ( .A1(a[249]), .A2(b[249]), .Z(p[249]) );
  XOR2D0 C1290 ( .A1(a[250]), .A2(b[250]), .Z(p[250]) );
  XOR2D0 C1289 ( .A1(a[251]), .A2(b[251]), .Z(p[251]) );
  XOR2D0 C1288 ( .A1(a[252]), .A2(b[252]), .Z(p[252]) );
  XOR2D0 C1287 ( .A1(a[253]), .A2(b[253]), .Z(p[253]) );
  XOR2D0 C1286 ( .A1(a[254]), .A2(b[254]), .Z(p[254]) );
  XOR2D0 C1285 ( .A1(a[255]), .A2(b[255]), .Z(p[255]) );
  AN2D0 C1284 ( .A1(a[0]), .A2(b[0]), .Z(g[0]) );
  AN2D0 C1283 ( .A1(a[1]), .A2(b[1]), .Z(g[1]) );
  AN2D0 C1282 ( .A1(a[2]), .A2(b[2]), .Z(g[2]) );
  AN2D0 C1281 ( .A1(a[3]), .A2(b[3]), .Z(g[3]) );
  AN2D0 C1280 ( .A1(a[4]), .A2(b[4]), .Z(g[4]) );
  AN2D0 C1279 ( .A1(a[5]), .A2(b[5]), .Z(g[5]) );
  AN2D0 C1278 ( .A1(a[6]), .A2(b[6]), .Z(g[6]) );
  AN2D0 C1277 ( .A1(a[7]), .A2(b[7]), .Z(g[7]) );
  AN2D0 C1276 ( .A1(a[8]), .A2(b[8]), .Z(g[8]) );
  AN2D0 C1275 ( .A1(a[9]), .A2(b[9]), .Z(g[9]) );
  AN2D0 C1274 ( .A1(a[10]), .A2(b[10]), .Z(g[10]) );
  AN2D0 C1273 ( .A1(a[11]), .A2(b[11]), .Z(g[11]) );
  AN2D0 C1272 ( .A1(a[12]), .A2(b[12]), .Z(g[12]) );
  AN2D0 C1271 ( .A1(a[13]), .A2(b[13]), .Z(g[13]) );
  AN2D0 C1270 ( .A1(a[14]), .A2(b[14]), .Z(g[14]) );
  AN2D0 C1269 ( .A1(a[15]), .A2(b[15]), .Z(g[15]) );
  AN2D0 C1268 ( .A1(a[16]), .A2(b[16]), .Z(g[16]) );
  AN2D0 C1267 ( .A1(a[17]), .A2(b[17]), .Z(g[17]) );
  AN2D0 C1266 ( .A1(a[18]), .A2(b[18]), .Z(g[18]) );
  AN2D0 C1265 ( .A1(a[19]), .A2(b[19]), .Z(g[19]) );
  AN2D0 C1264 ( .A1(a[20]), .A2(b[20]), .Z(g[20]) );
  AN2D0 C1263 ( .A1(a[21]), .A2(b[21]), .Z(g[21]) );
  AN2D0 C1262 ( .A1(a[22]), .A2(b[22]), .Z(g[22]) );
  AN2D0 C1261 ( .A1(a[23]), .A2(b[23]), .Z(g[23]) );
  AN2D0 C1260 ( .A1(a[24]), .A2(b[24]), .Z(g[24]) );
  AN2D0 C1259 ( .A1(a[25]), .A2(b[25]), .Z(g[25]) );
  AN2D0 C1258 ( .A1(a[26]), .A2(b[26]), .Z(g[26]) );
  AN2D0 C1257 ( .A1(a[27]), .A2(b[27]), .Z(g[27]) );
  AN2D0 C1256 ( .A1(a[28]), .A2(b[28]), .Z(g[28]) );
  AN2D0 C1255 ( .A1(a[29]), .A2(b[29]), .Z(g[29]) );
  AN2D0 C1254 ( .A1(a[30]), .A2(b[30]), .Z(g[30]) );
  AN2D0 C1253 ( .A1(a[31]), .A2(b[31]), .Z(g[31]) );
  AN2D0 C1252 ( .A1(a[32]), .A2(b[32]), .Z(g[32]) );
  AN2D0 C1251 ( .A1(a[33]), .A2(b[33]), .Z(g[33]) );
  AN2D0 C1250 ( .A1(a[34]), .A2(b[34]), .Z(g[34]) );
  AN2D0 C1249 ( .A1(a[35]), .A2(b[35]), .Z(g[35]) );
  AN2D0 C1248 ( .A1(a[36]), .A2(b[36]), .Z(g[36]) );
  AN2D0 C1247 ( .A1(a[37]), .A2(b[37]), .Z(g[37]) );
  AN2D0 C1246 ( .A1(a[38]), .A2(b[38]), .Z(g[38]) );
  AN2D0 C1245 ( .A1(a[39]), .A2(b[39]), .Z(g[39]) );
  AN2D0 C1244 ( .A1(a[40]), .A2(b[40]), .Z(g[40]) );
  AN2D0 C1243 ( .A1(a[41]), .A2(b[41]), .Z(g[41]) );
  AN2D0 C1242 ( .A1(a[42]), .A2(b[42]), .Z(g[42]) );
  AN2D0 C1241 ( .A1(a[43]), .A2(b[43]), .Z(g[43]) );
  AN2D0 C1240 ( .A1(a[44]), .A2(b[44]), .Z(g[44]) );
  AN2D0 C1239 ( .A1(a[45]), .A2(b[45]), .Z(g[45]) );
  AN2D0 C1238 ( .A1(a[46]), .A2(b[46]), .Z(g[46]) );
  AN2D0 C1237 ( .A1(a[47]), .A2(b[47]), .Z(g[47]) );
  AN2D0 C1236 ( .A1(a[48]), .A2(b[48]), .Z(g[48]) );
  AN2D0 C1235 ( .A1(a[49]), .A2(b[49]), .Z(g[49]) );
  AN2D0 C1234 ( .A1(a[50]), .A2(b[50]), .Z(g[50]) );
  AN2D0 C1233 ( .A1(a[51]), .A2(b[51]), .Z(g[51]) );
  AN2D0 C1232 ( .A1(a[52]), .A2(b[52]), .Z(g[52]) );
  AN2D0 C1231 ( .A1(a[53]), .A2(b[53]), .Z(g[53]) );
  AN2D0 C1230 ( .A1(a[54]), .A2(b[54]), .Z(g[54]) );
  AN2D0 C1229 ( .A1(a[55]), .A2(b[55]), .Z(g[55]) );
  AN2D0 C1228 ( .A1(a[56]), .A2(b[56]), .Z(g[56]) );
  AN2D0 C1227 ( .A1(a[57]), .A2(b[57]), .Z(g[57]) );
  AN2D0 C1226 ( .A1(a[58]), .A2(b[58]), .Z(g[58]) );
  AN2D0 C1225 ( .A1(a[59]), .A2(b[59]), .Z(g[59]) );
  AN2D0 C1224 ( .A1(a[60]), .A2(b[60]), .Z(g[60]) );
  AN2D0 C1223 ( .A1(a[61]), .A2(b[61]), .Z(g[61]) );
  AN2D0 C1222 ( .A1(a[62]), .A2(b[62]), .Z(g[62]) );
  AN2D0 C1221 ( .A1(a[63]), .A2(b[63]), .Z(g[63]) );
  AN2D0 C1220 ( .A1(a[64]), .A2(b[64]), .Z(g[64]) );
  AN2D0 C1219 ( .A1(a[65]), .A2(b[65]), .Z(g[65]) );
  AN2D0 C1218 ( .A1(a[66]), .A2(b[66]), .Z(g[66]) );
  AN2D0 C1217 ( .A1(a[67]), .A2(b[67]), .Z(g[67]) );
  AN2D0 C1216 ( .A1(a[68]), .A2(b[68]), .Z(g[68]) );
  AN2D0 C1215 ( .A1(a[69]), .A2(b[69]), .Z(g[69]) );
  AN2D0 C1214 ( .A1(a[70]), .A2(b[70]), .Z(g[70]) );
  AN2D0 C1213 ( .A1(a[71]), .A2(b[71]), .Z(g[71]) );
  AN2D0 C1212 ( .A1(a[72]), .A2(b[72]), .Z(g[72]) );
  AN2D0 C1211 ( .A1(a[73]), .A2(b[73]), .Z(g[73]) );
  AN2D0 C1210 ( .A1(a[74]), .A2(b[74]), .Z(g[74]) );
  AN2D0 C1209 ( .A1(a[75]), .A2(b[75]), .Z(g[75]) );
  AN2D0 C1208 ( .A1(a[76]), .A2(b[76]), .Z(g[76]) );
  AN2D0 C1207 ( .A1(a[77]), .A2(b[77]), .Z(g[77]) );
  AN2D0 C1206 ( .A1(a[78]), .A2(b[78]), .Z(g[78]) );
  AN2D0 C1205 ( .A1(a[79]), .A2(b[79]), .Z(g[79]) );
  AN2D0 C1204 ( .A1(a[80]), .A2(b[80]), .Z(g[80]) );
  AN2D0 C1203 ( .A1(a[81]), .A2(b[81]), .Z(g[81]) );
  AN2D0 C1202 ( .A1(a[82]), .A2(b[82]), .Z(g[82]) );
  AN2D0 C1201 ( .A1(a[83]), .A2(b[83]), .Z(g[83]) );
  AN2D0 C1200 ( .A1(a[84]), .A2(b[84]), .Z(g[84]) );
  AN2D0 C1199 ( .A1(a[85]), .A2(b[85]), .Z(g[85]) );
  AN2D0 C1198 ( .A1(a[86]), .A2(b[86]), .Z(g[86]) );
  AN2D0 C1197 ( .A1(a[87]), .A2(b[87]), .Z(g[87]) );
  AN2D0 C1196 ( .A1(a[88]), .A2(b[88]), .Z(g[88]) );
  AN2D0 C1195 ( .A1(a[89]), .A2(b[89]), .Z(g[89]) );
  AN2D0 C1194 ( .A1(a[90]), .A2(b[90]), .Z(g[90]) );
  AN2D0 C1193 ( .A1(a[91]), .A2(b[91]), .Z(g[91]) );
  AN2D0 C1192 ( .A1(a[92]), .A2(b[92]), .Z(g[92]) );
  AN2D0 C1191 ( .A1(a[93]), .A2(b[93]), .Z(g[93]) );
  AN2D0 C1190 ( .A1(a[94]), .A2(b[94]), .Z(g[94]) );
  AN2D0 C1189 ( .A1(a[95]), .A2(b[95]), .Z(g[95]) );
  AN2D0 C1188 ( .A1(a[96]), .A2(b[96]), .Z(g[96]) );
  AN2D0 C1187 ( .A1(a[97]), .A2(b[97]), .Z(g[97]) );
  AN2D0 C1186 ( .A1(a[98]), .A2(b[98]), .Z(g[98]) );
  AN2D0 C1185 ( .A1(a[99]), .A2(b[99]), .Z(g[99]) );
  AN2D0 C1184 ( .A1(a[100]), .A2(b[100]), .Z(g[100]) );
  AN2D0 C1183 ( .A1(a[101]), .A2(b[101]), .Z(g[101]) );
  AN2D0 C1182 ( .A1(a[102]), .A2(b[102]), .Z(g[102]) );
  AN2D0 C1181 ( .A1(a[103]), .A2(b[103]), .Z(g[103]) );
  AN2D0 C1180 ( .A1(a[104]), .A2(b[104]), .Z(g[104]) );
  AN2D0 C1179 ( .A1(a[105]), .A2(b[105]), .Z(g[105]) );
  AN2D0 C1178 ( .A1(a[106]), .A2(b[106]), .Z(g[106]) );
  AN2D0 C1177 ( .A1(a[107]), .A2(b[107]), .Z(g[107]) );
  AN2D0 C1176 ( .A1(a[108]), .A2(b[108]), .Z(g[108]) );
  AN2D0 C1175 ( .A1(a[109]), .A2(b[109]), .Z(g[109]) );
  AN2D0 C1174 ( .A1(a[110]), .A2(b[110]), .Z(g[110]) );
  AN2D0 C1173 ( .A1(a[111]), .A2(b[111]), .Z(g[111]) );
  AN2D0 C1172 ( .A1(a[112]), .A2(b[112]), .Z(g[112]) );
  AN2D0 C1171 ( .A1(a[113]), .A2(b[113]), .Z(g[113]) );
  AN2D0 C1170 ( .A1(a[114]), .A2(b[114]), .Z(g[114]) );
  AN2D0 C1169 ( .A1(a[115]), .A2(b[115]), .Z(g[115]) );
  AN2D0 C1168 ( .A1(a[116]), .A2(b[116]), .Z(g[116]) );
  AN2D0 C1167 ( .A1(a[117]), .A2(b[117]), .Z(g[117]) );
  AN2D0 C1166 ( .A1(a[118]), .A2(b[118]), .Z(g[118]) );
  AN2D0 C1165 ( .A1(a[119]), .A2(b[119]), .Z(g[119]) );
  AN2D0 C1164 ( .A1(a[120]), .A2(b[120]), .Z(g[120]) );
  AN2D0 C1163 ( .A1(a[121]), .A2(b[121]), .Z(g[121]) );
  AN2D0 C1162 ( .A1(a[122]), .A2(b[122]), .Z(g[122]) );
  AN2D0 C1161 ( .A1(a[123]), .A2(b[123]), .Z(g[123]) );
  AN2D0 C1160 ( .A1(a[124]), .A2(b[124]), .Z(g[124]) );
  AN2D0 C1159 ( .A1(a[125]), .A2(b[125]), .Z(g[125]) );
  AN2D0 C1158 ( .A1(a[126]), .A2(b[126]), .Z(g[126]) );
  AN2D0 C1157 ( .A1(a[127]), .A2(b[127]), .Z(g[127]) );
  AN2D0 C1156 ( .A1(a[128]), .A2(b[128]), .Z(g[128]) );
  AN2D0 C1155 ( .A1(a[129]), .A2(b[129]), .Z(g[129]) );
  AN2D0 C1154 ( .A1(a[130]), .A2(b[130]), .Z(g[130]) );
  AN2D0 C1153 ( .A1(a[131]), .A2(b[131]), .Z(g[131]) );
  AN2D0 C1152 ( .A1(a[132]), .A2(b[132]), .Z(g[132]) );
  AN2D0 C1151 ( .A1(a[133]), .A2(b[133]), .Z(g[133]) );
  AN2D0 C1150 ( .A1(a[134]), .A2(b[134]), .Z(g[134]) );
  AN2D0 C1149 ( .A1(a[135]), .A2(b[135]), .Z(g[135]) );
  AN2D0 C1148 ( .A1(a[136]), .A2(b[136]), .Z(g[136]) );
  AN2D0 C1147 ( .A1(a[137]), .A2(b[137]), .Z(g[137]) );
  AN2D0 C1146 ( .A1(a[138]), .A2(b[138]), .Z(g[138]) );
  AN2D0 C1145 ( .A1(a[139]), .A2(b[139]), .Z(g[139]) );
  AN2D0 C1144 ( .A1(a[140]), .A2(b[140]), .Z(g[140]) );
  AN2D0 C1143 ( .A1(a[141]), .A2(b[141]), .Z(g[141]) );
  AN2D0 C1142 ( .A1(a[142]), .A2(b[142]), .Z(g[142]) );
  AN2D0 C1141 ( .A1(a[143]), .A2(b[143]), .Z(g[143]) );
  AN2D0 C1140 ( .A1(a[144]), .A2(b[144]), .Z(g[144]) );
  AN2D0 C1139 ( .A1(a[145]), .A2(b[145]), .Z(g[145]) );
  AN2D0 C1138 ( .A1(a[146]), .A2(b[146]), .Z(g[146]) );
  AN2D0 C1137 ( .A1(a[147]), .A2(b[147]), .Z(g[147]) );
  AN2D0 C1136 ( .A1(a[148]), .A2(b[148]), .Z(g[148]) );
  AN2D0 C1135 ( .A1(a[149]), .A2(b[149]), .Z(g[149]) );
  AN2D0 C1134 ( .A1(a[150]), .A2(b[150]), .Z(g[150]) );
  AN2D0 C1133 ( .A1(a[151]), .A2(b[151]), .Z(g[151]) );
  AN2D0 C1132 ( .A1(a[152]), .A2(b[152]), .Z(g[152]) );
  AN2D0 C1131 ( .A1(a[153]), .A2(b[153]), .Z(g[153]) );
  AN2D0 C1130 ( .A1(a[154]), .A2(b[154]), .Z(g[154]) );
  AN2D0 C1129 ( .A1(a[155]), .A2(b[155]), .Z(g[155]) );
  AN2D0 C1128 ( .A1(a[156]), .A2(b[156]), .Z(g[156]) );
  AN2D0 C1127 ( .A1(a[157]), .A2(b[157]), .Z(g[157]) );
  AN2D0 C1126 ( .A1(a[158]), .A2(b[158]), .Z(g[158]) );
  AN2D0 C1125 ( .A1(a[159]), .A2(b[159]), .Z(g[159]) );
  AN2D0 C1124 ( .A1(a[160]), .A2(b[160]), .Z(g[160]) );
  AN2D0 C1123 ( .A1(a[161]), .A2(b[161]), .Z(g[161]) );
  AN2D0 C1122 ( .A1(a[162]), .A2(b[162]), .Z(g[162]) );
  AN2D0 C1121 ( .A1(a[163]), .A2(b[163]), .Z(g[163]) );
  AN2D0 C1120 ( .A1(a[164]), .A2(b[164]), .Z(g[164]) );
  AN2D0 C1119 ( .A1(a[165]), .A2(b[165]), .Z(g[165]) );
  AN2D0 C1118 ( .A1(a[166]), .A2(b[166]), .Z(g[166]) );
  AN2D0 C1117 ( .A1(a[167]), .A2(b[167]), .Z(g[167]) );
  AN2D0 C1116 ( .A1(a[168]), .A2(b[168]), .Z(g[168]) );
  AN2D0 C1115 ( .A1(a[169]), .A2(b[169]), .Z(g[169]) );
  AN2D0 C1114 ( .A1(a[170]), .A2(b[170]), .Z(g[170]) );
  AN2D0 C1113 ( .A1(a[171]), .A2(b[171]), .Z(g[171]) );
  AN2D0 C1112 ( .A1(a[172]), .A2(b[172]), .Z(g[172]) );
  AN2D0 C1111 ( .A1(a[173]), .A2(b[173]), .Z(g[173]) );
  AN2D0 C1110 ( .A1(a[174]), .A2(b[174]), .Z(g[174]) );
  AN2D0 C1109 ( .A1(a[175]), .A2(b[175]), .Z(g[175]) );
  AN2D0 C1108 ( .A1(a[176]), .A2(b[176]), .Z(g[176]) );
  AN2D0 C1107 ( .A1(a[177]), .A2(b[177]), .Z(g[177]) );
  AN2D0 C1106 ( .A1(a[178]), .A2(b[178]), .Z(g[178]) );
  AN2D0 C1105 ( .A1(a[179]), .A2(b[179]), .Z(g[179]) );
  AN2D0 C1104 ( .A1(a[180]), .A2(b[180]), .Z(g[180]) );
  AN2D0 C1103 ( .A1(a[181]), .A2(b[181]), .Z(g[181]) );
  AN2D0 C1102 ( .A1(a[182]), .A2(b[182]), .Z(g[182]) );
  AN2D0 C1101 ( .A1(a[183]), .A2(b[183]), .Z(g[183]) );
  AN2D0 C1100 ( .A1(a[184]), .A2(b[184]), .Z(g[184]) );
  AN2D0 C1099 ( .A1(a[185]), .A2(b[185]), .Z(g[185]) );
  AN2D0 C1098 ( .A1(a[186]), .A2(b[186]), .Z(g[186]) );
  AN2D0 C1097 ( .A1(a[187]), .A2(b[187]), .Z(g[187]) );
  AN2D0 C1096 ( .A1(a[188]), .A2(b[188]), .Z(g[188]) );
  AN2D0 C1095 ( .A1(a[189]), .A2(b[189]), .Z(g[189]) );
  AN2D0 C1094 ( .A1(a[190]), .A2(b[190]), .Z(g[190]) );
  AN2D0 C1093 ( .A1(a[191]), .A2(b[191]), .Z(g[191]) );
  AN2D0 C1092 ( .A1(a[192]), .A2(b[192]), .Z(g[192]) );
  AN2D0 C1091 ( .A1(a[193]), .A2(b[193]), .Z(g[193]) );
  AN2D0 C1090 ( .A1(a[194]), .A2(b[194]), .Z(g[194]) );
  AN2D0 C1089 ( .A1(a[195]), .A2(b[195]), .Z(g[195]) );
  AN2D0 C1088 ( .A1(a[196]), .A2(b[196]), .Z(g[196]) );
  AN2D0 C1087 ( .A1(a[197]), .A2(b[197]), .Z(g[197]) );
  AN2D0 C1086 ( .A1(a[198]), .A2(b[198]), .Z(g[198]) );
  AN2D0 C1085 ( .A1(a[199]), .A2(b[199]), .Z(g[199]) );
  AN2D0 C1084 ( .A1(a[200]), .A2(b[200]), .Z(g[200]) );
  AN2D0 C1083 ( .A1(a[201]), .A2(b[201]), .Z(g[201]) );
  AN2D0 C1082 ( .A1(a[202]), .A2(b[202]), .Z(g[202]) );
  AN2D0 C1081 ( .A1(a[203]), .A2(b[203]), .Z(g[203]) );
  AN2D0 C1080 ( .A1(a[204]), .A2(b[204]), .Z(g[204]) );
  AN2D0 C1079 ( .A1(a[205]), .A2(b[205]), .Z(g[205]) );
  AN2D0 C1078 ( .A1(a[206]), .A2(b[206]), .Z(g[206]) );
  AN2D0 C1077 ( .A1(a[207]), .A2(b[207]), .Z(g[207]) );
  AN2D0 C1076 ( .A1(a[208]), .A2(b[208]), .Z(g[208]) );
  AN2D0 C1075 ( .A1(a[209]), .A2(b[209]), .Z(g[209]) );
  AN2D0 C1074 ( .A1(a[210]), .A2(b[210]), .Z(g[210]) );
  AN2D0 C1073 ( .A1(a[211]), .A2(b[211]), .Z(g[211]) );
  AN2D0 C1072 ( .A1(a[212]), .A2(b[212]), .Z(g[212]) );
  AN2D0 C1071 ( .A1(a[213]), .A2(b[213]), .Z(g[213]) );
  AN2D0 C1070 ( .A1(a[214]), .A2(b[214]), .Z(g[214]) );
  AN2D0 C1069 ( .A1(a[215]), .A2(b[215]), .Z(g[215]) );
  AN2D0 C1068 ( .A1(a[216]), .A2(b[216]), .Z(g[216]) );
  AN2D0 C1067 ( .A1(a[217]), .A2(b[217]), .Z(g[217]) );
  AN2D0 C1066 ( .A1(a[218]), .A2(b[218]), .Z(g[218]) );
  AN2D0 C1065 ( .A1(a[219]), .A2(b[219]), .Z(g[219]) );
  AN2D0 C1064 ( .A1(a[220]), .A2(b[220]), .Z(g[220]) );
  AN2D0 C1063 ( .A1(a[221]), .A2(b[221]), .Z(g[221]) );
  AN2D0 C1062 ( .A1(a[222]), .A2(b[222]), .Z(g[222]) );
  AN2D0 C1061 ( .A1(a[223]), .A2(b[223]), .Z(g[223]) );
  AN2D0 C1060 ( .A1(a[224]), .A2(b[224]), .Z(g[224]) );
  AN2D0 C1059 ( .A1(a[225]), .A2(b[225]), .Z(g[225]) );
  AN2D0 C1058 ( .A1(a[226]), .A2(b[226]), .Z(g[226]) );
  AN2D0 C1057 ( .A1(a[227]), .A2(b[227]), .Z(g[227]) );
  AN2D0 C1056 ( .A1(a[228]), .A2(b[228]), .Z(g[228]) );
  AN2D0 C1055 ( .A1(a[229]), .A2(b[229]), .Z(g[229]) );
  AN2D0 C1054 ( .A1(a[230]), .A2(b[230]), .Z(g[230]) );
  AN2D0 C1053 ( .A1(a[231]), .A2(b[231]), .Z(g[231]) );
  AN2D0 C1052 ( .A1(a[232]), .A2(b[232]), .Z(g[232]) );
  AN2D0 C1051 ( .A1(a[233]), .A2(b[233]), .Z(g[233]) );
  AN2D0 C1050 ( .A1(a[234]), .A2(b[234]), .Z(g[234]) );
  AN2D0 C1049 ( .A1(a[235]), .A2(b[235]), .Z(g[235]) );
  AN2D0 C1048 ( .A1(a[236]), .A2(b[236]), .Z(g[236]) );
  AN2D0 C1047 ( .A1(a[237]), .A2(b[237]), .Z(g[237]) );
  AN2D0 C1046 ( .A1(a[238]), .A2(b[238]), .Z(g[238]) );
  AN2D0 C1045 ( .A1(a[239]), .A2(b[239]), .Z(g[239]) );
  AN2D0 C1044 ( .A1(a[240]), .A2(b[240]), .Z(g[240]) );
  AN2D0 C1043 ( .A1(a[241]), .A2(b[241]), .Z(g[241]) );
  AN2D0 C1042 ( .A1(a[242]), .A2(b[242]), .Z(g[242]) );
  AN2D0 C1041 ( .A1(a[243]), .A2(b[243]), .Z(g[243]) );
  AN2D0 C1040 ( .A1(a[244]), .A2(b[244]), .Z(g[244]) );
  AN2D0 C1039 ( .A1(a[245]), .A2(b[245]), .Z(g[245]) );
  AN2D0 C1038 ( .A1(a[246]), .A2(b[246]), .Z(g[246]) );
  AN2D0 C1037 ( .A1(a[247]), .A2(b[247]), .Z(g[247]) );
  AN2D0 C1036 ( .A1(a[248]), .A2(b[248]), .Z(g[248]) );
  AN2D0 C1035 ( .A1(a[249]), .A2(b[249]), .Z(g[249]) );
  AN2D0 C1034 ( .A1(a[250]), .A2(b[250]), .Z(g[250]) );
  AN2D0 C1033 ( .A1(a[251]), .A2(b[251]), .Z(g[251]) );
  AN2D0 C1032 ( .A1(a[252]), .A2(b[252]), .Z(g[252]) );
  AN2D0 C1031 ( .A1(a[253]), .A2(b[253]), .Z(g[253]) );
  AN2D0 C1030 ( .A1(a[254]), .A2(b[254]), .Z(g[254]) );
endmodule

