
module gen_linear_part ( a, b, n, s );
  input [8:0] a;
  input [8:0] b;
  input [1011:0] n;
  output [8:0] s;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359;

  XOR3D0 U1 ( .A1(n1), .A2(n2), .A3(n[1011]), .Z(s[8]) );
  XOR4D0 U2 ( .A1(a[8]), .A2(n3), .A3(n[1006]), .A4(b[8]), .Z(n2) );
  XOR4D0 U3 ( .A1(n[1002]), .A2(n[1001]), .A3(n4), .A4(n5), .Z(n3) );
  XOR3D0 U4 ( .A1(n6), .A2(n7), .A3(n[1000]), .Z(n5) );
  XOR4D0 U5 ( .A1(n[992]), .A2(n8), .A3(n[994]), .A4(n[993]), .Z(n7) );
  XOR4D0 U6 ( .A1(n[987]), .A2(n[986]), .A3(n9), .A4(n10), .Z(n8) );
  XOR3D0 U7 ( .A1(n11), .A2(n12), .A3(n[985]), .Z(n10) );
  XOR4D0 U8 ( .A1(n[978]), .A2(n13), .A3(n[980]), .A4(n[979]), .Z(n12) );
  XOR4D0 U9 ( .A1(n[973]), .A2(n[972]), .A3(n14), .A4(n15), .Z(n13) );
  XOR3D0 U10 ( .A1(n16), .A2(n17), .A3(n[971]), .Z(n15) );
  XOR4D0 U11 ( .A1(n[964]), .A2(n18), .A3(n[966]), .A4(n[965]), .Z(n17) );
  XOR4D0 U12 ( .A1(n[959]), .A2(n[958]), .A3(n19), .A4(n20), .Z(n18) );
  XOR3D0 U13 ( .A1(n21), .A2(n22), .A3(n[957]), .Z(n20) );
  XOR4D0 U14 ( .A1(n[950]), .A2(n23), .A3(n[952]), .A4(n[951]), .Z(n22) );
  XOR4D0 U15 ( .A1(n[945]), .A2(n[944]), .A3(n24), .A4(n25), .Z(n23) );
  XOR3D0 U16 ( .A1(n26), .A2(n27), .A3(n[943]), .Z(n25) );
  XOR4D0 U17 ( .A1(n[936]), .A2(n28), .A3(n[938]), .A4(n[937]), .Z(n27) );
  XOR4D0 U18 ( .A1(n[931]), .A2(n[930]), .A3(n29), .A4(n30), .Z(n28) );
  XOR3D0 U19 ( .A1(n31), .A2(n32), .A3(n[929]), .Z(n30) );
  XOR4D0 U20 ( .A1(n[922]), .A2(n33), .A3(n[924]), .A4(n[923]), .Z(n32) );
  XOR4D0 U21 ( .A1(n[917]), .A2(n[916]), .A3(n34), .A4(n35), .Z(n33) );
  XOR3D0 U22 ( .A1(n36), .A2(n37), .A3(n[915]), .Z(n35) );
  XOR4D0 U23 ( .A1(n[908]), .A2(n38), .A3(n[910]), .A4(n[909]), .Z(n37) );
  XOR4D0 U24 ( .A1(n[903]), .A2(n[902]), .A3(n39), .A4(n40), .Z(n38) );
  XOR3D0 U25 ( .A1(n41), .A2(n42), .A3(n[901]), .Z(n40) );
  XOR4D0 U26 ( .A1(n[894]), .A2(n43), .A3(n[896]), .A4(n[895]), .Z(n42) );
  XOR4D0 U27 ( .A1(n[889]), .A2(n[888]), .A3(n44), .A4(n45), .Z(n43) );
  XOR3D0 U28 ( .A1(n46), .A2(n47), .A3(n[887]), .Z(n45) );
  XOR4D0 U29 ( .A1(n[880]), .A2(n48), .A3(n[882]), .A4(n[881]), .Z(n47) );
  XOR4D0 U30 ( .A1(n[875]), .A2(n[874]), .A3(n49), .A4(n50), .Z(n48) );
  XOR3D0 U31 ( .A1(n51), .A2(n52), .A3(n[873]), .Z(n50) );
  XOR4D0 U32 ( .A1(n[866]), .A2(n53), .A3(n[868]), .A4(n[867]), .Z(n52) );
  XOR4D0 U33 ( .A1(n[861]), .A2(n[860]), .A3(n54), .A4(n55), .Z(n53) );
  XOR3D0 U34 ( .A1(n56), .A2(n57), .A3(n[859]), .Z(n55) );
  XOR4D0 U35 ( .A1(n[852]), .A2(n58), .A3(n[854]), .A4(n[853]), .Z(n57) );
  XOR4D0 U36 ( .A1(n[847]), .A2(n[846]), .A3(n59), .A4(n60), .Z(n58) );
  XOR3D0 U37 ( .A1(n61), .A2(n62), .A3(n[845]), .Z(n60) );
  XOR4D0 U38 ( .A1(n[838]), .A2(n63), .A3(n[840]), .A4(n[839]), .Z(n62) );
  XOR4D0 U39 ( .A1(n[833]), .A2(n[832]), .A3(n64), .A4(n65), .Z(n63) );
  XOR3D0 U40 ( .A1(n66), .A2(n67), .A3(n[831]), .Z(n65) );
  XOR4D0 U41 ( .A1(n[824]), .A2(n68), .A3(n[826]), .A4(n[825]), .Z(n67) );
  XOR4D0 U42 ( .A1(n[819]), .A2(n[818]), .A3(n69), .A4(n70), .Z(n68) );
  XOR3D0 U43 ( .A1(n71), .A2(n72), .A3(n[817]), .Z(n70) );
  XOR4D0 U44 ( .A1(n[810]), .A2(n73), .A3(n[812]), .A4(n[811]), .Z(n72) );
  XOR4D0 U45 ( .A1(n[805]), .A2(n[804]), .A3(n74), .A4(n75), .Z(n73) );
  XOR3D0 U46 ( .A1(n76), .A2(n77), .A3(n[803]), .Z(n75) );
  XOR4D0 U47 ( .A1(n[796]), .A2(n78), .A3(n[798]), .A4(n[797]), .Z(n77) );
  XOR4D0 U48 ( .A1(n[791]), .A2(n[790]), .A3(n79), .A4(n80), .Z(n78) );
  XOR3D0 U49 ( .A1(n81), .A2(n82), .A3(n[789]), .Z(n80) );
  XOR4D0 U50 ( .A1(n[782]), .A2(n83), .A3(n[784]), .A4(n[783]), .Z(n82) );
  XOR4D0 U51 ( .A1(n[777]), .A2(n[776]), .A3(n84), .A4(n85), .Z(n83) );
  XOR3D0 U52 ( .A1(n86), .A2(n87), .A3(n[775]), .Z(n85) );
  XOR4D0 U53 ( .A1(n[768]), .A2(n88), .A3(n[770]), .A4(n[769]), .Z(n87) );
  XOR4D0 U54 ( .A1(n[763]), .A2(n[762]), .A3(n89), .A4(n90), .Z(n88) );
  XOR3D0 U55 ( .A1(n91), .A2(n92), .A3(n[761]), .Z(n90) );
  XOR4D0 U56 ( .A1(n[754]), .A2(n93), .A3(n[756]), .A4(n[755]), .Z(n92) );
  XOR4D0 U57 ( .A1(n[749]), .A2(n[748]), .A3(n94), .A4(n95), .Z(n93) );
  XOR3D0 U58 ( .A1(n96), .A2(n97), .A3(n[747]), .Z(n95) );
  XOR4D0 U59 ( .A1(n[740]), .A2(n98), .A3(n[742]), .A4(n[741]), .Z(n97) );
  XOR4D0 U60 ( .A1(n[735]), .A2(n[734]), .A3(n99), .A4(n100), .Z(n98) );
  XOR3D0 U61 ( .A1(n101), .A2(n102), .A3(n[733]), .Z(n100) );
  XOR4D0 U62 ( .A1(n[726]), .A2(n103), .A3(n[728]), .A4(n[727]), .Z(n102) );
  XOR4D0 U63 ( .A1(n[721]), .A2(n[720]), .A3(n104), .A4(n105), .Z(n103) );
  XOR3D0 U64 ( .A1(n106), .A2(n107), .A3(n[719]), .Z(n105) );
  XOR4D0 U65 ( .A1(n[712]), .A2(n108), .A3(n[714]), .A4(n[713]), .Z(n107) );
  XOR4D0 U66 ( .A1(n[707]), .A2(n[706]), .A3(n109), .A4(n110), .Z(n108) );
  XOR3D0 U67 ( .A1(n111), .A2(n112), .A3(n[705]), .Z(n110) );
  XOR4D0 U68 ( .A1(n[698]), .A2(n113), .A3(n[700]), .A4(n[699]), .Z(n112) );
  XOR4D0 U69 ( .A1(n[693]), .A2(n[692]), .A3(n114), .A4(n115), .Z(n113) );
  XOR3D0 U70 ( .A1(n116), .A2(n117), .A3(n[691]), .Z(n115) );
  XOR4D0 U71 ( .A1(n[684]), .A2(n118), .A3(n[686]), .A4(n[685]), .Z(n117) );
  XOR4D0 U72 ( .A1(n[679]), .A2(n[678]), .A3(n119), .A4(n120), .Z(n118) );
  XOR3D0 U73 ( .A1(n121), .A2(n122), .A3(n[677]), .Z(n120) );
  XOR4D0 U74 ( .A1(n[670]), .A2(n123), .A3(n[672]), .A4(n[671]), .Z(n122) );
  XOR4D0 U75 ( .A1(n[665]), .A2(n[664]), .A3(n124), .A4(n125), .Z(n123) );
  XOR3D0 U76 ( .A1(n126), .A2(n127), .A3(n[663]), .Z(n125) );
  XOR4D0 U77 ( .A1(n[656]), .A2(n128), .A3(n[658]), .A4(n[657]), .Z(n127) );
  XOR4D0 U78 ( .A1(n[651]), .A2(n[650]), .A3(n129), .A4(n130), .Z(n128) );
  XOR3D0 U79 ( .A1(n131), .A2(n132), .A3(n[649]), .Z(n130) );
  XOR4D0 U80 ( .A1(n[642]), .A2(n133), .A3(n[644]), .A4(n[643]), .Z(n132) );
  XOR4D0 U81 ( .A1(n[637]), .A2(n[636]), .A3(n134), .A4(n135), .Z(n133) );
  XOR3D0 U82 ( .A1(n136), .A2(n137), .A3(n[635]), .Z(n135) );
  XOR4D0 U83 ( .A1(n[628]), .A2(n138), .A3(n[630]), .A4(n[629]), .Z(n137) );
  XOR4D0 U84 ( .A1(n[623]), .A2(n[622]), .A3(n139), .A4(n140), .Z(n138) );
  XOR3D0 U85 ( .A1(n141), .A2(n142), .A3(n[621]), .Z(n140) );
  XOR4D0 U86 ( .A1(n[614]), .A2(n143), .A3(n[616]), .A4(n[615]), .Z(n142) );
  XOR4D0 U87 ( .A1(n[609]), .A2(n[608]), .A3(n144), .A4(n145), .Z(n143) );
  XOR3D0 U88 ( .A1(n146), .A2(n147), .A3(n[607]), .Z(n145) );
  XOR4D0 U89 ( .A1(n[600]), .A2(n148), .A3(n[602]), .A4(n[601]), .Z(n147) );
  XOR4D0 U90 ( .A1(n[595]), .A2(n[594]), .A3(n149), .A4(n150), .Z(n148) );
  XOR3D0 U91 ( .A1(n151), .A2(n152), .A3(n[593]), .Z(n150) );
  XOR4D0 U92 ( .A1(n[586]), .A2(n153), .A3(n[588]), .A4(n[587]), .Z(n152) );
  XOR4D0 U93 ( .A1(n[581]), .A2(n[580]), .A3(n154), .A4(n155), .Z(n153) );
  XOR3D0 U94 ( .A1(n156), .A2(n157), .A3(n[579]), .Z(n155) );
  XOR4D0 U95 ( .A1(n[572]), .A2(n158), .A3(n[574]), .A4(n[573]), .Z(n157) );
  XOR4D0 U96 ( .A1(n[567]), .A2(n[566]), .A3(n159), .A4(n160), .Z(n158) );
  XOR3D0 U97 ( .A1(n161), .A2(n162), .A3(n[565]), .Z(n160) );
  XOR4D0 U98 ( .A1(n[558]), .A2(n163), .A3(n[560]), .A4(n[559]), .Z(n162) );
  XOR4D0 U99 ( .A1(n[553]), .A2(n[552]), .A3(n164), .A4(n165), .Z(n163) );
  XOR3D0 U100 ( .A1(n166), .A2(n167), .A3(n[551]), .Z(n165) );
  XOR4D0 U101 ( .A1(n[544]), .A2(n168), .A3(n[546]), .A4(n[545]), .Z(n167) );
  XOR4D0 U102 ( .A1(n[539]), .A2(n[538]), .A3(n169), .A4(n170), .Z(n168) );
  XOR3D0 U103 ( .A1(n171), .A2(n172), .A3(n[537]), .Z(n170) );
  XOR4D0 U104 ( .A1(n[530]), .A2(n173), .A3(n[532]), .A4(n[531]), .Z(n172) );
  XOR4D0 U105 ( .A1(n[525]), .A2(n[524]), .A3(n174), .A4(n175), .Z(n173) );
  XOR3D0 U106 ( .A1(n176), .A2(n177), .A3(n[523]), .Z(n175) );
  XOR4D0 U107 ( .A1(n[516]), .A2(n178), .A3(n[518]), .A4(n[517]), .Z(n177) );
  XOR4D0 U108 ( .A1(n[511]), .A2(n[510]), .A3(n179), .A4(n180), .Z(n178) );
  XOR3D0 U109 ( .A1(n181), .A2(n182), .A3(n[509]), .Z(n180) );
  XOR4D0 U110 ( .A1(n[502]), .A2(n[501]), .A3(n[504]), .A4(n[503]), .Z(n182)
         );
  XOR4D0 U111 ( .A1(n[506]), .A2(n[505]), .A3(n[508]), .A4(n[507]), .Z(n181)
         );
  XOR4D0 U112 ( .A1(n[513]), .A2(n[512]), .A3(n[515]), .A4(n[514]), .Z(n179)
         );
  XOR4D0 U113 ( .A1(n[520]), .A2(n[519]), .A3(n[522]), .A4(n[521]), .Z(n176)
         );
  XOR4D0 U114 ( .A1(n[527]), .A2(n[526]), .A3(n[529]), .A4(n[528]), .Z(n174)
         );
  XOR4D0 U115 ( .A1(n[534]), .A2(n[533]), .A3(n[536]), .A4(n[535]), .Z(n171)
         );
  XOR4D0 U116 ( .A1(n[541]), .A2(n[540]), .A3(n[543]), .A4(n[542]), .Z(n169)
         );
  XOR4D0 U117 ( .A1(n[548]), .A2(n[547]), .A3(n[550]), .A4(n[549]), .Z(n166)
         );
  XOR4D0 U118 ( .A1(n[555]), .A2(n[554]), .A3(n[557]), .A4(n[556]), .Z(n164)
         );
  XOR4D0 U119 ( .A1(n[562]), .A2(n[561]), .A3(n[564]), .A4(n[563]), .Z(n161)
         );
  XOR4D0 U120 ( .A1(n[569]), .A2(n[568]), .A3(n[571]), .A4(n[570]), .Z(n159)
         );
  XOR4D0 U121 ( .A1(n[576]), .A2(n[575]), .A3(n[578]), .A4(n[577]), .Z(n156)
         );
  XOR4D0 U122 ( .A1(n[583]), .A2(n[582]), .A3(n[585]), .A4(n[584]), .Z(n154)
         );
  XOR4D0 U123 ( .A1(n[590]), .A2(n[589]), .A3(n[592]), .A4(n[591]), .Z(n151)
         );
  XOR4D0 U124 ( .A1(n[597]), .A2(n[596]), .A3(n[599]), .A4(n[598]), .Z(n149)
         );
  XOR4D0 U125 ( .A1(n[604]), .A2(n[603]), .A3(n[606]), .A4(n[605]), .Z(n146)
         );
  XOR4D0 U126 ( .A1(n[611]), .A2(n[610]), .A3(n[613]), .A4(n[612]), .Z(n144)
         );
  XOR4D0 U127 ( .A1(n[618]), .A2(n[617]), .A3(n[620]), .A4(n[619]), .Z(n141)
         );
  XOR4D0 U128 ( .A1(n[625]), .A2(n[624]), .A3(n[627]), .A4(n[626]), .Z(n139)
         );
  XOR4D0 U129 ( .A1(n[632]), .A2(n[631]), .A3(n[634]), .A4(n[633]), .Z(n136)
         );
  XOR4D0 U130 ( .A1(n[639]), .A2(n[638]), .A3(n[641]), .A4(n[640]), .Z(n134)
         );
  XOR4D0 U131 ( .A1(n[646]), .A2(n[645]), .A3(n[648]), .A4(n[647]), .Z(n131)
         );
  XOR4D0 U132 ( .A1(n[653]), .A2(n[652]), .A3(n[655]), .A4(n[654]), .Z(n129)
         );
  XOR4D0 U133 ( .A1(n[660]), .A2(n[659]), .A3(n[662]), .A4(n[661]), .Z(n126)
         );
  XOR4D0 U134 ( .A1(n[667]), .A2(n[666]), .A3(n[669]), .A4(n[668]), .Z(n124)
         );
  XOR4D0 U135 ( .A1(n[674]), .A2(n[673]), .A3(n[676]), .A4(n[675]), .Z(n121)
         );
  XOR4D0 U136 ( .A1(n[681]), .A2(n[680]), .A3(n[683]), .A4(n[682]), .Z(n119)
         );
  XOR4D0 U137 ( .A1(n[688]), .A2(n[687]), .A3(n[690]), .A4(n[689]), .Z(n116)
         );
  XOR4D0 U138 ( .A1(n[695]), .A2(n[694]), .A3(n[697]), .A4(n[696]), .Z(n114)
         );
  XOR4D0 U139 ( .A1(n[702]), .A2(n[701]), .A3(n[704]), .A4(n[703]), .Z(n111)
         );
  XOR4D0 U140 ( .A1(n[709]), .A2(n[708]), .A3(n[711]), .A4(n[710]), .Z(n109)
         );
  XOR4D0 U141 ( .A1(n[716]), .A2(n[715]), .A3(n[718]), .A4(n[717]), .Z(n106)
         );
  XOR4D0 U142 ( .A1(n[723]), .A2(n[722]), .A3(n[725]), .A4(n[724]), .Z(n104)
         );
  XOR4D0 U143 ( .A1(n[730]), .A2(n[729]), .A3(n[732]), .A4(n[731]), .Z(n101)
         );
  XOR4D0 U144 ( .A1(n[737]), .A2(n[736]), .A3(n[739]), .A4(n[738]), .Z(n99) );
  XOR4D0 U145 ( .A1(n[744]), .A2(n[743]), .A3(n[746]), .A4(n[745]), .Z(n96) );
  XOR4D0 U146 ( .A1(n[751]), .A2(n[750]), .A3(n[753]), .A4(n[752]), .Z(n94) );
  XOR4D0 U147 ( .A1(n[758]), .A2(n[757]), .A3(n[760]), .A4(n[759]), .Z(n91) );
  XOR4D0 U148 ( .A1(n[765]), .A2(n[764]), .A3(n[767]), .A4(n[766]), .Z(n89) );
  XOR4D0 U149 ( .A1(n[772]), .A2(n[771]), .A3(n[774]), .A4(n[773]), .Z(n86) );
  XOR4D0 U150 ( .A1(n[779]), .A2(n[778]), .A3(n[781]), .A4(n[780]), .Z(n84) );
  XOR4D0 U151 ( .A1(n[786]), .A2(n[785]), .A3(n[788]), .A4(n[787]), .Z(n81) );
  XOR4D0 U152 ( .A1(n[793]), .A2(n[792]), .A3(n[795]), .A4(n[794]), .Z(n79) );
  XOR4D0 U153 ( .A1(n[800]), .A2(n[799]), .A3(n[802]), .A4(n[801]), .Z(n76) );
  XOR4D0 U154 ( .A1(n[807]), .A2(n[806]), .A3(n[809]), .A4(n[808]), .Z(n74) );
  XOR4D0 U155 ( .A1(n[814]), .A2(n[813]), .A3(n[816]), .A4(n[815]), .Z(n71) );
  XOR4D0 U156 ( .A1(n[821]), .A2(n[820]), .A3(n[823]), .A4(n[822]), .Z(n69) );
  XOR4D0 U157 ( .A1(n[828]), .A2(n[827]), .A3(n[830]), .A4(n[829]), .Z(n66) );
  XOR4D0 U158 ( .A1(n[835]), .A2(n[834]), .A3(n[837]), .A4(n[836]), .Z(n64) );
  XOR4D0 U159 ( .A1(n[842]), .A2(n[841]), .A3(n[844]), .A4(n[843]), .Z(n61) );
  XOR4D0 U160 ( .A1(n[849]), .A2(n[848]), .A3(n[851]), .A4(n[850]), .Z(n59) );
  XOR4D0 U161 ( .A1(n[856]), .A2(n[855]), .A3(n[858]), .A4(n[857]), .Z(n56) );
  XOR4D0 U162 ( .A1(n[863]), .A2(n[862]), .A3(n[865]), .A4(n[864]), .Z(n54) );
  XOR4D0 U163 ( .A1(n[870]), .A2(n[869]), .A3(n[872]), .A4(n[871]), .Z(n51) );
  XOR4D0 U164 ( .A1(n[877]), .A2(n[876]), .A3(n[879]), .A4(n[878]), .Z(n49) );
  XOR4D0 U165 ( .A1(n[884]), .A2(n[883]), .A3(n[886]), .A4(n[885]), .Z(n46) );
  XOR4D0 U166 ( .A1(n[891]), .A2(n[890]), .A3(n[893]), .A4(n[892]), .Z(n44) );
  XOR4D0 U167 ( .A1(n[898]), .A2(n[897]), .A3(n[900]), .A4(n[899]), .Z(n41) );
  XOR4D0 U168 ( .A1(n[905]), .A2(n[904]), .A3(n[907]), .A4(n[906]), .Z(n39) );
  XOR4D0 U169 ( .A1(n[912]), .A2(n[911]), .A3(n[914]), .A4(n[913]), .Z(n36) );
  XOR4D0 U170 ( .A1(n[919]), .A2(n[918]), .A3(n[921]), .A4(n[920]), .Z(n34) );
  XOR4D0 U171 ( .A1(n[926]), .A2(n[925]), .A3(n[928]), .A4(n[927]), .Z(n31) );
  XOR4D0 U172 ( .A1(n[933]), .A2(n[932]), .A3(n[935]), .A4(n[934]), .Z(n29) );
  XOR4D0 U173 ( .A1(n[940]), .A2(n[939]), .A3(n[942]), .A4(n[941]), .Z(n26) );
  XOR4D0 U174 ( .A1(n[947]), .A2(n[946]), .A3(n[949]), .A4(n[948]), .Z(n24) );
  XOR4D0 U175 ( .A1(n[954]), .A2(n[953]), .A3(n[956]), .A4(n[955]), .Z(n21) );
  XOR4D0 U176 ( .A1(n[961]), .A2(n[960]), .A3(n[963]), .A4(n[962]), .Z(n19) );
  XOR4D0 U177 ( .A1(n[968]), .A2(n[967]), .A3(n[970]), .A4(n[969]), .Z(n16) );
  XOR4D0 U178 ( .A1(n[975]), .A2(n[974]), .A3(n[977]), .A4(n[976]), .Z(n14) );
  XOR4D0 U179 ( .A1(n[982]), .A2(n[981]), .A3(n[984]), .A4(n[983]), .Z(n11) );
  XOR4D0 U180 ( .A1(n[989]), .A2(n[988]), .A3(n[991]), .A4(n[990]), .Z(n9) );
  XOR4D0 U181 ( .A1(n[996]), .A2(n[995]), .A3(n[998]), .A4(n[997]), .Z(n6) );
  XOR4D0 U182 ( .A1(n[1004]), .A2(n[1003]), .A3(n[999]), .A4(n[1005]), .Z(n4)
         );
  XOR4D0 U183 ( .A1(n[1008]), .A2(n[1007]), .A3(n[1010]), .A4(n[1009]), .Z(n1)
         );
  XOR4D0 U184 ( .A1(n183), .A2(n184), .A3(n185), .A4(n[495]), .Z(s[7]) );
  XOR3D0 U185 ( .A1(n[498]), .A2(n[497]), .A3(n[496]), .Z(n185) );
  XOR4D0 U186 ( .A1(a[7]), .A2(n186), .A3(n[492]), .A4(b[7]), .Z(n184) );
  XOR4D0 U187 ( .A1(n[487]), .A2(n[486]), .A3(n187), .A4(n188), .Z(n186) );
  XOR3D0 U188 ( .A1(n189), .A2(n190), .A3(n[485]), .Z(n188) );
  XOR4D0 U189 ( .A1(n[478]), .A2(n191), .A3(n[480]), .A4(n[479]), .Z(n190) );
  XOR4D0 U190 ( .A1(n[473]), .A2(n[472]), .A3(n192), .A4(n193), .Z(n191) );
  XOR3D0 U191 ( .A1(n194), .A2(n195), .A3(n[471]), .Z(n193) );
  XOR4D0 U192 ( .A1(n[464]), .A2(n196), .A3(n[466]), .A4(n[465]), .Z(n195) );
  XOR4D0 U193 ( .A1(n[459]), .A2(n[458]), .A3(n197), .A4(n198), .Z(n196) );
  XOR3D0 U194 ( .A1(n199), .A2(n200), .A3(n[457]), .Z(n198) );
  XOR4D0 U195 ( .A1(n[450]), .A2(n201), .A3(n[452]), .A4(n[451]), .Z(n200) );
  XOR4D0 U196 ( .A1(n[445]), .A2(n[444]), .A3(n202), .A4(n203), .Z(n201) );
  XOR3D0 U197 ( .A1(n204), .A2(n205), .A3(n[443]), .Z(n203) );
  XOR4D0 U198 ( .A1(n[436]), .A2(n206), .A3(n[438]), .A4(n[437]), .Z(n205) );
  XOR4D0 U199 ( .A1(n[431]), .A2(n[430]), .A3(n207), .A4(n208), .Z(n206) );
  XOR3D0 U200 ( .A1(n209), .A2(n210), .A3(n[429]), .Z(n208) );
  XOR4D0 U201 ( .A1(n[422]), .A2(n211), .A3(n[424]), .A4(n[423]), .Z(n210) );
  XOR4D0 U202 ( .A1(n[417]), .A2(n[416]), .A3(n212), .A4(n213), .Z(n211) );
  XOR3D0 U203 ( .A1(n214), .A2(n215), .A3(n[415]), .Z(n213) );
  XOR4D0 U204 ( .A1(n[408]), .A2(n216), .A3(n[410]), .A4(n[409]), .Z(n215) );
  XOR4D0 U205 ( .A1(n[403]), .A2(n[402]), .A3(n217), .A4(n218), .Z(n216) );
  XOR3D0 U206 ( .A1(n219), .A2(n220), .A3(n[401]), .Z(n218) );
  XOR4D0 U207 ( .A1(n[394]), .A2(n221), .A3(n[396]), .A4(n[395]), .Z(n220) );
  XOR4D0 U208 ( .A1(n[389]), .A2(n[388]), .A3(n222), .A4(n223), .Z(n221) );
  XOR3D0 U209 ( .A1(n224), .A2(n225), .A3(n[387]), .Z(n223) );
  XOR4D0 U210 ( .A1(n[380]), .A2(n226), .A3(n[382]), .A4(n[381]), .Z(n225) );
  XOR4D0 U211 ( .A1(n[375]), .A2(n[374]), .A3(n227), .A4(n228), .Z(n226) );
  XOR3D0 U212 ( .A1(n229), .A2(n230), .A3(n[373]), .Z(n228) );
  XOR4D0 U213 ( .A1(n[366]), .A2(n231), .A3(n[368]), .A4(n[367]), .Z(n230) );
  XOR4D0 U214 ( .A1(n[361]), .A2(n[360]), .A3(n232), .A4(n233), .Z(n231) );
  XOR3D0 U215 ( .A1(n234), .A2(n235), .A3(n[359]), .Z(n233) );
  XOR4D0 U216 ( .A1(n[352]), .A2(n236), .A3(n[354]), .A4(n[353]), .Z(n235) );
  XOR4D0 U217 ( .A1(n[347]), .A2(n[346]), .A3(n237), .A4(n238), .Z(n236) );
  XOR3D0 U218 ( .A1(n239), .A2(n240), .A3(n[345]), .Z(n238) );
  XOR4D0 U219 ( .A1(n[338]), .A2(n241), .A3(n[340]), .A4(n[339]), .Z(n240) );
  XOR4D0 U220 ( .A1(n[333]), .A2(n[332]), .A3(n242), .A4(n243), .Z(n241) );
  XOR3D0 U221 ( .A1(n244), .A2(n245), .A3(n[331]), .Z(n243) );
  XOR4D0 U222 ( .A1(n[324]), .A2(n246), .A3(n[326]), .A4(n[325]), .Z(n245) );
  XOR4D0 U223 ( .A1(n[319]), .A2(n[318]), .A3(n247), .A4(n248), .Z(n246) );
  XOR3D0 U224 ( .A1(n249), .A2(n250), .A3(n[317]), .Z(n248) );
  XOR4D0 U225 ( .A1(n[310]), .A2(n251), .A3(n[312]), .A4(n[311]), .Z(n250) );
  XOR4D0 U226 ( .A1(n[305]), .A2(n[304]), .A3(n252), .A4(n253), .Z(n251) );
  XOR3D0 U227 ( .A1(n254), .A2(n255), .A3(n[303]), .Z(n253) );
  XOR4D0 U228 ( .A1(n[296]), .A2(n256), .A3(n[298]), .A4(n[297]), .Z(n255) );
  XOR4D0 U229 ( .A1(n[291]), .A2(n[290]), .A3(n257), .A4(n258), .Z(n256) );
  XOR3D0 U230 ( .A1(n259), .A2(n260), .A3(n[289]), .Z(n258) );
  XOR4D0 U231 ( .A1(n[282]), .A2(n261), .A3(n[284]), .A4(n[283]), .Z(n260) );
  XOR4D0 U232 ( .A1(n[277]), .A2(n[276]), .A3(n262), .A4(n263), .Z(n261) );
  XOR3D0 U233 ( .A1(n264), .A2(n265), .A3(n[275]), .Z(n263) );
  XOR4D0 U234 ( .A1(n[268]), .A2(n266), .A3(n[270]), .A4(n[269]), .Z(n265) );
  XOR4D0 U235 ( .A1(n[263]), .A2(n[262]), .A3(n267), .A4(n268), .Z(n266) );
  XOR3D0 U236 ( .A1(n269), .A2(n270), .A3(n[261]), .Z(n268) );
  XOR3D0 U237 ( .A1(n[256]), .A2(n[255]), .A3(n271), .Z(n270) );
  XOR3D0 U238 ( .A1(n272), .A2(n273), .A3(n[254]), .Z(n271) );
  XOR4D0 U239 ( .A1(n[247]), .A2(n[246]), .A3(n[249]), .A4(n[248]), .Z(n273)
         );
  XOR4D0 U240 ( .A1(n[251]), .A2(n[250]), .A3(n[253]), .A4(n[252]), .Z(n272)
         );
  XOR4D0 U241 ( .A1(n[258]), .A2(n[257]), .A3(n[260]), .A4(n[259]), .Z(n269)
         );
  XOR4D0 U242 ( .A1(n[265]), .A2(n[264]), .A3(n[267]), .A4(n[266]), .Z(n267)
         );
  XOR4D0 U243 ( .A1(n[272]), .A2(n[271]), .A3(n[274]), .A4(n[273]), .Z(n264)
         );
  XOR4D0 U244 ( .A1(n[279]), .A2(n[278]), .A3(n[281]), .A4(n[280]), .Z(n262)
         );
  XOR4D0 U245 ( .A1(n[286]), .A2(n[285]), .A3(n[288]), .A4(n[287]), .Z(n259)
         );
  XOR4D0 U246 ( .A1(n[293]), .A2(n[292]), .A3(n[295]), .A4(n[294]), .Z(n257)
         );
  XOR4D0 U247 ( .A1(n[300]), .A2(n[299]), .A3(n[302]), .A4(n[301]), .Z(n254)
         );
  XOR4D0 U248 ( .A1(n[307]), .A2(n[306]), .A3(n[309]), .A4(n[308]), .Z(n252)
         );
  XOR4D0 U249 ( .A1(n[314]), .A2(n[313]), .A3(n[316]), .A4(n[315]), .Z(n249)
         );
  XOR4D0 U250 ( .A1(n[321]), .A2(n[320]), .A3(n[323]), .A4(n[322]), .Z(n247)
         );
  XOR4D0 U251 ( .A1(n[328]), .A2(n[327]), .A3(n[330]), .A4(n[329]), .Z(n244)
         );
  XOR4D0 U252 ( .A1(n[335]), .A2(n[334]), .A3(n[337]), .A4(n[336]), .Z(n242)
         );
  XOR4D0 U253 ( .A1(n[342]), .A2(n[341]), .A3(n[344]), .A4(n[343]), .Z(n239)
         );
  XOR4D0 U254 ( .A1(n[349]), .A2(n[348]), .A3(n[351]), .A4(n[350]), .Z(n237)
         );
  XOR4D0 U255 ( .A1(n[356]), .A2(n[355]), .A3(n[358]), .A4(n[357]), .Z(n234)
         );
  XOR4D0 U256 ( .A1(n[363]), .A2(n[362]), .A3(n[365]), .A4(n[364]), .Z(n232)
         );
  XOR4D0 U257 ( .A1(n[370]), .A2(n[369]), .A3(n[372]), .A4(n[371]), .Z(n229)
         );
  XOR4D0 U258 ( .A1(n[377]), .A2(n[376]), .A3(n[379]), .A4(n[378]), .Z(n227)
         );
  XOR4D0 U259 ( .A1(n[384]), .A2(n[383]), .A3(n[386]), .A4(n[385]), .Z(n224)
         );
  XOR4D0 U260 ( .A1(n[391]), .A2(n[390]), .A3(n[393]), .A4(n[392]), .Z(n222)
         );
  XOR4D0 U261 ( .A1(n[398]), .A2(n[397]), .A3(n[400]), .A4(n[399]), .Z(n219)
         );
  XOR4D0 U262 ( .A1(n[405]), .A2(n[404]), .A3(n[407]), .A4(n[406]), .Z(n217)
         );
  XOR4D0 U263 ( .A1(n[412]), .A2(n[411]), .A3(n[414]), .A4(n[413]), .Z(n214)
         );
  XOR4D0 U264 ( .A1(n[419]), .A2(n[418]), .A3(n[421]), .A4(n[420]), .Z(n212)
         );
  XOR4D0 U265 ( .A1(n[426]), .A2(n[425]), .A3(n[428]), .A4(n[427]), .Z(n209)
         );
  XOR4D0 U266 ( .A1(n[433]), .A2(n[432]), .A3(n[435]), .A4(n[434]), .Z(n207)
         );
  XOR4D0 U267 ( .A1(n[440]), .A2(n[439]), .A3(n[442]), .A4(n[441]), .Z(n204)
         );
  XOR4D0 U268 ( .A1(n[447]), .A2(n[446]), .A3(n[449]), .A4(n[448]), .Z(n202)
         );
  XOR4D0 U269 ( .A1(n[454]), .A2(n[453]), .A3(n[456]), .A4(n[455]), .Z(n199)
         );
  XOR4D0 U270 ( .A1(n[461]), .A2(n[460]), .A3(n[463]), .A4(n[462]), .Z(n197)
         );
  XOR4D0 U271 ( .A1(n[468]), .A2(n[467]), .A3(n[470]), .A4(n[469]), .Z(n194)
         );
  XOR4D0 U272 ( .A1(n[475]), .A2(n[474]), .A3(n[477]), .A4(n[476]), .Z(n192)
         );
  XOR4D0 U273 ( .A1(n[482]), .A2(n[481]), .A3(n[484]), .A4(n[483]), .Z(n189)
         );
  XOR4D0 U274 ( .A1(n[489]), .A2(n[488]), .A3(n[491]), .A4(n[490]), .Z(n187)
         );
  XOR4D0 U275 ( .A1(n[494]), .A2(n[493]), .A3(n[500]), .A4(n[499]), .Z(n183)
         );
  XOR4D0 U276 ( .A1(b[6]), .A2(a[6]), .A3(n274), .A4(n275), .Z(s[6]) );
  XOR4D0 U277 ( .A1(n[239]), .A2(n276), .A3(n[241]), .A4(n[240]), .Z(n275) );
  XOR4D0 U278 ( .A1(n[234]), .A2(n[233]), .A3(n277), .A4(n278), .Z(n276) );
  XOR3D0 U279 ( .A1(n279), .A2(n280), .A3(n[232]), .Z(n278) );
  XOR4D0 U280 ( .A1(n[225]), .A2(n281), .A3(n[227]), .A4(n[226]), .Z(n280) );
  XOR4D0 U281 ( .A1(n[220]), .A2(n[219]), .A3(n282), .A4(n283), .Z(n281) );
  XOR3D0 U282 ( .A1(n284), .A2(n285), .A3(n[218]), .Z(n283) );
  XOR4D0 U283 ( .A1(n[211]), .A2(n286), .A3(n[213]), .A4(n[212]), .Z(n285) );
  XOR4D0 U284 ( .A1(n[206]), .A2(n[205]), .A3(n287), .A4(n288), .Z(n286) );
  XOR3D0 U285 ( .A1(n289), .A2(n290), .A3(n[204]), .Z(n288) );
  XOR4D0 U286 ( .A1(n[197]), .A2(n291), .A3(n[199]), .A4(n[198]), .Z(n290) );
  XOR4D0 U287 ( .A1(n[192]), .A2(n[191]), .A3(n292), .A4(n293), .Z(n291) );
  XOR3D0 U288 ( .A1(n294), .A2(n295), .A3(n[190]), .Z(n293) );
  XOR4D0 U289 ( .A1(n[183]), .A2(n296), .A3(n[185]), .A4(n[184]), .Z(n295) );
  XOR4D0 U290 ( .A1(n[178]), .A2(n[177]), .A3(n297), .A4(n298), .Z(n296) );
  XOR3D0 U291 ( .A1(n299), .A2(n300), .A3(n[176]), .Z(n298) );
  XOR4D0 U292 ( .A1(n[169]), .A2(n301), .A3(n[171]), .A4(n[170]), .Z(n300) );
  XOR4D0 U293 ( .A1(n[164]), .A2(n[163]), .A3(n302), .A4(n303), .Z(n301) );
  XOR3D0 U294 ( .A1(n304), .A2(n305), .A3(n[162]), .Z(n303) );
  XOR4D0 U295 ( .A1(n[155]), .A2(n306), .A3(n[157]), .A4(n[156]), .Z(n305) );
  XOR4D0 U296 ( .A1(n[150]), .A2(n[149]), .A3(n307), .A4(n308), .Z(n306) );
  XOR3D0 U297 ( .A1(n309), .A2(n310), .A3(n[148]), .Z(n308) );
  XOR4D0 U298 ( .A1(n[141]), .A2(n311), .A3(n[143]), .A4(n[142]), .Z(n310) );
  XOR4D0 U299 ( .A1(n[136]), .A2(n[135]), .A3(n312), .A4(n313), .Z(n311) );
  XOR3D0 U300 ( .A1(n314), .A2(n315), .A3(n[134]), .Z(n313) );
  XOR3D0 U301 ( .A1(n[129]), .A2(n[128]), .A3(n316), .Z(n315) );
  XOR3D0 U302 ( .A1(n317), .A2(n318), .A3(n[127]), .Z(n316) );
  XOR4D0 U303 ( .A1(n[120]), .A2(n[119]), .A3(n[122]), .A4(n[121]), .Z(n318)
         );
  XOR4D0 U304 ( .A1(n[124]), .A2(n[123]), .A3(n[126]), .A4(n[125]), .Z(n317)
         );
  XOR4D0 U305 ( .A1(n[131]), .A2(n[130]), .A3(n[133]), .A4(n[132]), .Z(n314)
         );
  XOR4D0 U306 ( .A1(n[138]), .A2(n[137]), .A3(n[140]), .A4(n[139]), .Z(n312)
         );
  XOR4D0 U307 ( .A1(n[145]), .A2(n[144]), .A3(n[147]), .A4(n[146]), .Z(n309)
         );
  XOR4D0 U308 ( .A1(n[152]), .A2(n[151]), .A3(n[154]), .A4(n[153]), .Z(n307)
         );
  XOR4D0 U309 ( .A1(n[159]), .A2(n[158]), .A3(n[161]), .A4(n[160]), .Z(n304)
         );
  XOR4D0 U310 ( .A1(n[166]), .A2(n[165]), .A3(n[168]), .A4(n[167]), .Z(n302)
         );
  XOR4D0 U311 ( .A1(n[173]), .A2(n[172]), .A3(n[175]), .A4(n[174]), .Z(n299)
         );
  XOR4D0 U312 ( .A1(n[180]), .A2(n[179]), .A3(n[182]), .A4(n[181]), .Z(n297)
         );
  XOR4D0 U313 ( .A1(n[187]), .A2(n[186]), .A3(n[189]), .A4(n[188]), .Z(n294)
         );
  XOR4D0 U314 ( .A1(n[194]), .A2(n[193]), .A3(n[196]), .A4(n[195]), .Z(n292)
         );
  XOR4D0 U315 ( .A1(n[201]), .A2(n[200]), .A3(n[203]), .A4(n[202]), .Z(n289)
         );
  XOR4D0 U316 ( .A1(n[208]), .A2(n[207]), .A3(n[210]), .A4(n[209]), .Z(n287)
         );
  XOR4D0 U317 ( .A1(n[215]), .A2(n[214]), .A3(n[217]), .A4(n[216]), .Z(n284)
         );
  XOR4D0 U318 ( .A1(n[222]), .A2(n[221]), .A3(n[224]), .A4(n[223]), .Z(n282)
         );
  XOR4D0 U319 ( .A1(n[229]), .A2(n[228]), .A3(n[231]), .A4(n[230]), .Z(n279)
         );
  XOR4D0 U320 ( .A1(n[236]), .A2(n[235]), .A3(n[238]), .A4(n[237]), .Z(n277)
         );
  XOR4D0 U321 ( .A1(n[243]), .A2(n[242]), .A3(n[245]), .A4(n[244]), .Z(n274)
         );
  XOR3D0 U322 ( .A1(n319), .A2(n320), .A3(n[118]), .Z(s[5]) );
  XOR4D0 U323 ( .A1(a[5]), .A2(n321), .A3(n[113]), .A4(b[5]), .Z(n320) );
  XOR4D0 U324 ( .A1(n[108]), .A2(n[107]), .A3(n322), .A4(n323), .Z(n321) );
  XOR3D0 U325 ( .A1(n324), .A2(n325), .A3(n[106]), .Z(n323) );
  XOR4D0 U326 ( .A1(n[100]), .A2(n326), .A3(n[102]), .A4(n[101]), .Z(n325) );
  XOR4D0 U327 ( .A1(n[94]), .A2(n[93]), .A3(n327), .A4(n328), .Z(n326) );
  XOR3D0 U328 ( .A1(n329), .A2(n330), .A3(n[92]), .Z(n328) );
  XOR4D0 U329 ( .A1(n[85]), .A2(n331), .A3(n[87]), .A4(n[86]), .Z(n330) );
  XOR4D0 U330 ( .A1(n[80]), .A2(n[79]), .A3(n332), .A4(n333), .Z(n331) );
  XOR3D0 U331 ( .A1(n334), .A2(n335), .A3(n[78]), .Z(n333) );
  XOR4D0 U332 ( .A1(n[71]), .A2(n336), .A3(n[73]), .A4(n[72]), .Z(n335) );
  XOR4D0 U333 ( .A1(n[66]), .A2(n[65]), .A3(n337), .A4(n338), .Z(n336) );
  XOR3D0 U334 ( .A1(n339), .A2(n340), .A3(n[64]), .Z(n338) );
  XOR4D0 U335 ( .A1(n[57]), .A2(n[56]), .A3(n[59]), .A4(n[58]), .Z(n340) );
  XOR4D0 U336 ( .A1(n[61]), .A2(n[60]), .A3(n[63]), .A4(n[62]), .Z(n339) );
  XOR4D0 U337 ( .A1(n[68]), .A2(n[67]), .A3(n[70]), .A4(n[69]), .Z(n337) );
  XOR4D0 U338 ( .A1(n[75]), .A2(n[74]), .A3(n[77]), .A4(n[76]), .Z(n334) );
  XOR4D0 U339 ( .A1(n[82]), .A2(n[81]), .A3(n[84]), .A4(n[83]), .Z(n332) );
  XOR4D0 U340 ( .A1(n[89]), .A2(n[88]), .A3(n[91]), .A4(n[90]), .Z(n329) );
  XOR4D0 U341 ( .A1(n[96]), .A2(n[95]), .A3(n[98]), .A4(n[97]), .Z(n327) );
  XOR4D0 U342 ( .A1(n[104]), .A2(n[103]), .A3(n[99]), .A4(n[105]), .Z(n324) );
  XOR4D0 U343 ( .A1(n[110]), .A2(n[109]), .A3(n[112]), .A4(n[111]), .Z(n322)
         );
  XOR4D0 U344 ( .A1(n[115]), .A2(n[114]), .A3(n[117]), .A4(n[116]), .Z(n319)
         );
  XOR4D0 U345 ( .A1(n341), .A2(n342), .A3(n343), .A4(n[50]), .Z(s[4]) );
  XOR3D0 U346 ( .A1(n[53]), .A2(n[52]), .A3(n[51]), .Z(n343) );
  XOR4D0 U347 ( .A1(a[4]), .A2(n344), .A3(n[47]), .A4(b[4]), .Z(n342) );
  XOR4D0 U348 ( .A1(n[42]), .A2(n[41]), .A3(n345), .A4(n346), .Z(n344) );
  XOR3D0 U349 ( .A1(n347), .A2(n348), .A3(n[40]), .Z(n346) );
  XOR3D0 U350 ( .A1(n[35]), .A2(n[34]), .A3(n349), .Z(n348) );
  XOR3D0 U351 ( .A1(n350), .A2(n351), .A3(n[33]), .Z(n349) );
  XOR4D0 U352 ( .A1(n[26]), .A2(n[25]), .A3(n[28]), .A4(n[27]), .Z(n351) );
  XOR4D0 U353 ( .A1(n[30]), .A2(n[29]), .A3(n[32]), .A4(n[31]), .Z(n350) );
  XOR4D0 U354 ( .A1(n[37]), .A2(n[36]), .A3(n[39]), .A4(n[38]), .Z(n347) );
  XOR4D0 U355 ( .A1(n[44]), .A2(n[43]), .A3(n[46]), .A4(n[45]), .Z(n345) );
  XOR4D0 U356 ( .A1(n[49]), .A2(n[48]), .A3(n[55]), .A4(n[54]), .Z(n341) );
  XOR4D0 U357 ( .A1(b[3]), .A2(a[3]), .A3(n352), .A4(n353), .Z(s[3]) );
  XOR3D0 U358 ( .A1(n[20]), .A2(n[19]), .A3(n354), .Z(n353) );
  XOR3D0 U359 ( .A1(n355), .A2(n356), .A3(n[18]), .Z(n354) );
  XOR4D0 U360 ( .A1(n[11]), .A2(n[10]), .A3(n[13]), .A4(n[12]), .Z(n356) );
  XOR4D0 U361 ( .A1(n[15]), .A2(n[14]), .A3(n[17]), .A4(n[16]), .Z(n355) );
  XOR4D0 U362 ( .A1(n[22]), .A2(n[21]), .A3(n[24]), .A4(n[23]), .Z(n352) );
  XOR3D0 U363 ( .A1(n357), .A2(n358), .A3(n[9]), .Z(s[2]) );
  XOR4D0 U364 ( .A1(b[2]), .A2(a[2]), .A3(n[4]), .A4(n[3]), .Z(n358) );
  XOR4D0 U365 ( .A1(n[6]), .A2(n[5]), .A3(n[8]), .A4(n[7]), .Z(n357) );
  XOR3D0 U366 ( .A1(b[1]), .A2(a[1]), .A3(n359), .Z(s[1]) );
  XOR3D0 U367 ( .A1(n[2]), .A2(n[1]), .A3(n[0]), .Z(n359) );
  XOR2D0 U368 ( .A1(b[0]), .A2(a[0]), .Z(s[0]) );
endmodule


module gen_nonlinear_part ( a, b, n );
  input [8:0] a;
  input [8:0] b;
  output [1011:0] n;


  INVD0 U2 ( .I(1'b1), .ZN(n[1]) );
  INVD0 U4 ( .I(1'b1), .ZN(n[2]) );
  INVD0 U6 ( .I(1'b1), .ZN(n[5]) );
  INVD0 U8 ( .I(1'b1), .ZN(n[6]) );
  INVD0 U10 ( .I(1'b1), .ZN(n[8]) );
  INVD0 U12 ( .I(1'b1), .ZN(n[9]) );
  INVD0 U14 ( .I(1'b1), .ZN(n[13]) );
  INVD0 U16 ( .I(1'b1), .ZN(n[14]) );
  INVD0 U18 ( .I(1'b1), .ZN(n[16]) );
  INVD0 U20 ( .I(1'b1), .ZN(n[17]) );
  INVD0 U22 ( .I(1'b1), .ZN(n[20]) );
  INVD0 U24 ( .I(1'b1), .ZN(n[21]) );
  INVD0 U26 ( .I(1'b1), .ZN(n[23]) );
  INVD0 U28 ( .I(1'b1), .ZN(n[24]) );
  INVD0 U30 ( .I(1'b1), .ZN(n[29]) );
  INVD0 U32 ( .I(1'b1), .ZN(n[30]) );
  INVD0 U34 ( .I(1'b1), .ZN(n[32]) );
  INVD0 U36 ( .I(1'b1), .ZN(n[33]) );
  INVD0 U38 ( .I(1'b1), .ZN(n[36]) );
  INVD0 U40 ( .I(1'b1), .ZN(n[37]) );
  INVD0 U42 ( .I(1'b1), .ZN(n[39]) );
  INVD0 U44 ( .I(1'b1), .ZN(n[40]) );
  INVD0 U46 ( .I(1'b1), .ZN(n[44]) );
  INVD0 U48 ( .I(1'b1), .ZN(n[45]) );
  INVD0 U50 ( .I(1'b1), .ZN(n[47]) );
  INVD0 U52 ( .I(1'b1), .ZN(n[48]) );
  INVD0 U54 ( .I(1'b1), .ZN(n[51]) );
  INVD0 U56 ( .I(1'b1), .ZN(n[52]) );
  INVD0 U58 ( .I(1'b1), .ZN(n[54]) );
  INVD0 U60 ( .I(1'b1), .ZN(n[55]) );
  INVD0 U62 ( .I(1'b1), .ZN(n[61]) );
  INVD0 U64 ( .I(1'b1), .ZN(n[62]) );
  INVD0 U66 ( .I(1'b1), .ZN(n[64]) );
  INVD0 U68 ( .I(1'b1), .ZN(n[65]) );
  INVD0 U70 ( .I(1'b1), .ZN(n[68]) );
  INVD0 U72 ( .I(1'b1), .ZN(n[69]) );
  INVD0 U74 ( .I(1'b1), .ZN(n[71]) );
  INVD0 U76 ( .I(1'b1), .ZN(n[72]) );
  INVD0 U78 ( .I(1'b1), .ZN(n[76]) );
  INVD0 U80 ( .I(1'b1), .ZN(n[77]) );
  INVD0 U82 ( .I(1'b1), .ZN(n[79]) );
  INVD0 U84 ( .I(1'b1), .ZN(n[80]) );
  INVD0 U86 ( .I(1'b1), .ZN(n[83]) );
  INVD0 U88 ( .I(1'b1), .ZN(n[84]) );
  INVD0 U90 ( .I(1'b1), .ZN(n[86]) );
  INVD0 U92 ( .I(1'b1), .ZN(n[87]) );
  INVD0 U94 ( .I(1'b1), .ZN(n[92]) );
  INVD0 U96 ( .I(1'b1), .ZN(n[93]) );
  INVD0 U98 ( .I(1'b1), .ZN(n[95]) );
  INVD0 U100 ( .I(1'b1), .ZN(n[96]) );
  INVD0 U102 ( .I(1'b1), .ZN(n[99]) );
  INVD0 U104 ( .I(1'b1), .ZN(n[100]) );
  INVD0 U106 ( .I(1'b1), .ZN(n[102]) );
  INVD0 U108 ( .I(1'b1), .ZN(n[103]) );
  INVD0 U110 ( .I(1'b1), .ZN(n[107]) );
  INVD0 U112 ( .I(1'b1), .ZN(n[108]) );
  INVD0 U114 ( .I(1'b1), .ZN(n[110]) );
  INVD0 U116 ( .I(1'b1), .ZN(n[111]) );
  INVD0 U118 ( .I(1'b1), .ZN(n[114]) );
  INVD0 U120 ( .I(1'b1), .ZN(n[115]) );
  INVD0 U122 ( .I(1'b1), .ZN(n[117]) );
  INVD0 U124 ( .I(1'b1), .ZN(n[118]) );
  INVD0 U126 ( .I(1'b1), .ZN(n[125]) );
  INVD0 U128 ( .I(1'b1), .ZN(n[126]) );
  INVD0 U130 ( .I(1'b1), .ZN(n[128]) );
  INVD0 U132 ( .I(1'b1), .ZN(n[129]) );
  INVD0 U134 ( .I(1'b1), .ZN(n[132]) );
  INVD0 U136 ( .I(1'b1), .ZN(n[133]) );
  INVD0 U138 ( .I(1'b1), .ZN(n[135]) );
  INVD0 U140 ( .I(1'b1), .ZN(n[136]) );
  INVD0 U142 ( .I(1'b1), .ZN(n[140]) );
  INVD0 U144 ( .I(1'b1), .ZN(n[141]) );
  INVD0 U146 ( .I(1'b1), .ZN(n[143]) );
  INVD0 U148 ( .I(1'b1), .ZN(n[144]) );
  INVD0 U150 ( .I(1'b1), .ZN(n[147]) );
  INVD0 U152 ( .I(1'b1), .ZN(n[148]) );
  INVD0 U154 ( .I(1'b1), .ZN(n[150]) );
  INVD0 U156 ( .I(1'b1), .ZN(n[151]) );
  INVD0 U158 ( .I(1'b1), .ZN(n[156]) );
  INVD0 U160 ( .I(1'b1), .ZN(n[157]) );
  INVD0 U162 ( .I(1'b1), .ZN(n[159]) );
  INVD0 U164 ( .I(1'b1), .ZN(n[160]) );
  INVD0 U166 ( .I(1'b1), .ZN(n[163]) );
  INVD0 U168 ( .I(1'b1), .ZN(n[164]) );
  INVD0 U170 ( .I(1'b1), .ZN(n[166]) );
  INVD0 U172 ( .I(1'b1), .ZN(n[167]) );
  INVD0 U174 ( .I(1'b1), .ZN(n[171]) );
  INVD0 U176 ( .I(1'b1), .ZN(n[172]) );
  INVD0 U178 ( .I(1'b1), .ZN(n[174]) );
  INVD0 U180 ( .I(1'b1), .ZN(n[175]) );
  INVD0 U182 ( .I(1'b1), .ZN(n[178]) );
  INVD0 U184 ( .I(1'b1), .ZN(n[179]) );
  INVD0 U186 ( .I(1'b1), .ZN(n[181]) );
  INVD0 U188 ( .I(1'b1), .ZN(n[182]) );
  INVD0 U190 ( .I(1'b1), .ZN(n[188]) );
  INVD0 U192 ( .I(1'b1), .ZN(n[189]) );
  INVD0 U194 ( .I(1'b1), .ZN(n[191]) );
  INVD0 U196 ( .I(1'b1), .ZN(n[192]) );
  INVD0 U198 ( .I(1'b1), .ZN(n[195]) );
  INVD0 U200 ( .I(1'b1), .ZN(n[196]) );
  INVD0 U202 ( .I(1'b1), .ZN(n[198]) );
  INVD0 U204 ( .I(1'b1), .ZN(n[199]) );
  INVD0 U206 ( .I(1'b1), .ZN(n[203]) );
  INVD0 U208 ( .I(1'b1), .ZN(n[204]) );
  INVD0 U210 ( .I(1'b1), .ZN(n[206]) );
  INVD0 U212 ( .I(1'b1), .ZN(n[207]) );
  INVD0 U214 ( .I(1'b1), .ZN(n[210]) );
  INVD0 U216 ( .I(1'b1), .ZN(n[211]) );
  INVD0 U218 ( .I(1'b1), .ZN(n[213]) );
  INVD0 U220 ( .I(1'b1), .ZN(n[214]) );
  INVD0 U222 ( .I(1'b1), .ZN(n[219]) );
  INVD0 U224 ( .I(1'b1), .ZN(n[220]) );
  INVD0 U226 ( .I(1'b1), .ZN(n[222]) );
  INVD0 U228 ( .I(1'b1), .ZN(n[223]) );
  INVD0 U230 ( .I(1'b1), .ZN(n[226]) );
  INVD0 U232 ( .I(1'b1), .ZN(n[227]) );
  INVD0 U234 ( .I(1'b1), .ZN(n[229]) );
  INVD0 U236 ( .I(1'b1), .ZN(n[230]) );
  INVD0 U238 ( .I(1'b1), .ZN(n[234]) );
  INVD0 U240 ( .I(1'b1), .ZN(n[235]) );
  INVD0 U242 ( .I(1'b1), .ZN(n[237]) );
  INVD0 U244 ( .I(1'b1), .ZN(n[238]) );
  INVD0 U246 ( .I(1'b1), .ZN(n[241]) );
  INVD0 U248 ( .I(1'b1), .ZN(n[242]) );
  INVD0 U250 ( .I(1'b1), .ZN(n[244]) );
  INVD0 U252 ( .I(1'b1), .ZN(n[245]) );
  INVD0 U254 ( .I(1'b1), .ZN(n[253]) );
  INVD0 U256 ( .I(1'b1), .ZN(n[254]) );
  INVD0 U258 ( .I(1'b1), .ZN(n[256]) );
  INVD0 U260 ( .I(1'b1), .ZN(n[257]) );
  INVD0 U262 ( .I(1'b1), .ZN(n[260]) );
  INVD0 U264 ( .I(1'b1), .ZN(n[261]) );
  INVD0 U266 ( .I(1'b1), .ZN(n[263]) );
  INVD0 U268 ( .I(1'b1), .ZN(n[264]) );
  INVD0 U270 ( .I(1'b1), .ZN(n[268]) );
  INVD0 U272 ( .I(1'b1), .ZN(n[269]) );
  INVD0 U274 ( .I(1'b1), .ZN(n[271]) );
  INVD0 U276 ( .I(1'b1), .ZN(n[272]) );
  INVD0 U278 ( .I(1'b1), .ZN(n[275]) );
  INVD0 U280 ( .I(1'b1), .ZN(n[276]) );
  INVD0 U282 ( .I(1'b1), .ZN(n[278]) );
  INVD0 U284 ( .I(1'b1), .ZN(n[279]) );
  INVD0 U286 ( .I(1'b1), .ZN(n[284]) );
  INVD0 U288 ( .I(1'b1), .ZN(n[285]) );
  INVD0 U290 ( .I(1'b1), .ZN(n[287]) );
  INVD0 U292 ( .I(1'b1), .ZN(n[288]) );
  INVD0 U294 ( .I(1'b1), .ZN(n[291]) );
  INVD0 U296 ( .I(1'b1), .ZN(n[292]) );
  INVD0 U298 ( .I(1'b1), .ZN(n[294]) );
  INVD0 U300 ( .I(1'b1), .ZN(n[295]) );
  INVD0 U302 ( .I(1'b1), .ZN(n[299]) );
  INVD0 U304 ( .I(1'b1), .ZN(n[300]) );
  INVD0 U306 ( .I(1'b1), .ZN(n[302]) );
  INVD0 U308 ( .I(1'b1), .ZN(n[303]) );
  INVD0 U310 ( .I(1'b1), .ZN(n[306]) );
  INVD0 U312 ( .I(1'b1), .ZN(n[307]) );
  INVD0 U314 ( .I(1'b1), .ZN(n[309]) );
  INVD0 U316 ( .I(1'b1), .ZN(n[310]) );
  INVD0 U318 ( .I(1'b1), .ZN(n[316]) );
  INVD0 U320 ( .I(1'b1), .ZN(n[317]) );
  INVD0 U322 ( .I(1'b1), .ZN(n[319]) );
  INVD0 U324 ( .I(1'b1), .ZN(n[320]) );
  INVD0 U326 ( .I(1'b1), .ZN(n[323]) );
  INVD0 U328 ( .I(1'b1), .ZN(n[324]) );
  INVD0 U330 ( .I(1'b1), .ZN(n[326]) );
  INVD0 U332 ( .I(1'b1), .ZN(n[327]) );
  INVD0 U334 ( .I(1'b1), .ZN(n[331]) );
  INVD0 U336 ( .I(1'b1), .ZN(n[332]) );
  INVD0 U338 ( .I(1'b1), .ZN(n[334]) );
  INVD0 U340 ( .I(1'b1), .ZN(n[335]) );
  INVD0 U342 ( .I(1'b1), .ZN(n[338]) );
  INVD0 U344 ( .I(1'b1), .ZN(n[339]) );
  INVD0 U346 ( .I(1'b1), .ZN(n[341]) );
  INVD0 U348 ( .I(1'b1), .ZN(n[342]) );
  INVD0 U350 ( .I(1'b1), .ZN(n[347]) );
  INVD0 U352 ( .I(1'b1), .ZN(n[348]) );
  INVD0 U354 ( .I(1'b1), .ZN(n[350]) );
  INVD0 U356 ( .I(1'b1), .ZN(n[351]) );
  INVD0 U358 ( .I(1'b1), .ZN(n[354]) );
  INVD0 U360 ( .I(1'b1), .ZN(n[355]) );
  INVD0 U362 ( .I(1'b1), .ZN(n[357]) );
  INVD0 U364 ( .I(1'b1), .ZN(n[358]) );
  INVD0 U366 ( .I(1'b1), .ZN(n[362]) );
  INVD0 U368 ( .I(1'b1), .ZN(n[363]) );
  INVD0 U370 ( .I(1'b1), .ZN(n[365]) );
  INVD0 U372 ( .I(1'b1), .ZN(n[366]) );
  INVD0 U374 ( .I(1'b1), .ZN(n[369]) );
  INVD0 U376 ( .I(1'b1), .ZN(n[370]) );
  INVD0 U378 ( .I(1'b1), .ZN(n[372]) );
  INVD0 U380 ( .I(1'b1), .ZN(n[373]) );
  INVD0 U382 ( .I(1'b1), .ZN(n[380]) );
  INVD0 U384 ( .I(1'b1), .ZN(n[381]) );
  INVD0 U386 ( .I(1'b1), .ZN(n[383]) );
  INVD0 U388 ( .I(1'b1), .ZN(n[384]) );
  INVD0 U390 ( .I(1'b1), .ZN(n[387]) );
  INVD0 U392 ( .I(1'b1), .ZN(n[388]) );
  INVD0 U394 ( .I(1'b1), .ZN(n[390]) );
  INVD0 U396 ( .I(1'b1), .ZN(n[391]) );
  INVD0 U398 ( .I(1'b1), .ZN(n[395]) );
  INVD0 U400 ( .I(1'b1), .ZN(n[396]) );
  INVD0 U402 ( .I(1'b1), .ZN(n[398]) );
  INVD0 U404 ( .I(1'b1), .ZN(n[399]) );
  INVD0 U406 ( .I(1'b1), .ZN(n[402]) );
  INVD0 U408 ( .I(1'b1), .ZN(n[403]) );
  INVD0 U410 ( .I(1'b1), .ZN(n[405]) );
  INVD0 U412 ( .I(1'b1), .ZN(n[406]) );
  INVD0 U414 ( .I(1'b1), .ZN(n[411]) );
  INVD0 U416 ( .I(1'b1), .ZN(n[412]) );
  INVD0 U418 ( .I(1'b1), .ZN(n[414]) );
  INVD0 U420 ( .I(1'b1), .ZN(n[415]) );
  INVD0 U422 ( .I(1'b1), .ZN(n[418]) );
  INVD0 U424 ( .I(1'b1), .ZN(n[419]) );
  INVD0 U426 ( .I(1'b1), .ZN(n[421]) );
  INVD0 U428 ( .I(1'b1), .ZN(n[422]) );
  INVD0 U430 ( .I(1'b1), .ZN(n[426]) );
  INVD0 U432 ( .I(1'b1), .ZN(n[427]) );
  INVD0 U434 ( .I(1'b1), .ZN(n[429]) );
  INVD0 U436 ( .I(1'b1), .ZN(n[430]) );
  INVD0 U438 ( .I(1'b1), .ZN(n[433]) );
  INVD0 U440 ( .I(1'b1), .ZN(n[434]) );
  INVD0 U442 ( .I(1'b1), .ZN(n[436]) );
  INVD0 U444 ( .I(1'b1), .ZN(n[437]) );
  INVD0 U446 ( .I(1'b1), .ZN(n[443]) );
  INVD0 U448 ( .I(1'b1), .ZN(n[444]) );
  INVD0 U450 ( .I(1'b1), .ZN(n[446]) );
  INVD0 U452 ( .I(1'b1), .ZN(n[447]) );
  INVD0 U454 ( .I(1'b1), .ZN(n[450]) );
  INVD0 U456 ( .I(1'b1), .ZN(n[451]) );
  INVD0 U458 ( .I(1'b1), .ZN(n[453]) );
  INVD0 U460 ( .I(1'b1), .ZN(n[454]) );
  INVD0 U462 ( .I(1'b1), .ZN(n[458]) );
  INVD0 U464 ( .I(1'b1), .ZN(n[459]) );
  INVD0 U466 ( .I(1'b1), .ZN(n[461]) );
  INVD0 U468 ( .I(1'b1), .ZN(n[462]) );
  INVD0 U470 ( .I(1'b1), .ZN(n[465]) );
  INVD0 U472 ( .I(1'b1), .ZN(n[466]) );
  INVD0 U474 ( .I(1'b1), .ZN(n[468]) );
  INVD0 U476 ( .I(1'b1), .ZN(n[469]) );
  INVD0 U478 ( .I(1'b1), .ZN(n[474]) );
  INVD0 U480 ( .I(1'b1), .ZN(n[475]) );
  INVD0 U482 ( .I(1'b1), .ZN(n[477]) );
  INVD0 U484 ( .I(1'b1), .ZN(n[478]) );
  INVD0 U486 ( .I(1'b1), .ZN(n[481]) );
  INVD0 U488 ( .I(1'b1), .ZN(n[482]) );
  INVD0 U490 ( .I(1'b1), .ZN(n[484]) );
  INVD0 U492 ( .I(1'b1), .ZN(n[485]) );
  INVD0 U494 ( .I(1'b1), .ZN(n[489]) );
  INVD0 U496 ( .I(1'b1), .ZN(n[490]) );
  INVD0 U498 ( .I(1'b1), .ZN(n[492]) );
  INVD0 U500 ( .I(1'b1), .ZN(n[493]) );
  INVD0 U502 ( .I(1'b1), .ZN(n[496]) );
  INVD0 U505 ( .I(1'b1), .ZN(n[497]) );
  INVD0 U507 ( .I(1'b1), .ZN(n[499]) );
  INVD0 U509 ( .I(1'b1), .ZN(n[500]) );
  INVD0 U511 ( .I(1'b1), .ZN(n[509]) );
  INVD0 U513 ( .I(1'b1), .ZN(n[510]) );
  INVD0 U515 ( .I(1'b1), .ZN(n[512]) );
  INVD0 U517 ( .I(1'b1), .ZN(n[513]) );
  INVD0 U519 ( .I(1'b1), .ZN(n[516]) );
  INVD0 U521 ( .I(1'b1), .ZN(n[517]) );
  INVD0 U523 ( .I(1'b1), .ZN(n[519]) );
  INVD0 U525 ( .I(1'b1), .ZN(n[520]) );
  INVD0 U527 ( .I(1'b1), .ZN(n[524]) );
  INVD0 U529 ( .I(1'b1), .ZN(n[525]) );
  INVD0 U531 ( .I(1'b1), .ZN(n[527]) );
  INVD0 U533 ( .I(1'b1), .ZN(n[528]) );
  INVD0 U535 ( .I(1'b1), .ZN(n[531]) );
  INVD0 U537 ( .I(1'b1), .ZN(n[532]) );
  INVD0 U539 ( .I(1'b1), .ZN(n[534]) );
  INVD0 U541 ( .I(1'b1), .ZN(n[535]) );
  INVD0 U543 ( .I(1'b1), .ZN(n[540]) );
  INVD0 U545 ( .I(1'b1), .ZN(n[541]) );
  INVD0 U547 ( .I(1'b1), .ZN(n[543]) );
  INVD0 U549 ( .I(1'b1), .ZN(n[544]) );
  INVD0 U551 ( .I(1'b1), .ZN(n[547]) );
  INVD0 U553 ( .I(1'b1), .ZN(n[548]) );
  INVD0 U555 ( .I(1'b1), .ZN(n[550]) );
  INVD0 U557 ( .I(1'b1), .ZN(n[551]) );
  INVD0 U559 ( .I(1'b1), .ZN(n[555]) );
  INVD0 U561 ( .I(1'b1), .ZN(n[556]) );
  INVD0 U563 ( .I(1'b1), .ZN(n[558]) );
  INVD0 U565 ( .I(1'b1), .ZN(n[559]) );
  INVD0 U567 ( .I(1'b1), .ZN(n[562]) );
  INVD0 U569 ( .I(1'b1), .ZN(n[563]) );
  INVD0 U571 ( .I(1'b1), .ZN(n[565]) );
  INVD0 U573 ( .I(1'b1), .ZN(n[566]) );
  INVD0 U575 ( .I(1'b1), .ZN(n[572]) );
  INVD0 U577 ( .I(1'b1), .ZN(n[573]) );
  INVD0 U579 ( .I(1'b1), .ZN(n[575]) );
  INVD0 U581 ( .I(1'b1), .ZN(n[576]) );
  INVD0 U583 ( .I(1'b1), .ZN(n[579]) );
  INVD0 U585 ( .I(1'b1), .ZN(n[580]) );
  INVD0 U587 ( .I(1'b1), .ZN(n[582]) );
  INVD0 U589 ( .I(1'b1), .ZN(n[583]) );
  INVD0 U591 ( .I(1'b1), .ZN(n[587]) );
  INVD0 U593 ( .I(1'b1), .ZN(n[588]) );
  INVD0 U595 ( .I(1'b1), .ZN(n[590]) );
  INVD0 U597 ( .I(1'b1), .ZN(n[591]) );
  INVD0 U599 ( .I(1'b1), .ZN(n[594]) );
  INVD0 U601 ( .I(1'b1), .ZN(n[595]) );
  INVD0 U603 ( .I(1'b1), .ZN(n[597]) );
  INVD0 U605 ( .I(1'b1), .ZN(n[598]) );
  INVD0 U607 ( .I(1'b1), .ZN(n[603]) );
  INVD0 U609 ( .I(1'b1), .ZN(n[604]) );
  INVD0 U611 ( .I(1'b1), .ZN(n[606]) );
  INVD0 U613 ( .I(1'b1), .ZN(n[607]) );
  INVD0 U615 ( .I(1'b1), .ZN(n[610]) );
  INVD0 U617 ( .I(1'b1), .ZN(n[611]) );
  INVD0 U619 ( .I(1'b1), .ZN(n[613]) );
  INVD0 U621 ( .I(1'b1), .ZN(n[614]) );
  INVD0 U623 ( .I(1'b1), .ZN(n[618]) );
  INVD0 U625 ( .I(1'b1), .ZN(n[619]) );
  INVD0 U627 ( .I(1'b1), .ZN(n[621]) );
  INVD0 U629 ( .I(1'b1), .ZN(n[622]) );
  INVD0 U631 ( .I(1'b1), .ZN(n[625]) );
  INVD0 U633 ( .I(1'b1), .ZN(n[626]) );
  INVD0 U635 ( .I(1'b1), .ZN(n[628]) );
  INVD0 U637 ( .I(1'b1), .ZN(n[629]) );
  INVD0 U639 ( .I(1'b1), .ZN(n[636]) );
  INVD0 U641 ( .I(1'b1), .ZN(n[637]) );
  INVD0 U643 ( .I(1'b1), .ZN(n[639]) );
  INVD0 U645 ( .I(1'b1), .ZN(n[640]) );
  INVD0 U647 ( .I(1'b1), .ZN(n[643]) );
  INVD0 U649 ( .I(1'b1), .ZN(n[644]) );
  INVD0 U651 ( .I(1'b1), .ZN(n[646]) );
  INVD0 U653 ( .I(1'b1), .ZN(n[647]) );
  INVD0 U655 ( .I(1'b1), .ZN(n[651]) );
  INVD0 U657 ( .I(1'b1), .ZN(n[652]) );
  INVD0 U659 ( .I(1'b1), .ZN(n[654]) );
  INVD0 U661 ( .I(1'b1), .ZN(n[655]) );
  INVD0 U663 ( .I(1'b1), .ZN(n[658]) );
  INVD0 U665 ( .I(1'b1), .ZN(n[659]) );
  INVD0 U667 ( .I(1'b1), .ZN(n[661]) );
  INVD0 U669 ( .I(1'b1), .ZN(n[662]) );
  INVD0 U671 ( .I(1'b1), .ZN(n[667]) );
  INVD0 U673 ( .I(1'b1), .ZN(n[668]) );
  INVD0 U675 ( .I(1'b1), .ZN(n[670]) );
  INVD0 U677 ( .I(1'b1), .ZN(n[671]) );
  INVD0 U679 ( .I(1'b1), .ZN(n[674]) );
  INVD0 U681 ( .I(1'b1), .ZN(n[675]) );
  INVD0 U683 ( .I(1'b1), .ZN(n[677]) );
  INVD0 U685 ( .I(1'b1), .ZN(n[678]) );
  INVD0 U687 ( .I(1'b1), .ZN(n[682]) );
  INVD0 U689 ( .I(1'b1), .ZN(n[683]) );
  INVD0 U691 ( .I(1'b1), .ZN(n[685]) );
  INVD0 U693 ( .I(1'b1), .ZN(n[686]) );
  INVD0 U695 ( .I(1'b1), .ZN(n[689]) );
  INVD0 U697 ( .I(1'b1), .ZN(n[690]) );
  INVD0 U699 ( .I(1'b1), .ZN(n[692]) );
  INVD0 U701 ( .I(1'b1), .ZN(n[693]) );
  INVD0 U703 ( .I(1'b1), .ZN(n[699]) );
  INVD0 U705 ( .I(1'b1), .ZN(n[700]) );
  INVD0 U707 ( .I(1'b1), .ZN(n[702]) );
  INVD0 U709 ( .I(1'b1), .ZN(n[703]) );
  INVD0 U711 ( .I(1'b1), .ZN(n[706]) );
  INVD0 U713 ( .I(1'b1), .ZN(n[707]) );
  INVD0 U715 ( .I(1'b1), .ZN(n[709]) );
  INVD0 U717 ( .I(1'b1), .ZN(n[710]) );
  INVD0 U719 ( .I(1'b1), .ZN(n[714]) );
  INVD0 U721 ( .I(1'b1), .ZN(n[715]) );
  INVD0 U723 ( .I(1'b1), .ZN(n[717]) );
  INVD0 U725 ( .I(1'b1), .ZN(n[718]) );
  INVD0 U727 ( .I(1'b1), .ZN(n[721]) );
  INVD0 U729 ( .I(1'b1), .ZN(n[722]) );
  INVD0 U731 ( .I(1'b1), .ZN(n[724]) );
  INVD0 U733 ( .I(1'b1), .ZN(n[725]) );
  INVD0 U735 ( .I(1'b1), .ZN(n[730]) );
  INVD0 U737 ( .I(1'b1), .ZN(n[731]) );
  INVD0 U739 ( .I(1'b1), .ZN(n[733]) );
  INVD0 U741 ( .I(1'b1), .ZN(n[734]) );
  INVD0 U743 ( .I(1'b1), .ZN(n[737]) );
  INVD0 U745 ( .I(1'b1), .ZN(n[738]) );
  INVD0 U747 ( .I(1'b1), .ZN(n[740]) );
  INVD0 U749 ( .I(1'b1), .ZN(n[741]) );
  INVD0 U751 ( .I(1'b1), .ZN(n[745]) );
  INVD0 U753 ( .I(1'b1), .ZN(n[746]) );
  INVD0 U755 ( .I(1'b1), .ZN(n[748]) );
  INVD0 U757 ( .I(1'b1), .ZN(n[749]) );
  INVD0 U759 ( .I(1'b1), .ZN(n[752]) );
  INVD0 U761 ( .I(1'b1), .ZN(n[753]) );
  INVD0 U763 ( .I(1'b1), .ZN(n[755]) );
  INVD0 U765 ( .I(1'b1), .ZN(n[756]) );
  INVD0 U767 ( .I(1'b1), .ZN(n[764]) );
  INVD0 U769 ( .I(1'b1), .ZN(n[765]) );
  INVD0 U771 ( .I(1'b1), .ZN(n[767]) );
  INVD0 U773 ( .I(1'b1), .ZN(n[768]) );
  INVD0 U775 ( .I(1'b1), .ZN(n[771]) );
  INVD0 U777 ( .I(1'b1), .ZN(n[772]) );
  INVD0 U779 ( .I(1'b1), .ZN(n[774]) );
  INVD0 U781 ( .I(1'b1), .ZN(n[775]) );
  INVD0 U783 ( .I(1'b1), .ZN(n[779]) );
  INVD0 U785 ( .I(1'b1), .ZN(n[780]) );
  INVD0 U787 ( .I(1'b1), .ZN(n[782]) );
  INVD0 U789 ( .I(1'b1), .ZN(n[783]) );
  INVD0 U791 ( .I(1'b1), .ZN(n[786]) );
  INVD0 U793 ( .I(1'b1), .ZN(n[787]) );
  INVD0 U795 ( .I(1'b1), .ZN(n[789]) );
  INVD0 U797 ( .I(1'b1), .ZN(n[790]) );
  INVD0 U799 ( .I(1'b1), .ZN(n[795]) );
  INVD0 U801 ( .I(1'b1), .ZN(n[796]) );
  INVD0 U803 ( .I(1'b1), .ZN(n[798]) );
  INVD0 U805 ( .I(1'b1), .ZN(n[799]) );
  INVD0 U807 ( .I(1'b1), .ZN(n[802]) );
  INVD0 U809 ( .I(1'b1), .ZN(n[803]) );
  INVD0 U811 ( .I(1'b1), .ZN(n[805]) );
  INVD0 U813 ( .I(1'b1), .ZN(n[806]) );
  INVD0 U815 ( .I(1'b1), .ZN(n[810]) );
  INVD0 U817 ( .I(1'b1), .ZN(n[811]) );
  INVD0 U819 ( .I(1'b1), .ZN(n[813]) );
  INVD0 U821 ( .I(1'b1), .ZN(n[814]) );
  INVD0 U823 ( .I(1'b1), .ZN(n[817]) );
  INVD0 U825 ( .I(1'b1), .ZN(n[818]) );
  INVD0 U827 ( .I(1'b1), .ZN(n[820]) );
  INVD0 U829 ( .I(1'b1), .ZN(n[821]) );
  INVD0 U831 ( .I(1'b1), .ZN(n[827]) );
  INVD0 U833 ( .I(1'b1), .ZN(n[828]) );
  INVD0 U835 ( .I(1'b1), .ZN(n[830]) );
  INVD0 U837 ( .I(1'b1), .ZN(n[831]) );
  INVD0 U839 ( .I(1'b1), .ZN(n[834]) );
  INVD0 U841 ( .I(1'b1), .ZN(n[835]) );
  INVD0 U843 ( .I(1'b1), .ZN(n[837]) );
  INVD0 U845 ( .I(1'b1), .ZN(n[838]) );
  INVD0 U847 ( .I(1'b1), .ZN(n[842]) );
  INVD0 U849 ( .I(1'b1), .ZN(n[843]) );
  INVD0 U851 ( .I(1'b1), .ZN(n[845]) );
  INVD0 U853 ( .I(1'b1), .ZN(n[846]) );
  INVD0 U855 ( .I(1'b1), .ZN(n[849]) );
  INVD0 U857 ( .I(1'b1), .ZN(n[850]) );
  INVD0 U859 ( .I(1'b1), .ZN(n[852]) );
  INVD0 U861 ( .I(1'b1), .ZN(n[853]) );
  INVD0 U863 ( .I(1'b1), .ZN(n[858]) );
  INVD0 U865 ( .I(1'b1), .ZN(n[859]) );
  INVD0 U867 ( .I(1'b1), .ZN(n[861]) );
  INVD0 U869 ( .I(1'b1), .ZN(n[862]) );
  INVD0 U871 ( .I(1'b1), .ZN(n[865]) );
  INVD0 U873 ( .I(1'b1), .ZN(n[866]) );
  INVD0 U875 ( .I(1'b1), .ZN(n[868]) );
  INVD0 U877 ( .I(1'b1), .ZN(n[869]) );
  INVD0 U879 ( .I(1'b1), .ZN(n[873]) );
  INVD0 U881 ( .I(1'b1), .ZN(n[874]) );
  INVD0 U883 ( .I(1'b1), .ZN(n[876]) );
  INVD0 U885 ( .I(1'b1), .ZN(n[877]) );
  INVD0 U887 ( .I(1'b1), .ZN(n[880]) );
  INVD0 U889 ( .I(1'b1), .ZN(n[881]) );
  INVD0 U891 ( .I(1'b1), .ZN(n[883]) );
  INVD0 U893 ( .I(1'b1), .ZN(n[884]) );
  INVD0 U895 ( .I(1'b1), .ZN(n[891]) );
  INVD0 U897 ( .I(1'b1), .ZN(n[892]) );
  INVD0 U899 ( .I(1'b1), .ZN(n[894]) );
  INVD0 U901 ( .I(1'b1), .ZN(n[895]) );
  INVD0 U903 ( .I(1'b1), .ZN(n[898]) );
  INVD0 U905 ( .I(1'b1), .ZN(n[899]) );
  INVD0 U907 ( .I(1'b1), .ZN(n[901]) );
  INVD0 U909 ( .I(1'b1), .ZN(n[902]) );
  INVD0 U911 ( .I(1'b1), .ZN(n[906]) );
  INVD0 U913 ( .I(1'b1), .ZN(n[907]) );
  INVD0 U915 ( .I(1'b1), .ZN(n[909]) );
  INVD0 U917 ( .I(1'b1), .ZN(n[910]) );
  INVD0 U919 ( .I(1'b1), .ZN(n[913]) );
  INVD0 U921 ( .I(1'b1), .ZN(n[914]) );
  INVD0 U923 ( .I(1'b1), .ZN(n[916]) );
  INVD0 U925 ( .I(1'b1), .ZN(n[917]) );
  INVD0 U927 ( .I(1'b1), .ZN(n[922]) );
  INVD0 U929 ( .I(1'b1), .ZN(n[923]) );
  INVD0 U931 ( .I(1'b1), .ZN(n[925]) );
  INVD0 U933 ( .I(1'b1), .ZN(n[926]) );
  INVD0 U935 ( .I(1'b1), .ZN(n[929]) );
  INVD0 U937 ( .I(1'b1), .ZN(n[930]) );
  INVD0 U939 ( .I(1'b1), .ZN(n[932]) );
  INVD0 U941 ( .I(1'b1), .ZN(n[933]) );
  INVD0 U943 ( .I(1'b1), .ZN(n[937]) );
  INVD0 U945 ( .I(1'b1), .ZN(n[938]) );
  INVD0 U947 ( .I(1'b1), .ZN(n[940]) );
  INVD0 U949 ( .I(1'b1), .ZN(n[941]) );
  INVD0 U951 ( .I(1'b1), .ZN(n[944]) );
  INVD0 U953 ( .I(1'b1), .ZN(n[945]) );
  INVD0 U955 ( .I(1'b1), .ZN(n[947]) );
  INVD0 U957 ( .I(1'b1), .ZN(n[948]) );
  INVD0 U959 ( .I(1'b1), .ZN(n[954]) );
  INVD0 U961 ( .I(1'b1), .ZN(n[955]) );
  INVD0 U963 ( .I(1'b1), .ZN(n[957]) );
  INVD0 U965 ( .I(1'b1), .ZN(n[958]) );
  INVD0 U967 ( .I(1'b1), .ZN(n[961]) );
  INVD0 U969 ( .I(1'b1), .ZN(n[962]) );
  INVD0 U971 ( .I(1'b1), .ZN(n[964]) );
  INVD0 U973 ( .I(1'b1), .ZN(n[965]) );
  INVD0 U975 ( .I(1'b1), .ZN(n[969]) );
  INVD0 U977 ( .I(1'b1), .ZN(n[970]) );
  INVD0 U979 ( .I(1'b1), .ZN(n[972]) );
  INVD0 U981 ( .I(1'b1), .ZN(n[973]) );
  INVD0 U983 ( .I(1'b1), .ZN(n[976]) );
  INVD0 U985 ( .I(1'b1), .ZN(n[977]) );
  INVD0 U987 ( .I(1'b1), .ZN(n[979]) );
  INVD0 U989 ( .I(1'b1), .ZN(n[980]) );
  INVD0 U991 ( .I(1'b1), .ZN(n[985]) );
  INVD0 U993 ( .I(1'b1), .ZN(n[986]) );
  INVD0 U995 ( .I(1'b1), .ZN(n[988]) );
  INVD0 U997 ( .I(1'b1), .ZN(n[989]) );
  INVD0 U999 ( .I(1'b1), .ZN(n[992]) );
  INVD0 U1001 ( .I(1'b1), .ZN(n[993]) );
  INVD0 U1003 ( .I(1'b1), .ZN(n[995]) );
  INVD0 U1005 ( .I(1'b1), .ZN(n[996]) );
  INVD0 U1007 ( .I(1'b1), .ZN(n[1000]) );
  INVD0 U1009 ( .I(1'b1), .ZN(n[1001]) );
  INVD0 U1011 ( .I(1'b1), .ZN(n[1003]) );
  INVD0 U1013 ( .I(1'b1), .ZN(n[1004]) );
  INVD0 U1015 ( .I(1'b1), .ZN(n[1007]) );
  INVD0 U1017 ( .I(1'b1), .ZN(n[1008]) );
  INVD0 U1019 ( .I(1'b1), .ZN(n[1010]) );
  INVD0 U1021 ( .I(1'b1), .ZN(n[1011]) );
  AN2D0 U1023 ( .A1(b[7]), .A2(n[488]), .Z(n[999]) );
  AN2D0 U1024 ( .A1(n[487]), .A2(b[7]), .Z(n[998]) );
  AN2D0 U1025 ( .A1(n[486]), .A2(b[7]), .Z(n[997]) );
  AN2D0 U1026 ( .A1(n[483]), .A2(b[7]), .Z(n[994]) );
  AN2D0 U1027 ( .A1(n[480]), .A2(b[7]), .Z(n[991]) );
  AN2D0 U1028 ( .A1(n[479]), .A2(b[7]), .Z(n[990]) );
  AN2D0 U1029 ( .A1(n[476]), .A2(b[7]), .Z(n[987]) );
  AN2D0 U1030 ( .A1(n[473]), .A2(b[7]), .Z(n[984]) );
  AN2D0 U1031 ( .A1(n[472]), .A2(b[7]), .Z(n[983]) );
  AN2D0 U1032 ( .A1(n[471]), .A2(b[7]), .Z(n[982]) );
  AN2D0 U1033 ( .A1(n[470]), .A2(b[7]), .Z(n[981]) );
  AN2D0 U1034 ( .A1(n[467]), .A2(b[7]), .Z(n[978]) );
  AN2D0 U1035 ( .A1(n[464]), .A2(b[7]), .Z(n[975]) );
  AN2D0 U1036 ( .A1(n[463]), .A2(b[7]), .Z(n[974]) );
  AN2D0 U1037 ( .A1(n[460]), .A2(b[7]), .Z(n[971]) );
  AN2D0 U1038 ( .A1(n[457]), .A2(b[7]), .Z(n[968]) );
  AN2D0 U1039 ( .A1(n[456]), .A2(b[7]), .Z(n[967]) );
  AN2D0 U1040 ( .A1(n[455]), .A2(b[7]), .Z(n[966]) );
  AN2D0 U1041 ( .A1(n[452]), .A2(b[7]), .Z(n[963]) );
  AN2D0 U1042 ( .A1(n[449]), .A2(b[7]), .Z(n[960]) );
  AN2D0 U1043 ( .A1(n[448]), .A2(b[7]), .Z(n[959]) );
  AN2D0 U1044 ( .A1(n[445]), .A2(b[7]), .Z(n[956]) );
  AN2D0 U1045 ( .A1(n[442]), .A2(b[7]), .Z(n[953]) );
  AN2D0 U1046 ( .A1(n[441]), .A2(b[7]), .Z(n[952]) );
  AN2D0 U1047 ( .A1(n[440]), .A2(b[7]), .Z(n[951]) );
  AN2D0 U1048 ( .A1(n[439]), .A2(b[7]), .Z(n[950]) );
  AN2D0 U1049 ( .A1(n[438]), .A2(b[7]), .Z(n[949]) );
  AN2D0 U1050 ( .A1(n[435]), .A2(b[7]), .Z(n[946]) );
  AN2D0 U1051 ( .A1(n[432]), .A2(b[7]), .Z(n[943]) );
  AN2D0 U1052 ( .A1(n[431]), .A2(b[7]), .Z(n[942]) );
  AN2D0 U1053 ( .A1(n[428]), .A2(b[7]), .Z(n[939]) );
  AN2D0 U1054 ( .A1(n[425]), .A2(b[7]), .Z(n[936]) );
  AN2D0 U1055 ( .A1(n[424]), .A2(b[7]), .Z(n[935]) );
  AN2D0 U1056 ( .A1(n[423]), .A2(b[7]), .Z(n[934]) );
  AN2D0 U1057 ( .A1(n[420]), .A2(b[7]), .Z(n[931]) );
  AN2D0 U1058 ( .A1(n[417]), .A2(b[7]), .Z(n[928]) );
  AN2D0 U1059 ( .A1(n[416]), .A2(b[7]), .Z(n[927]) );
  AN2D0 U1060 ( .A1(n[413]), .A2(b[7]), .Z(n[924]) );
  AN2D0 U1061 ( .A1(n[410]), .A2(b[7]), .Z(n[921]) );
  AN2D0 U1062 ( .A1(n[409]), .A2(b[7]), .Z(n[920]) );
  AN2D0 U1063 ( .A1(n[408]), .A2(b[7]), .Z(n[919]) );
  AN2D0 U1064 ( .A1(n[407]), .A2(b[7]), .Z(n[918]) );
  AN2D0 U1065 ( .A1(n[404]), .A2(b[7]), .Z(n[915]) );
  AN2D0 U1066 ( .A1(n[401]), .A2(b[7]), .Z(n[912]) );
  AN2D0 U1067 ( .A1(n[400]), .A2(b[7]), .Z(n[911]) );
  AN2D0 U1068 ( .A1(n[397]), .A2(b[7]), .Z(n[908]) );
  AN2D0 U1069 ( .A1(n[394]), .A2(b[7]), .Z(n[905]) );
  AN2D0 U1070 ( .A1(n[393]), .A2(b[7]), .Z(n[904]) );
  AN2D0 U1071 ( .A1(n[392]), .A2(b[7]), .Z(n[903]) );
  AN2D0 U1072 ( .A1(n[389]), .A2(b[7]), .Z(n[900]) );
  AN2D0 U1073 ( .A1(n[386]), .A2(b[7]), .Z(n[897]) );
  AN2D0 U1074 ( .A1(n[385]), .A2(b[7]), .Z(n[896]) );
  AN2D0 U1075 ( .A1(n[382]), .A2(b[7]), .Z(n[893]) );
  AN2D0 U1076 ( .A1(n[379]), .A2(b[7]), .Z(n[890]) );
  AN2D0 U1077 ( .A1(n[378]), .A2(b[7]), .Z(n[889]) );
  AN2D0 U1078 ( .A1(n[377]), .A2(b[7]), .Z(n[888]) );
  AN2D0 U1079 ( .A1(n[376]), .A2(b[7]), .Z(n[887]) );
  AN2D0 U1080 ( .A1(n[375]), .A2(b[7]), .Z(n[886]) );
  AN2D0 U1081 ( .A1(n[374]), .A2(b[7]), .Z(n[885]) );
  AN2D0 U1082 ( .A1(n[371]), .A2(b[7]), .Z(n[882]) );
  AN2D0 U1083 ( .A1(n[368]), .A2(b[7]), .Z(n[879]) );
  AN2D0 U1084 ( .A1(n[367]), .A2(b[7]), .Z(n[878]) );
  AN2D0 U1085 ( .A1(n[364]), .A2(b[7]), .Z(n[875]) );
  AN2D0 U1086 ( .A1(n[361]), .A2(b[7]), .Z(n[872]) );
  AN2D0 U1087 ( .A1(n[360]), .A2(b[7]), .Z(n[871]) );
  AN2D0 U1088 ( .A1(n[359]), .A2(b[7]), .Z(n[870]) );
  AN2D0 U1089 ( .A1(n[356]), .A2(b[7]), .Z(n[867]) );
  AN2D0 U1090 ( .A1(n[353]), .A2(b[7]), .Z(n[864]) );
  AN2D0 U1091 ( .A1(n[352]), .A2(b[7]), .Z(n[863]) );
  AN2D0 U1092 ( .A1(n[349]), .A2(b[7]), .Z(n[860]) );
  AN2D0 U1093 ( .A1(n[346]), .A2(b[7]), .Z(n[857]) );
  AN2D0 U1094 ( .A1(n[345]), .A2(b[7]), .Z(n[856]) );
  AN2D0 U1095 ( .A1(n[344]), .A2(b[7]), .Z(n[855]) );
  AN2D0 U1096 ( .A1(n[343]), .A2(b[7]), .Z(n[854]) );
  AN2D0 U1097 ( .A1(n[340]), .A2(b[7]), .Z(n[851]) );
  AN2D0 U1098 ( .A1(n[337]), .A2(b[7]), .Z(n[848]) );
  AN2D0 U1099 ( .A1(n[336]), .A2(b[7]), .Z(n[847]) );
  AN2D0 U1100 ( .A1(n[333]), .A2(b[7]), .Z(n[844]) );
  AN2D0 U1101 ( .A1(n[330]), .A2(b[7]), .Z(n[841]) );
  AN2D0 U1102 ( .A1(n[329]), .A2(b[7]), .Z(n[840]) );
  AN2D0 U1103 ( .A1(n[328]), .A2(b[7]), .Z(n[839]) );
  AN2D0 U1104 ( .A1(n[325]), .A2(b[7]), .Z(n[836]) );
  AN2D0 U1105 ( .A1(n[322]), .A2(b[7]), .Z(n[833]) );
  AN2D0 U1106 ( .A1(n[321]), .A2(b[7]), .Z(n[832]) );
  AN2D0 U1107 ( .A1(n[318]), .A2(b[7]), .Z(n[829]) );
  AN2D0 U1108 ( .A1(n[315]), .A2(b[7]), .Z(n[826]) );
  AN2D0 U1109 ( .A1(n[314]), .A2(b[7]), .Z(n[825]) );
  AN2D0 U1110 ( .A1(n[313]), .A2(b[7]), .Z(n[824]) );
  AN2D0 U1111 ( .A1(n[312]), .A2(b[7]), .Z(n[823]) );
  AN2D0 U1112 ( .A1(n[311]), .A2(b[7]), .Z(n[822]) );
  AN2D0 U1113 ( .A1(n[308]), .A2(b[7]), .Z(n[819]) );
  AN2D0 U1114 ( .A1(n[305]), .A2(b[7]), .Z(n[816]) );
  AN2D0 U1115 ( .A1(n[304]), .A2(b[7]), .Z(n[815]) );
  AN2D0 U1116 ( .A1(n[301]), .A2(b[7]), .Z(n[812]) );
  AN2D0 U1117 ( .A1(n[298]), .A2(b[7]), .Z(n[809]) );
  AN2D0 U1118 ( .A1(n[297]), .A2(b[7]), .Z(n[808]) );
  AN2D0 U1119 ( .A1(n[296]), .A2(b[7]), .Z(n[807]) );
  AN2D0 U1120 ( .A1(n[293]), .A2(b[7]), .Z(n[804]) );
  AN2D0 U1121 ( .A1(n[290]), .A2(b[7]), .Z(n[801]) );
  AN2D0 U1122 ( .A1(n[289]), .A2(b[7]), .Z(n[800]) );
  AN2D0 U1123 ( .A1(n[286]), .A2(b[7]), .Z(n[797]) );
  AN2D0 U1124 ( .A1(n[283]), .A2(b[7]), .Z(n[794]) );
  AN2D0 U1125 ( .A1(n[282]), .A2(b[7]), .Z(n[793]) );
  AN2D0 U1126 ( .A1(n[281]), .A2(b[7]), .Z(n[792]) );
  AN2D0 U1127 ( .A1(n[280]), .A2(b[7]), .Z(n[791]) );
  AN2D0 U1128 ( .A1(n[277]), .A2(b[7]), .Z(n[788]) );
  AN2D0 U1129 ( .A1(n[274]), .A2(b[7]), .Z(n[785]) );
  AN2D0 U1130 ( .A1(n[273]), .A2(b[7]), .Z(n[784]) );
  AN2D0 U1131 ( .A1(n[270]), .A2(b[7]), .Z(n[781]) );
  AN2D0 U1132 ( .A1(n[267]), .A2(b[7]), .Z(n[778]) );
  AN2D0 U1133 ( .A1(n[266]), .A2(b[7]), .Z(n[777]) );
  AN2D0 U1134 ( .A1(n[265]), .A2(b[7]), .Z(n[776]) );
  AN2D0 U1135 ( .A1(n[262]), .A2(b[7]), .Z(n[773]) );
  AN2D0 U1136 ( .A1(n[259]), .A2(b[7]), .Z(n[770]) );
  AN2D0 U1137 ( .A1(n[258]), .A2(b[7]), .Z(n[769]) );
  AN2D0 U1138 ( .A1(n[255]), .A2(b[7]), .Z(n[766]) );
  AN2D0 U1139 ( .A1(n[252]), .A2(b[7]), .Z(n[763]) );
  AN2D0 U1140 ( .A1(n[251]), .A2(b[7]), .Z(n[762]) );
  AN2D0 U1141 ( .A1(n[250]), .A2(b[7]), .Z(n[761]) );
  AN2D0 U1142 ( .A1(n[249]), .A2(b[7]), .Z(n[760]) );
  AN2D0 U1143 ( .A1(n[248]), .A2(b[7]), .Z(n[759]) );
  AN2D0 U1144 ( .A1(n[247]), .A2(b[7]), .Z(n[758]) );
  AN2D0 U1145 ( .A1(n[246]), .A2(b[7]), .Z(n[757]) );
  AN2D0 U1146 ( .A1(a[7]), .A2(n[498]), .Z(n[754]) );
  AN2D0 U1147 ( .A1(n[495]), .A2(a[7]), .Z(n[751]) );
  AN2D0 U1148 ( .A1(n[494]), .A2(a[7]), .Z(n[750]) );
  AN2D0 U1149 ( .A1(n[491]), .A2(a[7]), .Z(n[747]) );
  AN2D0 U1150 ( .A1(a[7]), .A2(n[488]), .Z(n[744]) );
  AN2D0 U1151 ( .A1(a[7]), .A2(n[487]), .Z(n[743]) );
  AN2D0 U1152 ( .A1(a[7]), .A2(n[486]), .Z(n[742]) );
  AN2D0 U1153 ( .A1(a[7]), .A2(n[483]), .Z(n[739]) );
  AN2D0 U1154 ( .A1(a[7]), .A2(n[480]), .Z(n[736]) );
  AN2D0 U1155 ( .A1(a[7]), .A2(n[479]), .Z(n[735]) );
  AN2D0 U1156 ( .A1(a[7]), .A2(n[476]), .Z(n[732]) );
  AN2D0 U1157 ( .A1(a[7]), .A2(n[473]), .Z(n[729]) );
  AN2D0 U1158 ( .A1(a[7]), .A2(n[472]), .Z(n[728]) );
  AN2D0 U1159 ( .A1(a[7]), .A2(n[471]), .Z(n[727]) );
  AN2D0 U1160 ( .A1(a[7]), .A2(n[470]), .Z(n[726]) );
  AN2D0 U1161 ( .A1(a[7]), .A2(n[467]), .Z(n[723]) );
  AN2D0 U1162 ( .A1(a[7]), .A2(n[464]), .Z(n[720]) );
  AN2D0 U1163 ( .A1(a[7]), .A2(n[463]), .Z(n[719]) );
  AN2D0 U1164 ( .A1(a[7]), .A2(n[460]), .Z(n[716]) );
  AN2D0 U1165 ( .A1(a[7]), .A2(n[457]), .Z(n[713]) );
  AN2D0 U1166 ( .A1(a[7]), .A2(n[456]), .Z(n[712]) );
  AN2D0 U1167 ( .A1(a[7]), .A2(n[455]), .Z(n[711]) );
  AN2D0 U1168 ( .A1(a[7]), .A2(n[452]), .Z(n[708]) );
  AN2D0 U1169 ( .A1(a[7]), .A2(n[449]), .Z(n[705]) );
  AN2D0 U1170 ( .A1(a[7]), .A2(n[448]), .Z(n[704]) );
  AN2D0 U1171 ( .A1(a[7]), .A2(n[445]), .Z(n[701]) );
  AN2D0 U1172 ( .A1(a[7]), .A2(n[442]), .Z(n[698]) );
  AN2D0 U1173 ( .A1(a[7]), .A2(n[441]), .Z(n[697]) );
  AN2D0 U1174 ( .A1(a[7]), .A2(n[440]), .Z(n[696]) );
  AN2D0 U1175 ( .A1(a[7]), .A2(n[439]), .Z(n[695]) );
  AN2D0 U1176 ( .A1(a[7]), .A2(n[438]), .Z(n[694]) );
  AN2D0 U1177 ( .A1(a[7]), .A2(n[435]), .Z(n[691]) );
  AN2D0 U1178 ( .A1(a[7]), .A2(n[432]), .Z(n[688]) );
  AN2D0 U1179 ( .A1(a[7]), .A2(n[431]), .Z(n[687]) );
  AN2D0 U1180 ( .A1(a[7]), .A2(n[428]), .Z(n[684]) );
  AN2D0 U1181 ( .A1(a[7]), .A2(n[425]), .Z(n[681]) );
  AN2D0 U1182 ( .A1(a[7]), .A2(n[424]), .Z(n[680]) );
  AN2D0 U1183 ( .A1(a[7]), .A2(n[423]), .Z(n[679]) );
  AN2D0 U1184 ( .A1(a[7]), .A2(n[420]), .Z(n[676]) );
  AN2D0 U1185 ( .A1(a[7]), .A2(n[417]), .Z(n[673]) );
  AN2D0 U1186 ( .A1(a[7]), .A2(n[416]), .Z(n[672]) );
  AN2D0 U1187 ( .A1(a[7]), .A2(n[413]), .Z(n[669]) );
  AN2D0 U1188 ( .A1(a[7]), .A2(n[410]), .Z(n[666]) );
  AN2D0 U1189 ( .A1(a[7]), .A2(n[409]), .Z(n[665]) );
  AN2D0 U1190 ( .A1(a[7]), .A2(n[408]), .Z(n[664]) );
  AN2D0 U1191 ( .A1(a[7]), .A2(n[407]), .Z(n[663]) );
  AN2D0 U1192 ( .A1(a[7]), .A2(n[404]), .Z(n[660]) );
  AN2D0 U1193 ( .A1(a[7]), .A2(n[401]), .Z(n[657]) );
  AN2D0 U1194 ( .A1(a[7]), .A2(n[400]), .Z(n[656]) );
  AN2D0 U1195 ( .A1(a[7]), .A2(n[397]), .Z(n[653]) );
  AN2D0 U1196 ( .A1(a[7]), .A2(n[394]), .Z(n[650]) );
  AN2D0 U1197 ( .A1(a[7]), .A2(n[393]), .Z(n[649]) );
  AN2D0 U1198 ( .A1(a[7]), .A2(n[392]), .Z(n[648]) );
  AN2D0 U1199 ( .A1(a[7]), .A2(n[389]), .Z(n[645]) );
  AN2D0 U1200 ( .A1(a[7]), .A2(n[386]), .Z(n[642]) );
  AN2D0 U1201 ( .A1(a[7]), .A2(n[385]), .Z(n[641]) );
  AN2D0 U1202 ( .A1(a[7]), .A2(n[382]), .Z(n[638]) );
  AN2D0 U1203 ( .A1(a[7]), .A2(n[379]), .Z(n[635]) );
  AN2D0 U1204 ( .A1(a[7]), .A2(n[378]), .Z(n[634]) );
  AN2D0 U1205 ( .A1(a[7]), .A2(n[377]), .Z(n[633]) );
  AN2D0 U1206 ( .A1(a[7]), .A2(n[376]), .Z(n[632]) );
  AN2D0 U1207 ( .A1(a[7]), .A2(n[375]), .Z(n[631]) );
  AN2D0 U1208 ( .A1(a[7]), .A2(n[374]), .Z(n[630]) );
  AN2D0 U1209 ( .A1(a[7]), .A2(n[371]), .Z(n[627]) );
  AN2D0 U1210 ( .A1(a[7]), .A2(n[368]), .Z(n[624]) );
  AN2D0 U1211 ( .A1(a[7]), .A2(n[367]), .Z(n[623]) );
  AN2D0 U1212 ( .A1(a[7]), .A2(n[364]), .Z(n[620]) );
  AN2D0 U1213 ( .A1(a[7]), .A2(n[361]), .Z(n[617]) );
  AN2D0 U1214 ( .A1(a[7]), .A2(n[360]), .Z(n[616]) );
  AN2D0 U1215 ( .A1(a[7]), .A2(n[359]), .Z(n[615]) );
  AN2D0 U1216 ( .A1(a[7]), .A2(n[356]), .Z(n[612]) );
  AN2D0 U1217 ( .A1(a[7]), .A2(n[353]), .Z(n[609]) );
  AN2D0 U1218 ( .A1(a[7]), .A2(n[352]), .Z(n[608]) );
  AN2D0 U1219 ( .A1(a[7]), .A2(n[349]), .Z(n[605]) );
  AN2D0 U1220 ( .A1(a[7]), .A2(n[346]), .Z(n[602]) );
  AN2D0 U1221 ( .A1(a[7]), .A2(n[345]), .Z(n[601]) );
  AN2D0 U1222 ( .A1(a[7]), .A2(n[344]), .Z(n[600]) );
  AN2D0 U1223 ( .A1(a[7]), .A2(n[343]), .Z(n[599]) );
  AN2D0 U1224 ( .A1(a[7]), .A2(n[340]), .Z(n[596]) );
  AN2D0 U1225 ( .A1(a[7]), .A2(n[337]), .Z(n[593]) );
  AN2D0 U1226 ( .A1(a[7]), .A2(n[336]), .Z(n[592]) );
  AN2D0 U1227 ( .A1(a[7]), .A2(n[333]), .Z(n[589]) );
  AN2D0 U1228 ( .A1(a[7]), .A2(n[330]), .Z(n[586]) );
  AN2D0 U1229 ( .A1(a[7]), .A2(n[329]), .Z(n[585]) );
  AN2D0 U1230 ( .A1(a[7]), .A2(n[328]), .Z(n[584]) );
  AN2D0 U1231 ( .A1(a[7]), .A2(n[325]), .Z(n[581]) );
  AN2D0 U1232 ( .A1(a[7]), .A2(n[322]), .Z(n[578]) );
  AN2D0 U1233 ( .A1(a[7]), .A2(n[321]), .Z(n[577]) );
  AN2D0 U1234 ( .A1(a[7]), .A2(n[318]), .Z(n[574]) );
  AN2D0 U1235 ( .A1(a[7]), .A2(n[315]), .Z(n[571]) );
  AN2D0 U1236 ( .A1(a[7]), .A2(n[314]), .Z(n[570]) );
  AN2D0 U1237 ( .A1(a[7]), .A2(n[313]), .Z(n[569]) );
  AN2D0 U1238 ( .A1(a[7]), .A2(n[312]), .Z(n[568]) );
  AN2D0 U1239 ( .A1(a[7]), .A2(n[311]), .Z(n[567]) );
  AN2D0 U1240 ( .A1(a[7]), .A2(n[308]), .Z(n[564]) );
  AN2D0 U1241 ( .A1(a[7]), .A2(n[305]), .Z(n[561]) );
  AN2D0 U1242 ( .A1(a[7]), .A2(n[304]), .Z(n[560]) );
  AN2D0 U1243 ( .A1(a[7]), .A2(n[301]), .Z(n[557]) );
  AN2D0 U1244 ( .A1(a[7]), .A2(n[298]), .Z(n[554]) );
  AN2D0 U1245 ( .A1(a[7]), .A2(n[297]), .Z(n[553]) );
  AN2D0 U1246 ( .A1(a[7]), .A2(n[296]), .Z(n[552]) );
  AN2D0 U1247 ( .A1(a[7]), .A2(n[293]), .Z(n[549]) );
  AN2D0 U1248 ( .A1(a[7]), .A2(n[290]), .Z(n[546]) );
  AN2D0 U1249 ( .A1(a[7]), .A2(n[289]), .Z(n[545]) );
  AN2D0 U1250 ( .A1(a[7]), .A2(n[286]), .Z(n[542]) );
  AN2D0 U1251 ( .A1(a[7]), .A2(n[283]), .Z(n[539]) );
  AN2D0 U1252 ( .A1(a[7]), .A2(n[282]), .Z(n[538]) );
  AN2D0 U1253 ( .A1(a[7]), .A2(n[281]), .Z(n[537]) );
  AN2D0 U1254 ( .A1(a[7]), .A2(n[280]), .Z(n[536]) );
  AN2D0 U1255 ( .A1(a[7]), .A2(n[277]), .Z(n[533]) );
  AN2D0 U1256 ( .A1(a[7]), .A2(n[274]), .Z(n[530]) );
  AN2D0 U1257 ( .A1(a[7]), .A2(n[273]), .Z(n[529]) );
  AN2D0 U1258 ( .A1(a[7]), .A2(n[270]), .Z(n[526]) );
  AN2D0 U1259 ( .A1(a[7]), .A2(n[267]), .Z(n[523]) );
  AN2D0 U1260 ( .A1(a[7]), .A2(n[266]), .Z(n[522]) );
  AN2D0 U1261 ( .A1(a[7]), .A2(n[265]), .Z(n[521]) );
  AN2D0 U1262 ( .A1(a[7]), .A2(n[262]), .Z(n[518]) );
  AN2D0 U1263 ( .A1(a[7]), .A2(n[259]), .Z(n[515]) );
  AN2D0 U1264 ( .A1(a[7]), .A2(n[258]), .Z(n[514]) );
  AN2D0 U1265 ( .A1(a[7]), .A2(n[255]), .Z(n[511]) );
  AN2D0 U1266 ( .A1(a[7]), .A2(n[252]), .Z(n[508]) );
  AN2D0 U1267 ( .A1(a[7]), .A2(n[251]), .Z(n[507]) );
  AN2D0 U1268 ( .A1(a[7]), .A2(n[250]), .Z(n[506]) );
  AN2D0 U1269 ( .A1(a[7]), .A2(n[249]), .Z(n[505]) );
  AN2D0 U1270 ( .A1(a[7]), .A2(n[248]), .Z(n[504]) );
  AN2D0 U1271 ( .A1(a[7]), .A2(n[247]), .Z(n[503]) );
  AN2D0 U1272 ( .A1(a[7]), .A2(n[246]), .Z(n[502]) );
  AN2D0 U1273 ( .A1(a[7]), .A2(b[7]), .Z(n[501]) );
  AN2D0 U1274 ( .A1(n[233]), .A2(b[6]), .Z(n[488]) );
  AN2D0 U1275 ( .A1(b[6]), .A2(n[232]), .Z(n[487]) );
  AN2D0 U1276 ( .A1(b[6]), .A2(n[231]), .Z(n[486]) );
  AN2D0 U1277 ( .A1(b[6]), .A2(n[228]), .Z(n[483]) );
  AN2D0 U1278 ( .A1(b[6]), .A2(n[225]), .Z(n[480]) );
  AN2D0 U1279 ( .A1(b[6]), .A2(n[224]), .Z(n[479]) );
  AN2D0 U1280 ( .A1(b[6]), .A2(n[221]), .Z(n[476]) );
  AN2D0 U1281 ( .A1(b[6]), .A2(n[218]), .Z(n[473]) );
  AN2D0 U1282 ( .A1(b[6]), .A2(n[217]), .Z(n[472]) );
  AN2D0 U1283 ( .A1(b[6]), .A2(n[216]), .Z(n[471]) );
  AN2D0 U1284 ( .A1(b[6]), .A2(n[215]), .Z(n[470]) );
  AN2D0 U1285 ( .A1(b[6]), .A2(n[212]), .Z(n[467]) );
  AN2D0 U1286 ( .A1(b[6]), .A2(n[209]), .Z(n[464]) );
  AN2D0 U1287 ( .A1(b[6]), .A2(n[208]), .Z(n[463]) );
  AN2D0 U1288 ( .A1(b[6]), .A2(n[205]), .Z(n[460]) );
  AN2D0 U1289 ( .A1(b[6]), .A2(n[202]), .Z(n[457]) );
  AN2D0 U1290 ( .A1(b[6]), .A2(n[201]), .Z(n[456]) );
  AN2D0 U1291 ( .A1(b[6]), .A2(n[200]), .Z(n[455]) );
  AN2D0 U1292 ( .A1(b[6]), .A2(n[197]), .Z(n[452]) );
  AN2D0 U1293 ( .A1(b[6]), .A2(n[194]), .Z(n[449]) );
  AN2D0 U1294 ( .A1(b[6]), .A2(n[193]), .Z(n[448]) );
  AN2D0 U1295 ( .A1(b[6]), .A2(n[190]), .Z(n[445]) );
  AN2D0 U1296 ( .A1(b[6]), .A2(n[187]), .Z(n[442]) );
  AN2D0 U1297 ( .A1(b[6]), .A2(n[186]), .Z(n[441]) );
  AN2D0 U1298 ( .A1(b[6]), .A2(n[185]), .Z(n[440]) );
  AN2D0 U1299 ( .A1(b[6]), .A2(n[184]), .Z(n[439]) );
  AN2D0 U1300 ( .A1(b[6]), .A2(n[183]), .Z(n[438]) );
  AN2D0 U1301 ( .A1(b[6]), .A2(n[180]), .Z(n[435]) );
  AN2D0 U1302 ( .A1(b[6]), .A2(n[177]), .Z(n[432]) );
  AN2D0 U1303 ( .A1(b[6]), .A2(n[176]), .Z(n[431]) );
  AN2D0 U1304 ( .A1(b[6]), .A2(n[173]), .Z(n[428]) );
  AN2D0 U1305 ( .A1(b[6]), .A2(n[170]), .Z(n[425]) );
  AN2D0 U1306 ( .A1(b[6]), .A2(n[169]), .Z(n[424]) );
  AN2D0 U1307 ( .A1(b[6]), .A2(n[168]), .Z(n[423]) );
  AN2D0 U1308 ( .A1(b[6]), .A2(n[165]), .Z(n[420]) );
  AN2D0 U1309 ( .A1(b[6]), .A2(n[162]), .Z(n[417]) );
  AN2D0 U1310 ( .A1(b[6]), .A2(n[161]), .Z(n[416]) );
  AN2D0 U1311 ( .A1(b[6]), .A2(n[158]), .Z(n[413]) );
  AN2D0 U1312 ( .A1(b[6]), .A2(n[155]), .Z(n[410]) );
  AN2D0 U1313 ( .A1(b[6]), .A2(n[154]), .Z(n[409]) );
  AN2D0 U1314 ( .A1(b[6]), .A2(n[153]), .Z(n[408]) );
  AN2D0 U1315 ( .A1(b[6]), .A2(n[152]), .Z(n[407]) );
  AN2D0 U1316 ( .A1(b[6]), .A2(n[149]), .Z(n[404]) );
  AN2D0 U1317 ( .A1(b[6]), .A2(n[146]), .Z(n[401]) );
  AN2D0 U1318 ( .A1(b[6]), .A2(n[145]), .Z(n[400]) );
  AN2D0 U1319 ( .A1(b[6]), .A2(n[142]), .Z(n[397]) );
  AN2D0 U1320 ( .A1(b[6]), .A2(n[139]), .Z(n[394]) );
  AN2D0 U1321 ( .A1(b[6]), .A2(n[138]), .Z(n[393]) );
  AN2D0 U1322 ( .A1(b[6]), .A2(n[137]), .Z(n[392]) );
  AN2D0 U1323 ( .A1(b[6]), .A2(n[134]), .Z(n[389]) );
  AN2D0 U1324 ( .A1(b[6]), .A2(n[131]), .Z(n[386]) );
  AN2D0 U1325 ( .A1(b[6]), .A2(n[130]), .Z(n[385]) );
  AN2D0 U1326 ( .A1(b[6]), .A2(n[127]), .Z(n[382]) );
  AN2D0 U1327 ( .A1(b[6]), .A2(n[124]), .Z(n[379]) );
  AN2D0 U1328 ( .A1(b[6]), .A2(n[123]), .Z(n[378]) );
  AN2D0 U1329 ( .A1(b[6]), .A2(n[122]), .Z(n[377]) );
  AN2D0 U1330 ( .A1(b[6]), .A2(n[121]), .Z(n[376]) );
  AN2D0 U1331 ( .A1(b[6]), .A2(n[120]), .Z(n[375]) );
  AN2D0 U1332 ( .A1(b[6]), .A2(n[119]), .Z(n[374]) );
  AN2D0 U1333 ( .A1(n[243]), .A2(a[6]), .Z(n[371]) );
  AN2D0 U1334 ( .A1(a[6]), .A2(n[240]), .Z(n[368]) );
  AN2D0 U1335 ( .A1(a[6]), .A2(n[239]), .Z(n[367]) );
  AN2D0 U1336 ( .A1(a[6]), .A2(n[236]), .Z(n[364]) );
  AN2D0 U1337 ( .A1(n[233]), .A2(a[6]), .Z(n[361]) );
  AN2D0 U1338 ( .A1(n[232]), .A2(a[6]), .Z(n[360]) );
  AN2D0 U1339 ( .A1(n[231]), .A2(a[6]), .Z(n[359]) );
  AN2D0 U1340 ( .A1(n[228]), .A2(a[6]), .Z(n[356]) );
  AN2D0 U1341 ( .A1(n[225]), .A2(a[6]), .Z(n[353]) );
  AN2D0 U1342 ( .A1(n[224]), .A2(a[6]), .Z(n[352]) );
  AN2D0 U1343 ( .A1(n[221]), .A2(a[6]), .Z(n[349]) );
  AN2D0 U1344 ( .A1(n[218]), .A2(a[6]), .Z(n[346]) );
  AN2D0 U1345 ( .A1(n[217]), .A2(a[6]), .Z(n[345]) );
  AN2D0 U1346 ( .A1(n[216]), .A2(a[6]), .Z(n[344]) );
  AN2D0 U1347 ( .A1(n[215]), .A2(a[6]), .Z(n[343]) );
  AN2D0 U1348 ( .A1(n[212]), .A2(a[6]), .Z(n[340]) );
  AN2D0 U1349 ( .A1(n[209]), .A2(a[6]), .Z(n[337]) );
  AN2D0 U1350 ( .A1(n[208]), .A2(a[6]), .Z(n[336]) );
  AN2D0 U1351 ( .A1(n[205]), .A2(a[6]), .Z(n[333]) );
  AN2D0 U1352 ( .A1(n[202]), .A2(a[6]), .Z(n[330]) );
  AN2D0 U1353 ( .A1(n[201]), .A2(a[6]), .Z(n[329]) );
  AN2D0 U1354 ( .A1(n[200]), .A2(a[6]), .Z(n[328]) );
  AN2D0 U1355 ( .A1(n[197]), .A2(a[6]), .Z(n[325]) );
  AN2D0 U1356 ( .A1(n[194]), .A2(a[6]), .Z(n[322]) );
  AN2D0 U1357 ( .A1(n[193]), .A2(a[6]), .Z(n[321]) );
  AN2D0 U1358 ( .A1(n[190]), .A2(a[6]), .Z(n[318]) );
  AN2D0 U1359 ( .A1(n[187]), .A2(a[6]), .Z(n[315]) );
  AN2D0 U1360 ( .A1(n[186]), .A2(a[6]), .Z(n[314]) );
  AN2D0 U1361 ( .A1(n[185]), .A2(a[6]), .Z(n[313]) );
  AN2D0 U1362 ( .A1(n[184]), .A2(a[6]), .Z(n[312]) );
  AN2D0 U1363 ( .A1(n[183]), .A2(a[6]), .Z(n[311]) );
  AN2D0 U1364 ( .A1(n[180]), .A2(a[6]), .Z(n[308]) );
  AN2D0 U1365 ( .A1(n[177]), .A2(a[6]), .Z(n[305]) );
  AN2D0 U1366 ( .A1(n[176]), .A2(a[6]), .Z(n[304]) );
  AN2D0 U1367 ( .A1(n[173]), .A2(a[6]), .Z(n[301]) );
  AN2D0 U1368 ( .A1(n[170]), .A2(a[6]), .Z(n[298]) );
  AN2D0 U1369 ( .A1(n[169]), .A2(a[6]), .Z(n[297]) );
  AN2D0 U1370 ( .A1(n[168]), .A2(a[6]), .Z(n[296]) );
  AN2D0 U1371 ( .A1(n[165]), .A2(a[6]), .Z(n[293]) );
  AN2D0 U1372 ( .A1(n[162]), .A2(a[6]), .Z(n[290]) );
  AN2D0 U1373 ( .A1(n[161]), .A2(a[6]), .Z(n[289]) );
  AN2D0 U1374 ( .A1(n[158]), .A2(a[6]), .Z(n[286]) );
  AN2D0 U1375 ( .A1(n[155]), .A2(a[6]), .Z(n[283]) );
  AN2D0 U1376 ( .A1(n[154]), .A2(a[6]), .Z(n[282]) );
  AN2D0 U1377 ( .A1(n[153]), .A2(a[6]), .Z(n[281]) );
  AN2D0 U1378 ( .A1(n[152]), .A2(a[6]), .Z(n[280]) );
  AN2D0 U1379 ( .A1(n[149]), .A2(a[6]), .Z(n[277]) );
  AN2D0 U1380 ( .A1(n[146]), .A2(a[6]), .Z(n[274]) );
  AN2D0 U1381 ( .A1(n[145]), .A2(a[6]), .Z(n[273]) );
  AN2D0 U1382 ( .A1(n[142]), .A2(a[6]), .Z(n[270]) );
  AN2D0 U1383 ( .A1(n[139]), .A2(a[6]), .Z(n[267]) );
  AN2D0 U1384 ( .A1(n[138]), .A2(a[6]), .Z(n[266]) );
  AN2D0 U1385 ( .A1(n[137]), .A2(a[6]), .Z(n[265]) );
  AN2D0 U1386 ( .A1(n[134]), .A2(a[6]), .Z(n[262]) );
  AN2D0 U1387 ( .A1(n[131]), .A2(a[6]), .Z(n[259]) );
  AN2D0 U1388 ( .A1(n[130]), .A2(a[6]), .Z(n[258]) );
  AN2D0 U1389 ( .A1(n[127]), .A2(a[6]), .Z(n[255]) );
  AN2D0 U1390 ( .A1(n[124]), .A2(a[6]), .Z(n[252]) );
  AN2D0 U1391 ( .A1(n[123]), .A2(a[6]), .Z(n[251]) );
  AN2D0 U1392 ( .A1(n[122]), .A2(a[6]), .Z(n[250]) );
  AN2D0 U1393 ( .A1(n[121]), .A2(a[6]), .Z(n[249]) );
  AN2D0 U1394 ( .A1(n[120]), .A2(a[6]), .Z(n[248]) );
  AN2D0 U1395 ( .A1(n[119]), .A2(a[6]), .Z(n[247]) );
  AN2D0 U1396 ( .A1(b[6]), .A2(a[6]), .Z(n[246]) );
  AN2D0 U1397 ( .A1(n[106]), .A2(b[5]), .Z(n[233]) );
  AN2D0 U1398 ( .A1(b[5]), .A2(n[105]), .Z(n[232]) );
  AN2D0 U1399 ( .A1(b[5]), .A2(n[104]), .Z(n[231]) );
  AN2D0 U1400 ( .A1(b[5]), .A2(n[101]), .Z(n[228]) );
  AN2D0 U1401 ( .A1(b[5]), .A2(n[98]), .Z(n[225]) );
  AN2D0 U1402 ( .A1(b[5]), .A2(n[97]), .Z(n[224]) );
  AN2D0 U1403 ( .A1(b[5]), .A2(n[94]), .Z(n[221]) );
  AN2D0 U1404 ( .A1(b[5]), .A2(n[91]), .Z(n[218]) );
  AN2D0 U1405 ( .A1(b[5]), .A2(n[90]), .Z(n[217]) );
  AN2D0 U1406 ( .A1(b[5]), .A2(n[89]), .Z(n[216]) );
  AN2D0 U1407 ( .A1(b[5]), .A2(n[88]), .Z(n[215]) );
  AN2D0 U1408 ( .A1(b[5]), .A2(n[85]), .Z(n[212]) );
  AN2D0 U1409 ( .A1(b[5]), .A2(n[82]), .Z(n[209]) );
  AN2D0 U1410 ( .A1(b[5]), .A2(n[81]), .Z(n[208]) );
  AN2D0 U1411 ( .A1(b[5]), .A2(n[78]), .Z(n[205]) );
  AN2D0 U1412 ( .A1(b[5]), .A2(n[75]), .Z(n[202]) );
  AN2D0 U1413 ( .A1(b[5]), .A2(n[74]), .Z(n[201]) );
  AN2D0 U1414 ( .A1(b[5]), .A2(n[73]), .Z(n[200]) );
  AN2D0 U1415 ( .A1(b[5]), .A2(n[70]), .Z(n[197]) );
  AN2D0 U1416 ( .A1(b[5]), .A2(n[67]), .Z(n[194]) );
  AN2D0 U1417 ( .A1(b[5]), .A2(n[66]), .Z(n[193]) );
  AN2D0 U1418 ( .A1(b[5]), .A2(n[63]), .Z(n[190]) );
  AN2D0 U1419 ( .A1(b[5]), .A2(n[60]), .Z(n[187]) );
  AN2D0 U1420 ( .A1(b[5]), .A2(n[59]), .Z(n[186]) );
  AN2D0 U1421 ( .A1(b[5]), .A2(n[58]), .Z(n[185]) );
  AN2D0 U1422 ( .A1(b[5]), .A2(n[57]), .Z(n[184]) );
  AN2D0 U1423 ( .A1(b[5]), .A2(n[56]), .Z(n[183]) );
  AN2D0 U1424 ( .A1(n[116]), .A2(a[5]), .Z(n[180]) );
  AN2D0 U1425 ( .A1(a[5]), .A2(n[113]), .Z(n[177]) );
  AN2D0 U1426 ( .A1(a[5]), .A2(n[112]), .Z(n[176]) );
  AN2D0 U1427 ( .A1(a[5]), .A2(n[109]), .Z(n[173]) );
  AN2D0 U1428 ( .A1(n[106]), .A2(a[5]), .Z(n[170]) );
  AN2D0 U1429 ( .A1(n[105]), .A2(a[5]), .Z(n[169]) );
  AN2D0 U1430 ( .A1(n[104]), .A2(a[5]), .Z(n[168]) );
  AN2D0 U1431 ( .A1(n[101]), .A2(a[5]), .Z(n[165]) );
  AN2D0 U1432 ( .A1(n[98]), .A2(a[5]), .Z(n[162]) );
  AN2D0 U1433 ( .A1(b[4]), .A2(n[35]), .Z(n[98]) );
  AN2D0 U1434 ( .A1(n[97]), .A2(a[5]), .Z(n[161]) );
  AN2D0 U1435 ( .A1(b[4]), .A2(n[34]), .Z(n[97]) );
  AN2D0 U1436 ( .A1(n[94]), .A2(a[5]), .Z(n[158]) );
  AN2D0 U1437 ( .A1(b[4]), .A2(n[31]), .Z(n[94]) );
  AN2D0 U1438 ( .A1(n[91]), .A2(a[5]), .Z(n[155]) );
  AN2D0 U1439 ( .A1(b[4]), .A2(n[28]), .Z(n[91]) );
  AN2D0 U1440 ( .A1(n[90]), .A2(a[5]), .Z(n[154]) );
  AN2D0 U1441 ( .A1(b[4]), .A2(n[27]), .Z(n[90]) );
  AN2D0 U1442 ( .A1(n[89]), .A2(a[5]), .Z(n[153]) );
  AN2D0 U1443 ( .A1(b[4]), .A2(n[26]), .Z(n[89]) );
  AN2D0 U1444 ( .A1(n[88]), .A2(a[5]), .Z(n[152]) );
  AN2D0 U1445 ( .A1(b[4]), .A2(n[25]), .Z(n[88]) );
  AN2D0 U1446 ( .A1(n[85]), .A2(a[5]), .Z(n[149]) );
  AN2D0 U1447 ( .A1(n[53]), .A2(a[4]), .Z(n[85]) );
  AN2D0 U1448 ( .A1(n[82]), .A2(a[5]), .Z(n[146]) );
  AN2D0 U1449 ( .A1(a[4]), .A2(n[50]), .Z(n[82]) );
  AN2D0 U1450 ( .A1(n[81]), .A2(a[5]), .Z(n[145]) );
  AN2D0 U1451 ( .A1(a[4]), .A2(n[49]), .Z(n[81]) );
  AN2D0 U1452 ( .A1(n[78]), .A2(a[5]), .Z(n[142]) );
  AN2D0 U1453 ( .A1(a[4]), .A2(n[46]), .Z(n[78]) );
  AN2D0 U1454 ( .A1(n[75]), .A2(a[5]), .Z(n[139]) );
  AN2D0 U1455 ( .A1(n[43]), .A2(a[4]), .Z(n[75]) );
  AN2D0 U1456 ( .A1(n[74]), .A2(a[5]), .Z(n[138]) );
  AN2D0 U1457 ( .A1(n[42]), .A2(a[4]), .Z(n[74]) );
  AN2D0 U1458 ( .A1(n[73]), .A2(a[5]), .Z(n[137]) );
  AN2D0 U1459 ( .A1(n[41]), .A2(a[4]), .Z(n[73]) );
  AN2D0 U1460 ( .A1(n[70]), .A2(a[5]), .Z(n[134]) );
  AN2D0 U1461 ( .A1(n[38]), .A2(a[4]), .Z(n[70]) );
  AN2D0 U1462 ( .A1(n[67]), .A2(a[5]), .Z(n[131]) );
  AN2D0 U1463 ( .A1(n[35]), .A2(a[4]), .Z(n[67]) );
  AN2D0 U1464 ( .A1(a[3]), .A2(n[19]), .Z(n[35]) );
  AN2D0 U1465 ( .A1(n[66]), .A2(a[5]), .Z(n[130]) );
  AN2D0 U1466 ( .A1(n[34]), .A2(a[4]), .Z(n[66]) );
  AN2D0 U1467 ( .A1(a[3]), .A2(n[18]), .Z(n[34]) );
  AN2D0 U1468 ( .A1(n[63]), .A2(a[5]), .Z(n[127]) );
  AN2D0 U1469 ( .A1(n[31]), .A2(a[4]), .Z(n[63]) );
  AN2D0 U1470 ( .A1(a[3]), .A2(n[15]), .Z(n[31]) );
  AN2D0 U1471 ( .A1(n[60]), .A2(a[5]), .Z(n[124]) );
  AN2D0 U1472 ( .A1(n[28]), .A2(a[4]), .Z(n[60]) );
  AN2D0 U1473 ( .A1(n[12]), .A2(a[3]), .Z(n[28]) );
  AN2D0 U1474 ( .A1(n[59]), .A2(a[5]), .Z(n[123]) );
  AN2D0 U1475 ( .A1(n[27]), .A2(a[4]), .Z(n[59]) );
  AN2D0 U1476 ( .A1(n[11]), .A2(a[3]), .Z(n[27]) );
  AN2D0 U1477 ( .A1(n[58]), .A2(a[5]), .Z(n[122]) );
  AN2D0 U1478 ( .A1(n[26]), .A2(a[4]), .Z(n[58]) );
  AN2D0 U1479 ( .A1(n[10]), .A2(a[3]), .Z(n[26]) );
  AN2D0 U1480 ( .A1(n[57]), .A2(a[5]), .Z(n[121]) );
  AN2D0 U1481 ( .A1(n[25]), .A2(a[4]), .Z(n[57]) );
  AN2D0 U1482 ( .A1(b[3]), .A2(a[3]), .Z(n[25]) );
  AN2D0 U1483 ( .A1(n[56]), .A2(a[5]), .Z(n[120]) );
  AN2D0 U1484 ( .A1(b[4]), .A2(a[4]), .Z(n[56]) );
  AN2D0 U1485 ( .A1(b[5]), .A2(a[5]), .Z(n[119]) );
  AN2D0 U1486 ( .A1(n[43]), .A2(b[4]), .Z(n[106]) );
  AN2D0 U1487 ( .A1(n[12]), .A2(b[3]), .Z(n[43]) );
  AN2D0 U1488 ( .A1(n[4]), .A2(a[2]), .Z(n[12]) );
  AN2D0 U1489 ( .A1(b[4]), .A2(n[42]), .Z(n[105]) );
  AN2D0 U1490 ( .A1(b[3]), .A2(n[11]), .Z(n[42]) );
  AN2D0 U1491 ( .A1(a[2]), .A2(n[3]), .Z(n[11]) );
  AN2D0 U1492 ( .A1(b[4]), .A2(n[41]), .Z(n[104]) );
  AN2D0 U1493 ( .A1(b[3]), .A2(n[10]), .Z(n[41]) );
  AN2D0 U1494 ( .A1(a[2]), .A2(b[2]), .Z(n[10]) );
  AN2D0 U1495 ( .A1(b[4]), .A2(n[38]), .Z(n[101]) );
  AN2D0 U1496 ( .A1(n[22]), .A2(a[3]), .Z(n[38]) );
  AN2D0 U1497 ( .A1(n[498]), .A2(b[7]), .Z(n[1009]) );
  AN2D0 U1498 ( .A1(b[6]), .A2(n[243]), .Z(n[498]) );
  AN2D0 U1499 ( .A1(b[5]), .A2(n[116]), .Z(n[243]) );
  AN2D0 U1500 ( .A1(b[4]), .A2(n[53]), .Z(n[116]) );
  AN2D0 U1501 ( .A1(b[3]), .A2(n[22]), .Z(n[53]) );
  AN2D0 U1502 ( .A1(b[2]), .A2(n[7]), .Z(n[22]) );
  AN2D0 U1503 ( .A1(n[495]), .A2(b[7]), .Z(n[1006]) );
  AN2D0 U1504 ( .A1(b[6]), .A2(n[240]), .Z(n[495]) );
  AN2D0 U1505 ( .A1(b[5]), .A2(n[113]), .Z(n[240]) );
  AN2D0 U1506 ( .A1(b[4]), .A2(n[50]), .Z(n[113]) );
  AN2D0 U1507 ( .A1(b[3]), .A2(n[19]), .Z(n[50]) );
  AN2D0 U1508 ( .A1(n[4]), .A2(b[2]), .Z(n[19]) );
  AN2D0 U1509 ( .A1(n[0]), .A2(a[1]), .Z(n[4]) );
  AN2D0 U1510 ( .A1(n[494]), .A2(b[7]), .Z(n[1005]) );
  AN2D0 U1511 ( .A1(b[6]), .A2(n[239]), .Z(n[494]) );
  AN2D0 U1512 ( .A1(b[5]), .A2(n[112]), .Z(n[239]) );
  AN2D0 U1513 ( .A1(b[4]), .A2(n[49]), .Z(n[112]) );
  AN2D0 U1514 ( .A1(b[3]), .A2(n[18]), .Z(n[49]) );
  AN2D0 U1515 ( .A1(n[3]), .A2(b[2]), .Z(n[18]) );
  AN2D0 U1516 ( .A1(a[1]), .A2(b[1]), .Z(n[3]) );
  AN2D0 U1517 ( .A1(n[491]), .A2(b[7]), .Z(n[1002]) );
  AN2D0 U1518 ( .A1(b[6]), .A2(n[236]), .Z(n[491]) );
  AN2D0 U1519 ( .A1(b[5]), .A2(n[109]), .Z(n[236]) );
  AN2D0 U1520 ( .A1(b[4]), .A2(n[46]), .Z(n[109]) );
  AN2D0 U1521 ( .A1(b[3]), .A2(n[15]), .Z(n[46]) );
  AN2D0 U1522 ( .A1(a[2]), .A2(n[7]), .Z(n[15]) );
  AN2D0 U1523 ( .A1(n[0]), .A2(b[1]), .Z(n[7]) );
  AN2D0 U1524 ( .A1(b[0]), .A2(a[0]), .Z(n[0]) );
endmodule


module gen_cla_decomposed ( a, b, s );
  input [8:0] a;
  input [8:0] b;
  output [8:0] s;

  wire   [1011:0] n;

  gen_nonlinear_part NLIN ( .a(a), .b(b), .n(n) );
  gen_linear_part LIN ( .a(a), .b(b), .n({1'b0, 1'b0, n[1009], 1'b0, 1'b0, 
        n[1006:1005], 1'b0, 1'b0, n[1002], 1'b0, 1'b0, n[999:997], 1'b0, 1'b0, 
        n[994], 1'b0, 1'b0, n[991:990], 1'b0, 1'b0, n[987], 1'b0, 1'b0, 
        n[984:981], 1'b0, 1'b0, n[978], 1'b0, 1'b0, n[975:974], 1'b0, 1'b0, 
        n[971], 1'b0, 1'b0, n[968:966], 1'b0, 1'b0, n[963], 1'b0, 1'b0, 
        n[960:959], 1'b0, 1'b0, n[956], 1'b0, 1'b0, n[953:949], 1'b0, 1'b0, 
        n[946], 1'b0, 1'b0, n[943:942], 1'b0, 1'b0, n[939], 1'b0, 1'b0, 
        n[936:934], 1'b0, 1'b0, n[931], 1'b0, 1'b0, n[928:927], 1'b0, 1'b0, 
        n[924], 1'b0, 1'b0, n[921:918], 1'b0, 1'b0, n[915], 1'b0, 1'b0, 
        n[912:911], 1'b0, 1'b0, n[908], 1'b0, 1'b0, n[905:903], 1'b0, 1'b0, 
        n[900], 1'b0, 1'b0, n[897:896], 1'b0, 1'b0, n[893], 1'b0, 1'b0, 
        n[890:885], 1'b0, 1'b0, n[882], 1'b0, 1'b0, n[879:878], 1'b0, 1'b0, 
        n[875], 1'b0, 1'b0, n[872:870], 1'b0, 1'b0, n[867], 1'b0, 1'b0, 
        n[864:863], 1'b0, 1'b0, n[860], 1'b0, 1'b0, n[857:854], 1'b0, 1'b0, 
        n[851], 1'b0, 1'b0, n[848:847], 1'b0, 1'b0, n[844], 1'b0, 1'b0, 
        n[841:839], 1'b0, 1'b0, n[836], 1'b0, 1'b0, n[833:832], 1'b0, 1'b0, 
        n[829], 1'b0, 1'b0, n[826:822], 1'b0, 1'b0, n[819], 1'b0, 1'b0, 
        n[816:815], 1'b0, 1'b0, n[812], 1'b0, 1'b0, n[809:807], 1'b0, 1'b0, 
        n[804], 1'b0, 1'b0, n[801:800], 1'b0, 1'b0, n[797], 1'b0, 1'b0, 
        n[794:791], 1'b0, 1'b0, n[788], 1'b0, 1'b0, n[785:784], 1'b0, 1'b0, 
        n[781], 1'b0, 1'b0, n[778:776], 1'b0, 1'b0, n[773], 1'b0, 1'b0, 
        n[770:769], 1'b0, 1'b0, n[766], 1'b0, 1'b0, n[763:757], 1'b0, 1'b0, 
        n[754], 1'b0, 1'b0, n[751:750], 1'b0, 1'b0, n[747], 1'b0, 1'b0, 
        n[744:742], 1'b0, 1'b0, n[739], 1'b0, 1'b0, n[736:735], 1'b0, 1'b0, 
        n[732], 1'b0, 1'b0, n[729:726], 1'b0, 1'b0, n[723], 1'b0, 1'b0, 
        n[720:719], 1'b0, 1'b0, n[716], 1'b0, 1'b0, n[713:711], 1'b0, 1'b0, 
        n[708], 1'b0, 1'b0, n[705:704], 1'b0, 1'b0, n[701], 1'b0, 1'b0, 
        n[698:694], 1'b0, 1'b0, n[691], 1'b0, 1'b0, n[688:687], 1'b0, 1'b0, 
        n[684], 1'b0, 1'b0, n[681:679], 1'b0, 1'b0, n[676], 1'b0, 1'b0, 
        n[673:672], 1'b0, 1'b0, n[669], 1'b0, 1'b0, n[666:663], 1'b0, 1'b0, 
        n[660], 1'b0, 1'b0, n[657:656], 1'b0, 1'b0, n[653], 1'b0, 1'b0, 
        n[650:648], 1'b0, 1'b0, n[645], 1'b0, 1'b0, n[642:641], 1'b0, 1'b0, 
        n[638], 1'b0, 1'b0, n[635:630], 1'b0, 1'b0, n[627], 1'b0, 1'b0, 
        n[624:623], 1'b0, 1'b0, n[620], 1'b0, 1'b0, n[617:615], 1'b0, 1'b0, 
        n[612], 1'b0, 1'b0, n[609:608], 1'b0, 1'b0, n[605], 1'b0, 1'b0, 
        n[602:599], 1'b0, 1'b0, n[596], 1'b0, 1'b0, n[593:592], 1'b0, 1'b0, 
        n[589], 1'b0, 1'b0, n[586:584], 1'b0, 1'b0, n[581], 1'b0, 1'b0, 
        n[578:577], 1'b0, 1'b0, n[574], 1'b0, 1'b0, n[571:567], 1'b0, 1'b0, 
        n[564], 1'b0, 1'b0, n[561:560], 1'b0, 1'b0, n[557], 1'b0, 1'b0, 
        n[554:552], 1'b0, 1'b0, n[549], 1'b0, 1'b0, n[546:545], 1'b0, 1'b0, 
        n[542], 1'b0, 1'b0, n[539:536], 1'b0, 1'b0, n[533], 1'b0, 1'b0, 
        n[530:529], 1'b0, 1'b0, n[526], 1'b0, 1'b0, n[523:521], 1'b0, 1'b0, 
        n[518], 1'b0, 1'b0, n[515:514], 1'b0, 1'b0, n[511], 1'b0, 1'b0, 
        n[508:501], 1'b0, 1'b0, n[498], 1'b0, 1'b0, n[495:494], 1'b0, 1'b0, 
        n[491], 1'b0, 1'b0, n[488:486], 1'b0, 1'b0, n[483], 1'b0, 1'b0, 
        n[480:479], 1'b0, 1'b0, n[476], 1'b0, 1'b0, n[473:470], 1'b0, 1'b0, 
        n[467], 1'b0, 1'b0, n[464:463], 1'b0, 1'b0, n[460], 1'b0, 1'b0, 
        n[457:455], 1'b0, 1'b0, n[452], 1'b0, 1'b0, n[449:448], 1'b0, 1'b0, 
        n[445], 1'b0, 1'b0, n[442:438], 1'b0, 1'b0, n[435], 1'b0, 1'b0, 
        n[432:431], 1'b0, 1'b0, n[428], 1'b0, 1'b0, n[425:423], 1'b0, 1'b0, 
        n[420], 1'b0, 1'b0, n[417:416], 1'b0, 1'b0, n[413], 1'b0, 1'b0, 
        n[410:407], 1'b0, 1'b0, n[404], 1'b0, 1'b0, n[401:400], 1'b0, 1'b0, 
        n[397], 1'b0, 1'b0, n[394:392], 1'b0, 1'b0, n[389], 1'b0, 1'b0, 
        n[386:385], 1'b0, 1'b0, n[382], 1'b0, 1'b0, n[379:374], 1'b0, 1'b0, 
        n[371], 1'b0, 1'b0, n[368:367], 1'b0, 1'b0, n[364], 1'b0, 1'b0, 
        n[361:359], 1'b0, 1'b0, n[356], 1'b0, 1'b0, n[353:352], 1'b0, 1'b0, 
        n[349], 1'b0, 1'b0, n[346:343], 1'b0, 1'b0, n[340], 1'b0, 1'b0, 
        n[337:336], 1'b0, 1'b0, n[333], 1'b0, 1'b0, n[330:328], 1'b0, 1'b0, 
        n[325], 1'b0, 1'b0, n[322:321], 1'b0, 1'b0, n[318], 1'b0, 1'b0, 
        n[315:311], 1'b0, 1'b0, n[308], 1'b0, 1'b0, n[305:304], 1'b0, 1'b0, 
        n[301], 1'b0, 1'b0, n[298:296], 1'b0, 1'b0, n[293], 1'b0, 1'b0, 
        n[290:289], 1'b0, 1'b0, n[286], 1'b0, 1'b0, n[283:280], 1'b0, 1'b0, 
        n[277], 1'b0, 1'b0, n[274:273], 1'b0, 1'b0, n[270], 1'b0, 1'b0, 
        n[267:265], 1'b0, 1'b0, n[262], 1'b0, 1'b0, n[259:258], 1'b0, 1'b0, 
        n[255], 1'b0, 1'b0, n[252:246], 1'b0, 1'b0, n[243], 1'b0, 1'b0, 
        n[240:239], 1'b0, 1'b0, n[236], 1'b0, 1'b0, n[233:231], 1'b0, 1'b0, 
        n[228], 1'b0, 1'b0, n[225:224], 1'b0, 1'b0, n[221], 1'b0, 1'b0, 
        n[218:215], 1'b0, 1'b0, n[212], 1'b0, 1'b0, n[209:208], 1'b0, 1'b0, 
        n[205], 1'b0, 1'b0, n[202:200], 1'b0, 1'b0, n[197], 1'b0, 1'b0, 
        n[194:193], 1'b0, 1'b0, n[190], 1'b0, 1'b0, n[187:183], 1'b0, 1'b0, 
        n[180], 1'b0, 1'b0, n[177:176], 1'b0, 1'b0, n[173], 1'b0, 1'b0, 
        n[170:168], 1'b0, 1'b0, n[165], 1'b0, 1'b0, n[162:161], 1'b0, 1'b0, 
        n[158], 1'b0, 1'b0, n[155:152], 1'b0, 1'b0, n[149], 1'b0, 1'b0, 
        n[146:145], 1'b0, 1'b0, n[142], 1'b0, 1'b0, n[139:137], 1'b0, 1'b0, 
        n[134], 1'b0, 1'b0, n[131:130], 1'b0, 1'b0, n[127], 1'b0, 1'b0, 
        n[124:119], 1'b0, 1'b0, n[116], 1'b0, 1'b0, n[113:112], 1'b0, 1'b0, 
        n[109], 1'b0, 1'b0, n[106:104], 1'b0, 1'b0, n[101], 1'b0, 1'b0, 
        n[98:97], 1'b0, 1'b0, n[94], 1'b0, 1'b0, n[91:88], 1'b0, 1'b0, n[85], 
        1'b0, 1'b0, n[82:81], 1'b0, 1'b0, n[78], 1'b0, 1'b0, n[75:73], 1'b0, 
        1'b0, n[70], 1'b0, 1'b0, n[67:66], 1'b0, 1'b0, n[63], 1'b0, 1'b0, 
        n[60:56], 1'b0, 1'b0, n[53], 1'b0, 1'b0, n[50:49], 1'b0, 1'b0, n[46], 
        1'b0, 1'b0, n[43:41], 1'b0, 1'b0, n[38], 1'b0, 1'b0, n[35:34], 1'b0, 
        1'b0, n[31], 1'b0, 1'b0, n[28:25], 1'b0, 1'b0, n[22], 1'b0, 1'b0, 
        n[19:18], 1'b0, 1'b0, n[15], 1'b0, 1'b0, n[12:10], 1'b0, 1'b0, n[7], 
        1'b0, 1'b0, n[4:3], 1'b0, 1'b0, n[0]}), .s(s) );
endmodule

