module gen_nonlinear_part(a,b,n);
input  [7:0] a, b; //adder inputs
output [500:0] n; // non-linear outputs

wire [501:0] g;

assign g[0] = 0;
//Assigning outputs for input bit 0
assign g[1] = a[0] & b[0];
assign g[2] = a[0] & g[0];
assign g[3] = b[0] & g[0];
//Assigning outputs for input bit 1
assign g[4] = a[1] & b[1];
assign g[5] = a[1] & g[1];
assign g[8] = b[1] & g[1];
assign g[6] = a[1] & g[2];
assign g[9] = b[1] & g[2];
assign g[7] = a[1] & g[3];
assign g[10] = b[1] & g[3];
//Assigning outputs for input bit 2
assign g[11] = a[2] & b[2];
assign g[12] = a[2] & g[4];
assign g[19] = b[2] & g[4];
assign g[13] = a[2] & g[5];
assign g[20] = b[2] & g[5];
assign g[14] = a[2] & g[6];
assign g[21] = b[2] & g[6];
assign g[15] = a[2] & g[7];
assign g[22] = b[2] & g[7];
assign g[16] = a[2] & g[8];
assign g[23] = b[2] & g[8];
assign g[17] = a[2] & g[9];
assign g[24] = b[2] & g[9];
assign g[18] = a[2] & g[10];
assign g[25] = b[2] & g[10];
//Assigning outputs for input bit 3
assign g[26] = a[3] & b[3];
assign g[27] = a[3] & g[11];
assign g[42] = b[3] & g[11];
assign g[28] = a[3] & g[12];
assign g[43] = b[3] & g[12];
assign g[29] = a[3] & g[13];
assign g[44] = b[3] & g[13];
assign g[30] = a[3] & g[14];
assign g[45] = b[3] & g[14];
assign g[31] = a[3] & g[15];
assign g[46] = b[3] & g[15];
assign g[32] = a[3] & g[16];
assign g[47] = b[3] & g[16];
assign g[33] = a[3] & g[17];
assign g[48] = b[3] & g[17];
assign g[34] = a[3] & g[18];
assign g[49] = b[3] & g[18];
assign g[35] = a[3] & g[19];
assign g[50] = b[3] & g[19];
assign g[36] = a[3] & g[20];
assign g[51] = b[3] & g[20];
assign g[37] = a[3] & g[21];
assign g[52] = b[3] & g[21];
assign g[38] = a[3] & g[22];
assign g[53] = b[3] & g[22];
assign g[39] = a[3] & g[23];
assign g[54] = b[3] & g[23];
assign g[40] = a[3] & g[24];
assign g[55] = b[3] & g[24];
assign g[41] = a[3] & g[25];
assign g[56] = b[3] & g[25];
//Assigning outputs for input bit 4
assign g[57] = a[4] & b[4];
assign g[58] = a[4] & g[26];
assign g[89] = b[4] & g[26];
assign g[59] = a[4] & g[27];
assign g[90] = b[4] & g[27];
assign g[60] = a[4] & g[28];
assign g[91] = b[4] & g[28];
assign g[61] = a[4] & g[29];
assign g[92] = b[4] & g[29];
assign g[62] = a[4] & g[30];
assign g[93] = b[4] & g[30];
assign g[63] = a[4] & g[31];
assign g[94] = b[4] & g[31];
assign g[64] = a[4] & g[32];
assign g[95] = b[4] & g[32];
assign g[65] = a[4] & g[33];
assign g[96] = b[4] & g[33];
assign g[66] = a[4] & g[34];
assign g[97] = b[4] & g[34];
assign g[67] = a[4] & g[35];
assign g[98] = b[4] & g[35];
assign g[68] = a[4] & g[36];
assign g[99] = b[4] & g[36];
assign g[69] = a[4] & g[37];
assign g[100] = b[4] & g[37];
assign g[70] = a[4] & g[38];
assign g[101] = b[4] & g[38];
assign g[71] = a[4] & g[39];
assign g[102] = b[4] & g[39];
assign g[72] = a[4] & g[40];
assign g[103] = b[4] & g[40];
assign g[73] = a[4] & g[41];
assign g[104] = b[4] & g[41];
assign g[74] = a[4] & g[42];
assign g[105] = b[4] & g[42];
assign g[75] = a[4] & g[43];
assign g[106] = b[4] & g[43];
assign g[76] = a[4] & g[44];
assign g[107] = b[4] & g[44];
assign g[77] = a[4] & g[45];
assign g[108] = b[4] & g[45];
assign g[78] = a[4] & g[46];
assign g[109] = b[4] & g[46];
assign g[79] = a[4] & g[47];
assign g[110] = b[4] & g[47];
assign g[80] = a[4] & g[48];
assign g[111] = b[4] & g[48];
assign g[81] = a[4] & g[49];
assign g[112] = b[4] & g[49];
assign g[82] = a[4] & g[50];
assign g[113] = b[4] & g[50];
assign g[83] = a[4] & g[51];
assign g[114] = b[4] & g[51];
assign g[84] = a[4] & g[52];
assign g[115] = b[4] & g[52];
assign g[85] = a[4] & g[53];
assign g[116] = b[4] & g[53];
assign g[86] = a[4] & g[54];
assign g[117] = b[4] & g[54];
assign g[87] = a[4] & g[55];
assign g[118] = b[4] & g[55];
assign g[88] = a[4] & g[56];
assign g[119] = b[4] & g[56];
//Assigning outputs for input bit 5
assign g[120] = a[5] & b[5];
assign g[121] = a[5] & g[57];
assign g[184] = b[5] & g[57];
assign g[122] = a[5] & g[58];
assign g[185] = b[5] & g[58];
assign g[123] = a[5] & g[59];
assign g[186] = b[5] & g[59];
assign g[124] = a[5] & g[60];
assign g[187] = b[5] & g[60];
assign g[125] = a[5] & g[61];
assign g[188] = b[5] & g[61];
assign g[126] = a[5] & g[62];
assign g[189] = b[5] & g[62];
assign g[127] = a[5] & g[63];
assign g[190] = b[5] & g[63];
assign g[128] = a[5] & g[64];
assign g[191] = b[5] & g[64];
assign g[129] = a[5] & g[65];
assign g[192] = b[5] & g[65];
assign g[130] = a[5] & g[66];
assign g[193] = b[5] & g[66];
assign g[131] = a[5] & g[67];
assign g[194] = b[5] & g[67];
assign g[132] = a[5] & g[68];
assign g[195] = b[5] & g[68];
assign g[133] = a[5] & g[69];
assign g[196] = b[5] & g[69];
assign g[134] = a[5] & g[70];
assign g[197] = b[5] & g[70];
assign g[135] = a[5] & g[71];
assign g[198] = b[5] & g[71];
assign g[136] = a[5] & g[72];
assign g[199] = b[5] & g[72];
assign g[137] = a[5] & g[73];
assign g[200] = b[5] & g[73];
assign g[138] = a[5] & g[74];
assign g[201] = b[5] & g[74];
assign g[139] = a[5] & g[75];
assign g[202] = b[5] & g[75];
assign g[140] = a[5] & g[76];
assign g[203] = b[5] & g[76];
assign g[141] = a[5] & g[77];
assign g[204] = b[5] & g[77];
assign g[142] = a[5] & g[78];
assign g[205] = b[5] & g[78];
assign g[143] = a[5] & g[79];
assign g[206] = b[5] & g[79];
assign g[144] = a[5] & g[80];
assign g[207] = b[5] & g[80];
assign g[145] = a[5] & g[81];
assign g[208] = b[5] & g[81];
assign g[146] = a[5] & g[82];
assign g[209] = b[5] & g[82];
assign g[147] = a[5] & g[83];
assign g[210] = b[5] & g[83];
assign g[148] = a[5] & g[84];
assign g[211] = b[5] & g[84];
assign g[149] = a[5] & g[85];
assign g[212] = b[5] & g[85];
assign g[150] = a[5] & g[86];
assign g[213] = b[5] & g[86];
assign g[151] = a[5] & g[87];
assign g[214] = b[5] & g[87];
assign g[152] = a[5] & g[88];
assign g[215] = b[5] & g[88];
assign g[153] = a[5] & g[89];
assign g[216] = b[5] & g[89];
assign g[154] = a[5] & g[90];
assign g[217] = b[5] & g[90];
assign g[155] = a[5] & g[91];
assign g[218] = b[5] & g[91];
assign g[156] = a[5] & g[92];
assign g[219] = b[5] & g[92];
assign g[157] = a[5] & g[93];
assign g[220] = b[5] & g[93];
assign g[158] = a[5] & g[94];
assign g[221] = b[5] & g[94];
assign g[159] = a[5] & g[95];
assign g[222] = b[5] & g[95];
assign g[160] = a[5] & g[96];
assign g[223] = b[5] & g[96];
assign g[161] = a[5] & g[97];
assign g[224] = b[5] & g[97];
assign g[162] = a[5] & g[98];
assign g[225] = b[5] & g[98];
assign g[163] = a[5] & g[99];
assign g[226] = b[5] & g[99];
assign g[164] = a[5] & g[100];
assign g[227] = b[5] & g[100];
assign g[165] = a[5] & g[101];
assign g[228] = b[5] & g[101];
assign g[166] = a[5] & g[102];
assign g[229] = b[5] & g[102];
assign g[167] = a[5] & g[103];
assign g[230] = b[5] & g[103];
assign g[168] = a[5] & g[104];
assign g[231] = b[5] & g[104];
assign g[169] = a[5] & g[105];
assign g[232] = b[5] & g[105];
assign g[170] = a[5] & g[106];
assign g[233] = b[5] & g[106];
assign g[171] = a[5] & g[107];
assign g[234] = b[5] & g[107];
assign g[172] = a[5] & g[108];
assign g[235] = b[5] & g[108];
assign g[173] = a[5] & g[109];
assign g[236] = b[5] & g[109];
assign g[174] = a[5] & g[110];
assign g[237] = b[5] & g[110];
assign g[175] = a[5] & g[111];
assign g[238] = b[5] & g[111];
assign g[176] = a[5] & g[112];
assign g[239] = b[5] & g[112];
assign g[177] = a[5] & g[113];
assign g[240] = b[5] & g[113];
assign g[178] = a[5] & g[114];
assign g[241] = b[5] & g[114];
assign g[179] = a[5] & g[115];
assign g[242] = b[5] & g[115];
assign g[180] = a[5] & g[116];
assign g[243] = b[5] & g[116];
assign g[181] = a[5] & g[117];
assign g[244] = b[5] & g[117];
assign g[182] = a[5] & g[118];
assign g[245] = b[5] & g[118];
assign g[183] = a[5] & g[119];
assign g[246] = b[5] & g[119];
//Assigning outputs for input bit 6
assign g[247] = a[6] & b[6];
assign g[248] = a[6] & g[120];
assign g[375] = b[6] & g[120];
assign g[249] = a[6] & g[121];
assign g[376] = b[6] & g[121];
assign g[250] = a[6] & g[122];
assign g[377] = b[6] & g[122];
assign g[251] = a[6] & g[123];
assign g[378] = b[6] & g[123];
assign g[252] = a[6] & g[124];
assign g[379] = b[6] & g[124];
assign g[253] = a[6] & g[125];
assign g[380] = b[6] & g[125];
assign g[254] = a[6] & g[126];
assign g[381] = b[6] & g[126];
assign g[255] = a[6] & g[127];
assign g[382] = b[6] & g[127];
assign g[256] = a[6] & g[128];
assign g[383] = b[6] & g[128];
assign g[257] = a[6] & g[129];
assign g[384] = b[6] & g[129];
assign g[258] = a[6] & g[130];
assign g[385] = b[6] & g[130];
assign g[259] = a[6] & g[131];
assign g[386] = b[6] & g[131];
assign g[260] = a[6] & g[132];
assign g[387] = b[6] & g[132];
assign g[261] = a[6] & g[133];
assign g[388] = b[6] & g[133];
assign g[262] = a[6] & g[134];
assign g[389] = b[6] & g[134];
assign g[263] = a[6] & g[135];
assign g[390] = b[6] & g[135];
assign g[264] = a[6] & g[136];
assign g[391] = b[6] & g[136];
assign g[265] = a[6] & g[137];
assign g[392] = b[6] & g[137];
assign g[266] = a[6] & g[138];
assign g[393] = b[6] & g[138];
assign g[267] = a[6] & g[139];
assign g[394] = b[6] & g[139];
assign g[268] = a[6] & g[140];
assign g[395] = b[6] & g[140];
assign g[269] = a[6] & g[141];
assign g[396] = b[6] & g[141];
assign g[270] = a[6] & g[142];
assign g[397] = b[6] & g[142];
assign g[271] = a[6] & g[143];
assign g[398] = b[6] & g[143];
assign g[272] = a[6] & g[144];
assign g[399] = b[6] & g[144];
assign g[273] = a[6] & g[145];
assign g[400] = b[6] & g[145];
assign g[274] = a[6] & g[146];
assign g[401] = b[6] & g[146];
assign g[275] = a[6] & g[147];
assign g[402] = b[6] & g[147];
assign g[276] = a[6] & g[148];
assign g[403] = b[6] & g[148];
assign g[277] = a[6] & g[149];
assign g[404] = b[6] & g[149];
assign g[278] = a[6] & g[150];
assign g[405] = b[6] & g[150];
assign g[279] = a[6] & g[151];
assign g[406] = b[6] & g[151];
assign g[280] = a[6] & g[152];
assign g[407] = b[6] & g[152];
assign g[281] = a[6] & g[153];
assign g[408] = b[6] & g[153];
assign g[282] = a[6] & g[154];
assign g[409] = b[6] & g[154];
assign g[283] = a[6] & g[155];
assign g[410] = b[6] & g[155];
assign g[284] = a[6] & g[156];
assign g[411] = b[6] & g[156];
assign g[285] = a[6] & g[157];
assign g[412] = b[6] & g[157];
assign g[286] = a[6] & g[158];
assign g[413] = b[6] & g[158];
assign g[287] = a[6] & g[159];
assign g[414] = b[6] & g[159];
assign g[288] = a[6] & g[160];
assign g[415] = b[6] & g[160];
assign g[289] = a[6] & g[161];
assign g[416] = b[6] & g[161];
assign g[290] = a[6] & g[162];
assign g[417] = b[6] & g[162];
assign g[291] = a[6] & g[163];
assign g[418] = b[6] & g[163];
assign g[292] = a[6] & g[164];
assign g[419] = b[6] & g[164];
assign g[293] = a[6] & g[165];
assign g[420] = b[6] & g[165];
assign g[294] = a[6] & g[166];
assign g[421] = b[6] & g[166];
assign g[295] = a[6] & g[167];
assign g[422] = b[6] & g[167];
assign g[296] = a[6] & g[168];
assign g[423] = b[6] & g[168];
assign g[297] = a[6] & g[169];
assign g[424] = b[6] & g[169];
assign g[298] = a[6] & g[170];
assign g[425] = b[6] & g[170];
assign g[299] = a[6] & g[171];
assign g[426] = b[6] & g[171];
assign g[300] = a[6] & g[172];
assign g[427] = b[6] & g[172];
assign g[301] = a[6] & g[173];
assign g[428] = b[6] & g[173];
assign g[302] = a[6] & g[174];
assign g[429] = b[6] & g[174];
assign g[303] = a[6] & g[175];
assign g[430] = b[6] & g[175];
assign g[304] = a[6] & g[176];
assign g[431] = b[6] & g[176];
assign g[305] = a[6] & g[177];
assign g[432] = b[6] & g[177];
assign g[306] = a[6] & g[178];
assign g[433] = b[6] & g[178];
assign g[307] = a[6] & g[179];
assign g[434] = b[6] & g[179];
assign g[308] = a[6] & g[180];
assign g[435] = b[6] & g[180];
assign g[309] = a[6] & g[181];
assign g[436] = b[6] & g[181];
assign g[310] = a[6] & g[182];
assign g[437] = b[6] & g[182];
assign g[311] = a[6] & g[183];
assign g[438] = b[6] & g[183];
assign g[312] = a[6] & g[184];
assign g[439] = b[6] & g[184];
assign g[313] = a[6] & g[185];
assign g[440] = b[6] & g[185];
assign g[314] = a[6] & g[186];
assign g[441] = b[6] & g[186];
assign g[315] = a[6] & g[187];
assign g[442] = b[6] & g[187];
assign g[316] = a[6] & g[188];
assign g[443] = b[6] & g[188];
assign g[317] = a[6] & g[189];
assign g[444] = b[6] & g[189];
assign g[318] = a[6] & g[190];
assign g[445] = b[6] & g[190];
assign g[319] = a[6] & g[191];
assign g[446] = b[6] & g[191];
assign g[320] = a[6] & g[192];
assign g[447] = b[6] & g[192];
assign g[321] = a[6] & g[193];
assign g[448] = b[6] & g[193];
assign g[322] = a[6] & g[194];
assign g[449] = b[6] & g[194];
assign g[323] = a[6] & g[195];
assign g[450] = b[6] & g[195];
assign g[324] = a[6] & g[196];
assign g[451] = b[6] & g[196];
assign g[325] = a[6] & g[197];
assign g[452] = b[6] & g[197];
assign g[326] = a[6] & g[198];
assign g[453] = b[6] & g[198];
assign g[327] = a[6] & g[199];
assign g[454] = b[6] & g[199];
assign g[328] = a[6] & g[200];
assign g[455] = b[6] & g[200];
assign g[329] = a[6] & g[201];
assign g[456] = b[6] & g[201];
assign g[330] = a[6] & g[202];
assign g[457] = b[6] & g[202];
assign g[331] = a[6] & g[203];
assign g[458] = b[6] & g[203];
assign g[332] = a[6] & g[204];
assign g[459] = b[6] & g[204];
assign g[333] = a[6] & g[205];
assign g[460] = b[6] & g[205];
assign g[334] = a[6] & g[206];
assign g[461] = b[6] & g[206];
assign g[335] = a[6] & g[207];
assign g[462] = b[6] & g[207];
assign g[336] = a[6] & g[208];
assign g[463] = b[6] & g[208];
assign g[337] = a[6] & g[209];
assign g[464] = b[6] & g[209];
assign g[338] = a[6] & g[210];
assign g[465] = b[6] & g[210];
assign g[339] = a[6] & g[211];
assign g[466] = b[6] & g[211];
assign g[340] = a[6] & g[212];
assign g[467] = b[6] & g[212];
assign g[341] = a[6] & g[213];
assign g[468] = b[6] & g[213];
assign g[342] = a[6] & g[214];
assign g[469] = b[6] & g[214];
assign g[343] = a[6] & g[215];
assign g[470] = b[6] & g[215];
assign g[344] = a[6] & g[216];
assign g[471] = b[6] & g[216];
assign g[345] = a[6] & g[217];
assign g[472] = b[6] & g[217];
assign g[346] = a[6] & g[218];
assign g[473] = b[6] & g[218];
assign g[347] = a[6] & g[219];
assign g[474] = b[6] & g[219];
assign g[348] = a[6] & g[220];
assign g[475] = b[6] & g[220];
assign g[349] = a[6] & g[221];
assign g[476] = b[6] & g[221];
assign g[350] = a[6] & g[222];
assign g[477] = b[6] & g[222];
assign g[351] = a[6] & g[223];
assign g[478] = b[6] & g[223];
assign g[352] = a[6] & g[224];
assign g[479] = b[6] & g[224];
assign g[353] = a[6] & g[225];
assign g[480] = b[6] & g[225];
assign g[354] = a[6] & g[226];
assign g[481] = b[6] & g[226];
assign g[355] = a[6] & g[227];
assign g[482] = b[6] & g[227];
assign g[356] = a[6] & g[228];
assign g[483] = b[6] & g[228];
assign g[357] = a[6] & g[229];
assign g[484] = b[6] & g[229];
assign g[358] = a[6] & g[230];
assign g[485] = b[6] & g[230];
assign g[359] = a[6] & g[231];
assign g[486] = b[6] & g[231];
assign g[360] = a[6] & g[232];
assign g[487] = b[6] & g[232];
assign g[361] = a[6] & g[233];
assign g[488] = b[6] & g[233];
assign g[362] = a[6] & g[234];
assign g[489] = b[6] & g[234];
assign g[363] = a[6] & g[235];
assign g[490] = b[6] & g[235];
assign g[364] = a[6] & g[236];
assign g[491] = b[6] & g[236];
assign g[365] = a[6] & g[237];
assign g[492] = b[6] & g[237];
assign g[366] = a[6] & g[238];
assign g[493] = b[6] & g[238];
assign g[367] = a[6] & g[239];
assign g[494] = b[6] & g[239];
assign g[368] = a[6] & g[240];
assign g[495] = b[6] & g[240];
assign g[369] = a[6] & g[241];
assign g[496] = b[6] & g[241];
assign g[370] = a[6] & g[242];
assign g[497] = b[6] & g[242];
assign g[371] = a[6] & g[243];
assign g[498] = b[6] & g[243];
assign g[372] = a[6] & g[244];
assign g[499] = b[6] & g[244];
assign g[373] = a[6] & g[245];
assign g[500] = b[6] & g[245];
assign g[374] = a[6] & g[246];
assign g[501] = b[6] & g[246];
assign n = g[501:1]; //assign outputs
endmodule