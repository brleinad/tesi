module dec_lut (enc_s,dec_s);
`include "constants.v"

input [NBIT:0]  enc_s;
output reg [NBIT:0]  dec_s;
always @(*)
begin
    case(enc_s)
	0 : dec_s = 0;
	256 : dec_s = 1;
	128 : dec_s = 2;
	384 : dec_s = 3;
	64 : dec_s = 4;
	320 : dec_s = 5;
	288 : dec_s = 6;
	448 : dec_s = 7;
	32 : dec_s = 8;
	272 : dec_s = 9;
	264 : dec_s = 10;
	416 : dec_s = 11;
	260 : dec_s = 12;
	400 : dec_s = 13;
	392 : dec_s = 14;
	480 : dec_s = 15;
	8 : dec_s = 16;
	258 : dec_s = 17;
	257 : dec_s = 18;
	388 : dec_s = 19;
	192 : dec_s = 20;
	386 : dec_s = 21;
	385 : dec_s = 22;
	464 : dec_s = 23;
	160 : dec_s = 24;
	352 : dec_s = 25;
	336 : dec_s = 26;
	456 : dec_s = 27;
	328 : dec_s = 28;
	452 : dec_s = 29;
	450 : dec_s = 30;
	496 : dec_s = 31;
	16 : dec_s = 32;
	144 : dec_s = 33;
	136 : dec_s = 34;
	324 : dec_s = 35;
	132 : dec_s = 36;
	322 : dec_s = 37;
	321 : dec_s = 38;
	449 : dec_s = 39;
	130 : dec_s = 40;
	304 : dec_s = 41;
	296 : dec_s = 42;
	432 : dec_s = 43;
	292 : dec_s = 44;
	424 : dec_s = 45;
	420 : dec_s = 46;
	488 : dec_s = 47;
	129 : dec_s = 48;
	290 : dec_s = 49;
	289 : dec_s = 50;
	418 : dec_s = 51;
	280 : dec_s = 52;
	417 : dec_s = 53;
	408 : dec_s = 54;
	484 : dec_s = 55;
	276 : dec_s = 56;
	404 : dec_s = 57;
	402 : dec_s = 58;
	482 : dec_s = 59;
	401 : dec_s = 60;
	481 : dec_s = 61;
	472 : dec_s = 62;
	504 : dec_s = 63;
	4 : dec_s = 64;
	96 : dec_s = 65;
	80 : dec_s = 66;
	274 : dec_s = 67;
	72 : dec_s = 68;
	273 : dec_s = 69;
	268 : dec_s = 70;
	396 : dec_s = 71;
	68 : dec_s = 72;
	266 : dec_s = 73;
	265 : dec_s = 74;
	394 : dec_s = 75;
	262 : dec_s = 76;
	393 : dec_s = 77;
	390 : dec_s = 78;
	468 : dec_s = 79;
	66 : dec_s = 80;
	261 : dec_s = 81;
	259 : dec_s = 82;
	389 : dec_s = 83;
	224 : dec_s = 84;
	387 : dec_s = 85;
	368 : dec_s = 86;
	466 : dec_s = 87;
	208 : dec_s = 88;
	360 : dec_s = 89;
	356 : dec_s = 90;
	465 : dec_s = 91;
	354 : dec_s = 92;
	460 : dec_s = 93;
	458 : dec_s = 94;
	500 : dec_s = 95;
	65 : dec_s = 96;
	200 : dec_s = 97;
	196 : dec_s = 98;
	353 : dec_s = 99;
	194 : dec_s = 100;
	344 : dec_s = 101;
	340 : dec_s = 102;
	457 : dec_s = 103;
	193 : dec_s = 104;
	338 : dec_s = 105;
	337 : dec_s = 106;
	454 : dec_s = 107;
	332 : dec_s = 108;
	453 : dec_s = 109;
	451 : dec_s = 110;
	498 : dec_s = 111;
	176 : dec_s = 112;
	330 : dec_s = 113;
	329 : dec_s = 114;
	440 : dec_s = 115;
	326 : dec_s = 116;
	436 : dec_s = 117;
	434 : dec_s = 118;
	497 : dec_s = 119;
	325 : dec_s = 120;
	433 : dec_s = 121;
	428 : dec_s = 122;
	492 : dec_s = 123;
	426 : dec_s = 124;
	490 : dec_s = 125;
	489 : dec_s = 126;
	508 : dec_s = 127;
	2 : dec_s = 128;
	48 : dec_s = 129;
	40 : dec_s = 130;
	168 : dec_s = 131;
	36 : dec_s = 132;
	164 : dec_s = 133;
	162 : dec_s = 134;
	323 : dec_s = 135;
	34 : dec_s = 136;
	161 : dec_s = 137;
	152 : dec_s = 138;
	312 : dec_s = 139;
	148 : dec_s = 140;
	308 : dec_s = 141;
	306 : dec_s = 142;
	425 : dec_s = 143;
	33 : dec_s = 144;
	146 : dec_s = 145;
	145 : dec_s = 146;
	305 : dec_s = 147;
	140 : dec_s = 148;
	300 : dec_s = 149;
	298 : dec_s = 150;
	422 : dec_s = 151;
	138 : dec_s = 152;
	297 : dec_s = 153;
	294 : dec_s = 154;
	421 : dec_s = 155;
	293 : dec_s = 156;
	419 : dec_s = 157;
	412 : dec_s = 158;
	486 : dec_s = 159;
	24 : dec_s = 160;
	137 : dec_s = 161;
	134 : dec_s = 162;
	291 : dec_s = 163;
	133 : dec_s = 164;
	284 : dec_s = 165;
	282 : dec_s = 166;
	410 : dec_s = 167;
	131 : dec_s = 168;
	281 : dec_s = 169;
	278 : dec_s = 170;
	409 : dec_s = 171;
	277 : dec_s = 172;
	406 : dec_s = 173;
	405 : dec_s = 174;
	485 : dec_s = 175;
	112 : dec_s = 176;
	275 : dec_s = 177;
	270 : dec_s = 178;
	403 : dec_s = 179;
	269 : dec_s = 180;
	398 : dec_s = 181;
	397 : dec_s = 182;
	483 : dec_s = 183;
	267 : dec_s = 184;
	395 : dec_s = 185;
	391 : dec_s = 186;
	476 : dec_s = 187;
	376 : dec_s = 188;
	474 : dec_s = 189;
	473 : dec_s = 190;
	506 : dec_s = 191;
	20 : dec_s = 192;
	104 : dec_s = 193;
	100 : dec_s = 194;
	263 : dec_s = 195;
	98 : dec_s = 196;
	240 : dec_s = 197;
	232 : dec_s = 198;
	372 : dec_s = 199;
	97 : dec_s = 200;
	228 : dec_s = 201;
	226 : dec_s = 202;
	370 : dec_s = 203;
	225 : dec_s = 204;
	369 : dec_s = 205;
	364 : dec_s = 206;
	470 : dec_s = 207;
	88 : dec_s = 208;
	216 : dec_s = 209;
	212 : dec_s = 210;
	362 : dec_s = 211;
	210 : dec_s = 212;
	361 : dec_s = 213;
	358 : dec_s = 214;
	469 : dec_s = 215;
	209 : dec_s = 216;
	357 : dec_s = 217;
	355 : dec_s = 218;
	467 : dec_s = 219;
	348 : dec_s = 220;
	462 : dec_s = 221;
	461 : dec_s = 222;
	505 : dec_s = 223;
	84 : dec_s = 224;
	204 : dec_s = 225;
	202 : dec_s = 226;
	346 : dec_s = 227;
	201 : dec_s = 228;
	345 : dec_s = 229;
	342 : dec_s = 230;
	459 : dec_s = 231;
	198 : dec_s = 232;
	341 : dec_s = 233;
	339 : dec_s = 234;
	455 : dec_s = 235;
	334 : dec_s = 236;
	444 : dec_s = 237;
	442 : dec_s = 238;
	502 : dec_s = 239;
	197 : dec_s = 240;
	333 : dec_s = 241;
	331 : dec_s = 242;
	441 : dec_s = 243;
	327 : dec_s = 244;
	438 : dec_s = 245;
	437 : dec_s = 246;
	501 : dec_s = 247;
	316 : dec_s = 248;
	435 : dec_s = 249;
	430 : dec_s = 250;
	499 : dec_s = 251;
	429 : dec_s = 252;
	494 : dec_s = 253;
	493 : dec_s = 254;
	510 : dec_s = 255;
	1 : dec_s = 256;
	18 : dec_s = 257;
	17 : dec_s = 258;
	82 : dec_s = 259;
	12 : dec_s = 260;
	81 : dec_s = 261;
	76 : dec_s = 262;
	195 : dec_s = 263;
	10 : dec_s = 264;
	74 : dec_s = 265;
	73 : dec_s = 266;
	184 : dec_s = 267;
	70 : dec_s = 268;
	180 : dec_s = 269;
	178 : dec_s = 270;
	314 : dec_s = 271;
	9 : dec_s = 272;
	69 : dec_s = 273;
	67 : dec_s = 274;
	177 : dec_s = 275;
	56 : dec_s = 276;
	172 : dec_s = 277;
	170 : dec_s = 278;
	313 : dec_s = 279;
	52 : dec_s = 280;
	169 : dec_s = 281;
	166 : dec_s = 282;
	310 : dec_s = 283;
	165 : dec_s = 284;
	309 : dec_s = 285;
	307 : dec_s = 286;
	427 : dec_s = 287;
	6 : dec_s = 288;
	50 : dec_s = 289;
	49 : dec_s = 290;
	163 : dec_s = 291;
	44 : dec_s = 292;
	156 : dec_s = 293;
	154 : dec_s = 294;
	302 : dec_s = 295;
	42 : dec_s = 296;
	153 : dec_s = 297;
	150 : dec_s = 298;
	301 : dec_s = 299;
	149 : dec_s = 300;
	299 : dec_s = 301;
	295 : dec_s = 302;
	423 : dec_s = 303;
	41 : dec_s = 304;
	147 : dec_s = 305;
	142 : dec_s = 306;
	286 : dec_s = 307;
	141 : dec_s = 308;
	285 : dec_s = 309;
	283 : dec_s = 310;
	414 : dec_s = 311;
	139 : dec_s = 312;
	279 : dec_s = 313;
	271 : dec_s = 314;
	413 : dec_s = 315;
	248 : dec_s = 316;
	411 : dec_s = 317;
	407 : dec_s = 318;
	491 : dec_s = 319;
	5 : dec_s = 320;
	38 : dec_s = 321;
	37 : dec_s = 322;
	135 : dec_s = 323;
	35 : dec_s = 324;
	120 : dec_s = 325;
	116 : dec_s = 326;
	244 : dec_s = 327;
	28 : dec_s = 328;
	114 : dec_s = 329;
	113 : dec_s = 330;
	242 : dec_s = 331;
	108 : dec_s = 332;
	241 : dec_s = 333;
	236 : dec_s = 334;
	399 : dec_s = 335;
	26 : dec_s = 336;
	106 : dec_s = 337;
	105 : dec_s = 338;
	234 : dec_s = 339;
	102 : dec_s = 340;
	233 : dec_s = 341;
	230 : dec_s = 342;
	380 : dec_s = 343;
	101 : dec_s = 344;
	229 : dec_s = 345;
	227 : dec_s = 346;
	378 : dec_s = 347;
	220 : dec_s = 348;
	377 : dec_s = 349;
	374 : dec_s = 350;
	487 : dec_s = 351;
	25 : dec_s = 352;
	99 : dec_s = 353;
	92 : dec_s = 354;
	218 : dec_s = 355;
	90 : dec_s = 356;
	217 : dec_s = 357;
	214 : dec_s = 358;
	373 : dec_s = 359;
	89 : dec_s = 360;
	213 : dec_s = 361;
	211 : dec_s = 362;
	371 : dec_s = 363;
	206 : dec_s = 364;
	366 : dec_s = 365;
	365 : dec_s = 366;
	478 : dec_s = 367;
	86 : dec_s = 368;
	205 : dec_s = 369;
	203 : dec_s = 370;
	363 : dec_s = 371;
	199 : dec_s = 372;
	359 : dec_s = 373;
	350 : dec_s = 374;
	477 : dec_s = 375;
	188 : dec_s = 376;
	349 : dec_s = 377;
	347 : dec_s = 378;
	475 : dec_s = 379;
	343 : dec_s = 380;
	471 : dec_s = 381;
	463 : dec_s = 382;
	509 : dec_s = 383;
	3 : dec_s = 384;
	22 : dec_s = 385;
	21 : dec_s = 386;
	85 : dec_s = 387;
	19 : dec_s = 388;
	83 : dec_s = 389;
	78 : dec_s = 390;
	186 : dec_s = 391;
	14 : dec_s = 392;
	77 : dec_s = 393;
	75 : dec_s = 394;
	185 : dec_s = 395;
	71 : dec_s = 396;
	182 : dec_s = 397;
	181 : dec_s = 398;
	335 : dec_s = 399;
	13 : dec_s = 400;
	60 : dec_s = 401;
	58 : dec_s = 402;
	179 : dec_s = 403;
	57 : dec_s = 404;
	174 : dec_s = 405;
	173 : dec_s = 406;
	318 : dec_s = 407;
	54 : dec_s = 408;
	171 : dec_s = 409;
	167 : dec_s = 410;
	317 : dec_s = 411;
	158 : dec_s = 412;
	315 : dec_s = 413;
	311 : dec_s = 414;
	446 : dec_s = 415;
	11 : dec_s = 416;
	53 : dec_s = 417;
	51 : dec_s = 418;
	157 : dec_s = 419;
	46 : dec_s = 420;
	155 : dec_s = 421;
	151 : dec_s = 422;
	303 : dec_s = 423;
	45 : dec_s = 424;
	143 : dec_s = 425;
	124 : dec_s = 426;
	287 : dec_s = 427;
	122 : dec_s = 428;
	252 : dec_s = 429;
	250 : dec_s = 430;
	445 : dec_s = 431;
	43 : dec_s = 432;
	121 : dec_s = 433;
	118 : dec_s = 434;
	249 : dec_s = 435;
	117 : dec_s = 436;
	246 : dec_s = 437;
	245 : dec_s = 438;
	443 : dec_s = 439;
	115 : dec_s = 440;
	243 : dec_s = 441;
	238 : dec_s = 442;
	439 : dec_s = 443;
	237 : dec_s = 444;
	431 : dec_s = 445;
	415 : dec_s = 446;
	507 : dec_s = 447;
	7 : dec_s = 448;
	39 : dec_s = 449;
	30 : dec_s = 450;
	110 : dec_s = 451;
	29 : dec_s = 452;
	109 : dec_s = 453;
	107 : dec_s = 454;
	235 : dec_s = 455;
	27 : dec_s = 456;
	103 : dec_s = 457;
	94 : dec_s = 458;
	231 : dec_s = 459;
	93 : dec_s = 460;
	222 : dec_s = 461;
	221 : dec_s = 462;
	382 : dec_s = 463;
	23 : dec_s = 464;
	91 : dec_s = 465;
	87 : dec_s = 466;
	219 : dec_s = 467;
	79 : dec_s = 468;
	215 : dec_s = 469;
	207 : dec_s = 470;
	381 : dec_s = 471;
	62 : dec_s = 472;
	190 : dec_s = 473;
	189 : dec_s = 474;
	379 : dec_s = 475;
	187 : dec_s = 476;
	375 : dec_s = 477;
	367 : dec_s = 478;
	503 : dec_s = 479;
	15 : dec_s = 480;
	61 : dec_s = 481;
	59 : dec_s = 482;
	183 : dec_s = 483;
	55 : dec_s = 484;
	175 : dec_s = 485;
	159 : dec_s = 486;
	351 : dec_s = 487;
	47 : dec_s = 488;
	126 : dec_s = 489;
	125 : dec_s = 490;
	319 : dec_s = 491;
	123 : dec_s = 492;
	254 : dec_s = 493;
	253 : dec_s = 494;
	479 : dec_s = 495;
	31 : dec_s = 496;
	119 : dec_s = 497;
	111 : dec_s = 498;
	251 : dec_s = 499;
	95 : dec_s = 500;
	247 : dec_s = 501;
	239 : dec_s = 502;
	495 : dec_s = 503;
	63 : dec_s = 504;
	223 : dec_s = 505;
	191 : dec_s = 506;
	447 : dec_s = 507;
	127 : dec_s = 508;
	383 : dec_s = 509;
	255 : dec_s = 510;
	default : dec_s = 0;
    endcase
end
endmodule
