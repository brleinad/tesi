module gen_linear_part(a,b,n,s);

input  [15:0] a, b; //adder inputs
input [65518:0] n; // non-linear outputs
output [15:0] s;

wire [65518:0] t; // non-linear outputs
//asigning bit 0
assign s[0] = a[0] ^ b[0];
assign t[0] = n[0];

//asigning bit 1
assign s[1] = ( a[1] ^ b [1] ) ^ t[0];

assign t[1] = n[1];
assign t[2] = t[1] ^ n[2];
assign t[3] = t[2] ^ n[3];

//asigning bit 2
assign s[2] = ( a[2] ^ b [2] ) ^ t[3];

assign t[4] = n[4];
assign t[5] = t[4] ^ n[5];
assign t[6] = t[5] ^ n[6];
assign t[7] = t[6] ^ n[7];
assign t[8] = t[7] ^ n[8];
assign t[9] = t[8] ^ n[9];
assign t[10] = t[9] ^ n[10];

//asigning bit 3
assign s[3] = ( a[3] ^ b [3] ) ^ t[10];

assign t[11] = n[11];
assign t[12] = t[11] ^ n[12];
assign t[13] = t[12] ^ n[13];
assign t[14] = t[13] ^ n[14];
assign t[15] = t[14] ^ n[15];
assign t[16] = t[15] ^ n[16];
assign t[17] = t[16] ^ n[17];
assign t[18] = t[17] ^ n[18];
assign t[19] = t[18] ^ n[19];
assign t[20] = t[19] ^ n[20];
assign t[21] = t[20] ^ n[21];
assign t[22] = t[21] ^ n[22];
assign t[23] = t[22] ^ n[23];
assign t[24] = t[23] ^ n[24];
assign t[25] = t[24] ^ n[25];

//asigning bit 4
assign s[4] = ( a[4] ^ b [4] ) ^ t[25];

assign t[26] = n[26];
assign t[27] = t[26] ^ n[27];
assign t[28] = t[27] ^ n[28];
assign t[29] = t[28] ^ n[29];
assign t[30] = t[29] ^ n[30];
assign t[31] = t[30] ^ n[31];
assign t[32] = t[31] ^ n[32];
assign t[33] = t[32] ^ n[33];
assign t[34] = t[33] ^ n[34];
assign t[35] = t[34] ^ n[35];
assign t[36] = t[35] ^ n[36];
assign t[37] = t[36] ^ n[37];
assign t[38] = t[37] ^ n[38];
assign t[39] = t[38] ^ n[39];
assign t[40] = t[39] ^ n[40];
assign t[41] = t[40] ^ n[41];
assign t[42] = t[41] ^ n[42];
assign t[43] = t[42] ^ n[43];
assign t[44] = t[43] ^ n[44];
assign t[45] = t[44] ^ n[45];
assign t[46] = t[45] ^ n[46];
assign t[47] = t[46] ^ n[47];
assign t[48] = t[47] ^ n[48];
assign t[49] = t[48] ^ n[49];
assign t[50] = t[49] ^ n[50];
assign t[51] = t[50] ^ n[51];
assign t[52] = t[51] ^ n[52];
assign t[53] = t[52] ^ n[53];
assign t[54] = t[53] ^ n[54];
assign t[55] = t[54] ^ n[55];
assign t[56] = t[55] ^ n[56];

//asigning bit 5
assign s[5] = ( a[5] ^ b [5] ) ^ t[56];

assign t[57] = n[57];
assign t[58] = t[57] ^ n[58];
assign t[59] = t[58] ^ n[59];
assign t[60] = t[59] ^ n[60];
assign t[61] = t[60] ^ n[61];
assign t[62] = t[61] ^ n[62];
assign t[63] = t[62] ^ n[63];
assign t[64] = t[63] ^ n[64];
assign t[65] = t[64] ^ n[65];
assign t[66] = t[65] ^ n[66];
assign t[67] = t[66] ^ n[67];
assign t[68] = t[67] ^ n[68];
assign t[69] = t[68] ^ n[69];
assign t[70] = t[69] ^ n[70];
assign t[71] = t[70] ^ n[71];
assign t[72] = t[71] ^ n[72];
assign t[73] = t[72] ^ n[73];
assign t[74] = t[73] ^ n[74];
assign t[75] = t[74] ^ n[75];
assign t[76] = t[75] ^ n[76];
assign t[77] = t[76] ^ n[77];
assign t[78] = t[77] ^ n[78];
assign t[79] = t[78] ^ n[79];
assign t[80] = t[79] ^ n[80];
assign t[81] = t[80] ^ n[81];
assign t[82] = t[81] ^ n[82];
assign t[83] = t[82] ^ n[83];
assign t[84] = t[83] ^ n[84];
assign t[85] = t[84] ^ n[85];
assign t[86] = t[85] ^ n[86];
assign t[87] = t[86] ^ n[87];
assign t[88] = t[87] ^ n[88];
assign t[89] = t[88] ^ n[89];
assign t[90] = t[89] ^ n[90];
assign t[91] = t[90] ^ n[91];
assign t[92] = t[91] ^ n[92];
assign t[93] = t[92] ^ n[93];
assign t[94] = t[93] ^ n[94];
assign t[95] = t[94] ^ n[95];
assign t[96] = t[95] ^ n[96];
assign t[97] = t[96] ^ n[97];
assign t[98] = t[97] ^ n[98];
assign t[99] = t[98] ^ n[99];
assign t[100] = t[99] ^ n[100];
assign t[101] = t[100] ^ n[101];
assign t[102] = t[101] ^ n[102];
assign t[103] = t[102] ^ n[103];
assign t[104] = t[103] ^ n[104];
assign t[105] = t[104] ^ n[105];
assign t[106] = t[105] ^ n[106];
assign t[107] = t[106] ^ n[107];
assign t[108] = t[107] ^ n[108];
assign t[109] = t[108] ^ n[109];
assign t[110] = t[109] ^ n[110];
assign t[111] = t[110] ^ n[111];
assign t[112] = t[111] ^ n[112];
assign t[113] = t[112] ^ n[113];
assign t[114] = t[113] ^ n[114];
assign t[115] = t[114] ^ n[115];
assign t[116] = t[115] ^ n[116];
assign t[117] = t[116] ^ n[117];
assign t[118] = t[117] ^ n[118];
assign t[119] = t[118] ^ n[119];

//asigning bit 6
assign s[6] = ( a[6] ^ b [6] ) ^ t[119];

assign t[120] = n[120];
assign t[121] = t[120] ^ n[121];
assign t[122] = t[121] ^ n[122];
assign t[123] = t[122] ^ n[123];
assign t[124] = t[123] ^ n[124];
assign t[125] = t[124] ^ n[125];
assign t[126] = t[125] ^ n[126];
assign t[127] = t[126] ^ n[127];
assign t[128] = t[127] ^ n[128];
assign t[129] = t[128] ^ n[129];
assign t[130] = t[129] ^ n[130];
assign t[131] = t[130] ^ n[131];
assign t[132] = t[131] ^ n[132];
assign t[133] = t[132] ^ n[133];
assign t[134] = t[133] ^ n[134];
assign t[135] = t[134] ^ n[135];
assign t[136] = t[135] ^ n[136];
assign t[137] = t[136] ^ n[137];
assign t[138] = t[137] ^ n[138];
assign t[139] = t[138] ^ n[139];
assign t[140] = t[139] ^ n[140];
assign t[141] = t[140] ^ n[141];
assign t[142] = t[141] ^ n[142];
assign t[143] = t[142] ^ n[143];
assign t[144] = t[143] ^ n[144];
assign t[145] = t[144] ^ n[145];
assign t[146] = t[145] ^ n[146];
assign t[147] = t[146] ^ n[147];
assign t[148] = t[147] ^ n[148];
assign t[149] = t[148] ^ n[149];
assign t[150] = t[149] ^ n[150];
assign t[151] = t[150] ^ n[151];
assign t[152] = t[151] ^ n[152];
assign t[153] = t[152] ^ n[153];
assign t[154] = t[153] ^ n[154];
assign t[155] = t[154] ^ n[155];
assign t[156] = t[155] ^ n[156];
assign t[157] = t[156] ^ n[157];
assign t[158] = t[157] ^ n[158];
assign t[159] = t[158] ^ n[159];
assign t[160] = t[159] ^ n[160];
assign t[161] = t[160] ^ n[161];
assign t[162] = t[161] ^ n[162];
assign t[163] = t[162] ^ n[163];
assign t[164] = t[163] ^ n[164];
assign t[165] = t[164] ^ n[165];
assign t[166] = t[165] ^ n[166];
assign t[167] = t[166] ^ n[167];
assign t[168] = t[167] ^ n[168];
assign t[169] = t[168] ^ n[169];
assign t[170] = t[169] ^ n[170];
assign t[171] = t[170] ^ n[171];
assign t[172] = t[171] ^ n[172];
assign t[173] = t[172] ^ n[173];
assign t[174] = t[173] ^ n[174];
assign t[175] = t[174] ^ n[175];
assign t[176] = t[175] ^ n[176];
assign t[177] = t[176] ^ n[177];
assign t[178] = t[177] ^ n[178];
assign t[179] = t[178] ^ n[179];
assign t[180] = t[179] ^ n[180];
assign t[181] = t[180] ^ n[181];
assign t[182] = t[181] ^ n[182];
assign t[183] = t[182] ^ n[183];
assign t[184] = t[183] ^ n[184];
assign t[185] = t[184] ^ n[185];
assign t[186] = t[185] ^ n[186];
assign t[187] = t[186] ^ n[187];
assign t[188] = t[187] ^ n[188];
assign t[189] = t[188] ^ n[189];
assign t[190] = t[189] ^ n[190];
assign t[191] = t[190] ^ n[191];
assign t[192] = t[191] ^ n[192];
assign t[193] = t[192] ^ n[193];
assign t[194] = t[193] ^ n[194];
assign t[195] = t[194] ^ n[195];
assign t[196] = t[195] ^ n[196];
assign t[197] = t[196] ^ n[197];
assign t[198] = t[197] ^ n[198];
assign t[199] = t[198] ^ n[199];
assign t[200] = t[199] ^ n[200];
assign t[201] = t[200] ^ n[201];
assign t[202] = t[201] ^ n[202];
assign t[203] = t[202] ^ n[203];
assign t[204] = t[203] ^ n[204];
assign t[205] = t[204] ^ n[205];
assign t[206] = t[205] ^ n[206];
assign t[207] = t[206] ^ n[207];
assign t[208] = t[207] ^ n[208];
assign t[209] = t[208] ^ n[209];
assign t[210] = t[209] ^ n[210];
assign t[211] = t[210] ^ n[211];
assign t[212] = t[211] ^ n[212];
assign t[213] = t[212] ^ n[213];
assign t[214] = t[213] ^ n[214];
assign t[215] = t[214] ^ n[215];
assign t[216] = t[215] ^ n[216];
assign t[217] = t[216] ^ n[217];
assign t[218] = t[217] ^ n[218];
assign t[219] = t[218] ^ n[219];
assign t[220] = t[219] ^ n[220];
assign t[221] = t[220] ^ n[221];
assign t[222] = t[221] ^ n[222];
assign t[223] = t[222] ^ n[223];
assign t[224] = t[223] ^ n[224];
assign t[225] = t[224] ^ n[225];
assign t[226] = t[225] ^ n[226];
assign t[227] = t[226] ^ n[227];
assign t[228] = t[227] ^ n[228];
assign t[229] = t[228] ^ n[229];
assign t[230] = t[229] ^ n[230];
assign t[231] = t[230] ^ n[231];
assign t[232] = t[231] ^ n[232];
assign t[233] = t[232] ^ n[233];
assign t[234] = t[233] ^ n[234];
assign t[235] = t[234] ^ n[235];
assign t[236] = t[235] ^ n[236];
assign t[237] = t[236] ^ n[237];
assign t[238] = t[237] ^ n[238];
assign t[239] = t[238] ^ n[239];
assign t[240] = t[239] ^ n[240];
assign t[241] = t[240] ^ n[241];
assign t[242] = t[241] ^ n[242];
assign t[243] = t[242] ^ n[243];
assign t[244] = t[243] ^ n[244];
assign t[245] = t[244] ^ n[245];
assign t[246] = t[245] ^ n[246];

//asigning bit 7
assign s[7] = ( a[7] ^ b [7] ) ^ t[246];

assign t[247] = n[247];
assign t[248] = t[247] ^ n[248];
assign t[249] = t[248] ^ n[249];
assign t[250] = t[249] ^ n[250];
assign t[251] = t[250] ^ n[251];
assign t[252] = t[251] ^ n[252];
assign t[253] = t[252] ^ n[253];
assign t[254] = t[253] ^ n[254];
assign t[255] = t[254] ^ n[255];
assign t[256] = t[255] ^ n[256];
assign t[257] = t[256] ^ n[257];
assign t[258] = t[257] ^ n[258];
assign t[259] = t[258] ^ n[259];
assign t[260] = t[259] ^ n[260];
assign t[261] = t[260] ^ n[261];
assign t[262] = t[261] ^ n[262];
assign t[263] = t[262] ^ n[263];
assign t[264] = t[263] ^ n[264];
assign t[265] = t[264] ^ n[265];
assign t[266] = t[265] ^ n[266];
assign t[267] = t[266] ^ n[267];
assign t[268] = t[267] ^ n[268];
assign t[269] = t[268] ^ n[269];
assign t[270] = t[269] ^ n[270];
assign t[271] = t[270] ^ n[271];
assign t[272] = t[271] ^ n[272];
assign t[273] = t[272] ^ n[273];
assign t[274] = t[273] ^ n[274];
assign t[275] = t[274] ^ n[275];
assign t[276] = t[275] ^ n[276];
assign t[277] = t[276] ^ n[277];
assign t[278] = t[277] ^ n[278];
assign t[279] = t[278] ^ n[279];
assign t[280] = t[279] ^ n[280];
assign t[281] = t[280] ^ n[281];
assign t[282] = t[281] ^ n[282];
assign t[283] = t[282] ^ n[283];
assign t[284] = t[283] ^ n[284];
assign t[285] = t[284] ^ n[285];
assign t[286] = t[285] ^ n[286];
assign t[287] = t[286] ^ n[287];
assign t[288] = t[287] ^ n[288];
assign t[289] = t[288] ^ n[289];
assign t[290] = t[289] ^ n[290];
assign t[291] = t[290] ^ n[291];
assign t[292] = t[291] ^ n[292];
assign t[293] = t[292] ^ n[293];
assign t[294] = t[293] ^ n[294];
assign t[295] = t[294] ^ n[295];
assign t[296] = t[295] ^ n[296];
assign t[297] = t[296] ^ n[297];
assign t[298] = t[297] ^ n[298];
assign t[299] = t[298] ^ n[299];
assign t[300] = t[299] ^ n[300];
assign t[301] = t[300] ^ n[301];
assign t[302] = t[301] ^ n[302];
assign t[303] = t[302] ^ n[303];
assign t[304] = t[303] ^ n[304];
assign t[305] = t[304] ^ n[305];
assign t[306] = t[305] ^ n[306];
assign t[307] = t[306] ^ n[307];
assign t[308] = t[307] ^ n[308];
assign t[309] = t[308] ^ n[309];
assign t[310] = t[309] ^ n[310];
assign t[311] = t[310] ^ n[311];
assign t[312] = t[311] ^ n[312];
assign t[313] = t[312] ^ n[313];
assign t[314] = t[313] ^ n[314];
assign t[315] = t[314] ^ n[315];
assign t[316] = t[315] ^ n[316];
assign t[317] = t[316] ^ n[317];
assign t[318] = t[317] ^ n[318];
assign t[319] = t[318] ^ n[319];
assign t[320] = t[319] ^ n[320];
assign t[321] = t[320] ^ n[321];
assign t[322] = t[321] ^ n[322];
assign t[323] = t[322] ^ n[323];
assign t[324] = t[323] ^ n[324];
assign t[325] = t[324] ^ n[325];
assign t[326] = t[325] ^ n[326];
assign t[327] = t[326] ^ n[327];
assign t[328] = t[327] ^ n[328];
assign t[329] = t[328] ^ n[329];
assign t[330] = t[329] ^ n[330];
assign t[331] = t[330] ^ n[331];
assign t[332] = t[331] ^ n[332];
assign t[333] = t[332] ^ n[333];
assign t[334] = t[333] ^ n[334];
assign t[335] = t[334] ^ n[335];
assign t[336] = t[335] ^ n[336];
assign t[337] = t[336] ^ n[337];
assign t[338] = t[337] ^ n[338];
assign t[339] = t[338] ^ n[339];
assign t[340] = t[339] ^ n[340];
assign t[341] = t[340] ^ n[341];
assign t[342] = t[341] ^ n[342];
assign t[343] = t[342] ^ n[343];
assign t[344] = t[343] ^ n[344];
assign t[345] = t[344] ^ n[345];
assign t[346] = t[345] ^ n[346];
assign t[347] = t[346] ^ n[347];
assign t[348] = t[347] ^ n[348];
assign t[349] = t[348] ^ n[349];
assign t[350] = t[349] ^ n[350];
assign t[351] = t[350] ^ n[351];
assign t[352] = t[351] ^ n[352];
assign t[353] = t[352] ^ n[353];
assign t[354] = t[353] ^ n[354];
assign t[355] = t[354] ^ n[355];
assign t[356] = t[355] ^ n[356];
assign t[357] = t[356] ^ n[357];
assign t[358] = t[357] ^ n[358];
assign t[359] = t[358] ^ n[359];
assign t[360] = t[359] ^ n[360];
assign t[361] = t[360] ^ n[361];
assign t[362] = t[361] ^ n[362];
assign t[363] = t[362] ^ n[363];
assign t[364] = t[363] ^ n[364];
assign t[365] = t[364] ^ n[365];
assign t[366] = t[365] ^ n[366];
assign t[367] = t[366] ^ n[367];
assign t[368] = t[367] ^ n[368];
assign t[369] = t[368] ^ n[369];
assign t[370] = t[369] ^ n[370];
assign t[371] = t[370] ^ n[371];
assign t[372] = t[371] ^ n[372];
assign t[373] = t[372] ^ n[373];
assign t[374] = t[373] ^ n[374];
assign t[375] = t[374] ^ n[375];
assign t[376] = t[375] ^ n[376];
assign t[377] = t[376] ^ n[377];
assign t[378] = t[377] ^ n[378];
assign t[379] = t[378] ^ n[379];
assign t[380] = t[379] ^ n[380];
assign t[381] = t[380] ^ n[381];
assign t[382] = t[381] ^ n[382];
assign t[383] = t[382] ^ n[383];
assign t[384] = t[383] ^ n[384];
assign t[385] = t[384] ^ n[385];
assign t[386] = t[385] ^ n[386];
assign t[387] = t[386] ^ n[387];
assign t[388] = t[387] ^ n[388];
assign t[389] = t[388] ^ n[389];
assign t[390] = t[389] ^ n[390];
assign t[391] = t[390] ^ n[391];
assign t[392] = t[391] ^ n[392];
assign t[393] = t[392] ^ n[393];
assign t[394] = t[393] ^ n[394];
assign t[395] = t[394] ^ n[395];
assign t[396] = t[395] ^ n[396];
assign t[397] = t[396] ^ n[397];
assign t[398] = t[397] ^ n[398];
assign t[399] = t[398] ^ n[399];
assign t[400] = t[399] ^ n[400];
assign t[401] = t[400] ^ n[401];
assign t[402] = t[401] ^ n[402];
assign t[403] = t[402] ^ n[403];
assign t[404] = t[403] ^ n[404];
assign t[405] = t[404] ^ n[405];
assign t[406] = t[405] ^ n[406];
assign t[407] = t[406] ^ n[407];
assign t[408] = t[407] ^ n[408];
assign t[409] = t[408] ^ n[409];
assign t[410] = t[409] ^ n[410];
assign t[411] = t[410] ^ n[411];
assign t[412] = t[411] ^ n[412];
assign t[413] = t[412] ^ n[413];
assign t[414] = t[413] ^ n[414];
assign t[415] = t[414] ^ n[415];
assign t[416] = t[415] ^ n[416];
assign t[417] = t[416] ^ n[417];
assign t[418] = t[417] ^ n[418];
assign t[419] = t[418] ^ n[419];
assign t[420] = t[419] ^ n[420];
assign t[421] = t[420] ^ n[421];
assign t[422] = t[421] ^ n[422];
assign t[423] = t[422] ^ n[423];
assign t[424] = t[423] ^ n[424];
assign t[425] = t[424] ^ n[425];
assign t[426] = t[425] ^ n[426];
assign t[427] = t[426] ^ n[427];
assign t[428] = t[427] ^ n[428];
assign t[429] = t[428] ^ n[429];
assign t[430] = t[429] ^ n[430];
assign t[431] = t[430] ^ n[431];
assign t[432] = t[431] ^ n[432];
assign t[433] = t[432] ^ n[433];
assign t[434] = t[433] ^ n[434];
assign t[435] = t[434] ^ n[435];
assign t[436] = t[435] ^ n[436];
assign t[437] = t[436] ^ n[437];
assign t[438] = t[437] ^ n[438];
assign t[439] = t[438] ^ n[439];
assign t[440] = t[439] ^ n[440];
assign t[441] = t[440] ^ n[441];
assign t[442] = t[441] ^ n[442];
assign t[443] = t[442] ^ n[443];
assign t[444] = t[443] ^ n[444];
assign t[445] = t[444] ^ n[445];
assign t[446] = t[445] ^ n[446];
assign t[447] = t[446] ^ n[447];
assign t[448] = t[447] ^ n[448];
assign t[449] = t[448] ^ n[449];
assign t[450] = t[449] ^ n[450];
assign t[451] = t[450] ^ n[451];
assign t[452] = t[451] ^ n[452];
assign t[453] = t[452] ^ n[453];
assign t[454] = t[453] ^ n[454];
assign t[455] = t[454] ^ n[455];
assign t[456] = t[455] ^ n[456];
assign t[457] = t[456] ^ n[457];
assign t[458] = t[457] ^ n[458];
assign t[459] = t[458] ^ n[459];
assign t[460] = t[459] ^ n[460];
assign t[461] = t[460] ^ n[461];
assign t[462] = t[461] ^ n[462];
assign t[463] = t[462] ^ n[463];
assign t[464] = t[463] ^ n[464];
assign t[465] = t[464] ^ n[465];
assign t[466] = t[465] ^ n[466];
assign t[467] = t[466] ^ n[467];
assign t[468] = t[467] ^ n[468];
assign t[469] = t[468] ^ n[469];
assign t[470] = t[469] ^ n[470];
assign t[471] = t[470] ^ n[471];
assign t[472] = t[471] ^ n[472];
assign t[473] = t[472] ^ n[473];
assign t[474] = t[473] ^ n[474];
assign t[475] = t[474] ^ n[475];
assign t[476] = t[475] ^ n[476];
assign t[477] = t[476] ^ n[477];
assign t[478] = t[477] ^ n[478];
assign t[479] = t[478] ^ n[479];
assign t[480] = t[479] ^ n[480];
assign t[481] = t[480] ^ n[481];
assign t[482] = t[481] ^ n[482];
assign t[483] = t[482] ^ n[483];
assign t[484] = t[483] ^ n[484];
assign t[485] = t[484] ^ n[485];
assign t[486] = t[485] ^ n[486];
assign t[487] = t[486] ^ n[487];
assign t[488] = t[487] ^ n[488];
assign t[489] = t[488] ^ n[489];
assign t[490] = t[489] ^ n[490];
assign t[491] = t[490] ^ n[491];
assign t[492] = t[491] ^ n[492];
assign t[493] = t[492] ^ n[493];
assign t[494] = t[493] ^ n[494];
assign t[495] = t[494] ^ n[495];
assign t[496] = t[495] ^ n[496];
assign t[497] = t[496] ^ n[497];
assign t[498] = t[497] ^ n[498];
assign t[499] = t[498] ^ n[499];
assign t[500] = t[499] ^ n[500];
assign t[501] = t[500] ^ n[501];

//asigning bit 8
assign s[8] = ( a[8] ^ b [8] ) ^ t[501];

assign t[502] = n[502];
assign t[503] = t[502] ^ n[503];
assign t[504] = t[503] ^ n[504];
assign t[505] = t[504] ^ n[505];
assign t[506] = t[505] ^ n[506];
assign t[507] = t[506] ^ n[507];
assign t[508] = t[507] ^ n[508];
assign t[509] = t[508] ^ n[509];
assign t[510] = t[509] ^ n[510];
assign t[511] = t[510] ^ n[511];
assign t[512] = t[511] ^ n[512];
assign t[513] = t[512] ^ n[513];
assign t[514] = t[513] ^ n[514];
assign t[515] = t[514] ^ n[515];
assign t[516] = t[515] ^ n[516];
assign t[517] = t[516] ^ n[517];
assign t[518] = t[517] ^ n[518];
assign t[519] = t[518] ^ n[519];
assign t[520] = t[519] ^ n[520];
assign t[521] = t[520] ^ n[521];
assign t[522] = t[521] ^ n[522];
assign t[523] = t[522] ^ n[523];
assign t[524] = t[523] ^ n[524];
assign t[525] = t[524] ^ n[525];
assign t[526] = t[525] ^ n[526];
assign t[527] = t[526] ^ n[527];
assign t[528] = t[527] ^ n[528];
assign t[529] = t[528] ^ n[529];
assign t[530] = t[529] ^ n[530];
assign t[531] = t[530] ^ n[531];
assign t[532] = t[531] ^ n[532];
assign t[533] = t[532] ^ n[533];
assign t[534] = t[533] ^ n[534];
assign t[535] = t[534] ^ n[535];
assign t[536] = t[535] ^ n[536];
assign t[537] = t[536] ^ n[537];
assign t[538] = t[537] ^ n[538];
assign t[539] = t[538] ^ n[539];
assign t[540] = t[539] ^ n[540];
assign t[541] = t[540] ^ n[541];
assign t[542] = t[541] ^ n[542];
assign t[543] = t[542] ^ n[543];
assign t[544] = t[543] ^ n[544];
assign t[545] = t[544] ^ n[545];
assign t[546] = t[545] ^ n[546];
assign t[547] = t[546] ^ n[547];
assign t[548] = t[547] ^ n[548];
assign t[549] = t[548] ^ n[549];
assign t[550] = t[549] ^ n[550];
assign t[551] = t[550] ^ n[551];
assign t[552] = t[551] ^ n[552];
assign t[553] = t[552] ^ n[553];
assign t[554] = t[553] ^ n[554];
assign t[555] = t[554] ^ n[555];
assign t[556] = t[555] ^ n[556];
assign t[557] = t[556] ^ n[557];
assign t[558] = t[557] ^ n[558];
assign t[559] = t[558] ^ n[559];
assign t[560] = t[559] ^ n[560];
assign t[561] = t[560] ^ n[561];
assign t[562] = t[561] ^ n[562];
assign t[563] = t[562] ^ n[563];
assign t[564] = t[563] ^ n[564];
assign t[565] = t[564] ^ n[565];
assign t[566] = t[565] ^ n[566];
assign t[567] = t[566] ^ n[567];
assign t[568] = t[567] ^ n[568];
assign t[569] = t[568] ^ n[569];
assign t[570] = t[569] ^ n[570];
assign t[571] = t[570] ^ n[571];
assign t[572] = t[571] ^ n[572];
assign t[573] = t[572] ^ n[573];
assign t[574] = t[573] ^ n[574];
assign t[575] = t[574] ^ n[575];
assign t[576] = t[575] ^ n[576];
assign t[577] = t[576] ^ n[577];
assign t[578] = t[577] ^ n[578];
assign t[579] = t[578] ^ n[579];
assign t[580] = t[579] ^ n[580];
assign t[581] = t[580] ^ n[581];
assign t[582] = t[581] ^ n[582];
assign t[583] = t[582] ^ n[583];
assign t[584] = t[583] ^ n[584];
assign t[585] = t[584] ^ n[585];
assign t[586] = t[585] ^ n[586];
assign t[587] = t[586] ^ n[587];
assign t[588] = t[587] ^ n[588];
assign t[589] = t[588] ^ n[589];
assign t[590] = t[589] ^ n[590];
assign t[591] = t[590] ^ n[591];
assign t[592] = t[591] ^ n[592];
assign t[593] = t[592] ^ n[593];
assign t[594] = t[593] ^ n[594];
assign t[595] = t[594] ^ n[595];
assign t[596] = t[595] ^ n[596];
assign t[597] = t[596] ^ n[597];
assign t[598] = t[597] ^ n[598];
assign t[599] = t[598] ^ n[599];
assign t[600] = t[599] ^ n[600];
assign t[601] = t[600] ^ n[601];
assign t[602] = t[601] ^ n[602];
assign t[603] = t[602] ^ n[603];
assign t[604] = t[603] ^ n[604];
assign t[605] = t[604] ^ n[605];
assign t[606] = t[605] ^ n[606];
assign t[607] = t[606] ^ n[607];
assign t[608] = t[607] ^ n[608];
assign t[609] = t[608] ^ n[609];
assign t[610] = t[609] ^ n[610];
assign t[611] = t[610] ^ n[611];
assign t[612] = t[611] ^ n[612];
assign t[613] = t[612] ^ n[613];
assign t[614] = t[613] ^ n[614];
assign t[615] = t[614] ^ n[615];
assign t[616] = t[615] ^ n[616];
assign t[617] = t[616] ^ n[617];
assign t[618] = t[617] ^ n[618];
assign t[619] = t[618] ^ n[619];
assign t[620] = t[619] ^ n[620];
assign t[621] = t[620] ^ n[621];
assign t[622] = t[621] ^ n[622];
assign t[623] = t[622] ^ n[623];
assign t[624] = t[623] ^ n[624];
assign t[625] = t[624] ^ n[625];
assign t[626] = t[625] ^ n[626];
assign t[627] = t[626] ^ n[627];
assign t[628] = t[627] ^ n[628];
assign t[629] = t[628] ^ n[629];
assign t[630] = t[629] ^ n[630];
assign t[631] = t[630] ^ n[631];
assign t[632] = t[631] ^ n[632];
assign t[633] = t[632] ^ n[633];
assign t[634] = t[633] ^ n[634];
assign t[635] = t[634] ^ n[635];
assign t[636] = t[635] ^ n[636];
assign t[637] = t[636] ^ n[637];
assign t[638] = t[637] ^ n[638];
assign t[639] = t[638] ^ n[639];
assign t[640] = t[639] ^ n[640];
assign t[641] = t[640] ^ n[641];
assign t[642] = t[641] ^ n[642];
assign t[643] = t[642] ^ n[643];
assign t[644] = t[643] ^ n[644];
assign t[645] = t[644] ^ n[645];
assign t[646] = t[645] ^ n[646];
assign t[647] = t[646] ^ n[647];
assign t[648] = t[647] ^ n[648];
assign t[649] = t[648] ^ n[649];
assign t[650] = t[649] ^ n[650];
assign t[651] = t[650] ^ n[651];
assign t[652] = t[651] ^ n[652];
assign t[653] = t[652] ^ n[653];
assign t[654] = t[653] ^ n[654];
assign t[655] = t[654] ^ n[655];
assign t[656] = t[655] ^ n[656];
assign t[657] = t[656] ^ n[657];
assign t[658] = t[657] ^ n[658];
assign t[659] = t[658] ^ n[659];
assign t[660] = t[659] ^ n[660];
assign t[661] = t[660] ^ n[661];
assign t[662] = t[661] ^ n[662];
assign t[663] = t[662] ^ n[663];
assign t[664] = t[663] ^ n[664];
assign t[665] = t[664] ^ n[665];
assign t[666] = t[665] ^ n[666];
assign t[667] = t[666] ^ n[667];
assign t[668] = t[667] ^ n[668];
assign t[669] = t[668] ^ n[669];
assign t[670] = t[669] ^ n[670];
assign t[671] = t[670] ^ n[671];
assign t[672] = t[671] ^ n[672];
assign t[673] = t[672] ^ n[673];
assign t[674] = t[673] ^ n[674];
assign t[675] = t[674] ^ n[675];
assign t[676] = t[675] ^ n[676];
assign t[677] = t[676] ^ n[677];
assign t[678] = t[677] ^ n[678];
assign t[679] = t[678] ^ n[679];
assign t[680] = t[679] ^ n[680];
assign t[681] = t[680] ^ n[681];
assign t[682] = t[681] ^ n[682];
assign t[683] = t[682] ^ n[683];
assign t[684] = t[683] ^ n[684];
assign t[685] = t[684] ^ n[685];
assign t[686] = t[685] ^ n[686];
assign t[687] = t[686] ^ n[687];
assign t[688] = t[687] ^ n[688];
assign t[689] = t[688] ^ n[689];
assign t[690] = t[689] ^ n[690];
assign t[691] = t[690] ^ n[691];
assign t[692] = t[691] ^ n[692];
assign t[693] = t[692] ^ n[693];
assign t[694] = t[693] ^ n[694];
assign t[695] = t[694] ^ n[695];
assign t[696] = t[695] ^ n[696];
assign t[697] = t[696] ^ n[697];
assign t[698] = t[697] ^ n[698];
assign t[699] = t[698] ^ n[699];
assign t[700] = t[699] ^ n[700];
assign t[701] = t[700] ^ n[701];
assign t[702] = t[701] ^ n[702];
assign t[703] = t[702] ^ n[703];
assign t[704] = t[703] ^ n[704];
assign t[705] = t[704] ^ n[705];
assign t[706] = t[705] ^ n[706];
assign t[707] = t[706] ^ n[707];
assign t[708] = t[707] ^ n[708];
assign t[709] = t[708] ^ n[709];
assign t[710] = t[709] ^ n[710];
assign t[711] = t[710] ^ n[711];
assign t[712] = t[711] ^ n[712];
assign t[713] = t[712] ^ n[713];
assign t[714] = t[713] ^ n[714];
assign t[715] = t[714] ^ n[715];
assign t[716] = t[715] ^ n[716];
assign t[717] = t[716] ^ n[717];
assign t[718] = t[717] ^ n[718];
assign t[719] = t[718] ^ n[719];
assign t[720] = t[719] ^ n[720];
assign t[721] = t[720] ^ n[721];
assign t[722] = t[721] ^ n[722];
assign t[723] = t[722] ^ n[723];
assign t[724] = t[723] ^ n[724];
assign t[725] = t[724] ^ n[725];
assign t[726] = t[725] ^ n[726];
assign t[727] = t[726] ^ n[727];
assign t[728] = t[727] ^ n[728];
assign t[729] = t[728] ^ n[729];
assign t[730] = t[729] ^ n[730];
assign t[731] = t[730] ^ n[731];
assign t[732] = t[731] ^ n[732];
assign t[733] = t[732] ^ n[733];
assign t[734] = t[733] ^ n[734];
assign t[735] = t[734] ^ n[735];
assign t[736] = t[735] ^ n[736];
assign t[737] = t[736] ^ n[737];
assign t[738] = t[737] ^ n[738];
assign t[739] = t[738] ^ n[739];
assign t[740] = t[739] ^ n[740];
assign t[741] = t[740] ^ n[741];
assign t[742] = t[741] ^ n[742];
assign t[743] = t[742] ^ n[743];
assign t[744] = t[743] ^ n[744];
assign t[745] = t[744] ^ n[745];
assign t[746] = t[745] ^ n[746];
assign t[747] = t[746] ^ n[747];
assign t[748] = t[747] ^ n[748];
assign t[749] = t[748] ^ n[749];
assign t[750] = t[749] ^ n[750];
assign t[751] = t[750] ^ n[751];
assign t[752] = t[751] ^ n[752];
assign t[753] = t[752] ^ n[753];
assign t[754] = t[753] ^ n[754];
assign t[755] = t[754] ^ n[755];
assign t[756] = t[755] ^ n[756];
assign t[757] = t[756] ^ n[757];
assign t[758] = t[757] ^ n[758];
assign t[759] = t[758] ^ n[759];
assign t[760] = t[759] ^ n[760];
assign t[761] = t[760] ^ n[761];
assign t[762] = t[761] ^ n[762];
assign t[763] = t[762] ^ n[763];
assign t[764] = t[763] ^ n[764];
assign t[765] = t[764] ^ n[765];
assign t[766] = t[765] ^ n[766];
assign t[767] = t[766] ^ n[767];
assign t[768] = t[767] ^ n[768];
assign t[769] = t[768] ^ n[769];
assign t[770] = t[769] ^ n[770];
assign t[771] = t[770] ^ n[771];
assign t[772] = t[771] ^ n[772];
assign t[773] = t[772] ^ n[773];
assign t[774] = t[773] ^ n[774];
assign t[775] = t[774] ^ n[775];
assign t[776] = t[775] ^ n[776];
assign t[777] = t[776] ^ n[777];
assign t[778] = t[777] ^ n[778];
assign t[779] = t[778] ^ n[779];
assign t[780] = t[779] ^ n[780];
assign t[781] = t[780] ^ n[781];
assign t[782] = t[781] ^ n[782];
assign t[783] = t[782] ^ n[783];
assign t[784] = t[783] ^ n[784];
assign t[785] = t[784] ^ n[785];
assign t[786] = t[785] ^ n[786];
assign t[787] = t[786] ^ n[787];
assign t[788] = t[787] ^ n[788];
assign t[789] = t[788] ^ n[789];
assign t[790] = t[789] ^ n[790];
assign t[791] = t[790] ^ n[791];
assign t[792] = t[791] ^ n[792];
assign t[793] = t[792] ^ n[793];
assign t[794] = t[793] ^ n[794];
assign t[795] = t[794] ^ n[795];
assign t[796] = t[795] ^ n[796];
assign t[797] = t[796] ^ n[797];
assign t[798] = t[797] ^ n[798];
assign t[799] = t[798] ^ n[799];
assign t[800] = t[799] ^ n[800];
assign t[801] = t[800] ^ n[801];
assign t[802] = t[801] ^ n[802];
assign t[803] = t[802] ^ n[803];
assign t[804] = t[803] ^ n[804];
assign t[805] = t[804] ^ n[805];
assign t[806] = t[805] ^ n[806];
assign t[807] = t[806] ^ n[807];
assign t[808] = t[807] ^ n[808];
assign t[809] = t[808] ^ n[809];
assign t[810] = t[809] ^ n[810];
assign t[811] = t[810] ^ n[811];
assign t[812] = t[811] ^ n[812];
assign t[813] = t[812] ^ n[813];
assign t[814] = t[813] ^ n[814];
assign t[815] = t[814] ^ n[815];
assign t[816] = t[815] ^ n[816];
assign t[817] = t[816] ^ n[817];
assign t[818] = t[817] ^ n[818];
assign t[819] = t[818] ^ n[819];
assign t[820] = t[819] ^ n[820];
assign t[821] = t[820] ^ n[821];
assign t[822] = t[821] ^ n[822];
assign t[823] = t[822] ^ n[823];
assign t[824] = t[823] ^ n[824];
assign t[825] = t[824] ^ n[825];
assign t[826] = t[825] ^ n[826];
assign t[827] = t[826] ^ n[827];
assign t[828] = t[827] ^ n[828];
assign t[829] = t[828] ^ n[829];
assign t[830] = t[829] ^ n[830];
assign t[831] = t[830] ^ n[831];
assign t[832] = t[831] ^ n[832];
assign t[833] = t[832] ^ n[833];
assign t[834] = t[833] ^ n[834];
assign t[835] = t[834] ^ n[835];
assign t[836] = t[835] ^ n[836];
assign t[837] = t[836] ^ n[837];
assign t[838] = t[837] ^ n[838];
assign t[839] = t[838] ^ n[839];
assign t[840] = t[839] ^ n[840];
assign t[841] = t[840] ^ n[841];
assign t[842] = t[841] ^ n[842];
assign t[843] = t[842] ^ n[843];
assign t[844] = t[843] ^ n[844];
assign t[845] = t[844] ^ n[845];
assign t[846] = t[845] ^ n[846];
assign t[847] = t[846] ^ n[847];
assign t[848] = t[847] ^ n[848];
assign t[849] = t[848] ^ n[849];
assign t[850] = t[849] ^ n[850];
assign t[851] = t[850] ^ n[851];
assign t[852] = t[851] ^ n[852];
assign t[853] = t[852] ^ n[853];
assign t[854] = t[853] ^ n[854];
assign t[855] = t[854] ^ n[855];
assign t[856] = t[855] ^ n[856];
assign t[857] = t[856] ^ n[857];
assign t[858] = t[857] ^ n[858];
assign t[859] = t[858] ^ n[859];
assign t[860] = t[859] ^ n[860];
assign t[861] = t[860] ^ n[861];
assign t[862] = t[861] ^ n[862];
assign t[863] = t[862] ^ n[863];
assign t[864] = t[863] ^ n[864];
assign t[865] = t[864] ^ n[865];
assign t[866] = t[865] ^ n[866];
assign t[867] = t[866] ^ n[867];
assign t[868] = t[867] ^ n[868];
assign t[869] = t[868] ^ n[869];
assign t[870] = t[869] ^ n[870];
assign t[871] = t[870] ^ n[871];
assign t[872] = t[871] ^ n[872];
assign t[873] = t[872] ^ n[873];
assign t[874] = t[873] ^ n[874];
assign t[875] = t[874] ^ n[875];
assign t[876] = t[875] ^ n[876];
assign t[877] = t[876] ^ n[877];
assign t[878] = t[877] ^ n[878];
assign t[879] = t[878] ^ n[879];
assign t[880] = t[879] ^ n[880];
assign t[881] = t[880] ^ n[881];
assign t[882] = t[881] ^ n[882];
assign t[883] = t[882] ^ n[883];
assign t[884] = t[883] ^ n[884];
assign t[885] = t[884] ^ n[885];
assign t[886] = t[885] ^ n[886];
assign t[887] = t[886] ^ n[887];
assign t[888] = t[887] ^ n[888];
assign t[889] = t[888] ^ n[889];
assign t[890] = t[889] ^ n[890];
assign t[891] = t[890] ^ n[891];
assign t[892] = t[891] ^ n[892];
assign t[893] = t[892] ^ n[893];
assign t[894] = t[893] ^ n[894];
assign t[895] = t[894] ^ n[895];
assign t[896] = t[895] ^ n[896];
assign t[897] = t[896] ^ n[897];
assign t[898] = t[897] ^ n[898];
assign t[899] = t[898] ^ n[899];
assign t[900] = t[899] ^ n[900];
assign t[901] = t[900] ^ n[901];
assign t[902] = t[901] ^ n[902];
assign t[903] = t[902] ^ n[903];
assign t[904] = t[903] ^ n[904];
assign t[905] = t[904] ^ n[905];
assign t[906] = t[905] ^ n[906];
assign t[907] = t[906] ^ n[907];
assign t[908] = t[907] ^ n[908];
assign t[909] = t[908] ^ n[909];
assign t[910] = t[909] ^ n[910];
assign t[911] = t[910] ^ n[911];
assign t[912] = t[911] ^ n[912];
assign t[913] = t[912] ^ n[913];
assign t[914] = t[913] ^ n[914];
assign t[915] = t[914] ^ n[915];
assign t[916] = t[915] ^ n[916];
assign t[917] = t[916] ^ n[917];
assign t[918] = t[917] ^ n[918];
assign t[919] = t[918] ^ n[919];
assign t[920] = t[919] ^ n[920];
assign t[921] = t[920] ^ n[921];
assign t[922] = t[921] ^ n[922];
assign t[923] = t[922] ^ n[923];
assign t[924] = t[923] ^ n[924];
assign t[925] = t[924] ^ n[925];
assign t[926] = t[925] ^ n[926];
assign t[927] = t[926] ^ n[927];
assign t[928] = t[927] ^ n[928];
assign t[929] = t[928] ^ n[929];
assign t[930] = t[929] ^ n[930];
assign t[931] = t[930] ^ n[931];
assign t[932] = t[931] ^ n[932];
assign t[933] = t[932] ^ n[933];
assign t[934] = t[933] ^ n[934];
assign t[935] = t[934] ^ n[935];
assign t[936] = t[935] ^ n[936];
assign t[937] = t[936] ^ n[937];
assign t[938] = t[937] ^ n[938];
assign t[939] = t[938] ^ n[939];
assign t[940] = t[939] ^ n[940];
assign t[941] = t[940] ^ n[941];
assign t[942] = t[941] ^ n[942];
assign t[943] = t[942] ^ n[943];
assign t[944] = t[943] ^ n[944];
assign t[945] = t[944] ^ n[945];
assign t[946] = t[945] ^ n[946];
assign t[947] = t[946] ^ n[947];
assign t[948] = t[947] ^ n[948];
assign t[949] = t[948] ^ n[949];
assign t[950] = t[949] ^ n[950];
assign t[951] = t[950] ^ n[951];
assign t[952] = t[951] ^ n[952];
assign t[953] = t[952] ^ n[953];
assign t[954] = t[953] ^ n[954];
assign t[955] = t[954] ^ n[955];
assign t[956] = t[955] ^ n[956];
assign t[957] = t[956] ^ n[957];
assign t[958] = t[957] ^ n[958];
assign t[959] = t[958] ^ n[959];
assign t[960] = t[959] ^ n[960];
assign t[961] = t[960] ^ n[961];
assign t[962] = t[961] ^ n[962];
assign t[963] = t[962] ^ n[963];
assign t[964] = t[963] ^ n[964];
assign t[965] = t[964] ^ n[965];
assign t[966] = t[965] ^ n[966];
assign t[967] = t[966] ^ n[967];
assign t[968] = t[967] ^ n[968];
assign t[969] = t[968] ^ n[969];
assign t[970] = t[969] ^ n[970];
assign t[971] = t[970] ^ n[971];
assign t[972] = t[971] ^ n[972];
assign t[973] = t[972] ^ n[973];
assign t[974] = t[973] ^ n[974];
assign t[975] = t[974] ^ n[975];
assign t[976] = t[975] ^ n[976];
assign t[977] = t[976] ^ n[977];
assign t[978] = t[977] ^ n[978];
assign t[979] = t[978] ^ n[979];
assign t[980] = t[979] ^ n[980];
assign t[981] = t[980] ^ n[981];
assign t[982] = t[981] ^ n[982];
assign t[983] = t[982] ^ n[983];
assign t[984] = t[983] ^ n[984];
assign t[985] = t[984] ^ n[985];
assign t[986] = t[985] ^ n[986];
assign t[987] = t[986] ^ n[987];
assign t[988] = t[987] ^ n[988];
assign t[989] = t[988] ^ n[989];
assign t[990] = t[989] ^ n[990];
assign t[991] = t[990] ^ n[991];
assign t[992] = t[991] ^ n[992];
assign t[993] = t[992] ^ n[993];
assign t[994] = t[993] ^ n[994];
assign t[995] = t[994] ^ n[995];
assign t[996] = t[995] ^ n[996];
assign t[997] = t[996] ^ n[997];
assign t[998] = t[997] ^ n[998];
assign t[999] = t[998] ^ n[999];
assign t[1000] = t[999] ^ n[1000];
assign t[1001] = t[1000] ^ n[1001];
assign t[1002] = t[1001] ^ n[1002];
assign t[1003] = t[1002] ^ n[1003];
assign t[1004] = t[1003] ^ n[1004];
assign t[1005] = t[1004] ^ n[1005];
assign t[1006] = t[1005] ^ n[1006];
assign t[1007] = t[1006] ^ n[1007];
assign t[1008] = t[1007] ^ n[1008];
assign t[1009] = t[1008] ^ n[1009];
assign t[1010] = t[1009] ^ n[1010];
assign t[1011] = t[1010] ^ n[1011];
assign t[1012] = t[1011] ^ n[1012];

//asigning bit 9
assign s[9] = ( a[9] ^ b [9] ) ^ t[1012];

assign t[1013] = n[1013];
assign t[1014] = t[1013] ^ n[1014];
assign t[1015] = t[1014] ^ n[1015];
assign t[1016] = t[1015] ^ n[1016];
assign t[1017] = t[1016] ^ n[1017];
assign t[1018] = t[1017] ^ n[1018];
assign t[1019] = t[1018] ^ n[1019];
assign t[1020] = t[1019] ^ n[1020];
assign t[1021] = t[1020] ^ n[1021];
assign t[1022] = t[1021] ^ n[1022];
assign t[1023] = t[1022] ^ n[1023];
assign t[1024] = t[1023] ^ n[1024];
assign t[1025] = t[1024] ^ n[1025];
assign t[1026] = t[1025] ^ n[1026];
assign t[1027] = t[1026] ^ n[1027];
assign t[1028] = t[1027] ^ n[1028];
assign t[1029] = t[1028] ^ n[1029];
assign t[1030] = t[1029] ^ n[1030];
assign t[1031] = t[1030] ^ n[1031];
assign t[1032] = t[1031] ^ n[1032];
assign t[1033] = t[1032] ^ n[1033];
assign t[1034] = t[1033] ^ n[1034];
assign t[1035] = t[1034] ^ n[1035];
assign t[1036] = t[1035] ^ n[1036];
assign t[1037] = t[1036] ^ n[1037];
assign t[1038] = t[1037] ^ n[1038];
assign t[1039] = t[1038] ^ n[1039];
assign t[1040] = t[1039] ^ n[1040];
assign t[1041] = t[1040] ^ n[1041];
assign t[1042] = t[1041] ^ n[1042];
assign t[1043] = t[1042] ^ n[1043];
assign t[1044] = t[1043] ^ n[1044];
assign t[1045] = t[1044] ^ n[1045];
assign t[1046] = t[1045] ^ n[1046];
assign t[1047] = t[1046] ^ n[1047];
assign t[1048] = t[1047] ^ n[1048];
assign t[1049] = t[1048] ^ n[1049];
assign t[1050] = t[1049] ^ n[1050];
assign t[1051] = t[1050] ^ n[1051];
assign t[1052] = t[1051] ^ n[1052];
assign t[1053] = t[1052] ^ n[1053];
assign t[1054] = t[1053] ^ n[1054];
assign t[1055] = t[1054] ^ n[1055];
assign t[1056] = t[1055] ^ n[1056];
assign t[1057] = t[1056] ^ n[1057];
assign t[1058] = t[1057] ^ n[1058];
assign t[1059] = t[1058] ^ n[1059];
assign t[1060] = t[1059] ^ n[1060];
assign t[1061] = t[1060] ^ n[1061];
assign t[1062] = t[1061] ^ n[1062];
assign t[1063] = t[1062] ^ n[1063];
assign t[1064] = t[1063] ^ n[1064];
assign t[1065] = t[1064] ^ n[1065];
assign t[1066] = t[1065] ^ n[1066];
assign t[1067] = t[1066] ^ n[1067];
assign t[1068] = t[1067] ^ n[1068];
assign t[1069] = t[1068] ^ n[1069];
assign t[1070] = t[1069] ^ n[1070];
assign t[1071] = t[1070] ^ n[1071];
assign t[1072] = t[1071] ^ n[1072];
assign t[1073] = t[1072] ^ n[1073];
assign t[1074] = t[1073] ^ n[1074];
assign t[1075] = t[1074] ^ n[1075];
assign t[1076] = t[1075] ^ n[1076];
assign t[1077] = t[1076] ^ n[1077];
assign t[1078] = t[1077] ^ n[1078];
assign t[1079] = t[1078] ^ n[1079];
assign t[1080] = t[1079] ^ n[1080];
assign t[1081] = t[1080] ^ n[1081];
assign t[1082] = t[1081] ^ n[1082];
assign t[1083] = t[1082] ^ n[1083];
assign t[1084] = t[1083] ^ n[1084];
assign t[1085] = t[1084] ^ n[1085];
assign t[1086] = t[1085] ^ n[1086];
assign t[1087] = t[1086] ^ n[1087];
assign t[1088] = t[1087] ^ n[1088];
assign t[1089] = t[1088] ^ n[1089];
assign t[1090] = t[1089] ^ n[1090];
assign t[1091] = t[1090] ^ n[1091];
assign t[1092] = t[1091] ^ n[1092];
assign t[1093] = t[1092] ^ n[1093];
assign t[1094] = t[1093] ^ n[1094];
assign t[1095] = t[1094] ^ n[1095];
assign t[1096] = t[1095] ^ n[1096];
assign t[1097] = t[1096] ^ n[1097];
assign t[1098] = t[1097] ^ n[1098];
assign t[1099] = t[1098] ^ n[1099];
assign t[1100] = t[1099] ^ n[1100];
assign t[1101] = t[1100] ^ n[1101];
assign t[1102] = t[1101] ^ n[1102];
assign t[1103] = t[1102] ^ n[1103];
assign t[1104] = t[1103] ^ n[1104];
assign t[1105] = t[1104] ^ n[1105];
assign t[1106] = t[1105] ^ n[1106];
assign t[1107] = t[1106] ^ n[1107];
assign t[1108] = t[1107] ^ n[1108];
assign t[1109] = t[1108] ^ n[1109];
assign t[1110] = t[1109] ^ n[1110];
assign t[1111] = t[1110] ^ n[1111];
assign t[1112] = t[1111] ^ n[1112];
assign t[1113] = t[1112] ^ n[1113];
assign t[1114] = t[1113] ^ n[1114];
assign t[1115] = t[1114] ^ n[1115];
assign t[1116] = t[1115] ^ n[1116];
assign t[1117] = t[1116] ^ n[1117];
assign t[1118] = t[1117] ^ n[1118];
assign t[1119] = t[1118] ^ n[1119];
assign t[1120] = t[1119] ^ n[1120];
assign t[1121] = t[1120] ^ n[1121];
assign t[1122] = t[1121] ^ n[1122];
assign t[1123] = t[1122] ^ n[1123];
assign t[1124] = t[1123] ^ n[1124];
assign t[1125] = t[1124] ^ n[1125];
assign t[1126] = t[1125] ^ n[1126];
assign t[1127] = t[1126] ^ n[1127];
assign t[1128] = t[1127] ^ n[1128];
assign t[1129] = t[1128] ^ n[1129];
assign t[1130] = t[1129] ^ n[1130];
assign t[1131] = t[1130] ^ n[1131];
assign t[1132] = t[1131] ^ n[1132];
assign t[1133] = t[1132] ^ n[1133];
assign t[1134] = t[1133] ^ n[1134];
assign t[1135] = t[1134] ^ n[1135];
assign t[1136] = t[1135] ^ n[1136];
assign t[1137] = t[1136] ^ n[1137];
assign t[1138] = t[1137] ^ n[1138];
assign t[1139] = t[1138] ^ n[1139];
assign t[1140] = t[1139] ^ n[1140];
assign t[1141] = t[1140] ^ n[1141];
assign t[1142] = t[1141] ^ n[1142];
assign t[1143] = t[1142] ^ n[1143];
assign t[1144] = t[1143] ^ n[1144];
assign t[1145] = t[1144] ^ n[1145];
assign t[1146] = t[1145] ^ n[1146];
assign t[1147] = t[1146] ^ n[1147];
assign t[1148] = t[1147] ^ n[1148];
assign t[1149] = t[1148] ^ n[1149];
assign t[1150] = t[1149] ^ n[1150];
assign t[1151] = t[1150] ^ n[1151];
assign t[1152] = t[1151] ^ n[1152];
assign t[1153] = t[1152] ^ n[1153];
assign t[1154] = t[1153] ^ n[1154];
assign t[1155] = t[1154] ^ n[1155];
assign t[1156] = t[1155] ^ n[1156];
assign t[1157] = t[1156] ^ n[1157];
assign t[1158] = t[1157] ^ n[1158];
assign t[1159] = t[1158] ^ n[1159];
assign t[1160] = t[1159] ^ n[1160];
assign t[1161] = t[1160] ^ n[1161];
assign t[1162] = t[1161] ^ n[1162];
assign t[1163] = t[1162] ^ n[1163];
assign t[1164] = t[1163] ^ n[1164];
assign t[1165] = t[1164] ^ n[1165];
assign t[1166] = t[1165] ^ n[1166];
assign t[1167] = t[1166] ^ n[1167];
assign t[1168] = t[1167] ^ n[1168];
assign t[1169] = t[1168] ^ n[1169];
assign t[1170] = t[1169] ^ n[1170];
assign t[1171] = t[1170] ^ n[1171];
assign t[1172] = t[1171] ^ n[1172];
assign t[1173] = t[1172] ^ n[1173];
assign t[1174] = t[1173] ^ n[1174];
assign t[1175] = t[1174] ^ n[1175];
assign t[1176] = t[1175] ^ n[1176];
assign t[1177] = t[1176] ^ n[1177];
assign t[1178] = t[1177] ^ n[1178];
assign t[1179] = t[1178] ^ n[1179];
assign t[1180] = t[1179] ^ n[1180];
assign t[1181] = t[1180] ^ n[1181];
assign t[1182] = t[1181] ^ n[1182];
assign t[1183] = t[1182] ^ n[1183];
assign t[1184] = t[1183] ^ n[1184];
assign t[1185] = t[1184] ^ n[1185];
assign t[1186] = t[1185] ^ n[1186];
assign t[1187] = t[1186] ^ n[1187];
assign t[1188] = t[1187] ^ n[1188];
assign t[1189] = t[1188] ^ n[1189];
assign t[1190] = t[1189] ^ n[1190];
assign t[1191] = t[1190] ^ n[1191];
assign t[1192] = t[1191] ^ n[1192];
assign t[1193] = t[1192] ^ n[1193];
assign t[1194] = t[1193] ^ n[1194];
assign t[1195] = t[1194] ^ n[1195];
assign t[1196] = t[1195] ^ n[1196];
assign t[1197] = t[1196] ^ n[1197];
assign t[1198] = t[1197] ^ n[1198];
assign t[1199] = t[1198] ^ n[1199];
assign t[1200] = t[1199] ^ n[1200];
assign t[1201] = t[1200] ^ n[1201];
assign t[1202] = t[1201] ^ n[1202];
assign t[1203] = t[1202] ^ n[1203];
assign t[1204] = t[1203] ^ n[1204];
assign t[1205] = t[1204] ^ n[1205];
assign t[1206] = t[1205] ^ n[1206];
assign t[1207] = t[1206] ^ n[1207];
assign t[1208] = t[1207] ^ n[1208];
assign t[1209] = t[1208] ^ n[1209];
assign t[1210] = t[1209] ^ n[1210];
assign t[1211] = t[1210] ^ n[1211];
assign t[1212] = t[1211] ^ n[1212];
assign t[1213] = t[1212] ^ n[1213];
assign t[1214] = t[1213] ^ n[1214];
assign t[1215] = t[1214] ^ n[1215];
assign t[1216] = t[1215] ^ n[1216];
assign t[1217] = t[1216] ^ n[1217];
assign t[1218] = t[1217] ^ n[1218];
assign t[1219] = t[1218] ^ n[1219];
assign t[1220] = t[1219] ^ n[1220];
assign t[1221] = t[1220] ^ n[1221];
assign t[1222] = t[1221] ^ n[1222];
assign t[1223] = t[1222] ^ n[1223];
assign t[1224] = t[1223] ^ n[1224];
assign t[1225] = t[1224] ^ n[1225];
assign t[1226] = t[1225] ^ n[1226];
assign t[1227] = t[1226] ^ n[1227];
assign t[1228] = t[1227] ^ n[1228];
assign t[1229] = t[1228] ^ n[1229];
assign t[1230] = t[1229] ^ n[1230];
assign t[1231] = t[1230] ^ n[1231];
assign t[1232] = t[1231] ^ n[1232];
assign t[1233] = t[1232] ^ n[1233];
assign t[1234] = t[1233] ^ n[1234];
assign t[1235] = t[1234] ^ n[1235];
assign t[1236] = t[1235] ^ n[1236];
assign t[1237] = t[1236] ^ n[1237];
assign t[1238] = t[1237] ^ n[1238];
assign t[1239] = t[1238] ^ n[1239];
assign t[1240] = t[1239] ^ n[1240];
assign t[1241] = t[1240] ^ n[1241];
assign t[1242] = t[1241] ^ n[1242];
assign t[1243] = t[1242] ^ n[1243];
assign t[1244] = t[1243] ^ n[1244];
assign t[1245] = t[1244] ^ n[1245];
assign t[1246] = t[1245] ^ n[1246];
assign t[1247] = t[1246] ^ n[1247];
assign t[1248] = t[1247] ^ n[1248];
assign t[1249] = t[1248] ^ n[1249];
assign t[1250] = t[1249] ^ n[1250];
assign t[1251] = t[1250] ^ n[1251];
assign t[1252] = t[1251] ^ n[1252];
assign t[1253] = t[1252] ^ n[1253];
assign t[1254] = t[1253] ^ n[1254];
assign t[1255] = t[1254] ^ n[1255];
assign t[1256] = t[1255] ^ n[1256];
assign t[1257] = t[1256] ^ n[1257];
assign t[1258] = t[1257] ^ n[1258];
assign t[1259] = t[1258] ^ n[1259];
assign t[1260] = t[1259] ^ n[1260];
assign t[1261] = t[1260] ^ n[1261];
assign t[1262] = t[1261] ^ n[1262];
assign t[1263] = t[1262] ^ n[1263];
assign t[1264] = t[1263] ^ n[1264];
assign t[1265] = t[1264] ^ n[1265];
assign t[1266] = t[1265] ^ n[1266];
assign t[1267] = t[1266] ^ n[1267];
assign t[1268] = t[1267] ^ n[1268];
assign t[1269] = t[1268] ^ n[1269];
assign t[1270] = t[1269] ^ n[1270];
assign t[1271] = t[1270] ^ n[1271];
assign t[1272] = t[1271] ^ n[1272];
assign t[1273] = t[1272] ^ n[1273];
assign t[1274] = t[1273] ^ n[1274];
assign t[1275] = t[1274] ^ n[1275];
assign t[1276] = t[1275] ^ n[1276];
assign t[1277] = t[1276] ^ n[1277];
assign t[1278] = t[1277] ^ n[1278];
assign t[1279] = t[1278] ^ n[1279];
assign t[1280] = t[1279] ^ n[1280];
assign t[1281] = t[1280] ^ n[1281];
assign t[1282] = t[1281] ^ n[1282];
assign t[1283] = t[1282] ^ n[1283];
assign t[1284] = t[1283] ^ n[1284];
assign t[1285] = t[1284] ^ n[1285];
assign t[1286] = t[1285] ^ n[1286];
assign t[1287] = t[1286] ^ n[1287];
assign t[1288] = t[1287] ^ n[1288];
assign t[1289] = t[1288] ^ n[1289];
assign t[1290] = t[1289] ^ n[1290];
assign t[1291] = t[1290] ^ n[1291];
assign t[1292] = t[1291] ^ n[1292];
assign t[1293] = t[1292] ^ n[1293];
assign t[1294] = t[1293] ^ n[1294];
assign t[1295] = t[1294] ^ n[1295];
assign t[1296] = t[1295] ^ n[1296];
assign t[1297] = t[1296] ^ n[1297];
assign t[1298] = t[1297] ^ n[1298];
assign t[1299] = t[1298] ^ n[1299];
assign t[1300] = t[1299] ^ n[1300];
assign t[1301] = t[1300] ^ n[1301];
assign t[1302] = t[1301] ^ n[1302];
assign t[1303] = t[1302] ^ n[1303];
assign t[1304] = t[1303] ^ n[1304];
assign t[1305] = t[1304] ^ n[1305];
assign t[1306] = t[1305] ^ n[1306];
assign t[1307] = t[1306] ^ n[1307];
assign t[1308] = t[1307] ^ n[1308];
assign t[1309] = t[1308] ^ n[1309];
assign t[1310] = t[1309] ^ n[1310];
assign t[1311] = t[1310] ^ n[1311];
assign t[1312] = t[1311] ^ n[1312];
assign t[1313] = t[1312] ^ n[1313];
assign t[1314] = t[1313] ^ n[1314];
assign t[1315] = t[1314] ^ n[1315];
assign t[1316] = t[1315] ^ n[1316];
assign t[1317] = t[1316] ^ n[1317];
assign t[1318] = t[1317] ^ n[1318];
assign t[1319] = t[1318] ^ n[1319];
assign t[1320] = t[1319] ^ n[1320];
assign t[1321] = t[1320] ^ n[1321];
assign t[1322] = t[1321] ^ n[1322];
assign t[1323] = t[1322] ^ n[1323];
assign t[1324] = t[1323] ^ n[1324];
assign t[1325] = t[1324] ^ n[1325];
assign t[1326] = t[1325] ^ n[1326];
assign t[1327] = t[1326] ^ n[1327];
assign t[1328] = t[1327] ^ n[1328];
assign t[1329] = t[1328] ^ n[1329];
assign t[1330] = t[1329] ^ n[1330];
assign t[1331] = t[1330] ^ n[1331];
assign t[1332] = t[1331] ^ n[1332];
assign t[1333] = t[1332] ^ n[1333];
assign t[1334] = t[1333] ^ n[1334];
assign t[1335] = t[1334] ^ n[1335];
assign t[1336] = t[1335] ^ n[1336];
assign t[1337] = t[1336] ^ n[1337];
assign t[1338] = t[1337] ^ n[1338];
assign t[1339] = t[1338] ^ n[1339];
assign t[1340] = t[1339] ^ n[1340];
assign t[1341] = t[1340] ^ n[1341];
assign t[1342] = t[1341] ^ n[1342];
assign t[1343] = t[1342] ^ n[1343];
assign t[1344] = t[1343] ^ n[1344];
assign t[1345] = t[1344] ^ n[1345];
assign t[1346] = t[1345] ^ n[1346];
assign t[1347] = t[1346] ^ n[1347];
assign t[1348] = t[1347] ^ n[1348];
assign t[1349] = t[1348] ^ n[1349];
assign t[1350] = t[1349] ^ n[1350];
assign t[1351] = t[1350] ^ n[1351];
assign t[1352] = t[1351] ^ n[1352];
assign t[1353] = t[1352] ^ n[1353];
assign t[1354] = t[1353] ^ n[1354];
assign t[1355] = t[1354] ^ n[1355];
assign t[1356] = t[1355] ^ n[1356];
assign t[1357] = t[1356] ^ n[1357];
assign t[1358] = t[1357] ^ n[1358];
assign t[1359] = t[1358] ^ n[1359];
assign t[1360] = t[1359] ^ n[1360];
assign t[1361] = t[1360] ^ n[1361];
assign t[1362] = t[1361] ^ n[1362];
assign t[1363] = t[1362] ^ n[1363];
assign t[1364] = t[1363] ^ n[1364];
assign t[1365] = t[1364] ^ n[1365];
assign t[1366] = t[1365] ^ n[1366];
assign t[1367] = t[1366] ^ n[1367];
assign t[1368] = t[1367] ^ n[1368];
assign t[1369] = t[1368] ^ n[1369];
assign t[1370] = t[1369] ^ n[1370];
assign t[1371] = t[1370] ^ n[1371];
assign t[1372] = t[1371] ^ n[1372];
assign t[1373] = t[1372] ^ n[1373];
assign t[1374] = t[1373] ^ n[1374];
assign t[1375] = t[1374] ^ n[1375];
assign t[1376] = t[1375] ^ n[1376];
assign t[1377] = t[1376] ^ n[1377];
assign t[1378] = t[1377] ^ n[1378];
assign t[1379] = t[1378] ^ n[1379];
assign t[1380] = t[1379] ^ n[1380];
assign t[1381] = t[1380] ^ n[1381];
assign t[1382] = t[1381] ^ n[1382];
assign t[1383] = t[1382] ^ n[1383];
assign t[1384] = t[1383] ^ n[1384];
assign t[1385] = t[1384] ^ n[1385];
assign t[1386] = t[1385] ^ n[1386];
assign t[1387] = t[1386] ^ n[1387];
assign t[1388] = t[1387] ^ n[1388];
assign t[1389] = t[1388] ^ n[1389];
assign t[1390] = t[1389] ^ n[1390];
assign t[1391] = t[1390] ^ n[1391];
assign t[1392] = t[1391] ^ n[1392];
assign t[1393] = t[1392] ^ n[1393];
assign t[1394] = t[1393] ^ n[1394];
assign t[1395] = t[1394] ^ n[1395];
assign t[1396] = t[1395] ^ n[1396];
assign t[1397] = t[1396] ^ n[1397];
assign t[1398] = t[1397] ^ n[1398];
assign t[1399] = t[1398] ^ n[1399];
assign t[1400] = t[1399] ^ n[1400];
assign t[1401] = t[1400] ^ n[1401];
assign t[1402] = t[1401] ^ n[1402];
assign t[1403] = t[1402] ^ n[1403];
assign t[1404] = t[1403] ^ n[1404];
assign t[1405] = t[1404] ^ n[1405];
assign t[1406] = t[1405] ^ n[1406];
assign t[1407] = t[1406] ^ n[1407];
assign t[1408] = t[1407] ^ n[1408];
assign t[1409] = t[1408] ^ n[1409];
assign t[1410] = t[1409] ^ n[1410];
assign t[1411] = t[1410] ^ n[1411];
assign t[1412] = t[1411] ^ n[1412];
assign t[1413] = t[1412] ^ n[1413];
assign t[1414] = t[1413] ^ n[1414];
assign t[1415] = t[1414] ^ n[1415];
assign t[1416] = t[1415] ^ n[1416];
assign t[1417] = t[1416] ^ n[1417];
assign t[1418] = t[1417] ^ n[1418];
assign t[1419] = t[1418] ^ n[1419];
assign t[1420] = t[1419] ^ n[1420];
assign t[1421] = t[1420] ^ n[1421];
assign t[1422] = t[1421] ^ n[1422];
assign t[1423] = t[1422] ^ n[1423];
assign t[1424] = t[1423] ^ n[1424];
assign t[1425] = t[1424] ^ n[1425];
assign t[1426] = t[1425] ^ n[1426];
assign t[1427] = t[1426] ^ n[1427];
assign t[1428] = t[1427] ^ n[1428];
assign t[1429] = t[1428] ^ n[1429];
assign t[1430] = t[1429] ^ n[1430];
assign t[1431] = t[1430] ^ n[1431];
assign t[1432] = t[1431] ^ n[1432];
assign t[1433] = t[1432] ^ n[1433];
assign t[1434] = t[1433] ^ n[1434];
assign t[1435] = t[1434] ^ n[1435];
assign t[1436] = t[1435] ^ n[1436];
assign t[1437] = t[1436] ^ n[1437];
assign t[1438] = t[1437] ^ n[1438];
assign t[1439] = t[1438] ^ n[1439];
assign t[1440] = t[1439] ^ n[1440];
assign t[1441] = t[1440] ^ n[1441];
assign t[1442] = t[1441] ^ n[1442];
assign t[1443] = t[1442] ^ n[1443];
assign t[1444] = t[1443] ^ n[1444];
assign t[1445] = t[1444] ^ n[1445];
assign t[1446] = t[1445] ^ n[1446];
assign t[1447] = t[1446] ^ n[1447];
assign t[1448] = t[1447] ^ n[1448];
assign t[1449] = t[1448] ^ n[1449];
assign t[1450] = t[1449] ^ n[1450];
assign t[1451] = t[1450] ^ n[1451];
assign t[1452] = t[1451] ^ n[1452];
assign t[1453] = t[1452] ^ n[1453];
assign t[1454] = t[1453] ^ n[1454];
assign t[1455] = t[1454] ^ n[1455];
assign t[1456] = t[1455] ^ n[1456];
assign t[1457] = t[1456] ^ n[1457];
assign t[1458] = t[1457] ^ n[1458];
assign t[1459] = t[1458] ^ n[1459];
assign t[1460] = t[1459] ^ n[1460];
assign t[1461] = t[1460] ^ n[1461];
assign t[1462] = t[1461] ^ n[1462];
assign t[1463] = t[1462] ^ n[1463];
assign t[1464] = t[1463] ^ n[1464];
assign t[1465] = t[1464] ^ n[1465];
assign t[1466] = t[1465] ^ n[1466];
assign t[1467] = t[1466] ^ n[1467];
assign t[1468] = t[1467] ^ n[1468];
assign t[1469] = t[1468] ^ n[1469];
assign t[1470] = t[1469] ^ n[1470];
assign t[1471] = t[1470] ^ n[1471];
assign t[1472] = t[1471] ^ n[1472];
assign t[1473] = t[1472] ^ n[1473];
assign t[1474] = t[1473] ^ n[1474];
assign t[1475] = t[1474] ^ n[1475];
assign t[1476] = t[1475] ^ n[1476];
assign t[1477] = t[1476] ^ n[1477];
assign t[1478] = t[1477] ^ n[1478];
assign t[1479] = t[1478] ^ n[1479];
assign t[1480] = t[1479] ^ n[1480];
assign t[1481] = t[1480] ^ n[1481];
assign t[1482] = t[1481] ^ n[1482];
assign t[1483] = t[1482] ^ n[1483];
assign t[1484] = t[1483] ^ n[1484];
assign t[1485] = t[1484] ^ n[1485];
assign t[1486] = t[1485] ^ n[1486];
assign t[1487] = t[1486] ^ n[1487];
assign t[1488] = t[1487] ^ n[1488];
assign t[1489] = t[1488] ^ n[1489];
assign t[1490] = t[1489] ^ n[1490];
assign t[1491] = t[1490] ^ n[1491];
assign t[1492] = t[1491] ^ n[1492];
assign t[1493] = t[1492] ^ n[1493];
assign t[1494] = t[1493] ^ n[1494];
assign t[1495] = t[1494] ^ n[1495];
assign t[1496] = t[1495] ^ n[1496];
assign t[1497] = t[1496] ^ n[1497];
assign t[1498] = t[1497] ^ n[1498];
assign t[1499] = t[1498] ^ n[1499];
assign t[1500] = t[1499] ^ n[1500];
assign t[1501] = t[1500] ^ n[1501];
assign t[1502] = t[1501] ^ n[1502];
assign t[1503] = t[1502] ^ n[1503];
assign t[1504] = t[1503] ^ n[1504];
assign t[1505] = t[1504] ^ n[1505];
assign t[1506] = t[1505] ^ n[1506];
assign t[1507] = t[1506] ^ n[1507];
assign t[1508] = t[1507] ^ n[1508];
assign t[1509] = t[1508] ^ n[1509];
assign t[1510] = t[1509] ^ n[1510];
assign t[1511] = t[1510] ^ n[1511];
assign t[1512] = t[1511] ^ n[1512];
assign t[1513] = t[1512] ^ n[1513];
assign t[1514] = t[1513] ^ n[1514];
assign t[1515] = t[1514] ^ n[1515];
assign t[1516] = t[1515] ^ n[1516];
assign t[1517] = t[1516] ^ n[1517];
assign t[1518] = t[1517] ^ n[1518];
assign t[1519] = t[1518] ^ n[1519];
assign t[1520] = t[1519] ^ n[1520];
assign t[1521] = t[1520] ^ n[1521];
assign t[1522] = t[1521] ^ n[1522];
assign t[1523] = t[1522] ^ n[1523];
assign t[1524] = t[1523] ^ n[1524];
assign t[1525] = t[1524] ^ n[1525];
assign t[1526] = t[1525] ^ n[1526];
assign t[1527] = t[1526] ^ n[1527];
assign t[1528] = t[1527] ^ n[1528];
assign t[1529] = t[1528] ^ n[1529];
assign t[1530] = t[1529] ^ n[1530];
assign t[1531] = t[1530] ^ n[1531];
assign t[1532] = t[1531] ^ n[1532];
assign t[1533] = t[1532] ^ n[1533];
assign t[1534] = t[1533] ^ n[1534];
assign t[1535] = t[1534] ^ n[1535];
assign t[1536] = t[1535] ^ n[1536];
assign t[1537] = t[1536] ^ n[1537];
assign t[1538] = t[1537] ^ n[1538];
assign t[1539] = t[1538] ^ n[1539];
assign t[1540] = t[1539] ^ n[1540];
assign t[1541] = t[1540] ^ n[1541];
assign t[1542] = t[1541] ^ n[1542];
assign t[1543] = t[1542] ^ n[1543];
assign t[1544] = t[1543] ^ n[1544];
assign t[1545] = t[1544] ^ n[1545];
assign t[1546] = t[1545] ^ n[1546];
assign t[1547] = t[1546] ^ n[1547];
assign t[1548] = t[1547] ^ n[1548];
assign t[1549] = t[1548] ^ n[1549];
assign t[1550] = t[1549] ^ n[1550];
assign t[1551] = t[1550] ^ n[1551];
assign t[1552] = t[1551] ^ n[1552];
assign t[1553] = t[1552] ^ n[1553];
assign t[1554] = t[1553] ^ n[1554];
assign t[1555] = t[1554] ^ n[1555];
assign t[1556] = t[1555] ^ n[1556];
assign t[1557] = t[1556] ^ n[1557];
assign t[1558] = t[1557] ^ n[1558];
assign t[1559] = t[1558] ^ n[1559];
assign t[1560] = t[1559] ^ n[1560];
assign t[1561] = t[1560] ^ n[1561];
assign t[1562] = t[1561] ^ n[1562];
assign t[1563] = t[1562] ^ n[1563];
assign t[1564] = t[1563] ^ n[1564];
assign t[1565] = t[1564] ^ n[1565];
assign t[1566] = t[1565] ^ n[1566];
assign t[1567] = t[1566] ^ n[1567];
assign t[1568] = t[1567] ^ n[1568];
assign t[1569] = t[1568] ^ n[1569];
assign t[1570] = t[1569] ^ n[1570];
assign t[1571] = t[1570] ^ n[1571];
assign t[1572] = t[1571] ^ n[1572];
assign t[1573] = t[1572] ^ n[1573];
assign t[1574] = t[1573] ^ n[1574];
assign t[1575] = t[1574] ^ n[1575];
assign t[1576] = t[1575] ^ n[1576];
assign t[1577] = t[1576] ^ n[1577];
assign t[1578] = t[1577] ^ n[1578];
assign t[1579] = t[1578] ^ n[1579];
assign t[1580] = t[1579] ^ n[1580];
assign t[1581] = t[1580] ^ n[1581];
assign t[1582] = t[1581] ^ n[1582];
assign t[1583] = t[1582] ^ n[1583];
assign t[1584] = t[1583] ^ n[1584];
assign t[1585] = t[1584] ^ n[1585];
assign t[1586] = t[1585] ^ n[1586];
assign t[1587] = t[1586] ^ n[1587];
assign t[1588] = t[1587] ^ n[1588];
assign t[1589] = t[1588] ^ n[1589];
assign t[1590] = t[1589] ^ n[1590];
assign t[1591] = t[1590] ^ n[1591];
assign t[1592] = t[1591] ^ n[1592];
assign t[1593] = t[1592] ^ n[1593];
assign t[1594] = t[1593] ^ n[1594];
assign t[1595] = t[1594] ^ n[1595];
assign t[1596] = t[1595] ^ n[1596];
assign t[1597] = t[1596] ^ n[1597];
assign t[1598] = t[1597] ^ n[1598];
assign t[1599] = t[1598] ^ n[1599];
assign t[1600] = t[1599] ^ n[1600];
assign t[1601] = t[1600] ^ n[1601];
assign t[1602] = t[1601] ^ n[1602];
assign t[1603] = t[1602] ^ n[1603];
assign t[1604] = t[1603] ^ n[1604];
assign t[1605] = t[1604] ^ n[1605];
assign t[1606] = t[1605] ^ n[1606];
assign t[1607] = t[1606] ^ n[1607];
assign t[1608] = t[1607] ^ n[1608];
assign t[1609] = t[1608] ^ n[1609];
assign t[1610] = t[1609] ^ n[1610];
assign t[1611] = t[1610] ^ n[1611];
assign t[1612] = t[1611] ^ n[1612];
assign t[1613] = t[1612] ^ n[1613];
assign t[1614] = t[1613] ^ n[1614];
assign t[1615] = t[1614] ^ n[1615];
assign t[1616] = t[1615] ^ n[1616];
assign t[1617] = t[1616] ^ n[1617];
assign t[1618] = t[1617] ^ n[1618];
assign t[1619] = t[1618] ^ n[1619];
assign t[1620] = t[1619] ^ n[1620];
assign t[1621] = t[1620] ^ n[1621];
assign t[1622] = t[1621] ^ n[1622];
assign t[1623] = t[1622] ^ n[1623];
assign t[1624] = t[1623] ^ n[1624];
assign t[1625] = t[1624] ^ n[1625];
assign t[1626] = t[1625] ^ n[1626];
assign t[1627] = t[1626] ^ n[1627];
assign t[1628] = t[1627] ^ n[1628];
assign t[1629] = t[1628] ^ n[1629];
assign t[1630] = t[1629] ^ n[1630];
assign t[1631] = t[1630] ^ n[1631];
assign t[1632] = t[1631] ^ n[1632];
assign t[1633] = t[1632] ^ n[1633];
assign t[1634] = t[1633] ^ n[1634];
assign t[1635] = t[1634] ^ n[1635];
assign t[1636] = t[1635] ^ n[1636];
assign t[1637] = t[1636] ^ n[1637];
assign t[1638] = t[1637] ^ n[1638];
assign t[1639] = t[1638] ^ n[1639];
assign t[1640] = t[1639] ^ n[1640];
assign t[1641] = t[1640] ^ n[1641];
assign t[1642] = t[1641] ^ n[1642];
assign t[1643] = t[1642] ^ n[1643];
assign t[1644] = t[1643] ^ n[1644];
assign t[1645] = t[1644] ^ n[1645];
assign t[1646] = t[1645] ^ n[1646];
assign t[1647] = t[1646] ^ n[1647];
assign t[1648] = t[1647] ^ n[1648];
assign t[1649] = t[1648] ^ n[1649];
assign t[1650] = t[1649] ^ n[1650];
assign t[1651] = t[1650] ^ n[1651];
assign t[1652] = t[1651] ^ n[1652];
assign t[1653] = t[1652] ^ n[1653];
assign t[1654] = t[1653] ^ n[1654];
assign t[1655] = t[1654] ^ n[1655];
assign t[1656] = t[1655] ^ n[1656];
assign t[1657] = t[1656] ^ n[1657];
assign t[1658] = t[1657] ^ n[1658];
assign t[1659] = t[1658] ^ n[1659];
assign t[1660] = t[1659] ^ n[1660];
assign t[1661] = t[1660] ^ n[1661];
assign t[1662] = t[1661] ^ n[1662];
assign t[1663] = t[1662] ^ n[1663];
assign t[1664] = t[1663] ^ n[1664];
assign t[1665] = t[1664] ^ n[1665];
assign t[1666] = t[1665] ^ n[1666];
assign t[1667] = t[1666] ^ n[1667];
assign t[1668] = t[1667] ^ n[1668];
assign t[1669] = t[1668] ^ n[1669];
assign t[1670] = t[1669] ^ n[1670];
assign t[1671] = t[1670] ^ n[1671];
assign t[1672] = t[1671] ^ n[1672];
assign t[1673] = t[1672] ^ n[1673];
assign t[1674] = t[1673] ^ n[1674];
assign t[1675] = t[1674] ^ n[1675];
assign t[1676] = t[1675] ^ n[1676];
assign t[1677] = t[1676] ^ n[1677];
assign t[1678] = t[1677] ^ n[1678];
assign t[1679] = t[1678] ^ n[1679];
assign t[1680] = t[1679] ^ n[1680];
assign t[1681] = t[1680] ^ n[1681];
assign t[1682] = t[1681] ^ n[1682];
assign t[1683] = t[1682] ^ n[1683];
assign t[1684] = t[1683] ^ n[1684];
assign t[1685] = t[1684] ^ n[1685];
assign t[1686] = t[1685] ^ n[1686];
assign t[1687] = t[1686] ^ n[1687];
assign t[1688] = t[1687] ^ n[1688];
assign t[1689] = t[1688] ^ n[1689];
assign t[1690] = t[1689] ^ n[1690];
assign t[1691] = t[1690] ^ n[1691];
assign t[1692] = t[1691] ^ n[1692];
assign t[1693] = t[1692] ^ n[1693];
assign t[1694] = t[1693] ^ n[1694];
assign t[1695] = t[1694] ^ n[1695];
assign t[1696] = t[1695] ^ n[1696];
assign t[1697] = t[1696] ^ n[1697];
assign t[1698] = t[1697] ^ n[1698];
assign t[1699] = t[1698] ^ n[1699];
assign t[1700] = t[1699] ^ n[1700];
assign t[1701] = t[1700] ^ n[1701];
assign t[1702] = t[1701] ^ n[1702];
assign t[1703] = t[1702] ^ n[1703];
assign t[1704] = t[1703] ^ n[1704];
assign t[1705] = t[1704] ^ n[1705];
assign t[1706] = t[1705] ^ n[1706];
assign t[1707] = t[1706] ^ n[1707];
assign t[1708] = t[1707] ^ n[1708];
assign t[1709] = t[1708] ^ n[1709];
assign t[1710] = t[1709] ^ n[1710];
assign t[1711] = t[1710] ^ n[1711];
assign t[1712] = t[1711] ^ n[1712];
assign t[1713] = t[1712] ^ n[1713];
assign t[1714] = t[1713] ^ n[1714];
assign t[1715] = t[1714] ^ n[1715];
assign t[1716] = t[1715] ^ n[1716];
assign t[1717] = t[1716] ^ n[1717];
assign t[1718] = t[1717] ^ n[1718];
assign t[1719] = t[1718] ^ n[1719];
assign t[1720] = t[1719] ^ n[1720];
assign t[1721] = t[1720] ^ n[1721];
assign t[1722] = t[1721] ^ n[1722];
assign t[1723] = t[1722] ^ n[1723];
assign t[1724] = t[1723] ^ n[1724];
assign t[1725] = t[1724] ^ n[1725];
assign t[1726] = t[1725] ^ n[1726];
assign t[1727] = t[1726] ^ n[1727];
assign t[1728] = t[1727] ^ n[1728];
assign t[1729] = t[1728] ^ n[1729];
assign t[1730] = t[1729] ^ n[1730];
assign t[1731] = t[1730] ^ n[1731];
assign t[1732] = t[1731] ^ n[1732];
assign t[1733] = t[1732] ^ n[1733];
assign t[1734] = t[1733] ^ n[1734];
assign t[1735] = t[1734] ^ n[1735];
assign t[1736] = t[1735] ^ n[1736];
assign t[1737] = t[1736] ^ n[1737];
assign t[1738] = t[1737] ^ n[1738];
assign t[1739] = t[1738] ^ n[1739];
assign t[1740] = t[1739] ^ n[1740];
assign t[1741] = t[1740] ^ n[1741];
assign t[1742] = t[1741] ^ n[1742];
assign t[1743] = t[1742] ^ n[1743];
assign t[1744] = t[1743] ^ n[1744];
assign t[1745] = t[1744] ^ n[1745];
assign t[1746] = t[1745] ^ n[1746];
assign t[1747] = t[1746] ^ n[1747];
assign t[1748] = t[1747] ^ n[1748];
assign t[1749] = t[1748] ^ n[1749];
assign t[1750] = t[1749] ^ n[1750];
assign t[1751] = t[1750] ^ n[1751];
assign t[1752] = t[1751] ^ n[1752];
assign t[1753] = t[1752] ^ n[1753];
assign t[1754] = t[1753] ^ n[1754];
assign t[1755] = t[1754] ^ n[1755];
assign t[1756] = t[1755] ^ n[1756];
assign t[1757] = t[1756] ^ n[1757];
assign t[1758] = t[1757] ^ n[1758];
assign t[1759] = t[1758] ^ n[1759];
assign t[1760] = t[1759] ^ n[1760];
assign t[1761] = t[1760] ^ n[1761];
assign t[1762] = t[1761] ^ n[1762];
assign t[1763] = t[1762] ^ n[1763];
assign t[1764] = t[1763] ^ n[1764];
assign t[1765] = t[1764] ^ n[1765];
assign t[1766] = t[1765] ^ n[1766];
assign t[1767] = t[1766] ^ n[1767];
assign t[1768] = t[1767] ^ n[1768];
assign t[1769] = t[1768] ^ n[1769];
assign t[1770] = t[1769] ^ n[1770];
assign t[1771] = t[1770] ^ n[1771];
assign t[1772] = t[1771] ^ n[1772];
assign t[1773] = t[1772] ^ n[1773];
assign t[1774] = t[1773] ^ n[1774];
assign t[1775] = t[1774] ^ n[1775];
assign t[1776] = t[1775] ^ n[1776];
assign t[1777] = t[1776] ^ n[1777];
assign t[1778] = t[1777] ^ n[1778];
assign t[1779] = t[1778] ^ n[1779];
assign t[1780] = t[1779] ^ n[1780];
assign t[1781] = t[1780] ^ n[1781];
assign t[1782] = t[1781] ^ n[1782];
assign t[1783] = t[1782] ^ n[1783];
assign t[1784] = t[1783] ^ n[1784];
assign t[1785] = t[1784] ^ n[1785];
assign t[1786] = t[1785] ^ n[1786];
assign t[1787] = t[1786] ^ n[1787];
assign t[1788] = t[1787] ^ n[1788];
assign t[1789] = t[1788] ^ n[1789];
assign t[1790] = t[1789] ^ n[1790];
assign t[1791] = t[1790] ^ n[1791];
assign t[1792] = t[1791] ^ n[1792];
assign t[1793] = t[1792] ^ n[1793];
assign t[1794] = t[1793] ^ n[1794];
assign t[1795] = t[1794] ^ n[1795];
assign t[1796] = t[1795] ^ n[1796];
assign t[1797] = t[1796] ^ n[1797];
assign t[1798] = t[1797] ^ n[1798];
assign t[1799] = t[1798] ^ n[1799];
assign t[1800] = t[1799] ^ n[1800];
assign t[1801] = t[1800] ^ n[1801];
assign t[1802] = t[1801] ^ n[1802];
assign t[1803] = t[1802] ^ n[1803];
assign t[1804] = t[1803] ^ n[1804];
assign t[1805] = t[1804] ^ n[1805];
assign t[1806] = t[1805] ^ n[1806];
assign t[1807] = t[1806] ^ n[1807];
assign t[1808] = t[1807] ^ n[1808];
assign t[1809] = t[1808] ^ n[1809];
assign t[1810] = t[1809] ^ n[1810];
assign t[1811] = t[1810] ^ n[1811];
assign t[1812] = t[1811] ^ n[1812];
assign t[1813] = t[1812] ^ n[1813];
assign t[1814] = t[1813] ^ n[1814];
assign t[1815] = t[1814] ^ n[1815];
assign t[1816] = t[1815] ^ n[1816];
assign t[1817] = t[1816] ^ n[1817];
assign t[1818] = t[1817] ^ n[1818];
assign t[1819] = t[1818] ^ n[1819];
assign t[1820] = t[1819] ^ n[1820];
assign t[1821] = t[1820] ^ n[1821];
assign t[1822] = t[1821] ^ n[1822];
assign t[1823] = t[1822] ^ n[1823];
assign t[1824] = t[1823] ^ n[1824];
assign t[1825] = t[1824] ^ n[1825];
assign t[1826] = t[1825] ^ n[1826];
assign t[1827] = t[1826] ^ n[1827];
assign t[1828] = t[1827] ^ n[1828];
assign t[1829] = t[1828] ^ n[1829];
assign t[1830] = t[1829] ^ n[1830];
assign t[1831] = t[1830] ^ n[1831];
assign t[1832] = t[1831] ^ n[1832];
assign t[1833] = t[1832] ^ n[1833];
assign t[1834] = t[1833] ^ n[1834];
assign t[1835] = t[1834] ^ n[1835];
assign t[1836] = t[1835] ^ n[1836];
assign t[1837] = t[1836] ^ n[1837];
assign t[1838] = t[1837] ^ n[1838];
assign t[1839] = t[1838] ^ n[1839];
assign t[1840] = t[1839] ^ n[1840];
assign t[1841] = t[1840] ^ n[1841];
assign t[1842] = t[1841] ^ n[1842];
assign t[1843] = t[1842] ^ n[1843];
assign t[1844] = t[1843] ^ n[1844];
assign t[1845] = t[1844] ^ n[1845];
assign t[1846] = t[1845] ^ n[1846];
assign t[1847] = t[1846] ^ n[1847];
assign t[1848] = t[1847] ^ n[1848];
assign t[1849] = t[1848] ^ n[1849];
assign t[1850] = t[1849] ^ n[1850];
assign t[1851] = t[1850] ^ n[1851];
assign t[1852] = t[1851] ^ n[1852];
assign t[1853] = t[1852] ^ n[1853];
assign t[1854] = t[1853] ^ n[1854];
assign t[1855] = t[1854] ^ n[1855];
assign t[1856] = t[1855] ^ n[1856];
assign t[1857] = t[1856] ^ n[1857];
assign t[1858] = t[1857] ^ n[1858];
assign t[1859] = t[1858] ^ n[1859];
assign t[1860] = t[1859] ^ n[1860];
assign t[1861] = t[1860] ^ n[1861];
assign t[1862] = t[1861] ^ n[1862];
assign t[1863] = t[1862] ^ n[1863];
assign t[1864] = t[1863] ^ n[1864];
assign t[1865] = t[1864] ^ n[1865];
assign t[1866] = t[1865] ^ n[1866];
assign t[1867] = t[1866] ^ n[1867];
assign t[1868] = t[1867] ^ n[1868];
assign t[1869] = t[1868] ^ n[1869];
assign t[1870] = t[1869] ^ n[1870];
assign t[1871] = t[1870] ^ n[1871];
assign t[1872] = t[1871] ^ n[1872];
assign t[1873] = t[1872] ^ n[1873];
assign t[1874] = t[1873] ^ n[1874];
assign t[1875] = t[1874] ^ n[1875];
assign t[1876] = t[1875] ^ n[1876];
assign t[1877] = t[1876] ^ n[1877];
assign t[1878] = t[1877] ^ n[1878];
assign t[1879] = t[1878] ^ n[1879];
assign t[1880] = t[1879] ^ n[1880];
assign t[1881] = t[1880] ^ n[1881];
assign t[1882] = t[1881] ^ n[1882];
assign t[1883] = t[1882] ^ n[1883];
assign t[1884] = t[1883] ^ n[1884];
assign t[1885] = t[1884] ^ n[1885];
assign t[1886] = t[1885] ^ n[1886];
assign t[1887] = t[1886] ^ n[1887];
assign t[1888] = t[1887] ^ n[1888];
assign t[1889] = t[1888] ^ n[1889];
assign t[1890] = t[1889] ^ n[1890];
assign t[1891] = t[1890] ^ n[1891];
assign t[1892] = t[1891] ^ n[1892];
assign t[1893] = t[1892] ^ n[1893];
assign t[1894] = t[1893] ^ n[1894];
assign t[1895] = t[1894] ^ n[1895];
assign t[1896] = t[1895] ^ n[1896];
assign t[1897] = t[1896] ^ n[1897];
assign t[1898] = t[1897] ^ n[1898];
assign t[1899] = t[1898] ^ n[1899];
assign t[1900] = t[1899] ^ n[1900];
assign t[1901] = t[1900] ^ n[1901];
assign t[1902] = t[1901] ^ n[1902];
assign t[1903] = t[1902] ^ n[1903];
assign t[1904] = t[1903] ^ n[1904];
assign t[1905] = t[1904] ^ n[1905];
assign t[1906] = t[1905] ^ n[1906];
assign t[1907] = t[1906] ^ n[1907];
assign t[1908] = t[1907] ^ n[1908];
assign t[1909] = t[1908] ^ n[1909];
assign t[1910] = t[1909] ^ n[1910];
assign t[1911] = t[1910] ^ n[1911];
assign t[1912] = t[1911] ^ n[1912];
assign t[1913] = t[1912] ^ n[1913];
assign t[1914] = t[1913] ^ n[1914];
assign t[1915] = t[1914] ^ n[1915];
assign t[1916] = t[1915] ^ n[1916];
assign t[1917] = t[1916] ^ n[1917];
assign t[1918] = t[1917] ^ n[1918];
assign t[1919] = t[1918] ^ n[1919];
assign t[1920] = t[1919] ^ n[1920];
assign t[1921] = t[1920] ^ n[1921];
assign t[1922] = t[1921] ^ n[1922];
assign t[1923] = t[1922] ^ n[1923];
assign t[1924] = t[1923] ^ n[1924];
assign t[1925] = t[1924] ^ n[1925];
assign t[1926] = t[1925] ^ n[1926];
assign t[1927] = t[1926] ^ n[1927];
assign t[1928] = t[1927] ^ n[1928];
assign t[1929] = t[1928] ^ n[1929];
assign t[1930] = t[1929] ^ n[1930];
assign t[1931] = t[1930] ^ n[1931];
assign t[1932] = t[1931] ^ n[1932];
assign t[1933] = t[1932] ^ n[1933];
assign t[1934] = t[1933] ^ n[1934];
assign t[1935] = t[1934] ^ n[1935];
assign t[1936] = t[1935] ^ n[1936];
assign t[1937] = t[1936] ^ n[1937];
assign t[1938] = t[1937] ^ n[1938];
assign t[1939] = t[1938] ^ n[1939];
assign t[1940] = t[1939] ^ n[1940];
assign t[1941] = t[1940] ^ n[1941];
assign t[1942] = t[1941] ^ n[1942];
assign t[1943] = t[1942] ^ n[1943];
assign t[1944] = t[1943] ^ n[1944];
assign t[1945] = t[1944] ^ n[1945];
assign t[1946] = t[1945] ^ n[1946];
assign t[1947] = t[1946] ^ n[1947];
assign t[1948] = t[1947] ^ n[1948];
assign t[1949] = t[1948] ^ n[1949];
assign t[1950] = t[1949] ^ n[1950];
assign t[1951] = t[1950] ^ n[1951];
assign t[1952] = t[1951] ^ n[1952];
assign t[1953] = t[1952] ^ n[1953];
assign t[1954] = t[1953] ^ n[1954];
assign t[1955] = t[1954] ^ n[1955];
assign t[1956] = t[1955] ^ n[1956];
assign t[1957] = t[1956] ^ n[1957];
assign t[1958] = t[1957] ^ n[1958];
assign t[1959] = t[1958] ^ n[1959];
assign t[1960] = t[1959] ^ n[1960];
assign t[1961] = t[1960] ^ n[1961];
assign t[1962] = t[1961] ^ n[1962];
assign t[1963] = t[1962] ^ n[1963];
assign t[1964] = t[1963] ^ n[1964];
assign t[1965] = t[1964] ^ n[1965];
assign t[1966] = t[1965] ^ n[1966];
assign t[1967] = t[1966] ^ n[1967];
assign t[1968] = t[1967] ^ n[1968];
assign t[1969] = t[1968] ^ n[1969];
assign t[1970] = t[1969] ^ n[1970];
assign t[1971] = t[1970] ^ n[1971];
assign t[1972] = t[1971] ^ n[1972];
assign t[1973] = t[1972] ^ n[1973];
assign t[1974] = t[1973] ^ n[1974];
assign t[1975] = t[1974] ^ n[1975];
assign t[1976] = t[1975] ^ n[1976];
assign t[1977] = t[1976] ^ n[1977];
assign t[1978] = t[1977] ^ n[1978];
assign t[1979] = t[1978] ^ n[1979];
assign t[1980] = t[1979] ^ n[1980];
assign t[1981] = t[1980] ^ n[1981];
assign t[1982] = t[1981] ^ n[1982];
assign t[1983] = t[1982] ^ n[1983];
assign t[1984] = t[1983] ^ n[1984];
assign t[1985] = t[1984] ^ n[1985];
assign t[1986] = t[1985] ^ n[1986];
assign t[1987] = t[1986] ^ n[1987];
assign t[1988] = t[1987] ^ n[1988];
assign t[1989] = t[1988] ^ n[1989];
assign t[1990] = t[1989] ^ n[1990];
assign t[1991] = t[1990] ^ n[1991];
assign t[1992] = t[1991] ^ n[1992];
assign t[1993] = t[1992] ^ n[1993];
assign t[1994] = t[1993] ^ n[1994];
assign t[1995] = t[1994] ^ n[1995];
assign t[1996] = t[1995] ^ n[1996];
assign t[1997] = t[1996] ^ n[1997];
assign t[1998] = t[1997] ^ n[1998];
assign t[1999] = t[1998] ^ n[1999];
assign t[2000] = t[1999] ^ n[2000];
assign t[2001] = t[2000] ^ n[2001];
assign t[2002] = t[2001] ^ n[2002];
assign t[2003] = t[2002] ^ n[2003];
assign t[2004] = t[2003] ^ n[2004];
assign t[2005] = t[2004] ^ n[2005];
assign t[2006] = t[2005] ^ n[2006];
assign t[2007] = t[2006] ^ n[2007];
assign t[2008] = t[2007] ^ n[2008];
assign t[2009] = t[2008] ^ n[2009];
assign t[2010] = t[2009] ^ n[2010];
assign t[2011] = t[2010] ^ n[2011];
assign t[2012] = t[2011] ^ n[2012];
assign t[2013] = t[2012] ^ n[2013];
assign t[2014] = t[2013] ^ n[2014];
assign t[2015] = t[2014] ^ n[2015];
assign t[2016] = t[2015] ^ n[2016];
assign t[2017] = t[2016] ^ n[2017];
assign t[2018] = t[2017] ^ n[2018];
assign t[2019] = t[2018] ^ n[2019];
assign t[2020] = t[2019] ^ n[2020];
assign t[2021] = t[2020] ^ n[2021];
assign t[2022] = t[2021] ^ n[2022];
assign t[2023] = t[2022] ^ n[2023];
assign t[2024] = t[2023] ^ n[2024];
assign t[2025] = t[2024] ^ n[2025];
assign t[2026] = t[2025] ^ n[2026];
assign t[2027] = t[2026] ^ n[2027];
assign t[2028] = t[2027] ^ n[2028];
assign t[2029] = t[2028] ^ n[2029];
assign t[2030] = t[2029] ^ n[2030];
assign t[2031] = t[2030] ^ n[2031];
assign t[2032] = t[2031] ^ n[2032];
assign t[2033] = t[2032] ^ n[2033];
assign t[2034] = t[2033] ^ n[2034];
assign t[2035] = t[2034] ^ n[2035];

//asigning bit 10
assign s[10] = ( a[10] ^ b [10] ) ^ t[2035];

assign t[2036] = n[2036];
assign t[2037] = t[2036] ^ n[2037];
assign t[2038] = t[2037] ^ n[2038];
assign t[2039] = t[2038] ^ n[2039];
assign t[2040] = t[2039] ^ n[2040];
assign t[2041] = t[2040] ^ n[2041];
assign t[2042] = t[2041] ^ n[2042];
assign t[2043] = t[2042] ^ n[2043];
assign t[2044] = t[2043] ^ n[2044];
assign t[2045] = t[2044] ^ n[2045];
assign t[2046] = t[2045] ^ n[2046];
assign t[2047] = t[2046] ^ n[2047];
assign t[2048] = t[2047] ^ n[2048];
assign t[2049] = t[2048] ^ n[2049];
assign t[2050] = t[2049] ^ n[2050];
assign t[2051] = t[2050] ^ n[2051];
assign t[2052] = t[2051] ^ n[2052];
assign t[2053] = t[2052] ^ n[2053];
assign t[2054] = t[2053] ^ n[2054];
assign t[2055] = t[2054] ^ n[2055];
assign t[2056] = t[2055] ^ n[2056];
assign t[2057] = t[2056] ^ n[2057];
assign t[2058] = t[2057] ^ n[2058];
assign t[2059] = t[2058] ^ n[2059];
assign t[2060] = t[2059] ^ n[2060];
assign t[2061] = t[2060] ^ n[2061];
assign t[2062] = t[2061] ^ n[2062];
assign t[2063] = t[2062] ^ n[2063];
assign t[2064] = t[2063] ^ n[2064];
assign t[2065] = t[2064] ^ n[2065];
assign t[2066] = t[2065] ^ n[2066];
assign t[2067] = t[2066] ^ n[2067];
assign t[2068] = t[2067] ^ n[2068];
assign t[2069] = t[2068] ^ n[2069];
assign t[2070] = t[2069] ^ n[2070];
assign t[2071] = t[2070] ^ n[2071];
assign t[2072] = t[2071] ^ n[2072];
assign t[2073] = t[2072] ^ n[2073];
assign t[2074] = t[2073] ^ n[2074];
assign t[2075] = t[2074] ^ n[2075];
assign t[2076] = t[2075] ^ n[2076];
assign t[2077] = t[2076] ^ n[2077];
assign t[2078] = t[2077] ^ n[2078];
assign t[2079] = t[2078] ^ n[2079];
assign t[2080] = t[2079] ^ n[2080];
assign t[2081] = t[2080] ^ n[2081];
assign t[2082] = t[2081] ^ n[2082];
assign t[2083] = t[2082] ^ n[2083];
assign t[2084] = t[2083] ^ n[2084];
assign t[2085] = t[2084] ^ n[2085];
assign t[2086] = t[2085] ^ n[2086];
assign t[2087] = t[2086] ^ n[2087];
assign t[2088] = t[2087] ^ n[2088];
assign t[2089] = t[2088] ^ n[2089];
assign t[2090] = t[2089] ^ n[2090];
assign t[2091] = t[2090] ^ n[2091];
assign t[2092] = t[2091] ^ n[2092];
assign t[2093] = t[2092] ^ n[2093];
assign t[2094] = t[2093] ^ n[2094];
assign t[2095] = t[2094] ^ n[2095];
assign t[2096] = t[2095] ^ n[2096];
assign t[2097] = t[2096] ^ n[2097];
assign t[2098] = t[2097] ^ n[2098];
assign t[2099] = t[2098] ^ n[2099];
assign t[2100] = t[2099] ^ n[2100];
assign t[2101] = t[2100] ^ n[2101];
assign t[2102] = t[2101] ^ n[2102];
assign t[2103] = t[2102] ^ n[2103];
assign t[2104] = t[2103] ^ n[2104];
assign t[2105] = t[2104] ^ n[2105];
assign t[2106] = t[2105] ^ n[2106];
assign t[2107] = t[2106] ^ n[2107];
assign t[2108] = t[2107] ^ n[2108];
assign t[2109] = t[2108] ^ n[2109];
assign t[2110] = t[2109] ^ n[2110];
assign t[2111] = t[2110] ^ n[2111];
assign t[2112] = t[2111] ^ n[2112];
assign t[2113] = t[2112] ^ n[2113];
assign t[2114] = t[2113] ^ n[2114];
assign t[2115] = t[2114] ^ n[2115];
assign t[2116] = t[2115] ^ n[2116];
assign t[2117] = t[2116] ^ n[2117];
assign t[2118] = t[2117] ^ n[2118];
assign t[2119] = t[2118] ^ n[2119];
assign t[2120] = t[2119] ^ n[2120];
assign t[2121] = t[2120] ^ n[2121];
assign t[2122] = t[2121] ^ n[2122];
assign t[2123] = t[2122] ^ n[2123];
assign t[2124] = t[2123] ^ n[2124];
assign t[2125] = t[2124] ^ n[2125];
assign t[2126] = t[2125] ^ n[2126];
assign t[2127] = t[2126] ^ n[2127];
assign t[2128] = t[2127] ^ n[2128];
assign t[2129] = t[2128] ^ n[2129];
assign t[2130] = t[2129] ^ n[2130];
assign t[2131] = t[2130] ^ n[2131];
assign t[2132] = t[2131] ^ n[2132];
assign t[2133] = t[2132] ^ n[2133];
assign t[2134] = t[2133] ^ n[2134];
assign t[2135] = t[2134] ^ n[2135];
assign t[2136] = t[2135] ^ n[2136];
assign t[2137] = t[2136] ^ n[2137];
assign t[2138] = t[2137] ^ n[2138];
assign t[2139] = t[2138] ^ n[2139];
assign t[2140] = t[2139] ^ n[2140];
assign t[2141] = t[2140] ^ n[2141];
assign t[2142] = t[2141] ^ n[2142];
assign t[2143] = t[2142] ^ n[2143];
assign t[2144] = t[2143] ^ n[2144];
assign t[2145] = t[2144] ^ n[2145];
assign t[2146] = t[2145] ^ n[2146];
assign t[2147] = t[2146] ^ n[2147];
assign t[2148] = t[2147] ^ n[2148];
assign t[2149] = t[2148] ^ n[2149];
assign t[2150] = t[2149] ^ n[2150];
assign t[2151] = t[2150] ^ n[2151];
assign t[2152] = t[2151] ^ n[2152];
assign t[2153] = t[2152] ^ n[2153];
assign t[2154] = t[2153] ^ n[2154];
assign t[2155] = t[2154] ^ n[2155];
assign t[2156] = t[2155] ^ n[2156];
assign t[2157] = t[2156] ^ n[2157];
assign t[2158] = t[2157] ^ n[2158];
assign t[2159] = t[2158] ^ n[2159];
assign t[2160] = t[2159] ^ n[2160];
assign t[2161] = t[2160] ^ n[2161];
assign t[2162] = t[2161] ^ n[2162];
assign t[2163] = t[2162] ^ n[2163];
assign t[2164] = t[2163] ^ n[2164];
assign t[2165] = t[2164] ^ n[2165];
assign t[2166] = t[2165] ^ n[2166];
assign t[2167] = t[2166] ^ n[2167];
assign t[2168] = t[2167] ^ n[2168];
assign t[2169] = t[2168] ^ n[2169];
assign t[2170] = t[2169] ^ n[2170];
assign t[2171] = t[2170] ^ n[2171];
assign t[2172] = t[2171] ^ n[2172];
assign t[2173] = t[2172] ^ n[2173];
assign t[2174] = t[2173] ^ n[2174];
assign t[2175] = t[2174] ^ n[2175];
assign t[2176] = t[2175] ^ n[2176];
assign t[2177] = t[2176] ^ n[2177];
assign t[2178] = t[2177] ^ n[2178];
assign t[2179] = t[2178] ^ n[2179];
assign t[2180] = t[2179] ^ n[2180];
assign t[2181] = t[2180] ^ n[2181];
assign t[2182] = t[2181] ^ n[2182];
assign t[2183] = t[2182] ^ n[2183];
assign t[2184] = t[2183] ^ n[2184];
assign t[2185] = t[2184] ^ n[2185];
assign t[2186] = t[2185] ^ n[2186];
assign t[2187] = t[2186] ^ n[2187];
assign t[2188] = t[2187] ^ n[2188];
assign t[2189] = t[2188] ^ n[2189];
assign t[2190] = t[2189] ^ n[2190];
assign t[2191] = t[2190] ^ n[2191];
assign t[2192] = t[2191] ^ n[2192];
assign t[2193] = t[2192] ^ n[2193];
assign t[2194] = t[2193] ^ n[2194];
assign t[2195] = t[2194] ^ n[2195];
assign t[2196] = t[2195] ^ n[2196];
assign t[2197] = t[2196] ^ n[2197];
assign t[2198] = t[2197] ^ n[2198];
assign t[2199] = t[2198] ^ n[2199];
assign t[2200] = t[2199] ^ n[2200];
assign t[2201] = t[2200] ^ n[2201];
assign t[2202] = t[2201] ^ n[2202];
assign t[2203] = t[2202] ^ n[2203];
assign t[2204] = t[2203] ^ n[2204];
assign t[2205] = t[2204] ^ n[2205];
assign t[2206] = t[2205] ^ n[2206];
assign t[2207] = t[2206] ^ n[2207];
assign t[2208] = t[2207] ^ n[2208];
assign t[2209] = t[2208] ^ n[2209];
assign t[2210] = t[2209] ^ n[2210];
assign t[2211] = t[2210] ^ n[2211];
assign t[2212] = t[2211] ^ n[2212];
assign t[2213] = t[2212] ^ n[2213];
assign t[2214] = t[2213] ^ n[2214];
assign t[2215] = t[2214] ^ n[2215];
assign t[2216] = t[2215] ^ n[2216];
assign t[2217] = t[2216] ^ n[2217];
assign t[2218] = t[2217] ^ n[2218];
assign t[2219] = t[2218] ^ n[2219];
assign t[2220] = t[2219] ^ n[2220];
assign t[2221] = t[2220] ^ n[2221];
assign t[2222] = t[2221] ^ n[2222];
assign t[2223] = t[2222] ^ n[2223];
assign t[2224] = t[2223] ^ n[2224];
assign t[2225] = t[2224] ^ n[2225];
assign t[2226] = t[2225] ^ n[2226];
assign t[2227] = t[2226] ^ n[2227];
assign t[2228] = t[2227] ^ n[2228];
assign t[2229] = t[2228] ^ n[2229];
assign t[2230] = t[2229] ^ n[2230];
assign t[2231] = t[2230] ^ n[2231];
assign t[2232] = t[2231] ^ n[2232];
assign t[2233] = t[2232] ^ n[2233];
assign t[2234] = t[2233] ^ n[2234];
assign t[2235] = t[2234] ^ n[2235];
assign t[2236] = t[2235] ^ n[2236];
assign t[2237] = t[2236] ^ n[2237];
assign t[2238] = t[2237] ^ n[2238];
assign t[2239] = t[2238] ^ n[2239];
assign t[2240] = t[2239] ^ n[2240];
assign t[2241] = t[2240] ^ n[2241];
assign t[2242] = t[2241] ^ n[2242];
assign t[2243] = t[2242] ^ n[2243];
assign t[2244] = t[2243] ^ n[2244];
assign t[2245] = t[2244] ^ n[2245];
assign t[2246] = t[2245] ^ n[2246];
assign t[2247] = t[2246] ^ n[2247];
assign t[2248] = t[2247] ^ n[2248];
assign t[2249] = t[2248] ^ n[2249];
assign t[2250] = t[2249] ^ n[2250];
assign t[2251] = t[2250] ^ n[2251];
assign t[2252] = t[2251] ^ n[2252];
assign t[2253] = t[2252] ^ n[2253];
assign t[2254] = t[2253] ^ n[2254];
assign t[2255] = t[2254] ^ n[2255];
assign t[2256] = t[2255] ^ n[2256];
assign t[2257] = t[2256] ^ n[2257];
assign t[2258] = t[2257] ^ n[2258];
assign t[2259] = t[2258] ^ n[2259];
assign t[2260] = t[2259] ^ n[2260];
assign t[2261] = t[2260] ^ n[2261];
assign t[2262] = t[2261] ^ n[2262];
assign t[2263] = t[2262] ^ n[2263];
assign t[2264] = t[2263] ^ n[2264];
assign t[2265] = t[2264] ^ n[2265];
assign t[2266] = t[2265] ^ n[2266];
assign t[2267] = t[2266] ^ n[2267];
assign t[2268] = t[2267] ^ n[2268];
assign t[2269] = t[2268] ^ n[2269];
assign t[2270] = t[2269] ^ n[2270];
assign t[2271] = t[2270] ^ n[2271];
assign t[2272] = t[2271] ^ n[2272];
assign t[2273] = t[2272] ^ n[2273];
assign t[2274] = t[2273] ^ n[2274];
assign t[2275] = t[2274] ^ n[2275];
assign t[2276] = t[2275] ^ n[2276];
assign t[2277] = t[2276] ^ n[2277];
assign t[2278] = t[2277] ^ n[2278];
assign t[2279] = t[2278] ^ n[2279];
assign t[2280] = t[2279] ^ n[2280];
assign t[2281] = t[2280] ^ n[2281];
assign t[2282] = t[2281] ^ n[2282];
assign t[2283] = t[2282] ^ n[2283];
assign t[2284] = t[2283] ^ n[2284];
assign t[2285] = t[2284] ^ n[2285];
assign t[2286] = t[2285] ^ n[2286];
assign t[2287] = t[2286] ^ n[2287];
assign t[2288] = t[2287] ^ n[2288];
assign t[2289] = t[2288] ^ n[2289];
assign t[2290] = t[2289] ^ n[2290];
assign t[2291] = t[2290] ^ n[2291];
assign t[2292] = t[2291] ^ n[2292];
assign t[2293] = t[2292] ^ n[2293];
assign t[2294] = t[2293] ^ n[2294];
assign t[2295] = t[2294] ^ n[2295];
assign t[2296] = t[2295] ^ n[2296];
assign t[2297] = t[2296] ^ n[2297];
assign t[2298] = t[2297] ^ n[2298];
assign t[2299] = t[2298] ^ n[2299];
assign t[2300] = t[2299] ^ n[2300];
assign t[2301] = t[2300] ^ n[2301];
assign t[2302] = t[2301] ^ n[2302];
assign t[2303] = t[2302] ^ n[2303];
assign t[2304] = t[2303] ^ n[2304];
assign t[2305] = t[2304] ^ n[2305];
assign t[2306] = t[2305] ^ n[2306];
assign t[2307] = t[2306] ^ n[2307];
assign t[2308] = t[2307] ^ n[2308];
assign t[2309] = t[2308] ^ n[2309];
assign t[2310] = t[2309] ^ n[2310];
assign t[2311] = t[2310] ^ n[2311];
assign t[2312] = t[2311] ^ n[2312];
assign t[2313] = t[2312] ^ n[2313];
assign t[2314] = t[2313] ^ n[2314];
assign t[2315] = t[2314] ^ n[2315];
assign t[2316] = t[2315] ^ n[2316];
assign t[2317] = t[2316] ^ n[2317];
assign t[2318] = t[2317] ^ n[2318];
assign t[2319] = t[2318] ^ n[2319];
assign t[2320] = t[2319] ^ n[2320];
assign t[2321] = t[2320] ^ n[2321];
assign t[2322] = t[2321] ^ n[2322];
assign t[2323] = t[2322] ^ n[2323];
assign t[2324] = t[2323] ^ n[2324];
assign t[2325] = t[2324] ^ n[2325];
assign t[2326] = t[2325] ^ n[2326];
assign t[2327] = t[2326] ^ n[2327];
assign t[2328] = t[2327] ^ n[2328];
assign t[2329] = t[2328] ^ n[2329];
assign t[2330] = t[2329] ^ n[2330];
assign t[2331] = t[2330] ^ n[2331];
assign t[2332] = t[2331] ^ n[2332];
assign t[2333] = t[2332] ^ n[2333];
assign t[2334] = t[2333] ^ n[2334];
assign t[2335] = t[2334] ^ n[2335];
assign t[2336] = t[2335] ^ n[2336];
assign t[2337] = t[2336] ^ n[2337];
assign t[2338] = t[2337] ^ n[2338];
assign t[2339] = t[2338] ^ n[2339];
assign t[2340] = t[2339] ^ n[2340];
assign t[2341] = t[2340] ^ n[2341];
assign t[2342] = t[2341] ^ n[2342];
assign t[2343] = t[2342] ^ n[2343];
assign t[2344] = t[2343] ^ n[2344];
assign t[2345] = t[2344] ^ n[2345];
assign t[2346] = t[2345] ^ n[2346];
assign t[2347] = t[2346] ^ n[2347];
assign t[2348] = t[2347] ^ n[2348];
assign t[2349] = t[2348] ^ n[2349];
assign t[2350] = t[2349] ^ n[2350];
assign t[2351] = t[2350] ^ n[2351];
assign t[2352] = t[2351] ^ n[2352];
assign t[2353] = t[2352] ^ n[2353];
assign t[2354] = t[2353] ^ n[2354];
assign t[2355] = t[2354] ^ n[2355];
assign t[2356] = t[2355] ^ n[2356];
assign t[2357] = t[2356] ^ n[2357];
assign t[2358] = t[2357] ^ n[2358];
assign t[2359] = t[2358] ^ n[2359];
assign t[2360] = t[2359] ^ n[2360];
assign t[2361] = t[2360] ^ n[2361];
assign t[2362] = t[2361] ^ n[2362];
assign t[2363] = t[2362] ^ n[2363];
assign t[2364] = t[2363] ^ n[2364];
assign t[2365] = t[2364] ^ n[2365];
assign t[2366] = t[2365] ^ n[2366];
assign t[2367] = t[2366] ^ n[2367];
assign t[2368] = t[2367] ^ n[2368];
assign t[2369] = t[2368] ^ n[2369];
assign t[2370] = t[2369] ^ n[2370];
assign t[2371] = t[2370] ^ n[2371];
assign t[2372] = t[2371] ^ n[2372];
assign t[2373] = t[2372] ^ n[2373];
assign t[2374] = t[2373] ^ n[2374];
assign t[2375] = t[2374] ^ n[2375];
assign t[2376] = t[2375] ^ n[2376];
assign t[2377] = t[2376] ^ n[2377];
assign t[2378] = t[2377] ^ n[2378];
assign t[2379] = t[2378] ^ n[2379];
assign t[2380] = t[2379] ^ n[2380];
assign t[2381] = t[2380] ^ n[2381];
assign t[2382] = t[2381] ^ n[2382];
assign t[2383] = t[2382] ^ n[2383];
assign t[2384] = t[2383] ^ n[2384];
assign t[2385] = t[2384] ^ n[2385];
assign t[2386] = t[2385] ^ n[2386];
assign t[2387] = t[2386] ^ n[2387];
assign t[2388] = t[2387] ^ n[2388];
assign t[2389] = t[2388] ^ n[2389];
assign t[2390] = t[2389] ^ n[2390];
assign t[2391] = t[2390] ^ n[2391];
assign t[2392] = t[2391] ^ n[2392];
assign t[2393] = t[2392] ^ n[2393];
assign t[2394] = t[2393] ^ n[2394];
assign t[2395] = t[2394] ^ n[2395];
assign t[2396] = t[2395] ^ n[2396];
assign t[2397] = t[2396] ^ n[2397];
assign t[2398] = t[2397] ^ n[2398];
assign t[2399] = t[2398] ^ n[2399];
assign t[2400] = t[2399] ^ n[2400];
assign t[2401] = t[2400] ^ n[2401];
assign t[2402] = t[2401] ^ n[2402];
assign t[2403] = t[2402] ^ n[2403];
assign t[2404] = t[2403] ^ n[2404];
assign t[2405] = t[2404] ^ n[2405];
assign t[2406] = t[2405] ^ n[2406];
assign t[2407] = t[2406] ^ n[2407];
assign t[2408] = t[2407] ^ n[2408];
assign t[2409] = t[2408] ^ n[2409];
assign t[2410] = t[2409] ^ n[2410];
assign t[2411] = t[2410] ^ n[2411];
assign t[2412] = t[2411] ^ n[2412];
assign t[2413] = t[2412] ^ n[2413];
assign t[2414] = t[2413] ^ n[2414];
assign t[2415] = t[2414] ^ n[2415];
assign t[2416] = t[2415] ^ n[2416];
assign t[2417] = t[2416] ^ n[2417];
assign t[2418] = t[2417] ^ n[2418];
assign t[2419] = t[2418] ^ n[2419];
assign t[2420] = t[2419] ^ n[2420];
assign t[2421] = t[2420] ^ n[2421];
assign t[2422] = t[2421] ^ n[2422];
assign t[2423] = t[2422] ^ n[2423];
assign t[2424] = t[2423] ^ n[2424];
assign t[2425] = t[2424] ^ n[2425];
assign t[2426] = t[2425] ^ n[2426];
assign t[2427] = t[2426] ^ n[2427];
assign t[2428] = t[2427] ^ n[2428];
assign t[2429] = t[2428] ^ n[2429];
assign t[2430] = t[2429] ^ n[2430];
assign t[2431] = t[2430] ^ n[2431];
assign t[2432] = t[2431] ^ n[2432];
assign t[2433] = t[2432] ^ n[2433];
assign t[2434] = t[2433] ^ n[2434];
assign t[2435] = t[2434] ^ n[2435];
assign t[2436] = t[2435] ^ n[2436];
assign t[2437] = t[2436] ^ n[2437];
assign t[2438] = t[2437] ^ n[2438];
assign t[2439] = t[2438] ^ n[2439];
assign t[2440] = t[2439] ^ n[2440];
assign t[2441] = t[2440] ^ n[2441];
assign t[2442] = t[2441] ^ n[2442];
assign t[2443] = t[2442] ^ n[2443];
assign t[2444] = t[2443] ^ n[2444];
assign t[2445] = t[2444] ^ n[2445];
assign t[2446] = t[2445] ^ n[2446];
assign t[2447] = t[2446] ^ n[2447];
assign t[2448] = t[2447] ^ n[2448];
assign t[2449] = t[2448] ^ n[2449];
assign t[2450] = t[2449] ^ n[2450];
assign t[2451] = t[2450] ^ n[2451];
assign t[2452] = t[2451] ^ n[2452];
assign t[2453] = t[2452] ^ n[2453];
assign t[2454] = t[2453] ^ n[2454];
assign t[2455] = t[2454] ^ n[2455];
assign t[2456] = t[2455] ^ n[2456];
assign t[2457] = t[2456] ^ n[2457];
assign t[2458] = t[2457] ^ n[2458];
assign t[2459] = t[2458] ^ n[2459];
assign t[2460] = t[2459] ^ n[2460];
assign t[2461] = t[2460] ^ n[2461];
assign t[2462] = t[2461] ^ n[2462];
assign t[2463] = t[2462] ^ n[2463];
assign t[2464] = t[2463] ^ n[2464];
assign t[2465] = t[2464] ^ n[2465];
assign t[2466] = t[2465] ^ n[2466];
assign t[2467] = t[2466] ^ n[2467];
assign t[2468] = t[2467] ^ n[2468];
assign t[2469] = t[2468] ^ n[2469];
assign t[2470] = t[2469] ^ n[2470];
assign t[2471] = t[2470] ^ n[2471];
assign t[2472] = t[2471] ^ n[2472];
assign t[2473] = t[2472] ^ n[2473];
assign t[2474] = t[2473] ^ n[2474];
assign t[2475] = t[2474] ^ n[2475];
assign t[2476] = t[2475] ^ n[2476];
assign t[2477] = t[2476] ^ n[2477];
assign t[2478] = t[2477] ^ n[2478];
assign t[2479] = t[2478] ^ n[2479];
assign t[2480] = t[2479] ^ n[2480];
assign t[2481] = t[2480] ^ n[2481];
assign t[2482] = t[2481] ^ n[2482];
assign t[2483] = t[2482] ^ n[2483];
assign t[2484] = t[2483] ^ n[2484];
assign t[2485] = t[2484] ^ n[2485];
assign t[2486] = t[2485] ^ n[2486];
assign t[2487] = t[2486] ^ n[2487];
assign t[2488] = t[2487] ^ n[2488];
assign t[2489] = t[2488] ^ n[2489];
assign t[2490] = t[2489] ^ n[2490];
assign t[2491] = t[2490] ^ n[2491];
assign t[2492] = t[2491] ^ n[2492];
assign t[2493] = t[2492] ^ n[2493];
assign t[2494] = t[2493] ^ n[2494];
assign t[2495] = t[2494] ^ n[2495];
assign t[2496] = t[2495] ^ n[2496];
assign t[2497] = t[2496] ^ n[2497];
assign t[2498] = t[2497] ^ n[2498];
assign t[2499] = t[2498] ^ n[2499];
assign t[2500] = t[2499] ^ n[2500];
assign t[2501] = t[2500] ^ n[2501];
assign t[2502] = t[2501] ^ n[2502];
assign t[2503] = t[2502] ^ n[2503];
assign t[2504] = t[2503] ^ n[2504];
assign t[2505] = t[2504] ^ n[2505];
assign t[2506] = t[2505] ^ n[2506];
assign t[2507] = t[2506] ^ n[2507];
assign t[2508] = t[2507] ^ n[2508];
assign t[2509] = t[2508] ^ n[2509];
assign t[2510] = t[2509] ^ n[2510];
assign t[2511] = t[2510] ^ n[2511];
assign t[2512] = t[2511] ^ n[2512];
assign t[2513] = t[2512] ^ n[2513];
assign t[2514] = t[2513] ^ n[2514];
assign t[2515] = t[2514] ^ n[2515];
assign t[2516] = t[2515] ^ n[2516];
assign t[2517] = t[2516] ^ n[2517];
assign t[2518] = t[2517] ^ n[2518];
assign t[2519] = t[2518] ^ n[2519];
assign t[2520] = t[2519] ^ n[2520];
assign t[2521] = t[2520] ^ n[2521];
assign t[2522] = t[2521] ^ n[2522];
assign t[2523] = t[2522] ^ n[2523];
assign t[2524] = t[2523] ^ n[2524];
assign t[2525] = t[2524] ^ n[2525];
assign t[2526] = t[2525] ^ n[2526];
assign t[2527] = t[2526] ^ n[2527];
assign t[2528] = t[2527] ^ n[2528];
assign t[2529] = t[2528] ^ n[2529];
assign t[2530] = t[2529] ^ n[2530];
assign t[2531] = t[2530] ^ n[2531];
assign t[2532] = t[2531] ^ n[2532];
assign t[2533] = t[2532] ^ n[2533];
assign t[2534] = t[2533] ^ n[2534];
assign t[2535] = t[2534] ^ n[2535];
assign t[2536] = t[2535] ^ n[2536];
assign t[2537] = t[2536] ^ n[2537];
assign t[2538] = t[2537] ^ n[2538];
assign t[2539] = t[2538] ^ n[2539];
assign t[2540] = t[2539] ^ n[2540];
assign t[2541] = t[2540] ^ n[2541];
assign t[2542] = t[2541] ^ n[2542];
assign t[2543] = t[2542] ^ n[2543];
assign t[2544] = t[2543] ^ n[2544];
assign t[2545] = t[2544] ^ n[2545];
assign t[2546] = t[2545] ^ n[2546];
assign t[2547] = t[2546] ^ n[2547];
assign t[2548] = t[2547] ^ n[2548];
assign t[2549] = t[2548] ^ n[2549];
assign t[2550] = t[2549] ^ n[2550];
assign t[2551] = t[2550] ^ n[2551];
assign t[2552] = t[2551] ^ n[2552];
assign t[2553] = t[2552] ^ n[2553];
assign t[2554] = t[2553] ^ n[2554];
assign t[2555] = t[2554] ^ n[2555];
assign t[2556] = t[2555] ^ n[2556];
assign t[2557] = t[2556] ^ n[2557];
assign t[2558] = t[2557] ^ n[2558];
assign t[2559] = t[2558] ^ n[2559];
assign t[2560] = t[2559] ^ n[2560];
assign t[2561] = t[2560] ^ n[2561];
assign t[2562] = t[2561] ^ n[2562];
assign t[2563] = t[2562] ^ n[2563];
assign t[2564] = t[2563] ^ n[2564];
assign t[2565] = t[2564] ^ n[2565];
assign t[2566] = t[2565] ^ n[2566];
assign t[2567] = t[2566] ^ n[2567];
assign t[2568] = t[2567] ^ n[2568];
assign t[2569] = t[2568] ^ n[2569];
assign t[2570] = t[2569] ^ n[2570];
assign t[2571] = t[2570] ^ n[2571];
assign t[2572] = t[2571] ^ n[2572];
assign t[2573] = t[2572] ^ n[2573];
assign t[2574] = t[2573] ^ n[2574];
assign t[2575] = t[2574] ^ n[2575];
assign t[2576] = t[2575] ^ n[2576];
assign t[2577] = t[2576] ^ n[2577];
assign t[2578] = t[2577] ^ n[2578];
assign t[2579] = t[2578] ^ n[2579];
assign t[2580] = t[2579] ^ n[2580];
assign t[2581] = t[2580] ^ n[2581];
assign t[2582] = t[2581] ^ n[2582];
assign t[2583] = t[2582] ^ n[2583];
assign t[2584] = t[2583] ^ n[2584];
assign t[2585] = t[2584] ^ n[2585];
assign t[2586] = t[2585] ^ n[2586];
assign t[2587] = t[2586] ^ n[2587];
assign t[2588] = t[2587] ^ n[2588];
assign t[2589] = t[2588] ^ n[2589];
assign t[2590] = t[2589] ^ n[2590];
assign t[2591] = t[2590] ^ n[2591];
assign t[2592] = t[2591] ^ n[2592];
assign t[2593] = t[2592] ^ n[2593];
assign t[2594] = t[2593] ^ n[2594];
assign t[2595] = t[2594] ^ n[2595];
assign t[2596] = t[2595] ^ n[2596];
assign t[2597] = t[2596] ^ n[2597];
assign t[2598] = t[2597] ^ n[2598];
assign t[2599] = t[2598] ^ n[2599];
assign t[2600] = t[2599] ^ n[2600];
assign t[2601] = t[2600] ^ n[2601];
assign t[2602] = t[2601] ^ n[2602];
assign t[2603] = t[2602] ^ n[2603];
assign t[2604] = t[2603] ^ n[2604];
assign t[2605] = t[2604] ^ n[2605];
assign t[2606] = t[2605] ^ n[2606];
assign t[2607] = t[2606] ^ n[2607];
assign t[2608] = t[2607] ^ n[2608];
assign t[2609] = t[2608] ^ n[2609];
assign t[2610] = t[2609] ^ n[2610];
assign t[2611] = t[2610] ^ n[2611];
assign t[2612] = t[2611] ^ n[2612];
assign t[2613] = t[2612] ^ n[2613];
assign t[2614] = t[2613] ^ n[2614];
assign t[2615] = t[2614] ^ n[2615];
assign t[2616] = t[2615] ^ n[2616];
assign t[2617] = t[2616] ^ n[2617];
assign t[2618] = t[2617] ^ n[2618];
assign t[2619] = t[2618] ^ n[2619];
assign t[2620] = t[2619] ^ n[2620];
assign t[2621] = t[2620] ^ n[2621];
assign t[2622] = t[2621] ^ n[2622];
assign t[2623] = t[2622] ^ n[2623];
assign t[2624] = t[2623] ^ n[2624];
assign t[2625] = t[2624] ^ n[2625];
assign t[2626] = t[2625] ^ n[2626];
assign t[2627] = t[2626] ^ n[2627];
assign t[2628] = t[2627] ^ n[2628];
assign t[2629] = t[2628] ^ n[2629];
assign t[2630] = t[2629] ^ n[2630];
assign t[2631] = t[2630] ^ n[2631];
assign t[2632] = t[2631] ^ n[2632];
assign t[2633] = t[2632] ^ n[2633];
assign t[2634] = t[2633] ^ n[2634];
assign t[2635] = t[2634] ^ n[2635];
assign t[2636] = t[2635] ^ n[2636];
assign t[2637] = t[2636] ^ n[2637];
assign t[2638] = t[2637] ^ n[2638];
assign t[2639] = t[2638] ^ n[2639];
assign t[2640] = t[2639] ^ n[2640];
assign t[2641] = t[2640] ^ n[2641];
assign t[2642] = t[2641] ^ n[2642];
assign t[2643] = t[2642] ^ n[2643];
assign t[2644] = t[2643] ^ n[2644];
assign t[2645] = t[2644] ^ n[2645];
assign t[2646] = t[2645] ^ n[2646];
assign t[2647] = t[2646] ^ n[2647];
assign t[2648] = t[2647] ^ n[2648];
assign t[2649] = t[2648] ^ n[2649];
assign t[2650] = t[2649] ^ n[2650];
assign t[2651] = t[2650] ^ n[2651];
assign t[2652] = t[2651] ^ n[2652];
assign t[2653] = t[2652] ^ n[2653];
assign t[2654] = t[2653] ^ n[2654];
assign t[2655] = t[2654] ^ n[2655];
assign t[2656] = t[2655] ^ n[2656];
assign t[2657] = t[2656] ^ n[2657];
assign t[2658] = t[2657] ^ n[2658];
assign t[2659] = t[2658] ^ n[2659];
assign t[2660] = t[2659] ^ n[2660];
assign t[2661] = t[2660] ^ n[2661];
assign t[2662] = t[2661] ^ n[2662];
assign t[2663] = t[2662] ^ n[2663];
assign t[2664] = t[2663] ^ n[2664];
assign t[2665] = t[2664] ^ n[2665];
assign t[2666] = t[2665] ^ n[2666];
assign t[2667] = t[2666] ^ n[2667];
assign t[2668] = t[2667] ^ n[2668];
assign t[2669] = t[2668] ^ n[2669];
assign t[2670] = t[2669] ^ n[2670];
assign t[2671] = t[2670] ^ n[2671];
assign t[2672] = t[2671] ^ n[2672];
assign t[2673] = t[2672] ^ n[2673];
assign t[2674] = t[2673] ^ n[2674];
assign t[2675] = t[2674] ^ n[2675];
assign t[2676] = t[2675] ^ n[2676];
assign t[2677] = t[2676] ^ n[2677];
assign t[2678] = t[2677] ^ n[2678];
assign t[2679] = t[2678] ^ n[2679];
assign t[2680] = t[2679] ^ n[2680];
assign t[2681] = t[2680] ^ n[2681];
assign t[2682] = t[2681] ^ n[2682];
assign t[2683] = t[2682] ^ n[2683];
assign t[2684] = t[2683] ^ n[2684];
assign t[2685] = t[2684] ^ n[2685];
assign t[2686] = t[2685] ^ n[2686];
assign t[2687] = t[2686] ^ n[2687];
assign t[2688] = t[2687] ^ n[2688];
assign t[2689] = t[2688] ^ n[2689];
assign t[2690] = t[2689] ^ n[2690];
assign t[2691] = t[2690] ^ n[2691];
assign t[2692] = t[2691] ^ n[2692];
assign t[2693] = t[2692] ^ n[2693];
assign t[2694] = t[2693] ^ n[2694];
assign t[2695] = t[2694] ^ n[2695];
assign t[2696] = t[2695] ^ n[2696];
assign t[2697] = t[2696] ^ n[2697];
assign t[2698] = t[2697] ^ n[2698];
assign t[2699] = t[2698] ^ n[2699];
assign t[2700] = t[2699] ^ n[2700];
assign t[2701] = t[2700] ^ n[2701];
assign t[2702] = t[2701] ^ n[2702];
assign t[2703] = t[2702] ^ n[2703];
assign t[2704] = t[2703] ^ n[2704];
assign t[2705] = t[2704] ^ n[2705];
assign t[2706] = t[2705] ^ n[2706];
assign t[2707] = t[2706] ^ n[2707];
assign t[2708] = t[2707] ^ n[2708];
assign t[2709] = t[2708] ^ n[2709];
assign t[2710] = t[2709] ^ n[2710];
assign t[2711] = t[2710] ^ n[2711];
assign t[2712] = t[2711] ^ n[2712];
assign t[2713] = t[2712] ^ n[2713];
assign t[2714] = t[2713] ^ n[2714];
assign t[2715] = t[2714] ^ n[2715];
assign t[2716] = t[2715] ^ n[2716];
assign t[2717] = t[2716] ^ n[2717];
assign t[2718] = t[2717] ^ n[2718];
assign t[2719] = t[2718] ^ n[2719];
assign t[2720] = t[2719] ^ n[2720];
assign t[2721] = t[2720] ^ n[2721];
assign t[2722] = t[2721] ^ n[2722];
assign t[2723] = t[2722] ^ n[2723];
assign t[2724] = t[2723] ^ n[2724];
assign t[2725] = t[2724] ^ n[2725];
assign t[2726] = t[2725] ^ n[2726];
assign t[2727] = t[2726] ^ n[2727];
assign t[2728] = t[2727] ^ n[2728];
assign t[2729] = t[2728] ^ n[2729];
assign t[2730] = t[2729] ^ n[2730];
assign t[2731] = t[2730] ^ n[2731];
assign t[2732] = t[2731] ^ n[2732];
assign t[2733] = t[2732] ^ n[2733];
assign t[2734] = t[2733] ^ n[2734];
assign t[2735] = t[2734] ^ n[2735];
assign t[2736] = t[2735] ^ n[2736];
assign t[2737] = t[2736] ^ n[2737];
assign t[2738] = t[2737] ^ n[2738];
assign t[2739] = t[2738] ^ n[2739];
assign t[2740] = t[2739] ^ n[2740];
assign t[2741] = t[2740] ^ n[2741];
assign t[2742] = t[2741] ^ n[2742];
assign t[2743] = t[2742] ^ n[2743];
assign t[2744] = t[2743] ^ n[2744];
assign t[2745] = t[2744] ^ n[2745];
assign t[2746] = t[2745] ^ n[2746];
assign t[2747] = t[2746] ^ n[2747];
assign t[2748] = t[2747] ^ n[2748];
assign t[2749] = t[2748] ^ n[2749];
assign t[2750] = t[2749] ^ n[2750];
assign t[2751] = t[2750] ^ n[2751];
assign t[2752] = t[2751] ^ n[2752];
assign t[2753] = t[2752] ^ n[2753];
assign t[2754] = t[2753] ^ n[2754];
assign t[2755] = t[2754] ^ n[2755];
assign t[2756] = t[2755] ^ n[2756];
assign t[2757] = t[2756] ^ n[2757];
assign t[2758] = t[2757] ^ n[2758];
assign t[2759] = t[2758] ^ n[2759];
assign t[2760] = t[2759] ^ n[2760];
assign t[2761] = t[2760] ^ n[2761];
assign t[2762] = t[2761] ^ n[2762];
assign t[2763] = t[2762] ^ n[2763];
assign t[2764] = t[2763] ^ n[2764];
assign t[2765] = t[2764] ^ n[2765];
assign t[2766] = t[2765] ^ n[2766];
assign t[2767] = t[2766] ^ n[2767];
assign t[2768] = t[2767] ^ n[2768];
assign t[2769] = t[2768] ^ n[2769];
assign t[2770] = t[2769] ^ n[2770];
assign t[2771] = t[2770] ^ n[2771];
assign t[2772] = t[2771] ^ n[2772];
assign t[2773] = t[2772] ^ n[2773];
assign t[2774] = t[2773] ^ n[2774];
assign t[2775] = t[2774] ^ n[2775];
assign t[2776] = t[2775] ^ n[2776];
assign t[2777] = t[2776] ^ n[2777];
assign t[2778] = t[2777] ^ n[2778];
assign t[2779] = t[2778] ^ n[2779];
assign t[2780] = t[2779] ^ n[2780];
assign t[2781] = t[2780] ^ n[2781];
assign t[2782] = t[2781] ^ n[2782];
assign t[2783] = t[2782] ^ n[2783];
assign t[2784] = t[2783] ^ n[2784];
assign t[2785] = t[2784] ^ n[2785];
assign t[2786] = t[2785] ^ n[2786];
assign t[2787] = t[2786] ^ n[2787];
assign t[2788] = t[2787] ^ n[2788];
assign t[2789] = t[2788] ^ n[2789];
assign t[2790] = t[2789] ^ n[2790];
assign t[2791] = t[2790] ^ n[2791];
assign t[2792] = t[2791] ^ n[2792];
assign t[2793] = t[2792] ^ n[2793];
assign t[2794] = t[2793] ^ n[2794];
assign t[2795] = t[2794] ^ n[2795];
assign t[2796] = t[2795] ^ n[2796];
assign t[2797] = t[2796] ^ n[2797];
assign t[2798] = t[2797] ^ n[2798];
assign t[2799] = t[2798] ^ n[2799];
assign t[2800] = t[2799] ^ n[2800];
assign t[2801] = t[2800] ^ n[2801];
assign t[2802] = t[2801] ^ n[2802];
assign t[2803] = t[2802] ^ n[2803];
assign t[2804] = t[2803] ^ n[2804];
assign t[2805] = t[2804] ^ n[2805];
assign t[2806] = t[2805] ^ n[2806];
assign t[2807] = t[2806] ^ n[2807];
assign t[2808] = t[2807] ^ n[2808];
assign t[2809] = t[2808] ^ n[2809];
assign t[2810] = t[2809] ^ n[2810];
assign t[2811] = t[2810] ^ n[2811];
assign t[2812] = t[2811] ^ n[2812];
assign t[2813] = t[2812] ^ n[2813];
assign t[2814] = t[2813] ^ n[2814];
assign t[2815] = t[2814] ^ n[2815];
assign t[2816] = t[2815] ^ n[2816];
assign t[2817] = t[2816] ^ n[2817];
assign t[2818] = t[2817] ^ n[2818];
assign t[2819] = t[2818] ^ n[2819];
assign t[2820] = t[2819] ^ n[2820];
assign t[2821] = t[2820] ^ n[2821];
assign t[2822] = t[2821] ^ n[2822];
assign t[2823] = t[2822] ^ n[2823];
assign t[2824] = t[2823] ^ n[2824];
assign t[2825] = t[2824] ^ n[2825];
assign t[2826] = t[2825] ^ n[2826];
assign t[2827] = t[2826] ^ n[2827];
assign t[2828] = t[2827] ^ n[2828];
assign t[2829] = t[2828] ^ n[2829];
assign t[2830] = t[2829] ^ n[2830];
assign t[2831] = t[2830] ^ n[2831];
assign t[2832] = t[2831] ^ n[2832];
assign t[2833] = t[2832] ^ n[2833];
assign t[2834] = t[2833] ^ n[2834];
assign t[2835] = t[2834] ^ n[2835];
assign t[2836] = t[2835] ^ n[2836];
assign t[2837] = t[2836] ^ n[2837];
assign t[2838] = t[2837] ^ n[2838];
assign t[2839] = t[2838] ^ n[2839];
assign t[2840] = t[2839] ^ n[2840];
assign t[2841] = t[2840] ^ n[2841];
assign t[2842] = t[2841] ^ n[2842];
assign t[2843] = t[2842] ^ n[2843];
assign t[2844] = t[2843] ^ n[2844];
assign t[2845] = t[2844] ^ n[2845];
assign t[2846] = t[2845] ^ n[2846];
assign t[2847] = t[2846] ^ n[2847];
assign t[2848] = t[2847] ^ n[2848];
assign t[2849] = t[2848] ^ n[2849];
assign t[2850] = t[2849] ^ n[2850];
assign t[2851] = t[2850] ^ n[2851];
assign t[2852] = t[2851] ^ n[2852];
assign t[2853] = t[2852] ^ n[2853];
assign t[2854] = t[2853] ^ n[2854];
assign t[2855] = t[2854] ^ n[2855];
assign t[2856] = t[2855] ^ n[2856];
assign t[2857] = t[2856] ^ n[2857];
assign t[2858] = t[2857] ^ n[2858];
assign t[2859] = t[2858] ^ n[2859];
assign t[2860] = t[2859] ^ n[2860];
assign t[2861] = t[2860] ^ n[2861];
assign t[2862] = t[2861] ^ n[2862];
assign t[2863] = t[2862] ^ n[2863];
assign t[2864] = t[2863] ^ n[2864];
assign t[2865] = t[2864] ^ n[2865];
assign t[2866] = t[2865] ^ n[2866];
assign t[2867] = t[2866] ^ n[2867];
assign t[2868] = t[2867] ^ n[2868];
assign t[2869] = t[2868] ^ n[2869];
assign t[2870] = t[2869] ^ n[2870];
assign t[2871] = t[2870] ^ n[2871];
assign t[2872] = t[2871] ^ n[2872];
assign t[2873] = t[2872] ^ n[2873];
assign t[2874] = t[2873] ^ n[2874];
assign t[2875] = t[2874] ^ n[2875];
assign t[2876] = t[2875] ^ n[2876];
assign t[2877] = t[2876] ^ n[2877];
assign t[2878] = t[2877] ^ n[2878];
assign t[2879] = t[2878] ^ n[2879];
assign t[2880] = t[2879] ^ n[2880];
assign t[2881] = t[2880] ^ n[2881];
assign t[2882] = t[2881] ^ n[2882];
assign t[2883] = t[2882] ^ n[2883];
assign t[2884] = t[2883] ^ n[2884];
assign t[2885] = t[2884] ^ n[2885];
assign t[2886] = t[2885] ^ n[2886];
assign t[2887] = t[2886] ^ n[2887];
assign t[2888] = t[2887] ^ n[2888];
assign t[2889] = t[2888] ^ n[2889];
assign t[2890] = t[2889] ^ n[2890];
assign t[2891] = t[2890] ^ n[2891];
assign t[2892] = t[2891] ^ n[2892];
assign t[2893] = t[2892] ^ n[2893];
assign t[2894] = t[2893] ^ n[2894];
assign t[2895] = t[2894] ^ n[2895];
assign t[2896] = t[2895] ^ n[2896];
assign t[2897] = t[2896] ^ n[2897];
assign t[2898] = t[2897] ^ n[2898];
assign t[2899] = t[2898] ^ n[2899];
assign t[2900] = t[2899] ^ n[2900];
assign t[2901] = t[2900] ^ n[2901];
assign t[2902] = t[2901] ^ n[2902];
assign t[2903] = t[2902] ^ n[2903];
assign t[2904] = t[2903] ^ n[2904];
assign t[2905] = t[2904] ^ n[2905];
assign t[2906] = t[2905] ^ n[2906];
assign t[2907] = t[2906] ^ n[2907];
assign t[2908] = t[2907] ^ n[2908];
assign t[2909] = t[2908] ^ n[2909];
assign t[2910] = t[2909] ^ n[2910];
assign t[2911] = t[2910] ^ n[2911];
assign t[2912] = t[2911] ^ n[2912];
assign t[2913] = t[2912] ^ n[2913];
assign t[2914] = t[2913] ^ n[2914];
assign t[2915] = t[2914] ^ n[2915];
assign t[2916] = t[2915] ^ n[2916];
assign t[2917] = t[2916] ^ n[2917];
assign t[2918] = t[2917] ^ n[2918];
assign t[2919] = t[2918] ^ n[2919];
assign t[2920] = t[2919] ^ n[2920];
assign t[2921] = t[2920] ^ n[2921];
assign t[2922] = t[2921] ^ n[2922];
assign t[2923] = t[2922] ^ n[2923];
assign t[2924] = t[2923] ^ n[2924];
assign t[2925] = t[2924] ^ n[2925];
assign t[2926] = t[2925] ^ n[2926];
assign t[2927] = t[2926] ^ n[2927];
assign t[2928] = t[2927] ^ n[2928];
assign t[2929] = t[2928] ^ n[2929];
assign t[2930] = t[2929] ^ n[2930];
assign t[2931] = t[2930] ^ n[2931];
assign t[2932] = t[2931] ^ n[2932];
assign t[2933] = t[2932] ^ n[2933];
assign t[2934] = t[2933] ^ n[2934];
assign t[2935] = t[2934] ^ n[2935];
assign t[2936] = t[2935] ^ n[2936];
assign t[2937] = t[2936] ^ n[2937];
assign t[2938] = t[2937] ^ n[2938];
assign t[2939] = t[2938] ^ n[2939];
assign t[2940] = t[2939] ^ n[2940];
assign t[2941] = t[2940] ^ n[2941];
assign t[2942] = t[2941] ^ n[2942];
assign t[2943] = t[2942] ^ n[2943];
assign t[2944] = t[2943] ^ n[2944];
assign t[2945] = t[2944] ^ n[2945];
assign t[2946] = t[2945] ^ n[2946];
assign t[2947] = t[2946] ^ n[2947];
assign t[2948] = t[2947] ^ n[2948];
assign t[2949] = t[2948] ^ n[2949];
assign t[2950] = t[2949] ^ n[2950];
assign t[2951] = t[2950] ^ n[2951];
assign t[2952] = t[2951] ^ n[2952];
assign t[2953] = t[2952] ^ n[2953];
assign t[2954] = t[2953] ^ n[2954];
assign t[2955] = t[2954] ^ n[2955];
assign t[2956] = t[2955] ^ n[2956];
assign t[2957] = t[2956] ^ n[2957];
assign t[2958] = t[2957] ^ n[2958];
assign t[2959] = t[2958] ^ n[2959];
assign t[2960] = t[2959] ^ n[2960];
assign t[2961] = t[2960] ^ n[2961];
assign t[2962] = t[2961] ^ n[2962];
assign t[2963] = t[2962] ^ n[2963];
assign t[2964] = t[2963] ^ n[2964];
assign t[2965] = t[2964] ^ n[2965];
assign t[2966] = t[2965] ^ n[2966];
assign t[2967] = t[2966] ^ n[2967];
assign t[2968] = t[2967] ^ n[2968];
assign t[2969] = t[2968] ^ n[2969];
assign t[2970] = t[2969] ^ n[2970];
assign t[2971] = t[2970] ^ n[2971];
assign t[2972] = t[2971] ^ n[2972];
assign t[2973] = t[2972] ^ n[2973];
assign t[2974] = t[2973] ^ n[2974];
assign t[2975] = t[2974] ^ n[2975];
assign t[2976] = t[2975] ^ n[2976];
assign t[2977] = t[2976] ^ n[2977];
assign t[2978] = t[2977] ^ n[2978];
assign t[2979] = t[2978] ^ n[2979];
assign t[2980] = t[2979] ^ n[2980];
assign t[2981] = t[2980] ^ n[2981];
assign t[2982] = t[2981] ^ n[2982];
assign t[2983] = t[2982] ^ n[2983];
assign t[2984] = t[2983] ^ n[2984];
assign t[2985] = t[2984] ^ n[2985];
assign t[2986] = t[2985] ^ n[2986];
assign t[2987] = t[2986] ^ n[2987];
assign t[2988] = t[2987] ^ n[2988];
assign t[2989] = t[2988] ^ n[2989];
assign t[2990] = t[2989] ^ n[2990];
assign t[2991] = t[2990] ^ n[2991];
assign t[2992] = t[2991] ^ n[2992];
assign t[2993] = t[2992] ^ n[2993];
assign t[2994] = t[2993] ^ n[2994];
assign t[2995] = t[2994] ^ n[2995];
assign t[2996] = t[2995] ^ n[2996];
assign t[2997] = t[2996] ^ n[2997];
assign t[2998] = t[2997] ^ n[2998];
assign t[2999] = t[2998] ^ n[2999];
assign t[3000] = t[2999] ^ n[3000];
assign t[3001] = t[3000] ^ n[3001];
assign t[3002] = t[3001] ^ n[3002];
assign t[3003] = t[3002] ^ n[3003];
assign t[3004] = t[3003] ^ n[3004];
assign t[3005] = t[3004] ^ n[3005];
assign t[3006] = t[3005] ^ n[3006];
assign t[3007] = t[3006] ^ n[3007];
assign t[3008] = t[3007] ^ n[3008];
assign t[3009] = t[3008] ^ n[3009];
assign t[3010] = t[3009] ^ n[3010];
assign t[3011] = t[3010] ^ n[3011];
assign t[3012] = t[3011] ^ n[3012];
assign t[3013] = t[3012] ^ n[3013];
assign t[3014] = t[3013] ^ n[3014];
assign t[3015] = t[3014] ^ n[3015];
assign t[3016] = t[3015] ^ n[3016];
assign t[3017] = t[3016] ^ n[3017];
assign t[3018] = t[3017] ^ n[3018];
assign t[3019] = t[3018] ^ n[3019];
assign t[3020] = t[3019] ^ n[3020];
assign t[3021] = t[3020] ^ n[3021];
assign t[3022] = t[3021] ^ n[3022];
assign t[3023] = t[3022] ^ n[3023];
assign t[3024] = t[3023] ^ n[3024];
assign t[3025] = t[3024] ^ n[3025];
assign t[3026] = t[3025] ^ n[3026];
assign t[3027] = t[3026] ^ n[3027];
assign t[3028] = t[3027] ^ n[3028];
assign t[3029] = t[3028] ^ n[3029];
assign t[3030] = t[3029] ^ n[3030];
assign t[3031] = t[3030] ^ n[3031];
assign t[3032] = t[3031] ^ n[3032];
assign t[3033] = t[3032] ^ n[3033];
assign t[3034] = t[3033] ^ n[3034];
assign t[3035] = t[3034] ^ n[3035];
assign t[3036] = t[3035] ^ n[3036];
assign t[3037] = t[3036] ^ n[3037];
assign t[3038] = t[3037] ^ n[3038];
assign t[3039] = t[3038] ^ n[3039];
assign t[3040] = t[3039] ^ n[3040];
assign t[3041] = t[3040] ^ n[3041];
assign t[3042] = t[3041] ^ n[3042];
assign t[3043] = t[3042] ^ n[3043];
assign t[3044] = t[3043] ^ n[3044];
assign t[3045] = t[3044] ^ n[3045];
assign t[3046] = t[3045] ^ n[3046];
assign t[3047] = t[3046] ^ n[3047];
assign t[3048] = t[3047] ^ n[3048];
assign t[3049] = t[3048] ^ n[3049];
assign t[3050] = t[3049] ^ n[3050];
assign t[3051] = t[3050] ^ n[3051];
assign t[3052] = t[3051] ^ n[3052];
assign t[3053] = t[3052] ^ n[3053];
assign t[3054] = t[3053] ^ n[3054];
assign t[3055] = t[3054] ^ n[3055];
assign t[3056] = t[3055] ^ n[3056];
assign t[3057] = t[3056] ^ n[3057];
assign t[3058] = t[3057] ^ n[3058];
assign t[3059] = t[3058] ^ n[3059];
assign t[3060] = t[3059] ^ n[3060];
assign t[3061] = t[3060] ^ n[3061];
assign t[3062] = t[3061] ^ n[3062];
assign t[3063] = t[3062] ^ n[3063];
assign t[3064] = t[3063] ^ n[3064];
assign t[3065] = t[3064] ^ n[3065];
assign t[3066] = t[3065] ^ n[3066];
assign t[3067] = t[3066] ^ n[3067];
assign t[3068] = t[3067] ^ n[3068];
assign t[3069] = t[3068] ^ n[3069];
assign t[3070] = t[3069] ^ n[3070];
assign t[3071] = t[3070] ^ n[3071];
assign t[3072] = t[3071] ^ n[3072];
assign t[3073] = t[3072] ^ n[3073];
assign t[3074] = t[3073] ^ n[3074];
assign t[3075] = t[3074] ^ n[3075];
assign t[3076] = t[3075] ^ n[3076];
assign t[3077] = t[3076] ^ n[3077];
assign t[3078] = t[3077] ^ n[3078];
assign t[3079] = t[3078] ^ n[3079];
assign t[3080] = t[3079] ^ n[3080];
assign t[3081] = t[3080] ^ n[3081];
assign t[3082] = t[3081] ^ n[3082];
assign t[3083] = t[3082] ^ n[3083];
assign t[3084] = t[3083] ^ n[3084];
assign t[3085] = t[3084] ^ n[3085];
assign t[3086] = t[3085] ^ n[3086];
assign t[3087] = t[3086] ^ n[3087];
assign t[3088] = t[3087] ^ n[3088];
assign t[3089] = t[3088] ^ n[3089];
assign t[3090] = t[3089] ^ n[3090];
assign t[3091] = t[3090] ^ n[3091];
assign t[3092] = t[3091] ^ n[3092];
assign t[3093] = t[3092] ^ n[3093];
assign t[3094] = t[3093] ^ n[3094];
assign t[3095] = t[3094] ^ n[3095];
assign t[3096] = t[3095] ^ n[3096];
assign t[3097] = t[3096] ^ n[3097];
assign t[3098] = t[3097] ^ n[3098];
assign t[3099] = t[3098] ^ n[3099];
assign t[3100] = t[3099] ^ n[3100];
assign t[3101] = t[3100] ^ n[3101];
assign t[3102] = t[3101] ^ n[3102];
assign t[3103] = t[3102] ^ n[3103];
assign t[3104] = t[3103] ^ n[3104];
assign t[3105] = t[3104] ^ n[3105];
assign t[3106] = t[3105] ^ n[3106];
assign t[3107] = t[3106] ^ n[3107];
assign t[3108] = t[3107] ^ n[3108];
assign t[3109] = t[3108] ^ n[3109];
assign t[3110] = t[3109] ^ n[3110];
assign t[3111] = t[3110] ^ n[3111];
assign t[3112] = t[3111] ^ n[3112];
assign t[3113] = t[3112] ^ n[3113];
assign t[3114] = t[3113] ^ n[3114];
assign t[3115] = t[3114] ^ n[3115];
assign t[3116] = t[3115] ^ n[3116];
assign t[3117] = t[3116] ^ n[3117];
assign t[3118] = t[3117] ^ n[3118];
assign t[3119] = t[3118] ^ n[3119];
assign t[3120] = t[3119] ^ n[3120];
assign t[3121] = t[3120] ^ n[3121];
assign t[3122] = t[3121] ^ n[3122];
assign t[3123] = t[3122] ^ n[3123];
assign t[3124] = t[3123] ^ n[3124];
assign t[3125] = t[3124] ^ n[3125];
assign t[3126] = t[3125] ^ n[3126];
assign t[3127] = t[3126] ^ n[3127];
assign t[3128] = t[3127] ^ n[3128];
assign t[3129] = t[3128] ^ n[3129];
assign t[3130] = t[3129] ^ n[3130];
assign t[3131] = t[3130] ^ n[3131];
assign t[3132] = t[3131] ^ n[3132];
assign t[3133] = t[3132] ^ n[3133];
assign t[3134] = t[3133] ^ n[3134];
assign t[3135] = t[3134] ^ n[3135];
assign t[3136] = t[3135] ^ n[3136];
assign t[3137] = t[3136] ^ n[3137];
assign t[3138] = t[3137] ^ n[3138];
assign t[3139] = t[3138] ^ n[3139];
assign t[3140] = t[3139] ^ n[3140];
assign t[3141] = t[3140] ^ n[3141];
assign t[3142] = t[3141] ^ n[3142];
assign t[3143] = t[3142] ^ n[3143];
assign t[3144] = t[3143] ^ n[3144];
assign t[3145] = t[3144] ^ n[3145];
assign t[3146] = t[3145] ^ n[3146];
assign t[3147] = t[3146] ^ n[3147];
assign t[3148] = t[3147] ^ n[3148];
assign t[3149] = t[3148] ^ n[3149];
assign t[3150] = t[3149] ^ n[3150];
assign t[3151] = t[3150] ^ n[3151];
assign t[3152] = t[3151] ^ n[3152];
assign t[3153] = t[3152] ^ n[3153];
assign t[3154] = t[3153] ^ n[3154];
assign t[3155] = t[3154] ^ n[3155];
assign t[3156] = t[3155] ^ n[3156];
assign t[3157] = t[3156] ^ n[3157];
assign t[3158] = t[3157] ^ n[3158];
assign t[3159] = t[3158] ^ n[3159];
assign t[3160] = t[3159] ^ n[3160];
assign t[3161] = t[3160] ^ n[3161];
assign t[3162] = t[3161] ^ n[3162];
assign t[3163] = t[3162] ^ n[3163];
assign t[3164] = t[3163] ^ n[3164];
assign t[3165] = t[3164] ^ n[3165];
assign t[3166] = t[3165] ^ n[3166];
assign t[3167] = t[3166] ^ n[3167];
assign t[3168] = t[3167] ^ n[3168];
assign t[3169] = t[3168] ^ n[3169];
assign t[3170] = t[3169] ^ n[3170];
assign t[3171] = t[3170] ^ n[3171];
assign t[3172] = t[3171] ^ n[3172];
assign t[3173] = t[3172] ^ n[3173];
assign t[3174] = t[3173] ^ n[3174];
assign t[3175] = t[3174] ^ n[3175];
assign t[3176] = t[3175] ^ n[3176];
assign t[3177] = t[3176] ^ n[3177];
assign t[3178] = t[3177] ^ n[3178];
assign t[3179] = t[3178] ^ n[3179];
assign t[3180] = t[3179] ^ n[3180];
assign t[3181] = t[3180] ^ n[3181];
assign t[3182] = t[3181] ^ n[3182];
assign t[3183] = t[3182] ^ n[3183];
assign t[3184] = t[3183] ^ n[3184];
assign t[3185] = t[3184] ^ n[3185];
assign t[3186] = t[3185] ^ n[3186];
assign t[3187] = t[3186] ^ n[3187];
assign t[3188] = t[3187] ^ n[3188];
assign t[3189] = t[3188] ^ n[3189];
assign t[3190] = t[3189] ^ n[3190];
assign t[3191] = t[3190] ^ n[3191];
assign t[3192] = t[3191] ^ n[3192];
assign t[3193] = t[3192] ^ n[3193];
assign t[3194] = t[3193] ^ n[3194];
assign t[3195] = t[3194] ^ n[3195];
assign t[3196] = t[3195] ^ n[3196];
assign t[3197] = t[3196] ^ n[3197];
assign t[3198] = t[3197] ^ n[3198];
assign t[3199] = t[3198] ^ n[3199];
assign t[3200] = t[3199] ^ n[3200];
assign t[3201] = t[3200] ^ n[3201];
assign t[3202] = t[3201] ^ n[3202];
assign t[3203] = t[3202] ^ n[3203];
assign t[3204] = t[3203] ^ n[3204];
assign t[3205] = t[3204] ^ n[3205];
assign t[3206] = t[3205] ^ n[3206];
assign t[3207] = t[3206] ^ n[3207];
assign t[3208] = t[3207] ^ n[3208];
assign t[3209] = t[3208] ^ n[3209];
assign t[3210] = t[3209] ^ n[3210];
assign t[3211] = t[3210] ^ n[3211];
assign t[3212] = t[3211] ^ n[3212];
assign t[3213] = t[3212] ^ n[3213];
assign t[3214] = t[3213] ^ n[3214];
assign t[3215] = t[3214] ^ n[3215];
assign t[3216] = t[3215] ^ n[3216];
assign t[3217] = t[3216] ^ n[3217];
assign t[3218] = t[3217] ^ n[3218];
assign t[3219] = t[3218] ^ n[3219];
assign t[3220] = t[3219] ^ n[3220];
assign t[3221] = t[3220] ^ n[3221];
assign t[3222] = t[3221] ^ n[3222];
assign t[3223] = t[3222] ^ n[3223];
assign t[3224] = t[3223] ^ n[3224];
assign t[3225] = t[3224] ^ n[3225];
assign t[3226] = t[3225] ^ n[3226];
assign t[3227] = t[3226] ^ n[3227];
assign t[3228] = t[3227] ^ n[3228];
assign t[3229] = t[3228] ^ n[3229];
assign t[3230] = t[3229] ^ n[3230];
assign t[3231] = t[3230] ^ n[3231];
assign t[3232] = t[3231] ^ n[3232];
assign t[3233] = t[3232] ^ n[3233];
assign t[3234] = t[3233] ^ n[3234];
assign t[3235] = t[3234] ^ n[3235];
assign t[3236] = t[3235] ^ n[3236];
assign t[3237] = t[3236] ^ n[3237];
assign t[3238] = t[3237] ^ n[3238];
assign t[3239] = t[3238] ^ n[3239];
assign t[3240] = t[3239] ^ n[3240];
assign t[3241] = t[3240] ^ n[3241];
assign t[3242] = t[3241] ^ n[3242];
assign t[3243] = t[3242] ^ n[3243];
assign t[3244] = t[3243] ^ n[3244];
assign t[3245] = t[3244] ^ n[3245];
assign t[3246] = t[3245] ^ n[3246];
assign t[3247] = t[3246] ^ n[3247];
assign t[3248] = t[3247] ^ n[3248];
assign t[3249] = t[3248] ^ n[3249];
assign t[3250] = t[3249] ^ n[3250];
assign t[3251] = t[3250] ^ n[3251];
assign t[3252] = t[3251] ^ n[3252];
assign t[3253] = t[3252] ^ n[3253];
assign t[3254] = t[3253] ^ n[3254];
assign t[3255] = t[3254] ^ n[3255];
assign t[3256] = t[3255] ^ n[3256];
assign t[3257] = t[3256] ^ n[3257];
assign t[3258] = t[3257] ^ n[3258];
assign t[3259] = t[3258] ^ n[3259];
assign t[3260] = t[3259] ^ n[3260];
assign t[3261] = t[3260] ^ n[3261];
assign t[3262] = t[3261] ^ n[3262];
assign t[3263] = t[3262] ^ n[3263];
assign t[3264] = t[3263] ^ n[3264];
assign t[3265] = t[3264] ^ n[3265];
assign t[3266] = t[3265] ^ n[3266];
assign t[3267] = t[3266] ^ n[3267];
assign t[3268] = t[3267] ^ n[3268];
assign t[3269] = t[3268] ^ n[3269];
assign t[3270] = t[3269] ^ n[3270];
assign t[3271] = t[3270] ^ n[3271];
assign t[3272] = t[3271] ^ n[3272];
assign t[3273] = t[3272] ^ n[3273];
assign t[3274] = t[3273] ^ n[3274];
assign t[3275] = t[3274] ^ n[3275];
assign t[3276] = t[3275] ^ n[3276];
assign t[3277] = t[3276] ^ n[3277];
assign t[3278] = t[3277] ^ n[3278];
assign t[3279] = t[3278] ^ n[3279];
assign t[3280] = t[3279] ^ n[3280];
assign t[3281] = t[3280] ^ n[3281];
assign t[3282] = t[3281] ^ n[3282];
assign t[3283] = t[3282] ^ n[3283];
assign t[3284] = t[3283] ^ n[3284];
assign t[3285] = t[3284] ^ n[3285];
assign t[3286] = t[3285] ^ n[3286];
assign t[3287] = t[3286] ^ n[3287];
assign t[3288] = t[3287] ^ n[3288];
assign t[3289] = t[3288] ^ n[3289];
assign t[3290] = t[3289] ^ n[3290];
assign t[3291] = t[3290] ^ n[3291];
assign t[3292] = t[3291] ^ n[3292];
assign t[3293] = t[3292] ^ n[3293];
assign t[3294] = t[3293] ^ n[3294];
assign t[3295] = t[3294] ^ n[3295];
assign t[3296] = t[3295] ^ n[3296];
assign t[3297] = t[3296] ^ n[3297];
assign t[3298] = t[3297] ^ n[3298];
assign t[3299] = t[3298] ^ n[3299];
assign t[3300] = t[3299] ^ n[3300];
assign t[3301] = t[3300] ^ n[3301];
assign t[3302] = t[3301] ^ n[3302];
assign t[3303] = t[3302] ^ n[3303];
assign t[3304] = t[3303] ^ n[3304];
assign t[3305] = t[3304] ^ n[3305];
assign t[3306] = t[3305] ^ n[3306];
assign t[3307] = t[3306] ^ n[3307];
assign t[3308] = t[3307] ^ n[3308];
assign t[3309] = t[3308] ^ n[3309];
assign t[3310] = t[3309] ^ n[3310];
assign t[3311] = t[3310] ^ n[3311];
assign t[3312] = t[3311] ^ n[3312];
assign t[3313] = t[3312] ^ n[3313];
assign t[3314] = t[3313] ^ n[3314];
assign t[3315] = t[3314] ^ n[3315];
assign t[3316] = t[3315] ^ n[3316];
assign t[3317] = t[3316] ^ n[3317];
assign t[3318] = t[3317] ^ n[3318];
assign t[3319] = t[3318] ^ n[3319];
assign t[3320] = t[3319] ^ n[3320];
assign t[3321] = t[3320] ^ n[3321];
assign t[3322] = t[3321] ^ n[3322];
assign t[3323] = t[3322] ^ n[3323];
assign t[3324] = t[3323] ^ n[3324];
assign t[3325] = t[3324] ^ n[3325];
assign t[3326] = t[3325] ^ n[3326];
assign t[3327] = t[3326] ^ n[3327];
assign t[3328] = t[3327] ^ n[3328];
assign t[3329] = t[3328] ^ n[3329];
assign t[3330] = t[3329] ^ n[3330];
assign t[3331] = t[3330] ^ n[3331];
assign t[3332] = t[3331] ^ n[3332];
assign t[3333] = t[3332] ^ n[3333];
assign t[3334] = t[3333] ^ n[3334];
assign t[3335] = t[3334] ^ n[3335];
assign t[3336] = t[3335] ^ n[3336];
assign t[3337] = t[3336] ^ n[3337];
assign t[3338] = t[3337] ^ n[3338];
assign t[3339] = t[3338] ^ n[3339];
assign t[3340] = t[3339] ^ n[3340];
assign t[3341] = t[3340] ^ n[3341];
assign t[3342] = t[3341] ^ n[3342];
assign t[3343] = t[3342] ^ n[3343];
assign t[3344] = t[3343] ^ n[3344];
assign t[3345] = t[3344] ^ n[3345];
assign t[3346] = t[3345] ^ n[3346];
assign t[3347] = t[3346] ^ n[3347];
assign t[3348] = t[3347] ^ n[3348];
assign t[3349] = t[3348] ^ n[3349];
assign t[3350] = t[3349] ^ n[3350];
assign t[3351] = t[3350] ^ n[3351];
assign t[3352] = t[3351] ^ n[3352];
assign t[3353] = t[3352] ^ n[3353];
assign t[3354] = t[3353] ^ n[3354];
assign t[3355] = t[3354] ^ n[3355];
assign t[3356] = t[3355] ^ n[3356];
assign t[3357] = t[3356] ^ n[3357];
assign t[3358] = t[3357] ^ n[3358];
assign t[3359] = t[3358] ^ n[3359];
assign t[3360] = t[3359] ^ n[3360];
assign t[3361] = t[3360] ^ n[3361];
assign t[3362] = t[3361] ^ n[3362];
assign t[3363] = t[3362] ^ n[3363];
assign t[3364] = t[3363] ^ n[3364];
assign t[3365] = t[3364] ^ n[3365];
assign t[3366] = t[3365] ^ n[3366];
assign t[3367] = t[3366] ^ n[3367];
assign t[3368] = t[3367] ^ n[3368];
assign t[3369] = t[3368] ^ n[3369];
assign t[3370] = t[3369] ^ n[3370];
assign t[3371] = t[3370] ^ n[3371];
assign t[3372] = t[3371] ^ n[3372];
assign t[3373] = t[3372] ^ n[3373];
assign t[3374] = t[3373] ^ n[3374];
assign t[3375] = t[3374] ^ n[3375];
assign t[3376] = t[3375] ^ n[3376];
assign t[3377] = t[3376] ^ n[3377];
assign t[3378] = t[3377] ^ n[3378];
assign t[3379] = t[3378] ^ n[3379];
assign t[3380] = t[3379] ^ n[3380];
assign t[3381] = t[3380] ^ n[3381];
assign t[3382] = t[3381] ^ n[3382];
assign t[3383] = t[3382] ^ n[3383];
assign t[3384] = t[3383] ^ n[3384];
assign t[3385] = t[3384] ^ n[3385];
assign t[3386] = t[3385] ^ n[3386];
assign t[3387] = t[3386] ^ n[3387];
assign t[3388] = t[3387] ^ n[3388];
assign t[3389] = t[3388] ^ n[3389];
assign t[3390] = t[3389] ^ n[3390];
assign t[3391] = t[3390] ^ n[3391];
assign t[3392] = t[3391] ^ n[3392];
assign t[3393] = t[3392] ^ n[3393];
assign t[3394] = t[3393] ^ n[3394];
assign t[3395] = t[3394] ^ n[3395];
assign t[3396] = t[3395] ^ n[3396];
assign t[3397] = t[3396] ^ n[3397];
assign t[3398] = t[3397] ^ n[3398];
assign t[3399] = t[3398] ^ n[3399];
assign t[3400] = t[3399] ^ n[3400];
assign t[3401] = t[3400] ^ n[3401];
assign t[3402] = t[3401] ^ n[3402];
assign t[3403] = t[3402] ^ n[3403];
assign t[3404] = t[3403] ^ n[3404];
assign t[3405] = t[3404] ^ n[3405];
assign t[3406] = t[3405] ^ n[3406];
assign t[3407] = t[3406] ^ n[3407];
assign t[3408] = t[3407] ^ n[3408];
assign t[3409] = t[3408] ^ n[3409];
assign t[3410] = t[3409] ^ n[3410];
assign t[3411] = t[3410] ^ n[3411];
assign t[3412] = t[3411] ^ n[3412];
assign t[3413] = t[3412] ^ n[3413];
assign t[3414] = t[3413] ^ n[3414];
assign t[3415] = t[3414] ^ n[3415];
assign t[3416] = t[3415] ^ n[3416];
assign t[3417] = t[3416] ^ n[3417];
assign t[3418] = t[3417] ^ n[3418];
assign t[3419] = t[3418] ^ n[3419];
assign t[3420] = t[3419] ^ n[3420];
assign t[3421] = t[3420] ^ n[3421];
assign t[3422] = t[3421] ^ n[3422];
assign t[3423] = t[3422] ^ n[3423];
assign t[3424] = t[3423] ^ n[3424];
assign t[3425] = t[3424] ^ n[3425];
assign t[3426] = t[3425] ^ n[3426];
assign t[3427] = t[3426] ^ n[3427];
assign t[3428] = t[3427] ^ n[3428];
assign t[3429] = t[3428] ^ n[3429];
assign t[3430] = t[3429] ^ n[3430];
assign t[3431] = t[3430] ^ n[3431];
assign t[3432] = t[3431] ^ n[3432];
assign t[3433] = t[3432] ^ n[3433];
assign t[3434] = t[3433] ^ n[3434];
assign t[3435] = t[3434] ^ n[3435];
assign t[3436] = t[3435] ^ n[3436];
assign t[3437] = t[3436] ^ n[3437];
assign t[3438] = t[3437] ^ n[3438];
assign t[3439] = t[3438] ^ n[3439];
assign t[3440] = t[3439] ^ n[3440];
assign t[3441] = t[3440] ^ n[3441];
assign t[3442] = t[3441] ^ n[3442];
assign t[3443] = t[3442] ^ n[3443];
assign t[3444] = t[3443] ^ n[3444];
assign t[3445] = t[3444] ^ n[3445];
assign t[3446] = t[3445] ^ n[3446];
assign t[3447] = t[3446] ^ n[3447];
assign t[3448] = t[3447] ^ n[3448];
assign t[3449] = t[3448] ^ n[3449];
assign t[3450] = t[3449] ^ n[3450];
assign t[3451] = t[3450] ^ n[3451];
assign t[3452] = t[3451] ^ n[3452];
assign t[3453] = t[3452] ^ n[3453];
assign t[3454] = t[3453] ^ n[3454];
assign t[3455] = t[3454] ^ n[3455];
assign t[3456] = t[3455] ^ n[3456];
assign t[3457] = t[3456] ^ n[3457];
assign t[3458] = t[3457] ^ n[3458];
assign t[3459] = t[3458] ^ n[3459];
assign t[3460] = t[3459] ^ n[3460];
assign t[3461] = t[3460] ^ n[3461];
assign t[3462] = t[3461] ^ n[3462];
assign t[3463] = t[3462] ^ n[3463];
assign t[3464] = t[3463] ^ n[3464];
assign t[3465] = t[3464] ^ n[3465];
assign t[3466] = t[3465] ^ n[3466];
assign t[3467] = t[3466] ^ n[3467];
assign t[3468] = t[3467] ^ n[3468];
assign t[3469] = t[3468] ^ n[3469];
assign t[3470] = t[3469] ^ n[3470];
assign t[3471] = t[3470] ^ n[3471];
assign t[3472] = t[3471] ^ n[3472];
assign t[3473] = t[3472] ^ n[3473];
assign t[3474] = t[3473] ^ n[3474];
assign t[3475] = t[3474] ^ n[3475];
assign t[3476] = t[3475] ^ n[3476];
assign t[3477] = t[3476] ^ n[3477];
assign t[3478] = t[3477] ^ n[3478];
assign t[3479] = t[3478] ^ n[3479];
assign t[3480] = t[3479] ^ n[3480];
assign t[3481] = t[3480] ^ n[3481];
assign t[3482] = t[3481] ^ n[3482];
assign t[3483] = t[3482] ^ n[3483];
assign t[3484] = t[3483] ^ n[3484];
assign t[3485] = t[3484] ^ n[3485];
assign t[3486] = t[3485] ^ n[3486];
assign t[3487] = t[3486] ^ n[3487];
assign t[3488] = t[3487] ^ n[3488];
assign t[3489] = t[3488] ^ n[3489];
assign t[3490] = t[3489] ^ n[3490];
assign t[3491] = t[3490] ^ n[3491];
assign t[3492] = t[3491] ^ n[3492];
assign t[3493] = t[3492] ^ n[3493];
assign t[3494] = t[3493] ^ n[3494];
assign t[3495] = t[3494] ^ n[3495];
assign t[3496] = t[3495] ^ n[3496];
assign t[3497] = t[3496] ^ n[3497];
assign t[3498] = t[3497] ^ n[3498];
assign t[3499] = t[3498] ^ n[3499];
assign t[3500] = t[3499] ^ n[3500];
assign t[3501] = t[3500] ^ n[3501];
assign t[3502] = t[3501] ^ n[3502];
assign t[3503] = t[3502] ^ n[3503];
assign t[3504] = t[3503] ^ n[3504];
assign t[3505] = t[3504] ^ n[3505];
assign t[3506] = t[3505] ^ n[3506];
assign t[3507] = t[3506] ^ n[3507];
assign t[3508] = t[3507] ^ n[3508];
assign t[3509] = t[3508] ^ n[3509];
assign t[3510] = t[3509] ^ n[3510];
assign t[3511] = t[3510] ^ n[3511];
assign t[3512] = t[3511] ^ n[3512];
assign t[3513] = t[3512] ^ n[3513];
assign t[3514] = t[3513] ^ n[3514];
assign t[3515] = t[3514] ^ n[3515];
assign t[3516] = t[3515] ^ n[3516];
assign t[3517] = t[3516] ^ n[3517];
assign t[3518] = t[3517] ^ n[3518];
assign t[3519] = t[3518] ^ n[3519];
assign t[3520] = t[3519] ^ n[3520];
assign t[3521] = t[3520] ^ n[3521];
assign t[3522] = t[3521] ^ n[3522];
assign t[3523] = t[3522] ^ n[3523];
assign t[3524] = t[3523] ^ n[3524];
assign t[3525] = t[3524] ^ n[3525];
assign t[3526] = t[3525] ^ n[3526];
assign t[3527] = t[3526] ^ n[3527];
assign t[3528] = t[3527] ^ n[3528];
assign t[3529] = t[3528] ^ n[3529];
assign t[3530] = t[3529] ^ n[3530];
assign t[3531] = t[3530] ^ n[3531];
assign t[3532] = t[3531] ^ n[3532];
assign t[3533] = t[3532] ^ n[3533];
assign t[3534] = t[3533] ^ n[3534];
assign t[3535] = t[3534] ^ n[3535];
assign t[3536] = t[3535] ^ n[3536];
assign t[3537] = t[3536] ^ n[3537];
assign t[3538] = t[3537] ^ n[3538];
assign t[3539] = t[3538] ^ n[3539];
assign t[3540] = t[3539] ^ n[3540];
assign t[3541] = t[3540] ^ n[3541];
assign t[3542] = t[3541] ^ n[3542];
assign t[3543] = t[3542] ^ n[3543];
assign t[3544] = t[3543] ^ n[3544];
assign t[3545] = t[3544] ^ n[3545];
assign t[3546] = t[3545] ^ n[3546];
assign t[3547] = t[3546] ^ n[3547];
assign t[3548] = t[3547] ^ n[3548];
assign t[3549] = t[3548] ^ n[3549];
assign t[3550] = t[3549] ^ n[3550];
assign t[3551] = t[3550] ^ n[3551];
assign t[3552] = t[3551] ^ n[3552];
assign t[3553] = t[3552] ^ n[3553];
assign t[3554] = t[3553] ^ n[3554];
assign t[3555] = t[3554] ^ n[3555];
assign t[3556] = t[3555] ^ n[3556];
assign t[3557] = t[3556] ^ n[3557];
assign t[3558] = t[3557] ^ n[3558];
assign t[3559] = t[3558] ^ n[3559];
assign t[3560] = t[3559] ^ n[3560];
assign t[3561] = t[3560] ^ n[3561];
assign t[3562] = t[3561] ^ n[3562];
assign t[3563] = t[3562] ^ n[3563];
assign t[3564] = t[3563] ^ n[3564];
assign t[3565] = t[3564] ^ n[3565];
assign t[3566] = t[3565] ^ n[3566];
assign t[3567] = t[3566] ^ n[3567];
assign t[3568] = t[3567] ^ n[3568];
assign t[3569] = t[3568] ^ n[3569];
assign t[3570] = t[3569] ^ n[3570];
assign t[3571] = t[3570] ^ n[3571];
assign t[3572] = t[3571] ^ n[3572];
assign t[3573] = t[3572] ^ n[3573];
assign t[3574] = t[3573] ^ n[3574];
assign t[3575] = t[3574] ^ n[3575];
assign t[3576] = t[3575] ^ n[3576];
assign t[3577] = t[3576] ^ n[3577];
assign t[3578] = t[3577] ^ n[3578];
assign t[3579] = t[3578] ^ n[3579];
assign t[3580] = t[3579] ^ n[3580];
assign t[3581] = t[3580] ^ n[3581];
assign t[3582] = t[3581] ^ n[3582];
assign t[3583] = t[3582] ^ n[3583];
assign t[3584] = t[3583] ^ n[3584];
assign t[3585] = t[3584] ^ n[3585];
assign t[3586] = t[3585] ^ n[3586];
assign t[3587] = t[3586] ^ n[3587];
assign t[3588] = t[3587] ^ n[3588];
assign t[3589] = t[3588] ^ n[3589];
assign t[3590] = t[3589] ^ n[3590];
assign t[3591] = t[3590] ^ n[3591];
assign t[3592] = t[3591] ^ n[3592];
assign t[3593] = t[3592] ^ n[3593];
assign t[3594] = t[3593] ^ n[3594];
assign t[3595] = t[3594] ^ n[3595];
assign t[3596] = t[3595] ^ n[3596];
assign t[3597] = t[3596] ^ n[3597];
assign t[3598] = t[3597] ^ n[3598];
assign t[3599] = t[3598] ^ n[3599];
assign t[3600] = t[3599] ^ n[3600];
assign t[3601] = t[3600] ^ n[3601];
assign t[3602] = t[3601] ^ n[3602];
assign t[3603] = t[3602] ^ n[3603];
assign t[3604] = t[3603] ^ n[3604];
assign t[3605] = t[3604] ^ n[3605];
assign t[3606] = t[3605] ^ n[3606];
assign t[3607] = t[3606] ^ n[3607];
assign t[3608] = t[3607] ^ n[3608];
assign t[3609] = t[3608] ^ n[3609];
assign t[3610] = t[3609] ^ n[3610];
assign t[3611] = t[3610] ^ n[3611];
assign t[3612] = t[3611] ^ n[3612];
assign t[3613] = t[3612] ^ n[3613];
assign t[3614] = t[3613] ^ n[3614];
assign t[3615] = t[3614] ^ n[3615];
assign t[3616] = t[3615] ^ n[3616];
assign t[3617] = t[3616] ^ n[3617];
assign t[3618] = t[3617] ^ n[3618];
assign t[3619] = t[3618] ^ n[3619];
assign t[3620] = t[3619] ^ n[3620];
assign t[3621] = t[3620] ^ n[3621];
assign t[3622] = t[3621] ^ n[3622];
assign t[3623] = t[3622] ^ n[3623];
assign t[3624] = t[3623] ^ n[3624];
assign t[3625] = t[3624] ^ n[3625];
assign t[3626] = t[3625] ^ n[3626];
assign t[3627] = t[3626] ^ n[3627];
assign t[3628] = t[3627] ^ n[3628];
assign t[3629] = t[3628] ^ n[3629];
assign t[3630] = t[3629] ^ n[3630];
assign t[3631] = t[3630] ^ n[3631];
assign t[3632] = t[3631] ^ n[3632];
assign t[3633] = t[3632] ^ n[3633];
assign t[3634] = t[3633] ^ n[3634];
assign t[3635] = t[3634] ^ n[3635];
assign t[3636] = t[3635] ^ n[3636];
assign t[3637] = t[3636] ^ n[3637];
assign t[3638] = t[3637] ^ n[3638];
assign t[3639] = t[3638] ^ n[3639];
assign t[3640] = t[3639] ^ n[3640];
assign t[3641] = t[3640] ^ n[3641];
assign t[3642] = t[3641] ^ n[3642];
assign t[3643] = t[3642] ^ n[3643];
assign t[3644] = t[3643] ^ n[3644];
assign t[3645] = t[3644] ^ n[3645];
assign t[3646] = t[3645] ^ n[3646];
assign t[3647] = t[3646] ^ n[3647];
assign t[3648] = t[3647] ^ n[3648];
assign t[3649] = t[3648] ^ n[3649];
assign t[3650] = t[3649] ^ n[3650];
assign t[3651] = t[3650] ^ n[3651];
assign t[3652] = t[3651] ^ n[3652];
assign t[3653] = t[3652] ^ n[3653];
assign t[3654] = t[3653] ^ n[3654];
assign t[3655] = t[3654] ^ n[3655];
assign t[3656] = t[3655] ^ n[3656];
assign t[3657] = t[3656] ^ n[3657];
assign t[3658] = t[3657] ^ n[3658];
assign t[3659] = t[3658] ^ n[3659];
assign t[3660] = t[3659] ^ n[3660];
assign t[3661] = t[3660] ^ n[3661];
assign t[3662] = t[3661] ^ n[3662];
assign t[3663] = t[3662] ^ n[3663];
assign t[3664] = t[3663] ^ n[3664];
assign t[3665] = t[3664] ^ n[3665];
assign t[3666] = t[3665] ^ n[3666];
assign t[3667] = t[3666] ^ n[3667];
assign t[3668] = t[3667] ^ n[3668];
assign t[3669] = t[3668] ^ n[3669];
assign t[3670] = t[3669] ^ n[3670];
assign t[3671] = t[3670] ^ n[3671];
assign t[3672] = t[3671] ^ n[3672];
assign t[3673] = t[3672] ^ n[3673];
assign t[3674] = t[3673] ^ n[3674];
assign t[3675] = t[3674] ^ n[3675];
assign t[3676] = t[3675] ^ n[3676];
assign t[3677] = t[3676] ^ n[3677];
assign t[3678] = t[3677] ^ n[3678];
assign t[3679] = t[3678] ^ n[3679];
assign t[3680] = t[3679] ^ n[3680];
assign t[3681] = t[3680] ^ n[3681];
assign t[3682] = t[3681] ^ n[3682];
assign t[3683] = t[3682] ^ n[3683];
assign t[3684] = t[3683] ^ n[3684];
assign t[3685] = t[3684] ^ n[3685];
assign t[3686] = t[3685] ^ n[3686];
assign t[3687] = t[3686] ^ n[3687];
assign t[3688] = t[3687] ^ n[3688];
assign t[3689] = t[3688] ^ n[3689];
assign t[3690] = t[3689] ^ n[3690];
assign t[3691] = t[3690] ^ n[3691];
assign t[3692] = t[3691] ^ n[3692];
assign t[3693] = t[3692] ^ n[3693];
assign t[3694] = t[3693] ^ n[3694];
assign t[3695] = t[3694] ^ n[3695];
assign t[3696] = t[3695] ^ n[3696];
assign t[3697] = t[3696] ^ n[3697];
assign t[3698] = t[3697] ^ n[3698];
assign t[3699] = t[3698] ^ n[3699];
assign t[3700] = t[3699] ^ n[3700];
assign t[3701] = t[3700] ^ n[3701];
assign t[3702] = t[3701] ^ n[3702];
assign t[3703] = t[3702] ^ n[3703];
assign t[3704] = t[3703] ^ n[3704];
assign t[3705] = t[3704] ^ n[3705];
assign t[3706] = t[3705] ^ n[3706];
assign t[3707] = t[3706] ^ n[3707];
assign t[3708] = t[3707] ^ n[3708];
assign t[3709] = t[3708] ^ n[3709];
assign t[3710] = t[3709] ^ n[3710];
assign t[3711] = t[3710] ^ n[3711];
assign t[3712] = t[3711] ^ n[3712];
assign t[3713] = t[3712] ^ n[3713];
assign t[3714] = t[3713] ^ n[3714];
assign t[3715] = t[3714] ^ n[3715];
assign t[3716] = t[3715] ^ n[3716];
assign t[3717] = t[3716] ^ n[3717];
assign t[3718] = t[3717] ^ n[3718];
assign t[3719] = t[3718] ^ n[3719];
assign t[3720] = t[3719] ^ n[3720];
assign t[3721] = t[3720] ^ n[3721];
assign t[3722] = t[3721] ^ n[3722];
assign t[3723] = t[3722] ^ n[3723];
assign t[3724] = t[3723] ^ n[3724];
assign t[3725] = t[3724] ^ n[3725];
assign t[3726] = t[3725] ^ n[3726];
assign t[3727] = t[3726] ^ n[3727];
assign t[3728] = t[3727] ^ n[3728];
assign t[3729] = t[3728] ^ n[3729];
assign t[3730] = t[3729] ^ n[3730];
assign t[3731] = t[3730] ^ n[3731];
assign t[3732] = t[3731] ^ n[3732];
assign t[3733] = t[3732] ^ n[3733];
assign t[3734] = t[3733] ^ n[3734];
assign t[3735] = t[3734] ^ n[3735];
assign t[3736] = t[3735] ^ n[3736];
assign t[3737] = t[3736] ^ n[3737];
assign t[3738] = t[3737] ^ n[3738];
assign t[3739] = t[3738] ^ n[3739];
assign t[3740] = t[3739] ^ n[3740];
assign t[3741] = t[3740] ^ n[3741];
assign t[3742] = t[3741] ^ n[3742];
assign t[3743] = t[3742] ^ n[3743];
assign t[3744] = t[3743] ^ n[3744];
assign t[3745] = t[3744] ^ n[3745];
assign t[3746] = t[3745] ^ n[3746];
assign t[3747] = t[3746] ^ n[3747];
assign t[3748] = t[3747] ^ n[3748];
assign t[3749] = t[3748] ^ n[3749];
assign t[3750] = t[3749] ^ n[3750];
assign t[3751] = t[3750] ^ n[3751];
assign t[3752] = t[3751] ^ n[3752];
assign t[3753] = t[3752] ^ n[3753];
assign t[3754] = t[3753] ^ n[3754];
assign t[3755] = t[3754] ^ n[3755];
assign t[3756] = t[3755] ^ n[3756];
assign t[3757] = t[3756] ^ n[3757];
assign t[3758] = t[3757] ^ n[3758];
assign t[3759] = t[3758] ^ n[3759];
assign t[3760] = t[3759] ^ n[3760];
assign t[3761] = t[3760] ^ n[3761];
assign t[3762] = t[3761] ^ n[3762];
assign t[3763] = t[3762] ^ n[3763];
assign t[3764] = t[3763] ^ n[3764];
assign t[3765] = t[3764] ^ n[3765];
assign t[3766] = t[3765] ^ n[3766];
assign t[3767] = t[3766] ^ n[3767];
assign t[3768] = t[3767] ^ n[3768];
assign t[3769] = t[3768] ^ n[3769];
assign t[3770] = t[3769] ^ n[3770];
assign t[3771] = t[3770] ^ n[3771];
assign t[3772] = t[3771] ^ n[3772];
assign t[3773] = t[3772] ^ n[3773];
assign t[3774] = t[3773] ^ n[3774];
assign t[3775] = t[3774] ^ n[3775];
assign t[3776] = t[3775] ^ n[3776];
assign t[3777] = t[3776] ^ n[3777];
assign t[3778] = t[3777] ^ n[3778];
assign t[3779] = t[3778] ^ n[3779];
assign t[3780] = t[3779] ^ n[3780];
assign t[3781] = t[3780] ^ n[3781];
assign t[3782] = t[3781] ^ n[3782];
assign t[3783] = t[3782] ^ n[3783];
assign t[3784] = t[3783] ^ n[3784];
assign t[3785] = t[3784] ^ n[3785];
assign t[3786] = t[3785] ^ n[3786];
assign t[3787] = t[3786] ^ n[3787];
assign t[3788] = t[3787] ^ n[3788];
assign t[3789] = t[3788] ^ n[3789];
assign t[3790] = t[3789] ^ n[3790];
assign t[3791] = t[3790] ^ n[3791];
assign t[3792] = t[3791] ^ n[3792];
assign t[3793] = t[3792] ^ n[3793];
assign t[3794] = t[3793] ^ n[3794];
assign t[3795] = t[3794] ^ n[3795];
assign t[3796] = t[3795] ^ n[3796];
assign t[3797] = t[3796] ^ n[3797];
assign t[3798] = t[3797] ^ n[3798];
assign t[3799] = t[3798] ^ n[3799];
assign t[3800] = t[3799] ^ n[3800];
assign t[3801] = t[3800] ^ n[3801];
assign t[3802] = t[3801] ^ n[3802];
assign t[3803] = t[3802] ^ n[3803];
assign t[3804] = t[3803] ^ n[3804];
assign t[3805] = t[3804] ^ n[3805];
assign t[3806] = t[3805] ^ n[3806];
assign t[3807] = t[3806] ^ n[3807];
assign t[3808] = t[3807] ^ n[3808];
assign t[3809] = t[3808] ^ n[3809];
assign t[3810] = t[3809] ^ n[3810];
assign t[3811] = t[3810] ^ n[3811];
assign t[3812] = t[3811] ^ n[3812];
assign t[3813] = t[3812] ^ n[3813];
assign t[3814] = t[3813] ^ n[3814];
assign t[3815] = t[3814] ^ n[3815];
assign t[3816] = t[3815] ^ n[3816];
assign t[3817] = t[3816] ^ n[3817];
assign t[3818] = t[3817] ^ n[3818];
assign t[3819] = t[3818] ^ n[3819];
assign t[3820] = t[3819] ^ n[3820];
assign t[3821] = t[3820] ^ n[3821];
assign t[3822] = t[3821] ^ n[3822];
assign t[3823] = t[3822] ^ n[3823];
assign t[3824] = t[3823] ^ n[3824];
assign t[3825] = t[3824] ^ n[3825];
assign t[3826] = t[3825] ^ n[3826];
assign t[3827] = t[3826] ^ n[3827];
assign t[3828] = t[3827] ^ n[3828];
assign t[3829] = t[3828] ^ n[3829];
assign t[3830] = t[3829] ^ n[3830];
assign t[3831] = t[3830] ^ n[3831];
assign t[3832] = t[3831] ^ n[3832];
assign t[3833] = t[3832] ^ n[3833];
assign t[3834] = t[3833] ^ n[3834];
assign t[3835] = t[3834] ^ n[3835];
assign t[3836] = t[3835] ^ n[3836];
assign t[3837] = t[3836] ^ n[3837];
assign t[3838] = t[3837] ^ n[3838];
assign t[3839] = t[3838] ^ n[3839];
assign t[3840] = t[3839] ^ n[3840];
assign t[3841] = t[3840] ^ n[3841];
assign t[3842] = t[3841] ^ n[3842];
assign t[3843] = t[3842] ^ n[3843];
assign t[3844] = t[3843] ^ n[3844];
assign t[3845] = t[3844] ^ n[3845];
assign t[3846] = t[3845] ^ n[3846];
assign t[3847] = t[3846] ^ n[3847];
assign t[3848] = t[3847] ^ n[3848];
assign t[3849] = t[3848] ^ n[3849];
assign t[3850] = t[3849] ^ n[3850];
assign t[3851] = t[3850] ^ n[3851];
assign t[3852] = t[3851] ^ n[3852];
assign t[3853] = t[3852] ^ n[3853];
assign t[3854] = t[3853] ^ n[3854];
assign t[3855] = t[3854] ^ n[3855];
assign t[3856] = t[3855] ^ n[3856];
assign t[3857] = t[3856] ^ n[3857];
assign t[3858] = t[3857] ^ n[3858];
assign t[3859] = t[3858] ^ n[3859];
assign t[3860] = t[3859] ^ n[3860];
assign t[3861] = t[3860] ^ n[3861];
assign t[3862] = t[3861] ^ n[3862];
assign t[3863] = t[3862] ^ n[3863];
assign t[3864] = t[3863] ^ n[3864];
assign t[3865] = t[3864] ^ n[3865];
assign t[3866] = t[3865] ^ n[3866];
assign t[3867] = t[3866] ^ n[3867];
assign t[3868] = t[3867] ^ n[3868];
assign t[3869] = t[3868] ^ n[3869];
assign t[3870] = t[3869] ^ n[3870];
assign t[3871] = t[3870] ^ n[3871];
assign t[3872] = t[3871] ^ n[3872];
assign t[3873] = t[3872] ^ n[3873];
assign t[3874] = t[3873] ^ n[3874];
assign t[3875] = t[3874] ^ n[3875];
assign t[3876] = t[3875] ^ n[3876];
assign t[3877] = t[3876] ^ n[3877];
assign t[3878] = t[3877] ^ n[3878];
assign t[3879] = t[3878] ^ n[3879];
assign t[3880] = t[3879] ^ n[3880];
assign t[3881] = t[3880] ^ n[3881];
assign t[3882] = t[3881] ^ n[3882];
assign t[3883] = t[3882] ^ n[3883];
assign t[3884] = t[3883] ^ n[3884];
assign t[3885] = t[3884] ^ n[3885];
assign t[3886] = t[3885] ^ n[3886];
assign t[3887] = t[3886] ^ n[3887];
assign t[3888] = t[3887] ^ n[3888];
assign t[3889] = t[3888] ^ n[3889];
assign t[3890] = t[3889] ^ n[3890];
assign t[3891] = t[3890] ^ n[3891];
assign t[3892] = t[3891] ^ n[3892];
assign t[3893] = t[3892] ^ n[3893];
assign t[3894] = t[3893] ^ n[3894];
assign t[3895] = t[3894] ^ n[3895];
assign t[3896] = t[3895] ^ n[3896];
assign t[3897] = t[3896] ^ n[3897];
assign t[3898] = t[3897] ^ n[3898];
assign t[3899] = t[3898] ^ n[3899];
assign t[3900] = t[3899] ^ n[3900];
assign t[3901] = t[3900] ^ n[3901];
assign t[3902] = t[3901] ^ n[3902];
assign t[3903] = t[3902] ^ n[3903];
assign t[3904] = t[3903] ^ n[3904];
assign t[3905] = t[3904] ^ n[3905];
assign t[3906] = t[3905] ^ n[3906];
assign t[3907] = t[3906] ^ n[3907];
assign t[3908] = t[3907] ^ n[3908];
assign t[3909] = t[3908] ^ n[3909];
assign t[3910] = t[3909] ^ n[3910];
assign t[3911] = t[3910] ^ n[3911];
assign t[3912] = t[3911] ^ n[3912];
assign t[3913] = t[3912] ^ n[3913];
assign t[3914] = t[3913] ^ n[3914];
assign t[3915] = t[3914] ^ n[3915];
assign t[3916] = t[3915] ^ n[3916];
assign t[3917] = t[3916] ^ n[3917];
assign t[3918] = t[3917] ^ n[3918];
assign t[3919] = t[3918] ^ n[3919];
assign t[3920] = t[3919] ^ n[3920];
assign t[3921] = t[3920] ^ n[3921];
assign t[3922] = t[3921] ^ n[3922];
assign t[3923] = t[3922] ^ n[3923];
assign t[3924] = t[3923] ^ n[3924];
assign t[3925] = t[3924] ^ n[3925];
assign t[3926] = t[3925] ^ n[3926];
assign t[3927] = t[3926] ^ n[3927];
assign t[3928] = t[3927] ^ n[3928];
assign t[3929] = t[3928] ^ n[3929];
assign t[3930] = t[3929] ^ n[3930];
assign t[3931] = t[3930] ^ n[3931];
assign t[3932] = t[3931] ^ n[3932];
assign t[3933] = t[3932] ^ n[3933];
assign t[3934] = t[3933] ^ n[3934];
assign t[3935] = t[3934] ^ n[3935];
assign t[3936] = t[3935] ^ n[3936];
assign t[3937] = t[3936] ^ n[3937];
assign t[3938] = t[3937] ^ n[3938];
assign t[3939] = t[3938] ^ n[3939];
assign t[3940] = t[3939] ^ n[3940];
assign t[3941] = t[3940] ^ n[3941];
assign t[3942] = t[3941] ^ n[3942];
assign t[3943] = t[3942] ^ n[3943];
assign t[3944] = t[3943] ^ n[3944];
assign t[3945] = t[3944] ^ n[3945];
assign t[3946] = t[3945] ^ n[3946];
assign t[3947] = t[3946] ^ n[3947];
assign t[3948] = t[3947] ^ n[3948];
assign t[3949] = t[3948] ^ n[3949];
assign t[3950] = t[3949] ^ n[3950];
assign t[3951] = t[3950] ^ n[3951];
assign t[3952] = t[3951] ^ n[3952];
assign t[3953] = t[3952] ^ n[3953];
assign t[3954] = t[3953] ^ n[3954];
assign t[3955] = t[3954] ^ n[3955];
assign t[3956] = t[3955] ^ n[3956];
assign t[3957] = t[3956] ^ n[3957];
assign t[3958] = t[3957] ^ n[3958];
assign t[3959] = t[3958] ^ n[3959];
assign t[3960] = t[3959] ^ n[3960];
assign t[3961] = t[3960] ^ n[3961];
assign t[3962] = t[3961] ^ n[3962];
assign t[3963] = t[3962] ^ n[3963];
assign t[3964] = t[3963] ^ n[3964];
assign t[3965] = t[3964] ^ n[3965];
assign t[3966] = t[3965] ^ n[3966];
assign t[3967] = t[3966] ^ n[3967];
assign t[3968] = t[3967] ^ n[3968];
assign t[3969] = t[3968] ^ n[3969];
assign t[3970] = t[3969] ^ n[3970];
assign t[3971] = t[3970] ^ n[3971];
assign t[3972] = t[3971] ^ n[3972];
assign t[3973] = t[3972] ^ n[3973];
assign t[3974] = t[3973] ^ n[3974];
assign t[3975] = t[3974] ^ n[3975];
assign t[3976] = t[3975] ^ n[3976];
assign t[3977] = t[3976] ^ n[3977];
assign t[3978] = t[3977] ^ n[3978];
assign t[3979] = t[3978] ^ n[3979];
assign t[3980] = t[3979] ^ n[3980];
assign t[3981] = t[3980] ^ n[3981];
assign t[3982] = t[3981] ^ n[3982];
assign t[3983] = t[3982] ^ n[3983];
assign t[3984] = t[3983] ^ n[3984];
assign t[3985] = t[3984] ^ n[3985];
assign t[3986] = t[3985] ^ n[3986];
assign t[3987] = t[3986] ^ n[3987];
assign t[3988] = t[3987] ^ n[3988];
assign t[3989] = t[3988] ^ n[3989];
assign t[3990] = t[3989] ^ n[3990];
assign t[3991] = t[3990] ^ n[3991];
assign t[3992] = t[3991] ^ n[3992];
assign t[3993] = t[3992] ^ n[3993];
assign t[3994] = t[3993] ^ n[3994];
assign t[3995] = t[3994] ^ n[3995];
assign t[3996] = t[3995] ^ n[3996];
assign t[3997] = t[3996] ^ n[3997];
assign t[3998] = t[3997] ^ n[3998];
assign t[3999] = t[3998] ^ n[3999];
assign t[4000] = t[3999] ^ n[4000];
assign t[4001] = t[4000] ^ n[4001];
assign t[4002] = t[4001] ^ n[4002];
assign t[4003] = t[4002] ^ n[4003];
assign t[4004] = t[4003] ^ n[4004];
assign t[4005] = t[4004] ^ n[4005];
assign t[4006] = t[4005] ^ n[4006];
assign t[4007] = t[4006] ^ n[4007];
assign t[4008] = t[4007] ^ n[4008];
assign t[4009] = t[4008] ^ n[4009];
assign t[4010] = t[4009] ^ n[4010];
assign t[4011] = t[4010] ^ n[4011];
assign t[4012] = t[4011] ^ n[4012];
assign t[4013] = t[4012] ^ n[4013];
assign t[4014] = t[4013] ^ n[4014];
assign t[4015] = t[4014] ^ n[4015];
assign t[4016] = t[4015] ^ n[4016];
assign t[4017] = t[4016] ^ n[4017];
assign t[4018] = t[4017] ^ n[4018];
assign t[4019] = t[4018] ^ n[4019];
assign t[4020] = t[4019] ^ n[4020];
assign t[4021] = t[4020] ^ n[4021];
assign t[4022] = t[4021] ^ n[4022];
assign t[4023] = t[4022] ^ n[4023];
assign t[4024] = t[4023] ^ n[4024];
assign t[4025] = t[4024] ^ n[4025];
assign t[4026] = t[4025] ^ n[4026];
assign t[4027] = t[4026] ^ n[4027];
assign t[4028] = t[4027] ^ n[4028];
assign t[4029] = t[4028] ^ n[4029];
assign t[4030] = t[4029] ^ n[4030];
assign t[4031] = t[4030] ^ n[4031];
assign t[4032] = t[4031] ^ n[4032];
assign t[4033] = t[4032] ^ n[4033];
assign t[4034] = t[4033] ^ n[4034];
assign t[4035] = t[4034] ^ n[4035];
assign t[4036] = t[4035] ^ n[4036];
assign t[4037] = t[4036] ^ n[4037];
assign t[4038] = t[4037] ^ n[4038];
assign t[4039] = t[4038] ^ n[4039];
assign t[4040] = t[4039] ^ n[4040];
assign t[4041] = t[4040] ^ n[4041];
assign t[4042] = t[4041] ^ n[4042];
assign t[4043] = t[4042] ^ n[4043];
assign t[4044] = t[4043] ^ n[4044];
assign t[4045] = t[4044] ^ n[4045];
assign t[4046] = t[4045] ^ n[4046];
assign t[4047] = t[4046] ^ n[4047];
assign t[4048] = t[4047] ^ n[4048];
assign t[4049] = t[4048] ^ n[4049];
assign t[4050] = t[4049] ^ n[4050];
assign t[4051] = t[4050] ^ n[4051];
assign t[4052] = t[4051] ^ n[4052];
assign t[4053] = t[4052] ^ n[4053];
assign t[4054] = t[4053] ^ n[4054];
assign t[4055] = t[4054] ^ n[4055];
assign t[4056] = t[4055] ^ n[4056];
assign t[4057] = t[4056] ^ n[4057];
assign t[4058] = t[4057] ^ n[4058];
assign t[4059] = t[4058] ^ n[4059];
assign t[4060] = t[4059] ^ n[4060];
assign t[4061] = t[4060] ^ n[4061];
assign t[4062] = t[4061] ^ n[4062];
assign t[4063] = t[4062] ^ n[4063];
assign t[4064] = t[4063] ^ n[4064];
assign t[4065] = t[4064] ^ n[4065];
assign t[4066] = t[4065] ^ n[4066];
assign t[4067] = t[4066] ^ n[4067];
assign t[4068] = t[4067] ^ n[4068];
assign t[4069] = t[4068] ^ n[4069];
assign t[4070] = t[4069] ^ n[4070];
assign t[4071] = t[4070] ^ n[4071];
assign t[4072] = t[4071] ^ n[4072];
assign t[4073] = t[4072] ^ n[4073];
assign t[4074] = t[4073] ^ n[4074];
assign t[4075] = t[4074] ^ n[4075];
assign t[4076] = t[4075] ^ n[4076];
assign t[4077] = t[4076] ^ n[4077];
assign t[4078] = t[4077] ^ n[4078];
assign t[4079] = t[4078] ^ n[4079];
assign t[4080] = t[4079] ^ n[4080];
assign t[4081] = t[4080] ^ n[4081];
assign t[4082] = t[4081] ^ n[4082];

//asigning bit 11
assign s[11] = ( a[11] ^ b [11] ) ^ t[4082];

assign t[4083] = n[4083];
assign t[4084] = t[4083] ^ n[4084];
assign t[4085] = t[4084] ^ n[4085];
assign t[4086] = t[4085] ^ n[4086];
assign t[4087] = t[4086] ^ n[4087];
assign t[4088] = t[4087] ^ n[4088];
assign t[4089] = t[4088] ^ n[4089];
assign t[4090] = t[4089] ^ n[4090];
assign t[4091] = t[4090] ^ n[4091];
assign t[4092] = t[4091] ^ n[4092];
assign t[4093] = t[4092] ^ n[4093];
assign t[4094] = t[4093] ^ n[4094];
assign t[4095] = t[4094] ^ n[4095];
assign t[4096] = t[4095] ^ n[4096];
assign t[4097] = t[4096] ^ n[4097];
assign t[4098] = t[4097] ^ n[4098];
assign t[4099] = t[4098] ^ n[4099];
assign t[4100] = t[4099] ^ n[4100];
assign t[4101] = t[4100] ^ n[4101];
assign t[4102] = t[4101] ^ n[4102];
assign t[4103] = t[4102] ^ n[4103];
assign t[4104] = t[4103] ^ n[4104];
assign t[4105] = t[4104] ^ n[4105];
assign t[4106] = t[4105] ^ n[4106];
assign t[4107] = t[4106] ^ n[4107];
assign t[4108] = t[4107] ^ n[4108];
assign t[4109] = t[4108] ^ n[4109];
assign t[4110] = t[4109] ^ n[4110];
assign t[4111] = t[4110] ^ n[4111];
assign t[4112] = t[4111] ^ n[4112];
assign t[4113] = t[4112] ^ n[4113];
assign t[4114] = t[4113] ^ n[4114];
assign t[4115] = t[4114] ^ n[4115];
assign t[4116] = t[4115] ^ n[4116];
assign t[4117] = t[4116] ^ n[4117];
assign t[4118] = t[4117] ^ n[4118];
assign t[4119] = t[4118] ^ n[4119];
assign t[4120] = t[4119] ^ n[4120];
assign t[4121] = t[4120] ^ n[4121];
assign t[4122] = t[4121] ^ n[4122];
assign t[4123] = t[4122] ^ n[4123];
assign t[4124] = t[4123] ^ n[4124];
assign t[4125] = t[4124] ^ n[4125];
assign t[4126] = t[4125] ^ n[4126];
assign t[4127] = t[4126] ^ n[4127];
assign t[4128] = t[4127] ^ n[4128];
assign t[4129] = t[4128] ^ n[4129];
assign t[4130] = t[4129] ^ n[4130];
assign t[4131] = t[4130] ^ n[4131];
assign t[4132] = t[4131] ^ n[4132];
assign t[4133] = t[4132] ^ n[4133];
assign t[4134] = t[4133] ^ n[4134];
assign t[4135] = t[4134] ^ n[4135];
assign t[4136] = t[4135] ^ n[4136];
assign t[4137] = t[4136] ^ n[4137];
assign t[4138] = t[4137] ^ n[4138];
assign t[4139] = t[4138] ^ n[4139];
assign t[4140] = t[4139] ^ n[4140];
assign t[4141] = t[4140] ^ n[4141];
assign t[4142] = t[4141] ^ n[4142];
assign t[4143] = t[4142] ^ n[4143];
assign t[4144] = t[4143] ^ n[4144];
assign t[4145] = t[4144] ^ n[4145];
assign t[4146] = t[4145] ^ n[4146];
assign t[4147] = t[4146] ^ n[4147];
assign t[4148] = t[4147] ^ n[4148];
assign t[4149] = t[4148] ^ n[4149];
assign t[4150] = t[4149] ^ n[4150];
assign t[4151] = t[4150] ^ n[4151];
assign t[4152] = t[4151] ^ n[4152];
assign t[4153] = t[4152] ^ n[4153];
assign t[4154] = t[4153] ^ n[4154];
assign t[4155] = t[4154] ^ n[4155];
assign t[4156] = t[4155] ^ n[4156];
assign t[4157] = t[4156] ^ n[4157];
assign t[4158] = t[4157] ^ n[4158];
assign t[4159] = t[4158] ^ n[4159];
assign t[4160] = t[4159] ^ n[4160];
assign t[4161] = t[4160] ^ n[4161];
assign t[4162] = t[4161] ^ n[4162];
assign t[4163] = t[4162] ^ n[4163];
assign t[4164] = t[4163] ^ n[4164];
assign t[4165] = t[4164] ^ n[4165];
assign t[4166] = t[4165] ^ n[4166];
assign t[4167] = t[4166] ^ n[4167];
assign t[4168] = t[4167] ^ n[4168];
assign t[4169] = t[4168] ^ n[4169];
assign t[4170] = t[4169] ^ n[4170];
assign t[4171] = t[4170] ^ n[4171];
assign t[4172] = t[4171] ^ n[4172];
assign t[4173] = t[4172] ^ n[4173];
assign t[4174] = t[4173] ^ n[4174];
assign t[4175] = t[4174] ^ n[4175];
assign t[4176] = t[4175] ^ n[4176];
assign t[4177] = t[4176] ^ n[4177];
assign t[4178] = t[4177] ^ n[4178];
assign t[4179] = t[4178] ^ n[4179];
assign t[4180] = t[4179] ^ n[4180];
assign t[4181] = t[4180] ^ n[4181];
assign t[4182] = t[4181] ^ n[4182];
assign t[4183] = t[4182] ^ n[4183];
assign t[4184] = t[4183] ^ n[4184];
assign t[4185] = t[4184] ^ n[4185];
assign t[4186] = t[4185] ^ n[4186];
assign t[4187] = t[4186] ^ n[4187];
assign t[4188] = t[4187] ^ n[4188];
assign t[4189] = t[4188] ^ n[4189];
assign t[4190] = t[4189] ^ n[4190];
assign t[4191] = t[4190] ^ n[4191];
assign t[4192] = t[4191] ^ n[4192];
assign t[4193] = t[4192] ^ n[4193];
assign t[4194] = t[4193] ^ n[4194];
assign t[4195] = t[4194] ^ n[4195];
assign t[4196] = t[4195] ^ n[4196];
assign t[4197] = t[4196] ^ n[4197];
assign t[4198] = t[4197] ^ n[4198];
assign t[4199] = t[4198] ^ n[4199];
assign t[4200] = t[4199] ^ n[4200];
assign t[4201] = t[4200] ^ n[4201];
assign t[4202] = t[4201] ^ n[4202];
assign t[4203] = t[4202] ^ n[4203];
assign t[4204] = t[4203] ^ n[4204];
assign t[4205] = t[4204] ^ n[4205];
assign t[4206] = t[4205] ^ n[4206];
assign t[4207] = t[4206] ^ n[4207];
assign t[4208] = t[4207] ^ n[4208];
assign t[4209] = t[4208] ^ n[4209];
assign t[4210] = t[4209] ^ n[4210];
assign t[4211] = t[4210] ^ n[4211];
assign t[4212] = t[4211] ^ n[4212];
assign t[4213] = t[4212] ^ n[4213];
assign t[4214] = t[4213] ^ n[4214];
assign t[4215] = t[4214] ^ n[4215];
assign t[4216] = t[4215] ^ n[4216];
assign t[4217] = t[4216] ^ n[4217];
assign t[4218] = t[4217] ^ n[4218];
assign t[4219] = t[4218] ^ n[4219];
assign t[4220] = t[4219] ^ n[4220];
assign t[4221] = t[4220] ^ n[4221];
assign t[4222] = t[4221] ^ n[4222];
assign t[4223] = t[4222] ^ n[4223];
assign t[4224] = t[4223] ^ n[4224];
assign t[4225] = t[4224] ^ n[4225];
assign t[4226] = t[4225] ^ n[4226];
assign t[4227] = t[4226] ^ n[4227];
assign t[4228] = t[4227] ^ n[4228];
assign t[4229] = t[4228] ^ n[4229];
assign t[4230] = t[4229] ^ n[4230];
assign t[4231] = t[4230] ^ n[4231];
assign t[4232] = t[4231] ^ n[4232];
assign t[4233] = t[4232] ^ n[4233];
assign t[4234] = t[4233] ^ n[4234];
assign t[4235] = t[4234] ^ n[4235];
assign t[4236] = t[4235] ^ n[4236];
assign t[4237] = t[4236] ^ n[4237];
assign t[4238] = t[4237] ^ n[4238];
assign t[4239] = t[4238] ^ n[4239];
assign t[4240] = t[4239] ^ n[4240];
assign t[4241] = t[4240] ^ n[4241];
assign t[4242] = t[4241] ^ n[4242];
assign t[4243] = t[4242] ^ n[4243];
assign t[4244] = t[4243] ^ n[4244];
assign t[4245] = t[4244] ^ n[4245];
assign t[4246] = t[4245] ^ n[4246];
assign t[4247] = t[4246] ^ n[4247];
assign t[4248] = t[4247] ^ n[4248];
assign t[4249] = t[4248] ^ n[4249];
assign t[4250] = t[4249] ^ n[4250];
assign t[4251] = t[4250] ^ n[4251];
assign t[4252] = t[4251] ^ n[4252];
assign t[4253] = t[4252] ^ n[4253];
assign t[4254] = t[4253] ^ n[4254];
assign t[4255] = t[4254] ^ n[4255];
assign t[4256] = t[4255] ^ n[4256];
assign t[4257] = t[4256] ^ n[4257];
assign t[4258] = t[4257] ^ n[4258];
assign t[4259] = t[4258] ^ n[4259];
assign t[4260] = t[4259] ^ n[4260];
assign t[4261] = t[4260] ^ n[4261];
assign t[4262] = t[4261] ^ n[4262];
assign t[4263] = t[4262] ^ n[4263];
assign t[4264] = t[4263] ^ n[4264];
assign t[4265] = t[4264] ^ n[4265];
assign t[4266] = t[4265] ^ n[4266];
assign t[4267] = t[4266] ^ n[4267];
assign t[4268] = t[4267] ^ n[4268];
assign t[4269] = t[4268] ^ n[4269];
assign t[4270] = t[4269] ^ n[4270];
assign t[4271] = t[4270] ^ n[4271];
assign t[4272] = t[4271] ^ n[4272];
assign t[4273] = t[4272] ^ n[4273];
assign t[4274] = t[4273] ^ n[4274];
assign t[4275] = t[4274] ^ n[4275];
assign t[4276] = t[4275] ^ n[4276];
assign t[4277] = t[4276] ^ n[4277];
assign t[4278] = t[4277] ^ n[4278];
assign t[4279] = t[4278] ^ n[4279];
assign t[4280] = t[4279] ^ n[4280];
assign t[4281] = t[4280] ^ n[4281];
assign t[4282] = t[4281] ^ n[4282];
assign t[4283] = t[4282] ^ n[4283];
assign t[4284] = t[4283] ^ n[4284];
assign t[4285] = t[4284] ^ n[4285];
assign t[4286] = t[4285] ^ n[4286];
assign t[4287] = t[4286] ^ n[4287];
assign t[4288] = t[4287] ^ n[4288];
assign t[4289] = t[4288] ^ n[4289];
assign t[4290] = t[4289] ^ n[4290];
assign t[4291] = t[4290] ^ n[4291];
assign t[4292] = t[4291] ^ n[4292];
assign t[4293] = t[4292] ^ n[4293];
assign t[4294] = t[4293] ^ n[4294];
assign t[4295] = t[4294] ^ n[4295];
assign t[4296] = t[4295] ^ n[4296];
assign t[4297] = t[4296] ^ n[4297];
assign t[4298] = t[4297] ^ n[4298];
assign t[4299] = t[4298] ^ n[4299];
assign t[4300] = t[4299] ^ n[4300];
assign t[4301] = t[4300] ^ n[4301];
assign t[4302] = t[4301] ^ n[4302];
assign t[4303] = t[4302] ^ n[4303];
assign t[4304] = t[4303] ^ n[4304];
assign t[4305] = t[4304] ^ n[4305];
assign t[4306] = t[4305] ^ n[4306];
assign t[4307] = t[4306] ^ n[4307];
assign t[4308] = t[4307] ^ n[4308];
assign t[4309] = t[4308] ^ n[4309];
assign t[4310] = t[4309] ^ n[4310];
assign t[4311] = t[4310] ^ n[4311];
assign t[4312] = t[4311] ^ n[4312];
assign t[4313] = t[4312] ^ n[4313];
assign t[4314] = t[4313] ^ n[4314];
assign t[4315] = t[4314] ^ n[4315];
assign t[4316] = t[4315] ^ n[4316];
assign t[4317] = t[4316] ^ n[4317];
assign t[4318] = t[4317] ^ n[4318];
assign t[4319] = t[4318] ^ n[4319];
assign t[4320] = t[4319] ^ n[4320];
assign t[4321] = t[4320] ^ n[4321];
assign t[4322] = t[4321] ^ n[4322];
assign t[4323] = t[4322] ^ n[4323];
assign t[4324] = t[4323] ^ n[4324];
assign t[4325] = t[4324] ^ n[4325];
assign t[4326] = t[4325] ^ n[4326];
assign t[4327] = t[4326] ^ n[4327];
assign t[4328] = t[4327] ^ n[4328];
assign t[4329] = t[4328] ^ n[4329];
assign t[4330] = t[4329] ^ n[4330];
assign t[4331] = t[4330] ^ n[4331];
assign t[4332] = t[4331] ^ n[4332];
assign t[4333] = t[4332] ^ n[4333];
assign t[4334] = t[4333] ^ n[4334];
assign t[4335] = t[4334] ^ n[4335];
assign t[4336] = t[4335] ^ n[4336];
assign t[4337] = t[4336] ^ n[4337];
assign t[4338] = t[4337] ^ n[4338];
assign t[4339] = t[4338] ^ n[4339];
assign t[4340] = t[4339] ^ n[4340];
assign t[4341] = t[4340] ^ n[4341];
assign t[4342] = t[4341] ^ n[4342];
assign t[4343] = t[4342] ^ n[4343];
assign t[4344] = t[4343] ^ n[4344];
assign t[4345] = t[4344] ^ n[4345];
assign t[4346] = t[4345] ^ n[4346];
assign t[4347] = t[4346] ^ n[4347];
assign t[4348] = t[4347] ^ n[4348];
assign t[4349] = t[4348] ^ n[4349];
assign t[4350] = t[4349] ^ n[4350];
assign t[4351] = t[4350] ^ n[4351];
assign t[4352] = t[4351] ^ n[4352];
assign t[4353] = t[4352] ^ n[4353];
assign t[4354] = t[4353] ^ n[4354];
assign t[4355] = t[4354] ^ n[4355];
assign t[4356] = t[4355] ^ n[4356];
assign t[4357] = t[4356] ^ n[4357];
assign t[4358] = t[4357] ^ n[4358];
assign t[4359] = t[4358] ^ n[4359];
assign t[4360] = t[4359] ^ n[4360];
assign t[4361] = t[4360] ^ n[4361];
assign t[4362] = t[4361] ^ n[4362];
assign t[4363] = t[4362] ^ n[4363];
assign t[4364] = t[4363] ^ n[4364];
assign t[4365] = t[4364] ^ n[4365];
assign t[4366] = t[4365] ^ n[4366];
assign t[4367] = t[4366] ^ n[4367];
assign t[4368] = t[4367] ^ n[4368];
assign t[4369] = t[4368] ^ n[4369];
assign t[4370] = t[4369] ^ n[4370];
assign t[4371] = t[4370] ^ n[4371];
assign t[4372] = t[4371] ^ n[4372];
assign t[4373] = t[4372] ^ n[4373];
assign t[4374] = t[4373] ^ n[4374];
assign t[4375] = t[4374] ^ n[4375];
assign t[4376] = t[4375] ^ n[4376];
assign t[4377] = t[4376] ^ n[4377];
assign t[4378] = t[4377] ^ n[4378];
assign t[4379] = t[4378] ^ n[4379];
assign t[4380] = t[4379] ^ n[4380];
assign t[4381] = t[4380] ^ n[4381];
assign t[4382] = t[4381] ^ n[4382];
assign t[4383] = t[4382] ^ n[4383];
assign t[4384] = t[4383] ^ n[4384];
assign t[4385] = t[4384] ^ n[4385];
assign t[4386] = t[4385] ^ n[4386];
assign t[4387] = t[4386] ^ n[4387];
assign t[4388] = t[4387] ^ n[4388];
assign t[4389] = t[4388] ^ n[4389];
assign t[4390] = t[4389] ^ n[4390];
assign t[4391] = t[4390] ^ n[4391];
assign t[4392] = t[4391] ^ n[4392];
assign t[4393] = t[4392] ^ n[4393];
assign t[4394] = t[4393] ^ n[4394];
assign t[4395] = t[4394] ^ n[4395];
assign t[4396] = t[4395] ^ n[4396];
assign t[4397] = t[4396] ^ n[4397];
assign t[4398] = t[4397] ^ n[4398];
assign t[4399] = t[4398] ^ n[4399];
assign t[4400] = t[4399] ^ n[4400];
assign t[4401] = t[4400] ^ n[4401];
assign t[4402] = t[4401] ^ n[4402];
assign t[4403] = t[4402] ^ n[4403];
assign t[4404] = t[4403] ^ n[4404];
assign t[4405] = t[4404] ^ n[4405];
assign t[4406] = t[4405] ^ n[4406];
assign t[4407] = t[4406] ^ n[4407];
assign t[4408] = t[4407] ^ n[4408];
assign t[4409] = t[4408] ^ n[4409];
assign t[4410] = t[4409] ^ n[4410];
assign t[4411] = t[4410] ^ n[4411];
assign t[4412] = t[4411] ^ n[4412];
assign t[4413] = t[4412] ^ n[4413];
assign t[4414] = t[4413] ^ n[4414];
assign t[4415] = t[4414] ^ n[4415];
assign t[4416] = t[4415] ^ n[4416];
assign t[4417] = t[4416] ^ n[4417];
assign t[4418] = t[4417] ^ n[4418];
assign t[4419] = t[4418] ^ n[4419];
assign t[4420] = t[4419] ^ n[4420];
assign t[4421] = t[4420] ^ n[4421];
assign t[4422] = t[4421] ^ n[4422];
assign t[4423] = t[4422] ^ n[4423];
assign t[4424] = t[4423] ^ n[4424];
assign t[4425] = t[4424] ^ n[4425];
assign t[4426] = t[4425] ^ n[4426];
assign t[4427] = t[4426] ^ n[4427];
assign t[4428] = t[4427] ^ n[4428];
assign t[4429] = t[4428] ^ n[4429];
assign t[4430] = t[4429] ^ n[4430];
assign t[4431] = t[4430] ^ n[4431];
assign t[4432] = t[4431] ^ n[4432];
assign t[4433] = t[4432] ^ n[4433];
assign t[4434] = t[4433] ^ n[4434];
assign t[4435] = t[4434] ^ n[4435];
assign t[4436] = t[4435] ^ n[4436];
assign t[4437] = t[4436] ^ n[4437];
assign t[4438] = t[4437] ^ n[4438];
assign t[4439] = t[4438] ^ n[4439];
assign t[4440] = t[4439] ^ n[4440];
assign t[4441] = t[4440] ^ n[4441];
assign t[4442] = t[4441] ^ n[4442];
assign t[4443] = t[4442] ^ n[4443];
assign t[4444] = t[4443] ^ n[4444];
assign t[4445] = t[4444] ^ n[4445];
assign t[4446] = t[4445] ^ n[4446];
assign t[4447] = t[4446] ^ n[4447];
assign t[4448] = t[4447] ^ n[4448];
assign t[4449] = t[4448] ^ n[4449];
assign t[4450] = t[4449] ^ n[4450];
assign t[4451] = t[4450] ^ n[4451];
assign t[4452] = t[4451] ^ n[4452];
assign t[4453] = t[4452] ^ n[4453];
assign t[4454] = t[4453] ^ n[4454];
assign t[4455] = t[4454] ^ n[4455];
assign t[4456] = t[4455] ^ n[4456];
assign t[4457] = t[4456] ^ n[4457];
assign t[4458] = t[4457] ^ n[4458];
assign t[4459] = t[4458] ^ n[4459];
assign t[4460] = t[4459] ^ n[4460];
assign t[4461] = t[4460] ^ n[4461];
assign t[4462] = t[4461] ^ n[4462];
assign t[4463] = t[4462] ^ n[4463];
assign t[4464] = t[4463] ^ n[4464];
assign t[4465] = t[4464] ^ n[4465];
assign t[4466] = t[4465] ^ n[4466];
assign t[4467] = t[4466] ^ n[4467];
assign t[4468] = t[4467] ^ n[4468];
assign t[4469] = t[4468] ^ n[4469];
assign t[4470] = t[4469] ^ n[4470];
assign t[4471] = t[4470] ^ n[4471];
assign t[4472] = t[4471] ^ n[4472];
assign t[4473] = t[4472] ^ n[4473];
assign t[4474] = t[4473] ^ n[4474];
assign t[4475] = t[4474] ^ n[4475];
assign t[4476] = t[4475] ^ n[4476];
assign t[4477] = t[4476] ^ n[4477];
assign t[4478] = t[4477] ^ n[4478];
assign t[4479] = t[4478] ^ n[4479];
assign t[4480] = t[4479] ^ n[4480];
assign t[4481] = t[4480] ^ n[4481];
assign t[4482] = t[4481] ^ n[4482];
assign t[4483] = t[4482] ^ n[4483];
assign t[4484] = t[4483] ^ n[4484];
assign t[4485] = t[4484] ^ n[4485];
assign t[4486] = t[4485] ^ n[4486];
assign t[4487] = t[4486] ^ n[4487];
assign t[4488] = t[4487] ^ n[4488];
assign t[4489] = t[4488] ^ n[4489];
assign t[4490] = t[4489] ^ n[4490];
assign t[4491] = t[4490] ^ n[4491];
assign t[4492] = t[4491] ^ n[4492];
assign t[4493] = t[4492] ^ n[4493];
assign t[4494] = t[4493] ^ n[4494];
assign t[4495] = t[4494] ^ n[4495];
assign t[4496] = t[4495] ^ n[4496];
assign t[4497] = t[4496] ^ n[4497];
assign t[4498] = t[4497] ^ n[4498];
assign t[4499] = t[4498] ^ n[4499];
assign t[4500] = t[4499] ^ n[4500];
assign t[4501] = t[4500] ^ n[4501];
assign t[4502] = t[4501] ^ n[4502];
assign t[4503] = t[4502] ^ n[4503];
assign t[4504] = t[4503] ^ n[4504];
assign t[4505] = t[4504] ^ n[4505];
assign t[4506] = t[4505] ^ n[4506];
assign t[4507] = t[4506] ^ n[4507];
assign t[4508] = t[4507] ^ n[4508];
assign t[4509] = t[4508] ^ n[4509];
assign t[4510] = t[4509] ^ n[4510];
assign t[4511] = t[4510] ^ n[4511];
assign t[4512] = t[4511] ^ n[4512];
assign t[4513] = t[4512] ^ n[4513];
assign t[4514] = t[4513] ^ n[4514];
assign t[4515] = t[4514] ^ n[4515];
assign t[4516] = t[4515] ^ n[4516];
assign t[4517] = t[4516] ^ n[4517];
assign t[4518] = t[4517] ^ n[4518];
assign t[4519] = t[4518] ^ n[4519];
assign t[4520] = t[4519] ^ n[4520];
assign t[4521] = t[4520] ^ n[4521];
assign t[4522] = t[4521] ^ n[4522];
assign t[4523] = t[4522] ^ n[4523];
assign t[4524] = t[4523] ^ n[4524];
assign t[4525] = t[4524] ^ n[4525];
assign t[4526] = t[4525] ^ n[4526];
assign t[4527] = t[4526] ^ n[4527];
assign t[4528] = t[4527] ^ n[4528];
assign t[4529] = t[4528] ^ n[4529];
assign t[4530] = t[4529] ^ n[4530];
assign t[4531] = t[4530] ^ n[4531];
assign t[4532] = t[4531] ^ n[4532];
assign t[4533] = t[4532] ^ n[4533];
assign t[4534] = t[4533] ^ n[4534];
assign t[4535] = t[4534] ^ n[4535];
assign t[4536] = t[4535] ^ n[4536];
assign t[4537] = t[4536] ^ n[4537];
assign t[4538] = t[4537] ^ n[4538];
assign t[4539] = t[4538] ^ n[4539];
assign t[4540] = t[4539] ^ n[4540];
assign t[4541] = t[4540] ^ n[4541];
assign t[4542] = t[4541] ^ n[4542];
assign t[4543] = t[4542] ^ n[4543];
assign t[4544] = t[4543] ^ n[4544];
assign t[4545] = t[4544] ^ n[4545];
assign t[4546] = t[4545] ^ n[4546];
assign t[4547] = t[4546] ^ n[4547];
assign t[4548] = t[4547] ^ n[4548];
assign t[4549] = t[4548] ^ n[4549];
assign t[4550] = t[4549] ^ n[4550];
assign t[4551] = t[4550] ^ n[4551];
assign t[4552] = t[4551] ^ n[4552];
assign t[4553] = t[4552] ^ n[4553];
assign t[4554] = t[4553] ^ n[4554];
assign t[4555] = t[4554] ^ n[4555];
assign t[4556] = t[4555] ^ n[4556];
assign t[4557] = t[4556] ^ n[4557];
assign t[4558] = t[4557] ^ n[4558];
assign t[4559] = t[4558] ^ n[4559];
assign t[4560] = t[4559] ^ n[4560];
assign t[4561] = t[4560] ^ n[4561];
assign t[4562] = t[4561] ^ n[4562];
assign t[4563] = t[4562] ^ n[4563];
assign t[4564] = t[4563] ^ n[4564];
assign t[4565] = t[4564] ^ n[4565];
assign t[4566] = t[4565] ^ n[4566];
assign t[4567] = t[4566] ^ n[4567];
assign t[4568] = t[4567] ^ n[4568];
assign t[4569] = t[4568] ^ n[4569];
assign t[4570] = t[4569] ^ n[4570];
assign t[4571] = t[4570] ^ n[4571];
assign t[4572] = t[4571] ^ n[4572];
assign t[4573] = t[4572] ^ n[4573];
assign t[4574] = t[4573] ^ n[4574];
assign t[4575] = t[4574] ^ n[4575];
assign t[4576] = t[4575] ^ n[4576];
assign t[4577] = t[4576] ^ n[4577];
assign t[4578] = t[4577] ^ n[4578];
assign t[4579] = t[4578] ^ n[4579];
assign t[4580] = t[4579] ^ n[4580];
assign t[4581] = t[4580] ^ n[4581];
assign t[4582] = t[4581] ^ n[4582];
assign t[4583] = t[4582] ^ n[4583];
assign t[4584] = t[4583] ^ n[4584];
assign t[4585] = t[4584] ^ n[4585];
assign t[4586] = t[4585] ^ n[4586];
assign t[4587] = t[4586] ^ n[4587];
assign t[4588] = t[4587] ^ n[4588];
assign t[4589] = t[4588] ^ n[4589];
assign t[4590] = t[4589] ^ n[4590];
assign t[4591] = t[4590] ^ n[4591];
assign t[4592] = t[4591] ^ n[4592];
assign t[4593] = t[4592] ^ n[4593];
assign t[4594] = t[4593] ^ n[4594];
assign t[4595] = t[4594] ^ n[4595];
assign t[4596] = t[4595] ^ n[4596];
assign t[4597] = t[4596] ^ n[4597];
assign t[4598] = t[4597] ^ n[4598];
assign t[4599] = t[4598] ^ n[4599];
assign t[4600] = t[4599] ^ n[4600];
assign t[4601] = t[4600] ^ n[4601];
assign t[4602] = t[4601] ^ n[4602];
assign t[4603] = t[4602] ^ n[4603];
assign t[4604] = t[4603] ^ n[4604];
assign t[4605] = t[4604] ^ n[4605];
assign t[4606] = t[4605] ^ n[4606];
assign t[4607] = t[4606] ^ n[4607];
assign t[4608] = t[4607] ^ n[4608];
assign t[4609] = t[4608] ^ n[4609];
assign t[4610] = t[4609] ^ n[4610];
assign t[4611] = t[4610] ^ n[4611];
assign t[4612] = t[4611] ^ n[4612];
assign t[4613] = t[4612] ^ n[4613];
assign t[4614] = t[4613] ^ n[4614];
assign t[4615] = t[4614] ^ n[4615];
assign t[4616] = t[4615] ^ n[4616];
assign t[4617] = t[4616] ^ n[4617];
assign t[4618] = t[4617] ^ n[4618];
assign t[4619] = t[4618] ^ n[4619];
assign t[4620] = t[4619] ^ n[4620];
assign t[4621] = t[4620] ^ n[4621];
assign t[4622] = t[4621] ^ n[4622];
assign t[4623] = t[4622] ^ n[4623];
assign t[4624] = t[4623] ^ n[4624];
assign t[4625] = t[4624] ^ n[4625];
assign t[4626] = t[4625] ^ n[4626];
assign t[4627] = t[4626] ^ n[4627];
assign t[4628] = t[4627] ^ n[4628];
assign t[4629] = t[4628] ^ n[4629];
assign t[4630] = t[4629] ^ n[4630];
assign t[4631] = t[4630] ^ n[4631];
assign t[4632] = t[4631] ^ n[4632];
assign t[4633] = t[4632] ^ n[4633];
assign t[4634] = t[4633] ^ n[4634];
assign t[4635] = t[4634] ^ n[4635];
assign t[4636] = t[4635] ^ n[4636];
assign t[4637] = t[4636] ^ n[4637];
assign t[4638] = t[4637] ^ n[4638];
assign t[4639] = t[4638] ^ n[4639];
assign t[4640] = t[4639] ^ n[4640];
assign t[4641] = t[4640] ^ n[4641];
assign t[4642] = t[4641] ^ n[4642];
assign t[4643] = t[4642] ^ n[4643];
assign t[4644] = t[4643] ^ n[4644];
assign t[4645] = t[4644] ^ n[4645];
assign t[4646] = t[4645] ^ n[4646];
assign t[4647] = t[4646] ^ n[4647];
assign t[4648] = t[4647] ^ n[4648];
assign t[4649] = t[4648] ^ n[4649];
assign t[4650] = t[4649] ^ n[4650];
assign t[4651] = t[4650] ^ n[4651];
assign t[4652] = t[4651] ^ n[4652];
assign t[4653] = t[4652] ^ n[4653];
assign t[4654] = t[4653] ^ n[4654];
assign t[4655] = t[4654] ^ n[4655];
assign t[4656] = t[4655] ^ n[4656];
assign t[4657] = t[4656] ^ n[4657];
assign t[4658] = t[4657] ^ n[4658];
assign t[4659] = t[4658] ^ n[4659];
assign t[4660] = t[4659] ^ n[4660];
assign t[4661] = t[4660] ^ n[4661];
assign t[4662] = t[4661] ^ n[4662];
assign t[4663] = t[4662] ^ n[4663];
assign t[4664] = t[4663] ^ n[4664];
assign t[4665] = t[4664] ^ n[4665];
assign t[4666] = t[4665] ^ n[4666];
assign t[4667] = t[4666] ^ n[4667];
assign t[4668] = t[4667] ^ n[4668];
assign t[4669] = t[4668] ^ n[4669];
assign t[4670] = t[4669] ^ n[4670];
assign t[4671] = t[4670] ^ n[4671];
assign t[4672] = t[4671] ^ n[4672];
assign t[4673] = t[4672] ^ n[4673];
assign t[4674] = t[4673] ^ n[4674];
assign t[4675] = t[4674] ^ n[4675];
assign t[4676] = t[4675] ^ n[4676];
assign t[4677] = t[4676] ^ n[4677];
assign t[4678] = t[4677] ^ n[4678];
assign t[4679] = t[4678] ^ n[4679];
assign t[4680] = t[4679] ^ n[4680];
assign t[4681] = t[4680] ^ n[4681];
assign t[4682] = t[4681] ^ n[4682];
assign t[4683] = t[4682] ^ n[4683];
assign t[4684] = t[4683] ^ n[4684];
assign t[4685] = t[4684] ^ n[4685];
assign t[4686] = t[4685] ^ n[4686];
assign t[4687] = t[4686] ^ n[4687];
assign t[4688] = t[4687] ^ n[4688];
assign t[4689] = t[4688] ^ n[4689];
assign t[4690] = t[4689] ^ n[4690];
assign t[4691] = t[4690] ^ n[4691];
assign t[4692] = t[4691] ^ n[4692];
assign t[4693] = t[4692] ^ n[4693];
assign t[4694] = t[4693] ^ n[4694];
assign t[4695] = t[4694] ^ n[4695];
assign t[4696] = t[4695] ^ n[4696];
assign t[4697] = t[4696] ^ n[4697];
assign t[4698] = t[4697] ^ n[4698];
assign t[4699] = t[4698] ^ n[4699];
assign t[4700] = t[4699] ^ n[4700];
assign t[4701] = t[4700] ^ n[4701];
assign t[4702] = t[4701] ^ n[4702];
assign t[4703] = t[4702] ^ n[4703];
assign t[4704] = t[4703] ^ n[4704];
assign t[4705] = t[4704] ^ n[4705];
assign t[4706] = t[4705] ^ n[4706];
assign t[4707] = t[4706] ^ n[4707];
assign t[4708] = t[4707] ^ n[4708];
assign t[4709] = t[4708] ^ n[4709];
assign t[4710] = t[4709] ^ n[4710];
assign t[4711] = t[4710] ^ n[4711];
assign t[4712] = t[4711] ^ n[4712];
assign t[4713] = t[4712] ^ n[4713];
assign t[4714] = t[4713] ^ n[4714];
assign t[4715] = t[4714] ^ n[4715];
assign t[4716] = t[4715] ^ n[4716];
assign t[4717] = t[4716] ^ n[4717];
assign t[4718] = t[4717] ^ n[4718];
assign t[4719] = t[4718] ^ n[4719];
assign t[4720] = t[4719] ^ n[4720];
assign t[4721] = t[4720] ^ n[4721];
assign t[4722] = t[4721] ^ n[4722];
assign t[4723] = t[4722] ^ n[4723];
assign t[4724] = t[4723] ^ n[4724];
assign t[4725] = t[4724] ^ n[4725];
assign t[4726] = t[4725] ^ n[4726];
assign t[4727] = t[4726] ^ n[4727];
assign t[4728] = t[4727] ^ n[4728];
assign t[4729] = t[4728] ^ n[4729];
assign t[4730] = t[4729] ^ n[4730];
assign t[4731] = t[4730] ^ n[4731];
assign t[4732] = t[4731] ^ n[4732];
assign t[4733] = t[4732] ^ n[4733];
assign t[4734] = t[4733] ^ n[4734];
assign t[4735] = t[4734] ^ n[4735];
assign t[4736] = t[4735] ^ n[4736];
assign t[4737] = t[4736] ^ n[4737];
assign t[4738] = t[4737] ^ n[4738];
assign t[4739] = t[4738] ^ n[4739];
assign t[4740] = t[4739] ^ n[4740];
assign t[4741] = t[4740] ^ n[4741];
assign t[4742] = t[4741] ^ n[4742];
assign t[4743] = t[4742] ^ n[4743];
assign t[4744] = t[4743] ^ n[4744];
assign t[4745] = t[4744] ^ n[4745];
assign t[4746] = t[4745] ^ n[4746];
assign t[4747] = t[4746] ^ n[4747];
assign t[4748] = t[4747] ^ n[4748];
assign t[4749] = t[4748] ^ n[4749];
assign t[4750] = t[4749] ^ n[4750];
assign t[4751] = t[4750] ^ n[4751];
assign t[4752] = t[4751] ^ n[4752];
assign t[4753] = t[4752] ^ n[4753];
assign t[4754] = t[4753] ^ n[4754];
assign t[4755] = t[4754] ^ n[4755];
assign t[4756] = t[4755] ^ n[4756];
assign t[4757] = t[4756] ^ n[4757];
assign t[4758] = t[4757] ^ n[4758];
assign t[4759] = t[4758] ^ n[4759];
assign t[4760] = t[4759] ^ n[4760];
assign t[4761] = t[4760] ^ n[4761];
assign t[4762] = t[4761] ^ n[4762];
assign t[4763] = t[4762] ^ n[4763];
assign t[4764] = t[4763] ^ n[4764];
assign t[4765] = t[4764] ^ n[4765];
assign t[4766] = t[4765] ^ n[4766];
assign t[4767] = t[4766] ^ n[4767];
assign t[4768] = t[4767] ^ n[4768];
assign t[4769] = t[4768] ^ n[4769];
assign t[4770] = t[4769] ^ n[4770];
assign t[4771] = t[4770] ^ n[4771];
assign t[4772] = t[4771] ^ n[4772];
assign t[4773] = t[4772] ^ n[4773];
assign t[4774] = t[4773] ^ n[4774];
assign t[4775] = t[4774] ^ n[4775];
assign t[4776] = t[4775] ^ n[4776];
assign t[4777] = t[4776] ^ n[4777];
assign t[4778] = t[4777] ^ n[4778];
assign t[4779] = t[4778] ^ n[4779];
assign t[4780] = t[4779] ^ n[4780];
assign t[4781] = t[4780] ^ n[4781];
assign t[4782] = t[4781] ^ n[4782];
assign t[4783] = t[4782] ^ n[4783];
assign t[4784] = t[4783] ^ n[4784];
assign t[4785] = t[4784] ^ n[4785];
assign t[4786] = t[4785] ^ n[4786];
assign t[4787] = t[4786] ^ n[4787];
assign t[4788] = t[4787] ^ n[4788];
assign t[4789] = t[4788] ^ n[4789];
assign t[4790] = t[4789] ^ n[4790];
assign t[4791] = t[4790] ^ n[4791];
assign t[4792] = t[4791] ^ n[4792];
assign t[4793] = t[4792] ^ n[4793];
assign t[4794] = t[4793] ^ n[4794];
assign t[4795] = t[4794] ^ n[4795];
assign t[4796] = t[4795] ^ n[4796];
assign t[4797] = t[4796] ^ n[4797];
assign t[4798] = t[4797] ^ n[4798];
assign t[4799] = t[4798] ^ n[4799];
assign t[4800] = t[4799] ^ n[4800];
assign t[4801] = t[4800] ^ n[4801];
assign t[4802] = t[4801] ^ n[4802];
assign t[4803] = t[4802] ^ n[4803];
assign t[4804] = t[4803] ^ n[4804];
assign t[4805] = t[4804] ^ n[4805];
assign t[4806] = t[4805] ^ n[4806];
assign t[4807] = t[4806] ^ n[4807];
assign t[4808] = t[4807] ^ n[4808];
assign t[4809] = t[4808] ^ n[4809];
assign t[4810] = t[4809] ^ n[4810];
assign t[4811] = t[4810] ^ n[4811];
assign t[4812] = t[4811] ^ n[4812];
assign t[4813] = t[4812] ^ n[4813];
assign t[4814] = t[4813] ^ n[4814];
assign t[4815] = t[4814] ^ n[4815];
assign t[4816] = t[4815] ^ n[4816];
assign t[4817] = t[4816] ^ n[4817];
assign t[4818] = t[4817] ^ n[4818];
assign t[4819] = t[4818] ^ n[4819];
assign t[4820] = t[4819] ^ n[4820];
assign t[4821] = t[4820] ^ n[4821];
assign t[4822] = t[4821] ^ n[4822];
assign t[4823] = t[4822] ^ n[4823];
assign t[4824] = t[4823] ^ n[4824];
assign t[4825] = t[4824] ^ n[4825];
assign t[4826] = t[4825] ^ n[4826];
assign t[4827] = t[4826] ^ n[4827];
assign t[4828] = t[4827] ^ n[4828];
assign t[4829] = t[4828] ^ n[4829];
assign t[4830] = t[4829] ^ n[4830];
assign t[4831] = t[4830] ^ n[4831];
assign t[4832] = t[4831] ^ n[4832];
assign t[4833] = t[4832] ^ n[4833];
assign t[4834] = t[4833] ^ n[4834];
assign t[4835] = t[4834] ^ n[4835];
assign t[4836] = t[4835] ^ n[4836];
assign t[4837] = t[4836] ^ n[4837];
assign t[4838] = t[4837] ^ n[4838];
assign t[4839] = t[4838] ^ n[4839];
assign t[4840] = t[4839] ^ n[4840];
assign t[4841] = t[4840] ^ n[4841];
assign t[4842] = t[4841] ^ n[4842];
assign t[4843] = t[4842] ^ n[4843];
assign t[4844] = t[4843] ^ n[4844];
assign t[4845] = t[4844] ^ n[4845];
assign t[4846] = t[4845] ^ n[4846];
assign t[4847] = t[4846] ^ n[4847];
assign t[4848] = t[4847] ^ n[4848];
assign t[4849] = t[4848] ^ n[4849];
assign t[4850] = t[4849] ^ n[4850];
assign t[4851] = t[4850] ^ n[4851];
assign t[4852] = t[4851] ^ n[4852];
assign t[4853] = t[4852] ^ n[4853];
assign t[4854] = t[4853] ^ n[4854];
assign t[4855] = t[4854] ^ n[4855];
assign t[4856] = t[4855] ^ n[4856];
assign t[4857] = t[4856] ^ n[4857];
assign t[4858] = t[4857] ^ n[4858];
assign t[4859] = t[4858] ^ n[4859];
assign t[4860] = t[4859] ^ n[4860];
assign t[4861] = t[4860] ^ n[4861];
assign t[4862] = t[4861] ^ n[4862];
assign t[4863] = t[4862] ^ n[4863];
assign t[4864] = t[4863] ^ n[4864];
assign t[4865] = t[4864] ^ n[4865];
assign t[4866] = t[4865] ^ n[4866];
assign t[4867] = t[4866] ^ n[4867];
assign t[4868] = t[4867] ^ n[4868];
assign t[4869] = t[4868] ^ n[4869];
assign t[4870] = t[4869] ^ n[4870];
assign t[4871] = t[4870] ^ n[4871];
assign t[4872] = t[4871] ^ n[4872];
assign t[4873] = t[4872] ^ n[4873];
assign t[4874] = t[4873] ^ n[4874];
assign t[4875] = t[4874] ^ n[4875];
assign t[4876] = t[4875] ^ n[4876];
assign t[4877] = t[4876] ^ n[4877];
assign t[4878] = t[4877] ^ n[4878];
assign t[4879] = t[4878] ^ n[4879];
assign t[4880] = t[4879] ^ n[4880];
assign t[4881] = t[4880] ^ n[4881];
assign t[4882] = t[4881] ^ n[4882];
assign t[4883] = t[4882] ^ n[4883];
assign t[4884] = t[4883] ^ n[4884];
assign t[4885] = t[4884] ^ n[4885];
assign t[4886] = t[4885] ^ n[4886];
assign t[4887] = t[4886] ^ n[4887];
assign t[4888] = t[4887] ^ n[4888];
assign t[4889] = t[4888] ^ n[4889];
assign t[4890] = t[4889] ^ n[4890];
assign t[4891] = t[4890] ^ n[4891];
assign t[4892] = t[4891] ^ n[4892];
assign t[4893] = t[4892] ^ n[4893];
assign t[4894] = t[4893] ^ n[4894];
assign t[4895] = t[4894] ^ n[4895];
assign t[4896] = t[4895] ^ n[4896];
assign t[4897] = t[4896] ^ n[4897];
assign t[4898] = t[4897] ^ n[4898];
assign t[4899] = t[4898] ^ n[4899];
assign t[4900] = t[4899] ^ n[4900];
assign t[4901] = t[4900] ^ n[4901];
assign t[4902] = t[4901] ^ n[4902];
assign t[4903] = t[4902] ^ n[4903];
assign t[4904] = t[4903] ^ n[4904];
assign t[4905] = t[4904] ^ n[4905];
assign t[4906] = t[4905] ^ n[4906];
assign t[4907] = t[4906] ^ n[4907];
assign t[4908] = t[4907] ^ n[4908];
assign t[4909] = t[4908] ^ n[4909];
assign t[4910] = t[4909] ^ n[4910];
assign t[4911] = t[4910] ^ n[4911];
assign t[4912] = t[4911] ^ n[4912];
assign t[4913] = t[4912] ^ n[4913];
assign t[4914] = t[4913] ^ n[4914];
assign t[4915] = t[4914] ^ n[4915];
assign t[4916] = t[4915] ^ n[4916];
assign t[4917] = t[4916] ^ n[4917];
assign t[4918] = t[4917] ^ n[4918];
assign t[4919] = t[4918] ^ n[4919];
assign t[4920] = t[4919] ^ n[4920];
assign t[4921] = t[4920] ^ n[4921];
assign t[4922] = t[4921] ^ n[4922];
assign t[4923] = t[4922] ^ n[4923];
assign t[4924] = t[4923] ^ n[4924];
assign t[4925] = t[4924] ^ n[4925];
assign t[4926] = t[4925] ^ n[4926];
assign t[4927] = t[4926] ^ n[4927];
assign t[4928] = t[4927] ^ n[4928];
assign t[4929] = t[4928] ^ n[4929];
assign t[4930] = t[4929] ^ n[4930];
assign t[4931] = t[4930] ^ n[4931];
assign t[4932] = t[4931] ^ n[4932];
assign t[4933] = t[4932] ^ n[4933];
assign t[4934] = t[4933] ^ n[4934];
assign t[4935] = t[4934] ^ n[4935];
assign t[4936] = t[4935] ^ n[4936];
assign t[4937] = t[4936] ^ n[4937];
assign t[4938] = t[4937] ^ n[4938];
assign t[4939] = t[4938] ^ n[4939];
assign t[4940] = t[4939] ^ n[4940];
assign t[4941] = t[4940] ^ n[4941];
assign t[4942] = t[4941] ^ n[4942];
assign t[4943] = t[4942] ^ n[4943];
assign t[4944] = t[4943] ^ n[4944];
assign t[4945] = t[4944] ^ n[4945];
assign t[4946] = t[4945] ^ n[4946];
assign t[4947] = t[4946] ^ n[4947];
assign t[4948] = t[4947] ^ n[4948];
assign t[4949] = t[4948] ^ n[4949];
assign t[4950] = t[4949] ^ n[4950];
assign t[4951] = t[4950] ^ n[4951];
assign t[4952] = t[4951] ^ n[4952];
assign t[4953] = t[4952] ^ n[4953];
assign t[4954] = t[4953] ^ n[4954];
assign t[4955] = t[4954] ^ n[4955];
assign t[4956] = t[4955] ^ n[4956];
assign t[4957] = t[4956] ^ n[4957];
assign t[4958] = t[4957] ^ n[4958];
assign t[4959] = t[4958] ^ n[4959];
assign t[4960] = t[4959] ^ n[4960];
assign t[4961] = t[4960] ^ n[4961];
assign t[4962] = t[4961] ^ n[4962];
assign t[4963] = t[4962] ^ n[4963];
assign t[4964] = t[4963] ^ n[4964];
assign t[4965] = t[4964] ^ n[4965];
assign t[4966] = t[4965] ^ n[4966];
assign t[4967] = t[4966] ^ n[4967];
assign t[4968] = t[4967] ^ n[4968];
assign t[4969] = t[4968] ^ n[4969];
assign t[4970] = t[4969] ^ n[4970];
assign t[4971] = t[4970] ^ n[4971];
assign t[4972] = t[4971] ^ n[4972];
assign t[4973] = t[4972] ^ n[4973];
assign t[4974] = t[4973] ^ n[4974];
assign t[4975] = t[4974] ^ n[4975];
assign t[4976] = t[4975] ^ n[4976];
assign t[4977] = t[4976] ^ n[4977];
assign t[4978] = t[4977] ^ n[4978];
assign t[4979] = t[4978] ^ n[4979];
assign t[4980] = t[4979] ^ n[4980];
assign t[4981] = t[4980] ^ n[4981];
assign t[4982] = t[4981] ^ n[4982];
assign t[4983] = t[4982] ^ n[4983];
assign t[4984] = t[4983] ^ n[4984];
assign t[4985] = t[4984] ^ n[4985];
assign t[4986] = t[4985] ^ n[4986];
assign t[4987] = t[4986] ^ n[4987];
assign t[4988] = t[4987] ^ n[4988];
assign t[4989] = t[4988] ^ n[4989];
assign t[4990] = t[4989] ^ n[4990];
assign t[4991] = t[4990] ^ n[4991];
assign t[4992] = t[4991] ^ n[4992];
assign t[4993] = t[4992] ^ n[4993];
assign t[4994] = t[4993] ^ n[4994];
assign t[4995] = t[4994] ^ n[4995];
assign t[4996] = t[4995] ^ n[4996];
assign t[4997] = t[4996] ^ n[4997];
assign t[4998] = t[4997] ^ n[4998];
assign t[4999] = t[4998] ^ n[4999];
assign t[5000] = t[4999] ^ n[5000];
assign t[5001] = t[5000] ^ n[5001];
assign t[5002] = t[5001] ^ n[5002];
assign t[5003] = t[5002] ^ n[5003];
assign t[5004] = t[5003] ^ n[5004];
assign t[5005] = t[5004] ^ n[5005];
assign t[5006] = t[5005] ^ n[5006];
assign t[5007] = t[5006] ^ n[5007];
assign t[5008] = t[5007] ^ n[5008];
assign t[5009] = t[5008] ^ n[5009];
assign t[5010] = t[5009] ^ n[5010];
assign t[5011] = t[5010] ^ n[5011];
assign t[5012] = t[5011] ^ n[5012];
assign t[5013] = t[5012] ^ n[5013];
assign t[5014] = t[5013] ^ n[5014];
assign t[5015] = t[5014] ^ n[5015];
assign t[5016] = t[5015] ^ n[5016];
assign t[5017] = t[5016] ^ n[5017];
assign t[5018] = t[5017] ^ n[5018];
assign t[5019] = t[5018] ^ n[5019];
assign t[5020] = t[5019] ^ n[5020];
assign t[5021] = t[5020] ^ n[5021];
assign t[5022] = t[5021] ^ n[5022];
assign t[5023] = t[5022] ^ n[5023];
assign t[5024] = t[5023] ^ n[5024];
assign t[5025] = t[5024] ^ n[5025];
assign t[5026] = t[5025] ^ n[5026];
assign t[5027] = t[5026] ^ n[5027];
assign t[5028] = t[5027] ^ n[5028];
assign t[5029] = t[5028] ^ n[5029];
assign t[5030] = t[5029] ^ n[5030];
assign t[5031] = t[5030] ^ n[5031];
assign t[5032] = t[5031] ^ n[5032];
assign t[5033] = t[5032] ^ n[5033];
assign t[5034] = t[5033] ^ n[5034];
assign t[5035] = t[5034] ^ n[5035];
assign t[5036] = t[5035] ^ n[5036];
assign t[5037] = t[5036] ^ n[5037];
assign t[5038] = t[5037] ^ n[5038];
assign t[5039] = t[5038] ^ n[5039];
assign t[5040] = t[5039] ^ n[5040];
assign t[5041] = t[5040] ^ n[5041];
assign t[5042] = t[5041] ^ n[5042];
assign t[5043] = t[5042] ^ n[5043];
assign t[5044] = t[5043] ^ n[5044];
assign t[5045] = t[5044] ^ n[5045];
assign t[5046] = t[5045] ^ n[5046];
assign t[5047] = t[5046] ^ n[5047];
assign t[5048] = t[5047] ^ n[5048];
assign t[5049] = t[5048] ^ n[5049];
assign t[5050] = t[5049] ^ n[5050];
assign t[5051] = t[5050] ^ n[5051];
assign t[5052] = t[5051] ^ n[5052];
assign t[5053] = t[5052] ^ n[5053];
assign t[5054] = t[5053] ^ n[5054];
assign t[5055] = t[5054] ^ n[5055];
assign t[5056] = t[5055] ^ n[5056];
assign t[5057] = t[5056] ^ n[5057];
assign t[5058] = t[5057] ^ n[5058];
assign t[5059] = t[5058] ^ n[5059];
assign t[5060] = t[5059] ^ n[5060];
assign t[5061] = t[5060] ^ n[5061];
assign t[5062] = t[5061] ^ n[5062];
assign t[5063] = t[5062] ^ n[5063];
assign t[5064] = t[5063] ^ n[5064];
assign t[5065] = t[5064] ^ n[5065];
assign t[5066] = t[5065] ^ n[5066];
assign t[5067] = t[5066] ^ n[5067];
assign t[5068] = t[5067] ^ n[5068];
assign t[5069] = t[5068] ^ n[5069];
assign t[5070] = t[5069] ^ n[5070];
assign t[5071] = t[5070] ^ n[5071];
assign t[5072] = t[5071] ^ n[5072];
assign t[5073] = t[5072] ^ n[5073];
assign t[5074] = t[5073] ^ n[5074];
assign t[5075] = t[5074] ^ n[5075];
assign t[5076] = t[5075] ^ n[5076];
assign t[5077] = t[5076] ^ n[5077];
assign t[5078] = t[5077] ^ n[5078];
assign t[5079] = t[5078] ^ n[5079];
assign t[5080] = t[5079] ^ n[5080];
assign t[5081] = t[5080] ^ n[5081];
assign t[5082] = t[5081] ^ n[5082];
assign t[5083] = t[5082] ^ n[5083];
assign t[5084] = t[5083] ^ n[5084];
assign t[5085] = t[5084] ^ n[5085];
assign t[5086] = t[5085] ^ n[5086];
assign t[5087] = t[5086] ^ n[5087];
assign t[5088] = t[5087] ^ n[5088];
assign t[5089] = t[5088] ^ n[5089];
assign t[5090] = t[5089] ^ n[5090];
assign t[5091] = t[5090] ^ n[5091];
assign t[5092] = t[5091] ^ n[5092];
assign t[5093] = t[5092] ^ n[5093];
assign t[5094] = t[5093] ^ n[5094];
assign t[5095] = t[5094] ^ n[5095];
assign t[5096] = t[5095] ^ n[5096];
assign t[5097] = t[5096] ^ n[5097];
assign t[5098] = t[5097] ^ n[5098];
assign t[5099] = t[5098] ^ n[5099];
assign t[5100] = t[5099] ^ n[5100];
assign t[5101] = t[5100] ^ n[5101];
assign t[5102] = t[5101] ^ n[5102];
assign t[5103] = t[5102] ^ n[5103];
assign t[5104] = t[5103] ^ n[5104];
assign t[5105] = t[5104] ^ n[5105];
assign t[5106] = t[5105] ^ n[5106];
assign t[5107] = t[5106] ^ n[5107];
assign t[5108] = t[5107] ^ n[5108];
assign t[5109] = t[5108] ^ n[5109];
assign t[5110] = t[5109] ^ n[5110];
assign t[5111] = t[5110] ^ n[5111];
assign t[5112] = t[5111] ^ n[5112];
assign t[5113] = t[5112] ^ n[5113];
assign t[5114] = t[5113] ^ n[5114];
assign t[5115] = t[5114] ^ n[5115];
assign t[5116] = t[5115] ^ n[5116];
assign t[5117] = t[5116] ^ n[5117];
assign t[5118] = t[5117] ^ n[5118];
assign t[5119] = t[5118] ^ n[5119];
assign t[5120] = t[5119] ^ n[5120];
assign t[5121] = t[5120] ^ n[5121];
assign t[5122] = t[5121] ^ n[5122];
assign t[5123] = t[5122] ^ n[5123];
assign t[5124] = t[5123] ^ n[5124];
assign t[5125] = t[5124] ^ n[5125];
assign t[5126] = t[5125] ^ n[5126];
assign t[5127] = t[5126] ^ n[5127];
assign t[5128] = t[5127] ^ n[5128];
assign t[5129] = t[5128] ^ n[5129];
assign t[5130] = t[5129] ^ n[5130];
assign t[5131] = t[5130] ^ n[5131];
assign t[5132] = t[5131] ^ n[5132];
assign t[5133] = t[5132] ^ n[5133];
assign t[5134] = t[5133] ^ n[5134];
assign t[5135] = t[5134] ^ n[5135];
assign t[5136] = t[5135] ^ n[5136];
assign t[5137] = t[5136] ^ n[5137];
assign t[5138] = t[5137] ^ n[5138];
assign t[5139] = t[5138] ^ n[5139];
assign t[5140] = t[5139] ^ n[5140];
assign t[5141] = t[5140] ^ n[5141];
assign t[5142] = t[5141] ^ n[5142];
assign t[5143] = t[5142] ^ n[5143];
assign t[5144] = t[5143] ^ n[5144];
assign t[5145] = t[5144] ^ n[5145];
assign t[5146] = t[5145] ^ n[5146];
assign t[5147] = t[5146] ^ n[5147];
assign t[5148] = t[5147] ^ n[5148];
assign t[5149] = t[5148] ^ n[5149];
assign t[5150] = t[5149] ^ n[5150];
assign t[5151] = t[5150] ^ n[5151];
assign t[5152] = t[5151] ^ n[5152];
assign t[5153] = t[5152] ^ n[5153];
assign t[5154] = t[5153] ^ n[5154];
assign t[5155] = t[5154] ^ n[5155];
assign t[5156] = t[5155] ^ n[5156];
assign t[5157] = t[5156] ^ n[5157];
assign t[5158] = t[5157] ^ n[5158];
assign t[5159] = t[5158] ^ n[5159];
assign t[5160] = t[5159] ^ n[5160];
assign t[5161] = t[5160] ^ n[5161];
assign t[5162] = t[5161] ^ n[5162];
assign t[5163] = t[5162] ^ n[5163];
assign t[5164] = t[5163] ^ n[5164];
assign t[5165] = t[5164] ^ n[5165];
assign t[5166] = t[5165] ^ n[5166];
assign t[5167] = t[5166] ^ n[5167];
assign t[5168] = t[5167] ^ n[5168];
assign t[5169] = t[5168] ^ n[5169];
assign t[5170] = t[5169] ^ n[5170];
assign t[5171] = t[5170] ^ n[5171];
assign t[5172] = t[5171] ^ n[5172];
assign t[5173] = t[5172] ^ n[5173];
assign t[5174] = t[5173] ^ n[5174];
assign t[5175] = t[5174] ^ n[5175];
assign t[5176] = t[5175] ^ n[5176];
assign t[5177] = t[5176] ^ n[5177];
assign t[5178] = t[5177] ^ n[5178];
assign t[5179] = t[5178] ^ n[5179];
assign t[5180] = t[5179] ^ n[5180];
assign t[5181] = t[5180] ^ n[5181];
assign t[5182] = t[5181] ^ n[5182];
assign t[5183] = t[5182] ^ n[5183];
assign t[5184] = t[5183] ^ n[5184];
assign t[5185] = t[5184] ^ n[5185];
assign t[5186] = t[5185] ^ n[5186];
assign t[5187] = t[5186] ^ n[5187];
assign t[5188] = t[5187] ^ n[5188];
assign t[5189] = t[5188] ^ n[5189];
assign t[5190] = t[5189] ^ n[5190];
assign t[5191] = t[5190] ^ n[5191];
assign t[5192] = t[5191] ^ n[5192];
assign t[5193] = t[5192] ^ n[5193];
assign t[5194] = t[5193] ^ n[5194];
assign t[5195] = t[5194] ^ n[5195];
assign t[5196] = t[5195] ^ n[5196];
assign t[5197] = t[5196] ^ n[5197];
assign t[5198] = t[5197] ^ n[5198];
assign t[5199] = t[5198] ^ n[5199];
assign t[5200] = t[5199] ^ n[5200];
assign t[5201] = t[5200] ^ n[5201];
assign t[5202] = t[5201] ^ n[5202];
assign t[5203] = t[5202] ^ n[5203];
assign t[5204] = t[5203] ^ n[5204];
assign t[5205] = t[5204] ^ n[5205];
assign t[5206] = t[5205] ^ n[5206];
assign t[5207] = t[5206] ^ n[5207];
assign t[5208] = t[5207] ^ n[5208];
assign t[5209] = t[5208] ^ n[5209];
assign t[5210] = t[5209] ^ n[5210];
assign t[5211] = t[5210] ^ n[5211];
assign t[5212] = t[5211] ^ n[5212];
assign t[5213] = t[5212] ^ n[5213];
assign t[5214] = t[5213] ^ n[5214];
assign t[5215] = t[5214] ^ n[5215];
assign t[5216] = t[5215] ^ n[5216];
assign t[5217] = t[5216] ^ n[5217];
assign t[5218] = t[5217] ^ n[5218];
assign t[5219] = t[5218] ^ n[5219];
assign t[5220] = t[5219] ^ n[5220];
assign t[5221] = t[5220] ^ n[5221];
assign t[5222] = t[5221] ^ n[5222];
assign t[5223] = t[5222] ^ n[5223];
assign t[5224] = t[5223] ^ n[5224];
assign t[5225] = t[5224] ^ n[5225];
assign t[5226] = t[5225] ^ n[5226];
assign t[5227] = t[5226] ^ n[5227];
assign t[5228] = t[5227] ^ n[5228];
assign t[5229] = t[5228] ^ n[5229];
assign t[5230] = t[5229] ^ n[5230];
assign t[5231] = t[5230] ^ n[5231];
assign t[5232] = t[5231] ^ n[5232];
assign t[5233] = t[5232] ^ n[5233];
assign t[5234] = t[5233] ^ n[5234];
assign t[5235] = t[5234] ^ n[5235];
assign t[5236] = t[5235] ^ n[5236];
assign t[5237] = t[5236] ^ n[5237];
assign t[5238] = t[5237] ^ n[5238];
assign t[5239] = t[5238] ^ n[5239];
assign t[5240] = t[5239] ^ n[5240];
assign t[5241] = t[5240] ^ n[5241];
assign t[5242] = t[5241] ^ n[5242];
assign t[5243] = t[5242] ^ n[5243];
assign t[5244] = t[5243] ^ n[5244];
assign t[5245] = t[5244] ^ n[5245];
assign t[5246] = t[5245] ^ n[5246];
assign t[5247] = t[5246] ^ n[5247];
assign t[5248] = t[5247] ^ n[5248];
assign t[5249] = t[5248] ^ n[5249];
assign t[5250] = t[5249] ^ n[5250];
assign t[5251] = t[5250] ^ n[5251];
assign t[5252] = t[5251] ^ n[5252];
assign t[5253] = t[5252] ^ n[5253];
assign t[5254] = t[5253] ^ n[5254];
assign t[5255] = t[5254] ^ n[5255];
assign t[5256] = t[5255] ^ n[5256];
assign t[5257] = t[5256] ^ n[5257];
assign t[5258] = t[5257] ^ n[5258];
assign t[5259] = t[5258] ^ n[5259];
assign t[5260] = t[5259] ^ n[5260];
assign t[5261] = t[5260] ^ n[5261];
assign t[5262] = t[5261] ^ n[5262];
assign t[5263] = t[5262] ^ n[5263];
assign t[5264] = t[5263] ^ n[5264];
assign t[5265] = t[5264] ^ n[5265];
assign t[5266] = t[5265] ^ n[5266];
assign t[5267] = t[5266] ^ n[5267];
assign t[5268] = t[5267] ^ n[5268];
assign t[5269] = t[5268] ^ n[5269];
assign t[5270] = t[5269] ^ n[5270];
assign t[5271] = t[5270] ^ n[5271];
assign t[5272] = t[5271] ^ n[5272];
assign t[5273] = t[5272] ^ n[5273];
assign t[5274] = t[5273] ^ n[5274];
assign t[5275] = t[5274] ^ n[5275];
assign t[5276] = t[5275] ^ n[5276];
assign t[5277] = t[5276] ^ n[5277];
assign t[5278] = t[5277] ^ n[5278];
assign t[5279] = t[5278] ^ n[5279];
assign t[5280] = t[5279] ^ n[5280];
assign t[5281] = t[5280] ^ n[5281];
assign t[5282] = t[5281] ^ n[5282];
assign t[5283] = t[5282] ^ n[5283];
assign t[5284] = t[5283] ^ n[5284];
assign t[5285] = t[5284] ^ n[5285];
assign t[5286] = t[5285] ^ n[5286];
assign t[5287] = t[5286] ^ n[5287];
assign t[5288] = t[5287] ^ n[5288];
assign t[5289] = t[5288] ^ n[5289];
assign t[5290] = t[5289] ^ n[5290];
assign t[5291] = t[5290] ^ n[5291];
assign t[5292] = t[5291] ^ n[5292];
assign t[5293] = t[5292] ^ n[5293];
assign t[5294] = t[5293] ^ n[5294];
assign t[5295] = t[5294] ^ n[5295];
assign t[5296] = t[5295] ^ n[5296];
assign t[5297] = t[5296] ^ n[5297];
assign t[5298] = t[5297] ^ n[5298];
assign t[5299] = t[5298] ^ n[5299];
assign t[5300] = t[5299] ^ n[5300];
assign t[5301] = t[5300] ^ n[5301];
assign t[5302] = t[5301] ^ n[5302];
assign t[5303] = t[5302] ^ n[5303];
assign t[5304] = t[5303] ^ n[5304];
assign t[5305] = t[5304] ^ n[5305];
assign t[5306] = t[5305] ^ n[5306];
assign t[5307] = t[5306] ^ n[5307];
assign t[5308] = t[5307] ^ n[5308];
assign t[5309] = t[5308] ^ n[5309];
assign t[5310] = t[5309] ^ n[5310];
assign t[5311] = t[5310] ^ n[5311];
assign t[5312] = t[5311] ^ n[5312];
assign t[5313] = t[5312] ^ n[5313];
assign t[5314] = t[5313] ^ n[5314];
assign t[5315] = t[5314] ^ n[5315];
assign t[5316] = t[5315] ^ n[5316];
assign t[5317] = t[5316] ^ n[5317];
assign t[5318] = t[5317] ^ n[5318];
assign t[5319] = t[5318] ^ n[5319];
assign t[5320] = t[5319] ^ n[5320];
assign t[5321] = t[5320] ^ n[5321];
assign t[5322] = t[5321] ^ n[5322];
assign t[5323] = t[5322] ^ n[5323];
assign t[5324] = t[5323] ^ n[5324];
assign t[5325] = t[5324] ^ n[5325];
assign t[5326] = t[5325] ^ n[5326];
assign t[5327] = t[5326] ^ n[5327];
assign t[5328] = t[5327] ^ n[5328];
assign t[5329] = t[5328] ^ n[5329];
assign t[5330] = t[5329] ^ n[5330];
assign t[5331] = t[5330] ^ n[5331];
assign t[5332] = t[5331] ^ n[5332];
assign t[5333] = t[5332] ^ n[5333];
assign t[5334] = t[5333] ^ n[5334];
assign t[5335] = t[5334] ^ n[5335];
assign t[5336] = t[5335] ^ n[5336];
assign t[5337] = t[5336] ^ n[5337];
assign t[5338] = t[5337] ^ n[5338];
assign t[5339] = t[5338] ^ n[5339];
assign t[5340] = t[5339] ^ n[5340];
assign t[5341] = t[5340] ^ n[5341];
assign t[5342] = t[5341] ^ n[5342];
assign t[5343] = t[5342] ^ n[5343];
assign t[5344] = t[5343] ^ n[5344];
assign t[5345] = t[5344] ^ n[5345];
assign t[5346] = t[5345] ^ n[5346];
assign t[5347] = t[5346] ^ n[5347];
assign t[5348] = t[5347] ^ n[5348];
assign t[5349] = t[5348] ^ n[5349];
assign t[5350] = t[5349] ^ n[5350];
assign t[5351] = t[5350] ^ n[5351];
assign t[5352] = t[5351] ^ n[5352];
assign t[5353] = t[5352] ^ n[5353];
assign t[5354] = t[5353] ^ n[5354];
assign t[5355] = t[5354] ^ n[5355];
assign t[5356] = t[5355] ^ n[5356];
assign t[5357] = t[5356] ^ n[5357];
assign t[5358] = t[5357] ^ n[5358];
assign t[5359] = t[5358] ^ n[5359];
assign t[5360] = t[5359] ^ n[5360];
assign t[5361] = t[5360] ^ n[5361];
assign t[5362] = t[5361] ^ n[5362];
assign t[5363] = t[5362] ^ n[5363];
assign t[5364] = t[5363] ^ n[5364];
assign t[5365] = t[5364] ^ n[5365];
assign t[5366] = t[5365] ^ n[5366];
assign t[5367] = t[5366] ^ n[5367];
assign t[5368] = t[5367] ^ n[5368];
assign t[5369] = t[5368] ^ n[5369];
assign t[5370] = t[5369] ^ n[5370];
assign t[5371] = t[5370] ^ n[5371];
assign t[5372] = t[5371] ^ n[5372];
assign t[5373] = t[5372] ^ n[5373];
assign t[5374] = t[5373] ^ n[5374];
assign t[5375] = t[5374] ^ n[5375];
assign t[5376] = t[5375] ^ n[5376];
assign t[5377] = t[5376] ^ n[5377];
assign t[5378] = t[5377] ^ n[5378];
assign t[5379] = t[5378] ^ n[5379];
assign t[5380] = t[5379] ^ n[5380];
assign t[5381] = t[5380] ^ n[5381];
assign t[5382] = t[5381] ^ n[5382];
assign t[5383] = t[5382] ^ n[5383];
assign t[5384] = t[5383] ^ n[5384];
assign t[5385] = t[5384] ^ n[5385];
assign t[5386] = t[5385] ^ n[5386];
assign t[5387] = t[5386] ^ n[5387];
assign t[5388] = t[5387] ^ n[5388];
assign t[5389] = t[5388] ^ n[5389];
assign t[5390] = t[5389] ^ n[5390];
assign t[5391] = t[5390] ^ n[5391];
assign t[5392] = t[5391] ^ n[5392];
assign t[5393] = t[5392] ^ n[5393];
assign t[5394] = t[5393] ^ n[5394];
assign t[5395] = t[5394] ^ n[5395];
assign t[5396] = t[5395] ^ n[5396];
assign t[5397] = t[5396] ^ n[5397];
assign t[5398] = t[5397] ^ n[5398];
assign t[5399] = t[5398] ^ n[5399];
assign t[5400] = t[5399] ^ n[5400];
assign t[5401] = t[5400] ^ n[5401];
assign t[5402] = t[5401] ^ n[5402];
assign t[5403] = t[5402] ^ n[5403];
assign t[5404] = t[5403] ^ n[5404];
assign t[5405] = t[5404] ^ n[5405];
assign t[5406] = t[5405] ^ n[5406];
assign t[5407] = t[5406] ^ n[5407];
assign t[5408] = t[5407] ^ n[5408];
assign t[5409] = t[5408] ^ n[5409];
assign t[5410] = t[5409] ^ n[5410];
assign t[5411] = t[5410] ^ n[5411];
assign t[5412] = t[5411] ^ n[5412];
assign t[5413] = t[5412] ^ n[5413];
assign t[5414] = t[5413] ^ n[5414];
assign t[5415] = t[5414] ^ n[5415];
assign t[5416] = t[5415] ^ n[5416];
assign t[5417] = t[5416] ^ n[5417];
assign t[5418] = t[5417] ^ n[5418];
assign t[5419] = t[5418] ^ n[5419];
assign t[5420] = t[5419] ^ n[5420];
assign t[5421] = t[5420] ^ n[5421];
assign t[5422] = t[5421] ^ n[5422];
assign t[5423] = t[5422] ^ n[5423];
assign t[5424] = t[5423] ^ n[5424];
assign t[5425] = t[5424] ^ n[5425];
assign t[5426] = t[5425] ^ n[5426];
assign t[5427] = t[5426] ^ n[5427];
assign t[5428] = t[5427] ^ n[5428];
assign t[5429] = t[5428] ^ n[5429];
assign t[5430] = t[5429] ^ n[5430];
assign t[5431] = t[5430] ^ n[5431];
assign t[5432] = t[5431] ^ n[5432];
assign t[5433] = t[5432] ^ n[5433];
assign t[5434] = t[5433] ^ n[5434];
assign t[5435] = t[5434] ^ n[5435];
assign t[5436] = t[5435] ^ n[5436];
assign t[5437] = t[5436] ^ n[5437];
assign t[5438] = t[5437] ^ n[5438];
assign t[5439] = t[5438] ^ n[5439];
assign t[5440] = t[5439] ^ n[5440];
assign t[5441] = t[5440] ^ n[5441];
assign t[5442] = t[5441] ^ n[5442];
assign t[5443] = t[5442] ^ n[5443];
assign t[5444] = t[5443] ^ n[5444];
assign t[5445] = t[5444] ^ n[5445];
assign t[5446] = t[5445] ^ n[5446];
assign t[5447] = t[5446] ^ n[5447];
assign t[5448] = t[5447] ^ n[5448];
assign t[5449] = t[5448] ^ n[5449];
assign t[5450] = t[5449] ^ n[5450];
assign t[5451] = t[5450] ^ n[5451];
assign t[5452] = t[5451] ^ n[5452];
assign t[5453] = t[5452] ^ n[5453];
assign t[5454] = t[5453] ^ n[5454];
assign t[5455] = t[5454] ^ n[5455];
assign t[5456] = t[5455] ^ n[5456];
assign t[5457] = t[5456] ^ n[5457];
assign t[5458] = t[5457] ^ n[5458];
assign t[5459] = t[5458] ^ n[5459];
assign t[5460] = t[5459] ^ n[5460];
assign t[5461] = t[5460] ^ n[5461];
assign t[5462] = t[5461] ^ n[5462];
assign t[5463] = t[5462] ^ n[5463];
assign t[5464] = t[5463] ^ n[5464];
assign t[5465] = t[5464] ^ n[5465];
assign t[5466] = t[5465] ^ n[5466];
assign t[5467] = t[5466] ^ n[5467];
assign t[5468] = t[5467] ^ n[5468];
assign t[5469] = t[5468] ^ n[5469];
assign t[5470] = t[5469] ^ n[5470];
assign t[5471] = t[5470] ^ n[5471];
assign t[5472] = t[5471] ^ n[5472];
assign t[5473] = t[5472] ^ n[5473];
assign t[5474] = t[5473] ^ n[5474];
assign t[5475] = t[5474] ^ n[5475];
assign t[5476] = t[5475] ^ n[5476];
assign t[5477] = t[5476] ^ n[5477];
assign t[5478] = t[5477] ^ n[5478];
assign t[5479] = t[5478] ^ n[5479];
assign t[5480] = t[5479] ^ n[5480];
assign t[5481] = t[5480] ^ n[5481];
assign t[5482] = t[5481] ^ n[5482];
assign t[5483] = t[5482] ^ n[5483];
assign t[5484] = t[5483] ^ n[5484];
assign t[5485] = t[5484] ^ n[5485];
assign t[5486] = t[5485] ^ n[5486];
assign t[5487] = t[5486] ^ n[5487];
assign t[5488] = t[5487] ^ n[5488];
assign t[5489] = t[5488] ^ n[5489];
assign t[5490] = t[5489] ^ n[5490];
assign t[5491] = t[5490] ^ n[5491];
assign t[5492] = t[5491] ^ n[5492];
assign t[5493] = t[5492] ^ n[5493];
assign t[5494] = t[5493] ^ n[5494];
assign t[5495] = t[5494] ^ n[5495];
assign t[5496] = t[5495] ^ n[5496];
assign t[5497] = t[5496] ^ n[5497];
assign t[5498] = t[5497] ^ n[5498];
assign t[5499] = t[5498] ^ n[5499];
assign t[5500] = t[5499] ^ n[5500];
assign t[5501] = t[5500] ^ n[5501];
assign t[5502] = t[5501] ^ n[5502];
assign t[5503] = t[5502] ^ n[5503];
assign t[5504] = t[5503] ^ n[5504];
assign t[5505] = t[5504] ^ n[5505];
assign t[5506] = t[5505] ^ n[5506];
assign t[5507] = t[5506] ^ n[5507];
assign t[5508] = t[5507] ^ n[5508];
assign t[5509] = t[5508] ^ n[5509];
assign t[5510] = t[5509] ^ n[5510];
assign t[5511] = t[5510] ^ n[5511];
assign t[5512] = t[5511] ^ n[5512];
assign t[5513] = t[5512] ^ n[5513];
assign t[5514] = t[5513] ^ n[5514];
assign t[5515] = t[5514] ^ n[5515];
assign t[5516] = t[5515] ^ n[5516];
assign t[5517] = t[5516] ^ n[5517];
assign t[5518] = t[5517] ^ n[5518];
assign t[5519] = t[5518] ^ n[5519];
assign t[5520] = t[5519] ^ n[5520];
assign t[5521] = t[5520] ^ n[5521];
assign t[5522] = t[5521] ^ n[5522];
assign t[5523] = t[5522] ^ n[5523];
assign t[5524] = t[5523] ^ n[5524];
assign t[5525] = t[5524] ^ n[5525];
assign t[5526] = t[5525] ^ n[5526];
assign t[5527] = t[5526] ^ n[5527];
assign t[5528] = t[5527] ^ n[5528];
assign t[5529] = t[5528] ^ n[5529];
assign t[5530] = t[5529] ^ n[5530];
assign t[5531] = t[5530] ^ n[5531];
assign t[5532] = t[5531] ^ n[5532];
assign t[5533] = t[5532] ^ n[5533];
assign t[5534] = t[5533] ^ n[5534];
assign t[5535] = t[5534] ^ n[5535];
assign t[5536] = t[5535] ^ n[5536];
assign t[5537] = t[5536] ^ n[5537];
assign t[5538] = t[5537] ^ n[5538];
assign t[5539] = t[5538] ^ n[5539];
assign t[5540] = t[5539] ^ n[5540];
assign t[5541] = t[5540] ^ n[5541];
assign t[5542] = t[5541] ^ n[5542];
assign t[5543] = t[5542] ^ n[5543];
assign t[5544] = t[5543] ^ n[5544];
assign t[5545] = t[5544] ^ n[5545];
assign t[5546] = t[5545] ^ n[5546];
assign t[5547] = t[5546] ^ n[5547];
assign t[5548] = t[5547] ^ n[5548];
assign t[5549] = t[5548] ^ n[5549];
assign t[5550] = t[5549] ^ n[5550];
assign t[5551] = t[5550] ^ n[5551];
assign t[5552] = t[5551] ^ n[5552];
assign t[5553] = t[5552] ^ n[5553];
assign t[5554] = t[5553] ^ n[5554];
assign t[5555] = t[5554] ^ n[5555];
assign t[5556] = t[5555] ^ n[5556];
assign t[5557] = t[5556] ^ n[5557];
assign t[5558] = t[5557] ^ n[5558];
assign t[5559] = t[5558] ^ n[5559];
assign t[5560] = t[5559] ^ n[5560];
assign t[5561] = t[5560] ^ n[5561];
assign t[5562] = t[5561] ^ n[5562];
assign t[5563] = t[5562] ^ n[5563];
assign t[5564] = t[5563] ^ n[5564];
assign t[5565] = t[5564] ^ n[5565];
assign t[5566] = t[5565] ^ n[5566];
assign t[5567] = t[5566] ^ n[5567];
assign t[5568] = t[5567] ^ n[5568];
assign t[5569] = t[5568] ^ n[5569];
assign t[5570] = t[5569] ^ n[5570];
assign t[5571] = t[5570] ^ n[5571];
assign t[5572] = t[5571] ^ n[5572];
assign t[5573] = t[5572] ^ n[5573];
assign t[5574] = t[5573] ^ n[5574];
assign t[5575] = t[5574] ^ n[5575];
assign t[5576] = t[5575] ^ n[5576];
assign t[5577] = t[5576] ^ n[5577];
assign t[5578] = t[5577] ^ n[5578];
assign t[5579] = t[5578] ^ n[5579];
assign t[5580] = t[5579] ^ n[5580];
assign t[5581] = t[5580] ^ n[5581];
assign t[5582] = t[5581] ^ n[5582];
assign t[5583] = t[5582] ^ n[5583];
assign t[5584] = t[5583] ^ n[5584];
assign t[5585] = t[5584] ^ n[5585];
assign t[5586] = t[5585] ^ n[5586];
assign t[5587] = t[5586] ^ n[5587];
assign t[5588] = t[5587] ^ n[5588];
assign t[5589] = t[5588] ^ n[5589];
assign t[5590] = t[5589] ^ n[5590];
assign t[5591] = t[5590] ^ n[5591];
assign t[5592] = t[5591] ^ n[5592];
assign t[5593] = t[5592] ^ n[5593];
assign t[5594] = t[5593] ^ n[5594];
assign t[5595] = t[5594] ^ n[5595];
assign t[5596] = t[5595] ^ n[5596];
assign t[5597] = t[5596] ^ n[5597];
assign t[5598] = t[5597] ^ n[5598];
assign t[5599] = t[5598] ^ n[5599];
assign t[5600] = t[5599] ^ n[5600];
assign t[5601] = t[5600] ^ n[5601];
assign t[5602] = t[5601] ^ n[5602];
assign t[5603] = t[5602] ^ n[5603];
assign t[5604] = t[5603] ^ n[5604];
assign t[5605] = t[5604] ^ n[5605];
assign t[5606] = t[5605] ^ n[5606];
assign t[5607] = t[5606] ^ n[5607];
assign t[5608] = t[5607] ^ n[5608];
assign t[5609] = t[5608] ^ n[5609];
assign t[5610] = t[5609] ^ n[5610];
assign t[5611] = t[5610] ^ n[5611];
assign t[5612] = t[5611] ^ n[5612];
assign t[5613] = t[5612] ^ n[5613];
assign t[5614] = t[5613] ^ n[5614];
assign t[5615] = t[5614] ^ n[5615];
assign t[5616] = t[5615] ^ n[5616];
assign t[5617] = t[5616] ^ n[5617];
assign t[5618] = t[5617] ^ n[5618];
assign t[5619] = t[5618] ^ n[5619];
assign t[5620] = t[5619] ^ n[5620];
assign t[5621] = t[5620] ^ n[5621];
assign t[5622] = t[5621] ^ n[5622];
assign t[5623] = t[5622] ^ n[5623];
assign t[5624] = t[5623] ^ n[5624];
assign t[5625] = t[5624] ^ n[5625];
assign t[5626] = t[5625] ^ n[5626];
assign t[5627] = t[5626] ^ n[5627];
assign t[5628] = t[5627] ^ n[5628];
assign t[5629] = t[5628] ^ n[5629];
assign t[5630] = t[5629] ^ n[5630];
assign t[5631] = t[5630] ^ n[5631];
assign t[5632] = t[5631] ^ n[5632];
assign t[5633] = t[5632] ^ n[5633];
assign t[5634] = t[5633] ^ n[5634];
assign t[5635] = t[5634] ^ n[5635];
assign t[5636] = t[5635] ^ n[5636];
assign t[5637] = t[5636] ^ n[5637];
assign t[5638] = t[5637] ^ n[5638];
assign t[5639] = t[5638] ^ n[5639];
assign t[5640] = t[5639] ^ n[5640];
assign t[5641] = t[5640] ^ n[5641];
assign t[5642] = t[5641] ^ n[5642];
assign t[5643] = t[5642] ^ n[5643];
assign t[5644] = t[5643] ^ n[5644];
assign t[5645] = t[5644] ^ n[5645];
assign t[5646] = t[5645] ^ n[5646];
assign t[5647] = t[5646] ^ n[5647];
assign t[5648] = t[5647] ^ n[5648];
assign t[5649] = t[5648] ^ n[5649];
assign t[5650] = t[5649] ^ n[5650];
assign t[5651] = t[5650] ^ n[5651];
assign t[5652] = t[5651] ^ n[5652];
assign t[5653] = t[5652] ^ n[5653];
assign t[5654] = t[5653] ^ n[5654];
assign t[5655] = t[5654] ^ n[5655];
assign t[5656] = t[5655] ^ n[5656];
assign t[5657] = t[5656] ^ n[5657];
assign t[5658] = t[5657] ^ n[5658];
assign t[5659] = t[5658] ^ n[5659];
assign t[5660] = t[5659] ^ n[5660];
assign t[5661] = t[5660] ^ n[5661];
assign t[5662] = t[5661] ^ n[5662];
assign t[5663] = t[5662] ^ n[5663];
assign t[5664] = t[5663] ^ n[5664];
assign t[5665] = t[5664] ^ n[5665];
assign t[5666] = t[5665] ^ n[5666];
assign t[5667] = t[5666] ^ n[5667];
assign t[5668] = t[5667] ^ n[5668];
assign t[5669] = t[5668] ^ n[5669];
assign t[5670] = t[5669] ^ n[5670];
assign t[5671] = t[5670] ^ n[5671];
assign t[5672] = t[5671] ^ n[5672];
assign t[5673] = t[5672] ^ n[5673];
assign t[5674] = t[5673] ^ n[5674];
assign t[5675] = t[5674] ^ n[5675];
assign t[5676] = t[5675] ^ n[5676];
assign t[5677] = t[5676] ^ n[5677];
assign t[5678] = t[5677] ^ n[5678];
assign t[5679] = t[5678] ^ n[5679];
assign t[5680] = t[5679] ^ n[5680];
assign t[5681] = t[5680] ^ n[5681];
assign t[5682] = t[5681] ^ n[5682];
assign t[5683] = t[5682] ^ n[5683];
assign t[5684] = t[5683] ^ n[5684];
assign t[5685] = t[5684] ^ n[5685];
assign t[5686] = t[5685] ^ n[5686];
assign t[5687] = t[5686] ^ n[5687];
assign t[5688] = t[5687] ^ n[5688];
assign t[5689] = t[5688] ^ n[5689];
assign t[5690] = t[5689] ^ n[5690];
assign t[5691] = t[5690] ^ n[5691];
assign t[5692] = t[5691] ^ n[5692];
assign t[5693] = t[5692] ^ n[5693];
assign t[5694] = t[5693] ^ n[5694];
assign t[5695] = t[5694] ^ n[5695];
assign t[5696] = t[5695] ^ n[5696];
assign t[5697] = t[5696] ^ n[5697];
assign t[5698] = t[5697] ^ n[5698];
assign t[5699] = t[5698] ^ n[5699];
assign t[5700] = t[5699] ^ n[5700];
assign t[5701] = t[5700] ^ n[5701];
assign t[5702] = t[5701] ^ n[5702];
assign t[5703] = t[5702] ^ n[5703];
assign t[5704] = t[5703] ^ n[5704];
assign t[5705] = t[5704] ^ n[5705];
assign t[5706] = t[5705] ^ n[5706];
assign t[5707] = t[5706] ^ n[5707];
assign t[5708] = t[5707] ^ n[5708];
assign t[5709] = t[5708] ^ n[5709];
assign t[5710] = t[5709] ^ n[5710];
assign t[5711] = t[5710] ^ n[5711];
assign t[5712] = t[5711] ^ n[5712];
assign t[5713] = t[5712] ^ n[5713];
assign t[5714] = t[5713] ^ n[5714];
assign t[5715] = t[5714] ^ n[5715];
assign t[5716] = t[5715] ^ n[5716];
assign t[5717] = t[5716] ^ n[5717];
assign t[5718] = t[5717] ^ n[5718];
assign t[5719] = t[5718] ^ n[5719];
assign t[5720] = t[5719] ^ n[5720];
assign t[5721] = t[5720] ^ n[5721];
assign t[5722] = t[5721] ^ n[5722];
assign t[5723] = t[5722] ^ n[5723];
assign t[5724] = t[5723] ^ n[5724];
assign t[5725] = t[5724] ^ n[5725];
assign t[5726] = t[5725] ^ n[5726];
assign t[5727] = t[5726] ^ n[5727];
assign t[5728] = t[5727] ^ n[5728];
assign t[5729] = t[5728] ^ n[5729];
assign t[5730] = t[5729] ^ n[5730];
assign t[5731] = t[5730] ^ n[5731];
assign t[5732] = t[5731] ^ n[5732];
assign t[5733] = t[5732] ^ n[5733];
assign t[5734] = t[5733] ^ n[5734];
assign t[5735] = t[5734] ^ n[5735];
assign t[5736] = t[5735] ^ n[5736];
assign t[5737] = t[5736] ^ n[5737];
assign t[5738] = t[5737] ^ n[5738];
assign t[5739] = t[5738] ^ n[5739];
assign t[5740] = t[5739] ^ n[5740];
assign t[5741] = t[5740] ^ n[5741];
assign t[5742] = t[5741] ^ n[5742];
assign t[5743] = t[5742] ^ n[5743];
assign t[5744] = t[5743] ^ n[5744];
assign t[5745] = t[5744] ^ n[5745];
assign t[5746] = t[5745] ^ n[5746];
assign t[5747] = t[5746] ^ n[5747];
assign t[5748] = t[5747] ^ n[5748];
assign t[5749] = t[5748] ^ n[5749];
assign t[5750] = t[5749] ^ n[5750];
assign t[5751] = t[5750] ^ n[5751];
assign t[5752] = t[5751] ^ n[5752];
assign t[5753] = t[5752] ^ n[5753];
assign t[5754] = t[5753] ^ n[5754];
assign t[5755] = t[5754] ^ n[5755];
assign t[5756] = t[5755] ^ n[5756];
assign t[5757] = t[5756] ^ n[5757];
assign t[5758] = t[5757] ^ n[5758];
assign t[5759] = t[5758] ^ n[5759];
assign t[5760] = t[5759] ^ n[5760];
assign t[5761] = t[5760] ^ n[5761];
assign t[5762] = t[5761] ^ n[5762];
assign t[5763] = t[5762] ^ n[5763];
assign t[5764] = t[5763] ^ n[5764];
assign t[5765] = t[5764] ^ n[5765];
assign t[5766] = t[5765] ^ n[5766];
assign t[5767] = t[5766] ^ n[5767];
assign t[5768] = t[5767] ^ n[5768];
assign t[5769] = t[5768] ^ n[5769];
assign t[5770] = t[5769] ^ n[5770];
assign t[5771] = t[5770] ^ n[5771];
assign t[5772] = t[5771] ^ n[5772];
assign t[5773] = t[5772] ^ n[5773];
assign t[5774] = t[5773] ^ n[5774];
assign t[5775] = t[5774] ^ n[5775];
assign t[5776] = t[5775] ^ n[5776];
assign t[5777] = t[5776] ^ n[5777];
assign t[5778] = t[5777] ^ n[5778];
assign t[5779] = t[5778] ^ n[5779];
assign t[5780] = t[5779] ^ n[5780];
assign t[5781] = t[5780] ^ n[5781];
assign t[5782] = t[5781] ^ n[5782];
assign t[5783] = t[5782] ^ n[5783];
assign t[5784] = t[5783] ^ n[5784];
assign t[5785] = t[5784] ^ n[5785];
assign t[5786] = t[5785] ^ n[5786];
assign t[5787] = t[5786] ^ n[5787];
assign t[5788] = t[5787] ^ n[5788];
assign t[5789] = t[5788] ^ n[5789];
assign t[5790] = t[5789] ^ n[5790];
assign t[5791] = t[5790] ^ n[5791];
assign t[5792] = t[5791] ^ n[5792];
assign t[5793] = t[5792] ^ n[5793];
assign t[5794] = t[5793] ^ n[5794];
assign t[5795] = t[5794] ^ n[5795];
assign t[5796] = t[5795] ^ n[5796];
assign t[5797] = t[5796] ^ n[5797];
assign t[5798] = t[5797] ^ n[5798];
assign t[5799] = t[5798] ^ n[5799];
assign t[5800] = t[5799] ^ n[5800];
assign t[5801] = t[5800] ^ n[5801];
assign t[5802] = t[5801] ^ n[5802];
assign t[5803] = t[5802] ^ n[5803];
assign t[5804] = t[5803] ^ n[5804];
assign t[5805] = t[5804] ^ n[5805];
assign t[5806] = t[5805] ^ n[5806];
assign t[5807] = t[5806] ^ n[5807];
assign t[5808] = t[5807] ^ n[5808];
assign t[5809] = t[5808] ^ n[5809];
assign t[5810] = t[5809] ^ n[5810];
assign t[5811] = t[5810] ^ n[5811];
assign t[5812] = t[5811] ^ n[5812];
assign t[5813] = t[5812] ^ n[5813];
assign t[5814] = t[5813] ^ n[5814];
assign t[5815] = t[5814] ^ n[5815];
assign t[5816] = t[5815] ^ n[5816];
assign t[5817] = t[5816] ^ n[5817];
assign t[5818] = t[5817] ^ n[5818];
assign t[5819] = t[5818] ^ n[5819];
assign t[5820] = t[5819] ^ n[5820];
assign t[5821] = t[5820] ^ n[5821];
assign t[5822] = t[5821] ^ n[5822];
assign t[5823] = t[5822] ^ n[5823];
assign t[5824] = t[5823] ^ n[5824];
assign t[5825] = t[5824] ^ n[5825];
assign t[5826] = t[5825] ^ n[5826];
assign t[5827] = t[5826] ^ n[5827];
assign t[5828] = t[5827] ^ n[5828];
assign t[5829] = t[5828] ^ n[5829];
assign t[5830] = t[5829] ^ n[5830];
assign t[5831] = t[5830] ^ n[5831];
assign t[5832] = t[5831] ^ n[5832];
assign t[5833] = t[5832] ^ n[5833];
assign t[5834] = t[5833] ^ n[5834];
assign t[5835] = t[5834] ^ n[5835];
assign t[5836] = t[5835] ^ n[5836];
assign t[5837] = t[5836] ^ n[5837];
assign t[5838] = t[5837] ^ n[5838];
assign t[5839] = t[5838] ^ n[5839];
assign t[5840] = t[5839] ^ n[5840];
assign t[5841] = t[5840] ^ n[5841];
assign t[5842] = t[5841] ^ n[5842];
assign t[5843] = t[5842] ^ n[5843];
assign t[5844] = t[5843] ^ n[5844];
assign t[5845] = t[5844] ^ n[5845];
assign t[5846] = t[5845] ^ n[5846];
assign t[5847] = t[5846] ^ n[5847];
assign t[5848] = t[5847] ^ n[5848];
assign t[5849] = t[5848] ^ n[5849];
assign t[5850] = t[5849] ^ n[5850];
assign t[5851] = t[5850] ^ n[5851];
assign t[5852] = t[5851] ^ n[5852];
assign t[5853] = t[5852] ^ n[5853];
assign t[5854] = t[5853] ^ n[5854];
assign t[5855] = t[5854] ^ n[5855];
assign t[5856] = t[5855] ^ n[5856];
assign t[5857] = t[5856] ^ n[5857];
assign t[5858] = t[5857] ^ n[5858];
assign t[5859] = t[5858] ^ n[5859];
assign t[5860] = t[5859] ^ n[5860];
assign t[5861] = t[5860] ^ n[5861];
assign t[5862] = t[5861] ^ n[5862];
assign t[5863] = t[5862] ^ n[5863];
assign t[5864] = t[5863] ^ n[5864];
assign t[5865] = t[5864] ^ n[5865];
assign t[5866] = t[5865] ^ n[5866];
assign t[5867] = t[5866] ^ n[5867];
assign t[5868] = t[5867] ^ n[5868];
assign t[5869] = t[5868] ^ n[5869];
assign t[5870] = t[5869] ^ n[5870];
assign t[5871] = t[5870] ^ n[5871];
assign t[5872] = t[5871] ^ n[5872];
assign t[5873] = t[5872] ^ n[5873];
assign t[5874] = t[5873] ^ n[5874];
assign t[5875] = t[5874] ^ n[5875];
assign t[5876] = t[5875] ^ n[5876];
assign t[5877] = t[5876] ^ n[5877];
assign t[5878] = t[5877] ^ n[5878];
assign t[5879] = t[5878] ^ n[5879];
assign t[5880] = t[5879] ^ n[5880];
assign t[5881] = t[5880] ^ n[5881];
assign t[5882] = t[5881] ^ n[5882];
assign t[5883] = t[5882] ^ n[5883];
assign t[5884] = t[5883] ^ n[5884];
assign t[5885] = t[5884] ^ n[5885];
assign t[5886] = t[5885] ^ n[5886];
assign t[5887] = t[5886] ^ n[5887];
assign t[5888] = t[5887] ^ n[5888];
assign t[5889] = t[5888] ^ n[5889];
assign t[5890] = t[5889] ^ n[5890];
assign t[5891] = t[5890] ^ n[5891];
assign t[5892] = t[5891] ^ n[5892];
assign t[5893] = t[5892] ^ n[5893];
assign t[5894] = t[5893] ^ n[5894];
assign t[5895] = t[5894] ^ n[5895];
assign t[5896] = t[5895] ^ n[5896];
assign t[5897] = t[5896] ^ n[5897];
assign t[5898] = t[5897] ^ n[5898];
assign t[5899] = t[5898] ^ n[5899];
assign t[5900] = t[5899] ^ n[5900];
assign t[5901] = t[5900] ^ n[5901];
assign t[5902] = t[5901] ^ n[5902];
assign t[5903] = t[5902] ^ n[5903];
assign t[5904] = t[5903] ^ n[5904];
assign t[5905] = t[5904] ^ n[5905];
assign t[5906] = t[5905] ^ n[5906];
assign t[5907] = t[5906] ^ n[5907];
assign t[5908] = t[5907] ^ n[5908];
assign t[5909] = t[5908] ^ n[5909];
assign t[5910] = t[5909] ^ n[5910];
assign t[5911] = t[5910] ^ n[5911];
assign t[5912] = t[5911] ^ n[5912];
assign t[5913] = t[5912] ^ n[5913];
assign t[5914] = t[5913] ^ n[5914];
assign t[5915] = t[5914] ^ n[5915];
assign t[5916] = t[5915] ^ n[5916];
assign t[5917] = t[5916] ^ n[5917];
assign t[5918] = t[5917] ^ n[5918];
assign t[5919] = t[5918] ^ n[5919];
assign t[5920] = t[5919] ^ n[5920];
assign t[5921] = t[5920] ^ n[5921];
assign t[5922] = t[5921] ^ n[5922];
assign t[5923] = t[5922] ^ n[5923];
assign t[5924] = t[5923] ^ n[5924];
assign t[5925] = t[5924] ^ n[5925];
assign t[5926] = t[5925] ^ n[5926];
assign t[5927] = t[5926] ^ n[5927];
assign t[5928] = t[5927] ^ n[5928];
assign t[5929] = t[5928] ^ n[5929];
assign t[5930] = t[5929] ^ n[5930];
assign t[5931] = t[5930] ^ n[5931];
assign t[5932] = t[5931] ^ n[5932];
assign t[5933] = t[5932] ^ n[5933];
assign t[5934] = t[5933] ^ n[5934];
assign t[5935] = t[5934] ^ n[5935];
assign t[5936] = t[5935] ^ n[5936];
assign t[5937] = t[5936] ^ n[5937];
assign t[5938] = t[5937] ^ n[5938];
assign t[5939] = t[5938] ^ n[5939];
assign t[5940] = t[5939] ^ n[5940];
assign t[5941] = t[5940] ^ n[5941];
assign t[5942] = t[5941] ^ n[5942];
assign t[5943] = t[5942] ^ n[5943];
assign t[5944] = t[5943] ^ n[5944];
assign t[5945] = t[5944] ^ n[5945];
assign t[5946] = t[5945] ^ n[5946];
assign t[5947] = t[5946] ^ n[5947];
assign t[5948] = t[5947] ^ n[5948];
assign t[5949] = t[5948] ^ n[5949];
assign t[5950] = t[5949] ^ n[5950];
assign t[5951] = t[5950] ^ n[5951];
assign t[5952] = t[5951] ^ n[5952];
assign t[5953] = t[5952] ^ n[5953];
assign t[5954] = t[5953] ^ n[5954];
assign t[5955] = t[5954] ^ n[5955];
assign t[5956] = t[5955] ^ n[5956];
assign t[5957] = t[5956] ^ n[5957];
assign t[5958] = t[5957] ^ n[5958];
assign t[5959] = t[5958] ^ n[5959];
assign t[5960] = t[5959] ^ n[5960];
assign t[5961] = t[5960] ^ n[5961];
assign t[5962] = t[5961] ^ n[5962];
assign t[5963] = t[5962] ^ n[5963];
assign t[5964] = t[5963] ^ n[5964];
assign t[5965] = t[5964] ^ n[5965];
assign t[5966] = t[5965] ^ n[5966];
assign t[5967] = t[5966] ^ n[5967];
assign t[5968] = t[5967] ^ n[5968];
assign t[5969] = t[5968] ^ n[5969];
assign t[5970] = t[5969] ^ n[5970];
assign t[5971] = t[5970] ^ n[5971];
assign t[5972] = t[5971] ^ n[5972];
assign t[5973] = t[5972] ^ n[5973];
assign t[5974] = t[5973] ^ n[5974];
assign t[5975] = t[5974] ^ n[5975];
assign t[5976] = t[5975] ^ n[5976];
assign t[5977] = t[5976] ^ n[5977];
assign t[5978] = t[5977] ^ n[5978];
assign t[5979] = t[5978] ^ n[5979];
assign t[5980] = t[5979] ^ n[5980];
assign t[5981] = t[5980] ^ n[5981];
assign t[5982] = t[5981] ^ n[5982];
assign t[5983] = t[5982] ^ n[5983];
assign t[5984] = t[5983] ^ n[5984];
assign t[5985] = t[5984] ^ n[5985];
assign t[5986] = t[5985] ^ n[5986];
assign t[5987] = t[5986] ^ n[5987];
assign t[5988] = t[5987] ^ n[5988];
assign t[5989] = t[5988] ^ n[5989];
assign t[5990] = t[5989] ^ n[5990];
assign t[5991] = t[5990] ^ n[5991];
assign t[5992] = t[5991] ^ n[5992];
assign t[5993] = t[5992] ^ n[5993];
assign t[5994] = t[5993] ^ n[5994];
assign t[5995] = t[5994] ^ n[5995];
assign t[5996] = t[5995] ^ n[5996];
assign t[5997] = t[5996] ^ n[5997];
assign t[5998] = t[5997] ^ n[5998];
assign t[5999] = t[5998] ^ n[5999];
assign t[6000] = t[5999] ^ n[6000];
assign t[6001] = t[6000] ^ n[6001];
assign t[6002] = t[6001] ^ n[6002];
assign t[6003] = t[6002] ^ n[6003];
assign t[6004] = t[6003] ^ n[6004];
assign t[6005] = t[6004] ^ n[6005];
assign t[6006] = t[6005] ^ n[6006];
assign t[6007] = t[6006] ^ n[6007];
assign t[6008] = t[6007] ^ n[6008];
assign t[6009] = t[6008] ^ n[6009];
assign t[6010] = t[6009] ^ n[6010];
assign t[6011] = t[6010] ^ n[6011];
assign t[6012] = t[6011] ^ n[6012];
assign t[6013] = t[6012] ^ n[6013];
assign t[6014] = t[6013] ^ n[6014];
assign t[6015] = t[6014] ^ n[6015];
assign t[6016] = t[6015] ^ n[6016];
assign t[6017] = t[6016] ^ n[6017];
assign t[6018] = t[6017] ^ n[6018];
assign t[6019] = t[6018] ^ n[6019];
assign t[6020] = t[6019] ^ n[6020];
assign t[6021] = t[6020] ^ n[6021];
assign t[6022] = t[6021] ^ n[6022];
assign t[6023] = t[6022] ^ n[6023];
assign t[6024] = t[6023] ^ n[6024];
assign t[6025] = t[6024] ^ n[6025];
assign t[6026] = t[6025] ^ n[6026];
assign t[6027] = t[6026] ^ n[6027];
assign t[6028] = t[6027] ^ n[6028];
assign t[6029] = t[6028] ^ n[6029];
assign t[6030] = t[6029] ^ n[6030];
assign t[6031] = t[6030] ^ n[6031];
assign t[6032] = t[6031] ^ n[6032];
assign t[6033] = t[6032] ^ n[6033];
assign t[6034] = t[6033] ^ n[6034];
assign t[6035] = t[6034] ^ n[6035];
assign t[6036] = t[6035] ^ n[6036];
assign t[6037] = t[6036] ^ n[6037];
assign t[6038] = t[6037] ^ n[6038];
assign t[6039] = t[6038] ^ n[6039];
assign t[6040] = t[6039] ^ n[6040];
assign t[6041] = t[6040] ^ n[6041];
assign t[6042] = t[6041] ^ n[6042];
assign t[6043] = t[6042] ^ n[6043];
assign t[6044] = t[6043] ^ n[6044];
assign t[6045] = t[6044] ^ n[6045];
assign t[6046] = t[6045] ^ n[6046];
assign t[6047] = t[6046] ^ n[6047];
assign t[6048] = t[6047] ^ n[6048];
assign t[6049] = t[6048] ^ n[6049];
assign t[6050] = t[6049] ^ n[6050];
assign t[6051] = t[6050] ^ n[6051];
assign t[6052] = t[6051] ^ n[6052];
assign t[6053] = t[6052] ^ n[6053];
assign t[6054] = t[6053] ^ n[6054];
assign t[6055] = t[6054] ^ n[6055];
assign t[6056] = t[6055] ^ n[6056];
assign t[6057] = t[6056] ^ n[6057];
assign t[6058] = t[6057] ^ n[6058];
assign t[6059] = t[6058] ^ n[6059];
assign t[6060] = t[6059] ^ n[6060];
assign t[6061] = t[6060] ^ n[6061];
assign t[6062] = t[6061] ^ n[6062];
assign t[6063] = t[6062] ^ n[6063];
assign t[6064] = t[6063] ^ n[6064];
assign t[6065] = t[6064] ^ n[6065];
assign t[6066] = t[6065] ^ n[6066];
assign t[6067] = t[6066] ^ n[6067];
assign t[6068] = t[6067] ^ n[6068];
assign t[6069] = t[6068] ^ n[6069];
assign t[6070] = t[6069] ^ n[6070];
assign t[6071] = t[6070] ^ n[6071];
assign t[6072] = t[6071] ^ n[6072];
assign t[6073] = t[6072] ^ n[6073];
assign t[6074] = t[6073] ^ n[6074];
assign t[6075] = t[6074] ^ n[6075];
assign t[6076] = t[6075] ^ n[6076];
assign t[6077] = t[6076] ^ n[6077];
assign t[6078] = t[6077] ^ n[6078];
assign t[6079] = t[6078] ^ n[6079];
assign t[6080] = t[6079] ^ n[6080];
assign t[6081] = t[6080] ^ n[6081];
assign t[6082] = t[6081] ^ n[6082];
assign t[6083] = t[6082] ^ n[6083];
assign t[6084] = t[6083] ^ n[6084];
assign t[6085] = t[6084] ^ n[6085];
assign t[6086] = t[6085] ^ n[6086];
assign t[6087] = t[6086] ^ n[6087];
assign t[6088] = t[6087] ^ n[6088];
assign t[6089] = t[6088] ^ n[6089];
assign t[6090] = t[6089] ^ n[6090];
assign t[6091] = t[6090] ^ n[6091];
assign t[6092] = t[6091] ^ n[6092];
assign t[6093] = t[6092] ^ n[6093];
assign t[6094] = t[6093] ^ n[6094];
assign t[6095] = t[6094] ^ n[6095];
assign t[6096] = t[6095] ^ n[6096];
assign t[6097] = t[6096] ^ n[6097];
assign t[6098] = t[6097] ^ n[6098];
assign t[6099] = t[6098] ^ n[6099];
assign t[6100] = t[6099] ^ n[6100];
assign t[6101] = t[6100] ^ n[6101];
assign t[6102] = t[6101] ^ n[6102];
assign t[6103] = t[6102] ^ n[6103];
assign t[6104] = t[6103] ^ n[6104];
assign t[6105] = t[6104] ^ n[6105];
assign t[6106] = t[6105] ^ n[6106];
assign t[6107] = t[6106] ^ n[6107];
assign t[6108] = t[6107] ^ n[6108];
assign t[6109] = t[6108] ^ n[6109];
assign t[6110] = t[6109] ^ n[6110];
assign t[6111] = t[6110] ^ n[6111];
assign t[6112] = t[6111] ^ n[6112];
assign t[6113] = t[6112] ^ n[6113];
assign t[6114] = t[6113] ^ n[6114];
assign t[6115] = t[6114] ^ n[6115];
assign t[6116] = t[6115] ^ n[6116];
assign t[6117] = t[6116] ^ n[6117];
assign t[6118] = t[6117] ^ n[6118];
assign t[6119] = t[6118] ^ n[6119];
assign t[6120] = t[6119] ^ n[6120];
assign t[6121] = t[6120] ^ n[6121];
assign t[6122] = t[6121] ^ n[6122];
assign t[6123] = t[6122] ^ n[6123];
assign t[6124] = t[6123] ^ n[6124];
assign t[6125] = t[6124] ^ n[6125];
assign t[6126] = t[6125] ^ n[6126];
assign t[6127] = t[6126] ^ n[6127];
assign t[6128] = t[6127] ^ n[6128];
assign t[6129] = t[6128] ^ n[6129];
assign t[6130] = t[6129] ^ n[6130];
assign t[6131] = t[6130] ^ n[6131];
assign t[6132] = t[6131] ^ n[6132];
assign t[6133] = t[6132] ^ n[6133];
assign t[6134] = t[6133] ^ n[6134];
assign t[6135] = t[6134] ^ n[6135];
assign t[6136] = t[6135] ^ n[6136];
assign t[6137] = t[6136] ^ n[6137];
assign t[6138] = t[6137] ^ n[6138];
assign t[6139] = t[6138] ^ n[6139];
assign t[6140] = t[6139] ^ n[6140];
assign t[6141] = t[6140] ^ n[6141];
assign t[6142] = t[6141] ^ n[6142];
assign t[6143] = t[6142] ^ n[6143];
assign t[6144] = t[6143] ^ n[6144];
assign t[6145] = t[6144] ^ n[6145];
assign t[6146] = t[6145] ^ n[6146];
assign t[6147] = t[6146] ^ n[6147];
assign t[6148] = t[6147] ^ n[6148];
assign t[6149] = t[6148] ^ n[6149];
assign t[6150] = t[6149] ^ n[6150];
assign t[6151] = t[6150] ^ n[6151];
assign t[6152] = t[6151] ^ n[6152];
assign t[6153] = t[6152] ^ n[6153];
assign t[6154] = t[6153] ^ n[6154];
assign t[6155] = t[6154] ^ n[6155];
assign t[6156] = t[6155] ^ n[6156];
assign t[6157] = t[6156] ^ n[6157];
assign t[6158] = t[6157] ^ n[6158];
assign t[6159] = t[6158] ^ n[6159];
assign t[6160] = t[6159] ^ n[6160];
assign t[6161] = t[6160] ^ n[6161];
assign t[6162] = t[6161] ^ n[6162];
assign t[6163] = t[6162] ^ n[6163];
assign t[6164] = t[6163] ^ n[6164];
assign t[6165] = t[6164] ^ n[6165];
assign t[6166] = t[6165] ^ n[6166];
assign t[6167] = t[6166] ^ n[6167];
assign t[6168] = t[6167] ^ n[6168];
assign t[6169] = t[6168] ^ n[6169];
assign t[6170] = t[6169] ^ n[6170];
assign t[6171] = t[6170] ^ n[6171];
assign t[6172] = t[6171] ^ n[6172];
assign t[6173] = t[6172] ^ n[6173];
assign t[6174] = t[6173] ^ n[6174];
assign t[6175] = t[6174] ^ n[6175];
assign t[6176] = t[6175] ^ n[6176];
assign t[6177] = t[6176] ^ n[6177];
assign t[6178] = t[6177] ^ n[6178];
assign t[6179] = t[6178] ^ n[6179];
assign t[6180] = t[6179] ^ n[6180];
assign t[6181] = t[6180] ^ n[6181];
assign t[6182] = t[6181] ^ n[6182];
assign t[6183] = t[6182] ^ n[6183];
assign t[6184] = t[6183] ^ n[6184];
assign t[6185] = t[6184] ^ n[6185];
assign t[6186] = t[6185] ^ n[6186];
assign t[6187] = t[6186] ^ n[6187];
assign t[6188] = t[6187] ^ n[6188];
assign t[6189] = t[6188] ^ n[6189];
assign t[6190] = t[6189] ^ n[6190];
assign t[6191] = t[6190] ^ n[6191];
assign t[6192] = t[6191] ^ n[6192];
assign t[6193] = t[6192] ^ n[6193];
assign t[6194] = t[6193] ^ n[6194];
assign t[6195] = t[6194] ^ n[6195];
assign t[6196] = t[6195] ^ n[6196];
assign t[6197] = t[6196] ^ n[6197];
assign t[6198] = t[6197] ^ n[6198];
assign t[6199] = t[6198] ^ n[6199];
assign t[6200] = t[6199] ^ n[6200];
assign t[6201] = t[6200] ^ n[6201];
assign t[6202] = t[6201] ^ n[6202];
assign t[6203] = t[6202] ^ n[6203];
assign t[6204] = t[6203] ^ n[6204];
assign t[6205] = t[6204] ^ n[6205];
assign t[6206] = t[6205] ^ n[6206];
assign t[6207] = t[6206] ^ n[6207];
assign t[6208] = t[6207] ^ n[6208];
assign t[6209] = t[6208] ^ n[6209];
assign t[6210] = t[6209] ^ n[6210];
assign t[6211] = t[6210] ^ n[6211];
assign t[6212] = t[6211] ^ n[6212];
assign t[6213] = t[6212] ^ n[6213];
assign t[6214] = t[6213] ^ n[6214];
assign t[6215] = t[6214] ^ n[6215];
assign t[6216] = t[6215] ^ n[6216];
assign t[6217] = t[6216] ^ n[6217];
assign t[6218] = t[6217] ^ n[6218];
assign t[6219] = t[6218] ^ n[6219];
assign t[6220] = t[6219] ^ n[6220];
assign t[6221] = t[6220] ^ n[6221];
assign t[6222] = t[6221] ^ n[6222];
assign t[6223] = t[6222] ^ n[6223];
assign t[6224] = t[6223] ^ n[6224];
assign t[6225] = t[6224] ^ n[6225];
assign t[6226] = t[6225] ^ n[6226];
assign t[6227] = t[6226] ^ n[6227];
assign t[6228] = t[6227] ^ n[6228];
assign t[6229] = t[6228] ^ n[6229];
assign t[6230] = t[6229] ^ n[6230];
assign t[6231] = t[6230] ^ n[6231];
assign t[6232] = t[6231] ^ n[6232];
assign t[6233] = t[6232] ^ n[6233];
assign t[6234] = t[6233] ^ n[6234];
assign t[6235] = t[6234] ^ n[6235];
assign t[6236] = t[6235] ^ n[6236];
assign t[6237] = t[6236] ^ n[6237];
assign t[6238] = t[6237] ^ n[6238];
assign t[6239] = t[6238] ^ n[6239];
assign t[6240] = t[6239] ^ n[6240];
assign t[6241] = t[6240] ^ n[6241];
assign t[6242] = t[6241] ^ n[6242];
assign t[6243] = t[6242] ^ n[6243];
assign t[6244] = t[6243] ^ n[6244];
assign t[6245] = t[6244] ^ n[6245];
assign t[6246] = t[6245] ^ n[6246];
assign t[6247] = t[6246] ^ n[6247];
assign t[6248] = t[6247] ^ n[6248];
assign t[6249] = t[6248] ^ n[6249];
assign t[6250] = t[6249] ^ n[6250];
assign t[6251] = t[6250] ^ n[6251];
assign t[6252] = t[6251] ^ n[6252];
assign t[6253] = t[6252] ^ n[6253];
assign t[6254] = t[6253] ^ n[6254];
assign t[6255] = t[6254] ^ n[6255];
assign t[6256] = t[6255] ^ n[6256];
assign t[6257] = t[6256] ^ n[6257];
assign t[6258] = t[6257] ^ n[6258];
assign t[6259] = t[6258] ^ n[6259];
assign t[6260] = t[6259] ^ n[6260];
assign t[6261] = t[6260] ^ n[6261];
assign t[6262] = t[6261] ^ n[6262];
assign t[6263] = t[6262] ^ n[6263];
assign t[6264] = t[6263] ^ n[6264];
assign t[6265] = t[6264] ^ n[6265];
assign t[6266] = t[6265] ^ n[6266];
assign t[6267] = t[6266] ^ n[6267];
assign t[6268] = t[6267] ^ n[6268];
assign t[6269] = t[6268] ^ n[6269];
assign t[6270] = t[6269] ^ n[6270];
assign t[6271] = t[6270] ^ n[6271];
assign t[6272] = t[6271] ^ n[6272];
assign t[6273] = t[6272] ^ n[6273];
assign t[6274] = t[6273] ^ n[6274];
assign t[6275] = t[6274] ^ n[6275];
assign t[6276] = t[6275] ^ n[6276];
assign t[6277] = t[6276] ^ n[6277];
assign t[6278] = t[6277] ^ n[6278];
assign t[6279] = t[6278] ^ n[6279];
assign t[6280] = t[6279] ^ n[6280];
assign t[6281] = t[6280] ^ n[6281];
assign t[6282] = t[6281] ^ n[6282];
assign t[6283] = t[6282] ^ n[6283];
assign t[6284] = t[6283] ^ n[6284];
assign t[6285] = t[6284] ^ n[6285];
assign t[6286] = t[6285] ^ n[6286];
assign t[6287] = t[6286] ^ n[6287];
assign t[6288] = t[6287] ^ n[6288];
assign t[6289] = t[6288] ^ n[6289];
assign t[6290] = t[6289] ^ n[6290];
assign t[6291] = t[6290] ^ n[6291];
assign t[6292] = t[6291] ^ n[6292];
assign t[6293] = t[6292] ^ n[6293];
assign t[6294] = t[6293] ^ n[6294];
assign t[6295] = t[6294] ^ n[6295];
assign t[6296] = t[6295] ^ n[6296];
assign t[6297] = t[6296] ^ n[6297];
assign t[6298] = t[6297] ^ n[6298];
assign t[6299] = t[6298] ^ n[6299];
assign t[6300] = t[6299] ^ n[6300];
assign t[6301] = t[6300] ^ n[6301];
assign t[6302] = t[6301] ^ n[6302];
assign t[6303] = t[6302] ^ n[6303];
assign t[6304] = t[6303] ^ n[6304];
assign t[6305] = t[6304] ^ n[6305];
assign t[6306] = t[6305] ^ n[6306];
assign t[6307] = t[6306] ^ n[6307];
assign t[6308] = t[6307] ^ n[6308];
assign t[6309] = t[6308] ^ n[6309];
assign t[6310] = t[6309] ^ n[6310];
assign t[6311] = t[6310] ^ n[6311];
assign t[6312] = t[6311] ^ n[6312];
assign t[6313] = t[6312] ^ n[6313];
assign t[6314] = t[6313] ^ n[6314];
assign t[6315] = t[6314] ^ n[6315];
assign t[6316] = t[6315] ^ n[6316];
assign t[6317] = t[6316] ^ n[6317];
assign t[6318] = t[6317] ^ n[6318];
assign t[6319] = t[6318] ^ n[6319];
assign t[6320] = t[6319] ^ n[6320];
assign t[6321] = t[6320] ^ n[6321];
assign t[6322] = t[6321] ^ n[6322];
assign t[6323] = t[6322] ^ n[6323];
assign t[6324] = t[6323] ^ n[6324];
assign t[6325] = t[6324] ^ n[6325];
assign t[6326] = t[6325] ^ n[6326];
assign t[6327] = t[6326] ^ n[6327];
assign t[6328] = t[6327] ^ n[6328];
assign t[6329] = t[6328] ^ n[6329];
assign t[6330] = t[6329] ^ n[6330];
assign t[6331] = t[6330] ^ n[6331];
assign t[6332] = t[6331] ^ n[6332];
assign t[6333] = t[6332] ^ n[6333];
assign t[6334] = t[6333] ^ n[6334];
assign t[6335] = t[6334] ^ n[6335];
assign t[6336] = t[6335] ^ n[6336];
assign t[6337] = t[6336] ^ n[6337];
assign t[6338] = t[6337] ^ n[6338];
assign t[6339] = t[6338] ^ n[6339];
assign t[6340] = t[6339] ^ n[6340];
assign t[6341] = t[6340] ^ n[6341];
assign t[6342] = t[6341] ^ n[6342];
assign t[6343] = t[6342] ^ n[6343];
assign t[6344] = t[6343] ^ n[6344];
assign t[6345] = t[6344] ^ n[6345];
assign t[6346] = t[6345] ^ n[6346];
assign t[6347] = t[6346] ^ n[6347];
assign t[6348] = t[6347] ^ n[6348];
assign t[6349] = t[6348] ^ n[6349];
assign t[6350] = t[6349] ^ n[6350];
assign t[6351] = t[6350] ^ n[6351];
assign t[6352] = t[6351] ^ n[6352];
assign t[6353] = t[6352] ^ n[6353];
assign t[6354] = t[6353] ^ n[6354];
assign t[6355] = t[6354] ^ n[6355];
assign t[6356] = t[6355] ^ n[6356];
assign t[6357] = t[6356] ^ n[6357];
assign t[6358] = t[6357] ^ n[6358];
assign t[6359] = t[6358] ^ n[6359];
assign t[6360] = t[6359] ^ n[6360];
assign t[6361] = t[6360] ^ n[6361];
assign t[6362] = t[6361] ^ n[6362];
assign t[6363] = t[6362] ^ n[6363];
assign t[6364] = t[6363] ^ n[6364];
assign t[6365] = t[6364] ^ n[6365];
assign t[6366] = t[6365] ^ n[6366];
assign t[6367] = t[6366] ^ n[6367];
assign t[6368] = t[6367] ^ n[6368];
assign t[6369] = t[6368] ^ n[6369];
assign t[6370] = t[6369] ^ n[6370];
assign t[6371] = t[6370] ^ n[6371];
assign t[6372] = t[6371] ^ n[6372];
assign t[6373] = t[6372] ^ n[6373];
assign t[6374] = t[6373] ^ n[6374];
assign t[6375] = t[6374] ^ n[6375];
assign t[6376] = t[6375] ^ n[6376];
assign t[6377] = t[6376] ^ n[6377];
assign t[6378] = t[6377] ^ n[6378];
assign t[6379] = t[6378] ^ n[6379];
assign t[6380] = t[6379] ^ n[6380];
assign t[6381] = t[6380] ^ n[6381];
assign t[6382] = t[6381] ^ n[6382];
assign t[6383] = t[6382] ^ n[6383];
assign t[6384] = t[6383] ^ n[6384];
assign t[6385] = t[6384] ^ n[6385];
assign t[6386] = t[6385] ^ n[6386];
assign t[6387] = t[6386] ^ n[6387];
assign t[6388] = t[6387] ^ n[6388];
assign t[6389] = t[6388] ^ n[6389];
assign t[6390] = t[6389] ^ n[6390];
assign t[6391] = t[6390] ^ n[6391];
assign t[6392] = t[6391] ^ n[6392];
assign t[6393] = t[6392] ^ n[6393];
assign t[6394] = t[6393] ^ n[6394];
assign t[6395] = t[6394] ^ n[6395];
assign t[6396] = t[6395] ^ n[6396];
assign t[6397] = t[6396] ^ n[6397];
assign t[6398] = t[6397] ^ n[6398];
assign t[6399] = t[6398] ^ n[6399];
assign t[6400] = t[6399] ^ n[6400];
assign t[6401] = t[6400] ^ n[6401];
assign t[6402] = t[6401] ^ n[6402];
assign t[6403] = t[6402] ^ n[6403];
assign t[6404] = t[6403] ^ n[6404];
assign t[6405] = t[6404] ^ n[6405];
assign t[6406] = t[6405] ^ n[6406];
assign t[6407] = t[6406] ^ n[6407];
assign t[6408] = t[6407] ^ n[6408];
assign t[6409] = t[6408] ^ n[6409];
assign t[6410] = t[6409] ^ n[6410];
assign t[6411] = t[6410] ^ n[6411];
assign t[6412] = t[6411] ^ n[6412];
assign t[6413] = t[6412] ^ n[6413];
assign t[6414] = t[6413] ^ n[6414];
assign t[6415] = t[6414] ^ n[6415];
assign t[6416] = t[6415] ^ n[6416];
assign t[6417] = t[6416] ^ n[6417];
assign t[6418] = t[6417] ^ n[6418];
assign t[6419] = t[6418] ^ n[6419];
assign t[6420] = t[6419] ^ n[6420];
assign t[6421] = t[6420] ^ n[6421];
assign t[6422] = t[6421] ^ n[6422];
assign t[6423] = t[6422] ^ n[6423];
assign t[6424] = t[6423] ^ n[6424];
assign t[6425] = t[6424] ^ n[6425];
assign t[6426] = t[6425] ^ n[6426];
assign t[6427] = t[6426] ^ n[6427];
assign t[6428] = t[6427] ^ n[6428];
assign t[6429] = t[6428] ^ n[6429];
assign t[6430] = t[6429] ^ n[6430];
assign t[6431] = t[6430] ^ n[6431];
assign t[6432] = t[6431] ^ n[6432];
assign t[6433] = t[6432] ^ n[6433];
assign t[6434] = t[6433] ^ n[6434];
assign t[6435] = t[6434] ^ n[6435];
assign t[6436] = t[6435] ^ n[6436];
assign t[6437] = t[6436] ^ n[6437];
assign t[6438] = t[6437] ^ n[6438];
assign t[6439] = t[6438] ^ n[6439];
assign t[6440] = t[6439] ^ n[6440];
assign t[6441] = t[6440] ^ n[6441];
assign t[6442] = t[6441] ^ n[6442];
assign t[6443] = t[6442] ^ n[6443];
assign t[6444] = t[6443] ^ n[6444];
assign t[6445] = t[6444] ^ n[6445];
assign t[6446] = t[6445] ^ n[6446];
assign t[6447] = t[6446] ^ n[6447];
assign t[6448] = t[6447] ^ n[6448];
assign t[6449] = t[6448] ^ n[6449];
assign t[6450] = t[6449] ^ n[6450];
assign t[6451] = t[6450] ^ n[6451];
assign t[6452] = t[6451] ^ n[6452];
assign t[6453] = t[6452] ^ n[6453];
assign t[6454] = t[6453] ^ n[6454];
assign t[6455] = t[6454] ^ n[6455];
assign t[6456] = t[6455] ^ n[6456];
assign t[6457] = t[6456] ^ n[6457];
assign t[6458] = t[6457] ^ n[6458];
assign t[6459] = t[6458] ^ n[6459];
assign t[6460] = t[6459] ^ n[6460];
assign t[6461] = t[6460] ^ n[6461];
assign t[6462] = t[6461] ^ n[6462];
assign t[6463] = t[6462] ^ n[6463];
assign t[6464] = t[6463] ^ n[6464];
assign t[6465] = t[6464] ^ n[6465];
assign t[6466] = t[6465] ^ n[6466];
assign t[6467] = t[6466] ^ n[6467];
assign t[6468] = t[6467] ^ n[6468];
assign t[6469] = t[6468] ^ n[6469];
assign t[6470] = t[6469] ^ n[6470];
assign t[6471] = t[6470] ^ n[6471];
assign t[6472] = t[6471] ^ n[6472];
assign t[6473] = t[6472] ^ n[6473];
assign t[6474] = t[6473] ^ n[6474];
assign t[6475] = t[6474] ^ n[6475];
assign t[6476] = t[6475] ^ n[6476];
assign t[6477] = t[6476] ^ n[6477];
assign t[6478] = t[6477] ^ n[6478];
assign t[6479] = t[6478] ^ n[6479];
assign t[6480] = t[6479] ^ n[6480];
assign t[6481] = t[6480] ^ n[6481];
assign t[6482] = t[6481] ^ n[6482];
assign t[6483] = t[6482] ^ n[6483];
assign t[6484] = t[6483] ^ n[6484];
assign t[6485] = t[6484] ^ n[6485];
assign t[6486] = t[6485] ^ n[6486];
assign t[6487] = t[6486] ^ n[6487];
assign t[6488] = t[6487] ^ n[6488];
assign t[6489] = t[6488] ^ n[6489];
assign t[6490] = t[6489] ^ n[6490];
assign t[6491] = t[6490] ^ n[6491];
assign t[6492] = t[6491] ^ n[6492];
assign t[6493] = t[6492] ^ n[6493];
assign t[6494] = t[6493] ^ n[6494];
assign t[6495] = t[6494] ^ n[6495];
assign t[6496] = t[6495] ^ n[6496];
assign t[6497] = t[6496] ^ n[6497];
assign t[6498] = t[6497] ^ n[6498];
assign t[6499] = t[6498] ^ n[6499];
assign t[6500] = t[6499] ^ n[6500];
assign t[6501] = t[6500] ^ n[6501];
assign t[6502] = t[6501] ^ n[6502];
assign t[6503] = t[6502] ^ n[6503];
assign t[6504] = t[6503] ^ n[6504];
assign t[6505] = t[6504] ^ n[6505];
assign t[6506] = t[6505] ^ n[6506];
assign t[6507] = t[6506] ^ n[6507];
assign t[6508] = t[6507] ^ n[6508];
assign t[6509] = t[6508] ^ n[6509];
assign t[6510] = t[6509] ^ n[6510];
assign t[6511] = t[6510] ^ n[6511];
assign t[6512] = t[6511] ^ n[6512];
assign t[6513] = t[6512] ^ n[6513];
assign t[6514] = t[6513] ^ n[6514];
assign t[6515] = t[6514] ^ n[6515];
assign t[6516] = t[6515] ^ n[6516];
assign t[6517] = t[6516] ^ n[6517];
assign t[6518] = t[6517] ^ n[6518];
assign t[6519] = t[6518] ^ n[6519];
assign t[6520] = t[6519] ^ n[6520];
assign t[6521] = t[6520] ^ n[6521];
assign t[6522] = t[6521] ^ n[6522];
assign t[6523] = t[6522] ^ n[6523];
assign t[6524] = t[6523] ^ n[6524];
assign t[6525] = t[6524] ^ n[6525];
assign t[6526] = t[6525] ^ n[6526];
assign t[6527] = t[6526] ^ n[6527];
assign t[6528] = t[6527] ^ n[6528];
assign t[6529] = t[6528] ^ n[6529];
assign t[6530] = t[6529] ^ n[6530];
assign t[6531] = t[6530] ^ n[6531];
assign t[6532] = t[6531] ^ n[6532];
assign t[6533] = t[6532] ^ n[6533];
assign t[6534] = t[6533] ^ n[6534];
assign t[6535] = t[6534] ^ n[6535];
assign t[6536] = t[6535] ^ n[6536];
assign t[6537] = t[6536] ^ n[6537];
assign t[6538] = t[6537] ^ n[6538];
assign t[6539] = t[6538] ^ n[6539];
assign t[6540] = t[6539] ^ n[6540];
assign t[6541] = t[6540] ^ n[6541];
assign t[6542] = t[6541] ^ n[6542];
assign t[6543] = t[6542] ^ n[6543];
assign t[6544] = t[6543] ^ n[6544];
assign t[6545] = t[6544] ^ n[6545];
assign t[6546] = t[6545] ^ n[6546];
assign t[6547] = t[6546] ^ n[6547];
assign t[6548] = t[6547] ^ n[6548];
assign t[6549] = t[6548] ^ n[6549];
assign t[6550] = t[6549] ^ n[6550];
assign t[6551] = t[6550] ^ n[6551];
assign t[6552] = t[6551] ^ n[6552];
assign t[6553] = t[6552] ^ n[6553];
assign t[6554] = t[6553] ^ n[6554];
assign t[6555] = t[6554] ^ n[6555];
assign t[6556] = t[6555] ^ n[6556];
assign t[6557] = t[6556] ^ n[6557];
assign t[6558] = t[6557] ^ n[6558];
assign t[6559] = t[6558] ^ n[6559];
assign t[6560] = t[6559] ^ n[6560];
assign t[6561] = t[6560] ^ n[6561];
assign t[6562] = t[6561] ^ n[6562];
assign t[6563] = t[6562] ^ n[6563];
assign t[6564] = t[6563] ^ n[6564];
assign t[6565] = t[6564] ^ n[6565];
assign t[6566] = t[6565] ^ n[6566];
assign t[6567] = t[6566] ^ n[6567];
assign t[6568] = t[6567] ^ n[6568];
assign t[6569] = t[6568] ^ n[6569];
assign t[6570] = t[6569] ^ n[6570];
assign t[6571] = t[6570] ^ n[6571];
assign t[6572] = t[6571] ^ n[6572];
assign t[6573] = t[6572] ^ n[6573];
assign t[6574] = t[6573] ^ n[6574];
assign t[6575] = t[6574] ^ n[6575];
assign t[6576] = t[6575] ^ n[6576];
assign t[6577] = t[6576] ^ n[6577];
assign t[6578] = t[6577] ^ n[6578];
assign t[6579] = t[6578] ^ n[6579];
assign t[6580] = t[6579] ^ n[6580];
assign t[6581] = t[6580] ^ n[6581];
assign t[6582] = t[6581] ^ n[6582];
assign t[6583] = t[6582] ^ n[6583];
assign t[6584] = t[6583] ^ n[6584];
assign t[6585] = t[6584] ^ n[6585];
assign t[6586] = t[6585] ^ n[6586];
assign t[6587] = t[6586] ^ n[6587];
assign t[6588] = t[6587] ^ n[6588];
assign t[6589] = t[6588] ^ n[6589];
assign t[6590] = t[6589] ^ n[6590];
assign t[6591] = t[6590] ^ n[6591];
assign t[6592] = t[6591] ^ n[6592];
assign t[6593] = t[6592] ^ n[6593];
assign t[6594] = t[6593] ^ n[6594];
assign t[6595] = t[6594] ^ n[6595];
assign t[6596] = t[6595] ^ n[6596];
assign t[6597] = t[6596] ^ n[6597];
assign t[6598] = t[6597] ^ n[6598];
assign t[6599] = t[6598] ^ n[6599];
assign t[6600] = t[6599] ^ n[6600];
assign t[6601] = t[6600] ^ n[6601];
assign t[6602] = t[6601] ^ n[6602];
assign t[6603] = t[6602] ^ n[6603];
assign t[6604] = t[6603] ^ n[6604];
assign t[6605] = t[6604] ^ n[6605];
assign t[6606] = t[6605] ^ n[6606];
assign t[6607] = t[6606] ^ n[6607];
assign t[6608] = t[6607] ^ n[6608];
assign t[6609] = t[6608] ^ n[6609];
assign t[6610] = t[6609] ^ n[6610];
assign t[6611] = t[6610] ^ n[6611];
assign t[6612] = t[6611] ^ n[6612];
assign t[6613] = t[6612] ^ n[6613];
assign t[6614] = t[6613] ^ n[6614];
assign t[6615] = t[6614] ^ n[6615];
assign t[6616] = t[6615] ^ n[6616];
assign t[6617] = t[6616] ^ n[6617];
assign t[6618] = t[6617] ^ n[6618];
assign t[6619] = t[6618] ^ n[6619];
assign t[6620] = t[6619] ^ n[6620];
assign t[6621] = t[6620] ^ n[6621];
assign t[6622] = t[6621] ^ n[6622];
assign t[6623] = t[6622] ^ n[6623];
assign t[6624] = t[6623] ^ n[6624];
assign t[6625] = t[6624] ^ n[6625];
assign t[6626] = t[6625] ^ n[6626];
assign t[6627] = t[6626] ^ n[6627];
assign t[6628] = t[6627] ^ n[6628];
assign t[6629] = t[6628] ^ n[6629];
assign t[6630] = t[6629] ^ n[6630];
assign t[6631] = t[6630] ^ n[6631];
assign t[6632] = t[6631] ^ n[6632];
assign t[6633] = t[6632] ^ n[6633];
assign t[6634] = t[6633] ^ n[6634];
assign t[6635] = t[6634] ^ n[6635];
assign t[6636] = t[6635] ^ n[6636];
assign t[6637] = t[6636] ^ n[6637];
assign t[6638] = t[6637] ^ n[6638];
assign t[6639] = t[6638] ^ n[6639];
assign t[6640] = t[6639] ^ n[6640];
assign t[6641] = t[6640] ^ n[6641];
assign t[6642] = t[6641] ^ n[6642];
assign t[6643] = t[6642] ^ n[6643];
assign t[6644] = t[6643] ^ n[6644];
assign t[6645] = t[6644] ^ n[6645];
assign t[6646] = t[6645] ^ n[6646];
assign t[6647] = t[6646] ^ n[6647];
assign t[6648] = t[6647] ^ n[6648];
assign t[6649] = t[6648] ^ n[6649];
assign t[6650] = t[6649] ^ n[6650];
assign t[6651] = t[6650] ^ n[6651];
assign t[6652] = t[6651] ^ n[6652];
assign t[6653] = t[6652] ^ n[6653];
assign t[6654] = t[6653] ^ n[6654];
assign t[6655] = t[6654] ^ n[6655];
assign t[6656] = t[6655] ^ n[6656];
assign t[6657] = t[6656] ^ n[6657];
assign t[6658] = t[6657] ^ n[6658];
assign t[6659] = t[6658] ^ n[6659];
assign t[6660] = t[6659] ^ n[6660];
assign t[6661] = t[6660] ^ n[6661];
assign t[6662] = t[6661] ^ n[6662];
assign t[6663] = t[6662] ^ n[6663];
assign t[6664] = t[6663] ^ n[6664];
assign t[6665] = t[6664] ^ n[6665];
assign t[6666] = t[6665] ^ n[6666];
assign t[6667] = t[6666] ^ n[6667];
assign t[6668] = t[6667] ^ n[6668];
assign t[6669] = t[6668] ^ n[6669];
assign t[6670] = t[6669] ^ n[6670];
assign t[6671] = t[6670] ^ n[6671];
assign t[6672] = t[6671] ^ n[6672];
assign t[6673] = t[6672] ^ n[6673];
assign t[6674] = t[6673] ^ n[6674];
assign t[6675] = t[6674] ^ n[6675];
assign t[6676] = t[6675] ^ n[6676];
assign t[6677] = t[6676] ^ n[6677];
assign t[6678] = t[6677] ^ n[6678];
assign t[6679] = t[6678] ^ n[6679];
assign t[6680] = t[6679] ^ n[6680];
assign t[6681] = t[6680] ^ n[6681];
assign t[6682] = t[6681] ^ n[6682];
assign t[6683] = t[6682] ^ n[6683];
assign t[6684] = t[6683] ^ n[6684];
assign t[6685] = t[6684] ^ n[6685];
assign t[6686] = t[6685] ^ n[6686];
assign t[6687] = t[6686] ^ n[6687];
assign t[6688] = t[6687] ^ n[6688];
assign t[6689] = t[6688] ^ n[6689];
assign t[6690] = t[6689] ^ n[6690];
assign t[6691] = t[6690] ^ n[6691];
assign t[6692] = t[6691] ^ n[6692];
assign t[6693] = t[6692] ^ n[6693];
assign t[6694] = t[6693] ^ n[6694];
assign t[6695] = t[6694] ^ n[6695];
assign t[6696] = t[6695] ^ n[6696];
assign t[6697] = t[6696] ^ n[6697];
assign t[6698] = t[6697] ^ n[6698];
assign t[6699] = t[6698] ^ n[6699];
assign t[6700] = t[6699] ^ n[6700];
assign t[6701] = t[6700] ^ n[6701];
assign t[6702] = t[6701] ^ n[6702];
assign t[6703] = t[6702] ^ n[6703];
assign t[6704] = t[6703] ^ n[6704];
assign t[6705] = t[6704] ^ n[6705];
assign t[6706] = t[6705] ^ n[6706];
assign t[6707] = t[6706] ^ n[6707];
assign t[6708] = t[6707] ^ n[6708];
assign t[6709] = t[6708] ^ n[6709];
assign t[6710] = t[6709] ^ n[6710];
assign t[6711] = t[6710] ^ n[6711];
assign t[6712] = t[6711] ^ n[6712];
assign t[6713] = t[6712] ^ n[6713];
assign t[6714] = t[6713] ^ n[6714];
assign t[6715] = t[6714] ^ n[6715];
assign t[6716] = t[6715] ^ n[6716];
assign t[6717] = t[6716] ^ n[6717];
assign t[6718] = t[6717] ^ n[6718];
assign t[6719] = t[6718] ^ n[6719];
assign t[6720] = t[6719] ^ n[6720];
assign t[6721] = t[6720] ^ n[6721];
assign t[6722] = t[6721] ^ n[6722];
assign t[6723] = t[6722] ^ n[6723];
assign t[6724] = t[6723] ^ n[6724];
assign t[6725] = t[6724] ^ n[6725];
assign t[6726] = t[6725] ^ n[6726];
assign t[6727] = t[6726] ^ n[6727];
assign t[6728] = t[6727] ^ n[6728];
assign t[6729] = t[6728] ^ n[6729];
assign t[6730] = t[6729] ^ n[6730];
assign t[6731] = t[6730] ^ n[6731];
assign t[6732] = t[6731] ^ n[6732];
assign t[6733] = t[6732] ^ n[6733];
assign t[6734] = t[6733] ^ n[6734];
assign t[6735] = t[6734] ^ n[6735];
assign t[6736] = t[6735] ^ n[6736];
assign t[6737] = t[6736] ^ n[6737];
assign t[6738] = t[6737] ^ n[6738];
assign t[6739] = t[6738] ^ n[6739];
assign t[6740] = t[6739] ^ n[6740];
assign t[6741] = t[6740] ^ n[6741];
assign t[6742] = t[6741] ^ n[6742];
assign t[6743] = t[6742] ^ n[6743];
assign t[6744] = t[6743] ^ n[6744];
assign t[6745] = t[6744] ^ n[6745];
assign t[6746] = t[6745] ^ n[6746];
assign t[6747] = t[6746] ^ n[6747];
assign t[6748] = t[6747] ^ n[6748];
assign t[6749] = t[6748] ^ n[6749];
assign t[6750] = t[6749] ^ n[6750];
assign t[6751] = t[6750] ^ n[6751];
assign t[6752] = t[6751] ^ n[6752];
assign t[6753] = t[6752] ^ n[6753];
assign t[6754] = t[6753] ^ n[6754];
assign t[6755] = t[6754] ^ n[6755];
assign t[6756] = t[6755] ^ n[6756];
assign t[6757] = t[6756] ^ n[6757];
assign t[6758] = t[6757] ^ n[6758];
assign t[6759] = t[6758] ^ n[6759];
assign t[6760] = t[6759] ^ n[6760];
assign t[6761] = t[6760] ^ n[6761];
assign t[6762] = t[6761] ^ n[6762];
assign t[6763] = t[6762] ^ n[6763];
assign t[6764] = t[6763] ^ n[6764];
assign t[6765] = t[6764] ^ n[6765];
assign t[6766] = t[6765] ^ n[6766];
assign t[6767] = t[6766] ^ n[6767];
assign t[6768] = t[6767] ^ n[6768];
assign t[6769] = t[6768] ^ n[6769];
assign t[6770] = t[6769] ^ n[6770];
assign t[6771] = t[6770] ^ n[6771];
assign t[6772] = t[6771] ^ n[6772];
assign t[6773] = t[6772] ^ n[6773];
assign t[6774] = t[6773] ^ n[6774];
assign t[6775] = t[6774] ^ n[6775];
assign t[6776] = t[6775] ^ n[6776];
assign t[6777] = t[6776] ^ n[6777];
assign t[6778] = t[6777] ^ n[6778];
assign t[6779] = t[6778] ^ n[6779];
assign t[6780] = t[6779] ^ n[6780];
assign t[6781] = t[6780] ^ n[6781];
assign t[6782] = t[6781] ^ n[6782];
assign t[6783] = t[6782] ^ n[6783];
assign t[6784] = t[6783] ^ n[6784];
assign t[6785] = t[6784] ^ n[6785];
assign t[6786] = t[6785] ^ n[6786];
assign t[6787] = t[6786] ^ n[6787];
assign t[6788] = t[6787] ^ n[6788];
assign t[6789] = t[6788] ^ n[6789];
assign t[6790] = t[6789] ^ n[6790];
assign t[6791] = t[6790] ^ n[6791];
assign t[6792] = t[6791] ^ n[6792];
assign t[6793] = t[6792] ^ n[6793];
assign t[6794] = t[6793] ^ n[6794];
assign t[6795] = t[6794] ^ n[6795];
assign t[6796] = t[6795] ^ n[6796];
assign t[6797] = t[6796] ^ n[6797];
assign t[6798] = t[6797] ^ n[6798];
assign t[6799] = t[6798] ^ n[6799];
assign t[6800] = t[6799] ^ n[6800];
assign t[6801] = t[6800] ^ n[6801];
assign t[6802] = t[6801] ^ n[6802];
assign t[6803] = t[6802] ^ n[6803];
assign t[6804] = t[6803] ^ n[6804];
assign t[6805] = t[6804] ^ n[6805];
assign t[6806] = t[6805] ^ n[6806];
assign t[6807] = t[6806] ^ n[6807];
assign t[6808] = t[6807] ^ n[6808];
assign t[6809] = t[6808] ^ n[6809];
assign t[6810] = t[6809] ^ n[6810];
assign t[6811] = t[6810] ^ n[6811];
assign t[6812] = t[6811] ^ n[6812];
assign t[6813] = t[6812] ^ n[6813];
assign t[6814] = t[6813] ^ n[6814];
assign t[6815] = t[6814] ^ n[6815];
assign t[6816] = t[6815] ^ n[6816];
assign t[6817] = t[6816] ^ n[6817];
assign t[6818] = t[6817] ^ n[6818];
assign t[6819] = t[6818] ^ n[6819];
assign t[6820] = t[6819] ^ n[6820];
assign t[6821] = t[6820] ^ n[6821];
assign t[6822] = t[6821] ^ n[6822];
assign t[6823] = t[6822] ^ n[6823];
assign t[6824] = t[6823] ^ n[6824];
assign t[6825] = t[6824] ^ n[6825];
assign t[6826] = t[6825] ^ n[6826];
assign t[6827] = t[6826] ^ n[6827];
assign t[6828] = t[6827] ^ n[6828];
assign t[6829] = t[6828] ^ n[6829];
assign t[6830] = t[6829] ^ n[6830];
assign t[6831] = t[6830] ^ n[6831];
assign t[6832] = t[6831] ^ n[6832];
assign t[6833] = t[6832] ^ n[6833];
assign t[6834] = t[6833] ^ n[6834];
assign t[6835] = t[6834] ^ n[6835];
assign t[6836] = t[6835] ^ n[6836];
assign t[6837] = t[6836] ^ n[6837];
assign t[6838] = t[6837] ^ n[6838];
assign t[6839] = t[6838] ^ n[6839];
assign t[6840] = t[6839] ^ n[6840];
assign t[6841] = t[6840] ^ n[6841];
assign t[6842] = t[6841] ^ n[6842];
assign t[6843] = t[6842] ^ n[6843];
assign t[6844] = t[6843] ^ n[6844];
assign t[6845] = t[6844] ^ n[6845];
assign t[6846] = t[6845] ^ n[6846];
assign t[6847] = t[6846] ^ n[6847];
assign t[6848] = t[6847] ^ n[6848];
assign t[6849] = t[6848] ^ n[6849];
assign t[6850] = t[6849] ^ n[6850];
assign t[6851] = t[6850] ^ n[6851];
assign t[6852] = t[6851] ^ n[6852];
assign t[6853] = t[6852] ^ n[6853];
assign t[6854] = t[6853] ^ n[6854];
assign t[6855] = t[6854] ^ n[6855];
assign t[6856] = t[6855] ^ n[6856];
assign t[6857] = t[6856] ^ n[6857];
assign t[6858] = t[6857] ^ n[6858];
assign t[6859] = t[6858] ^ n[6859];
assign t[6860] = t[6859] ^ n[6860];
assign t[6861] = t[6860] ^ n[6861];
assign t[6862] = t[6861] ^ n[6862];
assign t[6863] = t[6862] ^ n[6863];
assign t[6864] = t[6863] ^ n[6864];
assign t[6865] = t[6864] ^ n[6865];
assign t[6866] = t[6865] ^ n[6866];
assign t[6867] = t[6866] ^ n[6867];
assign t[6868] = t[6867] ^ n[6868];
assign t[6869] = t[6868] ^ n[6869];
assign t[6870] = t[6869] ^ n[6870];
assign t[6871] = t[6870] ^ n[6871];
assign t[6872] = t[6871] ^ n[6872];
assign t[6873] = t[6872] ^ n[6873];
assign t[6874] = t[6873] ^ n[6874];
assign t[6875] = t[6874] ^ n[6875];
assign t[6876] = t[6875] ^ n[6876];
assign t[6877] = t[6876] ^ n[6877];
assign t[6878] = t[6877] ^ n[6878];
assign t[6879] = t[6878] ^ n[6879];
assign t[6880] = t[6879] ^ n[6880];
assign t[6881] = t[6880] ^ n[6881];
assign t[6882] = t[6881] ^ n[6882];
assign t[6883] = t[6882] ^ n[6883];
assign t[6884] = t[6883] ^ n[6884];
assign t[6885] = t[6884] ^ n[6885];
assign t[6886] = t[6885] ^ n[6886];
assign t[6887] = t[6886] ^ n[6887];
assign t[6888] = t[6887] ^ n[6888];
assign t[6889] = t[6888] ^ n[6889];
assign t[6890] = t[6889] ^ n[6890];
assign t[6891] = t[6890] ^ n[6891];
assign t[6892] = t[6891] ^ n[6892];
assign t[6893] = t[6892] ^ n[6893];
assign t[6894] = t[6893] ^ n[6894];
assign t[6895] = t[6894] ^ n[6895];
assign t[6896] = t[6895] ^ n[6896];
assign t[6897] = t[6896] ^ n[6897];
assign t[6898] = t[6897] ^ n[6898];
assign t[6899] = t[6898] ^ n[6899];
assign t[6900] = t[6899] ^ n[6900];
assign t[6901] = t[6900] ^ n[6901];
assign t[6902] = t[6901] ^ n[6902];
assign t[6903] = t[6902] ^ n[6903];
assign t[6904] = t[6903] ^ n[6904];
assign t[6905] = t[6904] ^ n[6905];
assign t[6906] = t[6905] ^ n[6906];
assign t[6907] = t[6906] ^ n[6907];
assign t[6908] = t[6907] ^ n[6908];
assign t[6909] = t[6908] ^ n[6909];
assign t[6910] = t[6909] ^ n[6910];
assign t[6911] = t[6910] ^ n[6911];
assign t[6912] = t[6911] ^ n[6912];
assign t[6913] = t[6912] ^ n[6913];
assign t[6914] = t[6913] ^ n[6914];
assign t[6915] = t[6914] ^ n[6915];
assign t[6916] = t[6915] ^ n[6916];
assign t[6917] = t[6916] ^ n[6917];
assign t[6918] = t[6917] ^ n[6918];
assign t[6919] = t[6918] ^ n[6919];
assign t[6920] = t[6919] ^ n[6920];
assign t[6921] = t[6920] ^ n[6921];
assign t[6922] = t[6921] ^ n[6922];
assign t[6923] = t[6922] ^ n[6923];
assign t[6924] = t[6923] ^ n[6924];
assign t[6925] = t[6924] ^ n[6925];
assign t[6926] = t[6925] ^ n[6926];
assign t[6927] = t[6926] ^ n[6927];
assign t[6928] = t[6927] ^ n[6928];
assign t[6929] = t[6928] ^ n[6929];
assign t[6930] = t[6929] ^ n[6930];
assign t[6931] = t[6930] ^ n[6931];
assign t[6932] = t[6931] ^ n[6932];
assign t[6933] = t[6932] ^ n[6933];
assign t[6934] = t[6933] ^ n[6934];
assign t[6935] = t[6934] ^ n[6935];
assign t[6936] = t[6935] ^ n[6936];
assign t[6937] = t[6936] ^ n[6937];
assign t[6938] = t[6937] ^ n[6938];
assign t[6939] = t[6938] ^ n[6939];
assign t[6940] = t[6939] ^ n[6940];
assign t[6941] = t[6940] ^ n[6941];
assign t[6942] = t[6941] ^ n[6942];
assign t[6943] = t[6942] ^ n[6943];
assign t[6944] = t[6943] ^ n[6944];
assign t[6945] = t[6944] ^ n[6945];
assign t[6946] = t[6945] ^ n[6946];
assign t[6947] = t[6946] ^ n[6947];
assign t[6948] = t[6947] ^ n[6948];
assign t[6949] = t[6948] ^ n[6949];
assign t[6950] = t[6949] ^ n[6950];
assign t[6951] = t[6950] ^ n[6951];
assign t[6952] = t[6951] ^ n[6952];
assign t[6953] = t[6952] ^ n[6953];
assign t[6954] = t[6953] ^ n[6954];
assign t[6955] = t[6954] ^ n[6955];
assign t[6956] = t[6955] ^ n[6956];
assign t[6957] = t[6956] ^ n[6957];
assign t[6958] = t[6957] ^ n[6958];
assign t[6959] = t[6958] ^ n[6959];
assign t[6960] = t[6959] ^ n[6960];
assign t[6961] = t[6960] ^ n[6961];
assign t[6962] = t[6961] ^ n[6962];
assign t[6963] = t[6962] ^ n[6963];
assign t[6964] = t[6963] ^ n[6964];
assign t[6965] = t[6964] ^ n[6965];
assign t[6966] = t[6965] ^ n[6966];
assign t[6967] = t[6966] ^ n[6967];
assign t[6968] = t[6967] ^ n[6968];
assign t[6969] = t[6968] ^ n[6969];
assign t[6970] = t[6969] ^ n[6970];
assign t[6971] = t[6970] ^ n[6971];
assign t[6972] = t[6971] ^ n[6972];
assign t[6973] = t[6972] ^ n[6973];
assign t[6974] = t[6973] ^ n[6974];
assign t[6975] = t[6974] ^ n[6975];
assign t[6976] = t[6975] ^ n[6976];
assign t[6977] = t[6976] ^ n[6977];
assign t[6978] = t[6977] ^ n[6978];
assign t[6979] = t[6978] ^ n[6979];
assign t[6980] = t[6979] ^ n[6980];
assign t[6981] = t[6980] ^ n[6981];
assign t[6982] = t[6981] ^ n[6982];
assign t[6983] = t[6982] ^ n[6983];
assign t[6984] = t[6983] ^ n[6984];
assign t[6985] = t[6984] ^ n[6985];
assign t[6986] = t[6985] ^ n[6986];
assign t[6987] = t[6986] ^ n[6987];
assign t[6988] = t[6987] ^ n[6988];
assign t[6989] = t[6988] ^ n[6989];
assign t[6990] = t[6989] ^ n[6990];
assign t[6991] = t[6990] ^ n[6991];
assign t[6992] = t[6991] ^ n[6992];
assign t[6993] = t[6992] ^ n[6993];
assign t[6994] = t[6993] ^ n[6994];
assign t[6995] = t[6994] ^ n[6995];
assign t[6996] = t[6995] ^ n[6996];
assign t[6997] = t[6996] ^ n[6997];
assign t[6998] = t[6997] ^ n[6998];
assign t[6999] = t[6998] ^ n[6999];
assign t[7000] = t[6999] ^ n[7000];
assign t[7001] = t[7000] ^ n[7001];
assign t[7002] = t[7001] ^ n[7002];
assign t[7003] = t[7002] ^ n[7003];
assign t[7004] = t[7003] ^ n[7004];
assign t[7005] = t[7004] ^ n[7005];
assign t[7006] = t[7005] ^ n[7006];
assign t[7007] = t[7006] ^ n[7007];
assign t[7008] = t[7007] ^ n[7008];
assign t[7009] = t[7008] ^ n[7009];
assign t[7010] = t[7009] ^ n[7010];
assign t[7011] = t[7010] ^ n[7011];
assign t[7012] = t[7011] ^ n[7012];
assign t[7013] = t[7012] ^ n[7013];
assign t[7014] = t[7013] ^ n[7014];
assign t[7015] = t[7014] ^ n[7015];
assign t[7016] = t[7015] ^ n[7016];
assign t[7017] = t[7016] ^ n[7017];
assign t[7018] = t[7017] ^ n[7018];
assign t[7019] = t[7018] ^ n[7019];
assign t[7020] = t[7019] ^ n[7020];
assign t[7021] = t[7020] ^ n[7021];
assign t[7022] = t[7021] ^ n[7022];
assign t[7023] = t[7022] ^ n[7023];
assign t[7024] = t[7023] ^ n[7024];
assign t[7025] = t[7024] ^ n[7025];
assign t[7026] = t[7025] ^ n[7026];
assign t[7027] = t[7026] ^ n[7027];
assign t[7028] = t[7027] ^ n[7028];
assign t[7029] = t[7028] ^ n[7029];
assign t[7030] = t[7029] ^ n[7030];
assign t[7031] = t[7030] ^ n[7031];
assign t[7032] = t[7031] ^ n[7032];
assign t[7033] = t[7032] ^ n[7033];
assign t[7034] = t[7033] ^ n[7034];
assign t[7035] = t[7034] ^ n[7035];
assign t[7036] = t[7035] ^ n[7036];
assign t[7037] = t[7036] ^ n[7037];
assign t[7038] = t[7037] ^ n[7038];
assign t[7039] = t[7038] ^ n[7039];
assign t[7040] = t[7039] ^ n[7040];
assign t[7041] = t[7040] ^ n[7041];
assign t[7042] = t[7041] ^ n[7042];
assign t[7043] = t[7042] ^ n[7043];
assign t[7044] = t[7043] ^ n[7044];
assign t[7045] = t[7044] ^ n[7045];
assign t[7046] = t[7045] ^ n[7046];
assign t[7047] = t[7046] ^ n[7047];
assign t[7048] = t[7047] ^ n[7048];
assign t[7049] = t[7048] ^ n[7049];
assign t[7050] = t[7049] ^ n[7050];
assign t[7051] = t[7050] ^ n[7051];
assign t[7052] = t[7051] ^ n[7052];
assign t[7053] = t[7052] ^ n[7053];
assign t[7054] = t[7053] ^ n[7054];
assign t[7055] = t[7054] ^ n[7055];
assign t[7056] = t[7055] ^ n[7056];
assign t[7057] = t[7056] ^ n[7057];
assign t[7058] = t[7057] ^ n[7058];
assign t[7059] = t[7058] ^ n[7059];
assign t[7060] = t[7059] ^ n[7060];
assign t[7061] = t[7060] ^ n[7061];
assign t[7062] = t[7061] ^ n[7062];
assign t[7063] = t[7062] ^ n[7063];
assign t[7064] = t[7063] ^ n[7064];
assign t[7065] = t[7064] ^ n[7065];
assign t[7066] = t[7065] ^ n[7066];
assign t[7067] = t[7066] ^ n[7067];
assign t[7068] = t[7067] ^ n[7068];
assign t[7069] = t[7068] ^ n[7069];
assign t[7070] = t[7069] ^ n[7070];
assign t[7071] = t[7070] ^ n[7071];
assign t[7072] = t[7071] ^ n[7072];
assign t[7073] = t[7072] ^ n[7073];
assign t[7074] = t[7073] ^ n[7074];
assign t[7075] = t[7074] ^ n[7075];
assign t[7076] = t[7075] ^ n[7076];
assign t[7077] = t[7076] ^ n[7077];
assign t[7078] = t[7077] ^ n[7078];
assign t[7079] = t[7078] ^ n[7079];
assign t[7080] = t[7079] ^ n[7080];
assign t[7081] = t[7080] ^ n[7081];
assign t[7082] = t[7081] ^ n[7082];
assign t[7083] = t[7082] ^ n[7083];
assign t[7084] = t[7083] ^ n[7084];
assign t[7085] = t[7084] ^ n[7085];
assign t[7086] = t[7085] ^ n[7086];
assign t[7087] = t[7086] ^ n[7087];
assign t[7088] = t[7087] ^ n[7088];
assign t[7089] = t[7088] ^ n[7089];
assign t[7090] = t[7089] ^ n[7090];
assign t[7091] = t[7090] ^ n[7091];
assign t[7092] = t[7091] ^ n[7092];
assign t[7093] = t[7092] ^ n[7093];
assign t[7094] = t[7093] ^ n[7094];
assign t[7095] = t[7094] ^ n[7095];
assign t[7096] = t[7095] ^ n[7096];
assign t[7097] = t[7096] ^ n[7097];
assign t[7098] = t[7097] ^ n[7098];
assign t[7099] = t[7098] ^ n[7099];
assign t[7100] = t[7099] ^ n[7100];
assign t[7101] = t[7100] ^ n[7101];
assign t[7102] = t[7101] ^ n[7102];
assign t[7103] = t[7102] ^ n[7103];
assign t[7104] = t[7103] ^ n[7104];
assign t[7105] = t[7104] ^ n[7105];
assign t[7106] = t[7105] ^ n[7106];
assign t[7107] = t[7106] ^ n[7107];
assign t[7108] = t[7107] ^ n[7108];
assign t[7109] = t[7108] ^ n[7109];
assign t[7110] = t[7109] ^ n[7110];
assign t[7111] = t[7110] ^ n[7111];
assign t[7112] = t[7111] ^ n[7112];
assign t[7113] = t[7112] ^ n[7113];
assign t[7114] = t[7113] ^ n[7114];
assign t[7115] = t[7114] ^ n[7115];
assign t[7116] = t[7115] ^ n[7116];
assign t[7117] = t[7116] ^ n[7117];
assign t[7118] = t[7117] ^ n[7118];
assign t[7119] = t[7118] ^ n[7119];
assign t[7120] = t[7119] ^ n[7120];
assign t[7121] = t[7120] ^ n[7121];
assign t[7122] = t[7121] ^ n[7122];
assign t[7123] = t[7122] ^ n[7123];
assign t[7124] = t[7123] ^ n[7124];
assign t[7125] = t[7124] ^ n[7125];
assign t[7126] = t[7125] ^ n[7126];
assign t[7127] = t[7126] ^ n[7127];
assign t[7128] = t[7127] ^ n[7128];
assign t[7129] = t[7128] ^ n[7129];
assign t[7130] = t[7129] ^ n[7130];
assign t[7131] = t[7130] ^ n[7131];
assign t[7132] = t[7131] ^ n[7132];
assign t[7133] = t[7132] ^ n[7133];
assign t[7134] = t[7133] ^ n[7134];
assign t[7135] = t[7134] ^ n[7135];
assign t[7136] = t[7135] ^ n[7136];
assign t[7137] = t[7136] ^ n[7137];
assign t[7138] = t[7137] ^ n[7138];
assign t[7139] = t[7138] ^ n[7139];
assign t[7140] = t[7139] ^ n[7140];
assign t[7141] = t[7140] ^ n[7141];
assign t[7142] = t[7141] ^ n[7142];
assign t[7143] = t[7142] ^ n[7143];
assign t[7144] = t[7143] ^ n[7144];
assign t[7145] = t[7144] ^ n[7145];
assign t[7146] = t[7145] ^ n[7146];
assign t[7147] = t[7146] ^ n[7147];
assign t[7148] = t[7147] ^ n[7148];
assign t[7149] = t[7148] ^ n[7149];
assign t[7150] = t[7149] ^ n[7150];
assign t[7151] = t[7150] ^ n[7151];
assign t[7152] = t[7151] ^ n[7152];
assign t[7153] = t[7152] ^ n[7153];
assign t[7154] = t[7153] ^ n[7154];
assign t[7155] = t[7154] ^ n[7155];
assign t[7156] = t[7155] ^ n[7156];
assign t[7157] = t[7156] ^ n[7157];
assign t[7158] = t[7157] ^ n[7158];
assign t[7159] = t[7158] ^ n[7159];
assign t[7160] = t[7159] ^ n[7160];
assign t[7161] = t[7160] ^ n[7161];
assign t[7162] = t[7161] ^ n[7162];
assign t[7163] = t[7162] ^ n[7163];
assign t[7164] = t[7163] ^ n[7164];
assign t[7165] = t[7164] ^ n[7165];
assign t[7166] = t[7165] ^ n[7166];
assign t[7167] = t[7166] ^ n[7167];
assign t[7168] = t[7167] ^ n[7168];
assign t[7169] = t[7168] ^ n[7169];
assign t[7170] = t[7169] ^ n[7170];
assign t[7171] = t[7170] ^ n[7171];
assign t[7172] = t[7171] ^ n[7172];
assign t[7173] = t[7172] ^ n[7173];
assign t[7174] = t[7173] ^ n[7174];
assign t[7175] = t[7174] ^ n[7175];
assign t[7176] = t[7175] ^ n[7176];
assign t[7177] = t[7176] ^ n[7177];
assign t[7178] = t[7177] ^ n[7178];
assign t[7179] = t[7178] ^ n[7179];
assign t[7180] = t[7179] ^ n[7180];
assign t[7181] = t[7180] ^ n[7181];
assign t[7182] = t[7181] ^ n[7182];
assign t[7183] = t[7182] ^ n[7183];
assign t[7184] = t[7183] ^ n[7184];
assign t[7185] = t[7184] ^ n[7185];
assign t[7186] = t[7185] ^ n[7186];
assign t[7187] = t[7186] ^ n[7187];
assign t[7188] = t[7187] ^ n[7188];
assign t[7189] = t[7188] ^ n[7189];
assign t[7190] = t[7189] ^ n[7190];
assign t[7191] = t[7190] ^ n[7191];
assign t[7192] = t[7191] ^ n[7192];
assign t[7193] = t[7192] ^ n[7193];
assign t[7194] = t[7193] ^ n[7194];
assign t[7195] = t[7194] ^ n[7195];
assign t[7196] = t[7195] ^ n[7196];
assign t[7197] = t[7196] ^ n[7197];
assign t[7198] = t[7197] ^ n[7198];
assign t[7199] = t[7198] ^ n[7199];
assign t[7200] = t[7199] ^ n[7200];
assign t[7201] = t[7200] ^ n[7201];
assign t[7202] = t[7201] ^ n[7202];
assign t[7203] = t[7202] ^ n[7203];
assign t[7204] = t[7203] ^ n[7204];
assign t[7205] = t[7204] ^ n[7205];
assign t[7206] = t[7205] ^ n[7206];
assign t[7207] = t[7206] ^ n[7207];
assign t[7208] = t[7207] ^ n[7208];
assign t[7209] = t[7208] ^ n[7209];
assign t[7210] = t[7209] ^ n[7210];
assign t[7211] = t[7210] ^ n[7211];
assign t[7212] = t[7211] ^ n[7212];
assign t[7213] = t[7212] ^ n[7213];
assign t[7214] = t[7213] ^ n[7214];
assign t[7215] = t[7214] ^ n[7215];
assign t[7216] = t[7215] ^ n[7216];
assign t[7217] = t[7216] ^ n[7217];
assign t[7218] = t[7217] ^ n[7218];
assign t[7219] = t[7218] ^ n[7219];
assign t[7220] = t[7219] ^ n[7220];
assign t[7221] = t[7220] ^ n[7221];
assign t[7222] = t[7221] ^ n[7222];
assign t[7223] = t[7222] ^ n[7223];
assign t[7224] = t[7223] ^ n[7224];
assign t[7225] = t[7224] ^ n[7225];
assign t[7226] = t[7225] ^ n[7226];
assign t[7227] = t[7226] ^ n[7227];
assign t[7228] = t[7227] ^ n[7228];
assign t[7229] = t[7228] ^ n[7229];
assign t[7230] = t[7229] ^ n[7230];
assign t[7231] = t[7230] ^ n[7231];
assign t[7232] = t[7231] ^ n[7232];
assign t[7233] = t[7232] ^ n[7233];
assign t[7234] = t[7233] ^ n[7234];
assign t[7235] = t[7234] ^ n[7235];
assign t[7236] = t[7235] ^ n[7236];
assign t[7237] = t[7236] ^ n[7237];
assign t[7238] = t[7237] ^ n[7238];
assign t[7239] = t[7238] ^ n[7239];
assign t[7240] = t[7239] ^ n[7240];
assign t[7241] = t[7240] ^ n[7241];
assign t[7242] = t[7241] ^ n[7242];
assign t[7243] = t[7242] ^ n[7243];
assign t[7244] = t[7243] ^ n[7244];
assign t[7245] = t[7244] ^ n[7245];
assign t[7246] = t[7245] ^ n[7246];
assign t[7247] = t[7246] ^ n[7247];
assign t[7248] = t[7247] ^ n[7248];
assign t[7249] = t[7248] ^ n[7249];
assign t[7250] = t[7249] ^ n[7250];
assign t[7251] = t[7250] ^ n[7251];
assign t[7252] = t[7251] ^ n[7252];
assign t[7253] = t[7252] ^ n[7253];
assign t[7254] = t[7253] ^ n[7254];
assign t[7255] = t[7254] ^ n[7255];
assign t[7256] = t[7255] ^ n[7256];
assign t[7257] = t[7256] ^ n[7257];
assign t[7258] = t[7257] ^ n[7258];
assign t[7259] = t[7258] ^ n[7259];
assign t[7260] = t[7259] ^ n[7260];
assign t[7261] = t[7260] ^ n[7261];
assign t[7262] = t[7261] ^ n[7262];
assign t[7263] = t[7262] ^ n[7263];
assign t[7264] = t[7263] ^ n[7264];
assign t[7265] = t[7264] ^ n[7265];
assign t[7266] = t[7265] ^ n[7266];
assign t[7267] = t[7266] ^ n[7267];
assign t[7268] = t[7267] ^ n[7268];
assign t[7269] = t[7268] ^ n[7269];
assign t[7270] = t[7269] ^ n[7270];
assign t[7271] = t[7270] ^ n[7271];
assign t[7272] = t[7271] ^ n[7272];
assign t[7273] = t[7272] ^ n[7273];
assign t[7274] = t[7273] ^ n[7274];
assign t[7275] = t[7274] ^ n[7275];
assign t[7276] = t[7275] ^ n[7276];
assign t[7277] = t[7276] ^ n[7277];
assign t[7278] = t[7277] ^ n[7278];
assign t[7279] = t[7278] ^ n[7279];
assign t[7280] = t[7279] ^ n[7280];
assign t[7281] = t[7280] ^ n[7281];
assign t[7282] = t[7281] ^ n[7282];
assign t[7283] = t[7282] ^ n[7283];
assign t[7284] = t[7283] ^ n[7284];
assign t[7285] = t[7284] ^ n[7285];
assign t[7286] = t[7285] ^ n[7286];
assign t[7287] = t[7286] ^ n[7287];
assign t[7288] = t[7287] ^ n[7288];
assign t[7289] = t[7288] ^ n[7289];
assign t[7290] = t[7289] ^ n[7290];
assign t[7291] = t[7290] ^ n[7291];
assign t[7292] = t[7291] ^ n[7292];
assign t[7293] = t[7292] ^ n[7293];
assign t[7294] = t[7293] ^ n[7294];
assign t[7295] = t[7294] ^ n[7295];
assign t[7296] = t[7295] ^ n[7296];
assign t[7297] = t[7296] ^ n[7297];
assign t[7298] = t[7297] ^ n[7298];
assign t[7299] = t[7298] ^ n[7299];
assign t[7300] = t[7299] ^ n[7300];
assign t[7301] = t[7300] ^ n[7301];
assign t[7302] = t[7301] ^ n[7302];
assign t[7303] = t[7302] ^ n[7303];
assign t[7304] = t[7303] ^ n[7304];
assign t[7305] = t[7304] ^ n[7305];
assign t[7306] = t[7305] ^ n[7306];
assign t[7307] = t[7306] ^ n[7307];
assign t[7308] = t[7307] ^ n[7308];
assign t[7309] = t[7308] ^ n[7309];
assign t[7310] = t[7309] ^ n[7310];
assign t[7311] = t[7310] ^ n[7311];
assign t[7312] = t[7311] ^ n[7312];
assign t[7313] = t[7312] ^ n[7313];
assign t[7314] = t[7313] ^ n[7314];
assign t[7315] = t[7314] ^ n[7315];
assign t[7316] = t[7315] ^ n[7316];
assign t[7317] = t[7316] ^ n[7317];
assign t[7318] = t[7317] ^ n[7318];
assign t[7319] = t[7318] ^ n[7319];
assign t[7320] = t[7319] ^ n[7320];
assign t[7321] = t[7320] ^ n[7321];
assign t[7322] = t[7321] ^ n[7322];
assign t[7323] = t[7322] ^ n[7323];
assign t[7324] = t[7323] ^ n[7324];
assign t[7325] = t[7324] ^ n[7325];
assign t[7326] = t[7325] ^ n[7326];
assign t[7327] = t[7326] ^ n[7327];
assign t[7328] = t[7327] ^ n[7328];
assign t[7329] = t[7328] ^ n[7329];
assign t[7330] = t[7329] ^ n[7330];
assign t[7331] = t[7330] ^ n[7331];
assign t[7332] = t[7331] ^ n[7332];
assign t[7333] = t[7332] ^ n[7333];
assign t[7334] = t[7333] ^ n[7334];
assign t[7335] = t[7334] ^ n[7335];
assign t[7336] = t[7335] ^ n[7336];
assign t[7337] = t[7336] ^ n[7337];
assign t[7338] = t[7337] ^ n[7338];
assign t[7339] = t[7338] ^ n[7339];
assign t[7340] = t[7339] ^ n[7340];
assign t[7341] = t[7340] ^ n[7341];
assign t[7342] = t[7341] ^ n[7342];
assign t[7343] = t[7342] ^ n[7343];
assign t[7344] = t[7343] ^ n[7344];
assign t[7345] = t[7344] ^ n[7345];
assign t[7346] = t[7345] ^ n[7346];
assign t[7347] = t[7346] ^ n[7347];
assign t[7348] = t[7347] ^ n[7348];
assign t[7349] = t[7348] ^ n[7349];
assign t[7350] = t[7349] ^ n[7350];
assign t[7351] = t[7350] ^ n[7351];
assign t[7352] = t[7351] ^ n[7352];
assign t[7353] = t[7352] ^ n[7353];
assign t[7354] = t[7353] ^ n[7354];
assign t[7355] = t[7354] ^ n[7355];
assign t[7356] = t[7355] ^ n[7356];
assign t[7357] = t[7356] ^ n[7357];
assign t[7358] = t[7357] ^ n[7358];
assign t[7359] = t[7358] ^ n[7359];
assign t[7360] = t[7359] ^ n[7360];
assign t[7361] = t[7360] ^ n[7361];
assign t[7362] = t[7361] ^ n[7362];
assign t[7363] = t[7362] ^ n[7363];
assign t[7364] = t[7363] ^ n[7364];
assign t[7365] = t[7364] ^ n[7365];
assign t[7366] = t[7365] ^ n[7366];
assign t[7367] = t[7366] ^ n[7367];
assign t[7368] = t[7367] ^ n[7368];
assign t[7369] = t[7368] ^ n[7369];
assign t[7370] = t[7369] ^ n[7370];
assign t[7371] = t[7370] ^ n[7371];
assign t[7372] = t[7371] ^ n[7372];
assign t[7373] = t[7372] ^ n[7373];
assign t[7374] = t[7373] ^ n[7374];
assign t[7375] = t[7374] ^ n[7375];
assign t[7376] = t[7375] ^ n[7376];
assign t[7377] = t[7376] ^ n[7377];
assign t[7378] = t[7377] ^ n[7378];
assign t[7379] = t[7378] ^ n[7379];
assign t[7380] = t[7379] ^ n[7380];
assign t[7381] = t[7380] ^ n[7381];
assign t[7382] = t[7381] ^ n[7382];
assign t[7383] = t[7382] ^ n[7383];
assign t[7384] = t[7383] ^ n[7384];
assign t[7385] = t[7384] ^ n[7385];
assign t[7386] = t[7385] ^ n[7386];
assign t[7387] = t[7386] ^ n[7387];
assign t[7388] = t[7387] ^ n[7388];
assign t[7389] = t[7388] ^ n[7389];
assign t[7390] = t[7389] ^ n[7390];
assign t[7391] = t[7390] ^ n[7391];
assign t[7392] = t[7391] ^ n[7392];
assign t[7393] = t[7392] ^ n[7393];
assign t[7394] = t[7393] ^ n[7394];
assign t[7395] = t[7394] ^ n[7395];
assign t[7396] = t[7395] ^ n[7396];
assign t[7397] = t[7396] ^ n[7397];
assign t[7398] = t[7397] ^ n[7398];
assign t[7399] = t[7398] ^ n[7399];
assign t[7400] = t[7399] ^ n[7400];
assign t[7401] = t[7400] ^ n[7401];
assign t[7402] = t[7401] ^ n[7402];
assign t[7403] = t[7402] ^ n[7403];
assign t[7404] = t[7403] ^ n[7404];
assign t[7405] = t[7404] ^ n[7405];
assign t[7406] = t[7405] ^ n[7406];
assign t[7407] = t[7406] ^ n[7407];
assign t[7408] = t[7407] ^ n[7408];
assign t[7409] = t[7408] ^ n[7409];
assign t[7410] = t[7409] ^ n[7410];
assign t[7411] = t[7410] ^ n[7411];
assign t[7412] = t[7411] ^ n[7412];
assign t[7413] = t[7412] ^ n[7413];
assign t[7414] = t[7413] ^ n[7414];
assign t[7415] = t[7414] ^ n[7415];
assign t[7416] = t[7415] ^ n[7416];
assign t[7417] = t[7416] ^ n[7417];
assign t[7418] = t[7417] ^ n[7418];
assign t[7419] = t[7418] ^ n[7419];
assign t[7420] = t[7419] ^ n[7420];
assign t[7421] = t[7420] ^ n[7421];
assign t[7422] = t[7421] ^ n[7422];
assign t[7423] = t[7422] ^ n[7423];
assign t[7424] = t[7423] ^ n[7424];
assign t[7425] = t[7424] ^ n[7425];
assign t[7426] = t[7425] ^ n[7426];
assign t[7427] = t[7426] ^ n[7427];
assign t[7428] = t[7427] ^ n[7428];
assign t[7429] = t[7428] ^ n[7429];
assign t[7430] = t[7429] ^ n[7430];
assign t[7431] = t[7430] ^ n[7431];
assign t[7432] = t[7431] ^ n[7432];
assign t[7433] = t[7432] ^ n[7433];
assign t[7434] = t[7433] ^ n[7434];
assign t[7435] = t[7434] ^ n[7435];
assign t[7436] = t[7435] ^ n[7436];
assign t[7437] = t[7436] ^ n[7437];
assign t[7438] = t[7437] ^ n[7438];
assign t[7439] = t[7438] ^ n[7439];
assign t[7440] = t[7439] ^ n[7440];
assign t[7441] = t[7440] ^ n[7441];
assign t[7442] = t[7441] ^ n[7442];
assign t[7443] = t[7442] ^ n[7443];
assign t[7444] = t[7443] ^ n[7444];
assign t[7445] = t[7444] ^ n[7445];
assign t[7446] = t[7445] ^ n[7446];
assign t[7447] = t[7446] ^ n[7447];
assign t[7448] = t[7447] ^ n[7448];
assign t[7449] = t[7448] ^ n[7449];
assign t[7450] = t[7449] ^ n[7450];
assign t[7451] = t[7450] ^ n[7451];
assign t[7452] = t[7451] ^ n[7452];
assign t[7453] = t[7452] ^ n[7453];
assign t[7454] = t[7453] ^ n[7454];
assign t[7455] = t[7454] ^ n[7455];
assign t[7456] = t[7455] ^ n[7456];
assign t[7457] = t[7456] ^ n[7457];
assign t[7458] = t[7457] ^ n[7458];
assign t[7459] = t[7458] ^ n[7459];
assign t[7460] = t[7459] ^ n[7460];
assign t[7461] = t[7460] ^ n[7461];
assign t[7462] = t[7461] ^ n[7462];
assign t[7463] = t[7462] ^ n[7463];
assign t[7464] = t[7463] ^ n[7464];
assign t[7465] = t[7464] ^ n[7465];
assign t[7466] = t[7465] ^ n[7466];
assign t[7467] = t[7466] ^ n[7467];
assign t[7468] = t[7467] ^ n[7468];
assign t[7469] = t[7468] ^ n[7469];
assign t[7470] = t[7469] ^ n[7470];
assign t[7471] = t[7470] ^ n[7471];
assign t[7472] = t[7471] ^ n[7472];
assign t[7473] = t[7472] ^ n[7473];
assign t[7474] = t[7473] ^ n[7474];
assign t[7475] = t[7474] ^ n[7475];
assign t[7476] = t[7475] ^ n[7476];
assign t[7477] = t[7476] ^ n[7477];
assign t[7478] = t[7477] ^ n[7478];
assign t[7479] = t[7478] ^ n[7479];
assign t[7480] = t[7479] ^ n[7480];
assign t[7481] = t[7480] ^ n[7481];
assign t[7482] = t[7481] ^ n[7482];
assign t[7483] = t[7482] ^ n[7483];
assign t[7484] = t[7483] ^ n[7484];
assign t[7485] = t[7484] ^ n[7485];
assign t[7486] = t[7485] ^ n[7486];
assign t[7487] = t[7486] ^ n[7487];
assign t[7488] = t[7487] ^ n[7488];
assign t[7489] = t[7488] ^ n[7489];
assign t[7490] = t[7489] ^ n[7490];
assign t[7491] = t[7490] ^ n[7491];
assign t[7492] = t[7491] ^ n[7492];
assign t[7493] = t[7492] ^ n[7493];
assign t[7494] = t[7493] ^ n[7494];
assign t[7495] = t[7494] ^ n[7495];
assign t[7496] = t[7495] ^ n[7496];
assign t[7497] = t[7496] ^ n[7497];
assign t[7498] = t[7497] ^ n[7498];
assign t[7499] = t[7498] ^ n[7499];
assign t[7500] = t[7499] ^ n[7500];
assign t[7501] = t[7500] ^ n[7501];
assign t[7502] = t[7501] ^ n[7502];
assign t[7503] = t[7502] ^ n[7503];
assign t[7504] = t[7503] ^ n[7504];
assign t[7505] = t[7504] ^ n[7505];
assign t[7506] = t[7505] ^ n[7506];
assign t[7507] = t[7506] ^ n[7507];
assign t[7508] = t[7507] ^ n[7508];
assign t[7509] = t[7508] ^ n[7509];
assign t[7510] = t[7509] ^ n[7510];
assign t[7511] = t[7510] ^ n[7511];
assign t[7512] = t[7511] ^ n[7512];
assign t[7513] = t[7512] ^ n[7513];
assign t[7514] = t[7513] ^ n[7514];
assign t[7515] = t[7514] ^ n[7515];
assign t[7516] = t[7515] ^ n[7516];
assign t[7517] = t[7516] ^ n[7517];
assign t[7518] = t[7517] ^ n[7518];
assign t[7519] = t[7518] ^ n[7519];
assign t[7520] = t[7519] ^ n[7520];
assign t[7521] = t[7520] ^ n[7521];
assign t[7522] = t[7521] ^ n[7522];
assign t[7523] = t[7522] ^ n[7523];
assign t[7524] = t[7523] ^ n[7524];
assign t[7525] = t[7524] ^ n[7525];
assign t[7526] = t[7525] ^ n[7526];
assign t[7527] = t[7526] ^ n[7527];
assign t[7528] = t[7527] ^ n[7528];
assign t[7529] = t[7528] ^ n[7529];
assign t[7530] = t[7529] ^ n[7530];
assign t[7531] = t[7530] ^ n[7531];
assign t[7532] = t[7531] ^ n[7532];
assign t[7533] = t[7532] ^ n[7533];
assign t[7534] = t[7533] ^ n[7534];
assign t[7535] = t[7534] ^ n[7535];
assign t[7536] = t[7535] ^ n[7536];
assign t[7537] = t[7536] ^ n[7537];
assign t[7538] = t[7537] ^ n[7538];
assign t[7539] = t[7538] ^ n[7539];
assign t[7540] = t[7539] ^ n[7540];
assign t[7541] = t[7540] ^ n[7541];
assign t[7542] = t[7541] ^ n[7542];
assign t[7543] = t[7542] ^ n[7543];
assign t[7544] = t[7543] ^ n[7544];
assign t[7545] = t[7544] ^ n[7545];
assign t[7546] = t[7545] ^ n[7546];
assign t[7547] = t[7546] ^ n[7547];
assign t[7548] = t[7547] ^ n[7548];
assign t[7549] = t[7548] ^ n[7549];
assign t[7550] = t[7549] ^ n[7550];
assign t[7551] = t[7550] ^ n[7551];
assign t[7552] = t[7551] ^ n[7552];
assign t[7553] = t[7552] ^ n[7553];
assign t[7554] = t[7553] ^ n[7554];
assign t[7555] = t[7554] ^ n[7555];
assign t[7556] = t[7555] ^ n[7556];
assign t[7557] = t[7556] ^ n[7557];
assign t[7558] = t[7557] ^ n[7558];
assign t[7559] = t[7558] ^ n[7559];
assign t[7560] = t[7559] ^ n[7560];
assign t[7561] = t[7560] ^ n[7561];
assign t[7562] = t[7561] ^ n[7562];
assign t[7563] = t[7562] ^ n[7563];
assign t[7564] = t[7563] ^ n[7564];
assign t[7565] = t[7564] ^ n[7565];
assign t[7566] = t[7565] ^ n[7566];
assign t[7567] = t[7566] ^ n[7567];
assign t[7568] = t[7567] ^ n[7568];
assign t[7569] = t[7568] ^ n[7569];
assign t[7570] = t[7569] ^ n[7570];
assign t[7571] = t[7570] ^ n[7571];
assign t[7572] = t[7571] ^ n[7572];
assign t[7573] = t[7572] ^ n[7573];
assign t[7574] = t[7573] ^ n[7574];
assign t[7575] = t[7574] ^ n[7575];
assign t[7576] = t[7575] ^ n[7576];
assign t[7577] = t[7576] ^ n[7577];
assign t[7578] = t[7577] ^ n[7578];
assign t[7579] = t[7578] ^ n[7579];
assign t[7580] = t[7579] ^ n[7580];
assign t[7581] = t[7580] ^ n[7581];
assign t[7582] = t[7581] ^ n[7582];
assign t[7583] = t[7582] ^ n[7583];
assign t[7584] = t[7583] ^ n[7584];
assign t[7585] = t[7584] ^ n[7585];
assign t[7586] = t[7585] ^ n[7586];
assign t[7587] = t[7586] ^ n[7587];
assign t[7588] = t[7587] ^ n[7588];
assign t[7589] = t[7588] ^ n[7589];
assign t[7590] = t[7589] ^ n[7590];
assign t[7591] = t[7590] ^ n[7591];
assign t[7592] = t[7591] ^ n[7592];
assign t[7593] = t[7592] ^ n[7593];
assign t[7594] = t[7593] ^ n[7594];
assign t[7595] = t[7594] ^ n[7595];
assign t[7596] = t[7595] ^ n[7596];
assign t[7597] = t[7596] ^ n[7597];
assign t[7598] = t[7597] ^ n[7598];
assign t[7599] = t[7598] ^ n[7599];
assign t[7600] = t[7599] ^ n[7600];
assign t[7601] = t[7600] ^ n[7601];
assign t[7602] = t[7601] ^ n[7602];
assign t[7603] = t[7602] ^ n[7603];
assign t[7604] = t[7603] ^ n[7604];
assign t[7605] = t[7604] ^ n[7605];
assign t[7606] = t[7605] ^ n[7606];
assign t[7607] = t[7606] ^ n[7607];
assign t[7608] = t[7607] ^ n[7608];
assign t[7609] = t[7608] ^ n[7609];
assign t[7610] = t[7609] ^ n[7610];
assign t[7611] = t[7610] ^ n[7611];
assign t[7612] = t[7611] ^ n[7612];
assign t[7613] = t[7612] ^ n[7613];
assign t[7614] = t[7613] ^ n[7614];
assign t[7615] = t[7614] ^ n[7615];
assign t[7616] = t[7615] ^ n[7616];
assign t[7617] = t[7616] ^ n[7617];
assign t[7618] = t[7617] ^ n[7618];
assign t[7619] = t[7618] ^ n[7619];
assign t[7620] = t[7619] ^ n[7620];
assign t[7621] = t[7620] ^ n[7621];
assign t[7622] = t[7621] ^ n[7622];
assign t[7623] = t[7622] ^ n[7623];
assign t[7624] = t[7623] ^ n[7624];
assign t[7625] = t[7624] ^ n[7625];
assign t[7626] = t[7625] ^ n[7626];
assign t[7627] = t[7626] ^ n[7627];
assign t[7628] = t[7627] ^ n[7628];
assign t[7629] = t[7628] ^ n[7629];
assign t[7630] = t[7629] ^ n[7630];
assign t[7631] = t[7630] ^ n[7631];
assign t[7632] = t[7631] ^ n[7632];
assign t[7633] = t[7632] ^ n[7633];
assign t[7634] = t[7633] ^ n[7634];
assign t[7635] = t[7634] ^ n[7635];
assign t[7636] = t[7635] ^ n[7636];
assign t[7637] = t[7636] ^ n[7637];
assign t[7638] = t[7637] ^ n[7638];
assign t[7639] = t[7638] ^ n[7639];
assign t[7640] = t[7639] ^ n[7640];
assign t[7641] = t[7640] ^ n[7641];
assign t[7642] = t[7641] ^ n[7642];
assign t[7643] = t[7642] ^ n[7643];
assign t[7644] = t[7643] ^ n[7644];
assign t[7645] = t[7644] ^ n[7645];
assign t[7646] = t[7645] ^ n[7646];
assign t[7647] = t[7646] ^ n[7647];
assign t[7648] = t[7647] ^ n[7648];
assign t[7649] = t[7648] ^ n[7649];
assign t[7650] = t[7649] ^ n[7650];
assign t[7651] = t[7650] ^ n[7651];
assign t[7652] = t[7651] ^ n[7652];
assign t[7653] = t[7652] ^ n[7653];
assign t[7654] = t[7653] ^ n[7654];
assign t[7655] = t[7654] ^ n[7655];
assign t[7656] = t[7655] ^ n[7656];
assign t[7657] = t[7656] ^ n[7657];
assign t[7658] = t[7657] ^ n[7658];
assign t[7659] = t[7658] ^ n[7659];
assign t[7660] = t[7659] ^ n[7660];
assign t[7661] = t[7660] ^ n[7661];
assign t[7662] = t[7661] ^ n[7662];
assign t[7663] = t[7662] ^ n[7663];
assign t[7664] = t[7663] ^ n[7664];
assign t[7665] = t[7664] ^ n[7665];
assign t[7666] = t[7665] ^ n[7666];
assign t[7667] = t[7666] ^ n[7667];
assign t[7668] = t[7667] ^ n[7668];
assign t[7669] = t[7668] ^ n[7669];
assign t[7670] = t[7669] ^ n[7670];
assign t[7671] = t[7670] ^ n[7671];
assign t[7672] = t[7671] ^ n[7672];
assign t[7673] = t[7672] ^ n[7673];
assign t[7674] = t[7673] ^ n[7674];
assign t[7675] = t[7674] ^ n[7675];
assign t[7676] = t[7675] ^ n[7676];
assign t[7677] = t[7676] ^ n[7677];
assign t[7678] = t[7677] ^ n[7678];
assign t[7679] = t[7678] ^ n[7679];
assign t[7680] = t[7679] ^ n[7680];
assign t[7681] = t[7680] ^ n[7681];
assign t[7682] = t[7681] ^ n[7682];
assign t[7683] = t[7682] ^ n[7683];
assign t[7684] = t[7683] ^ n[7684];
assign t[7685] = t[7684] ^ n[7685];
assign t[7686] = t[7685] ^ n[7686];
assign t[7687] = t[7686] ^ n[7687];
assign t[7688] = t[7687] ^ n[7688];
assign t[7689] = t[7688] ^ n[7689];
assign t[7690] = t[7689] ^ n[7690];
assign t[7691] = t[7690] ^ n[7691];
assign t[7692] = t[7691] ^ n[7692];
assign t[7693] = t[7692] ^ n[7693];
assign t[7694] = t[7693] ^ n[7694];
assign t[7695] = t[7694] ^ n[7695];
assign t[7696] = t[7695] ^ n[7696];
assign t[7697] = t[7696] ^ n[7697];
assign t[7698] = t[7697] ^ n[7698];
assign t[7699] = t[7698] ^ n[7699];
assign t[7700] = t[7699] ^ n[7700];
assign t[7701] = t[7700] ^ n[7701];
assign t[7702] = t[7701] ^ n[7702];
assign t[7703] = t[7702] ^ n[7703];
assign t[7704] = t[7703] ^ n[7704];
assign t[7705] = t[7704] ^ n[7705];
assign t[7706] = t[7705] ^ n[7706];
assign t[7707] = t[7706] ^ n[7707];
assign t[7708] = t[7707] ^ n[7708];
assign t[7709] = t[7708] ^ n[7709];
assign t[7710] = t[7709] ^ n[7710];
assign t[7711] = t[7710] ^ n[7711];
assign t[7712] = t[7711] ^ n[7712];
assign t[7713] = t[7712] ^ n[7713];
assign t[7714] = t[7713] ^ n[7714];
assign t[7715] = t[7714] ^ n[7715];
assign t[7716] = t[7715] ^ n[7716];
assign t[7717] = t[7716] ^ n[7717];
assign t[7718] = t[7717] ^ n[7718];
assign t[7719] = t[7718] ^ n[7719];
assign t[7720] = t[7719] ^ n[7720];
assign t[7721] = t[7720] ^ n[7721];
assign t[7722] = t[7721] ^ n[7722];
assign t[7723] = t[7722] ^ n[7723];
assign t[7724] = t[7723] ^ n[7724];
assign t[7725] = t[7724] ^ n[7725];
assign t[7726] = t[7725] ^ n[7726];
assign t[7727] = t[7726] ^ n[7727];
assign t[7728] = t[7727] ^ n[7728];
assign t[7729] = t[7728] ^ n[7729];
assign t[7730] = t[7729] ^ n[7730];
assign t[7731] = t[7730] ^ n[7731];
assign t[7732] = t[7731] ^ n[7732];
assign t[7733] = t[7732] ^ n[7733];
assign t[7734] = t[7733] ^ n[7734];
assign t[7735] = t[7734] ^ n[7735];
assign t[7736] = t[7735] ^ n[7736];
assign t[7737] = t[7736] ^ n[7737];
assign t[7738] = t[7737] ^ n[7738];
assign t[7739] = t[7738] ^ n[7739];
assign t[7740] = t[7739] ^ n[7740];
assign t[7741] = t[7740] ^ n[7741];
assign t[7742] = t[7741] ^ n[7742];
assign t[7743] = t[7742] ^ n[7743];
assign t[7744] = t[7743] ^ n[7744];
assign t[7745] = t[7744] ^ n[7745];
assign t[7746] = t[7745] ^ n[7746];
assign t[7747] = t[7746] ^ n[7747];
assign t[7748] = t[7747] ^ n[7748];
assign t[7749] = t[7748] ^ n[7749];
assign t[7750] = t[7749] ^ n[7750];
assign t[7751] = t[7750] ^ n[7751];
assign t[7752] = t[7751] ^ n[7752];
assign t[7753] = t[7752] ^ n[7753];
assign t[7754] = t[7753] ^ n[7754];
assign t[7755] = t[7754] ^ n[7755];
assign t[7756] = t[7755] ^ n[7756];
assign t[7757] = t[7756] ^ n[7757];
assign t[7758] = t[7757] ^ n[7758];
assign t[7759] = t[7758] ^ n[7759];
assign t[7760] = t[7759] ^ n[7760];
assign t[7761] = t[7760] ^ n[7761];
assign t[7762] = t[7761] ^ n[7762];
assign t[7763] = t[7762] ^ n[7763];
assign t[7764] = t[7763] ^ n[7764];
assign t[7765] = t[7764] ^ n[7765];
assign t[7766] = t[7765] ^ n[7766];
assign t[7767] = t[7766] ^ n[7767];
assign t[7768] = t[7767] ^ n[7768];
assign t[7769] = t[7768] ^ n[7769];
assign t[7770] = t[7769] ^ n[7770];
assign t[7771] = t[7770] ^ n[7771];
assign t[7772] = t[7771] ^ n[7772];
assign t[7773] = t[7772] ^ n[7773];
assign t[7774] = t[7773] ^ n[7774];
assign t[7775] = t[7774] ^ n[7775];
assign t[7776] = t[7775] ^ n[7776];
assign t[7777] = t[7776] ^ n[7777];
assign t[7778] = t[7777] ^ n[7778];
assign t[7779] = t[7778] ^ n[7779];
assign t[7780] = t[7779] ^ n[7780];
assign t[7781] = t[7780] ^ n[7781];
assign t[7782] = t[7781] ^ n[7782];
assign t[7783] = t[7782] ^ n[7783];
assign t[7784] = t[7783] ^ n[7784];
assign t[7785] = t[7784] ^ n[7785];
assign t[7786] = t[7785] ^ n[7786];
assign t[7787] = t[7786] ^ n[7787];
assign t[7788] = t[7787] ^ n[7788];
assign t[7789] = t[7788] ^ n[7789];
assign t[7790] = t[7789] ^ n[7790];
assign t[7791] = t[7790] ^ n[7791];
assign t[7792] = t[7791] ^ n[7792];
assign t[7793] = t[7792] ^ n[7793];
assign t[7794] = t[7793] ^ n[7794];
assign t[7795] = t[7794] ^ n[7795];
assign t[7796] = t[7795] ^ n[7796];
assign t[7797] = t[7796] ^ n[7797];
assign t[7798] = t[7797] ^ n[7798];
assign t[7799] = t[7798] ^ n[7799];
assign t[7800] = t[7799] ^ n[7800];
assign t[7801] = t[7800] ^ n[7801];
assign t[7802] = t[7801] ^ n[7802];
assign t[7803] = t[7802] ^ n[7803];
assign t[7804] = t[7803] ^ n[7804];
assign t[7805] = t[7804] ^ n[7805];
assign t[7806] = t[7805] ^ n[7806];
assign t[7807] = t[7806] ^ n[7807];
assign t[7808] = t[7807] ^ n[7808];
assign t[7809] = t[7808] ^ n[7809];
assign t[7810] = t[7809] ^ n[7810];
assign t[7811] = t[7810] ^ n[7811];
assign t[7812] = t[7811] ^ n[7812];
assign t[7813] = t[7812] ^ n[7813];
assign t[7814] = t[7813] ^ n[7814];
assign t[7815] = t[7814] ^ n[7815];
assign t[7816] = t[7815] ^ n[7816];
assign t[7817] = t[7816] ^ n[7817];
assign t[7818] = t[7817] ^ n[7818];
assign t[7819] = t[7818] ^ n[7819];
assign t[7820] = t[7819] ^ n[7820];
assign t[7821] = t[7820] ^ n[7821];
assign t[7822] = t[7821] ^ n[7822];
assign t[7823] = t[7822] ^ n[7823];
assign t[7824] = t[7823] ^ n[7824];
assign t[7825] = t[7824] ^ n[7825];
assign t[7826] = t[7825] ^ n[7826];
assign t[7827] = t[7826] ^ n[7827];
assign t[7828] = t[7827] ^ n[7828];
assign t[7829] = t[7828] ^ n[7829];
assign t[7830] = t[7829] ^ n[7830];
assign t[7831] = t[7830] ^ n[7831];
assign t[7832] = t[7831] ^ n[7832];
assign t[7833] = t[7832] ^ n[7833];
assign t[7834] = t[7833] ^ n[7834];
assign t[7835] = t[7834] ^ n[7835];
assign t[7836] = t[7835] ^ n[7836];
assign t[7837] = t[7836] ^ n[7837];
assign t[7838] = t[7837] ^ n[7838];
assign t[7839] = t[7838] ^ n[7839];
assign t[7840] = t[7839] ^ n[7840];
assign t[7841] = t[7840] ^ n[7841];
assign t[7842] = t[7841] ^ n[7842];
assign t[7843] = t[7842] ^ n[7843];
assign t[7844] = t[7843] ^ n[7844];
assign t[7845] = t[7844] ^ n[7845];
assign t[7846] = t[7845] ^ n[7846];
assign t[7847] = t[7846] ^ n[7847];
assign t[7848] = t[7847] ^ n[7848];
assign t[7849] = t[7848] ^ n[7849];
assign t[7850] = t[7849] ^ n[7850];
assign t[7851] = t[7850] ^ n[7851];
assign t[7852] = t[7851] ^ n[7852];
assign t[7853] = t[7852] ^ n[7853];
assign t[7854] = t[7853] ^ n[7854];
assign t[7855] = t[7854] ^ n[7855];
assign t[7856] = t[7855] ^ n[7856];
assign t[7857] = t[7856] ^ n[7857];
assign t[7858] = t[7857] ^ n[7858];
assign t[7859] = t[7858] ^ n[7859];
assign t[7860] = t[7859] ^ n[7860];
assign t[7861] = t[7860] ^ n[7861];
assign t[7862] = t[7861] ^ n[7862];
assign t[7863] = t[7862] ^ n[7863];
assign t[7864] = t[7863] ^ n[7864];
assign t[7865] = t[7864] ^ n[7865];
assign t[7866] = t[7865] ^ n[7866];
assign t[7867] = t[7866] ^ n[7867];
assign t[7868] = t[7867] ^ n[7868];
assign t[7869] = t[7868] ^ n[7869];
assign t[7870] = t[7869] ^ n[7870];
assign t[7871] = t[7870] ^ n[7871];
assign t[7872] = t[7871] ^ n[7872];
assign t[7873] = t[7872] ^ n[7873];
assign t[7874] = t[7873] ^ n[7874];
assign t[7875] = t[7874] ^ n[7875];
assign t[7876] = t[7875] ^ n[7876];
assign t[7877] = t[7876] ^ n[7877];
assign t[7878] = t[7877] ^ n[7878];
assign t[7879] = t[7878] ^ n[7879];
assign t[7880] = t[7879] ^ n[7880];
assign t[7881] = t[7880] ^ n[7881];
assign t[7882] = t[7881] ^ n[7882];
assign t[7883] = t[7882] ^ n[7883];
assign t[7884] = t[7883] ^ n[7884];
assign t[7885] = t[7884] ^ n[7885];
assign t[7886] = t[7885] ^ n[7886];
assign t[7887] = t[7886] ^ n[7887];
assign t[7888] = t[7887] ^ n[7888];
assign t[7889] = t[7888] ^ n[7889];
assign t[7890] = t[7889] ^ n[7890];
assign t[7891] = t[7890] ^ n[7891];
assign t[7892] = t[7891] ^ n[7892];
assign t[7893] = t[7892] ^ n[7893];
assign t[7894] = t[7893] ^ n[7894];
assign t[7895] = t[7894] ^ n[7895];
assign t[7896] = t[7895] ^ n[7896];
assign t[7897] = t[7896] ^ n[7897];
assign t[7898] = t[7897] ^ n[7898];
assign t[7899] = t[7898] ^ n[7899];
assign t[7900] = t[7899] ^ n[7900];
assign t[7901] = t[7900] ^ n[7901];
assign t[7902] = t[7901] ^ n[7902];
assign t[7903] = t[7902] ^ n[7903];
assign t[7904] = t[7903] ^ n[7904];
assign t[7905] = t[7904] ^ n[7905];
assign t[7906] = t[7905] ^ n[7906];
assign t[7907] = t[7906] ^ n[7907];
assign t[7908] = t[7907] ^ n[7908];
assign t[7909] = t[7908] ^ n[7909];
assign t[7910] = t[7909] ^ n[7910];
assign t[7911] = t[7910] ^ n[7911];
assign t[7912] = t[7911] ^ n[7912];
assign t[7913] = t[7912] ^ n[7913];
assign t[7914] = t[7913] ^ n[7914];
assign t[7915] = t[7914] ^ n[7915];
assign t[7916] = t[7915] ^ n[7916];
assign t[7917] = t[7916] ^ n[7917];
assign t[7918] = t[7917] ^ n[7918];
assign t[7919] = t[7918] ^ n[7919];
assign t[7920] = t[7919] ^ n[7920];
assign t[7921] = t[7920] ^ n[7921];
assign t[7922] = t[7921] ^ n[7922];
assign t[7923] = t[7922] ^ n[7923];
assign t[7924] = t[7923] ^ n[7924];
assign t[7925] = t[7924] ^ n[7925];
assign t[7926] = t[7925] ^ n[7926];
assign t[7927] = t[7926] ^ n[7927];
assign t[7928] = t[7927] ^ n[7928];
assign t[7929] = t[7928] ^ n[7929];
assign t[7930] = t[7929] ^ n[7930];
assign t[7931] = t[7930] ^ n[7931];
assign t[7932] = t[7931] ^ n[7932];
assign t[7933] = t[7932] ^ n[7933];
assign t[7934] = t[7933] ^ n[7934];
assign t[7935] = t[7934] ^ n[7935];
assign t[7936] = t[7935] ^ n[7936];
assign t[7937] = t[7936] ^ n[7937];
assign t[7938] = t[7937] ^ n[7938];
assign t[7939] = t[7938] ^ n[7939];
assign t[7940] = t[7939] ^ n[7940];
assign t[7941] = t[7940] ^ n[7941];
assign t[7942] = t[7941] ^ n[7942];
assign t[7943] = t[7942] ^ n[7943];
assign t[7944] = t[7943] ^ n[7944];
assign t[7945] = t[7944] ^ n[7945];
assign t[7946] = t[7945] ^ n[7946];
assign t[7947] = t[7946] ^ n[7947];
assign t[7948] = t[7947] ^ n[7948];
assign t[7949] = t[7948] ^ n[7949];
assign t[7950] = t[7949] ^ n[7950];
assign t[7951] = t[7950] ^ n[7951];
assign t[7952] = t[7951] ^ n[7952];
assign t[7953] = t[7952] ^ n[7953];
assign t[7954] = t[7953] ^ n[7954];
assign t[7955] = t[7954] ^ n[7955];
assign t[7956] = t[7955] ^ n[7956];
assign t[7957] = t[7956] ^ n[7957];
assign t[7958] = t[7957] ^ n[7958];
assign t[7959] = t[7958] ^ n[7959];
assign t[7960] = t[7959] ^ n[7960];
assign t[7961] = t[7960] ^ n[7961];
assign t[7962] = t[7961] ^ n[7962];
assign t[7963] = t[7962] ^ n[7963];
assign t[7964] = t[7963] ^ n[7964];
assign t[7965] = t[7964] ^ n[7965];
assign t[7966] = t[7965] ^ n[7966];
assign t[7967] = t[7966] ^ n[7967];
assign t[7968] = t[7967] ^ n[7968];
assign t[7969] = t[7968] ^ n[7969];
assign t[7970] = t[7969] ^ n[7970];
assign t[7971] = t[7970] ^ n[7971];
assign t[7972] = t[7971] ^ n[7972];
assign t[7973] = t[7972] ^ n[7973];
assign t[7974] = t[7973] ^ n[7974];
assign t[7975] = t[7974] ^ n[7975];
assign t[7976] = t[7975] ^ n[7976];
assign t[7977] = t[7976] ^ n[7977];
assign t[7978] = t[7977] ^ n[7978];
assign t[7979] = t[7978] ^ n[7979];
assign t[7980] = t[7979] ^ n[7980];
assign t[7981] = t[7980] ^ n[7981];
assign t[7982] = t[7981] ^ n[7982];
assign t[7983] = t[7982] ^ n[7983];
assign t[7984] = t[7983] ^ n[7984];
assign t[7985] = t[7984] ^ n[7985];
assign t[7986] = t[7985] ^ n[7986];
assign t[7987] = t[7986] ^ n[7987];
assign t[7988] = t[7987] ^ n[7988];
assign t[7989] = t[7988] ^ n[7989];
assign t[7990] = t[7989] ^ n[7990];
assign t[7991] = t[7990] ^ n[7991];
assign t[7992] = t[7991] ^ n[7992];
assign t[7993] = t[7992] ^ n[7993];
assign t[7994] = t[7993] ^ n[7994];
assign t[7995] = t[7994] ^ n[7995];
assign t[7996] = t[7995] ^ n[7996];
assign t[7997] = t[7996] ^ n[7997];
assign t[7998] = t[7997] ^ n[7998];
assign t[7999] = t[7998] ^ n[7999];
assign t[8000] = t[7999] ^ n[8000];
assign t[8001] = t[8000] ^ n[8001];
assign t[8002] = t[8001] ^ n[8002];
assign t[8003] = t[8002] ^ n[8003];
assign t[8004] = t[8003] ^ n[8004];
assign t[8005] = t[8004] ^ n[8005];
assign t[8006] = t[8005] ^ n[8006];
assign t[8007] = t[8006] ^ n[8007];
assign t[8008] = t[8007] ^ n[8008];
assign t[8009] = t[8008] ^ n[8009];
assign t[8010] = t[8009] ^ n[8010];
assign t[8011] = t[8010] ^ n[8011];
assign t[8012] = t[8011] ^ n[8012];
assign t[8013] = t[8012] ^ n[8013];
assign t[8014] = t[8013] ^ n[8014];
assign t[8015] = t[8014] ^ n[8015];
assign t[8016] = t[8015] ^ n[8016];
assign t[8017] = t[8016] ^ n[8017];
assign t[8018] = t[8017] ^ n[8018];
assign t[8019] = t[8018] ^ n[8019];
assign t[8020] = t[8019] ^ n[8020];
assign t[8021] = t[8020] ^ n[8021];
assign t[8022] = t[8021] ^ n[8022];
assign t[8023] = t[8022] ^ n[8023];
assign t[8024] = t[8023] ^ n[8024];
assign t[8025] = t[8024] ^ n[8025];
assign t[8026] = t[8025] ^ n[8026];
assign t[8027] = t[8026] ^ n[8027];
assign t[8028] = t[8027] ^ n[8028];
assign t[8029] = t[8028] ^ n[8029];
assign t[8030] = t[8029] ^ n[8030];
assign t[8031] = t[8030] ^ n[8031];
assign t[8032] = t[8031] ^ n[8032];
assign t[8033] = t[8032] ^ n[8033];
assign t[8034] = t[8033] ^ n[8034];
assign t[8035] = t[8034] ^ n[8035];
assign t[8036] = t[8035] ^ n[8036];
assign t[8037] = t[8036] ^ n[8037];
assign t[8038] = t[8037] ^ n[8038];
assign t[8039] = t[8038] ^ n[8039];
assign t[8040] = t[8039] ^ n[8040];
assign t[8041] = t[8040] ^ n[8041];
assign t[8042] = t[8041] ^ n[8042];
assign t[8043] = t[8042] ^ n[8043];
assign t[8044] = t[8043] ^ n[8044];
assign t[8045] = t[8044] ^ n[8045];
assign t[8046] = t[8045] ^ n[8046];
assign t[8047] = t[8046] ^ n[8047];
assign t[8048] = t[8047] ^ n[8048];
assign t[8049] = t[8048] ^ n[8049];
assign t[8050] = t[8049] ^ n[8050];
assign t[8051] = t[8050] ^ n[8051];
assign t[8052] = t[8051] ^ n[8052];
assign t[8053] = t[8052] ^ n[8053];
assign t[8054] = t[8053] ^ n[8054];
assign t[8055] = t[8054] ^ n[8055];
assign t[8056] = t[8055] ^ n[8056];
assign t[8057] = t[8056] ^ n[8057];
assign t[8058] = t[8057] ^ n[8058];
assign t[8059] = t[8058] ^ n[8059];
assign t[8060] = t[8059] ^ n[8060];
assign t[8061] = t[8060] ^ n[8061];
assign t[8062] = t[8061] ^ n[8062];
assign t[8063] = t[8062] ^ n[8063];
assign t[8064] = t[8063] ^ n[8064];
assign t[8065] = t[8064] ^ n[8065];
assign t[8066] = t[8065] ^ n[8066];
assign t[8067] = t[8066] ^ n[8067];
assign t[8068] = t[8067] ^ n[8068];
assign t[8069] = t[8068] ^ n[8069];
assign t[8070] = t[8069] ^ n[8070];
assign t[8071] = t[8070] ^ n[8071];
assign t[8072] = t[8071] ^ n[8072];
assign t[8073] = t[8072] ^ n[8073];
assign t[8074] = t[8073] ^ n[8074];
assign t[8075] = t[8074] ^ n[8075];
assign t[8076] = t[8075] ^ n[8076];
assign t[8077] = t[8076] ^ n[8077];
assign t[8078] = t[8077] ^ n[8078];
assign t[8079] = t[8078] ^ n[8079];
assign t[8080] = t[8079] ^ n[8080];
assign t[8081] = t[8080] ^ n[8081];
assign t[8082] = t[8081] ^ n[8082];
assign t[8083] = t[8082] ^ n[8083];
assign t[8084] = t[8083] ^ n[8084];
assign t[8085] = t[8084] ^ n[8085];
assign t[8086] = t[8085] ^ n[8086];
assign t[8087] = t[8086] ^ n[8087];
assign t[8088] = t[8087] ^ n[8088];
assign t[8089] = t[8088] ^ n[8089];
assign t[8090] = t[8089] ^ n[8090];
assign t[8091] = t[8090] ^ n[8091];
assign t[8092] = t[8091] ^ n[8092];
assign t[8093] = t[8092] ^ n[8093];
assign t[8094] = t[8093] ^ n[8094];
assign t[8095] = t[8094] ^ n[8095];
assign t[8096] = t[8095] ^ n[8096];
assign t[8097] = t[8096] ^ n[8097];
assign t[8098] = t[8097] ^ n[8098];
assign t[8099] = t[8098] ^ n[8099];
assign t[8100] = t[8099] ^ n[8100];
assign t[8101] = t[8100] ^ n[8101];
assign t[8102] = t[8101] ^ n[8102];
assign t[8103] = t[8102] ^ n[8103];
assign t[8104] = t[8103] ^ n[8104];
assign t[8105] = t[8104] ^ n[8105];
assign t[8106] = t[8105] ^ n[8106];
assign t[8107] = t[8106] ^ n[8107];
assign t[8108] = t[8107] ^ n[8108];
assign t[8109] = t[8108] ^ n[8109];
assign t[8110] = t[8109] ^ n[8110];
assign t[8111] = t[8110] ^ n[8111];
assign t[8112] = t[8111] ^ n[8112];
assign t[8113] = t[8112] ^ n[8113];
assign t[8114] = t[8113] ^ n[8114];
assign t[8115] = t[8114] ^ n[8115];
assign t[8116] = t[8115] ^ n[8116];
assign t[8117] = t[8116] ^ n[8117];
assign t[8118] = t[8117] ^ n[8118];
assign t[8119] = t[8118] ^ n[8119];
assign t[8120] = t[8119] ^ n[8120];
assign t[8121] = t[8120] ^ n[8121];
assign t[8122] = t[8121] ^ n[8122];
assign t[8123] = t[8122] ^ n[8123];
assign t[8124] = t[8123] ^ n[8124];
assign t[8125] = t[8124] ^ n[8125];
assign t[8126] = t[8125] ^ n[8126];
assign t[8127] = t[8126] ^ n[8127];
assign t[8128] = t[8127] ^ n[8128];
assign t[8129] = t[8128] ^ n[8129];
assign t[8130] = t[8129] ^ n[8130];
assign t[8131] = t[8130] ^ n[8131];
assign t[8132] = t[8131] ^ n[8132];
assign t[8133] = t[8132] ^ n[8133];
assign t[8134] = t[8133] ^ n[8134];
assign t[8135] = t[8134] ^ n[8135];
assign t[8136] = t[8135] ^ n[8136];
assign t[8137] = t[8136] ^ n[8137];
assign t[8138] = t[8137] ^ n[8138];
assign t[8139] = t[8138] ^ n[8139];
assign t[8140] = t[8139] ^ n[8140];
assign t[8141] = t[8140] ^ n[8141];
assign t[8142] = t[8141] ^ n[8142];
assign t[8143] = t[8142] ^ n[8143];
assign t[8144] = t[8143] ^ n[8144];
assign t[8145] = t[8144] ^ n[8145];
assign t[8146] = t[8145] ^ n[8146];
assign t[8147] = t[8146] ^ n[8147];
assign t[8148] = t[8147] ^ n[8148];
assign t[8149] = t[8148] ^ n[8149];
assign t[8150] = t[8149] ^ n[8150];
assign t[8151] = t[8150] ^ n[8151];
assign t[8152] = t[8151] ^ n[8152];
assign t[8153] = t[8152] ^ n[8153];
assign t[8154] = t[8153] ^ n[8154];
assign t[8155] = t[8154] ^ n[8155];
assign t[8156] = t[8155] ^ n[8156];
assign t[8157] = t[8156] ^ n[8157];
assign t[8158] = t[8157] ^ n[8158];
assign t[8159] = t[8158] ^ n[8159];
assign t[8160] = t[8159] ^ n[8160];
assign t[8161] = t[8160] ^ n[8161];
assign t[8162] = t[8161] ^ n[8162];
assign t[8163] = t[8162] ^ n[8163];
assign t[8164] = t[8163] ^ n[8164];
assign t[8165] = t[8164] ^ n[8165];
assign t[8166] = t[8165] ^ n[8166];
assign t[8167] = t[8166] ^ n[8167];
assign t[8168] = t[8167] ^ n[8168];
assign t[8169] = t[8168] ^ n[8169];
assign t[8170] = t[8169] ^ n[8170];
assign t[8171] = t[8170] ^ n[8171];
assign t[8172] = t[8171] ^ n[8172];
assign t[8173] = t[8172] ^ n[8173];
assign t[8174] = t[8173] ^ n[8174];
assign t[8175] = t[8174] ^ n[8175];
assign t[8176] = t[8175] ^ n[8176];
assign t[8177] = t[8176] ^ n[8177];

//asigning bit 12
assign s[12] = ( a[12] ^ b [12] ) ^ t[8177];

assign t[8178] = n[8178];
assign t[8179] = t[8178] ^ n[8179];
assign t[8180] = t[8179] ^ n[8180];
assign t[8181] = t[8180] ^ n[8181];
assign t[8182] = t[8181] ^ n[8182];
assign t[8183] = t[8182] ^ n[8183];
assign t[8184] = t[8183] ^ n[8184];
assign t[8185] = t[8184] ^ n[8185];
assign t[8186] = t[8185] ^ n[8186];
assign t[8187] = t[8186] ^ n[8187];
assign t[8188] = t[8187] ^ n[8188];
assign t[8189] = t[8188] ^ n[8189];
assign t[8190] = t[8189] ^ n[8190];
assign t[8191] = t[8190] ^ n[8191];
assign t[8192] = t[8191] ^ n[8192];
assign t[8193] = t[8192] ^ n[8193];
assign t[8194] = t[8193] ^ n[8194];
assign t[8195] = t[8194] ^ n[8195];
assign t[8196] = t[8195] ^ n[8196];
assign t[8197] = t[8196] ^ n[8197];
assign t[8198] = t[8197] ^ n[8198];
assign t[8199] = t[8198] ^ n[8199];
assign t[8200] = t[8199] ^ n[8200];
assign t[8201] = t[8200] ^ n[8201];
assign t[8202] = t[8201] ^ n[8202];
assign t[8203] = t[8202] ^ n[8203];
assign t[8204] = t[8203] ^ n[8204];
assign t[8205] = t[8204] ^ n[8205];
assign t[8206] = t[8205] ^ n[8206];
assign t[8207] = t[8206] ^ n[8207];
assign t[8208] = t[8207] ^ n[8208];
assign t[8209] = t[8208] ^ n[8209];
assign t[8210] = t[8209] ^ n[8210];
assign t[8211] = t[8210] ^ n[8211];
assign t[8212] = t[8211] ^ n[8212];
assign t[8213] = t[8212] ^ n[8213];
assign t[8214] = t[8213] ^ n[8214];
assign t[8215] = t[8214] ^ n[8215];
assign t[8216] = t[8215] ^ n[8216];
assign t[8217] = t[8216] ^ n[8217];
assign t[8218] = t[8217] ^ n[8218];
assign t[8219] = t[8218] ^ n[8219];
assign t[8220] = t[8219] ^ n[8220];
assign t[8221] = t[8220] ^ n[8221];
assign t[8222] = t[8221] ^ n[8222];
assign t[8223] = t[8222] ^ n[8223];
assign t[8224] = t[8223] ^ n[8224];
assign t[8225] = t[8224] ^ n[8225];
assign t[8226] = t[8225] ^ n[8226];
assign t[8227] = t[8226] ^ n[8227];
assign t[8228] = t[8227] ^ n[8228];
assign t[8229] = t[8228] ^ n[8229];
assign t[8230] = t[8229] ^ n[8230];
assign t[8231] = t[8230] ^ n[8231];
assign t[8232] = t[8231] ^ n[8232];
assign t[8233] = t[8232] ^ n[8233];
assign t[8234] = t[8233] ^ n[8234];
assign t[8235] = t[8234] ^ n[8235];
assign t[8236] = t[8235] ^ n[8236];
assign t[8237] = t[8236] ^ n[8237];
assign t[8238] = t[8237] ^ n[8238];
assign t[8239] = t[8238] ^ n[8239];
assign t[8240] = t[8239] ^ n[8240];
assign t[8241] = t[8240] ^ n[8241];
assign t[8242] = t[8241] ^ n[8242];
assign t[8243] = t[8242] ^ n[8243];
assign t[8244] = t[8243] ^ n[8244];
assign t[8245] = t[8244] ^ n[8245];
assign t[8246] = t[8245] ^ n[8246];
assign t[8247] = t[8246] ^ n[8247];
assign t[8248] = t[8247] ^ n[8248];
assign t[8249] = t[8248] ^ n[8249];
assign t[8250] = t[8249] ^ n[8250];
assign t[8251] = t[8250] ^ n[8251];
assign t[8252] = t[8251] ^ n[8252];
assign t[8253] = t[8252] ^ n[8253];
assign t[8254] = t[8253] ^ n[8254];
assign t[8255] = t[8254] ^ n[8255];
assign t[8256] = t[8255] ^ n[8256];
assign t[8257] = t[8256] ^ n[8257];
assign t[8258] = t[8257] ^ n[8258];
assign t[8259] = t[8258] ^ n[8259];
assign t[8260] = t[8259] ^ n[8260];
assign t[8261] = t[8260] ^ n[8261];
assign t[8262] = t[8261] ^ n[8262];
assign t[8263] = t[8262] ^ n[8263];
assign t[8264] = t[8263] ^ n[8264];
assign t[8265] = t[8264] ^ n[8265];
assign t[8266] = t[8265] ^ n[8266];
assign t[8267] = t[8266] ^ n[8267];
assign t[8268] = t[8267] ^ n[8268];
assign t[8269] = t[8268] ^ n[8269];
assign t[8270] = t[8269] ^ n[8270];
assign t[8271] = t[8270] ^ n[8271];
assign t[8272] = t[8271] ^ n[8272];
assign t[8273] = t[8272] ^ n[8273];
assign t[8274] = t[8273] ^ n[8274];
assign t[8275] = t[8274] ^ n[8275];
assign t[8276] = t[8275] ^ n[8276];
assign t[8277] = t[8276] ^ n[8277];
assign t[8278] = t[8277] ^ n[8278];
assign t[8279] = t[8278] ^ n[8279];
assign t[8280] = t[8279] ^ n[8280];
assign t[8281] = t[8280] ^ n[8281];
assign t[8282] = t[8281] ^ n[8282];
assign t[8283] = t[8282] ^ n[8283];
assign t[8284] = t[8283] ^ n[8284];
assign t[8285] = t[8284] ^ n[8285];
assign t[8286] = t[8285] ^ n[8286];
assign t[8287] = t[8286] ^ n[8287];
assign t[8288] = t[8287] ^ n[8288];
assign t[8289] = t[8288] ^ n[8289];
assign t[8290] = t[8289] ^ n[8290];
assign t[8291] = t[8290] ^ n[8291];
assign t[8292] = t[8291] ^ n[8292];
assign t[8293] = t[8292] ^ n[8293];
assign t[8294] = t[8293] ^ n[8294];
assign t[8295] = t[8294] ^ n[8295];
assign t[8296] = t[8295] ^ n[8296];
assign t[8297] = t[8296] ^ n[8297];
assign t[8298] = t[8297] ^ n[8298];
assign t[8299] = t[8298] ^ n[8299];
assign t[8300] = t[8299] ^ n[8300];
assign t[8301] = t[8300] ^ n[8301];
assign t[8302] = t[8301] ^ n[8302];
assign t[8303] = t[8302] ^ n[8303];
assign t[8304] = t[8303] ^ n[8304];
assign t[8305] = t[8304] ^ n[8305];
assign t[8306] = t[8305] ^ n[8306];
assign t[8307] = t[8306] ^ n[8307];
assign t[8308] = t[8307] ^ n[8308];
assign t[8309] = t[8308] ^ n[8309];
assign t[8310] = t[8309] ^ n[8310];
assign t[8311] = t[8310] ^ n[8311];
assign t[8312] = t[8311] ^ n[8312];
assign t[8313] = t[8312] ^ n[8313];
assign t[8314] = t[8313] ^ n[8314];
assign t[8315] = t[8314] ^ n[8315];
assign t[8316] = t[8315] ^ n[8316];
assign t[8317] = t[8316] ^ n[8317];
assign t[8318] = t[8317] ^ n[8318];
assign t[8319] = t[8318] ^ n[8319];
assign t[8320] = t[8319] ^ n[8320];
assign t[8321] = t[8320] ^ n[8321];
assign t[8322] = t[8321] ^ n[8322];
assign t[8323] = t[8322] ^ n[8323];
assign t[8324] = t[8323] ^ n[8324];
assign t[8325] = t[8324] ^ n[8325];
assign t[8326] = t[8325] ^ n[8326];
assign t[8327] = t[8326] ^ n[8327];
assign t[8328] = t[8327] ^ n[8328];
assign t[8329] = t[8328] ^ n[8329];
assign t[8330] = t[8329] ^ n[8330];
assign t[8331] = t[8330] ^ n[8331];
assign t[8332] = t[8331] ^ n[8332];
assign t[8333] = t[8332] ^ n[8333];
assign t[8334] = t[8333] ^ n[8334];
assign t[8335] = t[8334] ^ n[8335];
assign t[8336] = t[8335] ^ n[8336];
assign t[8337] = t[8336] ^ n[8337];
assign t[8338] = t[8337] ^ n[8338];
assign t[8339] = t[8338] ^ n[8339];
assign t[8340] = t[8339] ^ n[8340];
assign t[8341] = t[8340] ^ n[8341];
assign t[8342] = t[8341] ^ n[8342];
assign t[8343] = t[8342] ^ n[8343];
assign t[8344] = t[8343] ^ n[8344];
assign t[8345] = t[8344] ^ n[8345];
assign t[8346] = t[8345] ^ n[8346];
assign t[8347] = t[8346] ^ n[8347];
assign t[8348] = t[8347] ^ n[8348];
assign t[8349] = t[8348] ^ n[8349];
assign t[8350] = t[8349] ^ n[8350];
assign t[8351] = t[8350] ^ n[8351];
assign t[8352] = t[8351] ^ n[8352];
assign t[8353] = t[8352] ^ n[8353];
assign t[8354] = t[8353] ^ n[8354];
assign t[8355] = t[8354] ^ n[8355];
assign t[8356] = t[8355] ^ n[8356];
assign t[8357] = t[8356] ^ n[8357];
assign t[8358] = t[8357] ^ n[8358];
assign t[8359] = t[8358] ^ n[8359];
assign t[8360] = t[8359] ^ n[8360];
assign t[8361] = t[8360] ^ n[8361];
assign t[8362] = t[8361] ^ n[8362];
assign t[8363] = t[8362] ^ n[8363];
assign t[8364] = t[8363] ^ n[8364];
assign t[8365] = t[8364] ^ n[8365];
assign t[8366] = t[8365] ^ n[8366];
assign t[8367] = t[8366] ^ n[8367];
assign t[8368] = t[8367] ^ n[8368];
assign t[8369] = t[8368] ^ n[8369];
assign t[8370] = t[8369] ^ n[8370];
assign t[8371] = t[8370] ^ n[8371];
assign t[8372] = t[8371] ^ n[8372];
assign t[8373] = t[8372] ^ n[8373];
assign t[8374] = t[8373] ^ n[8374];
assign t[8375] = t[8374] ^ n[8375];
assign t[8376] = t[8375] ^ n[8376];
assign t[8377] = t[8376] ^ n[8377];
assign t[8378] = t[8377] ^ n[8378];
assign t[8379] = t[8378] ^ n[8379];
assign t[8380] = t[8379] ^ n[8380];
assign t[8381] = t[8380] ^ n[8381];
assign t[8382] = t[8381] ^ n[8382];
assign t[8383] = t[8382] ^ n[8383];
assign t[8384] = t[8383] ^ n[8384];
assign t[8385] = t[8384] ^ n[8385];
assign t[8386] = t[8385] ^ n[8386];
assign t[8387] = t[8386] ^ n[8387];
assign t[8388] = t[8387] ^ n[8388];
assign t[8389] = t[8388] ^ n[8389];
assign t[8390] = t[8389] ^ n[8390];
assign t[8391] = t[8390] ^ n[8391];
assign t[8392] = t[8391] ^ n[8392];
assign t[8393] = t[8392] ^ n[8393];
assign t[8394] = t[8393] ^ n[8394];
assign t[8395] = t[8394] ^ n[8395];
assign t[8396] = t[8395] ^ n[8396];
assign t[8397] = t[8396] ^ n[8397];
assign t[8398] = t[8397] ^ n[8398];
assign t[8399] = t[8398] ^ n[8399];
assign t[8400] = t[8399] ^ n[8400];
assign t[8401] = t[8400] ^ n[8401];
assign t[8402] = t[8401] ^ n[8402];
assign t[8403] = t[8402] ^ n[8403];
assign t[8404] = t[8403] ^ n[8404];
assign t[8405] = t[8404] ^ n[8405];
assign t[8406] = t[8405] ^ n[8406];
assign t[8407] = t[8406] ^ n[8407];
assign t[8408] = t[8407] ^ n[8408];
assign t[8409] = t[8408] ^ n[8409];
assign t[8410] = t[8409] ^ n[8410];
assign t[8411] = t[8410] ^ n[8411];
assign t[8412] = t[8411] ^ n[8412];
assign t[8413] = t[8412] ^ n[8413];
assign t[8414] = t[8413] ^ n[8414];
assign t[8415] = t[8414] ^ n[8415];
assign t[8416] = t[8415] ^ n[8416];
assign t[8417] = t[8416] ^ n[8417];
assign t[8418] = t[8417] ^ n[8418];
assign t[8419] = t[8418] ^ n[8419];
assign t[8420] = t[8419] ^ n[8420];
assign t[8421] = t[8420] ^ n[8421];
assign t[8422] = t[8421] ^ n[8422];
assign t[8423] = t[8422] ^ n[8423];
assign t[8424] = t[8423] ^ n[8424];
assign t[8425] = t[8424] ^ n[8425];
assign t[8426] = t[8425] ^ n[8426];
assign t[8427] = t[8426] ^ n[8427];
assign t[8428] = t[8427] ^ n[8428];
assign t[8429] = t[8428] ^ n[8429];
assign t[8430] = t[8429] ^ n[8430];
assign t[8431] = t[8430] ^ n[8431];
assign t[8432] = t[8431] ^ n[8432];
assign t[8433] = t[8432] ^ n[8433];
assign t[8434] = t[8433] ^ n[8434];
assign t[8435] = t[8434] ^ n[8435];
assign t[8436] = t[8435] ^ n[8436];
assign t[8437] = t[8436] ^ n[8437];
assign t[8438] = t[8437] ^ n[8438];
assign t[8439] = t[8438] ^ n[8439];
assign t[8440] = t[8439] ^ n[8440];
assign t[8441] = t[8440] ^ n[8441];
assign t[8442] = t[8441] ^ n[8442];
assign t[8443] = t[8442] ^ n[8443];
assign t[8444] = t[8443] ^ n[8444];
assign t[8445] = t[8444] ^ n[8445];
assign t[8446] = t[8445] ^ n[8446];
assign t[8447] = t[8446] ^ n[8447];
assign t[8448] = t[8447] ^ n[8448];
assign t[8449] = t[8448] ^ n[8449];
assign t[8450] = t[8449] ^ n[8450];
assign t[8451] = t[8450] ^ n[8451];
assign t[8452] = t[8451] ^ n[8452];
assign t[8453] = t[8452] ^ n[8453];
assign t[8454] = t[8453] ^ n[8454];
assign t[8455] = t[8454] ^ n[8455];
assign t[8456] = t[8455] ^ n[8456];
assign t[8457] = t[8456] ^ n[8457];
assign t[8458] = t[8457] ^ n[8458];
assign t[8459] = t[8458] ^ n[8459];
assign t[8460] = t[8459] ^ n[8460];
assign t[8461] = t[8460] ^ n[8461];
assign t[8462] = t[8461] ^ n[8462];
assign t[8463] = t[8462] ^ n[8463];
assign t[8464] = t[8463] ^ n[8464];
assign t[8465] = t[8464] ^ n[8465];
assign t[8466] = t[8465] ^ n[8466];
assign t[8467] = t[8466] ^ n[8467];
assign t[8468] = t[8467] ^ n[8468];
assign t[8469] = t[8468] ^ n[8469];
assign t[8470] = t[8469] ^ n[8470];
assign t[8471] = t[8470] ^ n[8471];
assign t[8472] = t[8471] ^ n[8472];
assign t[8473] = t[8472] ^ n[8473];
assign t[8474] = t[8473] ^ n[8474];
assign t[8475] = t[8474] ^ n[8475];
assign t[8476] = t[8475] ^ n[8476];
assign t[8477] = t[8476] ^ n[8477];
assign t[8478] = t[8477] ^ n[8478];
assign t[8479] = t[8478] ^ n[8479];
assign t[8480] = t[8479] ^ n[8480];
assign t[8481] = t[8480] ^ n[8481];
assign t[8482] = t[8481] ^ n[8482];
assign t[8483] = t[8482] ^ n[8483];
assign t[8484] = t[8483] ^ n[8484];
assign t[8485] = t[8484] ^ n[8485];
assign t[8486] = t[8485] ^ n[8486];
assign t[8487] = t[8486] ^ n[8487];
assign t[8488] = t[8487] ^ n[8488];
assign t[8489] = t[8488] ^ n[8489];
assign t[8490] = t[8489] ^ n[8490];
assign t[8491] = t[8490] ^ n[8491];
assign t[8492] = t[8491] ^ n[8492];
assign t[8493] = t[8492] ^ n[8493];
assign t[8494] = t[8493] ^ n[8494];
assign t[8495] = t[8494] ^ n[8495];
assign t[8496] = t[8495] ^ n[8496];
assign t[8497] = t[8496] ^ n[8497];
assign t[8498] = t[8497] ^ n[8498];
assign t[8499] = t[8498] ^ n[8499];
assign t[8500] = t[8499] ^ n[8500];
assign t[8501] = t[8500] ^ n[8501];
assign t[8502] = t[8501] ^ n[8502];
assign t[8503] = t[8502] ^ n[8503];
assign t[8504] = t[8503] ^ n[8504];
assign t[8505] = t[8504] ^ n[8505];
assign t[8506] = t[8505] ^ n[8506];
assign t[8507] = t[8506] ^ n[8507];
assign t[8508] = t[8507] ^ n[8508];
assign t[8509] = t[8508] ^ n[8509];
assign t[8510] = t[8509] ^ n[8510];
assign t[8511] = t[8510] ^ n[8511];
assign t[8512] = t[8511] ^ n[8512];
assign t[8513] = t[8512] ^ n[8513];
assign t[8514] = t[8513] ^ n[8514];
assign t[8515] = t[8514] ^ n[8515];
assign t[8516] = t[8515] ^ n[8516];
assign t[8517] = t[8516] ^ n[8517];
assign t[8518] = t[8517] ^ n[8518];
assign t[8519] = t[8518] ^ n[8519];
assign t[8520] = t[8519] ^ n[8520];
assign t[8521] = t[8520] ^ n[8521];
assign t[8522] = t[8521] ^ n[8522];
assign t[8523] = t[8522] ^ n[8523];
assign t[8524] = t[8523] ^ n[8524];
assign t[8525] = t[8524] ^ n[8525];
assign t[8526] = t[8525] ^ n[8526];
assign t[8527] = t[8526] ^ n[8527];
assign t[8528] = t[8527] ^ n[8528];
assign t[8529] = t[8528] ^ n[8529];
assign t[8530] = t[8529] ^ n[8530];
assign t[8531] = t[8530] ^ n[8531];
assign t[8532] = t[8531] ^ n[8532];
assign t[8533] = t[8532] ^ n[8533];
assign t[8534] = t[8533] ^ n[8534];
assign t[8535] = t[8534] ^ n[8535];
assign t[8536] = t[8535] ^ n[8536];
assign t[8537] = t[8536] ^ n[8537];
assign t[8538] = t[8537] ^ n[8538];
assign t[8539] = t[8538] ^ n[8539];
assign t[8540] = t[8539] ^ n[8540];
assign t[8541] = t[8540] ^ n[8541];
assign t[8542] = t[8541] ^ n[8542];
assign t[8543] = t[8542] ^ n[8543];
assign t[8544] = t[8543] ^ n[8544];
assign t[8545] = t[8544] ^ n[8545];
assign t[8546] = t[8545] ^ n[8546];
assign t[8547] = t[8546] ^ n[8547];
assign t[8548] = t[8547] ^ n[8548];
assign t[8549] = t[8548] ^ n[8549];
assign t[8550] = t[8549] ^ n[8550];
assign t[8551] = t[8550] ^ n[8551];
assign t[8552] = t[8551] ^ n[8552];
assign t[8553] = t[8552] ^ n[8553];
assign t[8554] = t[8553] ^ n[8554];
assign t[8555] = t[8554] ^ n[8555];
assign t[8556] = t[8555] ^ n[8556];
assign t[8557] = t[8556] ^ n[8557];
assign t[8558] = t[8557] ^ n[8558];
assign t[8559] = t[8558] ^ n[8559];
assign t[8560] = t[8559] ^ n[8560];
assign t[8561] = t[8560] ^ n[8561];
assign t[8562] = t[8561] ^ n[8562];
assign t[8563] = t[8562] ^ n[8563];
assign t[8564] = t[8563] ^ n[8564];
assign t[8565] = t[8564] ^ n[8565];
assign t[8566] = t[8565] ^ n[8566];
assign t[8567] = t[8566] ^ n[8567];
assign t[8568] = t[8567] ^ n[8568];
assign t[8569] = t[8568] ^ n[8569];
assign t[8570] = t[8569] ^ n[8570];
assign t[8571] = t[8570] ^ n[8571];
assign t[8572] = t[8571] ^ n[8572];
assign t[8573] = t[8572] ^ n[8573];
assign t[8574] = t[8573] ^ n[8574];
assign t[8575] = t[8574] ^ n[8575];
assign t[8576] = t[8575] ^ n[8576];
assign t[8577] = t[8576] ^ n[8577];
assign t[8578] = t[8577] ^ n[8578];
assign t[8579] = t[8578] ^ n[8579];
assign t[8580] = t[8579] ^ n[8580];
assign t[8581] = t[8580] ^ n[8581];
assign t[8582] = t[8581] ^ n[8582];
assign t[8583] = t[8582] ^ n[8583];
assign t[8584] = t[8583] ^ n[8584];
assign t[8585] = t[8584] ^ n[8585];
assign t[8586] = t[8585] ^ n[8586];
assign t[8587] = t[8586] ^ n[8587];
assign t[8588] = t[8587] ^ n[8588];
assign t[8589] = t[8588] ^ n[8589];
assign t[8590] = t[8589] ^ n[8590];
assign t[8591] = t[8590] ^ n[8591];
assign t[8592] = t[8591] ^ n[8592];
assign t[8593] = t[8592] ^ n[8593];
assign t[8594] = t[8593] ^ n[8594];
assign t[8595] = t[8594] ^ n[8595];
assign t[8596] = t[8595] ^ n[8596];
assign t[8597] = t[8596] ^ n[8597];
assign t[8598] = t[8597] ^ n[8598];
assign t[8599] = t[8598] ^ n[8599];
assign t[8600] = t[8599] ^ n[8600];
assign t[8601] = t[8600] ^ n[8601];
assign t[8602] = t[8601] ^ n[8602];
assign t[8603] = t[8602] ^ n[8603];
assign t[8604] = t[8603] ^ n[8604];
assign t[8605] = t[8604] ^ n[8605];
assign t[8606] = t[8605] ^ n[8606];
assign t[8607] = t[8606] ^ n[8607];
assign t[8608] = t[8607] ^ n[8608];
assign t[8609] = t[8608] ^ n[8609];
assign t[8610] = t[8609] ^ n[8610];
assign t[8611] = t[8610] ^ n[8611];
assign t[8612] = t[8611] ^ n[8612];
assign t[8613] = t[8612] ^ n[8613];
assign t[8614] = t[8613] ^ n[8614];
assign t[8615] = t[8614] ^ n[8615];
assign t[8616] = t[8615] ^ n[8616];
assign t[8617] = t[8616] ^ n[8617];
assign t[8618] = t[8617] ^ n[8618];
assign t[8619] = t[8618] ^ n[8619];
assign t[8620] = t[8619] ^ n[8620];
assign t[8621] = t[8620] ^ n[8621];
assign t[8622] = t[8621] ^ n[8622];
assign t[8623] = t[8622] ^ n[8623];
assign t[8624] = t[8623] ^ n[8624];
assign t[8625] = t[8624] ^ n[8625];
assign t[8626] = t[8625] ^ n[8626];
assign t[8627] = t[8626] ^ n[8627];
assign t[8628] = t[8627] ^ n[8628];
assign t[8629] = t[8628] ^ n[8629];
assign t[8630] = t[8629] ^ n[8630];
assign t[8631] = t[8630] ^ n[8631];
assign t[8632] = t[8631] ^ n[8632];
assign t[8633] = t[8632] ^ n[8633];
assign t[8634] = t[8633] ^ n[8634];
assign t[8635] = t[8634] ^ n[8635];
assign t[8636] = t[8635] ^ n[8636];
assign t[8637] = t[8636] ^ n[8637];
assign t[8638] = t[8637] ^ n[8638];
assign t[8639] = t[8638] ^ n[8639];
assign t[8640] = t[8639] ^ n[8640];
assign t[8641] = t[8640] ^ n[8641];
assign t[8642] = t[8641] ^ n[8642];
assign t[8643] = t[8642] ^ n[8643];
assign t[8644] = t[8643] ^ n[8644];
assign t[8645] = t[8644] ^ n[8645];
assign t[8646] = t[8645] ^ n[8646];
assign t[8647] = t[8646] ^ n[8647];
assign t[8648] = t[8647] ^ n[8648];
assign t[8649] = t[8648] ^ n[8649];
assign t[8650] = t[8649] ^ n[8650];
assign t[8651] = t[8650] ^ n[8651];
assign t[8652] = t[8651] ^ n[8652];
assign t[8653] = t[8652] ^ n[8653];
assign t[8654] = t[8653] ^ n[8654];
assign t[8655] = t[8654] ^ n[8655];
assign t[8656] = t[8655] ^ n[8656];
assign t[8657] = t[8656] ^ n[8657];
assign t[8658] = t[8657] ^ n[8658];
assign t[8659] = t[8658] ^ n[8659];
assign t[8660] = t[8659] ^ n[8660];
assign t[8661] = t[8660] ^ n[8661];
assign t[8662] = t[8661] ^ n[8662];
assign t[8663] = t[8662] ^ n[8663];
assign t[8664] = t[8663] ^ n[8664];
assign t[8665] = t[8664] ^ n[8665];
assign t[8666] = t[8665] ^ n[8666];
assign t[8667] = t[8666] ^ n[8667];
assign t[8668] = t[8667] ^ n[8668];
assign t[8669] = t[8668] ^ n[8669];
assign t[8670] = t[8669] ^ n[8670];
assign t[8671] = t[8670] ^ n[8671];
assign t[8672] = t[8671] ^ n[8672];
assign t[8673] = t[8672] ^ n[8673];
assign t[8674] = t[8673] ^ n[8674];
assign t[8675] = t[8674] ^ n[8675];
assign t[8676] = t[8675] ^ n[8676];
assign t[8677] = t[8676] ^ n[8677];
assign t[8678] = t[8677] ^ n[8678];
assign t[8679] = t[8678] ^ n[8679];
assign t[8680] = t[8679] ^ n[8680];
assign t[8681] = t[8680] ^ n[8681];
assign t[8682] = t[8681] ^ n[8682];
assign t[8683] = t[8682] ^ n[8683];
assign t[8684] = t[8683] ^ n[8684];
assign t[8685] = t[8684] ^ n[8685];
assign t[8686] = t[8685] ^ n[8686];
assign t[8687] = t[8686] ^ n[8687];
assign t[8688] = t[8687] ^ n[8688];
assign t[8689] = t[8688] ^ n[8689];
assign t[8690] = t[8689] ^ n[8690];
assign t[8691] = t[8690] ^ n[8691];
assign t[8692] = t[8691] ^ n[8692];
assign t[8693] = t[8692] ^ n[8693];
assign t[8694] = t[8693] ^ n[8694];
assign t[8695] = t[8694] ^ n[8695];
assign t[8696] = t[8695] ^ n[8696];
assign t[8697] = t[8696] ^ n[8697];
assign t[8698] = t[8697] ^ n[8698];
assign t[8699] = t[8698] ^ n[8699];
assign t[8700] = t[8699] ^ n[8700];
assign t[8701] = t[8700] ^ n[8701];
assign t[8702] = t[8701] ^ n[8702];
assign t[8703] = t[8702] ^ n[8703];
assign t[8704] = t[8703] ^ n[8704];
assign t[8705] = t[8704] ^ n[8705];
assign t[8706] = t[8705] ^ n[8706];
assign t[8707] = t[8706] ^ n[8707];
assign t[8708] = t[8707] ^ n[8708];
assign t[8709] = t[8708] ^ n[8709];
assign t[8710] = t[8709] ^ n[8710];
assign t[8711] = t[8710] ^ n[8711];
assign t[8712] = t[8711] ^ n[8712];
assign t[8713] = t[8712] ^ n[8713];
assign t[8714] = t[8713] ^ n[8714];
assign t[8715] = t[8714] ^ n[8715];
assign t[8716] = t[8715] ^ n[8716];
assign t[8717] = t[8716] ^ n[8717];
assign t[8718] = t[8717] ^ n[8718];
assign t[8719] = t[8718] ^ n[8719];
assign t[8720] = t[8719] ^ n[8720];
assign t[8721] = t[8720] ^ n[8721];
assign t[8722] = t[8721] ^ n[8722];
assign t[8723] = t[8722] ^ n[8723];
assign t[8724] = t[8723] ^ n[8724];
assign t[8725] = t[8724] ^ n[8725];
assign t[8726] = t[8725] ^ n[8726];
assign t[8727] = t[8726] ^ n[8727];
assign t[8728] = t[8727] ^ n[8728];
assign t[8729] = t[8728] ^ n[8729];
assign t[8730] = t[8729] ^ n[8730];
assign t[8731] = t[8730] ^ n[8731];
assign t[8732] = t[8731] ^ n[8732];
assign t[8733] = t[8732] ^ n[8733];
assign t[8734] = t[8733] ^ n[8734];
assign t[8735] = t[8734] ^ n[8735];
assign t[8736] = t[8735] ^ n[8736];
assign t[8737] = t[8736] ^ n[8737];
assign t[8738] = t[8737] ^ n[8738];
assign t[8739] = t[8738] ^ n[8739];
assign t[8740] = t[8739] ^ n[8740];
assign t[8741] = t[8740] ^ n[8741];
assign t[8742] = t[8741] ^ n[8742];
assign t[8743] = t[8742] ^ n[8743];
assign t[8744] = t[8743] ^ n[8744];
assign t[8745] = t[8744] ^ n[8745];
assign t[8746] = t[8745] ^ n[8746];
assign t[8747] = t[8746] ^ n[8747];
assign t[8748] = t[8747] ^ n[8748];
assign t[8749] = t[8748] ^ n[8749];
assign t[8750] = t[8749] ^ n[8750];
assign t[8751] = t[8750] ^ n[8751];
assign t[8752] = t[8751] ^ n[8752];
assign t[8753] = t[8752] ^ n[8753];
assign t[8754] = t[8753] ^ n[8754];
assign t[8755] = t[8754] ^ n[8755];
assign t[8756] = t[8755] ^ n[8756];
assign t[8757] = t[8756] ^ n[8757];
assign t[8758] = t[8757] ^ n[8758];
assign t[8759] = t[8758] ^ n[8759];
assign t[8760] = t[8759] ^ n[8760];
assign t[8761] = t[8760] ^ n[8761];
assign t[8762] = t[8761] ^ n[8762];
assign t[8763] = t[8762] ^ n[8763];
assign t[8764] = t[8763] ^ n[8764];
assign t[8765] = t[8764] ^ n[8765];
assign t[8766] = t[8765] ^ n[8766];
assign t[8767] = t[8766] ^ n[8767];
assign t[8768] = t[8767] ^ n[8768];
assign t[8769] = t[8768] ^ n[8769];
assign t[8770] = t[8769] ^ n[8770];
assign t[8771] = t[8770] ^ n[8771];
assign t[8772] = t[8771] ^ n[8772];
assign t[8773] = t[8772] ^ n[8773];
assign t[8774] = t[8773] ^ n[8774];
assign t[8775] = t[8774] ^ n[8775];
assign t[8776] = t[8775] ^ n[8776];
assign t[8777] = t[8776] ^ n[8777];
assign t[8778] = t[8777] ^ n[8778];
assign t[8779] = t[8778] ^ n[8779];
assign t[8780] = t[8779] ^ n[8780];
assign t[8781] = t[8780] ^ n[8781];
assign t[8782] = t[8781] ^ n[8782];
assign t[8783] = t[8782] ^ n[8783];
assign t[8784] = t[8783] ^ n[8784];
assign t[8785] = t[8784] ^ n[8785];
assign t[8786] = t[8785] ^ n[8786];
assign t[8787] = t[8786] ^ n[8787];
assign t[8788] = t[8787] ^ n[8788];
assign t[8789] = t[8788] ^ n[8789];
assign t[8790] = t[8789] ^ n[8790];
assign t[8791] = t[8790] ^ n[8791];
assign t[8792] = t[8791] ^ n[8792];
assign t[8793] = t[8792] ^ n[8793];
assign t[8794] = t[8793] ^ n[8794];
assign t[8795] = t[8794] ^ n[8795];
assign t[8796] = t[8795] ^ n[8796];
assign t[8797] = t[8796] ^ n[8797];
assign t[8798] = t[8797] ^ n[8798];
assign t[8799] = t[8798] ^ n[8799];
assign t[8800] = t[8799] ^ n[8800];
assign t[8801] = t[8800] ^ n[8801];
assign t[8802] = t[8801] ^ n[8802];
assign t[8803] = t[8802] ^ n[8803];
assign t[8804] = t[8803] ^ n[8804];
assign t[8805] = t[8804] ^ n[8805];
assign t[8806] = t[8805] ^ n[8806];
assign t[8807] = t[8806] ^ n[8807];
assign t[8808] = t[8807] ^ n[8808];
assign t[8809] = t[8808] ^ n[8809];
assign t[8810] = t[8809] ^ n[8810];
assign t[8811] = t[8810] ^ n[8811];
assign t[8812] = t[8811] ^ n[8812];
assign t[8813] = t[8812] ^ n[8813];
assign t[8814] = t[8813] ^ n[8814];
assign t[8815] = t[8814] ^ n[8815];
assign t[8816] = t[8815] ^ n[8816];
assign t[8817] = t[8816] ^ n[8817];
assign t[8818] = t[8817] ^ n[8818];
assign t[8819] = t[8818] ^ n[8819];
assign t[8820] = t[8819] ^ n[8820];
assign t[8821] = t[8820] ^ n[8821];
assign t[8822] = t[8821] ^ n[8822];
assign t[8823] = t[8822] ^ n[8823];
assign t[8824] = t[8823] ^ n[8824];
assign t[8825] = t[8824] ^ n[8825];
assign t[8826] = t[8825] ^ n[8826];
assign t[8827] = t[8826] ^ n[8827];
assign t[8828] = t[8827] ^ n[8828];
assign t[8829] = t[8828] ^ n[8829];
assign t[8830] = t[8829] ^ n[8830];
assign t[8831] = t[8830] ^ n[8831];
assign t[8832] = t[8831] ^ n[8832];
assign t[8833] = t[8832] ^ n[8833];
assign t[8834] = t[8833] ^ n[8834];
assign t[8835] = t[8834] ^ n[8835];
assign t[8836] = t[8835] ^ n[8836];
assign t[8837] = t[8836] ^ n[8837];
assign t[8838] = t[8837] ^ n[8838];
assign t[8839] = t[8838] ^ n[8839];
assign t[8840] = t[8839] ^ n[8840];
assign t[8841] = t[8840] ^ n[8841];
assign t[8842] = t[8841] ^ n[8842];
assign t[8843] = t[8842] ^ n[8843];
assign t[8844] = t[8843] ^ n[8844];
assign t[8845] = t[8844] ^ n[8845];
assign t[8846] = t[8845] ^ n[8846];
assign t[8847] = t[8846] ^ n[8847];
assign t[8848] = t[8847] ^ n[8848];
assign t[8849] = t[8848] ^ n[8849];
assign t[8850] = t[8849] ^ n[8850];
assign t[8851] = t[8850] ^ n[8851];
assign t[8852] = t[8851] ^ n[8852];
assign t[8853] = t[8852] ^ n[8853];
assign t[8854] = t[8853] ^ n[8854];
assign t[8855] = t[8854] ^ n[8855];
assign t[8856] = t[8855] ^ n[8856];
assign t[8857] = t[8856] ^ n[8857];
assign t[8858] = t[8857] ^ n[8858];
assign t[8859] = t[8858] ^ n[8859];
assign t[8860] = t[8859] ^ n[8860];
assign t[8861] = t[8860] ^ n[8861];
assign t[8862] = t[8861] ^ n[8862];
assign t[8863] = t[8862] ^ n[8863];
assign t[8864] = t[8863] ^ n[8864];
assign t[8865] = t[8864] ^ n[8865];
assign t[8866] = t[8865] ^ n[8866];
assign t[8867] = t[8866] ^ n[8867];
assign t[8868] = t[8867] ^ n[8868];
assign t[8869] = t[8868] ^ n[8869];
assign t[8870] = t[8869] ^ n[8870];
assign t[8871] = t[8870] ^ n[8871];
assign t[8872] = t[8871] ^ n[8872];
assign t[8873] = t[8872] ^ n[8873];
assign t[8874] = t[8873] ^ n[8874];
assign t[8875] = t[8874] ^ n[8875];
assign t[8876] = t[8875] ^ n[8876];
assign t[8877] = t[8876] ^ n[8877];
assign t[8878] = t[8877] ^ n[8878];
assign t[8879] = t[8878] ^ n[8879];
assign t[8880] = t[8879] ^ n[8880];
assign t[8881] = t[8880] ^ n[8881];
assign t[8882] = t[8881] ^ n[8882];
assign t[8883] = t[8882] ^ n[8883];
assign t[8884] = t[8883] ^ n[8884];
assign t[8885] = t[8884] ^ n[8885];
assign t[8886] = t[8885] ^ n[8886];
assign t[8887] = t[8886] ^ n[8887];
assign t[8888] = t[8887] ^ n[8888];
assign t[8889] = t[8888] ^ n[8889];
assign t[8890] = t[8889] ^ n[8890];
assign t[8891] = t[8890] ^ n[8891];
assign t[8892] = t[8891] ^ n[8892];
assign t[8893] = t[8892] ^ n[8893];
assign t[8894] = t[8893] ^ n[8894];
assign t[8895] = t[8894] ^ n[8895];
assign t[8896] = t[8895] ^ n[8896];
assign t[8897] = t[8896] ^ n[8897];
assign t[8898] = t[8897] ^ n[8898];
assign t[8899] = t[8898] ^ n[8899];
assign t[8900] = t[8899] ^ n[8900];
assign t[8901] = t[8900] ^ n[8901];
assign t[8902] = t[8901] ^ n[8902];
assign t[8903] = t[8902] ^ n[8903];
assign t[8904] = t[8903] ^ n[8904];
assign t[8905] = t[8904] ^ n[8905];
assign t[8906] = t[8905] ^ n[8906];
assign t[8907] = t[8906] ^ n[8907];
assign t[8908] = t[8907] ^ n[8908];
assign t[8909] = t[8908] ^ n[8909];
assign t[8910] = t[8909] ^ n[8910];
assign t[8911] = t[8910] ^ n[8911];
assign t[8912] = t[8911] ^ n[8912];
assign t[8913] = t[8912] ^ n[8913];
assign t[8914] = t[8913] ^ n[8914];
assign t[8915] = t[8914] ^ n[8915];
assign t[8916] = t[8915] ^ n[8916];
assign t[8917] = t[8916] ^ n[8917];
assign t[8918] = t[8917] ^ n[8918];
assign t[8919] = t[8918] ^ n[8919];
assign t[8920] = t[8919] ^ n[8920];
assign t[8921] = t[8920] ^ n[8921];
assign t[8922] = t[8921] ^ n[8922];
assign t[8923] = t[8922] ^ n[8923];
assign t[8924] = t[8923] ^ n[8924];
assign t[8925] = t[8924] ^ n[8925];
assign t[8926] = t[8925] ^ n[8926];
assign t[8927] = t[8926] ^ n[8927];
assign t[8928] = t[8927] ^ n[8928];
assign t[8929] = t[8928] ^ n[8929];
assign t[8930] = t[8929] ^ n[8930];
assign t[8931] = t[8930] ^ n[8931];
assign t[8932] = t[8931] ^ n[8932];
assign t[8933] = t[8932] ^ n[8933];
assign t[8934] = t[8933] ^ n[8934];
assign t[8935] = t[8934] ^ n[8935];
assign t[8936] = t[8935] ^ n[8936];
assign t[8937] = t[8936] ^ n[8937];
assign t[8938] = t[8937] ^ n[8938];
assign t[8939] = t[8938] ^ n[8939];
assign t[8940] = t[8939] ^ n[8940];
assign t[8941] = t[8940] ^ n[8941];
assign t[8942] = t[8941] ^ n[8942];
assign t[8943] = t[8942] ^ n[8943];
assign t[8944] = t[8943] ^ n[8944];
assign t[8945] = t[8944] ^ n[8945];
assign t[8946] = t[8945] ^ n[8946];
assign t[8947] = t[8946] ^ n[8947];
assign t[8948] = t[8947] ^ n[8948];
assign t[8949] = t[8948] ^ n[8949];
assign t[8950] = t[8949] ^ n[8950];
assign t[8951] = t[8950] ^ n[8951];
assign t[8952] = t[8951] ^ n[8952];
assign t[8953] = t[8952] ^ n[8953];
assign t[8954] = t[8953] ^ n[8954];
assign t[8955] = t[8954] ^ n[8955];
assign t[8956] = t[8955] ^ n[8956];
assign t[8957] = t[8956] ^ n[8957];
assign t[8958] = t[8957] ^ n[8958];
assign t[8959] = t[8958] ^ n[8959];
assign t[8960] = t[8959] ^ n[8960];
assign t[8961] = t[8960] ^ n[8961];
assign t[8962] = t[8961] ^ n[8962];
assign t[8963] = t[8962] ^ n[8963];
assign t[8964] = t[8963] ^ n[8964];
assign t[8965] = t[8964] ^ n[8965];
assign t[8966] = t[8965] ^ n[8966];
assign t[8967] = t[8966] ^ n[8967];
assign t[8968] = t[8967] ^ n[8968];
assign t[8969] = t[8968] ^ n[8969];
assign t[8970] = t[8969] ^ n[8970];
assign t[8971] = t[8970] ^ n[8971];
assign t[8972] = t[8971] ^ n[8972];
assign t[8973] = t[8972] ^ n[8973];
assign t[8974] = t[8973] ^ n[8974];
assign t[8975] = t[8974] ^ n[8975];
assign t[8976] = t[8975] ^ n[8976];
assign t[8977] = t[8976] ^ n[8977];
assign t[8978] = t[8977] ^ n[8978];
assign t[8979] = t[8978] ^ n[8979];
assign t[8980] = t[8979] ^ n[8980];
assign t[8981] = t[8980] ^ n[8981];
assign t[8982] = t[8981] ^ n[8982];
assign t[8983] = t[8982] ^ n[8983];
assign t[8984] = t[8983] ^ n[8984];
assign t[8985] = t[8984] ^ n[8985];
assign t[8986] = t[8985] ^ n[8986];
assign t[8987] = t[8986] ^ n[8987];
assign t[8988] = t[8987] ^ n[8988];
assign t[8989] = t[8988] ^ n[8989];
assign t[8990] = t[8989] ^ n[8990];
assign t[8991] = t[8990] ^ n[8991];
assign t[8992] = t[8991] ^ n[8992];
assign t[8993] = t[8992] ^ n[8993];
assign t[8994] = t[8993] ^ n[8994];
assign t[8995] = t[8994] ^ n[8995];
assign t[8996] = t[8995] ^ n[8996];
assign t[8997] = t[8996] ^ n[8997];
assign t[8998] = t[8997] ^ n[8998];
assign t[8999] = t[8998] ^ n[8999];
assign t[9000] = t[8999] ^ n[9000];
assign t[9001] = t[9000] ^ n[9001];
assign t[9002] = t[9001] ^ n[9002];
assign t[9003] = t[9002] ^ n[9003];
assign t[9004] = t[9003] ^ n[9004];
assign t[9005] = t[9004] ^ n[9005];
assign t[9006] = t[9005] ^ n[9006];
assign t[9007] = t[9006] ^ n[9007];
assign t[9008] = t[9007] ^ n[9008];
assign t[9009] = t[9008] ^ n[9009];
assign t[9010] = t[9009] ^ n[9010];
assign t[9011] = t[9010] ^ n[9011];
assign t[9012] = t[9011] ^ n[9012];
assign t[9013] = t[9012] ^ n[9013];
assign t[9014] = t[9013] ^ n[9014];
assign t[9015] = t[9014] ^ n[9015];
assign t[9016] = t[9015] ^ n[9016];
assign t[9017] = t[9016] ^ n[9017];
assign t[9018] = t[9017] ^ n[9018];
assign t[9019] = t[9018] ^ n[9019];
assign t[9020] = t[9019] ^ n[9020];
assign t[9021] = t[9020] ^ n[9021];
assign t[9022] = t[9021] ^ n[9022];
assign t[9023] = t[9022] ^ n[9023];
assign t[9024] = t[9023] ^ n[9024];
assign t[9025] = t[9024] ^ n[9025];
assign t[9026] = t[9025] ^ n[9026];
assign t[9027] = t[9026] ^ n[9027];
assign t[9028] = t[9027] ^ n[9028];
assign t[9029] = t[9028] ^ n[9029];
assign t[9030] = t[9029] ^ n[9030];
assign t[9031] = t[9030] ^ n[9031];
assign t[9032] = t[9031] ^ n[9032];
assign t[9033] = t[9032] ^ n[9033];
assign t[9034] = t[9033] ^ n[9034];
assign t[9035] = t[9034] ^ n[9035];
assign t[9036] = t[9035] ^ n[9036];
assign t[9037] = t[9036] ^ n[9037];
assign t[9038] = t[9037] ^ n[9038];
assign t[9039] = t[9038] ^ n[9039];
assign t[9040] = t[9039] ^ n[9040];
assign t[9041] = t[9040] ^ n[9041];
assign t[9042] = t[9041] ^ n[9042];
assign t[9043] = t[9042] ^ n[9043];
assign t[9044] = t[9043] ^ n[9044];
assign t[9045] = t[9044] ^ n[9045];
assign t[9046] = t[9045] ^ n[9046];
assign t[9047] = t[9046] ^ n[9047];
assign t[9048] = t[9047] ^ n[9048];
assign t[9049] = t[9048] ^ n[9049];
assign t[9050] = t[9049] ^ n[9050];
assign t[9051] = t[9050] ^ n[9051];
assign t[9052] = t[9051] ^ n[9052];
assign t[9053] = t[9052] ^ n[9053];
assign t[9054] = t[9053] ^ n[9054];
assign t[9055] = t[9054] ^ n[9055];
assign t[9056] = t[9055] ^ n[9056];
assign t[9057] = t[9056] ^ n[9057];
assign t[9058] = t[9057] ^ n[9058];
assign t[9059] = t[9058] ^ n[9059];
assign t[9060] = t[9059] ^ n[9060];
assign t[9061] = t[9060] ^ n[9061];
assign t[9062] = t[9061] ^ n[9062];
assign t[9063] = t[9062] ^ n[9063];
assign t[9064] = t[9063] ^ n[9064];
assign t[9065] = t[9064] ^ n[9065];
assign t[9066] = t[9065] ^ n[9066];
assign t[9067] = t[9066] ^ n[9067];
assign t[9068] = t[9067] ^ n[9068];
assign t[9069] = t[9068] ^ n[9069];
assign t[9070] = t[9069] ^ n[9070];
assign t[9071] = t[9070] ^ n[9071];
assign t[9072] = t[9071] ^ n[9072];
assign t[9073] = t[9072] ^ n[9073];
assign t[9074] = t[9073] ^ n[9074];
assign t[9075] = t[9074] ^ n[9075];
assign t[9076] = t[9075] ^ n[9076];
assign t[9077] = t[9076] ^ n[9077];
assign t[9078] = t[9077] ^ n[9078];
assign t[9079] = t[9078] ^ n[9079];
assign t[9080] = t[9079] ^ n[9080];
assign t[9081] = t[9080] ^ n[9081];
assign t[9082] = t[9081] ^ n[9082];
assign t[9083] = t[9082] ^ n[9083];
assign t[9084] = t[9083] ^ n[9084];
assign t[9085] = t[9084] ^ n[9085];
assign t[9086] = t[9085] ^ n[9086];
assign t[9087] = t[9086] ^ n[9087];
assign t[9088] = t[9087] ^ n[9088];
assign t[9089] = t[9088] ^ n[9089];
assign t[9090] = t[9089] ^ n[9090];
assign t[9091] = t[9090] ^ n[9091];
assign t[9092] = t[9091] ^ n[9092];
assign t[9093] = t[9092] ^ n[9093];
assign t[9094] = t[9093] ^ n[9094];
assign t[9095] = t[9094] ^ n[9095];
assign t[9096] = t[9095] ^ n[9096];
assign t[9097] = t[9096] ^ n[9097];
assign t[9098] = t[9097] ^ n[9098];
assign t[9099] = t[9098] ^ n[9099];
assign t[9100] = t[9099] ^ n[9100];
assign t[9101] = t[9100] ^ n[9101];
assign t[9102] = t[9101] ^ n[9102];
assign t[9103] = t[9102] ^ n[9103];
assign t[9104] = t[9103] ^ n[9104];
assign t[9105] = t[9104] ^ n[9105];
assign t[9106] = t[9105] ^ n[9106];
assign t[9107] = t[9106] ^ n[9107];
assign t[9108] = t[9107] ^ n[9108];
assign t[9109] = t[9108] ^ n[9109];
assign t[9110] = t[9109] ^ n[9110];
assign t[9111] = t[9110] ^ n[9111];
assign t[9112] = t[9111] ^ n[9112];
assign t[9113] = t[9112] ^ n[9113];
assign t[9114] = t[9113] ^ n[9114];
assign t[9115] = t[9114] ^ n[9115];
assign t[9116] = t[9115] ^ n[9116];
assign t[9117] = t[9116] ^ n[9117];
assign t[9118] = t[9117] ^ n[9118];
assign t[9119] = t[9118] ^ n[9119];
assign t[9120] = t[9119] ^ n[9120];
assign t[9121] = t[9120] ^ n[9121];
assign t[9122] = t[9121] ^ n[9122];
assign t[9123] = t[9122] ^ n[9123];
assign t[9124] = t[9123] ^ n[9124];
assign t[9125] = t[9124] ^ n[9125];
assign t[9126] = t[9125] ^ n[9126];
assign t[9127] = t[9126] ^ n[9127];
assign t[9128] = t[9127] ^ n[9128];
assign t[9129] = t[9128] ^ n[9129];
assign t[9130] = t[9129] ^ n[9130];
assign t[9131] = t[9130] ^ n[9131];
assign t[9132] = t[9131] ^ n[9132];
assign t[9133] = t[9132] ^ n[9133];
assign t[9134] = t[9133] ^ n[9134];
assign t[9135] = t[9134] ^ n[9135];
assign t[9136] = t[9135] ^ n[9136];
assign t[9137] = t[9136] ^ n[9137];
assign t[9138] = t[9137] ^ n[9138];
assign t[9139] = t[9138] ^ n[9139];
assign t[9140] = t[9139] ^ n[9140];
assign t[9141] = t[9140] ^ n[9141];
assign t[9142] = t[9141] ^ n[9142];
assign t[9143] = t[9142] ^ n[9143];
assign t[9144] = t[9143] ^ n[9144];
assign t[9145] = t[9144] ^ n[9145];
assign t[9146] = t[9145] ^ n[9146];
assign t[9147] = t[9146] ^ n[9147];
assign t[9148] = t[9147] ^ n[9148];
assign t[9149] = t[9148] ^ n[9149];
assign t[9150] = t[9149] ^ n[9150];
assign t[9151] = t[9150] ^ n[9151];
assign t[9152] = t[9151] ^ n[9152];
assign t[9153] = t[9152] ^ n[9153];
assign t[9154] = t[9153] ^ n[9154];
assign t[9155] = t[9154] ^ n[9155];
assign t[9156] = t[9155] ^ n[9156];
assign t[9157] = t[9156] ^ n[9157];
assign t[9158] = t[9157] ^ n[9158];
assign t[9159] = t[9158] ^ n[9159];
assign t[9160] = t[9159] ^ n[9160];
assign t[9161] = t[9160] ^ n[9161];
assign t[9162] = t[9161] ^ n[9162];
assign t[9163] = t[9162] ^ n[9163];
assign t[9164] = t[9163] ^ n[9164];
assign t[9165] = t[9164] ^ n[9165];
assign t[9166] = t[9165] ^ n[9166];
assign t[9167] = t[9166] ^ n[9167];
assign t[9168] = t[9167] ^ n[9168];
assign t[9169] = t[9168] ^ n[9169];
assign t[9170] = t[9169] ^ n[9170];
assign t[9171] = t[9170] ^ n[9171];
assign t[9172] = t[9171] ^ n[9172];
assign t[9173] = t[9172] ^ n[9173];
assign t[9174] = t[9173] ^ n[9174];
assign t[9175] = t[9174] ^ n[9175];
assign t[9176] = t[9175] ^ n[9176];
assign t[9177] = t[9176] ^ n[9177];
assign t[9178] = t[9177] ^ n[9178];
assign t[9179] = t[9178] ^ n[9179];
assign t[9180] = t[9179] ^ n[9180];
assign t[9181] = t[9180] ^ n[9181];
assign t[9182] = t[9181] ^ n[9182];
assign t[9183] = t[9182] ^ n[9183];
assign t[9184] = t[9183] ^ n[9184];
assign t[9185] = t[9184] ^ n[9185];
assign t[9186] = t[9185] ^ n[9186];
assign t[9187] = t[9186] ^ n[9187];
assign t[9188] = t[9187] ^ n[9188];
assign t[9189] = t[9188] ^ n[9189];
assign t[9190] = t[9189] ^ n[9190];
assign t[9191] = t[9190] ^ n[9191];
assign t[9192] = t[9191] ^ n[9192];
assign t[9193] = t[9192] ^ n[9193];
assign t[9194] = t[9193] ^ n[9194];
assign t[9195] = t[9194] ^ n[9195];
assign t[9196] = t[9195] ^ n[9196];
assign t[9197] = t[9196] ^ n[9197];
assign t[9198] = t[9197] ^ n[9198];
assign t[9199] = t[9198] ^ n[9199];
assign t[9200] = t[9199] ^ n[9200];
assign t[9201] = t[9200] ^ n[9201];
assign t[9202] = t[9201] ^ n[9202];
assign t[9203] = t[9202] ^ n[9203];
assign t[9204] = t[9203] ^ n[9204];
assign t[9205] = t[9204] ^ n[9205];
assign t[9206] = t[9205] ^ n[9206];
assign t[9207] = t[9206] ^ n[9207];
assign t[9208] = t[9207] ^ n[9208];
assign t[9209] = t[9208] ^ n[9209];
assign t[9210] = t[9209] ^ n[9210];
assign t[9211] = t[9210] ^ n[9211];
assign t[9212] = t[9211] ^ n[9212];
assign t[9213] = t[9212] ^ n[9213];
assign t[9214] = t[9213] ^ n[9214];
assign t[9215] = t[9214] ^ n[9215];
assign t[9216] = t[9215] ^ n[9216];
assign t[9217] = t[9216] ^ n[9217];
assign t[9218] = t[9217] ^ n[9218];
assign t[9219] = t[9218] ^ n[9219];
assign t[9220] = t[9219] ^ n[9220];
assign t[9221] = t[9220] ^ n[9221];
assign t[9222] = t[9221] ^ n[9222];
assign t[9223] = t[9222] ^ n[9223];
assign t[9224] = t[9223] ^ n[9224];
assign t[9225] = t[9224] ^ n[9225];
assign t[9226] = t[9225] ^ n[9226];
assign t[9227] = t[9226] ^ n[9227];
assign t[9228] = t[9227] ^ n[9228];
assign t[9229] = t[9228] ^ n[9229];
assign t[9230] = t[9229] ^ n[9230];
assign t[9231] = t[9230] ^ n[9231];
assign t[9232] = t[9231] ^ n[9232];
assign t[9233] = t[9232] ^ n[9233];
assign t[9234] = t[9233] ^ n[9234];
assign t[9235] = t[9234] ^ n[9235];
assign t[9236] = t[9235] ^ n[9236];
assign t[9237] = t[9236] ^ n[9237];
assign t[9238] = t[9237] ^ n[9238];
assign t[9239] = t[9238] ^ n[9239];
assign t[9240] = t[9239] ^ n[9240];
assign t[9241] = t[9240] ^ n[9241];
assign t[9242] = t[9241] ^ n[9242];
assign t[9243] = t[9242] ^ n[9243];
assign t[9244] = t[9243] ^ n[9244];
assign t[9245] = t[9244] ^ n[9245];
assign t[9246] = t[9245] ^ n[9246];
assign t[9247] = t[9246] ^ n[9247];
assign t[9248] = t[9247] ^ n[9248];
assign t[9249] = t[9248] ^ n[9249];
assign t[9250] = t[9249] ^ n[9250];
assign t[9251] = t[9250] ^ n[9251];
assign t[9252] = t[9251] ^ n[9252];
assign t[9253] = t[9252] ^ n[9253];
assign t[9254] = t[9253] ^ n[9254];
assign t[9255] = t[9254] ^ n[9255];
assign t[9256] = t[9255] ^ n[9256];
assign t[9257] = t[9256] ^ n[9257];
assign t[9258] = t[9257] ^ n[9258];
assign t[9259] = t[9258] ^ n[9259];
assign t[9260] = t[9259] ^ n[9260];
assign t[9261] = t[9260] ^ n[9261];
assign t[9262] = t[9261] ^ n[9262];
assign t[9263] = t[9262] ^ n[9263];
assign t[9264] = t[9263] ^ n[9264];
assign t[9265] = t[9264] ^ n[9265];
assign t[9266] = t[9265] ^ n[9266];
assign t[9267] = t[9266] ^ n[9267];
assign t[9268] = t[9267] ^ n[9268];
assign t[9269] = t[9268] ^ n[9269];
assign t[9270] = t[9269] ^ n[9270];
assign t[9271] = t[9270] ^ n[9271];
assign t[9272] = t[9271] ^ n[9272];
assign t[9273] = t[9272] ^ n[9273];
assign t[9274] = t[9273] ^ n[9274];
assign t[9275] = t[9274] ^ n[9275];
assign t[9276] = t[9275] ^ n[9276];
assign t[9277] = t[9276] ^ n[9277];
assign t[9278] = t[9277] ^ n[9278];
assign t[9279] = t[9278] ^ n[9279];
assign t[9280] = t[9279] ^ n[9280];
assign t[9281] = t[9280] ^ n[9281];
assign t[9282] = t[9281] ^ n[9282];
assign t[9283] = t[9282] ^ n[9283];
assign t[9284] = t[9283] ^ n[9284];
assign t[9285] = t[9284] ^ n[9285];
assign t[9286] = t[9285] ^ n[9286];
assign t[9287] = t[9286] ^ n[9287];
assign t[9288] = t[9287] ^ n[9288];
assign t[9289] = t[9288] ^ n[9289];
assign t[9290] = t[9289] ^ n[9290];
assign t[9291] = t[9290] ^ n[9291];
assign t[9292] = t[9291] ^ n[9292];
assign t[9293] = t[9292] ^ n[9293];
assign t[9294] = t[9293] ^ n[9294];
assign t[9295] = t[9294] ^ n[9295];
assign t[9296] = t[9295] ^ n[9296];
assign t[9297] = t[9296] ^ n[9297];
assign t[9298] = t[9297] ^ n[9298];
assign t[9299] = t[9298] ^ n[9299];
assign t[9300] = t[9299] ^ n[9300];
assign t[9301] = t[9300] ^ n[9301];
assign t[9302] = t[9301] ^ n[9302];
assign t[9303] = t[9302] ^ n[9303];
assign t[9304] = t[9303] ^ n[9304];
assign t[9305] = t[9304] ^ n[9305];
assign t[9306] = t[9305] ^ n[9306];
assign t[9307] = t[9306] ^ n[9307];
assign t[9308] = t[9307] ^ n[9308];
assign t[9309] = t[9308] ^ n[9309];
assign t[9310] = t[9309] ^ n[9310];
assign t[9311] = t[9310] ^ n[9311];
assign t[9312] = t[9311] ^ n[9312];
assign t[9313] = t[9312] ^ n[9313];
assign t[9314] = t[9313] ^ n[9314];
assign t[9315] = t[9314] ^ n[9315];
assign t[9316] = t[9315] ^ n[9316];
assign t[9317] = t[9316] ^ n[9317];
assign t[9318] = t[9317] ^ n[9318];
assign t[9319] = t[9318] ^ n[9319];
assign t[9320] = t[9319] ^ n[9320];
assign t[9321] = t[9320] ^ n[9321];
assign t[9322] = t[9321] ^ n[9322];
assign t[9323] = t[9322] ^ n[9323];
assign t[9324] = t[9323] ^ n[9324];
assign t[9325] = t[9324] ^ n[9325];
assign t[9326] = t[9325] ^ n[9326];
assign t[9327] = t[9326] ^ n[9327];
assign t[9328] = t[9327] ^ n[9328];
assign t[9329] = t[9328] ^ n[9329];
assign t[9330] = t[9329] ^ n[9330];
assign t[9331] = t[9330] ^ n[9331];
assign t[9332] = t[9331] ^ n[9332];
assign t[9333] = t[9332] ^ n[9333];
assign t[9334] = t[9333] ^ n[9334];
assign t[9335] = t[9334] ^ n[9335];
assign t[9336] = t[9335] ^ n[9336];
assign t[9337] = t[9336] ^ n[9337];
assign t[9338] = t[9337] ^ n[9338];
assign t[9339] = t[9338] ^ n[9339];
assign t[9340] = t[9339] ^ n[9340];
assign t[9341] = t[9340] ^ n[9341];
assign t[9342] = t[9341] ^ n[9342];
assign t[9343] = t[9342] ^ n[9343];
assign t[9344] = t[9343] ^ n[9344];
assign t[9345] = t[9344] ^ n[9345];
assign t[9346] = t[9345] ^ n[9346];
assign t[9347] = t[9346] ^ n[9347];
assign t[9348] = t[9347] ^ n[9348];
assign t[9349] = t[9348] ^ n[9349];
assign t[9350] = t[9349] ^ n[9350];
assign t[9351] = t[9350] ^ n[9351];
assign t[9352] = t[9351] ^ n[9352];
assign t[9353] = t[9352] ^ n[9353];
assign t[9354] = t[9353] ^ n[9354];
assign t[9355] = t[9354] ^ n[9355];
assign t[9356] = t[9355] ^ n[9356];
assign t[9357] = t[9356] ^ n[9357];
assign t[9358] = t[9357] ^ n[9358];
assign t[9359] = t[9358] ^ n[9359];
assign t[9360] = t[9359] ^ n[9360];
assign t[9361] = t[9360] ^ n[9361];
assign t[9362] = t[9361] ^ n[9362];
assign t[9363] = t[9362] ^ n[9363];
assign t[9364] = t[9363] ^ n[9364];
assign t[9365] = t[9364] ^ n[9365];
assign t[9366] = t[9365] ^ n[9366];
assign t[9367] = t[9366] ^ n[9367];
assign t[9368] = t[9367] ^ n[9368];
assign t[9369] = t[9368] ^ n[9369];
assign t[9370] = t[9369] ^ n[9370];
assign t[9371] = t[9370] ^ n[9371];
assign t[9372] = t[9371] ^ n[9372];
assign t[9373] = t[9372] ^ n[9373];
assign t[9374] = t[9373] ^ n[9374];
assign t[9375] = t[9374] ^ n[9375];
assign t[9376] = t[9375] ^ n[9376];
assign t[9377] = t[9376] ^ n[9377];
assign t[9378] = t[9377] ^ n[9378];
assign t[9379] = t[9378] ^ n[9379];
assign t[9380] = t[9379] ^ n[9380];
assign t[9381] = t[9380] ^ n[9381];
assign t[9382] = t[9381] ^ n[9382];
assign t[9383] = t[9382] ^ n[9383];
assign t[9384] = t[9383] ^ n[9384];
assign t[9385] = t[9384] ^ n[9385];
assign t[9386] = t[9385] ^ n[9386];
assign t[9387] = t[9386] ^ n[9387];
assign t[9388] = t[9387] ^ n[9388];
assign t[9389] = t[9388] ^ n[9389];
assign t[9390] = t[9389] ^ n[9390];
assign t[9391] = t[9390] ^ n[9391];
assign t[9392] = t[9391] ^ n[9392];
assign t[9393] = t[9392] ^ n[9393];
assign t[9394] = t[9393] ^ n[9394];
assign t[9395] = t[9394] ^ n[9395];
assign t[9396] = t[9395] ^ n[9396];
assign t[9397] = t[9396] ^ n[9397];
assign t[9398] = t[9397] ^ n[9398];
assign t[9399] = t[9398] ^ n[9399];
assign t[9400] = t[9399] ^ n[9400];
assign t[9401] = t[9400] ^ n[9401];
assign t[9402] = t[9401] ^ n[9402];
assign t[9403] = t[9402] ^ n[9403];
assign t[9404] = t[9403] ^ n[9404];
assign t[9405] = t[9404] ^ n[9405];
assign t[9406] = t[9405] ^ n[9406];
assign t[9407] = t[9406] ^ n[9407];
assign t[9408] = t[9407] ^ n[9408];
assign t[9409] = t[9408] ^ n[9409];
assign t[9410] = t[9409] ^ n[9410];
assign t[9411] = t[9410] ^ n[9411];
assign t[9412] = t[9411] ^ n[9412];
assign t[9413] = t[9412] ^ n[9413];
assign t[9414] = t[9413] ^ n[9414];
assign t[9415] = t[9414] ^ n[9415];
assign t[9416] = t[9415] ^ n[9416];
assign t[9417] = t[9416] ^ n[9417];
assign t[9418] = t[9417] ^ n[9418];
assign t[9419] = t[9418] ^ n[9419];
assign t[9420] = t[9419] ^ n[9420];
assign t[9421] = t[9420] ^ n[9421];
assign t[9422] = t[9421] ^ n[9422];
assign t[9423] = t[9422] ^ n[9423];
assign t[9424] = t[9423] ^ n[9424];
assign t[9425] = t[9424] ^ n[9425];
assign t[9426] = t[9425] ^ n[9426];
assign t[9427] = t[9426] ^ n[9427];
assign t[9428] = t[9427] ^ n[9428];
assign t[9429] = t[9428] ^ n[9429];
assign t[9430] = t[9429] ^ n[9430];
assign t[9431] = t[9430] ^ n[9431];
assign t[9432] = t[9431] ^ n[9432];
assign t[9433] = t[9432] ^ n[9433];
assign t[9434] = t[9433] ^ n[9434];
assign t[9435] = t[9434] ^ n[9435];
assign t[9436] = t[9435] ^ n[9436];
assign t[9437] = t[9436] ^ n[9437];
assign t[9438] = t[9437] ^ n[9438];
assign t[9439] = t[9438] ^ n[9439];
assign t[9440] = t[9439] ^ n[9440];
assign t[9441] = t[9440] ^ n[9441];
assign t[9442] = t[9441] ^ n[9442];
assign t[9443] = t[9442] ^ n[9443];
assign t[9444] = t[9443] ^ n[9444];
assign t[9445] = t[9444] ^ n[9445];
assign t[9446] = t[9445] ^ n[9446];
assign t[9447] = t[9446] ^ n[9447];
assign t[9448] = t[9447] ^ n[9448];
assign t[9449] = t[9448] ^ n[9449];
assign t[9450] = t[9449] ^ n[9450];
assign t[9451] = t[9450] ^ n[9451];
assign t[9452] = t[9451] ^ n[9452];
assign t[9453] = t[9452] ^ n[9453];
assign t[9454] = t[9453] ^ n[9454];
assign t[9455] = t[9454] ^ n[9455];
assign t[9456] = t[9455] ^ n[9456];
assign t[9457] = t[9456] ^ n[9457];
assign t[9458] = t[9457] ^ n[9458];
assign t[9459] = t[9458] ^ n[9459];
assign t[9460] = t[9459] ^ n[9460];
assign t[9461] = t[9460] ^ n[9461];
assign t[9462] = t[9461] ^ n[9462];
assign t[9463] = t[9462] ^ n[9463];
assign t[9464] = t[9463] ^ n[9464];
assign t[9465] = t[9464] ^ n[9465];
assign t[9466] = t[9465] ^ n[9466];
assign t[9467] = t[9466] ^ n[9467];
assign t[9468] = t[9467] ^ n[9468];
assign t[9469] = t[9468] ^ n[9469];
assign t[9470] = t[9469] ^ n[9470];
assign t[9471] = t[9470] ^ n[9471];
assign t[9472] = t[9471] ^ n[9472];
assign t[9473] = t[9472] ^ n[9473];
assign t[9474] = t[9473] ^ n[9474];
assign t[9475] = t[9474] ^ n[9475];
assign t[9476] = t[9475] ^ n[9476];
assign t[9477] = t[9476] ^ n[9477];
assign t[9478] = t[9477] ^ n[9478];
assign t[9479] = t[9478] ^ n[9479];
assign t[9480] = t[9479] ^ n[9480];
assign t[9481] = t[9480] ^ n[9481];
assign t[9482] = t[9481] ^ n[9482];
assign t[9483] = t[9482] ^ n[9483];
assign t[9484] = t[9483] ^ n[9484];
assign t[9485] = t[9484] ^ n[9485];
assign t[9486] = t[9485] ^ n[9486];
assign t[9487] = t[9486] ^ n[9487];
assign t[9488] = t[9487] ^ n[9488];
assign t[9489] = t[9488] ^ n[9489];
assign t[9490] = t[9489] ^ n[9490];
assign t[9491] = t[9490] ^ n[9491];
assign t[9492] = t[9491] ^ n[9492];
assign t[9493] = t[9492] ^ n[9493];
assign t[9494] = t[9493] ^ n[9494];
assign t[9495] = t[9494] ^ n[9495];
assign t[9496] = t[9495] ^ n[9496];
assign t[9497] = t[9496] ^ n[9497];
assign t[9498] = t[9497] ^ n[9498];
assign t[9499] = t[9498] ^ n[9499];
assign t[9500] = t[9499] ^ n[9500];
assign t[9501] = t[9500] ^ n[9501];
assign t[9502] = t[9501] ^ n[9502];
assign t[9503] = t[9502] ^ n[9503];
assign t[9504] = t[9503] ^ n[9504];
assign t[9505] = t[9504] ^ n[9505];
assign t[9506] = t[9505] ^ n[9506];
assign t[9507] = t[9506] ^ n[9507];
assign t[9508] = t[9507] ^ n[9508];
assign t[9509] = t[9508] ^ n[9509];
assign t[9510] = t[9509] ^ n[9510];
assign t[9511] = t[9510] ^ n[9511];
assign t[9512] = t[9511] ^ n[9512];
assign t[9513] = t[9512] ^ n[9513];
assign t[9514] = t[9513] ^ n[9514];
assign t[9515] = t[9514] ^ n[9515];
assign t[9516] = t[9515] ^ n[9516];
assign t[9517] = t[9516] ^ n[9517];
assign t[9518] = t[9517] ^ n[9518];
assign t[9519] = t[9518] ^ n[9519];
assign t[9520] = t[9519] ^ n[9520];
assign t[9521] = t[9520] ^ n[9521];
assign t[9522] = t[9521] ^ n[9522];
assign t[9523] = t[9522] ^ n[9523];
assign t[9524] = t[9523] ^ n[9524];
assign t[9525] = t[9524] ^ n[9525];
assign t[9526] = t[9525] ^ n[9526];
assign t[9527] = t[9526] ^ n[9527];
assign t[9528] = t[9527] ^ n[9528];
assign t[9529] = t[9528] ^ n[9529];
assign t[9530] = t[9529] ^ n[9530];
assign t[9531] = t[9530] ^ n[9531];
assign t[9532] = t[9531] ^ n[9532];
assign t[9533] = t[9532] ^ n[9533];
assign t[9534] = t[9533] ^ n[9534];
assign t[9535] = t[9534] ^ n[9535];
assign t[9536] = t[9535] ^ n[9536];
assign t[9537] = t[9536] ^ n[9537];
assign t[9538] = t[9537] ^ n[9538];
assign t[9539] = t[9538] ^ n[9539];
assign t[9540] = t[9539] ^ n[9540];
assign t[9541] = t[9540] ^ n[9541];
assign t[9542] = t[9541] ^ n[9542];
assign t[9543] = t[9542] ^ n[9543];
assign t[9544] = t[9543] ^ n[9544];
assign t[9545] = t[9544] ^ n[9545];
assign t[9546] = t[9545] ^ n[9546];
assign t[9547] = t[9546] ^ n[9547];
assign t[9548] = t[9547] ^ n[9548];
assign t[9549] = t[9548] ^ n[9549];
assign t[9550] = t[9549] ^ n[9550];
assign t[9551] = t[9550] ^ n[9551];
assign t[9552] = t[9551] ^ n[9552];
assign t[9553] = t[9552] ^ n[9553];
assign t[9554] = t[9553] ^ n[9554];
assign t[9555] = t[9554] ^ n[9555];
assign t[9556] = t[9555] ^ n[9556];
assign t[9557] = t[9556] ^ n[9557];
assign t[9558] = t[9557] ^ n[9558];
assign t[9559] = t[9558] ^ n[9559];
assign t[9560] = t[9559] ^ n[9560];
assign t[9561] = t[9560] ^ n[9561];
assign t[9562] = t[9561] ^ n[9562];
assign t[9563] = t[9562] ^ n[9563];
assign t[9564] = t[9563] ^ n[9564];
assign t[9565] = t[9564] ^ n[9565];
assign t[9566] = t[9565] ^ n[9566];
assign t[9567] = t[9566] ^ n[9567];
assign t[9568] = t[9567] ^ n[9568];
assign t[9569] = t[9568] ^ n[9569];
assign t[9570] = t[9569] ^ n[9570];
assign t[9571] = t[9570] ^ n[9571];
assign t[9572] = t[9571] ^ n[9572];
assign t[9573] = t[9572] ^ n[9573];
assign t[9574] = t[9573] ^ n[9574];
assign t[9575] = t[9574] ^ n[9575];
assign t[9576] = t[9575] ^ n[9576];
assign t[9577] = t[9576] ^ n[9577];
assign t[9578] = t[9577] ^ n[9578];
assign t[9579] = t[9578] ^ n[9579];
assign t[9580] = t[9579] ^ n[9580];
assign t[9581] = t[9580] ^ n[9581];
assign t[9582] = t[9581] ^ n[9582];
assign t[9583] = t[9582] ^ n[9583];
assign t[9584] = t[9583] ^ n[9584];
assign t[9585] = t[9584] ^ n[9585];
assign t[9586] = t[9585] ^ n[9586];
assign t[9587] = t[9586] ^ n[9587];
assign t[9588] = t[9587] ^ n[9588];
assign t[9589] = t[9588] ^ n[9589];
assign t[9590] = t[9589] ^ n[9590];
assign t[9591] = t[9590] ^ n[9591];
assign t[9592] = t[9591] ^ n[9592];
assign t[9593] = t[9592] ^ n[9593];
assign t[9594] = t[9593] ^ n[9594];
assign t[9595] = t[9594] ^ n[9595];
assign t[9596] = t[9595] ^ n[9596];
assign t[9597] = t[9596] ^ n[9597];
assign t[9598] = t[9597] ^ n[9598];
assign t[9599] = t[9598] ^ n[9599];
assign t[9600] = t[9599] ^ n[9600];
assign t[9601] = t[9600] ^ n[9601];
assign t[9602] = t[9601] ^ n[9602];
assign t[9603] = t[9602] ^ n[9603];
assign t[9604] = t[9603] ^ n[9604];
assign t[9605] = t[9604] ^ n[9605];
assign t[9606] = t[9605] ^ n[9606];
assign t[9607] = t[9606] ^ n[9607];
assign t[9608] = t[9607] ^ n[9608];
assign t[9609] = t[9608] ^ n[9609];
assign t[9610] = t[9609] ^ n[9610];
assign t[9611] = t[9610] ^ n[9611];
assign t[9612] = t[9611] ^ n[9612];
assign t[9613] = t[9612] ^ n[9613];
assign t[9614] = t[9613] ^ n[9614];
assign t[9615] = t[9614] ^ n[9615];
assign t[9616] = t[9615] ^ n[9616];
assign t[9617] = t[9616] ^ n[9617];
assign t[9618] = t[9617] ^ n[9618];
assign t[9619] = t[9618] ^ n[9619];
assign t[9620] = t[9619] ^ n[9620];
assign t[9621] = t[9620] ^ n[9621];
assign t[9622] = t[9621] ^ n[9622];
assign t[9623] = t[9622] ^ n[9623];
assign t[9624] = t[9623] ^ n[9624];
assign t[9625] = t[9624] ^ n[9625];
assign t[9626] = t[9625] ^ n[9626];
assign t[9627] = t[9626] ^ n[9627];
assign t[9628] = t[9627] ^ n[9628];
assign t[9629] = t[9628] ^ n[9629];
assign t[9630] = t[9629] ^ n[9630];
assign t[9631] = t[9630] ^ n[9631];
assign t[9632] = t[9631] ^ n[9632];
assign t[9633] = t[9632] ^ n[9633];
assign t[9634] = t[9633] ^ n[9634];
assign t[9635] = t[9634] ^ n[9635];
assign t[9636] = t[9635] ^ n[9636];
assign t[9637] = t[9636] ^ n[9637];
assign t[9638] = t[9637] ^ n[9638];
assign t[9639] = t[9638] ^ n[9639];
assign t[9640] = t[9639] ^ n[9640];
assign t[9641] = t[9640] ^ n[9641];
assign t[9642] = t[9641] ^ n[9642];
assign t[9643] = t[9642] ^ n[9643];
assign t[9644] = t[9643] ^ n[9644];
assign t[9645] = t[9644] ^ n[9645];
assign t[9646] = t[9645] ^ n[9646];
assign t[9647] = t[9646] ^ n[9647];
assign t[9648] = t[9647] ^ n[9648];
assign t[9649] = t[9648] ^ n[9649];
assign t[9650] = t[9649] ^ n[9650];
assign t[9651] = t[9650] ^ n[9651];
assign t[9652] = t[9651] ^ n[9652];
assign t[9653] = t[9652] ^ n[9653];
assign t[9654] = t[9653] ^ n[9654];
assign t[9655] = t[9654] ^ n[9655];
assign t[9656] = t[9655] ^ n[9656];
assign t[9657] = t[9656] ^ n[9657];
assign t[9658] = t[9657] ^ n[9658];
assign t[9659] = t[9658] ^ n[9659];
assign t[9660] = t[9659] ^ n[9660];
assign t[9661] = t[9660] ^ n[9661];
assign t[9662] = t[9661] ^ n[9662];
assign t[9663] = t[9662] ^ n[9663];
assign t[9664] = t[9663] ^ n[9664];
assign t[9665] = t[9664] ^ n[9665];
assign t[9666] = t[9665] ^ n[9666];
assign t[9667] = t[9666] ^ n[9667];
assign t[9668] = t[9667] ^ n[9668];
assign t[9669] = t[9668] ^ n[9669];
assign t[9670] = t[9669] ^ n[9670];
assign t[9671] = t[9670] ^ n[9671];
assign t[9672] = t[9671] ^ n[9672];
assign t[9673] = t[9672] ^ n[9673];
assign t[9674] = t[9673] ^ n[9674];
assign t[9675] = t[9674] ^ n[9675];
assign t[9676] = t[9675] ^ n[9676];
assign t[9677] = t[9676] ^ n[9677];
assign t[9678] = t[9677] ^ n[9678];
assign t[9679] = t[9678] ^ n[9679];
assign t[9680] = t[9679] ^ n[9680];
assign t[9681] = t[9680] ^ n[9681];
assign t[9682] = t[9681] ^ n[9682];
assign t[9683] = t[9682] ^ n[9683];
assign t[9684] = t[9683] ^ n[9684];
assign t[9685] = t[9684] ^ n[9685];
assign t[9686] = t[9685] ^ n[9686];
assign t[9687] = t[9686] ^ n[9687];
assign t[9688] = t[9687] ^ n[9688];
assign t[9689] = t[9688] ^ n[9689];
assign t[9690] = t[9689] ^ n[9690];
assign t[9691] = t[9690] ^ n[9691];
assign t[9692] = t[9691] ^ n[9692];
assign t[9693] = t[9692] ^ n[9693];
assign t[9694] = t[9693] ^ n[9694];
assign t[9695] = t[9694] ^ n[9695];
assign t[9696] = t[9695] ^ n[9696];
assign t[9697] = t[9696] ^ n[9697];
assign t[9698] = t[9697] ^ n[9698];
assign t[9699] = t[9698] ^ n[9699];
assign t[9700] = t[9699] ^ n[9700];
assign t[9701] = t[9700] ^ n[9701];
assign t[9702] = t[9701] ^ n[9702];
assign t[9703] = t[9702] ^ n[9703];
assign t[9704] = t[9703] ^ n[9704];
assign t[9705] = t[9704] ^ n[9705];
assign t[9706] = t[9705] ^ n[9706];
assign t[9707] = t[9706] ^ n[9707];
assign t[9708] = t[9707] ^ n[9708];
assign t[9709] = t[9708] ^ n[9709];
assign t[9710] = t[9709] ^ n[9710];
assign t[9711] = t[9710] ^ n[9711];
assign t[9712] = t[9711] ^ n[9712];
assign t[9713] = t[9712] ^ n[9713];
assign t[9714] = t[9713] ^ n[9714];
assign t[9715] = t[9714] ^ n[9715];
assign t[9716] = t[9715] ^ n[9716];
assign t[9717] = t[9716] ^ n[9717];
assign t[9718] = t[9717] ^ n[9718];
assign t[9719] = t[9718] ^ n[9719];
assign t[9720] = t[9719] ^ n[9720];
assign t[9721] = t[9720] ^ n[9721];
assign t[9722] = t[9721] ^ n[9722];
assign t[9723] = t[9722] ^ n[9723];
assign t[9724] = t[9723] ^ n[9724];
assign t[9725] = t[9724] ^ n[9725];
assign t[9726] = t[9725] ^ n[9726];
assign t[9727] = t[9726] ^ n[9727];
assign t[9728] = t[9727] ^ n[9728];
assign t[9729] = t[9728] ^ n[9729];
assign t[9730] = t[9729] ^ n[9730];
assign t[9731] = t[9730] ^ n[9731];
assign t[9732] = t[9731] ^ n[9732];
assign t[9733] = t[9732] ^ n[9733];
assign t[9734] = t[9733] ^ n[9734];
assign t[9735] = t[9734] ^ n[9735];
assign t[9736] = t[9735] ^ n[9736];
assign t[9737] = t[9736] ^ n[9737];
assign t[9738] = t[9737] ^ n[9738];
assign t[9739] = t[9738] ^ n[9739];
assign t[9740] = t[9739] ^ n[9740];
assign t[9741] = t[9740] ^ n[9741];
assign t[9742] = t[9741] ^ n[9742];
assign t[9743] = t[9742] ^ n[9743];
assign t[9744] = t[9743] ^ n[9744];
assign t[9745] = t[9744] ^ n[9745];
assign t[9746] = t[9745] ^ n[9746];
assign t[9747] = t[9746] ^ n[9747];
assign t[9748] = t[9747] ^ n[9748];
assign t[9749] = t[9748] ^ n[9749];
assign t[9750] = t[9749] ^ n[9750];
assign t[9751] = t[9750] ^ n[9751];
assign t[9752] = t[9751] ^ n[9752];
assign t[9753] = t[9752] ^ n[9753];
assign t[9754] = t[9753] ^ n[9754];
assign t[9755] = t[9754] ^ n[9755];
assign t[9756] = t[9755] ^ n[9756];
assign t[9757] = t[9756] ^ n[9757];
assign t[9758] = t[9757] ^ n[9758];
assign t[9759] = t[9758] ^ n[9759];
assign t[9760] = t[9759] ^ n[9760];
assign t[9761] = t[9760] ^ n[9761];
assign t[9762] = t[9761] ^ n[9762];
assign t[9763] = t[9762] ^ n[9763];
assign t[9764] = t[9763] ^ n[9764];
assign t[9765] = t[9764] ^ n[9765];
assign t[9766] = t[9765] ^ n[9766];
assign t[9767] = t[9766] ^ n[9767];
assign t[9768] = t[9767] ^ n[9768];
assign t[9769] = t[9768] ^ n[9769];
assign t[9770] = t[9769] ^ n[9770];
assign t[9771] = t[9770] ^ n[9771];
assign t[9772] = t[9771] ^ n[9772];
assign t[9773] = t[9772] ^ n[9773];
assign t[9774] = t[9773] ^ n[9774];
assign t[9775] = t[9774] ^ n[9775];
assign t[9776] = t[9775] ^ n[9776];
assign t[9777] = t[9776] ^ n[9777];
assign t[9778] = t[9777] ^ n[9778];
assign t[9779] = t[9778] ^ n[9779];
assign t[9780] = t[9779] ^ n[9780];
assign t[9781] = t[9780] ^ n[9781];
assign t[9782] = t[9781] ^ n[9782];
assign t[9783] = t[9782] ^ n[9783];
assign t[9784] = t[9783] ^ n[9784];
assign t[9785] = t[9784] ^ n[9785];
assign t[9786] = t[9785] ^ n[9786];
assign t[9787] = t[9786] ^ n[9787];
assign t[9788] = t[9787] ^ n[9788];
assign t[9789] = t[9788] ^ n[9789];
assign t[9790] = t[9789] ^ n[9790];
assign t[9791] = t[9790] ^ n[9791];
assign t[9792] = t[9791] ^ n[9792];
assign t[9793] = t[9792] ^ n[9793];
assign t[9794] = t[9793] ^ n[9794];
assign t[9795] = t[9794] ^ n[9795];
assign t[9796] = t[9795] ^ n[9796];
assign t[9797] = t[9796] ^ n[9797];
assign t[9798] = t[9797] ^ n[9798];
assign t[9799] = t[9798] ^ n[9799];
assign t[9800] = t[9799] ^ n[9800];
assign t[9801] = t[9800] ^ n[9801];
assign t[9802] = t[9801] ^ n[9802];
assign t[9803] = t[9802] ^ n[9803];
assign t[9804] = t[9803] ^ n[9804];
assign t[9805] = t[9804] ^ n[9805];
assign t[9806] = t[9805] ^ n[9806];
assign t[9807] = t[9806] ^ n[9807];
assign t[9808] = t[9807] ^ n[9808];
assign t[9809] = t[9808] ^ n[9809];
assign t[9810] = t[9809] ^ n[9810];
assign t[9811] = t[9810] ^ n[9811];
assign t[9812] = t[9811] ^ n[9812];
assign t[9813] = t[9812] ^ n[9813];
assign t[9814] = t[9813] ^ n[9814];
assign t[9815] = t[9814] ^ n[9815];
assign t[9816] = t[9815] ^ n[9816];
assign t[9817] = t[9816] ^ n[9817];
assign t[9818] = t[9817] ^ n[9818];
assign t[9819] = t[9818] ^ n[9819];
assign t[9820] = t[9819] ^ n[9820];
assign t[9821] = t[9820] ^ n[9821];
assign t[9822] = t[9821] ^ n[9822];
assign t[9823] = t[9822] ^ n[9823];
assign t[9824] = t[9823] ^ n[9824];
assign t[9825] = t[9824] ^ n[9825];
assign t[9826] = t[9825] ^ n[9826];
assign t[9827] = t[9826] ^ n[9827];
assign t[9828] = t[9827] ^ n[9828];
assign t[9829] = t[9828] ^ n[9829];
assign t[9830] = t[9829] ^ n[9830];
assign t[9831] = t[9830] ^ n[9831];
assign t[9832] = t[9831] ^ n[9832];
assign t[9833] = t[9832] ^ n[9833];
assign t[9834] = t[9833] ^ n[9834];
assign t[9835] = t[9834] ^ n[9835];
assign t[9836] = t[9835] ^ n[9836];
assign t[9837] = t[9836] ^ n[9837];
assign t[9838] = t[9837] ^ n[9838];
assign t[9839] = t[9838] ^ n[9839];
assign t[9840] = t[9839] ^ n[9840];
assign t[9841] = t[9840] ^ n[9841];
assign t[9842] = t[9841] ^ n[9842];
assign t[9843] = t[9842] ^ n[9843];
assign t[9844] = t[9843] ^ n[9844];
assign t[9845] = t[9844] ^ n[9845];
assign t[9846] = t[9845] ^ n[9846];
assign t[9847] = t[9846] ^ n[9847];
assign t[9848] = t[9847] ^ n[9848];
assign t[9849] = t[9848] ^ n[9849];
assign t[9850] = t[9849] ^ n[9850];
assign t[9851] = t[9850] ^ n[9851];
assign t[9852] = t[9851] ^ n[9852];
assign t[9853] = t[9852] ^ n[9853];
assign t[9854] = t[9853] ^ n[9854];
assign t[9855] = t[9854] ^ n[9855];
assign t[9856] = t[9855] ^ n[9856];
assign t[9857] = t[9856] ^ n[9857];
assign t[9858] = t[9857] ^ n[9858];
assign t[9859] = t[9858] ^ n[9859];
assign t[9860] = t[9859] ^ n[9860];
assign t[9861] = t[9860] ^ n[9861];
assign t[9862] = t[9861] ^ n[9862];
assign t[9863] = t[9862] ^ n[9863];
assign t[9864] = t[9863] ^ n[9864];
assign t[9865] = t[9864] ^ n[9865];
assign t[9866] = t[9865] ^ n[9866];
assign t[9867] = t[9866] ^ n[9867];
assign t[9868] = t[9867] ^ n[9868];
assign t[9869] = t[9868] ^ n[9869];
assign t[9870] = t[9869] ^ n[9870];
assign t[9871] = t[9870] ^ n[9871];
assign t[9872] = t[9871] ^ n[9872];
assign t[9873] = t[9872] ^ n[9873];
assign t[9874] = t[9873] ^ n[9874];
assign t[9875] = t[9874] ^ n[9875];
assign t[9876] = t[9875] ^ n[9876];
assign t[9877] = t[9876] ^ n[9877];
assign t[9878] = t[9877] ^ n[9878];
assign t[9879] = t[9878] ^ n[9879];
assign t[9880] = t[9879] ^ n[9880];
assign t[9881] = t[9880] ^ n[9881];
assign t[9882] = t[9881] ^ n[9882];
assign t[9883] = t[9882] ^ n[9883];
assign t[9884] = t[9883] ^ n[9884];
assign t[9885] = t[9884] ^ n[9885];
assign t[9886] = t[9885] ^ n[9886];
assign t[9887] = t[9886] ^ n[9887];
assign t[9888] = t[9887] ^ n[9888];
assign t[9889] = t[9888] ^ n[9889];
assign t[9890] = t[9889] ^ n[9890];
assign t[9891] = t[9890] ^ n[9891];
assign t[9892] = t[9891] ^ n[9892];
assign t[9893] = t[9892] ^ n[9893];
assign t[9894] = t[9893] ^ n[9894];
assign t[9895] = t[9894] ^ n[9895];
assign t[9896] = t[9895] ^ n[9896];
assign t[9897] = t[9896] ^ n[9897];
assign t[9898] = t[9897] ^ n[9898];
assign t[9899] = t[9898] ^ n[9899];
assign t[9900] = t[9899] ^ n[9900];
assign t[9901] = t[9900] ^ n[9901];
assign t[9902] = t[9901] ^ n[9902];
assign t[9903] = t[9902] ^ n[9903];
assign t[9904] = t[9903] ^ n[9904];
assign t[9905] = t[9904] ^ n[9905];
assign t[9906] = t[9905] ^ n[9906];
assign t[9907] = t[9906] ^ n[9907];
assign t[9908] = t[9907] ^ n[9908];
assign t[9909] = t[9908] ^ n[9909];
assign t[9910] = t[9909] ^ n[9910];
assign t[9911] = t[9910] ^ n[9911];
assign t[9912] = t[9911] ^ n[9912];
assign t[9913] = t[9912] ^ n[9913];
assign t[9914] = t[9913] ^ n[9914];
assign t[9915] = t[9914] ^ n[9915];
assign t[9916] = t[9915] ^ n[9916];
assign t[9917] = t[9916] ^ n[9917];
assign t[9918] = t[9917] ^ n[9918];
assign t[9919] = t[9918] ^ n[9919];
assign t[9920] = t[9919] ^ n[9920];
assign t[9921] = t[9920] ^ n[9921];
assign t[9922] = t[9921] ^ n[9922];
assign t[9923] = t[9922] ^ n[9923];
assign t[9924] = t[9923] ^ n[9924];
assign t[9925] = t[9924] ^ n[9925];
assign t[9926] = t[9925] ^ n[9926];
assign t[9927] = t[9926] ^ n[9927];
assign t[9928] = t[9927] ^ n[9928];
assign t[9929] = t[9928] ^ n[9929];
assign t[9930] = t[9929] ^ n[9930];
assign t[9931] = t[9930] ^ n[9931];
assign t[9932] = t[9931] ^ n[9932];
assign t[9933] = t[9932] ^ n[9933];
assign t[9934] = t[9933] ^ n[9934];
assign t[9935] = t[9934] ^ n[9935];
assign t[9936] = t[9935] ^ n[9936];
assign t[9937] = t[9936] ^ n[9937];
assign t[9938] = t[9937] ^ n[9938];
assign t[9939] = t[9938] ^ n[9939];
assign t[9940] = t[9939] ^ n[9940];
assign t[9941] = t[9940] ^ n[9941];
assign t[9942] = t[9941] ^ n[9942];
assign t[9943] = t[9942] ^ n[9943];
assign t[9944] = t[9943] ^ n[9944];
assign t[9945] = t[9944] ^ n[9945];
assign t[9946] = t[9945] ^ n[9946];
assign t[9947] = t[9946] ^ n[9947];
assign t[9948] = t[9947] ^ n[9948];
assign t[9949] = t[9948] ^ n[9949];
assign t[9950] = t[9949] ^ n[9950];
assign t[9951] = t[9950] ^ n[9951];
assign t[9952] = t[9951] ^ n[9952];
assign t[9953] = t[9952] ^ n[9953];
assign t[9954] = t[9953] ^ n[9954];
assign t[9955] = t[9954] ^ n[9955];
assign t[9956] = t[9955] ^ n[9956];
assign t[9957] = t[9956] ^ n[9957];
assign t[9958] = t[9957] ^ n[9958];
assign t[9959] = t[9958] ^ n[9959];
assign t[9960] = t[9959] ^ n[9960];
assign t[9961] = t[9960] ^ n[9961];
assign t[9962] = t[9961] ^ n[9962];
assign t[9963] = t[9962] ^ n[9963];
assign t[9964] = t[9963] ^ n[9964];
assign t[9965] = t[9964] ^ n[9965];
assign t[9966] = t[9965] ^ n[9966];
assign t[9967] = t[9966] ^ n[9967];
assign t[9968] = t[9967] ^ n[9968];
assign t[9969] = t[9968] ^ n[9969];
assign t[9970] = t[9969] ^ n[9970];
assign t[9971] = t[9970] ^ n[9971];
assign t[9972] = t[9971] ^ n[9972];
assign t[9973] = t[9972] ^ n[9973];
assign t[9974] = t[9973] ^ n[9974];
assign t[9975] = t[9974] ^ n[9975];
assign t[9976] = t[9975] ^ n[9976];
assign t[9977] = t[9976] ^ n[9977];
assign t[9978] = t[9977] ^ n[9978];
assign t[9979] = t[9978] ^ n[9979];
assign t[9980] = t[9979] ^ n[9980];
assign t[9981] = t[9980] ^ n[9981];
assign t[9982] = t[9981] ^ n[9982];
assign t[9983] = t[9982] ^ n[9983];
assign t[9984] = t[9983] ^ n[9984];
assign t[9985] = t[9984] ^ n[9985];
assign t[9986] = t[9985] ^ n[9986];
assign t[9987] = t[9986] ^ n[9987];
assign t[9988] = t[9987] ^ n[9988];
assign t[9989] = t[9988] ^ n[9989];
assign t[9990] = t[9989] ^ n[9990];
assign t[9991] = t[9990] ^ n[9991];
assign t[9992] = t[9991] ^ n[9992];
assign t[9993] = t[9992] ^ n[9993];
assign t[9994] = t[9993] ^ n[9994];
assign t[9995] = t[9994] ^ n[9995];
assign t[9996] = t[9995] ^ n[9996];
assign t[9997] = t[9996] ^ n[9997];
assign t[9998] = t[9997] ^ n[9998];
assign t[9999] = t[9998] ^ n[9999];
assign t[10000] = t[9999] ^ n[10000];
assign t[10001] = t[10000] ^ n[10001];
assign t[10002] = t[10001] ^ n[10002];
assign t[10003] = t[10002] ^ n[10003];
assign t[10004] = t[10003] ^ n[10004];
assign t[10005] = t[10004] ^ n[10005];
assign t[10006] = t[10005] ^ n[10006];
assign t[10007] = t[10006] ^ n[10007];
assign t[10008] = t[10007] ^ n[10008];
assign t[10009] = t[10008] ^ n[10009];
assign t[10010] = t[10009] ^ n[10010];
assign t[10011] = t[10010] ^ n[10011];
assign t[10012] = t[10011] ^ n[10012];
assign t[10013] = t[10012] ^ n[10013];
assign t[10014] = t[10013] ^ n[10014];
assign t[10015] = t[10014] ^ n[10015];
assign t[10016] = t[10015] ^ n[10016];
assign t[10017] = t[10016] ^ n[10017];
assign t[10018] = t[10017] ^ n[10018];
assign t[10019] = t[10018] ^ n[10019];
assign t[10020] = t[10019] ^ n[10020];
assign t[10021] = t[10020] ^ n[10021];
assign t[10022] = t[10021] ^ n[10022];
assign t[10023] = t[10022] ^ n[10023];
assign t[10024] = t[10023] ^ n[10024];
assign t[10025] = t[10024] ^ n[10025];
assign t[10026] = t[10025] ^ n[10026];
assign t[10027] = t[10026] ^ n[10027];
assign t[10028] = t[10027] ^ n[10028];
assign t[10029] = t[10028] ^ n[10029];
assign t[10030] = t[10029] ^ n[10030];
assign t[10031] = t[10030] ^ n[10031];
assign t[10032] = t[10031] ^ n[10032];
assign t[10033] = t[10032] ^ n[10033];
assign t[10034] = t[10033] ^ n[10034];
assign t[10035] = t[10034] ^ n[10035];
assign t[10036] = t[10035] ^ n[10036];
assign t[10037] = t[10036] ^ n[10037];
assign t[10038] = t[10037] ^ n[10038];
assign t[10039] = t[10038] ^ n[10039];
assign t[10040] = t[10039] ^ n[10040];
assign t[10041] = t[10040] ^ n[10041];
assign t[10042] = t[10041] ^ n[10042];
assign t[10043] = t[10042] ^ n[10043];
assign t[10044] = t[10043] ^ n[10044];
assign t[10045] = t[10044] ^ n[10045];
assign t[10046] = t[10045] ^ n[10046];
assign t[10047] = t[10046] ^ n[10047];
assign t[10048] = t[10047] ^ n[10048];
assign t[10049] = t[10048] ^ n[10049];
assign t[10050] = t[10049] ^ n[10050];
assign t[10051] = t[10050] ^ n[10051];
assign t[10052] = t[10051] ^ n[10052];
assign t[10053] = t[10052] ^ n[10053];
assign t[10054] = t[10053] ^ n[10054];
assign t[10055] = t[10054] ^ n[10055];
assign t[10056] = t[10055] ^ n[10056];
assign t[10057] = t[10056] ^ n[10057];
assign t[10058] = t[10057] ^ n[10058];
assign t[10059] = t[10058] ^ n[10059];
assign t[10060] = t[10059] ^ n[10060];
assign t[10061] = t[10060] ^ n[10061];
assign t[10062] = t[10061] ^ n[10062];
assign t[10063] = t[10062] ^ n[10063];
assign t[10064] = t[10063] ^ n[10064];
assign t[10065] = t[10064] ^ n[10065];
assign t[10066] = t[10065] ^ n[10066];
assign t[10067] = t[10066] ^ n[10067];
assign t[10068] = t[10067] ^ n[10068];
assign t[10069] = t[10068] ^ n[10069];
assign t[10070] = t[10069] ^ n[10070];
assign t[10071] = t[10070] ^ n[10071];
assign t[10072] = t[10071] ^ n[10072];
assign t[10073] = t[10072] ^ n[10073];
assign t[10074] = t[10073] ^ n[10074];
assign t[10075] = t[10074] ^ n[10075];
assign t[10076] = t[10075] ^ n[10076];
assign t[10077] = t[10076] ^ n[10077];
assign t[10078] = t[10077] ^ n[10078];
assign t[10079] = t[10078] ^ n[10079];
assign t[10080] = t[10079] ^ n[10080];
assign t[10081] = t[10080] ^ n[10081];
assign t[10082] = t[10081] ^ n[10082];
assign t[10083] = t[10082] ^ n[10083];
assign t[10084] = t[10083] ^ n[10084];
assign t[10085] = t[10084] ^ n[10085];
assign t[10086] = t[10085] ^ n[10086];
assign t[10087] = t[10086] ^ n[10087];
assign t[10088] = t[10087] ^ n[10088];
assign t[10089] = t[10088] ^ n[10089];
assign t[10090] = t[10089] ^ n[10090];
assign t[10091] = t[10090] ^ n[10091];
assign t[10092] = t[10091] ^ n[10092];
assign t[10093] = t[10092] ^ n[10093];
assign t[10094] = t[10093] ^ n[10094];
assign t[10095] = t[10094] ^ n[10095];
assign t[10096] = t[10095] ^ n[10096];
assign t[10097] = t[10096] ^ n[10097];
assign t[10098] = t[10097] ^ n[10098];
assign t[10099] = t[10098] ^ n[10099];
assign t[10100] = t[10099] ^ n[10100];
assign t[10101] = t[10100] ^ n[10101];
assign t[10102] = t[10101] ^ n[10102];
assign t[10103] = t[10102] ^ n[10103];
assign t[10104] = t[10103] ^ n[10104];
assign t[10105] = t[10104] ^ n[10105];
assign t[10106] = t[10105] ^ n[10106];
assign t[10107] = t[10106] ^ n[10107];
assign t[10108] = t[10107] ^ n[10108];
assign t[10109] = t[10108] ^ n[10109];
assign t[10110] = t[10109] ^ n[10110];
assign t[10111] = t[10110] ^ n[10111];
assign t[10112] = t[10111] ^ n[10112];
assign t[10113] = t[10112] ^ n[10113];
assign t[10114] = t[10113] ^ n[10114];
assign t[10115] = t[10114] ^ n[10115];
assign t[10116] = t[10115] ^ n[10116];
assign t[10117] = t[10116] ^ n[10117];
assign t[10118] = t[10117] ^ n[10118];
assign t[10119] = t[10118] ^ n[10119];
assign t[10120] = t[10119] ^ n[10120];
assign t[10121] = t[10120] ^ n[10121];
assign t[10122] = t[10121] ^ n[10122];
assign t[10123] = t[10122] ^ n[10123];
assign t[10124] = t[10123] ^ n[10124];
assign t[10125] = t[10124] ^ n[10125];
assign t[10126] = t[10125] ^ n[10126];
assign t[10127] = t[10126] ^ n[10127];
assign t[10128] = t[10127] ^ n[10128];
assign t[10129] = t[10128] ^ n[10129];
assign t[10130] = t[10129] ^ n[10130];
assign t[10131] = t[10130] ^ n[10131];
assign t[10132] = t[10131] ^ n[10132];
assign t[10133] = t[10132] ^ n[10133];
assign t[10134] = t[10133] ^ n[10134];
assign t[10135] = t[10134] ^ n[10135];
assign t[10136] = t[10135] ^ n[10136];
assign t[10137] = t[10136] ^ n[10137];
assign t[10138] = t[10137] ^ n[10138];
assign t[10139] = t[10138] ^ n[10139];
assign t[10140] = t[10139] ^ n[10140];
assign t[10141] = t[10140] ^ n[10141];
assign t[10142] = t[10141] ^ n[10142];
assign t[10143] = t[10142] ^ n[10143];
assign t[10144] = t[10143] ^ n[10144];
assign t[10145] = t[10144] ^ n[10145];
assign t[10146] = t[10145] ^ n[10146];
assign t[10147] = t[10146] ^ n[10147];
assign t[10148] = t[10147] ^ n[10148];
assign t[10149] = t[10148] ^ n[10149];
assign t[10150] = t[10149] ^ n[10150];
assign t[10151] = t[10150] ^ n[10151];
assign t[10152] = t[10151] ^ n[10152];
assign t[10153] = t[10152] ^ n[10153];
assign t[10154] = t[10153] ^ n[10154];
assign t[10155] = t[10154] ^ n[10155];
assign t[10156] = t[10155] ^ n[10156];
assign t[10157] = t[10156] ^ n[10157];
assign t[10158] = t[10157] ^ n[10158];
assign t[10159] = t[10158] ^ n[10159];
assign t[10160] = t[10159] ^ n[10160];
assign t[10161] = t[10160] ^ n[10161];
assign t[10162] = t[10161] ^ n[10162];
assign t[10163] = t[10162] ^ n[10163];
assign t[10164] = t[10163] ^ n[10164];
assign t[10165] = t[10164] ^ n[10165];
assign t[10166] = t[10165] ^ n[10166];
assign t[10167] = t[10166] ^ n[10167];
assign t[10168] = t[10167] ^ n[10168];
assign t[10169] = t[10168] ^ n[10169];
assign t[10170] = t[10169] ^ n[10170];
assign t[10171] = t[10170] ^ n[10171];
assign t[10172] = t[10171] ^ n[10172];
assign t[10173] = t[10172] ^ n[10173];
assign t[10174] = t[10173] ^ n[10174];
assign t[10175] = t[10174] ^ n[10175];
assign t[10176] = t[10175] ^ n[10176];
assign t[10177] = t[10176] ^ n[10177];
assign t[10178] = t[10177] ^ n[10178];
assign t[10179] = t[10178] ^ n[10179];
assign t[10180] = t[10179] ^ n[10180];
assign t[10181] = t[10180] ^ n[10181];
assign t[10182] = t[10181] ^ n[10182];
assign t[10183] = t[10182] ^ n[10183];
assign t[10184] = t[10183] ^ n[10184];
assign t[10185] = t[10184] ^ n[10185];
assign t[10186] = t[10185] ^ n[10186];
assign t[10187] = t[10186] ^ n[10187];
assign t[10188] = t[10187] ^ n[10188];
assign t[10189] = t[10188] ^ n[10189];
assign t[10190] = t[10189] ^ n[10190];
assign t[10191] = t[10190] ^ n[10191];
assign t[10192] = t[10191] ^ n[10192];
assign t[10193] = t[10192] ^ n[10193];
assign t[10194] = t[10193] ^ n[10194];
assign t[10195] = t[10194] ^ n[10195];
assign t[10196] = t[10195] ^ n[10196];
assign t[10197] = t[10196] ^ n[10197];
assign t[10198] = t[10197] ^ n[10198];
assign t[10199] = t[10198] ^ n[10199];
assign t[10200] = t[10199] ^ n[10200];
assign t[10201] = t[10200] ^ n[10201];
assign t[10202] = t[10201] ^ n[10202];
assign t[10203] = t[10202] ^ n[10203];
assign t[10204] = t[10203] ^ n[10204];
assign t[10205] = t[10204] ^ n[10205];
assign t[10206] = t[10205] ^ n[10206];
assign t[10207] = t[10206] ^ n[10207];
assign t[10208] = t[10207] ^ n[10208];
assign t[10209] = t[10208] ^ n[10209];
assign t[10210] = t[10209] ^ n[10210];
assign t[10211] = t[10210] ^ n[10211];
assign t[10212] = t[10211] ^ n[10212];
assign t[10213] = t[10212] ^ n[10213];
assign t[10214] = t[10213] ^ n[10214];
assign t[10215] = t[10214] ^ n[10215];
assign t[10216] = t[10215] ^ n[10216];
assign t[10217] = t[10216] ^ n[10217];
assign t[10218] = t[10217] ^ n[10218];
assign t[10219] = t[10218] ^ n[10219];
assign t[10220] = t[10219] ^ n[10220];
assign t[10221] = t[10220] ^ n[10221];
assign t[10222] = t[10221] ^ n[10222];
assign t[10223] = t[10222] ^ n[10223];
assign t[10224] = t[10223] ^ n[10224];
assign t[10225] = t[10224] ^ n[10225];
assign t[10226] = t[10225] ^ n[10226];
assign t[10227] = t[10226] ^ n[10227];
assign t[10228] = t[10227] ^ n[10228];
assign t[10229] = t[10228] ^ n[10229];
assign t[10230] = t[10229] ^ n[10230];
assign t[10231] = t[10230] ^ n[10231];
assign t[10232] = t[10231] ^ n[10232];
assign t[10233] = t[10232] ^ n[10233];
assign t[10234] = t[10233] ^ n[10234];
assign t[10235] = t[10234] ^ n[10235];
assign t[10236] = t[10235] ^ n[10236];
assign t[10237] = t[10236] ^ n[10237];
assign t[10238] = t[10237] ^ n[10238];
assign t[10239] = t[10238] ^ n[10239];
assign t[10240] = t[10239] ^ n[10240];
assign t[10241] = t[10240] ^ n[10241];
assign t[10242] = t[10241] ^ n[10242];
assign t[10243] = t[10242] ^ n[10243];
assign t[10244] = t[10243] ^ n[10244];
assign t[10245] = t[10244] ^ n[10245];
assign t[10246] = t[10245] ^ n[10246];
assign t[10247] = t[10246] ^ n[10247];
assign t[10248] = t[10247] ^ n[10248];
assign t[10249] = t[10248] ^ n[10249];
assign t[10250] = t[10249] ^ n[10250];
assign t[10251] = t[10250] ^ n[10251];
assign t[10252] = t[10251] ^ n[10252];
assign t[10253] = t[10252] ^ n[10253];
assign t[10254] = t[10253] ^ n[10254];
assign t[10255] = t[10254] ^ n[10255];
assign t[10256] = t[10255] ^ n[10256];
assign t[10257] = t[10256] ^ n[10257];
assign t[10258] = t[10257] ^ n[10258];
assign t[10259] = t[10258] ^ n[10259];
assign t[10260] = t[10259] ^ n[10260];
assign t[10261] = t[10260] ^ n[10261];
assign t[10262] = t[10261] ^ n[10262];
assign t[10263] = t[10262] ^ n[10263];
assign t[10264] = t[10263] ^ n[10264];
assign t[10265] = t[10264] ^ n[10265];
assign t[10266] = t[10265] ^ n[10266];
assign t[10267] = t[10266] ^ n[10267];
assign t[10268] = t[10267] ^ n[10268];
assign t[10269] = t[10268] ^ n[10269];
assign t[10270] = t[10269] ^ n[10270];
assign t[10271] = t[10270] ^ n[10271];
assign t[10272] = t[10271] ^ n[10272];
assign t[10273] = t[10272] ^ n[10273];
assign t[10274] = t[10273] ^ n[10274];
assign t[10275] = t[10274] ^ n[10275];
assign t[10276] = t[10275] ^ n[10276];
assign t[10277] = t[10276] ^ n[10277];
assign t[10278] = t[10277] ^ n[10278];
assign t[10279] = t[10278] ^ n[10279];
assign t[10280] = t[10279] ^ n[10280];
assign t[10281] = t[10280] ^ n[10281];
assign t[10282] = t[10281] ^ n[10282];
assign t[10283] = t[10282] ^ n[10283];
assign t[10284] = t[10283] ^ n[10284];
assign t[10285] = t[10284] ^ n[10285];
assign t[10286] = t[10285] ^ n[10286];
assign t[10287] = t[10286] ^ n[10287];
assign t[10288] = t[10287] ^ n[10288];
assign t[10289] = t[10288] ^ n[10289];
assign t[10290] = t[10289] ^ n[10290];
assign t[10291] = t[10290] ^ n[10291];
assign t[10292] = t[10291] ^ n[10292];
assign t[10293] = t[10292] ^ n[10293];
assign t[10294] = t[10293] ^ n[10294];
assign t[10295] = t[10294] ^ n[10295];
assign t[10296] = t[10295] ^ n[10296];
assign t[10297] = t[10296] ^ n[10297];
assign t[10298] = t[10297] ^ n[10298];
assign t[10299] = t[10298] ^ n[10299];
assign t[10300] = t[10299] ^ n[10300];
assign t[10301] = t[10300] ^ n[10301];
assign t[10302] = t[10301] ^ n[10302];
assign t[10303] = t[10302] ^ n[10303];
assign t[10304] = t[10303] ^ n[10304];
assign t[10305] = t[10304] ^ n[10305];
assign t[10306] = t[10305] ^ n[10306];
assign t[10307] = t[10306] ^ n[10307];
assign t[10308] = t[10307] ^ n[10308];
assign t[10309] = t[10308] ^ n[10309];
assign t[10310] = t[10309] ^ n[10310];
assign t[10311] = t[10310] ^ n[10311];
assign t[10312] = t[10311] ^ n[10312];
assign t[10313] = t[10312] ^ n[10313];
assign t[10314] = t[10313] ^ n[10314];
assign t[10315] = t[10314] ^ n[10315];
assign t[10316] = t[10315] ^ n[10316];
assign t[10317] = t[10316] ^ n[10317];
assign t[10318] = t[10317] ^ n[10318];
assign t[10319] = t[10318] ^ n[10319];
assign t[10320] = t[10319] ^ n[10320];
assign t[10321] = t[10320] ^ n[10321];
assign t[10322] = t[10321] ^ n[10322];
assign t[10323] = t[10322] ^ n[10323];
assign t[10324] = t[10323] ^ n[10324];
assign t[10325] = t[10324] ^ n[10325];
assign t[10326] = t[10325] ^ n[10326];
assign t[10327] = t[10326] ^ n[10327];
assign t[10328] = t[10327] ^ n[10328];
assign t[10329] = t[10328] ^ n[10329];
assign t[10330] = t[10329] ^ n[10330];
assign t[10331] = t[10330] ^ n[10331];
assign t[10332] = t[10331] ^ n[10332];
assign t[10333] = t[10332] ^ n[10333];
assign t[10334] = t[10333] ^ n[10334];
assign t[10335] = t[10334] ^ n[10335];
assign t[10336] = t[10335] ^ n[10336];
assign t[10337] = t[10336] ^ n[10337];
assign t[10338] = t[10337] ^ n[10338];
assign t[10339] = t[10338] ^ n[10339];
assign t[10340] = t[10339] ^ n[10340];
assign t[10341] = t[10340] ^ n[10341];
assign t[10342] = t[10341] ^ n[10342];
assign t[10343] = t[10342] ^ n[10343];
assign t[10344] = t[10343] ^ n[10344];
assign t[10345] = t[10344] ^ n[10345];
assign t[10346] = t[10345] ^ n[10346];
assign t[10347] = t[10346] ^ n[10347];
assign t[10348] = t[10347] ^ n[10348];
assign t[10349] = t[10348] ^ n[10349];
assign t[10350] = t[10349] ^ n[10350];
assign t[10351] = t[10350] ^ n[10351];
assign t[10352] = t[10351] ^ n[10352];
assign t[10353] = t[10352] ^ n[10353];
assign t[10354] = t[10353] ^ n[10354];
assign t[10355] = t[10354] ^ n[10355];
assign t[10356] = t[10355] ^ n[10356];
assign t[10357] = t[10356] ^ n[10357];
assign t[10358] = t[10357] ^ n[10358];
assign t[10359] = t[10358] ^ n[10359];
assign t[10360] = t[10359] ^ n[10360];
assign t[10361] = t[10360] ^ n[10361];
assign t[10362] = t[10361] ^ n[10362];
assign t[10363] = t[10362] ^ n[10363];
assign t[10364] = t[10363] ^ n[10364];
assign t[10365] = t[10364] ^ n[10365];
assign t[10366] = t[10365] ^ n[10366];
assign t[10367] = t[10366] ^ n[10367];
assign t[10368] = t[10367] ^ n[10368];
assign t[10369] = t[10368] ^ n[10369];
assign t[10370] = t[10369] ^ n[10370];
assign t[10371] = t[10370] ^ n[10371];
assign t[10372] = t[10371] ^ n[10372];
assign t[10373] = t[10372] ^ n[10373];
assign t[10374] = t[10373] ^ n[10374];
assign t[10375] = t[10374] ^ n[10375];
assign t[10376] = t[10375] ^ n[10376];
assign t[10377] = t[10376] ^ n[10377];
assign t[10378] = t[10377] ^ n[10378];
assign t[10379] = t[10378] ^ n[10379];
assign t[10380] = t[10379] ^ n[10380];
assign t[10381] = t[10380] ^ n[10381];
assign t[10382] = t[10381] ^ n[10382];
assign t[10383] = t[10382] ^ n[10383];
assign t[10384] = t[10383] ^ n[10384];
assign t[10385] = t[10384] ^ n[10385];
assign t[10386] = t[10385] ^ n[10386];
assign t[10387] = t[10386] ^ n[10387];
assign t[10388] = t[10387] ^ n[10388];
assign t[10389] = t[10388] ^ n[10389];
assign t[10390] = t[10389] ^ n[10390];
assign t[10391] = t[10390] ^ n[10391];
assign t[10392] = t[10391] ^ n[10392];
assign t[10393] = t[10392] ^ n[10393];
assign t[10394] = t[10393] ^ n[10394];
assign t[10395] = t[10394] ^ n[10395];
assign t[10396] = t[10395] ^ n[10396];
assign t[10397] = t[10396] ^ n[10397];
assign t[10398] = t[10397] ^ n[10398];
assign t[10399] = t[10398] ^ n[10399];
assign t[10400] = t[10399] ^ n[10400];
assign t[10401] = t[10400] ^ n[10401];
assign t[10402] = t[10401] ^ n[10402];
assign t[10403] = t[10402] ^ n[10403];
assign t[10404] = t[10403] ^ n[10404];
assign t[10405] = t[10404] ^ n[10405];
assign t[10406] = t[10405] ^ n[10406];
assign t[10407] = t[10406] ^ n[10407];
assign t[10408] = t[10407] ^ n[10408];
assign t[10409] = t[10408] ^ n[10409];
assign t[10410] = t[10409] ^ n[10410];
assign t[10411] = t[10410] ^ n[10411];
assign t[10412] = t[10411] ^ n[10412];
assign t[10413] = t[10412] ^ n[10413];
assign t[10414] = t[10413] ^ n[10414];
assign t[10415] = t[10414] ^ n[10415];
assign t[10416] = t[10415] ^ n[10416];
assign t[10417] = t[10416] ^ n[10417];
assign t[10418] = t[10417] ^ n[10418];
assign t[10419] = t[10418] ^ n[10419];
assign t[10420] = t[10419] ^ n[10420];
assign t[10421] = t[10420] ^ n[10421];
assign t[10422] = t[10421] ^ n[10422];
assign t[10423] = t[10422] ^ n[10423];
assign t[10424] = t[10423] ^ n[10424];
assign t[10425] = t[10424] ^ n[10425];
assign t[10426] = t[10425] ^ n[10426];
assign t[10427] = t[10426] ^ n[10427];
assign t[10428] = t[10427] ^ n[10428];
assign t[10429] = t[10428] ^ n[10429];
assign t[10430] = t[10429] ^ n[10430];
assign t[10431] = t[10430] ^ n[10431];
assign t[10432] = t[10431] ^ n[10432];
assign t[10433] = t[10432] ^ n[10433];
assign t[10434] = t[10433] ^ n[10434];
assign t[10435] = t[10434] ^ n[10435];
assign t[10436] = t[10435] ^ n[10436];
assign t[10437] = t[10436] ^ n[10437];
assign t[10438] = t[10437] ^ n[10438];
assign t[10439] = t[10438] ^ n[10439];
assign t[10440] = t[10439] ^ n[10440];
assign t[10441] = t[10440] ^ n[10441];
assign t[10442] = t[10441] ^ n[10442];
assign t[10443] = t[10442] ^ n[10443];
assign t[10444] = t[10443] ^ n[10444];
assign t[10445] = t[10444] ^ n[10445];
assign t[10446] = t[10445] ^ n[10446];
assign t[10447] = t[10446] ^ n[10447];
assign t[10448] = t[10447] ^ n[10448];
assign t[10449] = t[10448] ^ n[10449];
assign t[10450] = t[10449] ^ n[10450];
assign t[10451] = t[10450] ^ n[10451];
assign t[10452] = t[10451] ^ n[10452];
assign t[10453] = t[10452] ^ n[10453];
assign t[10454] = t[10453] ^ n[10454];
assign t[10455] = t[10454] ^ n[10455];
assign t[10456] = t[10455] ^ n[10456];
assign t[10457] = t[10456] ^ n[10457];
assign t[10458] = t[10457] ^ n[10458];
assign t[10459] = t[10458] ^ n[10459];
assign t[10460] = t[10459] ^ n[10460];
assign t[10461] = t[10460] ^ n[10461];
assign t[10462] = t[10461] ^ n[10462];
assign t[10463] = t[10462] ^ n[10463];
assign t[10464] = t[10463] ^ n[10464];
assign t[10465] = t[10464] ^ n[10465];
assign t[10466] = t[10465] ^ n[10466];
assign t[10467] = t[10466] ^ n[10467];
assign t[10468] = t[10467] ^ n[10468];
assign t[10469] = t[10468] ^ n[10469];
assign t[10470] = t[10469] ^ n[10470];
assign t[10471] = t[10470] ^ n[10471];
assign t[10472] = t[10471] ^ n[10472];
assign t[10473] = t[10472] ^ n[10473];
assign t[10474] = t[10473] ^ n[10474];
assign t[10475] = t[10474] ^ n[10475];
assign t[10476] = t[10475] ^ n[10476];
assign t[10477] = t[10476] ^ n[10477];
assign t[10478] = t[10477] ^ n[10478];
assign t[10479] = t[10478] ^ n[10479];
assign t[10480] = t[10479] ^ n[10480];
assign t[10481] = t[10480] ^ n[10481];
assign t[10482] = t[10481] ^ n[10482];
assign t[10483] = t[10482] ^ n[10483];
assign t[10484] = t[10483] ^ n[10484];
assign t[10485] = t[10484] ^ n[10485];
assign t[10486] = t[10485] ^ n[10486];
assign t[10487] = t[10486] ^ n[10487];
assign t[10488] = t[10487] ^ n[10488];
assign t[10489] = t[10488] ^ n[10489];
assign t[10490] = t[10489] ^ n[10490];
assign t[10491] = t[10490] ^ n[10491];
assign t[10492] = t[10491] ^ n[10492];
assign t[10493] = t[10492] ^ n[10493];
assign t[10494] = t[10493] ^ n[10494];
assign t[10495] = t[10494] ^ n[10495];
assign t[10496] = t[10495] ^ n[10496];
assign t[10497] = t[10496] ^ n[10497];
assign t[10498] = t[10497] ^ n[10498];
assign t[10499] = t[10498] ^ n[10499];
assign t[10500] = t[10499] ^ n[10500];
assign t[10501] = t[10500] ^ n[10501];
assign t[10502] = t[10501] ^ n[10502];
assign t[10503] = t[10502] ^ n[10503];
assign t[10504] = t[10503] ^ n[10504];
assign t[10505] = t[10504] ^ n[10505];
assign t[10506] = t[10505] ^ n[10506];
assign t[10507] = t[10506] ^ n[10507];
assign t[10508] = t[10507] ^ n[10508];
assign t[10509] = t[10508] ^ n[10509];
assign t[10510] = t[10509] ^ n[10510];
assign t[10511] = t[10510] ^ n[10511];
assign t[10512] = t[10511] ^ n[10512];
assign t[10513] = t[10512] ^ n[10513];
assign t[10514] = t[10513] ^ n[10514];
assign t[10515] = t[10514] ^ n[10515];
assign t[10516] = t[10515] ^ n[10516];
assign t[10517] = t[10516] ^ n[10517];
assign t[10518] = t[10517] ^ n[10518];
assign t[10519] = t[10518] ^ n[10519];
assign t[10520] = t[10519] ^ n[10520];
assign t[10521] = t[10520] ^ n[10521];
assign t[10522] = t[10521] ^ n[10522];
assign t[10523] = t[10522] ^ n[10523];
assign t[10524] = t[10523] ^ n[10524];
assign t[10525] = t[10524] ^ n[10525];
assign t[10526] = t[10525] ^ n[10526];
assign t[10527] = t[10526] ^ n[10527];
assign t[10528] = t[10527] ^ n[10528];
assign t[10529] = t[10528] ^ n[10529];
assign t[10530] = t[10529] ^ n[10530];
assign t[10531] = t[10530] ^ n[10531];
assign t[10532] = t[10531] ^ n[10532];
assign t[10533] = t[10532] ^ n[10533];
assign t[10534] = t[10533] ^ n[10534];
assign t[10535] = t[10534] ^ n[10535];
assign t[10536] = t[10535] ^ n[10536];
assign t[10537] = t[10536] ^ n[10537];
assign t[10538] = t[10537] ^ n[10538];
assign t[10539] = t[10538] ^ n[10539];
assign t[10540] = t[10539] ^ n[10540];
assign t[10541] = t[10540] ^ n[10541];
assign t[10542] = t[10541] ^ n[10542];
assign t[10543] = t[10542] ^ n[10543];
assign t[10544] = t[10543] ^ n[10544];
assign t[10545] = t[10544] ^ n[10545];
assign t[10546] = t[10545] ^ n[10546];
assign t[10547] = t[10546] ^ n[10547];
assign t[10548] = t[10547] ^ n[10548];
assign t[10549] = t[10548] ^ n[10549];
assign t[10550] = t[10549] ^ n[10550];
assign t[10551] = t[10550] ^ n[10551];
assign t[10552] = t[10551] ^ n[10552];
assign t[10553] = t[10552] ^ n[10553];
assign t[10554] = t[10553] ^ n[10554];
assign t[10555] = t[10554] ^ n[10555];
assign t[10556] = t[10555] ^ n[10556];
assign t[10557] = t[10556] ^ n[10557];
assign t[10558] = t[10557] ^ n[10558];
assign t[10559] = t[10558] ^ n[10559];
assign t[10560] = t[10559] ^ n[10560];
assign t[10561] = t[10560] ^ n[10561];
assign t[10562] = t[10561] ^ n[10562];
assign t[10563] = t[10562] ^ n[10563];
assign t[10564] = t[10563] ^ n[10564];
assign t[10565] = t[10564] ^ n[10565];
assign t[10566] = t[10565] ^ n[10566];
assign t[10567] = t[10566] ^ n[10567];
assign t[10568] = t[10567] ^ n[10568];
assign t[10569] = t[10568] ^ n[10569];
assign t[10570] = t[10569] ^ n[10570];
assign t[10571] = t[10570] ^ n[10571];
assign t[10572] = t[10571] ^ n[10572];
assign t[10573] = t[10572] ^ n[10573];
assign t[10574] = t[10573] ^ n[10574];
assign t[10575] = t[10574] ^ n[10575];
assign t[10576] = t[10575] ^ n[10576];
assign t[10577] = t[10576] ^ n[10577];
assign t[10578] = t[10577] ^ n[10578];
assign t[10579] = t[10578] ^ n[10579];
assign t[10580] = t[10579] ^ n[10580];
assign t[10581] = t[10580] ^ n[10581];
assign t[10582] = t[10581] ^ n[10582];
assign t[10583] = t[10582] ^ n[10583];
assign t[10584] = t[10583] ^ n[10584];
assign t[10585] = t[10584] ^ n[10585];
assign t[10586] = t[10585] ^ n[10586];
assign t[10587] = t[10586] ^ n[10587];
assign t[10588] = t[10587] ^ n[10588];
assign t[10589] = t[10588] ^ n[10589];
assign t[10590] = t[10589] ^ n[10590];
assign t[10591] = t[10590] ^ n[10591];
assign t[10592] = t[10591] ^ n[10592];
assign t[10593] = t[10592] ^ n[10593];
assign t[10594] = t[10593] ^ n[10594];
assign t[10595] = t[10594] ^ n[10595];
assign t[10596] = t[10595] ^ n[10596];
assign t[10597] = t[10596] ^ n[10597];
assign t[10598] = t[10597] ^ n[10598];
assign t[10599] = t[10598] ^ n[10599];
assign t[10600] = t[10599] ^ n[10600];
assign t[10601] = t[10600] ^ n[10601];
assign t[10602] = t[10601] ^ n[10602];
assign t[10603] = t[10602] ^ n[10603];
assign t[10604] = t[10603] ^ n[10604];
assign t[10605] = t[10604] ^ n[10605];
assign t[10606] = t[10605] ^ n[10606];
assign t[10607] = t[10606] ^ n[10607];
assign t[10608] = t[10607] ^ n[10608];
assign t[10609] = t[10608] ^ n[10609];
assign t[10610] = t[10609] ^ n[10610];
assign t[10611] = t[10610] ^ n[10611];
assign t[10612] = t[10611] ^ n[10612];
assign t[10613] = t[10612] ^ n[10613];
assign t[10614] = t[10613] ^ n[10614];
assign t[10615] = t[10614] ^ n[10615];
assign t[10616] = t[10615] ^ n[10616];
assign t[10617] = t[10616] ^ n[10617];
assign t[10618] = t[10617] ^ n[10618];
assign t[10619] = t[10618] ^ n[10619];
assign t[10620] = t[10619] ^ n[10620];
assign t[10621] = t[10620] ^ n[10621];
assign t[10622] = t[10621] ^ n[10622];
assign t[10623] = t[10622] ^ n[10623];
assign t[10624] = t[10623] ^ n[10624];
assign t[10625] = t[10624] ^ n[10625];
assign t[10626] = t[10625] ^ n[10626];
assign t[10627] = t[10626] ^ n[10627];
assign t[10628] = t[10627] ^ n[10628];
assign t[10629] = t[10628] ^ n[10629];
assign t[10630] = t[10629] ^ n[10630];
assign t[10631] = t[10630] ^ n[10631];
assign t[10632] = t[10631] ^ n[10632];
assign t[10633] = t[10632] ^ n[10633];
assign t[10634] = t[10633] ^ n[10634];
assign t[10635] = t[10634] ^ n[10635];
assign t[10636] = t[10635] ^ n[10636];
assign t[10637] = t[10636] ^ n[10637];
assign t[10638] = t[10637] ^ n[10638];
assign t[10639] = t[10638] ^ n[10639];
assign t[10640] = t[10639] ^ n[10640];
assign t[10641] = t[10640] ^ n[10641];
assign t[10642] = t[10641] ^ n[10642];
assign t[10643] = t[10642] ^ n[10643];
assign t[10644] = t[10643] ^ n[10644];
assign t[10645] = t[10644] ^ n[10645];
assign t[10646] = t[10645] ^ n[10646];
assign t[10647] = t[10646] ^ n[10647];
assign t[10648] = t[10647] ^ n[10648];
assign t[10649] = t[10648] ^ n[10649];
assign t[10650] = t[10649] ^ n[10650];
assign t[10651] = t[10650] ^ n[10651];
assign t[10652] = t[10651] ^ n[10652];
assign t[10653] = t[10652] ^ n[10653];
assign t[10654] = t[10653] ^ n[10654];
assign t[10655] = t[10654] ^ n[10655];
assign t[10656] = t[10655] ^ n[10656];
assign t[10657] = t[10656] ^ n[10657];
assign t[10658] = t[10657] ^ n[10658];
assign t[10659] = t[10658] ^ n[10659];
assign t[10660] = t[10659] ^ n[10660];
assign t[10661] = t[10660] ^ n[10661];
assign t[10662] = t[10661] ^ n[10662];
assign t[10663] = t[10662] ^ n[10663];
assign t[10664] = t[10663] ^ n[10664];
assign t[10665] = t[10664] ^ n[10665];
assign t[10666] = t[10665] ^ n[10666];
assign t[10667] = t[10666] ^ n[10667];
assign t[10668] = t[10667] ^ n[10668];
assign t[10669] = t[10668] ^ n[10669];
assign t[10670] = t[10669] ^ n[10670];
assign t[10671] = t[10670] ^ n[10671];
assign t[10672] = t[10671] ^ n[10672];
assign t[10673] = t[10672] ^ n[10673];
assign t[10674] = t[10673] ^ n[10674];
assign t[10675] = t[10674] ^ n[10675];
assign t[10676] = t[10675] ^ n[10676];
assign t[10677] = t[10676] ^ n[10677];
assign t[10678] = t[10677] ^ n[10678];
assign t[10679] = t[10678] ^ n[10679];
assign t[10680] = t[10679] ^ n[10680];
assign t[10681] = t[10680] ^ n[10681];
assign t[10682] = t[10681] ^ n[10682];
assign t[10683] = t[10682] ^ n[10683];
assign t[10684] = t[10683] ^ n[10684];
assign t[10685] = t[10684] ^ n[10685];
assign t[10686] = t[10685] ^ n[10686];
assign t[10687] = t[10686] ^ n[10687];
assign t[10688] = t[10687] ^ n[10688];
assign t[10689] = t[10688] ^ n[10689];
assign t[10690] = t[10689] ^ n[10690];
assign t[10691] = t[10690] ^ n[10691];
assign t[10692] = t[10691] ^ n[10692];
assign t[10693] = t[10692] ^ n[10693];
assign t[10694] = t[10693] ^ n[10694];
assign t[10695] = t[10694] ^ n[10695];
assign t[10696] = t[10695] ^ n[10696];
assign t[10697] = t[10696] ^ n[10697];
assign t[10698] = t[10697] ^ n[10698];
assign t[10699] = t[10698] ^ n[10699];
assign t[10700] = t[10699] ^ n[10700];
assign t[10701] = t[10700] ^ n[10701];
assign t[10702] = t[10701] ^ n[10702];
assign t[10703] = t[10702] ^ n[10703];
assign t[10704] = t[10703] ^ n[10704];
assign t[10705] = t[10704] ^ n[10705];
assign t[10706] = t[10705] ^ n[10706];
assign t[10707] = t[10706] ^ n[10707];
assign t[10708] = t[10707] ^ n[10708];
assign t[10709] = t[10708] ^ n[10709];
assign t[10710] = t[10709] ^ n[10710];
assign t[10711] = t[10710] ^ n[10711];
assign t[10712] = t[10711] ^ n[10712];
assign t[10713] = t[10712] ^ n[10713];
assign t[10714] = t[10713] ^ n[10714];
assign t[10715] = t[10714] ^ n[10715];
assign t[10716] = t[10715] ^ n[10716];
assign t[10717] = t[10716] ^ n[10717];
assign t[10718] = t[10717] ^ n[10718];
assign t[10719] = t[10718] ^ n[10719];
assign t[10720] = t[10719] ^ n[10720];
assign t[10721] = t[10720] ^ n[10721];
assign t[10722] = t[10721] ^ n[10722];
assign t[10723] = t[10722] ^ n[10723];
assign t[10724] = t[10723] ^ n[10724];
assign t[10725] = t[10724] ^ n[10725];
assign t[10726] = t[10725] ^ n[10726];
assign t[10727] = t[10726] ^ n[10727];
assign t[10728] = t[10727] ^ n[10728];
assign t[10729] = t[10728] ^ n[10729];
assign t[10730] = t[10729] ^ n[10730];
assign t[10731] = t[10730] ^ n[10731];
assign t[10732] = t[10731] ^ n[10732];
assign t[10733] = t[10732] ^ n[10733];
assign t[10734] = t[10733] ^ n[10734];
assign t[10735] = t[10734] ^ n[10735];
assign t[10736] = t[10735] ^ n[10736];
assign t[10737] = t[10736] ^ n[10737];
assign t[10738] = t[10737] ^ n[10738];
assign t[10739] = t[10738] ^ n[10739];
assign t[10740] = t[10739] ^ n[10740];
assign t[10741] = t[10740] ^ n[10741];
assign t[10742] = t[10741] ^ n[10742];
assign t[10743] = t[10742] ^ n[10743];
assign t[10744] = t[10743] ^ n[10744];
assign t[10745] = t[10744] ^ n[10745];
assign t[10746] = t[10745] ^ n[10746];
assign t[10747] = t[10746] ^ n[10747];
assign t[10748] = t[10747] ^ n[10748];
assign t[10749] = t[10748] ^ n[10749];
assign t[10750] = t[10749] ^ n[10750];
assign t[10751] = t[10750] ^ n[10751];
assign t[10752] = t[10751] ^ n[10752];
assign t[10753] = t[10752] ^ n[10753];
assign t[10754] = t[10753] ^ n[10754];
assign t[10755] = t[10754] ^ n[10755];
assign t[10756] = t[10755] ^ n[10756];
assign t[10757] = t[10756] ^ n[10757];
assign t[10758] = t[10757] ^ n[10758];
assign t[10759] = t[10758] ^ n[10759];
assign t[10760] = t[10759] ^ n[10760];
assign t[10761] = t[10760] ^ n[10761];
assign t[10762] = t[10761] ^ n[10762];
assign t[10763] = t[10762] ^ n[10763];
assign t[10764] = t[10763] ^ n[10764];
assign t[10765] = t[10764] ^ n[10765];
assign t[10766] = t[10765] ^ n[10766];
assign t[10767] = t[10766] ^ n[10767];
assign t[10768] = t[10767] ^ n[10768];
assign t[10769] = t[10768] ^ n[10769];
assign t[10770] = t[10769] ^ n[10770];
assign t[10771] = t[10770] ^ n[10771];
assign t[10772] = t[10771] ^ n[10772];
assign t[10773] = t[10772] ^ n[10773];
assign t[10774] = t[10773] ^ n[10774];
assign t[10775] = t[10774] ^ n[10775];
assign t[10776] = t[10775] ^ n[10776];
assign t[10777] = t[10776] ^ n[10777];
assign t[10778] = t[10777] ^ n[10778];
assign t[10779] = t[10778] ^ n[10779];
assign t[10780] = t[10779] ^ n[10780];
assign t[10781] = t[10780] ^ n[10781];
assign t[10782] = t[10781] ^ n[10782];
assign t[10783] = t[10782] ^ n[10783];
assign t[10784] = t[10783] ^ n[10784];
assign t[10785] = t[10784] ^ n[10785];
assign t[10786] = t[10785] ^ n[10786];
assign t[10787] = t[10786] ^ n[10787];
assign t[10788] = t[10787] ^ n[10788];
assign t[10789] = t[10788] ^ n[10789];
assign t[10790] = t[10789] ^ n[10790];
assign t[10791] = t[10790] ^ n[10791];
assign t[10792] = t[10791] ^ n[10792];
assign t[10793] = t[10792] ^ n[10793];
assign t[10794] = t[10793] ^ n[10794];
assign t[10795] = t[10794] ^ n[10795];
assign t[10796] = t[10795] ^ n[10796];
assign t[10797] = t[10796] ^ n[10797];
assign t[10798] = t[10797] ^ n[10798];
assign t[10799] = t[10798] ^ n[10799];
assign t[10800] = t[10799] ^ n[10800];
assign t[10801] = t[10800] ^ n[10801];
assign t[10802] = t[10801] ^ n[10802];
assign t[10803] = t[10802] ^ n[10803];
assign t[10804] = t[10803] ^ n[10804];
assign t[10805] = t[10804] ^ n[10805];
assign t[10806] = t[10805] ^ n[10806];
assign t[10807] = t[10806] ^ n[10807];
assign t[10808] = t[10807] ^ n[10808];
assign t[10809] = t[10808] ^ n[10809];
assign t[10810] = t[10809] ^ n[10810];
assign t[10811] = t[10810] ^ n[10811];
assign t[10812] = t[10811] ^ n[10812];
assign t[10813] = t[10812] ^ n[10813];
assign t[10814] = t[10813] ^ n[10814];
assign t[10815] = t[10814] ^ n[10815];
assign t[10816] = t[10815] ^ n[10816];
assign t[10817] = t[10816] ^ n[10817];
assign t[10818] = t[10817] ^ n[10818];
assign t[10819] = t[10818] ^ n[10819];
assign t[10820] = t[10819] ^ n[10820];
assign t[10821] = t[10820] ^ n[10821];
assign t[10822] = t[10821] ^ n[10822];
assign t[10823] = t[10822] ^ n[10823];
assign t[10824] = t[10823] ^ n[10824];
assign t[10825] = t[10824] ^ n[10825];
assign t[10826] = t[10825] ^ n[10826];
assign t[10827] = t[10826] ^ n[10827];
assign t[10828] = t[10827] ^ n[10828];
assign t[10829] = t[10828] ^ n[10829];
assign t[10830] = t[10829] ^ n[10830];
assign t[10831] = t[10830] ^ n[10831];
assign t[10832] = t[10831] ^ n[10832];
assign t[10833] = t[10832] ^ n[10833];
assign t[10834] = t[10833] ^ n[10834];
assign t[10835] = t[10834] ^ n[10835];
assign t[10836] = t[10835] ^ n[10836];
assign t[10837] = t[10836] ^ n[10837];
assign t[10838] = t[10837] ^ n[10838];
assign t[10839] = t[10838] ^ n[10839];
assign t[10840] = t[10839] ^ n[10840];
assign t[10841] = t[10840] ^ n[10841];
assign t[10842] = t[10841] ^ n[10842];
assign t[10843] = t[10842] ^ n[10843];
assign t[10844] = t[10843] ^ n[10844];
assign t[10845] = t[10844] ^ n[10845];
assign t[10846] = t[10845] ^ n[10846];
assign t[10847] = t[10846] ^ n[10847];
assign t[10848] = t[10847] ^ n[10848];
assign t[10849] = t[10848] ^ n[10849];
assign t[10850] = t[10849] ^ n[10850];
assign t[10851] = t[10850] ^ n[10851];
assign t[10852] = t[10851] ^ n[10852];
assign t[10853] = t[10852] ^ n[10853];
assign t[10854] = t[10853] ^ n[10854];
assign t[10855] = t[10854] ^ n[10855];
assign t[10856] = t[10855] ^ n[10856];
assign t[10857] = t[10856] ^ n[10857];
assign t[10858] = t[10857] ^ n[10858];
assign t[10859] = t[10858] ^ n[10859];
assign t[10860] = t[10859] ^ n[10860];
assign t[10861] = t[10860] ^ n[10861];
assign t[10862] = t[10861] ^ n[10862];
assign t[10863] = t[10862] ^ n[10863];
assign t[10864] = t[10863] ^ n[10864];
assign t[10865] = t[10864] ^ n[10865];
assign t[10866] = t[10865] ^ n[10866];
assign t[10867] = t[10866] ^ n[10867];
assign t[10868] = t[10867] ^ n[10868];
assign t[10869] = t[10868] ^ n[10869];
assign t[10870] = t[10869] ^ n[10870];
assign t[10871] = t[10870] ^ n[10871];
assign t[10872] = t[10871] ^ n[10872];
assign t[10873] = t[10872] ^ n[10873];
assign t[10874] = t[10873] ^ n[10874];
assign t[10875] = t[10874] ^ n[10875];
assign t[10876] = t[10875] ^ n[10876];
assign t[10877] = t[10876] ^ n[10877];
assign t[10878] = t[10877] ^ n[10878];
assign t[10879] = t[10878] ^ n[10879];
assign t[10880] = t[10879] ^ n[10880];
assign t[10881] = t[10880] ^ n[10881];
assign t[10882] = t[10881] ^ n[10882];
assign t[10883] = t[10882] ^ n[10883];
assign t[10884] = t[10883] ^ n[10884];
assign t[10885] = t[10884] ^ n[10885];
assign t[10886] = t[10885] ^ n[10886];
assign t[10887] = t[10886] ^ n[10887];
assign t[10888] = t[10887] ^ n[10888];
assign t[10889] = t[10888] ^ n[10889];
assign t[10890] = t[10889] ^ n[10890];
assign t[10891] = t[10890] ^ n[10891];
assign t[10892] = t[10891] ^ n[10892];
assign t[10893] = t[10892] ^ n[10893];
assign t[10894] = t[10893] ^ n[10894];
assign t[10895] = t[10894] ^ n[10895];
assign t[10896] = t[10895] ^ n[10896];
assign t[10897] = t[10896] ^ n[10897];
assign t[10898] = t[10897] ^ n[10898];
assign t[10899] = t[10898] ^ n[10899];
assign t[10900] = t[10899] ^ n[10900];
assign t[10901] = t[10900] ^ n[10901];
assign t[10902] = t[10901] ^ n[10902];
assign t[10903] = t[10902] ^ n[10903];
assign t[10904] = t[10903] ^ n[10904];
assign t[10905] = t[10904] ^ n[10905];
assign t[10906] = t[10905] ^ n[10906];
assign t[10907] = t[10906] ^ n[10907];
assign t[10908] = t[10907] ^ n[10908];
assign t[10909] = t[10908] ^ n[10909];
assign t[10910] = t[10909] ^ n[10910];
assign t[10911] = t[10910] ^ n[10911];
assign t[10912] = t[10911] ^ n[10912];
assign t[10913] = t[10912] ^ n[10913];
assign t[10914] = t[10913] ^ n[10914];
assign t[10915] = t[10914] ^ n[10915];
assign t[10916] = t[10915] ^ n[10916];
assign t[10917] = t[10916] ^ n[10917];
assign t[10918] = t[10917] ^ n[10918];
assign t[10919] = t[10918] ^ n[10919];
assign t[10920] = t[10919] ^ n[10920];
assign t[10921] = t[10920] ^ n[10921];
assign t[10922] = t[10921] ^ n[10922];
assign t[10923] = t[10922] ^ n[10923];
assign t[10924] = t[10923] ^ n[10924];
assign t[10925] = t[10924] ^ n[10925];
assign t[10926] = t[10925] ^ n[10926];
assign t[10927] = t[10926] ^ n[10927];
assign t[10928] = t[10927] ^ n[10928];
assign t[10929] = t[10928] ^ n[10929];
assign t[10930] = t[10929] ^ n[10930];
assign t[10931] = t[10930] ^ n[10931];
assign t[10932] = t[10931] ^ n[10932];
assign t[10933] = t[10932] ^ n[10933];
assign t[10934] = t[10933] ^ n[10934];
assign t[10935] = t[10934] ^ n[10935];
assign t[10936] = t[10935] ^ n[10936];
assign t[10937] = t[10936] ^ n[10937];
assign t[10938] = t[10937] ^ n[10938];
assign t[10939] = t[10938] ^ n[10939];
assign t[10940] = t[10939] ^ n[10940];
assign t[10941] = t[10940] ^ n[10941];
assign t[10942] = t[10941] ^ n[10942];
assign t[10943] = t[10942] ^ n[10943];
assign t[10944] = t[10943] ^ n[10944];
assign t[10945] = t[10944] ^ n[10945];
assign t[10946] = t[10945] ^ n[10946];
assign t[10947] = t[10946] ^ n[10947];
assign t[10948] = t[10947] ^ n[10948];
assign t[10949] = t[10948] ^ n[10949];
assign t[10950] = t[10949] ^ n[10950];
assign t[10951] = t[10950] ^ n[10951];
assign t[10952] = t[10951] ^ n[10952];
assign t[10953] = t[10952] ^ n[10953];
assign t[10954] = t[10953] ^ n[10954];
assign t[10955] = t[10954] ^ n[10955];
assign t[10956] = t[10955] ^ n[10956];
assign t[10957] = t[10956] ^ n[10957];
assign t[10958] = t[10957] ^ n[10958];
assign t[10959] = t[10958] ^ n[10959];
assign t[10960] = t[10959] ^ n[10960];
assign t[10961] = t[10960] ^ n[10961];
assign t[10962] = t[10961] ^ n[10962];
assign t[10963] = t[10962] ^ n[10963];
assign t[10964] = t[10963] ^ n[10964];
assign t[10965] = t[10964] ^ n[10965];
assign t[10966] = t[10965] ^ n[10966];
assign t[10967] = t[10966] ^ n[10967];
assign t[10968] = t[10967] ^ n[10968];
assign t[10969] = t[10968] ^ n[10969];
assign t[10970] = t[10969] ^ n[10970];
assign t[10971] = t[10970] ^ n[10971];
assign t[10972] = t[10971] ^ n[10972];
assign t[10973] = t[10972] ^ n[10973];
assign t[10974] = t[10973] ^ n[10974];
assign t[10975] = t[10974] ^ n[10975];
assign t[10976] = t[10975] ^ n[10976];
assign t[10977] = t[10976] ^ n[10977];
assign t[10978] = t[10977] ^ n[10978];
assign t[10979] = t[10978] ^ n[10979];
assign t[10980] = t[10979] ^ n[10980];
assign t[10981] = t[10980] ^ n[10981];
assign t[10982] = t[10981] ^ n[10982];
assign t[10983] = t[10982] ^ n[10983];
assign t[10984] = t[10983] ^ n[10984];
assign t[10985] = t[10984] ^ n[10985];
assign t[10986] = t[10985] ^ n[10986];
assign t[10987] = t[10986] ^ n[10987];
assign t[10988] = t[10987] ^ n[10988];
assign t[10989] = t[10988] ^ n[10989];
assign t[10990] = t[10989] ^ n[10990];
assign t[10991] = t[10990] ^ n[10991];
assign t[10992] = t[10991] ^ n[10992];
assign t[10993] = t[10992] ^ n[10993];
assign t[10994] = t[10993] ^ n[10994];
assign t[10995] = t[10994] ^ n[10995];
assign t[10996] = t[10995] ^ n[10996];
assign t[10997] = t[10996] ^ n[10997];
assign t[10998] = t[10997] ^ n[10998];
assign t[10999] = t[10998] ^ n[10999];
assign t[11000] = t[10999] ^ n[11000];
assign t[11001] = t[11000] ^ n[11001];
assign t[11002] = t[11001] ^ n[11002];
assign t[11003] = t[11002] ^ n[11003];
assign t[11004] = t[11003] ^ n[11004];
assign t[11005] = t[11004] ^ n[11005];
assign t[11006] = t[11005] ^ n[11006];
assign t[11007] = t[11006] ^ n[11007];
assign t[11008] = t[11007] ^ n[11008];
assign t[11009] = t[11008] ^ n[11009];
assign t[11010] = t[11009] ^ n[11010];
assign t[11011] = t[11010] ^ n[11011];
assign t[11012] = t[11011] ^ n[11012];
assign t[11013] = t[11012] ^ n[11013];
assign t[11014] = t[11013] ^ n[11014];
assign t[11015] = t[11014] ^ n[11015];
assign t[11016] = t[11015] ^ n[11016];
assign t[11017] = t[11016] ^ n[11017];
assign t[11018] = t[11017] ^ n[11018];
assign t[11019] = t[11018] ^ n[11019];
assign t[11020] = t[11019] ^ n[11020];
assign t[11021] = t[11020] ^ n[11021];
assign t[11022] = t[11021] ^ n[11022];
assign t[11023] = t[11022] ^ n[11023];
assign t[11024] = t[11023] ^ n[11024];
assign t[11025] = t[11024] ^ n[11025];
assign t[11026] = t[11025] ^ n[11026];
assign t[11027] = t[11026] ^ n[11027];
assign t[11028] = t[11027] ^ n[11028];
assign t[11029] = t[11028] ^ n[11029];
assign t[11030] = t[11029] ^ n[11030];
assign t[11031] = t[11030] ^ n[11031];
assign t[11032] = t[11031] ^ n[11032];
assign t[11033] = t[11032] ^ n[11033];
assign t[11034] = t[11033] ^ n[11034];
assign t[11035] = t[11034] ^ n[11035];
assign t[11036] = t[11035] ^ n[11036];
assign t[11037] = t[11036] ^ n[11037];
assign t[11038] = t[11037] ^ n[11038];
assign t[11039] = t[11038] ^ n[11039];
assign t[11040] = t[11039] ^ n[11040];
assign t[11041] = t[11040] ^ n[11041];
assign t[11042] = t[11041] ^ n[11042];
assign t[11043] = t[11042] ^ n[11043];
assign t[11044] = t[11043] ^ n[11044];
assign t[11045] = t[11044] ^ n[11045];
assign t[11046] = t[11045] ^ n[11046];
assign t[11047] = t[11046] ^ n[11047];
assign t[11048] = t[11047] ^ n[11048];
assign t[11049] = t[11048] ^ n[11049];
assign t[11050] = t[11049] ^ n[11050];
assign t[11051] = t[11050] ^ n[11051];
assign t[11052] = t[11051] ^ n[11052];
assign t[11053] = t[11052] ^ n[11053];
assign t[11054] = t[11053] ^ n[11054];
assign t[11055] = t[11054] ^ n[11055];
assign t[11056] = t[11055] ^ n[11056];
assign t[11057] = t[11056] ^ n[11057];
assign t[11058] = t[11057] ^ n[11058];
assign t[11059] = t[11058] ^ n[11059];
assign t[11060] = t[11059] ^ n[11060];
assign t[11061] = t[11060] ^ n[11061];
assign t[11062] = t[11061] ^ n[11062];
assign t[11063] = t[11062] ^ n[11063];
assign t[11064] = t[11063] ^ n[11064];
assign t[11065] = t[11064] ^ n[11065];
assign t[11066] = t[11065] ^ n[11066];
assign t[11067] = t[11066] ^ n[11067];
assign t[11068] = t[11067] ^ n[11068];
assign t[11069] = t[11068] ^ n[11069];
assign t[11070] = t[11069] ^ n[11070];
assign t[11071] = t[11070] ^ n[11071];
assign t[11072] = t[11071] ^ n[11072];
assign t[11073] = t[11072] ^ n[11073];
assign t[11074] = t[11073] ^ n[11074];
assign t[11075] = t[11074] ^ n[11075];
assign t[11076] = t[11075] ^ n[11076];
assign t[11077] = t[11076] ^ n[11077];
assign t[11078] = t[11077] ^ n[11078];
assign t[11079] = t[11078] ^ n[11079];
assign t[11080] = t[11079] ^ n[11080];
assign t[11081] = t[11080] ^ n[11081];
assign t[11082] = t[11081] ^ n[11082];
assign t[11083] = t[11082] ^ n[11083];
assign t[11084] = t[11083] ^ n[11084];
assign t[11085] = t[11084] ^ n[11085];
assign t[11086] = t[11085] ^ n[11086];
assign t[11087] = t[11086] ^ n[11087];
assign t[11088] = t[11087] ^ n[11088];
assign t[11089] = t[11088] ^ n[11089];
assign t[11090] = t[11089] ^ n[11090];
assign t[11091] = t[11090] ^ n[11091];
assign t[11092] = t[11091] ^ n[11092];
assign t[11093] = t[11092] ^ n[11093];
assign t[11094] = t[11093] ^ n[11094];
assign t[11095] = t[11094] ^ n[11095];
assign t[11096] = t[11095] ^ n[11096];
assign t[11097] = t[11096] ^ n[11097];
assign t[11098] = t[11097] ^ n[11098];
assign t[11099] = t[11098] ^ n[11099];
assign t[11100] = t[11099] ^ n[11100];
assign t[11101] = t[11100] ^ n[11101];
assign t[11102] = t[11101] ^ n[11102];
assign t[11103] = t[11102] ^ n[11103];
assign t[11104] = t[11103] ^ n[11104];
assign t[11105] = t[11104] ^ n[11105];
assign t[11106] = t[11105] ^ n[11106];
assign t[11107] = t[11106] ^ n[11107];
assign t[11108] = t[11107] ^ n[11108];
assign t[11109] = t[11108] ^ n[11109];
assign t[11110] = t[11109] ^ n[11110];
assign t[11111] = t[11110] ^ n[11111];
assign t[11112] = t[11111] ^ n[11112];
assign t[11113] = t[11112] ^ n[11113];
assign t[11114] = t[11113] ^ n[11114];
assign t[11115] = t[11114] ^ n[11115];
assign t[11116] = t[11115] ^ n[11116];
assign t[11117] = t[11116] ^ n[11117];
assign t[11118] = t[11117] ^ n[11118];
assign t[11119] = t[11118] ^ n[11119];
assign t[11120] = t[11119] ^ n[11120];
assign t[11121] = t[11120] ^ n[11121];
assign t[11122] = t[11121] ^ n[11122];
assign t[11123] = t[11122] ^ n[11123];
assign t[11124] = t[11123] ^ n[11124];
assign t[11125] = t[11124] ^ n[11125];
assign t[11126] = t[11125] ^ n[11126];
assign t[11127] = t[11126] ^ n[11127];
assign t[11128] = t[11127] ^ n[11128];
assign t[11129] = t[11128] ^ n[11129];
assign t[11130] = t[11129] ^ n[11130];
assign t[11131] = t[11130] ^ n[11131];
assign t[11132] = t[11131] ^ n[11132];
assign t[11133] = t[11132] ^ n[11133];
assign t[11134] = t[11133] ^ n[11134];
assign t[11135] = t[11134] ^ n[11135];
assign t[11136] = t[11135] ^ n[11136];
assign t[11137] = t[11136] ^ n[11137];
assign t[11138] = t[11137] ^ n[11138];
assign t[11139] = t[11138] ^ n[11139];
assign t[11140] = t[11139] ^ n[11140];
assign t[11141] = t[11140] ^ n[11141];
assign t[11142] = t[11141] ^ n[11142];
assign t[11143] = t[11142] ^ n[11143];
assign t[11144] = t[11143] ^ n[11144];
assign t[11145] = t[11144] ^ n[11145];
assign t[11146] = t[11145] ^ n[11146];
assign t[11147] = t[11146] ^ n[11147];
assign t[11148] = t[11147] ^ n[11148];
assign t[11149] = t[11148] ^ n[11149];
assign t[11150] = t[11149] ^ n[11150];
assign t[11151] = t[11150] ^ n[11151];
assign t[11152] = t[11151] ^ n[11152];
assign t[11153] = t[11152] ^ n[11153];
assign t[11154] = t[11153] ^ n[11154];
assign t[11155] = t[11154] ^ n[11155];
assign t[11156] = t[11155] ^ n[11156];
assign t[11157] = t[11156] ^ n[11157];
assign t[11158] = t[11157] ^ n[11158];
assign t[11159] = t[11158] ^ n[11159];
assign t[11160] = t[11159] ^ n[11160];
assign t[11161] = t[11160] ^ n[11161];
assign t[11162] = t[11161] ^ n[11162];
assign t[11163] = t[11162] ^ n[11163];
assign t[11164] = t[11163] ^ n[11164];
assign t[11165] = t[11164] ^ n[11165];
assign t[11166] = t[11165] ^ n[11166];
assign t[11167] = t[11166] ^ n[11167];
assign t[11168] = t[11167] ^ n[11168];
assign t[11169] = t[11168] ^ n[11169];
assign t[11170] = t[11169] ^ n[11170];
assign t[11171] = t[11170] ^ n[11171];
assign t[11172] = t[11171] ^ n[11172];
assign t[11173] = t[11172] ^ n[11173];
assign t[11174] = t[11173] ^ n[11174];
assign t[11175] = t[11174] ^ n[11175];
assign t[11176] = t[11175] ^ n[11176];
assign t[11177] = t[11176] ^ n[11177];
assign t[11178] = t[11177] ^ n[11178];
assign t[11179] = t[11178] ^ n[11179];
assign t[11180] = t[11179] ^ n[11180];
assign t[11181] = t[11180] ^ n[11181];
assign t[11182] = t[11181] ^ n[11182];
assign t[11183] = t[11182] ^ n[11183];
assign t[11184] = t[11183] ^ n[11184];
assign t[11185] = t[11184] ^ n[11185];
assign t[11186] = t[11185] ^ n[11186];
assign t[11187] = t[11186] ^ n[11187];
assign t[11188] = t[11187] ^ n[11188];
assign t[11189] = t[11188] ^ n[11189];
assign t[11190] = t[11189] ^ n[11190];
assign t[11191] = t[11190] ^ n[11191];
assign t[11192] = t[11191] ^ n[11192];
assign t[11193] = t[11192] ^ n[11193];
assign t[11194] = t[11193] ^ n[11194];
assign t[11195] = t[11194] ^ n[11195];
assign t[11196] = t[11195] ^ n[11196];
assign t[11197] = t[11196] ^ n[11197];
assign t[11198] = t[11197] ^ n[11198];
assign t[11199] = t[11198] ^ n[11199];
assign t[11200] = t[11199] ^ n[11200];
assign t[11201] = t[11200] ^ n[11201];
assign t[11202] = t[11201] ^ n[11202];
assign t[11203] = t[11202] ^ n[11203];
assign t[11204] = t[11203] ^ n[11204];
assign t[11205] = t[11204] ^ n[11205];
assign t[11206] = t[11205] ^ n[11206];
assign t[11207] = t[11206] ^ n[11207];
assign t[11208] = t[11207] ^ n[11208];
assign t[11209] = t[11208] ^ n[11209];
assign t[11210] = t[11209] ^ n[11210];
assign t[11211] = t[11210] ^ n[11211];
assign t[11212] = t[11211] ^ n[11212];
assign t[11213] = t[11212] ^ n[11213];
assign t[11214] = t[11213] ^ n[11214];
assign t[11215] = t[11214] ^ n[11215];
assign t[11216] = t[11215] ^ n[11216];
assign t[11217] = t[11216] ^ n[11217];
assign t[11218] = t[11217] ^ n[11218];
assign t[11219] = t[11218] ^ n[11219];
assign t[11220] = t[11219] ^ n[11220];
assign t[11221] = t[11220] ^ n[11221];
assign t[11222] = t[11221] ^ n[11222];
assign t[11223] = t[11222] ^ n[11223];
assign t[11224] = t[11223] ^ n[11224];
assign t[11225] = t[11224] ^ n[11225];
assign t[11226] = t[11225] ^ n[11226];
assign t[11227] = t[11226] ^ n[11227];
assign t[11228] = t[11227] ^ n[11228];
assign t[11229] = t[11228] ^ n[11229];
assign t[11230] = t[11229] ^ n[11230];
assign t[11231] = t[11230] ^ n[11231];
assign t[11232] = t[11231] ^ n[11232];
assign t[11233] = t[11232] ^ n[11233];
assign t[11234] = t[11233] ^ n[11234];
assign t[11235] = t[11234] ^ n[11235];
assign t[11236] = t[11235] ^ n[11236];
assign t[11237] = t[11236] ^ n[11237];
assign t[11238] = t[11237] ^ n[11238];
assign t[11239] = t[11238] ^ n[11239];
assign t[11240] = t[11239] ^ n[11240];
assign t[11241] = t[11240] ^ n[11241];
assign t[11242] = t[11241] ^ n[11242];
assign t[11243] = t[11242] ^ n[11243];
assign t[11244] = t[11243] ^ n[11244];
assign t[11245] = t[11244] ^ n[11245];
assign t[11246] = t[11245] ^ n[11246];
assign t[11247] = t[11246] ^ n[11247];
assign t[11248] = t[11247] ^ n[11248];
assign t[11249] = t[11248] ^ n[11249];
assign t[11250] = t[11249] ^ n[11250];
assign t[11251] = t[11250] ^ n[11251];
assign t[11252] = t[11251] ^ n[11252];
assign t[11253] = t[11252] ^ n[11253];
assign t[11254] = t[11253] ^ n[11254];
assign t[11255] = t[11254] ^ n[11255];
assign t[11256] = t[11255] ^ n[11256];
assign t[11257] = t[11256] ^ n[11257];
assign t[11258] = t[11257] ^ n[11258];
assign t[11259] = t[11258] ^ n[11259];
assign t[11260] = t[11259] ^ n[11260];
assign t[11261] = t[11260] ^ n[11261];
assign t[11262] = t[11261] ^ n[11262];
assign t[11263] = t[11262] ^ n[11263];
assign t[11264] = t[11263] ^ n[11264];
assign t[11265] = t[11264] ^ n[11265];
assign t[11266] = t[11265] ^ n[11266];
assign t[11267] = t[11266] ^ n[11267];
assign t[11268] = t[11267] ^ n[11268];
assign t[11269] = t[11268] ^ n[11269];
assign t[11270] = t[11269] ^ n[11270];
assign t[11271] = t[11270] ^ n[11271];
assign t[11272] = t[11271] ^ n[11272];
assign t[11273] = t[11272] ^ n[11273];
assign t[11274] = t[11273] ^ n[11274];
assign t[11275] = t[11274] ^ n[11275];
assign t[11276] = t[11275] ^ n[11276];
assign t[11277] = t[11276] ^ n[11277];
assign t[11278] = t[11277] ^ n[11278];
assign t[11279] = t[11278] ^ n[11279];
assign t[11280] = t[11279] ^ n[11280];
assign t[11281] = t[11280] ^ n[11281];
assign t[11282] = t[11281] ^ n[11282];
assign t[11283] = t[11282] ^ n[11283];
assign t[11284] = t[11283] ^ n[11284];
assign t[11285] = t[11284] ^ n[11285];
assign t[11286] = t[11285] ^ n[11286];
assign t[11287] = t[11286] ^ n[11287];
assign t[11288] = t[11287] ^ n[11288];
assign t[11289] = t[11288] ^ n[11289];
assign t[11290] = t[11289] ^ n[11290];
assign t[11291] = t[11290] ^ n[11291];
assign t[11292] = t[11291] ^ n[11292];
assign t[11293] = t[11292] ^ n[11293];
assign t[11294] = t[11293] ^ n[11294];
assign t[11295] = t[11294] ^ n[11295];
assign t[11296] = t[11295] ^ n[11296];
assign t[11297] = t[11296] ^ n[11297];
assign t[11298] = t[11297] ^ n[11298];
assign t[11299] = t[11298] ^ n[11299];
assign t[11300] = t[11299] ^ n[11300];
assign t[11301] = t[11300] ^ n[11301];
assign t[11302] = t[11301] ^ n[11302];
assign t[11303] = t[11302] ^ n[11303];
assign t[11304] = t[11303] ^ n[11304];
assign t[11305] = t[11304] ^ n[11305];
assign t[11306] = t[11305] ^ n[11306];
assign t[11307] = t[11306] ^ n[11307];
assign t[11308] = t[11307] ^ n[11308];
assign t[11309] = t[11308] ^ n[11309];
assign t[11310] = t[11309] ^ n[11310];
assign t[11311] = t[11310] ^ n[11311];
assign t[11312] = t[11311] ^ n[11312];
assign t[11313] = t[11312] ^ n[11313];
assign t[11314] = t[11313] ^ n[11314];
assign t[11315] = t[11314] ^ n[11315];
assign t[11316] = t[11315] ^ n[11316];
assign t[11317] = t[11316] ^ n[11317];
assign t[11318] = t[11317] ^ n[11318];
assign t[11319] = t[11318] ^ n[11319];
assign t[11320] = t[11319] ^ n[11320];
assign t[11321] = t[11320] ^ n[11321];
assign t[11322] = t[11321] ^ n[11322];
assign t[11323] = t[11322] ^ n[11323];
assign t[11324] = t[11323] ^ n[11324];
assign t[11325] = t[11324] ^ n[11325];
assign t[11326] = t[11325] ^ n[11326];
assign t[11327] = t[11326] ^ n[11327];
assign t[11328] = t[11327] ^ n[11328];
assign t[11329] = t[11328] ^ n[11329];
assign t[11330] = t[11329] ^ n[11330];
assign t[11331] = t[11330] ^ n[11331];
assign t[11332] = t[11331] ^ n[11332];
assign t[11333] = t[11332] ^ n[11333];
assign t[11334] = t[11333] ^ n[11334];
assign t[11335] = t[11334] ^ n[11335];
assign t[11336] = t[11335] ^ n[11336];
assign t[11337] = t[11336] ^ n[11337];
assign t[11338] = t[11337] ^ n[11338];
assign t[11339] = t[11338] ^ n[11339];
assign t[11340] = t[11339] ^ n[11340];
assign t[11341] = t[11340] ^ n[11341];
assign t[11342] = t[11341] ^ n[11342];
assign t[11343] = t[11342] ^ n[11343];
assign t[11344] = t[11343] ^ n[11344];
assign t[11345] = t[11344] ^ n[11345];
assign t[11346] = t[11345] ^ n[11346];
assign t[11347] = t[11346] ^ n[11347];
assign t[11348] = t[11347] ^ n[11348];
assign t[11349] = t[11348] ^ n[11349];
assign t[11350] = t[11349] ^ n[11350];
assign t[11351] = t[11350] ^ n[11351];
assign t[11352] = t[11351] ^ n[11352];
assign t[11353] = t[11352] ^ n[11353];
assign t[11354] = t[11353] ^ n[11354];
assign t[11355] = t[11354] ^ n[11355];
assign t[11356] = t[11355] ^ n[11356];
assign t[11357] = t[11356] ^ n[11357];
assign t[11358] = t[11357] ^ n[11358];
assign t[11359] = t[11358] ^ n[11359];
assign t[11360] = t[11359] ^ n[11360];
assign t[11361] = t[11360] ^ n[11361];
assign t[11362] = t[11361] ^ n[11362];
assign t[11363] = t[11362] ^ n[11363];
assign t[11364] = t[11363] ^ n[11364];
assign t[11365] = t[11364] ^ n[11365];
assign t[11366] = t[11365] ^ n[11366];
assign t[11367] = t[11366] ^ n[11367];
assign t[11368] = t[11367] ^ n[11368];
assign t[11369] = t[11368] ^ n[11369];
assign t[11370] = t[11369] ^ n[11370];
assign t[11371] = t[11370] ^ n[11371];
assign t[11372] = t[11371] ^ n[11372];
assign t[11373] = t[11372] ^ n[11373];
assign t[11374] = t[11373] ^ n[11374];
assign t[11375] = t[11374] ^ n[11375];
assign t[11376] = t[11375] ^ n[11376];
assign t[11377] = t[11376] ^ n[11377];
assign t[11378] = t[11377] ^ n[11378];
assign t[11379] = t[11378] ^ n[11379];
assign t[11380] = t[11379] ^ n[11380];
assign t[11381] = t[11380] ^ n[11381];
assign t[11382] = t[11381] ^ n[11382];
assign t[11383] = t[11382] ^ n[11383];
assign t[11384] = t[11383] ^ n[11384];
assign t[11385] = t[11384] ^ n[11385];
assign t[11386] = t[11385] ^ n[11386];
assign t[11387] = t[11386] ^ n[11387];
assign t[11388] = t[11387] ^ n[11388];
assign t[11389] = t[11388] ^ n[11389];
assign t[11390] = t[11389] ^ n[11390];
assign t[11391] = t[11390] ^ n[11391];
assign t[11392] = t[11391] ^ n[11392];
assign t[11393] = t[11392] ^ n[11393];
assign t[11394] = t[11393] ^ n[11394];
assign t[11395] = t[11394] ^ n[11395];
assign t[11396] = t[11395] ^ n[11396];
assign t[11397] = t[11396] ^ n[11397];
assign t[11398] = t[11397] ^ n[11398];
assign t[11399] = t[11398] ^ n[11399];
assign t[11400] = t[11399] ^ n[11400];
assign t[11401] = t[11400] ^ n[11401];
assign t[11402] = t[11401] ^ n[11402];
assign t[11403] = t[11402] ^ n[11403];
assign t[11404] = t[11403] ^ n[11404];
assign t[11405] = t[11404] ^ n[11405];
assign t[11406] = t[11405] ^ n[11406];
assign t[11407] = t[11406] ^ n[11407];
assign t[11408] = t[11407] ^ n[11408];
assign t[11409] = t[11408] ^ n[11409];
assign t[11410] = t[11409] ^ n[11410];
assign t[11411] = t[11410] ^ n[11411];
assign t[11412] = t[11411] ^ n[11412];
assign t[11413] = t[11412] ^ n[11413];
assign t[11414] = t[11413] ^ n[11414];
assign t[11415] = t[11414] ^ n[11415];
assign t[11416] = t[11415] ^ n[11416];
assign t[11417] = t[11416] ^ n[11417];
assign t[11418] = t[11417] ^ n[11418];
assign t[11419] = t[11418] ^ n[11419];
assign t[11420] = t[11419] ^ n[11420];
assign t[11421] = t[11420] ^ n[11421];
assign t[11422] = t[11421] ^ n[11422];
assign t[11423] = t[11422] ^ n[11423];
assign t[11424] = t[11423] ^ n[11424];
assign t[11425] = t[11424] ^ n[11425];
assign t[11426] = t[11425] ^ n[11426];
assign t[11427] = t[11426] ^ n[11427];
assign t[11428] = t[11427] ^ n[11428];
assign t[11429] = t[11428] ^ n[11429];
assign t[11430] = t[11429] ^ n[11430];
assign t[11431] = t[11430] ^ n[11431];
assign t[11432] = t[11431] ^ n[11432];
assign t[11433] = t[11432] ^ n[11433];
assign t[11434] = t[11433] ^ n[11434];
assign t[11435] = t[11434] ^ n[11435];
assign t[11436] = t[11435] ^ n[11436];
assign t[11437] = t[11436] ^ n[11437];
assign t[11438] = t[11437] ^ n[11438];
assign t[11439] = t[11438] ^ n[11439];
assign t[11440] = t[11439] ^ n[11440];
assign t[11441] = t[11440] ^ n[11441];
assign t[11442] = t[11441] ^ n[11442];
assign t[11443] = t[11442] ^ n[11443];
assign t[11444] = t[11443] ^ n[11444];
assign t[11445] = t[11444] ^ n[11445];
assign t[11446] = t[11445] ^ n[11446];
assign t[11447] = t[11446] ^ n[11447];
assign t[11448] = t[11447] ^ n[11448];
assign t[11449] = t[11448] ^ n[11449];
assign t[11450] = t[11449] ^ n[11450];
assign t[11451] = t[11450] ^ n[11451];
assign t[11452] = t[11451] ^ n[11452];
assign t[11453] = t[11452] ^ n[11453];
assign t[11454] = t[11453] ^ n[11454];
assign t[11455] = t[11454] ^ n[11455];
assign t[11456] = t[11455] ^ n[11456];
assign t[11457] = t[11456] ^ n[11457];
assign t[11458] = t[11457] ^ n[11458];
assign t[11459] = t[11458] ^ n[11459];
assign t[11460] = t[11459] ^ n[11460];
assign t[11461] = t[11460] ^ n[11461];
assign t[11462] = t[11461] ^ n[11462];
assign t[11463] = t[11462] ^ n[11463];
assign t[11464] = t[11463] ^ n[11464];
assign t[11465] = t[11464] ^ n[11465];
assign t[11466] = t[11465] ^ n[11466];
assign t[11467] = t[11466] ^ n[11467];
assign t[11468] = t[11467] ^ n[11468];
assign t[11469] = t[11468] ^ n[11469];
assign t[11470] = t[11469] ^ n[11470];
assign t[11471] = t[11470] ^ n[11471];
assign t[11472] = t[11471] ^ n[11472];
assign t[11473] = t[11472] ^ n[11473];
assign t[11474] = t[11473] ^ n[11474];
assign t[11475] = t[11474] ^ n[11475];
assign t[11476] = t[11475] ^ n[11476];
assign t[11477] = t[11476] ^ n[11477];
assign t[11478] = t[11477] ^ n[11478];
assign t[11479] = t[11478] ^ n[11479];
assign t[11480] = t[11479] ^ n[11480];
assign t[11481] = t[11480] ^ n[11481];
assign t[11482] = t[11481] ^ n[11482];
assign t[11483] = t[11482] ^ n[11483];
assign t[11484] = t[11483] ^ n[11484];
assign t[11485] = t[11484] ^ n[11485];
assign t[11486] = t[11485] ^ n[11486];
assign t[11487] = t[11486] ^ n[11487];
assign t[11488] = t[11487] ^ n[11488];
assign t[11489] = t[11488] ^ n[11489];
assign t[11490] = t[11489] ^ n[11490];
assign t[11491] = t[11490] ^ n[11491];
assign t[11492] = t[11491] ^ n[11492];
assign t[11493] = t[11492] ^ n[11493];
assign t[11494] = t[11493] ^ n[11494];
assign t[11495] = t[11494] ^ n[11495];
assign t[11496] = t[11495] ^ n[11496];
assign t[11497] = t[11496] ^ n[11497];
assign t[11498] = t[11497] ^ n[11498];
assign t[11499] = t[11498] ^ n[11499];
assign t[11500] = t[11499] ^ n[11500];
assign t[11501] = t[11500] ^ n[11501];
assign t[11502] = t[11501] ^ n[11502];
assign t[11503] = t[11502] ^ n[11503];
assign t[11504] = t[11503] ^ n[11504];
assign t[11505] = t[11504] ^ n[11505];
assign t[11506] = t[11505] ^ n[11506];
assign t[11507] = t[11506] ^ n[11507];
assign t[11508] = t[11507] ^ n[11508];
assign t[11509] = t[11508] ^ n[11509];
assign t[11510] = t[11509] ^ n[11510];
assign t[11511] = t[11510] ^ n[11511];
assign t[11512] = t[11511] ^ n[11512];
assign t[11513] = t[11512] ^ n[11513];
assign t[11514] = t[11513] ^ n[11514];
assign t[11515] = t[11514] ^ n[11515];
assign t[11516] = t[11515] ^ n[11516];
assign t[11517] = t[11516] ^ n[11517];
assign t[11518] = t[11517] ^ n[11518];
assign t[11519] = t[11518] ^ n[11519];
assign t[11520] = t[11519] ^ n[11520];
assign t[11521] = t[11520] ^ n[11521];
assign t[11522] = t[11521] ^ n[11522];
assign t[11523] = t[11522] ^ n[11523];
assign t[11524] = t[11523] ^ n[11524];
assign t[11525] = t[11524] ^ n[11525];
assign t[11526] = t[11525] ^ n[11526];
assign t[11527] = t[11526] ^ n[11527];
assign t[11528] = t[11527] ^ n[11528];
assign t[11529] = t[11528] ^ n[11529];
assign t[11530] = t[11529] ^ n[11530];
assign t[11531] = t[11530] ^ n[11531];
assign t[11532] = t[11531] ^ n[11532];
assign t[11533] = t[11532] ^ n[11533];
assign t[11534] = t[11533] ^ n[11534];
assign t[11535] = t[11534] ^ n[11535];
assign t[11536] = t[11535] ^ n[11536];
assign t[11537] = t[11536] ^ n[11537];
assign t[11538] = t[11537] ^ n[11538];
assign t[11539] = t[11538] ^ n[11539];
assign t[11540] = t[11539] ^ n[11540];
assign t[11541] = t[11540] ^ n[11541];
assign t[11542] = t[11541] ^ n[11542];
assign t[11543] = t[11542] ^ n[11543];
assign t[11544] = t[11543] ^ n[11544];
assign t[11545] = t[11544] ^ n[11545];
assign t[11546] = t[11545] ^ n[11546];
assign t[11547] = t[11546] ^ n[11547];
assign t[11548] = t[11547] ^ n[11548];
assign t[11549] = t[11548] ^ n[11549];
assign t[11550] = t[11549] ^ n[11550];
assign t[11551] = t[11550] ^ n[11551];
assign t[11552] = t[11551] ^ n[11552];
assign t[11553] = t[11552] ^ n[11553];
assign t[11554] = t[11553] ^ n[11554];
assign t[11555] = t[11554] ^ n[11555];
assign t[11556] = t[11555] ^ n[11556];
assign t[11557] = t[11556] ^ n[11557];
assign t[11558] = t[11557] ^ n[11558];
assign t[11559] = t[11558] ^ n[11559];
assign t[11560] = t[11559] ^ n[11560];
assign t[11561] = t[11560] ^ n[11561];
assign t[11562] = t[11561] ^ n[11562];
assign t[11563] = t[11562] ^ n[11563];
assign t[11564] = t[11563] ^ n[11564];
assign t[11565] = t[11564] ^ n[11565];
assign t[11566] = t[11565] ^ n[11566];
assign t[11567] = t[11566] ^ n[11567];
assign t[11568] = t[11567] ^ n[11568];
assign t[11569] = t[11568] ^ n[11569];
assign t[11570] = t[11569] ^ n[11570];
assign t[11571] = t[11570] ^ n[11571];
assign t[11572] = t[11571] ^ n[11572];
assign t[11573] = t[11572] ^ n[11573];
assign t[11574] = t[11573] ^ n[11574];
assign t[11575] = t[11574] ^ n[11575];
assign t[11576] = t[11575] ^ n[11576];
assign t[11577] = t[11576] ^ n[11577];
assign t[11578] = t[11577] ^ n[11578];
assign t[11579] = t[11578] ^ n[11579];
assign t[11580] = t[11579] ^ n[11580];
assign t[11581] = t[11580] ^ n[11581];
assign t[11582] = t[11581] ^ n[11582];
assign t[11583] = t[11582] ^ n[11583];
assign t[11584] = t[11583] ^ n[11584];
assign t[11585] = t[11584] ^ n[11585];
assign t[11586] = t[11585] ^ n[11586];
assign t[11587] = t[11586] ^ n[11587];
assign t[11588] = t[11587] ^ n[11588];
assign t[11589] = t[11588] ^ n[11589];
assign t[11590] = t[11589] ^ n[11590];
assign t[11591] = t[11590] ^ n[11591];
assign t[11592] = t[11591] ^ n[11592];
assign t[11593] = t[11592] ^ n[11593];
assign t[11594] = t[11593] ^ n[11594];
assign t[11595] = t[11594] ^ n[11595];
assign t[11596] = t[11595] ^ n[11596];
assign t[11597] = t[11596] ^ n[11597];
assign t[11598] = t[11597] ^ n[11598];
assign t[11599] = t[11598] ^ n[11599];
assign t[11600] = t[11599] ^ n[11600];
assign t[11601] = t[11600] ^ n[11601];
assign t[11602] = t[11601] ^ n[11602];
assign t[11603] = t[11602] ^ n[11603];
assign t[11604] = t[11603] ^ n[11604];
assign t[11605] = t[11604] ^ n[11605];
assign t[11606] = t[11605] ^ n[11606];
assign t[11607] = t[11606] ^ n[11607];
assign t[11608] = t[11607] ^ n[11608];
assign t[11609] = t[11608] ^ n[11609];
assign t[11610] = t[11609] ^ n[11610];
assign t[11611] = t[11610] ^ n[11611];
assign t[11612] = t[11611] ^ n[11612];
assign t[11613] = t[11612] ^ n[11613];
assign t[11614] = t[11613] ^ n[11614];
assign t[11615] = t[11614] ^ n[11615];
assign t[11616] = t[11615] ^ n[11616];
assign t[11617] = t[11616] ^ n[11617];
assign t[11618] = t[11617] ^ n[11618];
assign t[11619] = t[11618] ^ n[11619];
assign t[11620] = t[11619] ^ n[11620];
assign t[11621] = t[11620] ^ n[11621];
assign t[11622] = t[11621] ^ n[11622];
assign t[11623] = t[11622] ^ n[11623];
assign t[11624] = t[11623] ^ n[11624];
assign t[11625] = t[11624] ^ n[11625];
assign t[11626] = t[11625] ^ n[11626];
assign t[11627] = t[11626] ^ n[11627];
assign t[11628] = t[11627] ^ n[11628];
assign t[11629] = t[11628] ^ n[11629];
assign t[11630] = t[11629] ^ n[11630];
assign t[11631] = t[11630] ^ n[11631];
assign t[11632] = t[11631] ^ n[11632];
assign t[11633] = t[11632] ^ n[11633];
assign t[11634] = t[11633] ^ n[11634];
assign t[11635] = t[11634] ^ n[11635];
assign t[11636] = t[11635] ^ n[11636];
assign t[11637] = t[11636] ^ n[11637];
assign t[11638] = t[11637] ^ n[11638];
assign t[11639] = t[11638] ^ n[11639];
assign t[11640] = t[11639] ^ n[11640];
assign t[11641] = t[11640] ^ n[11641];
assign t[11642] = t[11641] ^ n[11642];
assign t[11643] = t[11642] ^ n[11643];
assign t[11644] = t[11643] ^ n[11644];
assign t[11645] = t[11644] ^ n[11645];
assign t[11646] = t[11645] ^ n[11646];
assign t[11647] = t[11646] ^ n[11647];
assign t[11648] = t[11647] ^ n[11648];
assign t[11649] = t[11648] ^ n[11649];
assign t[11650] = t[11649] ^ n[11650];
assign t[11651] = t[11650] ^ n[11651];
assign t[11652] = t[11651] ^ n[11652];
assign t[11653] = t[11652] ^ n[11653];
assign t[11654] = t[11653] ^ n[11654];
assign t[11655] = t[11654] ^ n[11655];
assign t[11656] = t[11655] ^ n[11656];
assign t[11657] = t[11656] ^ n[11657];
assign t[11658] = t[11657] ^ n[11658];
assign t[11659] = t[11658] ^ n[11659];
assign t[11660] = t[11659] ^ n[11660];
assign t[11661] = t[11660] ^ n[11661];
assign t[11662] = t[11661] ^ n[11662];
assign t[11663] = t[11662] ^ n[11663];
assign t[11664] = t[11663] ^ n[11664];
assign t[11665] = t[11664] ^ n[11665];
assign t[11666] = t[11665] ^ n[11666];
assign t[11667] = t[11666] ^ n[11667];
assign t[11668] = t[11667] ^ n[11668];
assign t[11669] = t[11668] ^ n[11669];
assign t[11670] = t[11669] ^ n[11670];
assign t[11671] = t[11670] ^ n[11671];
assign t[11672] = t[11671] ^ n[11672];
assign t[11673] = t[11672] ^ n[11673];
assign t[11674] = t[11673] ^ n[11674];
assign t[11675] = t[11674] ^ n[11675];
assign t[11676] = t[11675] ^ n[11676];
assign t[11677] = t[11676] ^ n[11677];
assign t[11678] = t[11677] ^ n[11678];
assign t[11679] = t[11678] ^ n[11679];
assign t[11680] = t[11679] ^ n[11680];
assign t[11681] = t[11680] ^ n[11681];
assign t[11682] = t[11681] ^ n[11682];
assign t[11683] = t[11682] ^ n[11683];
assign t[11684] = t[11683] ^ n[11684];
assign t[11685] = t[11684] ^ n[11685];
assign t[11686] = t[11685] ^ n[11686];
assign t[11687] = t[11686] ^ n[11687];
assign t[11688] = t[11687] ^ n[11688];
assign t[11689] = t[11688] ^ n[11689];
assign t[11690] = t[11689] ^ n[11690];
assign t[11691] = t[11690] ^ n[11691];
assign t[11692] = t[11691] ^ n[11692];
assign t[11693] = t[11692] ^ n[11693];
assign t[11694] = t[11693] ^ n[11694];
assign t[11695] = t[11694] ^ n[11695];
assign t[11696] = t[11695] ^ n[11696];
assign t[11697] = t[11696] ^ n[11697];
assign t[11698] = t[11697] ^ n[11698];
assign t[11699] = t[11698] ^ n[11699];
assign t[11700] = t[11699] ^ n[11700];
assign t[11701] = t[11700] ^ n[11701];
assign t[11702] = t[11701] ^ n[11702];
assign t[11703] = t[11702] ^ n[11703];
assign t[11704] = t[11703] ^ n[11704];
assign t[11705] = t[11704] ^ n[11705];
assign t[11706] = t[11705] ^ n[11706];
assign t[11707] = t[11706] ^ n[11707];
assign t[11708] = t[11707] ^ n[11708];
assign t[11709] = t[11708] ^ n[11709];
assign t[11710] = t[11709] ^ n[11710];
assign t[11711] = t[11710] ^ n[11711];
assign t[11712] = t[11711] ^ n[11712];
assign t[11713] = t[11712] ^ n[11713];
assign t[11714] = t[11713] ^ n[11714];
assign t[11715] = t[11714] ^ n[11715];
assign t[11716] = t[11715] ^ n[11716];
assign t[11717] = t[11716] ^ n[11717];
assign t[11718] = t[11717] ^ n[11718];
assign t[11719] = t[11718] ^ n[11719];
assign t[11720] = t[11719] ^ n[11720];
assign t[11721] = t[11720] ^ n[11721];
assign t[11722] = t[11721] ^ n[11722];
assign t[11723] = t[11722] ^ n[11723];
assign t[11724] = t[11723] ^ n[11724];
assign t[11725] = t[11724] ^ n[11725];
assign t[11726] = t[11725] ^ n[11726];
assign t[11727] = t[11726] ^ n[11727];
assign t[11728] = t[11727] ^ n[11728];
assign t[11729] = t[11728] ^ n[11729];
assign t[11730] = t[11729] ^ n[11730];
assign t[11731] = t[11730] ^ n[11731];
assign t[11732] = t[11731] ^ n[11732];
assign t[11733] = t[11732] ^ n[11733];
assign t[11734] = t[11733] ^ n[11734];
assign t[11735] = t[11734] ^ n[11735];
assign t[11736] = t[11735] ^ n[11736];
assign t[11737] = t[11736] ^ n[11737];
assign t[11738] = t[11737] ^ n[11738];
assign t[11739] = t[11738] ^ n[11739];
assign t[11740] = t[11739] ^ n[11740];
assign t[11741] = t[11740] ^ n[11741];
assign t[11742] = t[11741] ^ n[11742];
assign t[11743] = t[11742] ^ n[11743];
assign t[11744] = t[11743] ^ n[11744];
assign t[11745] = t[11744] ^ n[11745];
assign t[11746] = t[11745] ^ n[11746];
assign t[11747] = t[11746] ^ n[11747];
assign t[11748] = t[11747] ^ n[11748];
assign t[11749] = t[11748] ^ n[11749];
assign t[11750] = t[11749] ^ n[11750];
assign t[11751] = t[11750] ^ n[11751];
assign t[11752] = t[11751] ^ n[11752];
assign t[11753] = t[11752] ^ n[11753];
assign t[11754] = t[11753] ^ n[11754];
assign t[11755] = t[11754] ^ n[11755];
assign t[11756] = t[11755] ^ n[11756];
assign t[11757] = t[11756] ^ n[11757];
assign t[11758] = t[11757] ^ n[11758];
assign t[11759] = t[11758] ^ n[11759];
assign t[11760] = t[11759] ^ n[11760];
assign t[11761] = t[11760] ^ n[11761];
assign t[11762] = t[11761] ^ n[11762];
assign t[11763] = t[11762] ^ n[11763];
assign t[11764] = t[11763] ^ n[11764];
assign t[11765] = t[11764] ^ n[11765];
assign t[11766] = t[11765] ^ n[11766];
assign t[11767] = t[11766] ^ n[11767];
assign t[11768] = t[11767] ^ n[11768];
assign t[11769] = t[11768] ^ n[11769];
assign t[11770] = t[11769] ^ n[11770];
assign t[11771] = t[11770] ^ n[11771];
assign t[11772] = t[11771] ^ n[11772];
assign t[11773] = t[11772] ^ n[11773];
assign t[11774] = t[11773] ^ n[11774];
assign t[11775] = t[11774] ^ n[11775];
assign t[11776] = t[11775] ^ n[11776];
assign t[11777] = t[11776] ^ n[11777];
assign t[11778] = t[11777] ^ n[11778];
assign t[11779] = t[11778] ^ n[11779];
assign t[11780] = t[11779] ^ n[11780];
assign t[11781] = t[11780] ^ n[11781];
assign t[11782] = t[11781] ^ n[11782];
assign t[11783] = t[11782] ^ n[11783];
assign t[11784] = t[11783] ^ n[11784];
assign t[11785] = t[11784] ^ n[11785];
assign t[11786] = t[11785] ^ n[11786];
assign t[11787] = t[11786] ^ n[11787];
assign t[11788] = t[11787] ^ n[11788];
assign t[11789] = t[11788] ^ n[11789];
assign t[11790] = t[11789] ^ n[11790];
assign t[11791] = t[11790] ^ n[11791];
assign t[11792] = t[11791] ^ n[11792];
assign t[11793] = t[11792] ^ n[11793];
assign t[11794] = t[11793] ^ n[11794];
assign t[11795] = t[11794] ^ n[11795];
assign t[11796] = t[11795] ^ n[11796];
assign t[11797] = t[11796] ^ n[11797];
assign t[11798] = t[11797] ^ n[11798];
assign t[11799] = t[11798] ^ n[11799];
assign t[11800] = t[11799] ^ n[11800];
assign t[11801] = t[11800] ^ n[11801];
assign t[11802] = t[11801] ^ n[11802];
assign t[11803] = t[11802] ^ n[11803];
assign t[11804] = t[11803] ^ n[11804];
assign t[11805] = t[11804] ^ n[11805];
assign t[11806] = t[11805] ^ n[11806];
assign t[11807] = t[11806] ^ n[11807];
assign t[11808] = t[11807] ^ n[11808];
assign t[11809] = t[11808] ^ n[11809];
assign t[11810] = t[11809] ^ n[11810];
assign t[11811] = t[11810] ^ n[11811];
assign t[11812] = t[11811] ^ n[11812];
assign t[11813] = t[11812] ^ n[11813];
assign t[11814] = t[11813] ^ n[11814];
assign t[11815] = t[11814] ^ n[11815];
assign t[11816] = t[11815] ^ n[11816];
assign t[11817] = t[11816] ^ n[11817];
assign t[11818] = t[11817] ^ n[11818];
assign t[11819] = t[11818] ^ n[11819];
assign t[11820] = t[11819] ^ n[11820];
assign t[11821] = t[11820] ^ n[11821];
assign t[11822] = t[11821] ^ n[11822];
assign t[11823] = t[11822] ^ n[11823];
assign t[11824] = t[11823] ^ n[11824];
assign t[11825] = t[11824] ^ n[11825];
assign t[11826] = t[11825] ^ n[11826];
assign t[11827] = t[11826] ^ n[11827];
assign t[11828] = t[11827] ^ n[11828];
assign t[11829] = t[11828] ^ n[11829];
assign t[11830] = t[11829] ^ n[11830];
assign t[11831] = t[11830] ^ n[11831];
assign t[11832] = t[11831] ^ n[11832];
assign t[11833] = t[11832] ^ n[11833];
assign t[11834] = t[11833] ^ n[11834];
assign t[11835] = t[11834] ^ n[11835];
assign t[11836] = t[11835] ^ n[11836];
assign t[11837] = t[11836] ^ n[11837];
assign t[11838] = t[11837] ^ n[11838];
assign t[11839] = t[11838] ^ n[11839];
assign t[11840] = t[11839] ^ n[11840];
assign t[11841] = t[11840] ^ n[11841];
assign t[11842] = t[11841] ^ n[11842];
assign t[11843] = t[11842] ^ n[11843];
assign t[11844] = t[11843] ^ n[11844];
assign t[11845] = t[11844] ^ n[11845];
assign t[11846] = t[11845] ^ n[11846];
assign t[11847] = t[11846] ^ n[11847];
assign t[11848] = t[11847] ^ n[11848];
assign t[11849] = t[11848] ^ n[11849];
assign t[11850] = t[11849] ^ n[11850];
assign t[11851] = t[11850] ^ n[11851];
assign t[11852] = t[11851] ^ n[11852];
assign t[11853] = t[11852] ^ n[11853];
assign t[11854] = t[11853] ^ n[11854];
assign t[11855] = t[11854] ^ n[11855];
assign t[11856] = t[11855] ^ n[11856];
assign t[11857] = t[11856] ^ n[11857];
assign t[11858] = t[11857] ^ n[11858];
assign t[11859] = t[11858] ^ n[11859];
assign t[11860] = t[11859] ^ n[11860];
assign t[11861] = t[11860] ^ n[11861];
assign t[11862] = t[11861] ^ n[11862];
assign t[11863] = t[11862] ^ n[11863];
assign t[11864] = t[11863] ^ n[11864];
assign t[11865] = t[11864] ^ n[11865];
assign t[11866] = t[11865] ^ n[11866];
assign t[11867] = t[11866] ^ n[11867];
assign t[11868] = t[11867] ^ n[11868];
assign t[11869] = t[11868] ^ n[11869];
assign t[11870] = t[11869] ^ n[11870];
assign t[11871] = t[11870] ^ n[11871];
assign t[11872] = t[11871] ^ n[11872];
assign t[11873] = t[11872] ^ n[11873];
assign t[11874] = t[11873] ^ n[11874];
assign t[11875] = t[11874] ^ n[11875];
assign t[11876] = t[11875] ^ n[11876];
assign t[11877] = t[11876] ^ n[11877];
assign t[11878] = t[11877] ^ n[11878];
assign t[11879] = t[11878] ^ n[11879];
assign t[11880] = t[11879] ^ n[11880];
assign t[11881] = t[11880] ^ n[11881];
assign t[11882] = t[11881] ^ n[11882];
assign t[11883] = t[11882] ^ n[11883];
assign t[11884] = t[11883] ^ n[11884];
assign t[11885] = t[11884] ^ n[11885];
assign t[11886] = t[11885] ^ n[11886];
assign t[11887] = t[11886] ^ n[11887];
assign t[11888] = t[11887] ^ n[11888];
assign t[11889] = t[11888] ^ n[11889];
assign t[11890] = t[11889] ^ n[11890];
assign t[11891] = t[11890] ^ n[11891];
assign t[11892] = t[11891] ^ n[11892];
assign t[11893] = t[11892] ^ n[11893];
assign t[11894] = t[11893] ^ n[11894];
assign t[11895] = t[11894] ^ n[11895];
assign t[11896] = t[11895] ^ n[11896];
assign t[11897] = t[11896] ^ n[11897];
assign t[11898] = t[11897] ^ n[11898];
assign t[11899] = t[11898] ^ n[11899];
assign t[11900] = t[11899] ^ n[11900];
assign t[11901] = t[11900] ^ n[11901];
assign t[11902] = t[11901] ^ n[11902];
assign t[11903] = t[11902] ^ n[11903];
assign t[11904] = t[11903] ^ n[11904];
assign t[11905] = t[11904] ^ n[11905];
assign t[11906] = t[11905] ^ n[11906];
assign t[11907] = t[11906] ^ n[11907];
assign t[11908] = t[11907] ^ n[11908];
assign t[11909] = t[11908] ^ n[11909];
assign t[11910] = t[11909] ^ n[11910];
assign t[11911] = t[11910] ^ n[11911];
assign t[11912] = t[11911] ^ n[11912];
assign t[11913] = t[11912] ^ n[11913];
assign t[11914] = t[11913] ^ n[11914];
assign t[11915] = t[11914] ^ n[11915];
assign t[11916] = t[11915] ^ n[11916];
assign t[11917] = t[11916] ^ n[11917];
assign t[11918] = t[11917] ^ n[11918];
assign t[11919] = t[11918] ^ n[11919];
assign t[11920] = t[11919] ^ n[11920];
assign t[11921] = t[11920] ^ n[11921];
assign t[11922] = t[11921] ^ n[11922];
assign t[11923] = t[11922] ^ n[11923];
assign t[11924] = t[11923] ^ n[11924];
assign t[11925] = t[11924] ^ n[11925];
assign t[11926] = t[11925] ^ n[11926];
assign t[11927] = t[11926] ^ n[11927];
assign t[11928] = t[11927] ^ n[11928];
assign t[11929] = t[11928] ^ n[11929];
assign t[11930] = t[11929] ^ n[11930];
assign t[11931] = t[11930] ^ n[11931];
assign t[11932] = t[11931] ^ n[11932];
assign t[11933] = t[11932] ^ n[11933];
assign t[11934] = t[11933] ^ n[11934];
assign t[11935] = t[11934] ^ n[11935];
assign t[11936] = t[11935] ^ n[11936];
assign t[11937] = t[11936] ^ n[11937];
assign t[11938] = t[11937] ^ n[11938];
assign t[11939] = t[11938] ^ n[11939];
assign t[11940] = t[11939] ^ n[11940];
assign t[11941] = t[11940] ^ n[11941];
assign t[11942] = t[11941] ^ n[11942];
assign t[11943] = t[11942] ^ n[11943];
assign t[11944] = t[11943] ^ n[11944];
assign t[11945] = t[11944] ^ n[11945];
assign t[11946] = t[11945] ^ n[11946];
assign t[11947] = t[11946] ^ n[11947];
assign t[11948] = t[11947] ^ n[11948];
assign t[11949] = t[11948] ^ n[11949];
assign t[11950] = t[11949] ^ n[11950];
assign t[11951] = t[11950] ^ n[11951];
assign t[11952] = t[11951] ^ n[11952];
assign t[11953] = t[11952] ^ n[11953];
assign t[11954] = t[11953] ^ n[11954];
assign t[11955] = t[11954] ^ n[11955];
assign t[11956] = t[11955] ^ n[11956];
assign t[11957] = t[11956] ^ n[11957];
assign t[11958] = t[11957] ^ n[11958];
assign t[11959] = t[11958] ^ n[11959];
assign t[11960] = t[11959] ^ n[11960];
assign t[11961] = t[11960] ^ n[11961];
assign t[11962] = t[11961] ^ n[11962];
assign t[11963] = t[11962] ^ n[11963];
assign t[11964] = t[11963] ^ n[11964];
assign t[11965] = t[11964] ^ n[11965];
assign t[11966] = t[11965] ^ n[11966];
assign t[11967] = t[11966] ^ n[11967];
assign t[11968] = t[11967] ^ n[11968];
assign t[11969] = t[11968] ^ n[11969];
assign t[11970] = t[11969] ^ n[11970];
assign t[11971] = t[11970] ^ n[11971];
assign t[11972] = t[11971] ^ n[11972];
assign t[11973] = t[11972] ^ n[11973];
assign t[11974] = t[11973] ^ n[11974];
assign t[11975] = t[11974] ^ n[11975];
assign t[11976] = t[11975] ^ n[11976];
assign t[11977] = t[11976] ^ n[11977];
assign t[11978] = t[11977] ^ n[11978];
assign t[11979] = t[11978] ^ n[11979];
assign t[11980] = t[11979] ^ n[11980];
assign t[11981] = t[11980] ^ n[11981];
assign t[11982] = t[11981] ^ n[11982];
assign t[11983] = t[11982] ^ n[11983];
assign t[11984] = t[11983] ^ n[11984];
assign t[11985] = t[11984] ^ n[11985];
assign t[11986] = t[11985] ^ n[11986];
assign t[11987] = t[11986] ^ n[11987];
assign t[11988] = t[11987] ^ n[11988];
assign t[11989] = t[11988] ^ n[11989];
assign t[11990] = t[11989] ^ n[11990];
assign t[11991] = t[11990] ^ n[11991];
assign t[11992] = t[11991] ^ n[11992];
assign t[11993] = t[11992] ^ n[11993];
assign t[11994] = t[11993] ^ n[11994];
assign t[11995] = t[11994] ^ n[11995];
assign t[11996] = t[11995] ^ n[11996];
assign t[11997] = t[11996] ^ n[11997];
assign t[11998] = t[11997] ^ n[11998];
assign t[11999] = t[11998] ^ n[11999];
assign t[12000] = t[11999] ^ n[12000];
assign t[12001] = t[12000] ^ n[12001];
assign t[12002] = t[12001] ^ n[12002];
assign t[12003] = t[12002] ^ n[12003];
assign t[12004] = t[12003] ^ n[12004];
assign t[12005] = t[12004] ^ n[12005];
assign t[12006] = t[12005] ^ n[12006];
assign t[12007] = t[12006] ^ n[12007];
assign t[12008] = t[12007] ^ n[12008];
assign t[12009] = t[12008] ^ n[12009];
assign t[12010] = t[12009] ^ n[12010];
assign t[12011] = t[12010] ^ n[12011];
assign t[12012] = t[12011] ^ n[12012];
assign t[12013] = t[12012] ^ n[12013];
assign t[12014] = t[12013] ^ n[12014];
assign t[12015] = t[12014] ^ n[12015];
assign t[12016] = t[12015] ^ n[12016];
assign t[12017] = t[12016] ^ n[12017];
assign t[12018] = t[12017] ^ n[12018];
assign t[12019] = t[12018] ^ n[12019];
assign t[12020] = t[12019] ^ n[12020];
assign t[12021] = t[12020] ^ n[12021];
assign t[12022] = t[12021] ^ n[12022];
assign t[12023] = t[12022] ^ n[12023];
assign t[12024] = t[12023] ^ n[12024];
assign t[12025] = t[12024] ^ n[12025];
assign t[12026] = t[12025] ^ n[12026];
assign t[12027] = t[12026] ^ n[12027];
assign t[12028] = t[12027] ^ n[12028];
assign t[12029] = t[12028] ^ n[12029];
assign t[12030] = t[12029] ^ n[12030];
assign t[12031] = t[12030] ^ n[12031];
assign t[12032] = t[12031] ^ n[12032];
assign t[12033] = t[12032] ^ n[12033];
assign t[12034] = t[12033] ^ n[12034];
assign t[12035] = t[12034] ^ n[12035];
assign t[12036] = t[12035] ^ n[12036];
assign t[12037] = t[12036] ^ n[12037];
assign t[12038] = t[12037] ^ n[12038];
assign t[12039] = t[12038] ^ n[12039];
assign t[12040] = t[12039] ^ n[12040];
assign t[12041] = t[12040] ^ n[12041];
assign t[12042] = t[12041] ^ n[12042];
assign t[12043] = t[12042] ^ n[12043];
assign t[12044] = t[12043] ^ n[12044];
assign t[12045] = t[12044] ^ n[12045];
assign t[12046] = t[12045] ^ n[12046];
assign t[12047] = t[12046] ^ n[12047];
assign t[12048] = t[12047] ^ n[12048];
assign t[12049] = t[12048] ^ n[12049];
assign t[12050] = t[12049] ^ n[12050];
assign t[12051] = t[12050] ^ n[12051];
assign t[12052] = t[12051] ^ n[12052];
assign t[12053] = t[12052] ^ n[12053];
assign t[12054] = t[12053] ^ n[12054];
assign t[12055] = t[12054] ^ n[12055];
assign t[12056] = t[12055] ^ n[12056];
assign t[12057] = t[12056] ^ n[12057];
assign t[12058] = t[12057] ^ n[12058];
assign t[12059] = t[12058] ^ n[12059];
assign t[12060] = t[12059] ^ n[12060];
assign t[12061] = t[12060] ^ n[12061];
assign t[12062] = t[12061] ^ n[12062];
assign t[12063] = t[12062] ^ n[12063];
assign t[12064] = t[12063] ^ n[12064];
assign t[12065] = t[12064] ^ n[12065];
assign t[12066] = t[12065] ^ n[12066];
assign t[12067] = t[12066] ^ n[12067];
assign t[12068] = t[12067] ^ n[12068];
assign t[12069] = t[12068] ^ n[12069];
assign t[12070] = t[12069] ^ n[12070];
assign t[12071] = t[12070] ^ n[12071];
assign t[12072] = t[12071] ^ n[12072];
assign t[12073] = t[12072] ^ n[12073];
assign t[12074] = t[12073] ^ n[12074];
assign t[12075] = t[12074] ^ n[12075];
assign t[12076] = t[12075] ^ n[12076];
assign t[12077] = t[12076] ^ n[12077];
assign t[12078] = t[12077] ^ n[12078];
assign t[12079] = t[12078] ^ n[12079];
assign t[12080] = t[12079] ^ n[12080];
assign t[12081] = t[12080] ^ n[12081];
assign t[12082] = t[12081] ^ n[12082];
assign t[12083] = t[12082] ^ n[12083];
assign t[12084] = t[12083] ^ n[12084];
assign t[12085] = t[12084] ^ n[12085];
assign t[12086] = t[12085] ^ n[12086];
assign t[12087] = t[12086] ^ n[12087];
assign t[12088] = t[12087] ^ n[12088];
assign t[12089] = t[12088] ^ n[12089];
assign t[12090] = t[12089] ^ n[12090];
assign t[12091] = t[12090] ^ n[12091];
assign t[12092] = t[12091] ^ n[12092];
assign t[12093] = t[12092] ^ n[12093];
assign t[12094] = t[12093] ^ n[12094];
assign t[12095] = t[12094] ^ n[12095];
assign t[12096] = t[12095] ^ n[12096];
assign t[12097] = t[12096] ^ n[12097];
assign t[12098] = t[12097] ^ n[12098];
assign t[12099] = t[12098] ^ n[12099];
assign t[12100] = t[12099] ^ n[12100];
assign t[12101] = t[12100] ^ n[12101];
assign t[12102] = t[12101] ^ n[12102];
assign t[12103] = t[12102] ^ n[12103];
assign t[12104] = t[12103] ^ n[12104];
assign t[12105] = t[12104] ^ n[12105];
assign t[12106] = t[12105] ^ n[12106];
assign t[12107] = t[12106] ^ n[12107];
assign t[12108] = t[12107] ^ n[12108];
assign t[12109] = t[12108] ^ n[12109];
assign t[12110] = t[12109] ^ n[12110];
assign t[12111] = t[12110] ^ n[12111];
assign t[12112] = t[12111] ^ n[12112];
assign t[12113] = t[12112] ^ n[12113];
assign t[12114] = t[12113] ^ n[12114];
assign t[12115] = t[12114] ^ n[12115];
assign t[12116] = t[12115] ^ n[12116];
assign t[12117] = t[12116] ^ n[12117];
assign t[12118] = t[12117] ^ n[12118];
assign t[12119] = t[12118] ^ n[12119];
assign t[12120] = t[12119] ^ n[12120];
assign t[12121] = t[12120] ^ n[12121];
assign t[12122] = t[12121] ^ n[12122];
assign t[12123] = t[12122] ^ n[12123];
assign t[12124] = t[12123] ^ n[12124];
assign t[12125] = t[12124] ^ n[12125];
assign t[12126] = t[12125] ^ n[12126];
assign t[12127] = t[12126] ^ n[12127];
assign t[12128] = t[12127] ^ n[12128];
assign t[12129] = t[12128] ^ n[12129];
assign t[12130] = t[12129] ^ n[12130];
assign t[12131] = t[12130] ^ n[12131];
assign t[12132] = t[12131] ^ n[12132];
assign t[12133] = t[12132] ^ n[12133];
assign t[12134] = t[12133] ^ n[12134];
assign t[12135] = t[12134] ^ n[12135];
assign t[12136] = t[12135] ^ n[12136];
assign t[12137] = t[12136] ^ n[12137];
assign t[12138] = t[12137] ^ n[12138];
assign t[12139] = t[12138] ^ n[12139];
assign t[12140] = t[12139] ^ n[12140];
assign t[12141] = t[12140] ^ n[12141];
assign t[12142] = t[12141] ^ n[12142];
assign t[12143] = t[12142] ^ n[12143];
assign t[12144] = t[12143] ^ n[12144];
assign t[12145] = t[12144] ^ n[12145];
assign t[12146] = t[12145] ^ n[12146];
assign t[12147] = t[12146] ^ n[12147];
assign t[12148] = t[12147] ^ n[12148];
assign t[12149] = t[12148] ^ n[12149];
assign t[12150] = t[12149] ^ n[12150];
assign t[12151] = t[12150] ^ n[12151];
assign t[12152] = t[12151] ^ n[12152];
assign t[12153] = t[12152] ^ n[12153];
assign t[12154] = t[12153] ^ n[12154];
assign t[12155] = t[12154] ^ n[12155];
assign t[12156] = t[12155] ^ n[12156];
assign t[12157] = t[12156] ^ n[12157];
assign t[12158] = t[12157] ^ n[12158];
assign t[12159] = t[12158] ^ n[12159];
assign t[12160] = t[12159] ^ n[12160];
assign t[12161] = t[12160] ^ n[12161];
assign t[12162] = t[12161] ^ n[12162];
assign t[12163] = t[12162] ^ n[12163];
assign t[12164] = t[12163] ^ n[12164];
assign t[12165] = t[12164] ^ n[12165];
assign t[12166] = t[12165] ^ n[12166];
assign t[12167] = t[12166] ^ n[12167];
assign t[12168] = t[12167] ^ n[12168];
assign t[12169] = t[12168] ^ n[12169];
assign t[12170] = t[12169] ^ n[12170];
assign t[12171] = t[12170] ^ n[12171];
assign t[12172] = t[12171] ^ n[12172];
assign t[12173] = t[12172] ^ n[12173];
assign t[12174] = t[12173] ^ n[12174];
assign t[12175] = t[12174] ^ n[12175];
assign t[12176] = t[12175] ^ n[12176];
assign t[12177] = t[12176] ^ n[12177];
assign t[12178] = t[12177] ^ n[12178];
assign t[12179] = t[12178] ^ n[12179];
assign t[12180] = t[12179] ^ n[12180];
assign t[12181] = t[12180] ^ n[12181];
assign t[12182] = t[12181] ^ n[12182];
assign t[12183] = t[12182] ^ n[12183];
assign t[12184] = t[12183] ^ n[12184];
assign t[12185] = t[12184] ^ n[12185];
assign t[12186] = t[12185] ^ n[12186];
assign t[12187] = t[12186] ^ n[12187];
assign t[12188] = t[12187] ^ n[12188];
assign t[12189] = t[12188] ^ n[12189];
assign t[12190] = t[12189] ^ n[12190];
assign t[12191] = t[12190] ^ n[12191];
assign t[12192] = t[12191] ^ n[12192];
assign t[12193] = t[12192] ^ n[12193];
assign t[12194] = t[12193] ^ n[12194];
assign t[12195] = t[12194] ^ n[12195];
assign t[12196] = t[12195] ^ n[12196];
assign t[12197] = t[12196] ^ n[12197];
assign t[12198] = t[12197] ^ n[12198];
assign t[12199] = t[12198] ^ n[12199];
assign t[12200] = t[12199] ^ n[12200];
assign t[12201] = t[12200] ^ n[12201];
assign t[12202] = t[12201] ^ n[12202];
assign t[12203] = t[12202] ^ n[12203];
assign t[12204] = t[12203] ^ n[12204];
assign t[12205] = t[12204] ^ n[12205];
assign t[12206] = t[12205] ^ n[12206];
assign t[12207] = t[12206] ^ n[12207];
assign t[12208] = t[12207] ^ n[12208];
assign t[12209] = t[12208] ^ n[12209];
assign t[12210] = t[12209] ^ n[12210];
assign t[12211] = t[12210] ^ n[12211];
assign t[12212] = t[12211] ^ n[12212];
assign t[12213] = t[12212] ^ n[12213];
assign t[12214] = t[12213] ^ n[12214];
assign t[12215] = t[12214] ^ n[12215];
assign t[12216] = t[12215] ^ n[12216];
assign t[12217] = t[12216] ^ n[12217];
assign t[12218] = t[12217] ^ n[12218];
assign t[12219] = t[12218] ^ n[12219];
assign t[12220] = t[12219] ^ n[12220];
assign t[12221] = t[12220] ^ n[12221];
assign t[12222] = t[12221] ^ n[12222];
assign t[12223] = t[12222] ^ n[12223];
assign t[12224] = t[12223] ^ n[12224];
assign t[12225] = t[12224] ^ n[12225];
assign t[12226] = t[12225] ^ n[12226];
assign t[12227] = t[12226] ^ n[12227];
assign t[12228] = t[12227] ^ n[12228];
assign t[12229] = t[12228] ^ n[12229];
assign t[12230] = t[12229] ^ n[12230];
assign t[12231] = t[12230] ^ n[12231];
assign t[12232] = t[12231] ^ n[12232];
assign t[12233] = t[12232] ^ n[12233];
assign t[12234] = t[12233] ^ n[12234];
assign t[12235] = t[12234] ^ n[12235];
assign t[12236] = t[12235] ^ n[12236];
assign t[12237] = t[12236] ^ n[12237];
assign t[12238] = t[12237] ^ n[12238];
assign t[12239] = t[12238] ^ n[12239];
assign t[12240] = t[12239] ^ n[12240];
assign t[12241] = t[12240] ^ n[12241];
assign t[12242] = t[12241] ^ n[12242];
assign t[12243] = t[12242] ^ n[12243];
assign t[12244] = t[12243] ^ n[12244];
assign t[12245] = t[12244] ^ n[12245];
assign t[12246] = t[12245] ^ n[12246];
assign t[12247] = t[12246] ^ n[12247];
assign t[12248] = t[12247] ^ n[12248];
assign t[12249] = t[12248] ^ n[12249];
assign t[12250] = t[12249] ^ n[12250];
assign t[12251] = t[12250] ^ n[12251];
assign t[12252] = t[12251] ^ n[12252];
assign t[12253] = t[12252] ^ n[12253];
assign t[12254] = t[12253] ^ n[12254];
assign t[12255] = t[12254] ^ n[12255];
assign t[12256] = t[12255] ^ n[12256];
assign t[12257] = t[12256] ^ n[12257];
assign t[12258] = t[12257] ^ n[12258];
assign t[12259] = t[12258] ^ n[12259];
assign t[12260] = t[12259] ^ n[12260];
assign t[12261] = t[12260] ^ n[12261];
assign t[12262] = t[12261] ^ n[12262];
assign t[12263] = t[12262] ^ n[12263];
assign t[12264] = t[12263] ^ n[12264];
assign t[12265] = t[12264] ^ n[12265];
assign t[12266] = t[12265] ^ n[12266];
assign t[12267] = t[12266] ^ n[12267];
assign t[12268] = t[12267] ^ n[12268];
assign t[12269] = t[12268] ^ n[12269];
assign t[12270] = t[12269] ^ n[12270];
assign t[12271] = t[12270] ^ n[12271];
assign t[12272] = t[12271] ^ n[12272];
assign t[12273] = t[12272] ^ n[12273];
assign t[12274] = t[12273] ^ n[12274];
assign t[12275] = t[12274] ^ n[12275];
assign t[12276] = t[12275] ^ n[12276];
assign t[12277] = t[12276] ^ n[12277];
assign t[12278] = t[12277] ^ n[12278];
assign t[12279] = t[12278] ^ n[12279];
assign t[12280] = t[12279] ^ n[12280];
assign t[12281] = t[12280] ^ n[12281];
assign t[12282] = t[12281] ^ n[12282];
assign t[12283] = t[12282] ^ n[12283];
assign t[12284] = t[12283] ^ n[12284];
assign t[12285] = t[12284] ^ n[12285];
assign t[12286] = t[12285] ^ n[12286];
assign t[12287] = t[12286] ^ n[12287];
assign t[12288] = t[12287] ^ n[12288];
assign t[12289] = t[12288] ^ n[12289];
assign t[12290] = t[12289] ^ n[12290];
assign t[12291] = t[12290] ^ n[12291];
assign t[12292] = t[12291] ^ n[12292];
assign t[12293] = t[12292] ^ n[12293];
assign t[12294] = t[12293] ^ n[12294];
assign t[12295] = t[12294] ^ n[12295];
assign t[12296] = t[12295] ^ n[12296];
assign t[12297] = t[12296] ^ n[12297];
assign t[12298] = t[12297] ^ n[12298];
assign t[12299] = t[12298] ^ n[12299];
assign t[12300] = t[12299] ^ n[12300];
assign t[12301] = t[12300] ^ n[12301];
assign t[12302] = t[12301] ^ n[12302];
assign t[12303] = t[12302] ^ n[12303];
assign t[12304] = t[12303] ^ n[12304];
assign t[12305] = t[12304] ^ n[12305];
assign t[12306] = t[12305] ^ n[12306];
assign t[12307] = t[12306] ^ n[12307];
assign t[12308] = t[12307] ^ n[12308];
assign t[12309] = t[12308] ^ n[12309];
assign t[12310] = t[12309] ^ n[12310];
assign t[12311] = t[12310] ^ n[12311];
assign t[12312] = t[12311] ^ n[12312];
assign t[12313] = t[12312] ^ n[12313];
assign t[12314] = t[12313] ^ n[12314];
assign t[12315] = t[12314] ^ n[12315];
assign t[12316] = t[12315] ^ n[12316];
assign t[12317] = t[12316] ^ n[12317];
assign t[12318] = t[12317] ^ n[12318];
assign t[12319] = t[12318] ^ n[12319];
assign t[12320] = t[12319] ^ n[12320];
assign t[12321] = t[12320] ^ n[12321];
assign t[12322] = t[12321] ^ n[12322];
assign t[12323] = t[12322] ^ n[12323];
assign t[12324] = t[12323] ^ n[12324];
assign t[12325] = t[12324] ^ n[12325];
assign t[12326] = t[12325] ^ n[12326];
assign t[12327] = t[12326] ^ n[12327];
assign t[12328] = t[12327] ^ n[12328];
assign t[12329] = t[12328] ^ n[12329];
assign t[12330] = t[12329] ^ n[12330];
assign t[12331] = t[12330] ^ n[12331];
assign t[12332] = t[12331] ^ n[12332];
assign t[12333] = t[12332] ^ n[12333];
assign t[12334] = t[12333] ^ n[12334];
assign t[12335] = t[12334] ^ n[12335];
assign t[12336] = t[12335] ^ n[12336];
assign t[12337] = t[12336] ^ n[12337];
assign t[12338] = t[12337] ^ n[12338];
assign t[12339] = t[12338] ^ n[12339];
assign t[12340] = t[12339] ^ n[12340];
assign t[12341] = t[12340] ^ n[12341];
assign t[12342] = t[12341] ^ n[12342];
assign t[12343] = t[12342] ^ n[12343];
assign t[12344] = t[12343] ^ n[12344];
assign t[12345] = t[12344] ^ n[12345];
assign t[12346] = t[12345] ^ n[12346];
assign t[12347] = t[12346] ^ n[12347];
assign t[12348] = t[12347] ^ n[12348];
assign t[12349] = t[12348] ^ n[12349];
assign t[12350] = t[12349] ^ n[12350];
assign t[12351] = t[12350] ^ n[12351];
assign t[12352] = t[12351] ^ n[12352];
assign t[12353] = t[12352] ^ n[12353];
assign t[12354] = t[12353] ^ n[12354];
assign t[12355] = t[12354] ^ n[12355];
assign t[12356] = t[12355] ^ n[12356];
assign t[12357] = t[12356] ^ n[12357];
assign t[12358] = t[12357] ^ n[12358];
assign t[12359] = t[12358] ^ n[12359];
assign t[12360] = t[12359] ^ n[12360];
assign t[12361] = t[12360] ^ n[12361];
assign t[12362] = t[12361] ^ n[12362];
assign t[12363] = t[12362] ^ n[12363];
assign t[12364] = t[12363] ^ n[12364];
assign t[12365] = t[12364] ^ n[12365];
assign t[12366] = t[12365] ^ n[12366];
assign t[12367] = t[12366] ^ n[12367];
assign t[12368] = t[12367] ^ n[12368];
assign t[12369] = t[12368] ^ n[12369];
assign t[12370] = t[12369] ^ n[12370];
assign t[12371] = t[12370] ^ n[12371];
assign t[12372] = t[12371] ^ n[12372];
assign t[12373] = t[12372] ^ n[12373];
assign t[12374] = t[12373] ^ n[12374];
assign t[12375] = t[12374] ^ n[12375];
assign t[12376] = t[12375] ^ n[12376];
assign t[12377] = t[12376] ^ n[12377];
assign t[12378] = t[12377] ^ n[12378];
assign t[12379] = t[12378] ^ n[12379];
assign t[12380] = t[12379] ^ n[12380];
assign t[12381] = t[12380] ^ n[12381];
assign t[12382] = t[12381] ^ n[12382];
assign t[12383] = t[12382] ^ n[12383];
assign t[12384] = t[12383] ^ n[12384];
assign t[12385] = t[12384] ^ n[12385];
assign t[12386] = t[12385] ^ n[12386];
assign t[12387] = t[12386] ^ n[12387];
assign t[12388] = t[12387] ^ n[12388];
assign t[12389] = t[12388] ^ n[12389];
assign t[12390] = t[12389] ^ n[12390];
assign t[12391] = t[12390] ^ n[12391];
assign t[12392] = t[12391] ^ n[12392];
assign t[12393] = t[12392] ^ n[12393];
assign t[12394] = t[12393] ^ n[12394];
assign t[12395] = t[12394] ^ n[12395];
assign t[12396] = t[12395] ^ n[12396];
assign t[12397] = t[12396] ^ n[12397];
assign t[12398] = t[12397] ^ n[12398];
assign t[12399] = t[12398] ^ n[12399];
assign t[12400] = t[12399] ^ n[12400];
assign t[12401] = t[12400] ^ n[12401];
assign t[12402] = t[12401] ^ n[12402];
assign t[12403] = t[12402] ^ n[12403];
assign t[12404] = t[12403] ^ n[12404];
assign t[12405] = t[12404] ^ n[12405];
assign t[12406] = t[12405] ^ n[12406];
assign t[12407] = t[12406] ^ n[12407];
assign t[12408] = t[12407] ^ n[12408];
assign t[12409] = t[12408] ^ n[12409];
assign t[12410] = t[12409] ^ n[12410];
assign t[12411] = t[12410] ^ n[12411];
assign t[12412] = t[12411] ^ n[12412];
assign t[12413] = t[12412] ^ n[12413];
assign t[12414] = t[12413] ^ n[12414];
assign t[12415] = t[12414] ^ n[12415];
assign t[12416] = t[12415] ^ n[12416];
assign t[12417] = t[12416] ^ n[12417];
assign t[12418] = t[12417] ^ n[12418];
assign t[12419] = t[12418] ^ n[12419];
assign t[12420] = t[12419] ^ n[12420];
assign t[12421] = t[12420] ^ n[12421];
assign t[12422] = t[12421] ^ n[12422];
assign t[12423] = t[12422] ^ n[12423];
assign t[12424] = t[12423] ^ n[12424];
assign t[12425] = t[12424] ^ n[12425];
assign t[12426] = t[12425] ^ n[12426];
assign t[12427] = t[12426] ^ n[12427];
assign t[12428] = t[12427] ^ n[12428];
assign t[12429] = t[12428] ^ n[12429];
assign t[12430] = t[12429] ^ n[12430];
assign t[12431] = t[12430] ^ n[12431];
assign t[12432] = t[12431] ^ n[12432];
assign t[12433] = t[12432] ^ n[12433];
assign t[12434] = t[12433] ^ n[12434];
assign t[12435] = t[12434] ^ n[12435];
assign t[12436] = t[12435] ^ n[12436];
assign t[12437] = t[12436] ^ n[12437];
assign t[12438] = t[12437] ^ n[12438];
assign t[12439] = t[12438] ^ n[12439];
assign t[12440] = t[12439] ^ n[12440];
assign t[12441] = t[12440] ^ n[12441];
assign t[12442] = t[12441] ^ n[12442];
assign t[12443] = t[12442] ^ n[12443];
assign t[12444] = t[12443] ^ n[12444];
assign t[12445] = t[12444] ^ n[12445];
assign t[12446] = t[12445] ^ n[12446];
assign t[12447] = t[12446] ^ n[12447];
assign t[12448] = t[12447] ^ n[12448];
assign t[12449] = t[12448] ^ n[12449];
assign t[12450] = t[12449] ^ n[12450];
assign t[12451] = t[12450] ^ n[12451];
assign t[12452] = t[12451] ^ n[12452];
assign t[12453] = t[12452] ^ n[12453];
assign t[12454] = t[12453] ^ n[12454];
assign t[12455] = t[12454] ^ n[12455];
assign t[12456] = t[12455] ^ n[12456];
assign t[12457] = t[12456] ^ n[12457];
assign t[12458] = t[12457] ^ n[12458];
assign t[12459] = t[12458] ^ n[12459];
assign t[12460] = t[12459] ^ n[12460];
assign t[12461] = t[12460] ^ n[12461];
assign t[12462] = t[12461] ^ n[12462];
assign t[12463] = t[12462] ^ n[12463];
assign t[12464] = t[12463] ^ n[12464];
assign t[12465] = t[12464] ^ n[12465];
assign t[12466] = t[12465] ^ n[12466];
assign t[12467] = t[12466] ^ n[12467];
assign t[12468] = t[12467] ^ n[12468];
assign t[12469] = t[12468] ^ n[12469];
assign t[12470] = t[12469] ^ n[12470];
assign t[12471] = t[12470] ^ n[12471];
assign t[12472] = t[12471] ^ n[12472];
assign t[12473] = t[12472] ^ n[12473];
assign t[12474] = t[12473] ^ n[12474];
assign t[12475] = t[12474] ^ n[12475];
assign t[12476] = t[12475] ^ n[12476];
assign t[12477] = t[12476] ^ n[12477];
assign t[12478] = t[12477] ^ n[12478];
assign t[12479] = t[12478] ^ n[12479];
assign t[12480] = t[12479] ^ n[12480];
assign t[12481] = t[12480] ^ n[12481];
assign t[12482] = t[12481] ^ n[12482];
assign t[12483] = t[12482] ^ n[12483];
assign t[12484] = t[12483] ^ n[12484];
assign t[12485] = t[12484] ^ n[12485];
assign t[12486] = t[12485] ^ n[12486];
assign t[12487] = t[12486] ^ n[12487];
assign t[12488] = t[12487] ^ n[12488];
assign t[12489] = t[12488] ^ n[12489];
assign t[12490] = t[12489] ^ n[12490];
assign t[12491] = t[12490] ^ n[12491];
assign t[12492] = t[12491] ^ n[12492];
assign t[12493] = t[12492] ^ n[12493];
assign t[12494] = t[12493] ^ n[12494];
assign t[12495] = t[12494] ^ n[12495];
assign t[12496] = t[12495] ^ n[12496];
assign t[12497] = t[12496] ^ n[12497];
assign t[12498] = t[12497] ^ n[12498];
assign t[12499] = t[12498] ^ n[12499];
assign t[12500] = t[12499] ^ n[12500];
assign t[12501] = t[12500] ^ n[12501];
assign t[12502] = t[12501] ^ n[12502];
assign t[12503] = t[12502] ^ n[12503];
assign t[12504] = t[12503] ^ n[12504];
assign t[12505] = t[12504] ^ n[12505];
assign t[12506] = t[12505] ^ n[12506];
assign t[12507] = t[12506] ^ n[12507];
assign t[12508] = t[12507] ^ n[12508];
assign t[12509] = t[12508] ^ n[12509];
assign t[12510] = t[12509] ^ n[12510];
assign t[12511] = t[12510] ^ n[12511];
assign t[12512] = t[12511] ^ n[12512];
assign t[12513] = t[12512] ^ n[12513];
assign t[12514] = t[12513] ^ n[12514];
assign t[12515] = t[12514] ^ n[12515];
assign t[12516] = t[12515] ^ n[12516];
assign t[12517] = t[12516] ^ n[12517];
assign t[12518] = t[12517] ^ n[12518];
assign t[12519] = t[12518] ^ n[12519];
assign t[12520] = t[12519] ^ n[12520];
assign t[12521] = t[12520] ^ n[12521];
assign t[12522] = t[12521] ^ n[12522];
assign t[12523] = t[12522] ^ n[12523];
assign t[12524] = t[12523] ^ n[12524];
assign t[12525] = t[12524] ^ n[12525];
assign t[12526] = t[12525] ^ n[12526];
assign t[12527] = t[12526] ^ n[12527];
assign t[12528] = t[12527] ^ n[12528];
assign t[12529] = t[12528] ^ n[12529];
assign t[12530] = t[12529] ^ n[12530];
assign t[12531] = t[12530] ^ n[12531];
assign t[12532] = t[12531] ^ n[12532];
assign t[12533] = t[12532] ^ n[12533];
assign t[12534] = t[12533] ^ n[12534];
assign t[12535] = t[12534] ^ n[12535];
assign t[12536] = t[12535] ^ n[12536];
assign t[12537] = t[12536] ^ n[12537];
assign t[12538] = t[12537] ^ n[12538];
assign t[12539] = t[12538] ^ n[12539];
assign t[12540] = t[12539] ^ n[12540];
assign t[12541] = t[12540] ^ n[12541];
assign t[12542] = t[12541] ^ n[12542];
assign t[12543] = t[12542] ^ n[12543];
assign t[12544] = t[12543] ^ n[12544];
assign t[12545] = t[12544] ^ n[12545];
assign t[12546] = t[12545] ^ n[12546];
assign t[12547] = t[12546] ^ n[12547];
assign t[12548] = t[12547] ^ n[12548];
assign t[12549] = t[12548] ^ n[12549];
assign t[12550] = t[12549] ^ n[12550];
assign t[12551] = t[12550] ^ n[12551];
assign t[12552] = t[12551] ^ n[12552];
assign t[12553] = t[12552] ^ n[12553];
assign t[12554] = t[12553] ^ n[12554];
assign t[12555] = t[12554] ^ n[12555];
assign t[12556] = t[12555] ^ n[12556];
assign t[12557] = t[12556] ^ n[12557];
assign t[12558] = t[12557] ^ n[12558];
assign t[12559] = t[12558] ^ n[12559];
assign t[12560] = t[12559] ^ n[12560];
assign t[12561] = t[12560] ^ n[12561];
assign t[12562] = t[12561] ^ n[12562];
assign t[12563] = t[12562] ^ n[12563];
assign t[12564] = t[12563] ^ n[12564];
assign t[12565] = t[12564] ^ n[12565];
assign t[12566] = t[12565] ^ n[12566];
assign t[12567] = t[12566] ^ n[12567];
assign t[12568] = t[12567] ^ n[12568];
assign t[12569] = t[12568] ^ n[12569];
assign t[12570] = t[12569] ^ n[12570];
assign t[12571] = t[12570] ^ n[12571];
assign t[12572] = t[12571] ^ n[12572];
assign t[12573] = t[12572] ^ n[12573];
assign t[12574] = t[12573] ^ n[12574];
assign t[12575] = t[12574] ^ n[12575];
assign t[12576] = t[12575] ^ n[12576];
assign t[12577] = t[12576] ^ n[12577];
assign t[12578] = t[12577] ^ n[12578];
assign t[12579] = t[12578] ^ n[12579];
assign t[12580] = t[12579] ^ n[12580];
assign t[12581] = t[12580] ^ n[12581];
assign t[12582] = t[12581] ^ n[12582];
assign t[12583] = t[12582] ^ n[12583];
assign t[12584] = t[12583] ^ n[12584];
assign t[12585] = t[12584] ^ n[12585];
assign t[12586] = t[12585] ^ n[12586];
assign t[12587] = t[12586] ^ n[12587];
assign t[12588] = t[12587] ^ n[12588];
assign t[12589] = t[12588] ^ n[12589];
assign t[12590] = t[12589] ^ n[12590];
assign t[12591] = t[12590] ^ n[12591];
assign t[12592] = t[12591] ^ n[12592];
assign t[12593] = t[12592] ^ n[12593];
assign t[12594] = t[12593] ^ n[12594];
assign t[12595] = t[12594] ^ n[12595];
assign t[12596] = t[12595] ^ n[12596];
assign t[12597] = t[12596] ^ n[12597];
assign t[12598] = t[12597] ^ n[12598];
assign t[12599] = t[12598] ^ n[12599];
assign t[12600] = t[12599] ^ n[12600];
assign t[12601] = t[12600] ^ n[12601];
assign t[12602] = t[12601] ^ n[12602];
assign t[12603] = t[12602] ^ n[12603];
assign t[12604] = t[12603] ^ n[12604];
assign t[12605] = t[12604] ^ n[12605];
assign t[12606] = t[12605] ^ n[12606];
assign t[12607] = t[12606] ^ n[12607];
assign t[12608] = t[12607] ^ n[12608];
assign t[12609] = t[12608] ^ n[12609];
assign t[12610] = t[12609] ^ n[12610];
assign t[12611] = t[12610] ^ n[12611];
assign t[12612] = t[12611] ^ n[12612];
assign t[12613] = t[12612] ^ n[12613];
assign t[12614] = t[12613] ^ n[12614];
assign t[12615] = t[12614] ^ n[12615];
assign t[12616] = t[12615] ^ n[12616];
assign t[12617] = t[12616] ^ n[12617];
assign t[12618] = t[12617] ^ n[12618];
assign t[12619] = t[12618] ^ n[12619];
assign t[12620] = t[12619] ^ n[12620];
assign t[12621] = t[12620] ^ n[12621];
assign t[12622] = t[12621] ^ n[12622];
assign t[12623] = t[12622] ^ n[12623];
assign t[12624] = t[12623] ^ n[12624];
assign t[12625] = t[12624] ^ n[12625];
assign t[12626] = t[12625] ^ n[12626];
assign t[12627] = t[12626] ^ n[12627];
assign t[12628] = t[12627] ^ n[12628];
assign t[12629] = t[12628] ^ n[12629];
assign t[12630] = t[12629] ^ n[12630];
assign t[12631] = t[12630] ^ n[12631];
assign t[12632] = t[12631] ^ n[12632];
assign t[12633] = t[12632] ^ n[12633];
assign t[12634] = t[12633] ^ n[12634];
assign t[12635] = t[12634] ^ n[12635];
assign t[12636] = t[12635] ^ n[12636];
assign t[12637] = t[12636] ^ n[12637];
assign t[12638] = t[12637] ^ n[12638];
assign t[12639] = t[12638] ^ n[12639];
assign t[12640] = t[12639] ^ n[12640];
assign t[12641] = t[12640] ^ n[12641];
assign t[12642] = t[12641] ^ n[12642];
assign t[12643] = t[12642] ^ n[12643];
assign t[12644] = t[12643] ^ n[12644];
assign t[12645] = t[12644] ^ n[12645];
assign t[12646] = t[12645] ^ n[12646];
assign t[12647] = t[12646] ^ n[12647];
assign t[12648] = t[12647] ^ n[12648];
assign t[12649] = t[12648] ^ n[12649];
assign t[12650] = t[12649] ^ n[12650];
assign t[12651] = t[12650] ^ n[12651];
assign t[12652] = t[12651] ^ n[12652];
assign t[12653] = t[12652] ^ n[12653];
assign t[12654] = t[12653] ^ n[12654];
assign t[12655] = t[12654] ^ n[12655];
assign t[12656] = t[12655] ^ n[12656];
assign t[12657] = t[12656] ^ n[12657];
assign t[12658] = t[12657] ^ n[12658];
assign t[12659] = t[12658] ^ n[12659];
assign t[12660] = t[12659] ^ n[12660];
assign t[12661] = t[12660] ^ n[12661];
assign t[12662] = t[12661] ^ n[12662];
assign t[12663] = t[12662] ^ n[12663];
assign t[12664] = t[12663] ^ n[12664];
assign t[12665] = t[12664] ^ n[12665];
assign t[12666] = t[12665] ^ n[12666];
assign t[12667] = t[12666] ^ n[12667];
assign t[12668] = t[12667] ^ n[12668];
assign t[12669] = t[12668] ^ n[12669];
assign t[12670] = t[12669] ^ n[12670];
assign t[12671] = t[12670] ^ n[12671];
assign t[12672] = t[12671] ^ n[12672];
assign t[12673] = t[12672] ^ n[12673];
assign t[12674] = t[12673] ^ n[12674];
assign t[12675] = t[12674] ^ n[12675];
assign t[12676] = t[12675] ^ n[12676];
assign t[12677] = t[12676] ^ n[12677];
assign t[12678] = t[12677] ^ n[12678];
assign t[12679] = t[12678] ^ n[12679];
assign t[12680] = t[12679] ^ n[12680];
assign t[12681] = t[12680] ^ n[12681];
assign t[12682] = t[12681] ^ n[12682];
assign t[12683] = t[12682] ^ n[12683];
assign t[12684] = t[12683] ^ n[12684];
assign t[12685] = t[12684] ^ n[12685];
assign t[12686] = t[12685] ^ n[12686];
assign t[12687] = t[12686] ^ n[12687];
assign t[12688] = t[12687] ^ n[12688];
assign t[12689] = t[12688] ^ n[12689];
assign t[12690] = t[12689] ^ n[12690];
assign t[12691] = t[12690] ^ n[12691];
assign t[12692] = t[12691] ^ n[12692];
assign t[12693] = t[12692] ^ n[12693];
assign t[12694] = t[12693] ^ n[12694];
assign t[12695] = t[12694] ^ n[12695];
assign t[12696] = t[12695] ^ n[12696];
assign t[12697] = t[12696] ^ n[12697];
assign t[12698] = t[12697] ^ n[12698];
assign t[12699] = t[12698] ^ n[12699];
assign t[12700] = t[12699] ^ n[12700];
assign t[12701] = t[12700] ^ n[12701];
assign t[12702] = t[12701] ^ n[12702];
assign t[12703] = t[12702] ^ n[12703];
assign t[12704] = t[12703] ^ n[12704];
assign t[12705] = t[12704] ^ n[12705];
assign t[12706] = t[12705] ^ n[12706];
assign t[12707] = t[12706] ^ n[12707];
assign t[12708] = t[12707] ^ n[12708];
assign t[12709] = t[12708] ^ n[12709];
assign t[12710] = t[12709] ^ n[12710];
assign t[12711] = t[12710] ^ n[12711];
assign t[12712] = t[12711] ^ n[12712];
assign t[12713] = t[12712] ^ n[12713];
assign t[12714] = t[12713] ^ n[12714];
assign t[12715] = t[12714] ^ n[12715];
assign t[12716] = t[12715] ^ n[12716];
assign t[12717] = t[12716] ^ n[12717];
assign t[12718] = t[12717] ^ n[12718];
assign t[12719] = t[12718] ^ n[12719];
assign t[12720] = t[12719] ^ n[12720];
assign t[12721] = t[12720] ^ n[12721];
assign t[12722] = t[12721] ^ n[12722];
assign t[12723] = t[12722] ^ n[12723];
assign t[12724] = t[12723] ^ n[12724];
assign t[12725] = t[12724] ^ n[12725];
assign t[12726] = t[12725] ^ n[12726];
assign t[12727] = t[12726] ^ n[12727];
assign t[12728] = t[12727] ^ n[12728];
assign t[12729] = t[12728] ^ n[12729];
assign t[12730] = t[12729] ^ n[12730];
assign t[12731] = t[12730] ^ n[12731];
assign t[12732] = t[12731] ^ n[12732];
assign t[12733] = t[12732] ^ n[12733];
assign t[12734] = t[12733] ^ n[12734];
assign t[12735] = t[12734] ^ n[12735];
assign t[12736] = t[12735] ^ n[12736];
assign t[12737] = t[12736] ^ n[12737];
assign t[12738] = t[12737] ^ n[12738];
assign t[12739] = t[12738] ^ n[12739];
assign t[12740] = t[12739] ^ n[12740];
assign t[12741] = t[12740] ^ n[12741];
assign t[12742] = t[12741] ^ n[12742];
assign t[12743] = t[12742] ^ n[12743];
assign t[12744] = t[12743] ^ n[12744];
assign t[12745] = t[12744] ^ n[12745];
assign t[12746] = t[12745] ^ n[12746];
assign t[12747] = t[12746] ^ n[12747];
assign t[12748] = t[12747] ^ n[12748];
assign t[12749] = t[12748] ^ n[12749];
assign t[12750] = t[12749] ^ n[12750];
assign t[12751] = t[12750] ^ n[12751];
assign t[12752] = t[12751] ^ n[12752];
assign t[12753] = t[12752] ^ n[12753];
assign t[12754] = t[12753] ^ n[12754];
assign t[12755] = t[12754] ^ n[12755];
assign t[12756] = t[12755] ^ n[12756];
assign t[12757] = t[12756] ^ n[12757];
assign t[12758] = t[12757] ^ n[12758];
assign t[12759] = t[12758] ^ n[12759];
assign t[12760] = t[12759] ^ n[12760];
assign t[12761] = t[12760] ^ n[12761];
assign t[12762] = t[12761] ^ n[12762];
assign t[12763] = t[12762] ^ n[12763];
assign t[12764] = t[12763] ^ n[12764];
assign t[12765] = t[12764] ^ n[12765];
assign t[12766] = t[12765] ^ n[12766];
assign t[12767] = t[12766] ^ n[12767];
assign t[12768] = t[12767] ^ n[12768];
assign t[12769] = t[12768] ^ n[12769];
assign t[12770] = t[12769] ^ n[12770];
assign t[12771] = t[12770] ^ n[12771];
assign t[12772] = t[12771] ^ n[12772];
assign t[12773] = t[12772] ^ n[12773];
assign t[12774] = t[12773] ^ n[12774];
assign t[12775] = t[12774] ^ n[12775];
assign t[12776] = t[12775] ^ n[12776];
assign t[12777] = t[12776] ^ n[12777];
assign t[12778] = t[12777] ^ n[12778];
assign t[12779] = t[12778] ^ n[12779];
assign t[12780] = t[12779] ^ n[12780];
assign t[12781] = t[12780] ^ n[12781];
assign t[12782] = t[12781] ^ n[12782];
assign t[12783] = t[12782] ^ n[12783];
assign t[12784] = t[12783] ^ n[12784];
assign t[12785] = t[12784] ^ n[12785];
assign t[12786] = t[12785] ^ n[12786];
assign t[12787] = t[12786] ^ n[12787];
assign t[12788] = t[12787] ^ n[12788];
assign t[12789] = t[12788] ^ n[12789];
assign t[12790] = t[12789] ^ n[12790];
assign t[12791] = t[12790] ^ n[12791];
assign t[12792] = t[12791] ^ n[12792];
assign t[12793] = t[12792] ^ n[12793];
assign t[12794] = t[12793] ^ n[12794];
assign t[12795] = t[12794] ^ n[12795];
assign t[12796] = t[12795] ^ n[12796];
assign t[12797] = t[12796] ^ n[12797];
assign t[12798] = t[12797] ^ n[12798];
assign t[12799] = t[12798] ^ n[12799];
assign t[12800] = t[12799] ^ n[12800];
assign t[12801] = t[12800] ^ n[12801];
assign t[12802] = t[12801] ^ n[12802];
assign t[12803] = t[12802] ^ n[12803];
assign t[12804] = t[12803] ^ n[12804];
assign t[12805] = t[12804] ^ n[12805];
assign t[12806] = t[12805] ^ n[12806];
assign t[12807] = t[12806] ^ n[12807];
assign t[12808] = t[12807] ^ n[12808];
assign t[12809] = t[12808] ^ n[12809];
assign t[12810] = t[12809] ^ n[12810];
assign t[12811] = t[12810] ^ n[12811];
assign t[12812] = t[12811] ^ n[12812];
assign t[12813] = t[12812] ^ n[12813];
assign t[12814] = t[12813] ^ n[12814];
assign t[12815] = t[12814] ^ n[12815];
assign t[12816] = t[12815] ^ n[12816];
assign t[12817] = t[12816] ^ n[12817];
assign t[12818] = t[12817] ^ n[12818];
assign t[12819] = t[12818] ^ n[12819];
assign t[12820] = t[12819] ^ n[12820];
assign t[12821] = t[12820] ^ n[12821];
assign t[12822] = t[12821] ^ n[12822];
assign t[12823] = t[12822] ^ n[12823];
assign t[12824] = t[12823] ^ n[12824];
assign t[12825] = t[12824] ^ n[12825];
assign t[12826] = t[12825] ^ n[12826];
assign t[12827] = t[12826] ^ n[12827];
assign t[12828] = t[12827] ^ n[12828];
assign t[12829] = t[12828] ^ n[12829];
assign t[12830] = t[12829] ^ n[12830];
assign t[12831] = t[12830] ^ n[12831];
assign t[12832] = t[12831] ^ n[12832];
assign t[12833] = t[12832] ^ n[12833];
assign t[12834] = t[12833] ^ n[12834];
assign t[12835] = t[12834] ^ n[12835];
assign t[12836] = t[12835] ^ n[12836];
assign t[12837] = t[12836] ^ n[12837];
assign t[12838] = t[12837] ^ n[12838];
assign t[12839] = t[12838] ^ n[12839];
assign t[12840] = t[12839] ^ n[12840];
assign t[12841] = t[12840] ^ n[12841];
assign t[12842] = t[12841] ^ n[12842];
assign t[12843] = t[12842] ^ n[12843];
assign t[12844] = t[12843] ^ n[12844];
assign t[12845] = t[12844] ^ n[12845];
assign t[12846] = t[12845] ^ n[12846];
assign t[12847] = t[12846] ^ n[12847];
assign t[12848] = t[12847] ^ n[12848];
assign t[12849] = t[12848] ^ n[12849];
assign t[12850] = t[12849] ^ n[12850];
assign t[12851] = t[12850] ^ n[12851];
assign t[12852] = t[12851] ^ n[12852];
assign t[12853] = t[12852] ^ n[12853];
assign t[12854] = t[12853] ^ n[12854];
assign t[12855] = t[12854] ^ n[12855];
assign t[12856] = t[12855] ^ n[12856];
assign t[12857] = t[12856] ^ n[12857];
assign t[12858] = t[12857] ^ n[12858];
assign t[12859] = t[12858] ^ n[12859];
assign t[12860] = t[12859] ^ n[12860];
assign t[12861] = t[12860] ^ n[12861];
assign t[12862] = t[12861] ^ n[12862];
assign t[12863] = t[12862] ^ n[12863];
assign t[12864] = t[12863] ^ n[12864];
assign t[12865] = t[12864] ^ n[12865];
assign t[12866] = t[12865] ^ n[12866];
assign t[12867] = t[12866] ^ n[12867];
assign t[12868] = t[12867] ^ n[12868];
assign t[12869] = t[12868] ^ n[12869];
assign t[12870] = t[12869] ^ n[12870];
assign t[12871] = t[12870] ^ n[12871];
assign t[12872] = t[12871] ^ n[12872];
assign t[12873] = t[12872] ^ n[12873];
assign t[12874] = t[12873] ^ n[12874];
assign t[12875] = t[12874] ^ n[12875];
assign t[12876] = t[12875] ^ n[12876];
assign t[12877] = t[12876] ^ n[12877];
assign t[12878] = t[12877] ^ n[12878];
assign t[12879] = t[12878] ^ n[12879];
assign t[12880] = t[12879] ^ n[12880];
assign t[12881] = t[12880] ^ n[12881];
assign t[12882] = t[12881] ^ n[12882];
assign t[12883] = t[12882] ^ n[12883];
assign t[12884] = t[12883] ^ n[12884];
assign t[12885] = t[12884] ^ n[12885];
assign t[12886] = t[12885] ^ n[12886];
assign t[12887] = t[12886] ^ n[12887];
assign t[12888] = t[12887] ^ n[12888];
assign t[12889] = t[12888] ^ n[12889];
assign t[12890] = t[12889] ^ n[12890];
assign t[12891] = t[12890] ^ n[12891];
assign t[12892] = t[12891] ^ n[12892];
assign t[12893] = t[12892] ^ n[12893];
assign t[12894] = t[12893] ^ n[12894];
assign t[12895] = t[12894] ^ n[12895];
assign t[12896] = t[12895] ^ n[12896];
assign t[12897] = t[12896] ^ n[12897];
assign t[12898] = t[12897] ^ n[12898];
assign t[12899] = t[12898] ^ n[12899];
assign t[12900] = t[12899] ^ n[12900];
assign t[12901] = t[12900] ^ n[12901];
assign t[12902] = t[12901] ^ n[12902];
assign t[12903] = t[12902] ^ n[12903];
assign t[12904] = t[12903] ^ n[12904];
assign t[12905] = t[12904] ^ n[12905];
assign t[12906] = t[12905] ^ n[12906];
assign t[12907] = t[12906] ^ n[12907];
assign t[12908] = t[12907] ^ n[12908];
assign t[12909] = t[12908] ^ n[12909];
assign t[12910] = t[12909] ^ n[12910];
assign t[12911] = t[12910] ^ n[12911];
assign t[12912] = t[12911] ^ n[12912];
assign t[12913] = t[12912] ^ n[12913];
assign t[12914] = t[12913] ^ n[12914];
assign t[12915] = t[12914] ^ n[12915];
assign t[12916] = t[12915] ^ n[12916];
assign t[12917] = t[12916] ^ n[12917];
assign t[12918] = t[12917] ^ n[12918];
assign t[12919] = t[12918] ^ n[12919];
assign t[12920] = t[12919] ^ n[12920];
assign t[12921] = t[12920] ^ n[12921];
assign t[12922] = t[12921] ^ n[12922];
assign t[12923] = t[12922] ^ n[12923];
assign t[12924] = t[12923] ^ n[12924];
assign t[12925] = t[12924] ^ n[12925];
assign t[12926] = t[12925] ^ n[12926];
assign t[12927] = t[12926] ^ n[12927];
assign t[12928] = t[12927] ^ n[12928];
assign t[12929] = t[12928] ^ n[12929];
assign t[12930] = t[12929] ^ n[12930];
assign t[12931] = t[12930] ^ n[12931];
assign t[12932] = t[12931] ^ n[12932];
assign t[12933] = t[12932] ^ n[12933];
assign t[12934] = t[12933] ^ n[12934];
assign t[12935] = t[12934] ^ n[12935];
assign t[12936] = t[12935] ^ n[12936];
assign t[12937] = t[12936] ^ n[12937];
assign t[12938] = t[12937] ^ n[12938];
assign t[12939] = t[12938] ^ n[12939];
assign t[12940] = t[12939] ^ n[12940];
assign t[12941] = t[12940] ^ n[12941];
assign t[12942] = t[12941] ^ n[12942];
assign t[12943] = t[12942] ^ n[12943];
assign t[12944] = t[12943] ^ n[12944];
assign t[12945] = t[12944] ^ n[12945];
assign t[12946] = t[12945] ^ n[12946];
assign t[12947] = t[12946] ^ n[12947];
assign t[12948] = t[12947] ^ n[12948];
assign t[12949] = t[12948] ^ n[12949];
assign t[12950] = t[12949] ^ n[12950];
assign t[12951] = t[12950] ^ n[12951];
assign t[12952] = t[12951] ^ n[12952];
assign t[12953] = t[12952] ^ n[12953];
assign t[12954] = t[12953] ^ n[12954];
assign t[12955] = t[12954] ^ n[12955];
assign t[12956] = t[12955] ^ n[12956];
assign t[12957] = t[12956] ^ n[12957];
assign t[12958] = t[12957] ^ n[12958];
assign t[12959] = t[12958] ^ n[12959];
assign t[12960] = t[12959] ^ n[12960];
assign t[12961] = t[12960] ^ n[12961];
assign t[12962] = t[12961] ^ n[12962];
assign t[12963] = t[12962] ^ n[12963];
assign t[12964] = t[12963] ^ n[12964];
assign t[12965] = t[12964] ^ n[12965];
assign t[12966] = t[12965] ^ n[12966];
assign t[12967] = t[12966] ^ n[12967];
assign t[12968] = t[12967] ^ n[12968];
assign t[12969] = t[12968] ^ n[12969];
assign t[12970] = t[12969] ^ n[12970];
assign t[12971] = t[12970] ^ n[12971];
assign t[12972] = t[12971] ^ n[12972];
assign t[12973] = t[12972] ^ n[12973];
assign t[12974] = t[12973] ^ n[12974];
assign t[12975] = t[12974] ^ n[12975];
assign t[12976] = t[12975] ^ n[12976];
assign t[12977] = t[12976] ^ n[12977];
assign t[12978] = t[12977] ^ n[12978];
assign t[12979] = t[12978] ^ n[12979];
assign t[12980] = t[12979] ^ n[12980];
assign t[12981] = t[12980] ^ n[12981];
assign t[12982] = t[12981] ^ n[12982];
assign t[12983] = t[12982] ^ n[12983];
assign t[12984] = t[12983] ^ n[12984];
assign t[12985] = t[12984] ^ n[12985];
assign t[12986] = t[12985] ^ n[12986];
assign t[12987] = t[12986] ^ n[12987];
assign t[12988] = t[12987] ^ n[12988];
assign t[12989] = t[12988] ^ n[12989];
assign t[12990] = t[12989] ^ n[12990];
assign t[12991] = t[12990] ^ n[12991];
assign t[12992] = t[12991] ^ n[12992];
assign t[12993] = t[12992] ^ n[12993];
assign t[12994] = t[12993] ^ n[12994];
assign t[12995] = t[12994] ^ n[12995];
assign t[12996] = t[12995] ^ n[12996];
assign t[12997] = t[12996] ^ n[12997];
assign t[12998] = t[12997] ^ n[12998];
assign t[12999] = t[12998] ^ n[12999];
assign t[13000] = t[12999] ^ n[13000];
assign t[13001] = t[13000] ^ n[13001];
assign t[13002] = t[13001] ^ n[13002];
assign t[13003] = t[13002] ^ n[13003];
assign t[13004] = t[13003] ^ n[13004];
assign t[13005] = t[13004] ^ n[13005];
assign t[13006] = t[13005] ^ n[13006];
assign t[13007] = t[13006] ^ n[13007];
assign t[13008] = t[13007] ^ n[13008];
assign t[13009] = t[13008] ^ n[13009];
assign t[13010] = t[13009] ^ n[13010];
assign t[13011] = t[13010] ^ n[13011];
assign t[13012] = t[13011] ^ n[13012];
assign t[13013] = t[13012] ^ n[13013];
assign t[13014] = t[13013] ^ n[13014];
assign t[13015] = t[13014] ^ n[13015];
assign t[13016] = t[13015] ^ n[13016];
assign t[13017] = t[13016] ^ n[13017];
assign t[13018] = t[13017] ^ n[13018];
assign t[13019] = t[13018] ^ n[13019];
assign t[13020] = t[13019] ^ n[13020];
assign t[13021] = t[13020] ^ n[13021];
assign t[13022] = t[13021] ^ n[13022];
assign t[13023] = t[13022] ^ n[13023];
assign t[13024] = t[13023] ^ n[13024];
assign t[13025] = t[13024] ^ n[13025];
assign t[13026] = t[13025] ^ n[13026];
assign t[13027] = t[13026] ^ n[13027];
assign t[13028] = t[13027] ^ n[13028];
assign t[13029] = t[13028] ^ n[13029];
assign t[13030] = t[13029] ^ n[13030];
assign t[13031] = t[13030] ^ n[13031];
assign t[13032] = t[13031] ^ n[13032];
assign t[13033] = t[13032] ^ n[13033];
assign t[13034] = t[13033] ^ n[13034];
assign t[13035] = t[13034] ^ n[13035];
assign t[13036] = t[13035] ^ n[13036];
assign t[13037] = t[13036] ^ n[13037];
assign t[13038] = t[13037] ^ n[13038];
assign t[13039] = t[13038] ^ n[13039];
assign t[13040] = t[13039] ^ n[13040];
assign t[13041] = t[13040] ^ n[13041];
assign t[13042] = t[13041] ^ n[13042];
assign t[13043] = t[13042] ^ n[13043];
assign t[13044] = t[13043] ^ n[13044];
assign t[13045] = t[13044] ^ n[13045];
assign t[13046] = t[13045] ^ n[13046];
assign t[13047] = t[13046] ^ n[13047];
assign t[13048] = t[13047] ^ n[13048];
assign t[13049] = t[13048] ^ n[13049];
assign t[13050] = t[13049] ^ n[13050];
assign t[13051] = t[13050] ^ n[13051];
assign t[13052] = t[13051] ^ n[13052];
assign t[13053] = t[13052] ^ n[13053];
assign t[13054] = t[13053] ^ n[13054];
assign t[13055] = t[13054] ^ n[13055];
assign t[13056] = t[13055] ^ n[13056];
assign t[13057] = t[13056] ^ n[13057];
assign t[13058] = t[13057] ^ n[13058];
assign t[13059] = t[13058] ^ n[13059];
assign t[13060] = t[13059] ^ n[13060];
assign t[13061] = t[13060] ^ n[13061];
assign t[13062] = t[13061] ^ n[13062];
assign t[13063] = t[13062] ^ n[13063];
assign t[13064] = t[13063] ^ n[13064];
assign t[13065] = t[13064] ^ n[13065];
assign t[13066] = t[13065] ^ n[13066];
assign t[13067] = t[13066] ^ n[13067];
assign t[13068] = t[13067] ^ n[13068];
assign t[13069] = t[13068] ^ n[13069];
assign t[13070] = t[13069] ^ n[13070];
assign t[13071] = t[13070] ^ n[13071];
assign t[13072] = t[13071] ^ n[13072];
assign t[13073] = t[13072] ^ n[13073];
assign t[13074] = t[13073] ^ n[13074];
assign t[13075] = t[13074] ^ n[13075];
assign t[13076] = t[13075] ^ n[13076];
assign t[13077] = t[13076] ^ n[13077];
assign t[13078] = t[13077] ^ n[13078];
assign t[13079] = t[13078] ^ n[13079];
assign t[13080] = t[13079] ^ n[13080];
assign t[13081] = t[13080] ^ n[13081];
assign t[13082] = t[13081] ^ n[13082];
assign t[13083] = t[13082] ^ n[13083];
assign t[13084] = t[13083] ^ n[13084];
assign t[13085] = t[13084] ^ n[13085];
assign t[13086] = t[13085] ^ n[13086];
assign t[13087] = t[13086] ^ n[13087];
assign t[13088] = t[13087] ^ n[13088];
assign t[13089] = t[13088] ^ n[13089];
assign t[13090] = t[13089] ^ n[13090];
assign t[13091] = t[13090] ^ n[13091];
assign t[13092] = t[13091] ^ n[13092];
assign t[13093] = t[13092] ^ n[13093];
assign t[13094] = t[13093] ^ n[13094];
assign t[13095] = t[13094] ^ n[13095];
assign t[13096] = t[13095] ^ n[13096];
assign t[13097] = t[13096] ^ n[13097];
assign t[13098] = t[13097] ^ n[13098];
assign t[13099] = t[13098] ^ n[13099];
assign t[13100] = t[13099] ^ n[13100];
assign t[13101] = t[13100] ^ n[13101];
assign t[13102] = t[13101] ^ n[13102];
assign t[13103] = t[13102] ^ n[13103];
assign t[13104] = t[13103] ^ n[13104];
assign t[13105] = t[13104] ^ n[13105];
assign t[13106] = t[13105] ^ n[13106];
assign t[13107] = t[13106] ^ n[13107];
assign t[13108] = t[13107] ^ n[13108];
assign t[13109] = t[13108] ^ n[13109];
assign t[13110] = t[13109] ^ n[13110];
assign t[13111] = t[13110] ^ n[13111];
assign t[13112] = t[13111] ^ n[13112];
assign t[13113] = t[13112] ^ n[13113];
assign t[13114] = t[13113] ^ n[13114];
assign t[13115] = t[13114] ^ n[13115];
assign t[13116] = t[13115] ^ n[13116];
assign t[13117] = t[13116] ^ n[13117];
assign t[13118] = t[13117] ^ n[13118];
assign t[13119] = t[13118] ^ n[13119];
assign t[13120] = t[13119] ^ n[13120];
assign t[13121] = t[13120] ^ n[13121];
assign t[13122] = t[13121] ^ n[13122];
assign t[13123] = t[13122] ^ n[13123];
assign t[13124] = t[13123] ^ n[13124];
assign t[13125] = t[13124] ^ n[13125];
assign t[13126] = t[13125] ^ n[13126];
assign t[13127] = t[13126] ^ n[13127];
assign t[13128] = t[13127] ^ n[13128];
assign t[13129] = t[13128] ^ n[13129];
assign t[13130] = t[13129] ^ n[13130];
assign t[13131] = t[13130] ^ n[13131];
assign t[13132] = t[13131] ^ n[13132];
assign t[13133] = t[13132] ^ n[13133];
assign t[13134] = t[13133] ^ n[13134];
assign t[13135] = t[13134] ^ n[13135];
assign t[13136] = t[13135] ^ n[13136];
assign t[13137] = t[13136] ^ n[13137];
assign t[13138] = t[13137] ^ n[13138];
assign t[13139] = t[13138] ^ n[13139];
assign t[13140] = t[13139] ^ n[13140];
assign t[13141] = t[13140] ^ n[13141];
assign t[13142] = t[13141] ^ n[13142];
assign t[13143] = t[13142] ^ n[13143];
assign t[13144] = t[13143] ^ n[13144];
assign t[13145] = t[13144] ^ n[13145];
assign t[13146] = t[13145] ^ n[13146];
assign t[13147] = t[13146] ^ n[13147];
assign t[13148] = t[13147] ^ n[13148];
assign t[13149] = t[13148] ^ n[13149];
assign t[13150] = t[13149] ^ n[13150];
assign t[13151] = t[13150] ^ n[13151];
assign t[13152] = t[13151] ^ n[13152];
assign t[13153] = t[13152] ^ n[13153];
assign t[13154] = t[13153] ^ n[13154];
assign t[13155] = t[13154] ^ n[13155];
assign t[13156] = t[13155] ^ n[13156];
assign t[13157] = t[13156] ^ n[13157];
assign t[13158] = t[13157] ^ n[13158];
assign t[13159] = t[13158] ^ n[13159];
assign t[13160] = t[13159] ^ n[13160];
assign t[13161] = t[13160] ^ n[13161];
assign t[13162] = t[13161] ^ n[13162];
assign t[13163] = t[13162] ^ n[13163];
assign t[13164] = t[13163] ^ n[13164];
assign t[13165] = t[13164] ^ n[13165];
assign t[13166] = t[13165] ^ n[13166];
assign t[13167] = t[13166] ^ n[13167];
assign t[13168] = t[13167] ^ n[13168];
assign t[13169] = t[13168] ^ n[13169];
assign t[13170] = t[13169] ^ n[13170];
assign t[13171] = t[13170] ^ n[13171];
assign t[13172] = t[13171] ^ n[13172];
assign t[13173] = t[13172] ^ n[13173];
assign t[13174] = t[13173] ^ n[13174];
assign t[13175] = t[13174] ^ n[13175];
assign t[13176] = t[13175] ^ n[13176];
assign t[13177] = t[13176] ^ n[13177];
assign t[13178] = t[13177] ^ n[13178];
assign t[13179] = t[13178] ^ n[13179];
assign t[13180] = t[13179] ^ n[13180];
assign t[13181] = t[13180] ^ n[13181];
assign t[13182] = t[13181] ^ n[13182];
assign t[13183] = t[13182] ^ n[13183];
assign t[13184] = t[13183] ^ n[13184];
assign t[13185] = t[13184] ^ n[13185];
assign t[13186] = t[13185] ^ n[13186];
assign t[13187] = t[13186] ^ n[13187];
assign t[13188] = t[13187] ^ n[13188];
assign t[13189] = t[13188] ^ n[13189];
assign t[13190] = t[13189] ^ n[13190];
assign t[13191] = t[13190] ^ n[13191];
assign t[13192] = t[13191] ^ n[13192];
assign t[13193] = t[13192] ^ n[13193];
assign t[13194] = t[13193] ^ n[13194];
assign t[13195] = t[13194] ^ n[13195];
assign t[13196] = t[13195] ^ n[13196];
assign t[13197] = t[13196] ^ n[13197];
assign t[13198] = t[13197] ^ n[13198];
assign t[13199] = t[13198] ^ n[13199];
assign t[13200] = t[13199] ^ n[13200];
assign t[13201] = t[13200] ^ n[13201];
assign t[13202] = t[13201] ^ n[13202];
assign t[13203] = t[13202] ^ n[13203];
assign t[13204] = t[13203] ^ n[13204];
assign t[13205] = t[13204] ^ n[13205];
assign t[13206] = t[13205] ^ n[13206];
assign t[13207] = t[13206] ^ n[13207];
assign t[13208] = t[13207] ^ n[13208];
assign t[13209] = t[13208] ^ n[13209];
assign t[13210] = t[13209] ^ n[13210];
assign t[13211] = t[13210] ^ n[13211];
assign t[13212] = t[13211] ^ n[13212];
assign t[13213] = t[13212] ^ n[13213];
assign t[13214] = t[13213] ^ n[13214];
assign t[13215] = t[13214] ^ n[13215];
assign t[13216] = t[13215] ^ n[13216];
assign t[13217] = t[13216] ^ n[13217];
assign t[13218] = t[13217] ^ n[13218];
assign t[13219] = t[13218] ^ n[13219];
assign t[13220] = t[13219] ^ n[13220];
assign t[13221] = t[13220] ^ n[13221];
assign t[13222] = t[13221] ^ n[13222];
assign t[13223] = t[13222] ^ n[13223];
assign t[13224] = t[13223] ^ n[13224];
assign t[13225] = t[13224] ^ n[13225];
assign t[13226] = t[13225] ^ n[13226];
assign t[13227] = t[13226] ^ n[13227];
assign t[13228] = t[13227] ^ n[13228];
assign t[13229] = t[13228] ^ n[13229];
assign t[13230] = t[13229] ^ n[13230];
assign t[13231] = t[13230] ^ n[13231];
assign t[13232] = t[13231] ^ n[13232];
assign t[13233] = t[13232] ^ n[13233];
assign t[13234] = t[13233] ^ n[13234];
assign t[13235] = t[13234] ^ n[13235];
assign t[13236] = t[13235] ^ n[13236];
assign t[13237] = t[13236] ^ n[13237];
assign t[13238] = t[13237] ^ n[13238];
assign t[13239] = t[13238] ^ n[13239];
assign t[13240] = t[13239] ^ n[13240];
assign t[13241] = t[13240] ^ n[13241];
assign t[13242] = t[13241] ^ n[13242];
assign t[13243] = t[13242] ^ n[13243];
assign t[13244] = t[13243] ^ n[13244];
assign t[13245] = t[13244] ^ n[13245];
assign t[13246] = t[13245] ^ n[13246];
assign t[13247] = t[13246] ^ n[13247];
assign t[13248] = t[13247] ^ n[13248];
assign t[13249] = t[13248] ^ n[13249];
assign t[13250] = t[13249] ^ n[13250];
assign t[13251] = t[13250] ^ n[13251];
assign t[13252] = t[13251] ^ n[13252];
assign t[13253] = t[13252] ^ n[13253];
assign t[13254] = t[13253] ^ n[13254];
assign t[13255] = t[13254] ^ n[13255];
assign t[13256] = t[13255] ^ n[13256];
assign t[13257] = t[13256] ^ n[13257];
assign t[13258] = t[13257] ^ n[13258];
assign t[13259] = t[13258] ^ n[13259];
assign t[13260] = t[13259] ^ n[13260];
assign t[13261] = t[13260] ^ n[13261];
assign t[13262] = t[13261] ^ n[13262];
assign t[13263] = t[13262] ^ n[13263];
assign t[13264] = t[13263] ^ n[13264];
assign t[13265] = t[13264] ^ n[13265];
assign t[13266] = t[13265] ^ n[13266];
assign t[13267] = t[13266] ^ n[13267];
assign t[13268] = t[13267] ^ n[13268];
assign t[13269] = t[13268] ^ n[13269];
assign t[13270] = t[13269] ^ n[13270];
assign t[13271] = t[13270] ^ n[13271];
assign t[13272] = t[13271] ^ n[13272];
assign t[13273] = t[13272] ^ n[13273];
assign t[13274] = t[13273] ^ n[13274];
assign t[13275] = t[13274] ^ n[13275];
assign t[13276] = t[13275] ^ n[13276];
assign t[13277] = t[13276] ^ n[13277];
assign t[13278] = t[13277] ^ n[13278];
assign t[13279] = t[13278] ^ n[13279];
assign t[13280] = t[13279] ^ n[13280];
assign t[13281] = t[13280] ^ n[13281];
assign t[13282] = t[13281] ^ n[13282];
assign t[13283] = t[13282] ^ n[13283];
assign t[13284] = t[13283] ^ n[13284];
assign t[13285] = t[13284] ^ n[13285];
assign t[13286] = t[13285] ^ n[13286];
assign t[13287] = t[13286] ^ n[13287];
assign t[13288] = t[13287] ^ n[13288];
assign t[13289] = t[13288] ^ n[13289];
assign t[13290] = t[13289] ^ n[13290];
assign t[13291] = t[13290] ^ n[13291];
assign t[13292] = t[13291] ^ n[13292];
assign t[13293] = t[13292] ^ n[13293];
assign t[13294] = t[13293] ^ n[13294];
assign t[13295] = t[13294] ^ n[13295];
assign t[13296] = t[13295] ^ n[13296];
assign t[13297] = t[13296] ^ n[13297];
assign t[13298] = t[13297] ^ n[13298];
assign t[13299] = t[13298] ^ n[13299];
assign t[13300] = t[13299] ^ n[13300];
assign t[13301] = t[13300] ^ n[13301];
assign t[13302] = t[13301] ^ n[13302];
assign t[13303] = t[13302] ^ n[13303];
assign t[13304] = t[13303] ^ n[13304];
assign t[13305] = t[13304] ^ n[13305];
assign t[13306] = t[13305] ^ n[13306];
assign t[13307] = t[13306] ^ n[13307];
assign t[13308] = t[13307] ^ n[13308];
assign t[13309] = t[13308] ^ n[13309];
assign t[13310] = t[13309] ^ n[13310];
assign t[13311] = t[13310] ^ n[13311];
assign t[13312] = t[13311] ^ n[13312];
assign t[13313] = t[13312] ^ n[13313];
assign t[13314] = t[13313] ^ n[13314];
assign t[13315] = t[13314] ^ n[13315];
assign t[13316] = t[13315] ^ n[13316];
assign t[13317] = t[13316] ^ n[13317];
assign t[13318] = t[13317] ^ n[13318];
assign t[13319] = t[13318] ^ n[13319];
assign t[13320] = t[13319] ^ n[13320];
assign t[13321] = t[13320] ^ n[13321];
assign t[13322] = t[13321] ^ n[13322];
assign t[13323] = t[13322] ^ n[13323];
assign t[13324] = t[13323] ^ n[13324];
assign t[13325] = t[13324] ^ n[13325];
assign t[13326] = t[13325] ^ n[13326];
assign t[13327] = t[13326] ^ n[13327];
assign t[13328] = t[13327] ^ n[13328];
assign t[13329] = t[13328] ^ n[13329];
assign t[13330] = t[13329] ^ n[13330];
assign t[13331] = t[13330] ^ n[13331];
assign t[13332] = t[13331] ^ n[13332];
assign t[13333] = t[13332] ^ n[13333];
assign t[13334] = t[13333] ^ n[13334];
assign t[13335] = t[13334] ^ n[13335];
assign t[13336] = t[13335] ^ n[13336];
assign t[13337] = t[13336] ^ n[13337];
assign t[13338] = t[13337] ^ n[13338];
assign t[13339] = t[13338] ^ n[13339];
assign t[13340] = t[13339] ^ n[13340];
assign t[13341] = t[13340] ^ n[13341];
assign t[13342] = t[13341] ^ n[13342];
assign t[13343] = t[13342] ^ n[13343];
assign t[13344] = t[13343] ^ n[13344];
assign t[13345] = t[13344] ^ n[13345];
assign t[13346] = t[13345] ^ n[13346];
assign t[13347] = t[13346] ^ n[13347];
assign t[13348] = t[13347] ^ n[13348];
assign t[13349] = t[13348] ^ n[13349];
assign t[13350] = t[13349] ^ n[13350];
assign t[13351] = t[13350] ^ n[13351];
assign t[13352] = t[13351] ^ n[13352];
assign t[13353] = t[13352] ^ n[13353];
assign t[13354] = t[13353] ^ n[13354];
assign t[13355] = t[13354] ^ n[13355];
assign t[13356] = t[13355] ^ n[13356];
assign t[13357] = t[13356] ^ n[13357];
assign t[13358] = t[13357] ^ n[13358];
assign t[13359] = t[13358] ^ n[13359];
assign t[13360] = t[13359] ^ n[13360];
assign t[13361] = t[13360] ^ n[13361];
assign t[13362] = t[13361] ^ n[13362];
assign t[13363] = t[13362] ^ n[13363];
assign t[13364] = t[13363] ^ n[13364];
assign t[13365] = t[13364] ^ n[13365];
assign t[13366] = t[13365] ^ n[13366];
assign t[13367] = t[13366] ^ n[13367];
assign t[13368] = t[13367] ^ n[13368];
assign t[13369] = t[13368] ^ n[13369];
assign t[13370] = t[13369] ^ n[13370];
assign t[13371] = t[13370] ^ n[13371];
assign t[13372] = t[13371] ^ n[13372];
assign t[13373] = t[13372] ^ n[13373];
assign t[13374] = t[13373] ^ n[13374];
assign t[13375] = t[13374] ^ n[13375];
assign t[13376] = t[13375] ^ n[13376];
assign t[13377] = t[13376] ^ n[13377];
assign t[13378] = t[13377] ^ n[13378];
assign t[13379] = t[13378] ^ n[13379];
assign t[13380] = t[13379] ^ n[13380];
assign t[13381] = t[13380] ^ n[13381];
assign t[13382] = t[13381] ^ n[13382];
assign t[13383] = t[13382] ^ n[13383];
assign t[13384] = t[13383] ^ n[13384];
assign t[13385] = t[13384] ^ n[13385];
assign t[13386] = t[13385] ^ n[13386];
assign t[13387] = t[13386] ^ n[13387];
assign t[13388] = t[13387] ^ n[13388];
assign t[13389] = t[13388] ^ n[13389];
assign t[13390] = t[13389] ^ n[13390];
assign t[13391] = t[13390] ^ n[13391];
assign t[13392] = t[13391] ^ n[13392];
assign t[13393] = t[13392] ^ n[13393];
assign t[13394] = t[13393] ^ n[13394];
assign t[13395] = t[13394] ^ n[13395];
assign t[13396] = t[13395] ^ n[13396];
assign t[13397] = t[13396] ^ n[13397];
assign t[13398] = t[13397] ^ n[13398];
assign t[13399] = t[13398] ^ n[13399];
assign t[13400] = t[13399] ^ n[13400];
assign t[13401] = t[13400] ^ n[13401];
assign t[13402] = t[13401] ^ n[13402];
assign t[13403] = t[13402] ^ n[13403];
assign t[13404] = t[13403] ^ n[13404];
assign t[13405] = t[13404] ^ n[13405];
assign t[13406] = t[13405] ^ n[13406];
assign t[13407] = t[13406] ^ n[13407];
assign t[13408] = t[13407] ^ n[13408];
assign t[13409] = t[13408] ^ n[13409];
assign t[13410] = t[13409] ^ n[13410];
assign t[13411] = t[13410] ^ n[13411];
assign t[13412] = t[13411] ^ n[13412];
assign t[13413] = t[13412] ^ n[13413];
assign t[13414] = t[13413] ^ n[13414];
assign t[13415] = t[13414] ^ n[13415];
assign t[13416] = t[13415] ^ n[13416];
assign t[13417] = t[13416] ^ n[13417];
assign t[13418] = t[13417] ^ n[13418];
assign t[13419] = t[13418] ^ n[13419];
assign t[13420] = t[13419] ^ n[13420];
assign t[13421] = t[13420] ^ n[13421];
assign t[13422] = t[13421] ^ n[13422];
assign t[13423] = t[13422] ^ n[13423];
assign t[13424] = t[13423] ^ n[13424];
assign t[13425] = t[13424] ^ n[13425];
assign t[13426] = t[13425] ^ n[13426];
assign t[13427] = t[13426] ^ n[13427];
assign t[13428] = t[13427] ^ n[13428];
assign t[13429] = t[13428] ^ n[13429];
assign t[13430] = t[13429] ^ n[13430];
assign t[13431] = t[13430] ^ n[13431];
assign t[13432] = t[13431] ^ n[13432];
assign t[13433] = t[13432] ^ n[13433];
assign t[13434] = t[13433] ^ n[13434];
assign t[13435] = t[13434] ^ n[13435];
assign t[13436] = t[13435] ^ n[13436];
assign t[13437] = t[13436] ^ n[13437];
assign t[13438] = t[13437] ^ n[13438];
assign t[13439] = t[13438] ^ n[13439];
assign t[13440] = t[13439] ^ n[13440];
assign t[13441] = t[13440] ^ n[13441];
assign t[13442] = t[13441] ^ n[13442];
assign t[13443] = t[13442] ^ n[13443];
assign t[13444] = t[13443] ^ n[13444];
assign t[13445] = t[13444] ^ n[13445];
assign t[13446] = t[13445] ^ n[13446];
assign t[13447] = t[13446] ^ n[13447];
assign t[13448] = t[13447] ^ n[13448];
assign t[13449] = t[13448] ^ n[13449];
assign t[13450] = t[13449] ^ n[13450];
assign t[13451] = t[13450] ^ n[13451];
assign t[13452] = t[13451] ^ n[13452];
assign t[13453] = t[13452] ^ n[13453];
assign t[13454] = t[13453] ^ n[13454];
assign t[13455] = t[13454] ^ n[13455];
assign t[13456] = t[13455] ^ n[13456];
assign t[13457] = t[13456] ^ n[13457];
assign t[13458] = t[13457] ^ n[13458];
assign t[13459] = t[13458] ^ n[13459];
assign t[13460] = t[13459] ^ n[13460];
assign t[13461] = t[13460] ^ n[13461];
assign t[13462] = t[13461] ^ n[13462];
assign t[13463] = t[13462] ^ n[13463];
assign t[13464] = t[13463] ^ n[13464];
assign t[13465] = t[13464] ^ n[13465];
assign t[13466] = t[13465] ^ n[13466];
assign t[13467] = t[13466] ^ n[13467];
assign t[13468] = t[13467] ^ n[13468];
assign t[13469] = t[13468] ^ n[13469];
assign t[13470] = t[13469] ^ n[13470];
assign t[13471] = t[13470] ^ n[13471];
assign t[13472] = t[13471] ^ n[13472];
assign t[13473] = t[13472] ^ n[13473];
assign t[13474] = t[13473] ^ n[13474];
assign t[13475] = t[13474] ^ n[13475];
assign t[13476] = t[13475] ^ n[13476];
assign t[13477] = t[13476] ^ n[13477];
assign t[13478] = t[13477] ^ n[13478];
assign t[13479] = t[13478] ^ n[13479];
assign t[13480] = t[13479] ^ n[13480];
assign t[13481] = t[13480] ^ n[13481];
assign t[13482] = t[13481] ^ n[13482];
assign t[13483] = t[13482] ^ n[13483];
assign t[13484] = t[13483] ^ n[13484];
assign t[13485] = t[13484] ^ n[13485];
assign t[13486] = t[13485] ^ n[13486];
assign t[13487] = t[13486] ^ n[13487];
assign t[13488] = t[13487] ^ n[13488];
assign t[13489] = t[13488] ^ n[13489];
assign t[13490] = t[13489] ^ n[13490];
assign t[13491] = t[13490] ^ n[13491];
assign t[13492] = t[13491] ^ n[13492];
assign t[13493] = t[13492] ^ n[13493];
assign t[13494] = t[13493] ^ n[13494];
assign t[13495] = t[13494] ^ n[13495];
assign t[13496] = t[13495] ^ n[13496];
assign t[13497] = t[13496] ^ n[13497];
assign t[13498] = t[13497] ^ n[13498];
assign t[13499] = t[13498] ^ n[13499];
assign t[13500] = t[13499] ^ n[13500];
assign t[13501] = t[13500] ^ n[13501];
assign t[13502] = t[13501] ^ n[13502];
assign t[13503] = t[13502] ^ n[13503];
assign t[13504] = t[13503] ^ n[13504];
assign t[13505] = t[13504] ^ n[13505];
assign t[13506] = t[13505] ^ n[13506];
assign t[13507] = t[13506] ^ n[13507];
assign t[13508] = t[13507] ^ n[13508];
assign t[13509] = t[13508] ^ n[13509];
assign t[13510] = t[13509] ^ n[13510];
assign t[13511] = t[13510] ^ n[13511];
assign t[13512] = t[13511] ^ n[13512];
assign t[13513] = t[13512] ^ n[13513];
assign t[13514] = t[13513] ^ n[13514];
assign t[13515] = t[13514] ^ n[13515];
assign t[13516] = t[13515] ^ n[13516];
assign t[13517] = t[13516] ^ n[13517];
assign t[13518] = t[13517] ^ n[13518];
assign t[13519] = t[13518] ^ n[13519];
assign t[13520] = t[13519] ^ n[13520];
assign t[13521] = t[13520] ^ n[13521];
assign t[13522] = t[13521] ^ n[13522];
assign t[13523] = t[13522] ^ n[13523];
assign t[13524] = t[13523] ^ n[13524];
assign t[13525] = t[13524] ^ n[13525];
assign t[13526] = t[13525] ^ n[13526];
assign t[13527] = t[13526] ^ n[13527];
assign t[13528] = t[13527] ^ n[13528];
assign t[13529] = t[13528] ^ n[13529];
assign t[13530] = t[13529] ^ n[13530];
assign t[13531] = t[13530] ^ n[13531];
assign t[13532] = t[13531] ^ n[13532];
assign t[13533] = t[13532] ^ n[13533];
assign t[13534] = t[13533] ^ n[13534];
assign t[13535] = t[13534] ^ n[13535];
assign t[13536] = t[13535] ^ n[13536];
assign t[13537] = t[13536] ^ n[13537];
assign t[13538] = t[13537] ^ n[13538];
assign t[13539] = t[13538] ^ n[13539];
assign t[13540] = t[13539] ^ n[13540];
assign t[13541] = t[13540] ^ n[13541];
assign t[13542] = t[13541] ^ n[13542];
assign t[13543] = t[13542] ^ n[13543];
assign t[13544] = t[13543] ^ n[13544];
assign t[13545] = t[13544] ^ n[13545];
assign t[13546] = t[13545] ^ n[13546];
assign t[13547] = t[13546] ^ n[13547];
assign t[13548] = t[13547] ^ n[13548];
assign t[13549] = t[13548] ^ n[13549];
assign t[13550] = t[13549] ^ n[13550];
assign t[13551] = t[13550] ^ n[13551];
assign t[13552] = t[13551] ^ n[13552];
assign t[13553] = t[13552] ^ n[13553];
assign t[13554] = t[13553] ^ n[13554];
assign t[13555] = t[13554] ^ n[13555];
assign t[13556] = t[13555] ^ n[13556];
assign t[13557] = t[13556] ^ n[13557];
assign t[13558] = t[13557] ^ n[13558];
assign t[13559] = t[13558] ^ n[13559];
assign t[13560] = t[13559] ^ n[13560];
assign t[13561] = t[13560] ^ n[13561];
assign t[13562] = t[13561] ^ n[13562];
assign t[13563] = t[13562] ^ n[13563];
assign t[13564] = t[13563] ^ n[13564];
assign t[13565] = t[13564] ^ n[13565];
assign t[13566] = t[13565] ^ n[13566];
assign t[13567] = t[13566] ^ n[13567];
assign t[13568] = t[13567] ^ n[13568];
assign t[13569] = t[13568] ^ n[13569];
assign t[13570] = t[13569] ^ n[13570];
assign t[13571] = t[13570] ^ n[13571];
assign t[13572] = t[13571] ^ n[13572];
assign t[13573] = t[13572] ^ n[13573];
assign t[13574] = t[13573] ^ n[13574];
assign t[13575] = t[13574] ^ n[13575];
assign t[13576] = t[13575] ^ n[13576];
assign t[13577] = t[13576] ^ n[13577];
assign t[13578] = t[13577] ^ n[13578];
assign t[13579] = t[13578] ^ n[13579];
assign t[13580] = t[13579] ^ n[13580];
assign t[13581] = t[13580] ^ n[13581];
assign t[13582] = t[13581] ^ n[13582];
assign t[13583] = t[13582] ^ n[13583];
assign t[13584] = t[13583] ^ n[13584];
assign t[13585] = t[13584] ^ n[13585];
assign t[13586] = t[13585] ^ n[13586];
assign t[13587] = t[13586] ^ n[13587];
assign t[13588] = t[13587] ^ n[13588];
assign t[13589] = t[13588] ^ n[13589];
assign t[13590] = t[13589] ^ n[13590];
assign t[13591] = t[13590] ^ n[13591];
assign t[13592] = t[13591] ^ n[13592];
assign t[13593] = t[13592] ^ n[13593];
assign t[13594] = t[13593] ^ n[13594];
assign t[13595] = t[13594] ^ n[13595];
assign t[13596] = t[13595] ^ n[13596];
assign t[13597] = t[13596] ^ n[13597];
assign t[13598] = t[13597] ^ n[13598];
assign t[13599] = t[13598] ^ n[13599];
assign t[13600] = t[13599] ^ n[13600];
assign t[13601] = t[13600] ^ n[13601];
assign t[13602] = t[13601] ^ n[13602];
assign t[13603] = t[13602] ^ n[13603];
assign t[13604] = t[13603] ^ n[13604];
assign t[13605] = t[13604] ^ n[13605];
assign t[13606] = t[13605] ^ n[13606];
assign t[13607] = t[13606] ^ n[13607];
assign t[13608] = t[13607] ^ n[13608];
assign t[13609] = t[13608] ^ n[13609];
assign t[13610] = t[13609] ^ n[13610];
assign t[13611] = t[13610] ^ n[13611];
assign t[13612] = t[13611] ^ n[13612];
assign t[13613] = t[13612] ^ n[13613];
assign t[13614] = t[13613] ^ n[13614];
assign t[13615] = t[13614] ^ n[13615];
assign t[13616] = t[13615] ^ n[13616];
assign t[13617] = t[13616] ^ n[13617];
assign t[13618] = t[13617] ^ n[13618];
assign t[13619] = t[13618] ^ n[13619];
assign t[13620] = t[13619] ^ n[13620];
assign t[13621] = t[13620] ^ n[13621];
assign t[13622] = t[13621] ^ n[13622];
assign t[13623] = t[13622] ^ n[13623];
assign t[13624] = t[13623] ^ n[13624];
assign t[13625] = t[13624] ^ n[13625];
assign t[13626] = t[13625] ^ n[13626];
assign t[13627] = t[13626] ^ n[13627];
assign t[13628] = t[13627] ^ n[13628];
assign t[13629] = t[13628] ^ n[13629];
assign t[13630] = t[13629] ^ n[13630];
assign t[13631] = t[13630] ^ n[13631];
assign t[13632] = t[13631] ^ n[13632];
assign t[13633] = t[13632] ^ n[13633];
assign t[13634] = t[13633] ^ n[13634];
assign t[13635] = t[13634] ^ n[13635];
assign t[13636] = t[13635] ^ n[13636];
assign t[13637] = t[13636] ^ n[13637];
assign t[13638] = t[13637] ^ n[13638];
assign t[13639] = t[13638] ^ n[13639];
assign t[13640] = t[13639] ^ n[13640];
assign t[13641] = t[13640] ^ n[13641];
assign t[13642] = t[13641] ^ n[13642];
assign t[13643] = t[13642] ^ n[13643];
assign t[13644] = t[13643] ^ n[13644];
assign t[13645] = t[13644] ^ n[13645];
assign t[13646] = t[13645] ^ n[13646];
assign t[13647] = t[13646] ^ n[13647];
assign t[13648] = t[13647] ^ n[13648];
assign t[13649] = t[13648] ^ n[13649];
assign t[13650] = t[13649] ^ n[13650];
assign t[13651] = t[13650] ^ n[13651];
assign t[13652] = t[13651] ^ n[13652];
assign t[13653] = t[13652] ^ n[13653];
assign t[13654] = t[13653] ^ n[13654];
assign t[13655] = t[13654] ^ n[13655];
assign t[13656] = t[13655] ^ n[13656];
assign t[13657] = t[13656] ^ n[13657];
assign t[13658] = t[13657] ^ n[13658];
assign t[13659] = t[13658] ^ n[13659];
assign t[13660] = t[13659] ^ n[13660];
assign t[13661] = t[13660] ^ n[13661];
assign t[13662] = t[13661] ^ n[13662];
assign t[13663] = t[13662] ^ n[13663];
assign t[13664] = t[13663] ^ n[13664];
assign t[13665] = t[13664] ^ n[13665];
assign t[13666] = t[13665] ^ n[13666];
assign t[13667] = t[13666] ^ n[13667];
assign t[13668] = t[13667] ^ n[13668];
assign t[13669] = t[13668] ^ n[13669];
assign t[13670] = t[13669] ^ n[13670];
assign t[13671] = t[13670] ^ n[13671];
assign t[13672] = t[13671] ^ n[13672];
assign t[13673] = t[13672] ^ n[13673];
assign t[13674] = t[13673] ^ n[13674];
assign t[13675] = t[13674] ^ n[13675];
assign t[13676] = t[13675] ^ n[13676];
assign t[13677] = t[13676] ^ n[13677];
assign t[13678] = t[13677] ^ n[13678];
assign t[13679] = t[13678] ^ n[13679];
assign t[13680] = t[13679] ^ n[13680];
assign t[13681] = t[13680] ^ n[13681];
assign t[13682] = t[13681] ^ n[13682];
assign t[13683] = t[13682] ^ n[13683];
assign t[13684] = t[13683] ^ n[13684];
assign t[13685] = t[13684] ^ n[13685];
assign t[13686] = t[13685] ^ n[13686];
assign t[13687] = t[13686] ^ n[13687];
assign t[13688] = t[13687] ^ n[13688];
assign t[13689] = t[13688] ^ n[13689];
assign t[13690] = t[13689] ^ n[13690];
assign t[13691] = t[13690] ^ n[13691];
assign t[13692] = t[13691] ^ n[13692];
assign t[13693] = t[13692] ^ n[13693];
assign t[13694] = t[13693] ^ n[13694];
assign t[13695] = t[13694] ^ n[13695];
assign t[13696] = t[13695] ^ n[13696];
assign t[13697] = t[13696] ^ n[13697];
assign t[13698] = t[13697] ^ n[13698];
assign t[13699] = t[13698] ^ n[13699];
assign t[13700] = t[13699] ^ n[13700];
assign t[13701] = t[13700] ^ n[13701];
assign t[13702] = t[13701] ^ n[13702];
assign t[13703] = t[13702] ^ n[13703];
assign t[13704] = t[13703] ^ n[13704];
assign t[13705] = t[13704] ^ n[13705];
assign t[13706] = t[13705] ^ n[13706];
assign t[13707] = t[13706] ^ n[13707];
assign t[13708] = t[13707] ^ n[13708];
assign t[13709] = t[13708] ^ n[13709];
assign t[13710] = t[13709] ^ n[13710];
assign t[13711] = t[13710] ^ n[13711];
assign t[13712] = t[13711] ^ n[13712];
assign t[13713] = t[13712] ^ n[13713];
assign t[13714] = t[13713] ^ n[13714];
assign t[13715] = t[13714] ^ n[13715];
assign t[13716] = t[13715] ^ n[13716];
assign t[13717] = t[13716] ^ n[13717];
assign t[13718] = t[13717] ^ n[13718];
assign t[13719] = t[13718] ^ n[13719];
assign t[13720] = t[13719] ^ n[13720];
assign t[13721] = t[13720] ^ n[13721];
assign t[13722] = t[13721] ^ n[13722];
assign t[13723] = t[13722] ^ n[13723];
assign t[13724] = t[13723] ^ n[13724];
assign t[13725] = t[13724] ^ n[13725];
assign t[13726] = t[13725] ^ n[13726];
assign t[13727] = t[13726] ^ n[13727];
assign t[13728] = t[13727] ^ n[13728];
assign t[13729] = t[13728] ^ n[13729];
assign t[13730] = t[13729] ^ n[13730];
assign t[13731] = t[13730] ^ n[13731];
assign t[13732] = t[13731] ^ n[13732];
assign t[13733] = t[13732] ^ n[13733];
assign t[13734] = t[13733] ^ n[13734];
assign t[13735] = t[13734] ^ n[13735];
assign t[13736] = t[13735] ^ n[13736];
assign t[13737] = t[13736] ^ n[13737];
assign t[13738] = t[13737] ^ n[13738];
assign t[13739] = t[13738] ^ n[13739];
assign t[13740] = t[13739] ^ n[13740];
assign t[13741] = t[13740] ^ n[13741];
assign t[13742] = t[13741] ^ n[13742];
assign t[13743] = t[13742] ^ n[13743];
assign t[13744] = t[13743] ^ n[13744];
assign t[13745] = t[13744] ^ n[13745];
assign t[13746] = t[13745] ^ n[13746];
assign t[13747] = t[13746] ^ n[13747];
assign t[13748] = t[13747] ^ n[13748];
assign t[13749] = t[13748] ^ n[13749];
assign t[13750] = t[13749] ^ n[13750];
assign t[13751] = t[13750] ^ n[13751];
assign t[13752] = t[13751] ^ n[13752];
assign t[13753] = t[13752] ^ n[13753];
assign t[13754] = t[13753] ^ n[13754];
assign t[13755] = t[13754] ^ n[13755];
assign t[13756] = t[13755] ^ n[13756];
assign t[13757] = t[13756] ^ n[13757];
assign t[13758] = t[13757] ^ n[13758];
assign t[13759] = t[13758] ^ n[13759];
assign t[13760] = t[13759] ^ n[13760];
assign t[13761] = t[13760] ^ n[13761];
assign t[13762] = t[13761] ^ n[13762];
assign t[13763] = t[13762] ^ n[13763];
assign t[13764] = t[13763] ^ n[13764];
assign t[13765] = t[13764] ^ n[13765];
assign t[13766] = t[13765] ^ n[13766];
assign t[13767] = t[13766] ^ n[13767];
assign t[13768] = t[13767] ^ n[13768];
assign t[13769] = t[13768] ^ n[13769];
assign t[13770] = t[13769] ^ n[13770];
assign t[13771] = t[13770] ^ n[13771];
assign t[13772] = t[13771] ^ n[13772];
assign t[13773] = t[13772] ^ n[13773];
assign t[13774] = t[13773] ^ n[13774];
assign t[13775] = t[13774] ^ n[13775];
assign t[13776] = t[13775] ^ n[13776];
assign t[13777] = t[13776] ^ n[13777];
assign t[13778] = t[13777] ^ n[13778];
assign t[13779] = t[13778] ^ n[13779];
assign t[13780] = t[13779] ^ n[13780];
assign t[13781] = t[13780] ^ n[13781];
assign t[13782] = t[13781] ^ n[13782];
assign t[13783] = t[13782] ^ n[13783];
assign t[13784] = t[13783] ^ n[13784];
assign t[13785] = t[13784] ^ n[13785];
assign t[13786] = t[13785] ^ n[13786];
assign t[13787] = t[13786] ^ n[13787];
assign t[13788] = t[13787] ^ n[13788];
assign t[13789] = t[13788] ^ n[13789];
assign t[13790] = t[13789] ^ n[13790];
assign t[13791] = t[13790] ^ n[13791];
assign t[13792] = t[13791] ^ n[13792];
assign t[13793] = t[13792] ^ n[13793];
assign t[13794] = t[13793] ^ n[13794];
assign t[13795] = t[13794] ^ n[13795];
assign t[13796] = t[13795] ^ n[13796];
assign t[13797] = t[13796] ^ n[13797];
assign t[13798] = t[13797] ^ n[13798];
assign t[13799] = t[13798] ^ n[13799];
assign t[13800] = t[13799] ^ n[13800];
assign t[13801] = t[13800] ^ n[13801];
assign t[13802] = t[13801] ^ n[13802];
assign t[13803] = t[13802] ^ n[13803];
assign t[13804] = t[13803] ^ n[13804];
assign t[13805] = t[13804] ^ n[13805];
assign t[13806] = t[13805] ^ n[13806];
assign t[13807] = t[13806] ^ n[13807];
assign t[13808] = t[13807] ^ n[13808];
assign t[13809] = t[13808] ^ n[13809];
assign t[13810] = t[13809] ^ n[13810];
assign t[13811] = t[13810] ^ n[13811];
assign t[13812] = t[13811] ^ n[13812];
assign t[13813] = t[13812] ^ n[13813];
assign t[13814] = t[13813] ^ n[13814];
assign t[13815] = t[13814] ^ n[13815];
assign t[13816] = t[13815] ^ n[13816];
assign t[13817] = t[13816] ^ n[13817];
assign t[13818] = t[13817] ^ n[13818];
assign t[13819] = t[13818] ^ n[13819];
assign t[13820] = t[13819] ^ n[13820];
assign t[13821] = t[13820] ^ n[13821];
assign t[13822] = t[13821] ^ n[13822];
assign t[13823] = t[13822] ^ n[13823];
assign t[13824] = t[13823] ^ n[13824];
assign t[13825] = t[13824] ^ n[13825];
assign t[13826] = t[13825] ^ n[13826];
assign t[13827] = t[13826] ^ n[13827];
assign t[13828] = t[13827] ^ n[13828];
assign t[13829] = t[13828] ^ n[13829];
assign t[13830] = t[13829] ^ n[13830];
assign t[13831] = t[13830] ^ n[13831];
assign t[13832] = t[13831] ^ n[13832];
assign t[13833] = t[13832] ^ n[13833];
assign t[13834] = t[13833] ^ n[13834];
assign t[13835] = t[13834] ^ n[13835];
assign t[13836] = t[13835] ^ n[13836];
assign t[13837] = t[13836] ^ n[13837];
assign t[13838] = t[13837] ^ n[13838];
assign t[13839] = t[13838] ^ n[13839];
assign t[13840] = t[13839] ^ n[13840];
assign t[13841] = t[13840] ^ n[13841];
assign t[13842] = t[13841] ^ n[13842];
assign t[13843] = t[13842] ^ n[13843];
assign t[13844] = t[13843] ^ n[13844];
assign t[13845] = t[13844] ^ n[13845];
assign t[13846] = t[13845] ^ n[13846];
assign t[13847] = t[13846] ^ n[13847];
assign t[13848] = t[13847] ^ n[13848];
assign t[13849] = t[13848] ^ n[13849];
assign t[13850] = t[13849] ^ n[13850];
assign t[13851] = t[13850] ^ n[13851];
assign t[13852] = t[13851] ^ n[13852];
assign t[13853] = t[13852] ^ n[13853];
assign t[13854] = t[13853] ^ n[13854];
assign t[13855] = t[13854] ^ n[13855];
assign t[13856] = t[13855] ^ n[13856];
assign t[13857] = t[13856] ^ n[13857];
assign t[13858] = t[13857] ^ n[13858];
assign t[13859] = t[13858] ^ n[13859];
assign t[13860] = t[13859] ^ n[13860];
assign t[13861] = t[13860] ^ n[13861];
assign t[13862] = t[13861] ^ n[13862];
assign t[13863] = t[13862] ^ n[13863];
assign t[13864] = t[13863] ^ n[13864];
assign t[13865] = t[13864] ^ n[13865];
assign t[13866] = t[13865] ^ n[13866];
assign t[13867] = t[13866] ^ n[13867];
assign t[13868] = t[13867] ^ n[13868];
assign t[13869] = t[13868] ^ n[13869];
assign t[13870] = t[13869] ^ n[13870];
assign t[13871] = t[13870] ^ n[13871];
assign t[13872] = t[13871] ^ n[13872];
assign t[13873] = t[13872] ^ n[13873];
assign t[13874] = t[13873] ^ n[13874];
assign t[13875] = t[13874] ^ n[13875];
assign t[13876] = t[13875] ^ n[13876];
assign t[13877] = t[13876] ^ n[13877];
assign t[13878] = t[13877] ^ n[13878];
assign t[13879] = t[13878] ^ n[13879];
assign t[13880] = t[13879] ^ n[13880];
assign t[13881] = t[13880] ^ n[13881];
assign t[13882] = t[13881] ^ n[13882];
assign t[13883] = t[13882] ^ n[13883];
assign t[13884] = t[13883] ^ n[13884];
assign t[13885] = t[13884] ^ n[13885];
assign t[13886] = t[13885] ^ n[13886];
assign t[13887] = t[13886] ^ n[13887];
assign t[13888] = t[13887] ^ n[13888];
assign t[13889] = t[13888] ^ n[13889];
assign t[13890] = t[13889] ^ n[13890];
assign t[13891] = t[13890] ^ n[13891];
assign t[13892] = t[13891] ^ n[13892];
assign t[13893] = t[13892] ^ n[13893];
assign t[13894] = t[13893] ^ n[13894];
assign t[13895] = t[13894] ^ n[13895];
assign t[13896] = t[13895] ^ n[13896];
assign t[13897] = t[13896] ^ n[13897];
assign t[13898] = t[13897] ^ n[13898];
assign t[13899] = t[13898] ^ n[13899];
assign t[13900] = t[13899] ^ n[13900];
assign t[13901] = t[13900] ^ n[13901];
assign t[13902] = t[13901] ^ n[13902];
assign t[13903] = t[13902] ^ n[13903];
assign t[13904] = t[13903] ^ n[13904];
assign t[13905] = t[13904] ^ n[13905];
assign t[13906] = t[13905] ^ n[13906];
assign t[13907] = t[13906] ^ n[13907];
assign t[13908] = t[13907] ^ n[13908];
assign t[13909] = t[13908] ^ n[13909];
assign t[13910] = t[13909] ^ n[13910];
assign t[13911] = t[13910] ^ n[13911];
assign t[13912] = t[13911] ^ n[13912];
assign t[13913] = t[13912] ^ n[13913];
assign t[13914] = t[13913] ^ n[13914];
assign t[13915] = t[13914] ^ n[13915];
assign t[13916] = t[13915] ^ n[13916];
assign t[13917] = t[13916] ^ n[13917];
assign t[13918] = t[13917] ^ n[13918];
assign t[13919] = t[13918] ^ n[13919];
assign t[13920] = t[13919] ^ n[13920];
assign t[13921] = t[13920] ^ n[13921];
assign t[13922] = t[13921] ^ n[13922];
assign t[13923] = t[13922] ^ n[13923];
assign t[13924] = t[13923] ^ n[13924];
assign t[13925] = t[13924] ^ n[13925];
assign t[13926] = t[13925] ^ n[13926];
assign t[13927] = t[13926] ^ n[13927];
assign t[13928] = t[13927] ^ n[13928];
assign t[13929] = t[13928] ^ n[13929];
assign t[13930] = t[13929] ^ n[13930];
assign t[13931] = t[13930] ^ n[13931];
assign t[13932] = t[13931] ^ n[13932];
assign t[13933] = t[13932] ^ n[13933];
assign t[13934] = t[13933] ^ n[13934];
assign t[13935] = t[13934] ^ n[13935];
assign t[13936] = t[13935] ^ n[13936];
assign t[13937] = t[13936] ^ n[13937];
assign t[13938] = t[13937] ^ n[13938];
assign t[13939] = t[13938] ^ n[13939];
assign t[13940] = t[13939] ^ n[13940];
assign t[13941] = t[13940] ^ n[13941];
assign t[13942] = t[13941] ^ n[13942];
assign t[13943] = t[13942] ^ n[13943];
assign t[13944] = t[13943] ^ n[13944];
assign t[13945] = t[13944] ^ n[13945];
assign t[13946] = t[13945] ^ n[13946];
assign t[13947] = t[13946] ^ n[13947];
assign t[13948] = t[13947] ^ n[13948];
assign t[13949] = t[13948] ^ n[13949];
assign t[13950] = t[13949] ^ n[13950];
assign t[13951] = t[13950] ^ n[13951];
assign t[13952] = t[13951] ^ n[13952];
assign t[13953] = t[13952] ^ n[13953];
assign t[13954] = t[13953] ^ n[13954];
assign t[13955] = t[13954] ^ n[13955];
assign t[13956] = t[13955] ^ n[13956];
assign t[13957] = t[13956] ^ n[13957];
assign t[13958] = t[13957] ^ n[13958];
assign t[13959] = t[13958] ^ n[13959];
assign t[13960] = t[13959] ^ n[13960];
assign t[13961] = t[13960] ^ n[13961];
assign t[13962] = t[13961] ^ n[13962];
assign t[13963] = t[13962] ^ n[13963];
assign t[13964] = t[13963] ^ n[13964];
assign t[13965] = t[13964] ^ n[13965];
assign t[13966] = t[13965] ^ n[13966];
assign t[13967] = t[13966] ^ n[13967];
assign t[13968] = t[13967] ^ n[13968];
assign t[13969] = t[13968] ^ n[13969];
assign t[13970] = t[13969] ^ n[13970];
assign t[13971] = t[13970] ^ n[13971];
assign t[13972] = t[13971] ^ n[13972];
assign t[13973] = t[13972] ^ n[13973];
assign t[13974] = t[13973] ^ n[13974];
assign t[13975] = t[13974] ^ n[13975];
assign t[13976] = t[13975] ^ n[13976];
assign t[13977] = t[13976] ^ n[13977];
assign t[13978] = t[13977] ^ n[13978];
assign t[13979] = t[13978] ^ n[13979];
assign t[13980] = t[13979] ^ n[13980];
assign t[13981] = t[13980] ^ n[13981];
assign t[13982] = t[13981] ^ n[13982];
assign t[13983] = t[13982] ^ n[13983];
assign t[13984] = t[13983] ^ n[13984];
assign t[13985] = t[13984] ^ n[13985];
assign t[13986] = t[13985] ^ n[13986];
assign t[13987] = t[13986] ^ n[13987];
assign t[13988] = t[13987] ^ n[13988];
assign t[13989] = t[13988] ^ n[13989];
assign t[13990] = t[13989] ^ n[13990];
assign t[13991] = t[13990] ^ n[13991];
assign t[13992] = t[13991] ^ n[13992];
assign t[13993] = t[13992] ^ n[13993];
assign t[13994] = t[13993] ^ n[13994];
assign t[13995] = t[13994] ^ n[13995];
assign t[13996] = t[13995] ^ n[13996];
assign t[13997] = t[13996] ^ n[13997];
assign t[13998] = t[13997] ^ n[13998];
assign t[13999] = t[13998] ^ n[13999];
assign t[14000] = t[13999] ^ n[14000];
assign t[14001] = t[14000] ^ n[14001];
assign t[14002] = t[14001] ^ n[14002];
assign t[14003] = t[14002] ^ n[14003];
assign t[14004] = t[14003] ^ n[14004];
assign t[14005] = t[14004] ^ n[14005];
assign t[14006] = t[14005] ^ n[14006];
assign t[14007] = t[14006] ^ n[14007];
assign t[14008] = t[14007] ^ n[14008];
assign t[14009] = t[14008] ^ n[14009];
assign t[14010] = t[14009] ^ n[14010];
assign t[14011] = t[14010] ^ n[14011];
assign t[14012] = t[14011] ^ n[14012];
assign t[14013] = t[14012] ^ n[14013];
assign t[14014] = t[14013] ^ n[14014];
assign t[14015] = t[14014] ^ n[14015];
assign t[14016] = t[14015] ^ n[14016];
assign t[14017] = t[14016] ^ n[14017];
assign t[14018] = t[14017] ^ n[14018];
assign t[14019] = t[14018] ^ n[14019];
assign t[14020] = t[14019] ^ n[14020];
assign t[14021] = t[14020] ^ n[14021];
assign t[14022] = t[14021] ^ n[14022];
assign t[14023] = t[14022] ^ n[14023];
assign t[14024] = t[14023] ^ n[14024];
assign t[14025] = t[14024] ^ n[14025];
assign t[14026] = t[14025] ^ n[14026];
assign t[14027] = t[14026] ^ n[14027];
assign t[14028] = t[14027] ^ n[14028];
assign t[14029] = t[14028] ^ n[14029];
assign t[14030] = t[14029] ^ n[14030];
assign t[14031] = t[14030] ^ n[14031];
assign t[14032] = t[14031] ^ n[14032];
assign t[14033] = t[14032] ^ n[14033];
assign t[14034] = t[14033] ^ n[14034];
assign t[14035] = t[14034] ^ n[14035];
assign t[14036] = t[14035] ^ n[14036];
assign t[14037] = t[14036] ^ n[14037];
assign t[14038] = t[14037] ^ n[14038];
assign t[14039] = t[14038] ^ n[14039];
assign t[14040] = t[14039] ^ n[14040];
assign t[14041] = t[14040] ^ n[14041];
assign t[14042] = t[14041] ^ n[14042];
assign t[14043] = t[14042] ^ n[14043];
assign t[14044] = t[14043] ^ n[14044];
assign t[14045] = t[14044] ^ n[14045];
assign t[14046] = t[14045] ^ n[14046];
assign t[14047] = t[14046] ^ n[14047];
assign t[14048] = t[14047] ^ n[14048];
assign t[14049] = t[14048] ^ n[14049];
assign t[14050] = t[14049] ^ n[14050];
assign t[14051] = t[14050] ^ n[14051];
assign t[14052] = t[14051] ^ n[14052];
assign t[14053] = t[14052] ^ n[14053];
assign t[14054] = t[14053] ^ n[14054];
assign t[14055] = t[14054] ^ n[14055];
assign t[14056] = t[14055] ^ n[14056];
assign t[14057] = t[14056] ^ n[14057];
assign t[14058] = t[14057] ^ n[14058];
assign t[14059] = t[14058] ^ n[14059];
assign t[14060] = t[14059] ^ n[14060];
assign t[14061] = t[14060] ^ n[14061];
assign t[14062] = t[14061] ^ n[14062];
assign t[14063] = t[14062] ^ n[14063];
assign t[14064] = t[14063] ^ n[14064];
assign t[14065] = t[14064] ^ n[14065];
assign t[14066] = t[14065] ^ n[14066];
assign t[14067] = t[14066] ^ n[14067];
assign t[14068] = t[14067] ^ n[14068];
assign t[14069] = t[14068] ^ n[14069];
assign t[14070] = t[14069] ^ n[14070];
assign t[14071] = t[14070] ^ n[14071];
assign t[14072] = t[14071] ^ n[14072];
assign t[14073] = t[14072] ^ n[14073];
assign t[14074] = t[14073] ^ n[14074];
assign t[14075] = t[14074] ^ n[14075];
assign t[14076] = t[14075] ^ n[14076];
assign t[14077] = t[14076] ^ n[14077];
assign t[14078] = t[14077] ^ n[14078];
assign t[14079] = t[14078] ^ n[14079];
assign t[14080] = t[14079] ^ n[14080];
assign t[14081] = t[14080] ^ n[14081];
assign t[14082] = t[14081] ^ n[14082];
assign t[14083] = t[14082] ^ n[14083];
assign t[14084] = t[14083] ^ n[14084];
assign t[14085] = t[14084] ^ n[14085];
assign t[14086] = t[14085] ^ n[14086];
assign t[14087] = t[14086] ^ n[14087];
assign t[14088] = t[14087] ^ n[14088];
assign t[14089] = t[14088] ^ n[14089];
assign t[14090] = t[14089] ^ n[14090];
assign t[14091] = t[14090] ^ n[14091];
assign t[14092] = t[14091] ^ n[14092];
assign t[14093] = t[14092] ^ n[14093];
assign t[14094] = t[14093] ^ n[14094];
assign t[14095] = t[14094] ^ n[14095];
assign t[14096] = t[14095] ^ n[14096];
assign t[14097] = t[14096] ^ n[14097];
assign t[14098] = t[14097] ^ n[14098];
assign t[14099] = t[14098] ^ n[14099];
assign t[14100] = t[14099] ^ n[14100];
assign t[14101] = t[14100] ^ n[14101];
assign t[14102] = t[14101] ^ n[14102];
assign t[14103] = t[14102] ^ n[14103];
assign t[14104] = t[14103] ^ n[14104];
assign t[14105] = t[14104] ^ n[14105];
assign t[14106] = t[14105] ^ n[14106];
assign t[14107] = t[14106] ^ n[14107];
assign t[14108] = t[14107] ^ n[14108];
assign t[14109] = t[14108] ^ n[14109];
assign t[14110] = t[14109] ^ n[14110];
assign t[14111] = t[14110] ^ n[14111];
assign t[14112] = t[14111] ^ n[14112];
assign t[14113] = t[14112] ^ n[14113];
assign t[14114] = t[14113] ^ n[14114];
assign t[14115] = t[14114] ^ n[14115];
assign t[14116] = t[14115] ^ n[14116];
assign t[14117] = t[14116] ^ n[14117];
assign t[14118] = t[14117] ^ n[14118];
assign t[14119] = t[14118] ^ n[14119];
assign t[14120] = t[14119] ^ n[14120];
assign t[14121] = t[14120] ^ n[14121];
assign t[14122] = t[14121] ^ n[14122];
assign t[14123] = t[14122] ^ n[14123];
assign t[14124] = t[14123] ^ n[14124];
assign t[14125] = t[14124] ^ n[14125];
assign t[14126] = t[14125] ^ n[14126];
assign t[14127] = t[14126] ^ n[14127];
assign t[14128] = t[14127] ^ n[14128];
assign t[14129] = t[14128] ^ n[14129];
assign t[14130] = t[14129] ^ n[14130];
assign t[14131] = t[14130] ^ n[14131];
assign t[14132] = t[14131] ^ n[14132];
assign t[14133] = t[14132] ^ n[14133];
assign t[14134] = t[14133] ^ n[14134];
assign t[14135] = t[14134] ^ n[14135];
assign t[14136] = t[14135] ^ n[14136];
assign t[14137] = t[14136] ^ n[14137];
assign t[14138] = t[14137] ^ n[14138];
assign t[14139] = t[14138] ^ n[14139];
assign t[14140] = t[14139] ^ n[14140];
assign t[14141] = t[14140] ^ n[14141];
assign t[14142] = t[14141] ^ n[14142];
assign t[14143] = t[14142] ^ n[14143];
assign t[14144] = t[14143] ^ n[14144];
assign t[14145] = t[14144] ^ n[14145];
assign t[14146] = t[14145] ^ n[14146];
assign t[14147] = t[14146] ^ n[14147];
assign t[14148] = t[14147] ^ n[14148];
assign t[14149] = t[14148] ^ n[14149];
assign t[14150] = t[14149] ^ n[14150];
assign t[14151] = t[14150] ^ n[14151];
assign t[14152] = t[14151] ^ n[14152];
assign t[14153] = t[14152] ^ n[14153];
assign t[14154] = t[14153] ^ n[14154];
assign t[14155] = t[14154] ^ n[14155];
assign t[14156] = t[14155] ^ n[14156];
assign t[14157] = t[14156] ^ n[14157];
assign t[14158] = t[14157] ^ n[14158];
assign t[14159] = t[14158] ^ n[14159];
assign t[14160] = t[14159] ^ n[14160];
assign t[14161] = t[14160] ^ n[14161];
assign t[14162] = t[14161] ^ n[14162];
assign t[14163] = t[14162] ^ n[14163];
assign t[14164] = t[14163] ^ n[14164];
assign t[14165] = t[14164] ^ n[14165];
assign t[14166] = t[14165] ^ n[14166];
assign t[14167] = t[14166] ^ n[14167];
assign t[14168] = t[14167] ^ n[14168];
assign t[14169] = t[14168] ^ n[14169];
assign t[14170] = t[14169] ^ n[14170];
assign t[14171] = t[14170] ^ n[14171];
assign t[14172] = t[14171] ^ n[14172];
assign t[14173] = t[14172] ^ n[14173];
assign t[14174] = t[14173] ^ n[14174];
assign t[14175] = t[14174] ^ n[14175];
assign t[14176] = t[14175] ^ n[14176];
assign t[14177] = t[14176] ^ n[14177];
assign t[14178] = t[14177] ^ n[14178];
assign t[14179] = t[14178] ^ n[14179];
assign t[14180] = t[14179] ^ n[14180];
assign t[14181] = t[14180] ^ n[14181];
assign t[14182] = t[14181] ^ n[14182];
assign t[14183] = t[14182] ^ n[14183];
assign t[14184] = t[14183] ^ n[14184];
assign t[14185] = t[14184] ^ n[14185];
assign t[14186] = t[14185] ^ n[14186];
assign t[14187] = t[14186] ^ n[14187];
assign t[14188] = t[14187] ^ n[14188];
assign t[14189] = t[14188] ^ n[14189];
assign t[14190] = t[14189] ^ n[14190];
assign t[14191] = t[14190] ^ n[14191];
assign t[14192] = t[14191] ^ n[14192];
assign t[14193] = t[14192] ^ n[14193];
assign t[14194] = t[14193] ^ n[14194];
assign t[14195] = t[14194] ^ n[14195];
assign t[14196] = t[14195] ^ n[14196];
assign t[14197] = t[14196] ^ n[14197];
assign t[14198] = t[14197] ^ n[14198];
assign t[14199] = t[14198] ^ n[14199];
assign t[14200] = t[14199] ^ n[14200];
assign t[14201] = t[14200] ^ n[14201];
assign t[14202] = t[14201] ^ n[14202];
assign t[14203] = t[14202] ^ n[14203];
assign t[14204] = t[14203] ^ n[14204];
assign t[14205] = t[14204] ^ n[14205];
assign t[14206] = t[14205] ^ n[14206];
assign t[14207] = t[14206] ^ n[14207];
assign t[14208] = t[14207] ^ n[14208];
assign t[14209] = t[14208] ^ n[14209];
assign t[14210] = t[14209] ^ n[14210];
assign t[14211] = t[14210] ^ n[14211];
assign t[14212] = t[14211] ^ n[14212];
assign t[14213] = t[14212] ^ n[14213];
assign t[14214] = t[14213] ^ n[14214];
assign t[14215] = t[14214] ^ n[14215];
assign t[14216] = t[14215] ^ n[14216];
assign t[14217] = t[14216] ^ n[14217];
assign t[14218] = t[14217] ^ n[14218];
assign t[14219] = t[14218] ^ n[14219];
assign t[14220] = t[14219] ^ n[14220];
assign t[14221] = t[14220] ^ n[14221];
assign t[14222] = t[14221] ^ n[14222];
assign t[14223] = t[14222] ^ n[14223];
assign t[14224] = t[14223] ^ n[14224];
assign t[14225] = t[14224] ^ n[14225];
assign t[14226] = t[14225] ^ n[14226];
assign t[14227] = t[14226] ^ n[14227];
assign t[14228] = t[14227] ^ n[14228];
assign t[14229] = t[14228] ^ n[14229];
assign t[14230] = t[14229] ^ n[14230];
assign t[14231] = t[14230] ^ n[14231];
assign t[14232] = t[14231] ^ n[14232];
assign t[14233] = t[14232] ^ n[14233];
assign t[14234] = t[14233] ^ n[14234];
assign t[14235] = t[14234] ^ n[14235];
assign t[14236] = t[14235] ^ n[14236];
assign t[14237] = t[14236] ^ n[14237];
assign t[14238] = t[14237] ^ n[14238];
assign t[14239] = t[14238] ^ n[14239];
assign t[14240] = t[14239] ^ n[14240];
assign t[14241] = t[14240] ^ n[14241];
assign t[14242] = t[14241] ^ n[14242];
assign t[14243] = t[14242] ^ n[14243];
assign t[14244] = t[14243] ^ n[14244];
assign t[14245] = t[14244] ^ n[14245];
assign t[14246] = t[14245] ^ n[14246];
assign t[14247] = t[14246] ^ n[14247];
assign t[14248] = t[14247] ^ n[14248];
assign t[14249] = t[14248] ^ n[14249];
assign t[14250] = t[14249] ^ n[14250];
assign t[14251] = t[14250] ^ n[14251];
assign t[14252] = t[14251] ^ n[14252];
assign t[14253] = t[14252] ^ n[14253];
assign t[14254] = t[14253] ^ n[14254];
assign t[14255] = t[14254] ^ n[14255];
assign t[14256] = t[14255] ^ n[14256];
assign t[14257] = t[14256] ^ n[14257];
assign t[14258] = t[14257] ^ n[14258];
assign t[14259] = t[14258] ^ n[14259];
assign t[14260] = t[14259] ^ n[14260];
assign t[14261] = t[14260] ^ n[14261];
assign t[14262] = t[14261] ^ n[14262];
assign t[14263] = t[14262] ^ n[14263];
assign t[14264] = t[14263] ^ n[14264];
assign t[14265] = t[14264] ^ n[14265];
assign t[14266] = t[14265] ^ n[14266];
assign t[14267] = t[14266] ^ n[14267];
assign t[14268] = t[14267] ^ n[14268];
assign t[14269] = t[14268] ^ n[14269];
assign t[14270] = t[14269] ^ n[14270];
assign t[14271] = t[14270] ^ n[14271];
assign t[14272] = t[14271] ^ n[14272];
assign t[14273] = t[14272] ^ n[14273];
assign t[14274] = t[14273] ^ n[14274];
assign t[14275] = t[14274] ^ n[14275];
assign t[14276] = t[14275] ^ n[14276];
assign t[14277] = t[14276] ^ n[14277];
assign t[14278] = t[14277] ^ n[14278];
assign t[14279] = t[14278] ^ n[14279];
assign t[14280] = t[14279] ^ n[14280];
assign t[14281] = t[14280] ^ n[14281];
assign t[14282] = t[14281] ^ n[14282];
assign t[14283] = t[14282] ^ n[14283];
assign t[14284] = t[14283] ^ n[14284];
assign t[14285] = t[14284] ^ n[14285];
assign t[14286] = t[14285] ^ n[14286];
assign t[14287] = t[14286] ^ n[14287];
assign t[14288] = t[14287] ^ n[14288];
assign t[14289] = t[14288] ^ n[14289];
assign t[14290] = t[14289] ^ n[14290];
assign t[14291] = t[14290] ^ n[14291];
assign t[14292] = t[14291] ^ n[14292];
assign t[14293] = t[14292] ^ n[14293];
assign t[14294] = t[14293] ^ n[14294];
assign t[14295] = t[14294] ^ n[14295];
assign t[14296] = t[14295] ^ n[14296];
assign t[14297] = t[14296] ^ n[14297];
assign t[14298] = t[14297] ^ n[14298];
assign t[14299] = t[14298] ^ n[14299];
assign t[14300] = t[14299] ^ n[14300];
assign t[14301] = t[14300] ^ n[14301];
assign t[14302] = t[14301] ^ n[14302];
assign t[14303] = t[14302] ^ n[14303];
assign t[14304] = t[14303] ^ n[14304];
assign t[14305] = t[14304] ^ n[14305];
assign t[14306] = t[14305] ^ n[14306];
assign t[14307] = t[14306] ^ n[14307];
assign t[14308] = t[14307] ^ n[14308];
assign t[14309] = t[14308] ^ n[14309];
assign t[14310] = t[14309] ^ n[14310];
assign t[14311] = t[14310] ^ n[14311];
assign t[14312] = t[14311] ^ n[14312];
assign t[14313] = t[14312] ^ n[14313];
assign t[14314] = t[14313] ^ n[14314];
assign t[14315] = t[14314] ^ n[14315];
assign t[14316] = t[14315] ^ n[14316];
assign t[14317] = t[14316] ^ n[14317];
assign t[14318] = t[14317] ^ n[14318];
assign t[14319] = t[14318] ^ n[14319];
assign t[14320] = t[14319] ^ n[14320];
assign t[14321] = t[14320] ^ n[14321];
assign t[14322] = t[14321] ^ n[14322];
assign t[14323] = t[14322] ^ n[14323];
assign t[14324] = t[14323] ^ n[14324];
assign t[14325] = t[14324] ^ n[14325];
assign t[14326] = t[14325] ^ n[14326];
assign t[14327] = t[14326] ^ n[14327];
assign t[14328] = t[14327] ^ n[14328];
assign t[14329] = t[14328] ^ n[14329];
assign t[14330] = t[14329] ^ n[14330];
assign t[14331] = t[14330] ^ n[14331];
assign t[14332] = t[14331] ^ n[14332];
assign t[14333] = t[14332] ^ n[14333];
assign t[14334] = t[14333] ^ n[14334];
assign t[14335] = t[14334] ^ n[14335];
assign t[14336] = t[14335] ^ n[14336];
assign t[14337] = t[14336] ^ n[14337];
assign t[14338] = t[14337] ^ n[14338];
assign t[14339] = t[14338] ^ n[14339];
assign t[14340] = t[14339] ^ n[14340];
assign t[14341] = t[14340] ^ n[14341];
assign t[14342] = t[14341] ^ n[14342];
assign t[14343] = t[14342] ^ n[14343];
assign t[14344] = t[14343] ^ n[14344];
assign t[14345] = t[14344] ^ n[14345];
assign t[14346] = t[14345] ^ n[14346];
assign t[14347] = t[14346] ^ n[14347];
assign t[14348] = t[14347] ^ n[14348];
assign t[14349] = t[14348] ^ n[14349];
assign t[14350] = t[14349] ^ n[14350];
assign t[14351] = t[14350] ^ n[14351];
assign t[14352] = t[14351] ^ n[14352];
assign t[14353] = t[14352] ^ n[14353];
assign t[14354] = t[14353] ^ n[14354];
assign t[14355] = t[14354] ^ n[14355];
assign t[14356] = t[14355] ^ n[14356];
assign t[14357] = t[14356] ^ n[14357];
assign t[14358] = t[14357] ^ n[14358];
assign t[14359] = t[14358] ^ n[14359];
assign t[14360] = t[14359] ^ n[14360];
assign t[14361] = t[14360] ^ n[14361];
assign t[14362] = t[14361] ^ n[14362];
assign t[14363] = t[14362] ^ n[14363];
assign t[14364] = t[14363] ^ n[14364];
assign t[14365] = t[14364] ^ n[14365];
assign t[14366] = t[14365] ^ n[14366];
assign t[14367] = t[14366] ^ n[14367];
assign t[14368] = t[14367] ^ n[14368];
assign t[14369] = t[14368] ^ n[14369];
assign t[14370] = t[14369] ^ n[14370];
assign t[14371] = t[14370] ^ n[14371];
assign t[14372] = t[14371] ^ n[14372];
assign t[14373] = t[14372] ^ n[14373];
assign t[14374] = t[14373] ^ n[14374];
assign t[14375] = t[14374] ^ n[14375];
assign t[14376] = t[14375] ^ n[14376];
assign t[14377] = t[14376] ^ n[14377];
assign t[14378] = t[14377] ^ n[14378];
assign t[14379] = t[14378] ^ n[14379];
assign t[14380] = t[14379] ^ n[14380];
assign t[14381] = t[14380] ^ n[14381];
assign t[14382] = t[14381] ^ n[14382];
assign t[14383] = t[14382] ^ n[14383];
assign t[14384] = t[14383] ^ n[14384];
assign t[14385] = t[14384] ^ n[14385];
assign t[14386] = t[14385] ^ n[14386];
assign t[14387] = t[14386] ^ n[14387];
assign t[14388] = t[14387] ^ n[14388];
assign t[14389] = t[14388] ^ n[14389];
assign t[14390] = t[14389] ^ n[14390];
assign t[14391] = t[14390] ^ n[14391];
assign t[14392] = t[14391] ^ n[14392];
assign t[14393] = t[14392] ^ n[14393];
assign t[14394] = t[14393] ^ n[14394];
assign t[14395] = t[14394] ^ n[14395];
assign t[14396] = t[14395] ^ n[14396];
assign t[14397] = t[14396] ^ n[14397];
assign t[14398] = t[14397] ^ n[14398];
assign t[14399] = t[14398] ^ n[14399];
assign t[14400] = t[14399] ^ n[14400];
assign t[14401] = t[14400] ^ n[14401];
assign t[14402] = t[14401] ^ n[14402];
assign t[14403] = t[14402] ^ n[14403];
assign t[14404] = t[14403] ^ n[14404];
assign t[14405] = t[14404] ^ n[14405];
assign t[14406] = t[14405] ^ n[14406];
assign t[14407] = t[14406] ^ n[14407];
assign t[14408] = t[14407] ^ n[14408];
assign t[14409] = t[14408] ^ n[14409];
assign t[14410] = t[14409] ^ n[14410];
assign t[14411] = t[14410] ^ n[14411];
assign t[14412] = t[14411] ^ n[14412];
assign t[14413] = t[14412] ^ n[14413];
assign t[14414] = t[14413] ^ n[14414];
assign t[14415] = t[14414] ^ n[14415];
assign t[14416] = t[14415] ^ n[14416];
assign t[14417] = t[14416] ^ n[14417];
assign t[14418] = t[14417] ^ n[14418];
assign t[14419] = t[14418] ^ n[14419];
assign t[14420] = t[14419] ^ n[14420];
assign t[14421] = t[14420] ^ n[14421];
assign t[14422] = t[14421] ^ n[14422];
assign t[14423] = t[14422] ^ n[14423];
assign t[14424] = t[14423] ^ n[14424];
assign t[14425] = t[14424] ^ n[14425];
assign t[14426] = t[14425] ^ n[14426];
assign t[14427] = t[14426] ^ n[14427];
assign t[14428] = t[14427] ^ n[14428];
assign t[14429] = t[14428] ^ n[14429];
assign t[14430] = t[14429] ^ n[14430];
assign t[14431] = t[14430] ^ n[14431];
assign t[14432] = t[14431] ^ n[14432];
assign t[14433] = t[14432] ^ n[14433];
assign t[14434] = t[14433] ^ n[14434];
assign t[14435] = t[14434] ^ n[14435];
assign t[14436] = t[14435] ^ n[14436];
assign t[14437] = t[14436] ^ n[14437];
assign t[14438] = t[14437] ^ n[14438];
assign t[14439] = t[14438] ^ n[14439];
assign t[14440] = t[14439] ^ n[14440];
assign t[14441] = t[14440] ^ n[14441];
assign t[14442] = t[14441] ^ n[14442];
assign t[14443] = t[14442] ^ n[14443];
assign t[14444] = t[14443] ^ n[14444];
assign t[14445] = t[14444] ^ n[14445];
assign t[14446] = t[14445] ^ n[14446];
assign t[14447] = t[14446] ^ n[14447];
assign t[14448] = t[14447] ^ n[14448];
assign t[14449] = t[14448] ^ n[14449];
assign t[14450] = t[14449] ^ n[14450];
assign t[14451] = t[14450] ^ n[14451];
assign t[14452] = t[14451] ^ n[14452];
assign t[14453] = t[14452] ^ n[14453];
assign t[14454] = t[14453] ^ n[14454];
assign t[14455] = t[14454] ^ n[14455];
assign t[14456] = t[14455] ^ n[14456];
assign t[14457] = t[14456] ^ n[14457];
assign t[14458] = t[14457] ^ n[14458];
assign t[14459] = t[14458] ^ n[14459];
assign t[14460] = t[14459] ^ n[14460];
assign t[14461] = t[14460] ^ n[14461];
assign t[14462] = t[14461] ^ n[14462];
assign t[14463] = t[14462] ^ n[14463];
assign t[14464] = t[14463] ^ n[14464];
assign t[14465] = t[14464] ^ n[14465];
assign t[14466] = t[14465] ^ n[14466];
assign t[14467] = t[14466] ^ n[14467];
assign t[14468] = t[14467] ^ n[14468];
assign t[14469] = t[14468] ^ n[14469];
assign t[14470] = t[14469] ^ n[14470];
assign t[14471] = t[14470] ^ n[14471];
assign t[14472] = t[14471] ^ n[14472];
assign t[14473] = t[14472] ^ n[14473];
assign t[14474] = t[14473] ^ n[14474];
assign t[14475] = t[14474] ^ n[14475];
assign t[14476] = t[14475] ^ n[14476];
assign t[14477] = t[14476] ^ n[14477];
assign t[14478] = t[14477] ^ n[14478];
assign t[14479] = t[14478] ^ n[14479];
assign t[14480] = t[14479] ^ n[14480];
assign t[14481] = t[14480] ^ n[14481];
assign t[14482] = t[14481] ^ n[14482];
assign t[14483] = t[14482] ^ n[14483];
assign t[14484] = t[14483] ^ n[14484];
assign t[14485] = t[14484] ^ n[14485];
assign t[14486] = t[14485] ^ n[14486];
assign t[14487] = t[14486] ^ n[14487];
assign t[14488] = t[14487] ^ n[14488];
assign t[14489] = t[14488] ^ n[14489];
assign t[14490] = t[14489] ^ n[14490];
assign t[14491] = t[14490] ^ n[14491];
assign t[14492] = t[14491] ^ n[14492];
assign t[14493] = t[14492] ^ n[14493];
assign t[14494] = t[14493] ^ n[14494];
assign t[14495] = t[14494] ^ n[14495];
assign t[14496] = t[14495] ^ n[14496];
assign t[14497] = t[14496] ^ n[14497];
assign t[14498] = t[14497] ^ n[14498];
assign t[14499] = t[14498] ^ n[14499];
assign t[14500] = t[14499] ^ n[14500];
assign t[14501] = t[14500] ^ n[14501];
assign t[14502] = t[14501] ^ n[14502];
assign t[14503] = t[14502] ^ n[14503];
assign t[14504] = t[14503] ^ n[14504];
assign t[14505] = t[14504] ^ n[14505];
assign t[14506] = t[14505] ^ n[14506];
assign t[14507] = t[14506] ^ n[14507];
assign t[14508] = t[14507] ^ n[14508];
assign t[14509] = t[14508] ^ n[14509];
assign t[14510] = t[14509] ^ n[14510];
assign t[14511] = t[14510] ^ n[14511];
assign t[14512] = t[14511] ^ n[14512];
assign t[14513] = t[14512] ^ n[14513];
assign t[14514] = t[14513] ^ n[14514];
assign t[14515] = t[14514] ^ n[14515];
assign t[14516] = t[14515] ^ n[14516];
assign t[14517] = t[14516] ^ n[14517];
assign t[14518] = t[14517] ^ n[14518];
assign t[14519] = t[14518] ^ n[14519];
assign t[14520] = t[14519] ^ n[14520];
assign t[14521] = t[14520] ^ n[14521];
assign t[14522] = t[14521] ^ n[14522];
assign t[14523] = t[14522] ^ n[14523];
assign t[14524] = t[14523] ^ n[14524];
assign t[14525] = t[14524] ^ n[14525];
assign t[14526] = t[14525] ^ n[14526];
assign t[14527] = t[14526] ^ n[14527];
assign t[14528] = t[14527] ^ n[14528];
assign t[14529] = t[14528] ^ n[14529];
assign t[14530] = t[14529] ^ n[14530];
assign t[14531] = t[14530] ^ n[14531];
assign t[14532] = t[14531] ^ n[14532];
assign t[14533] = t[14532] ^ n[14533];
assign t[14534] = t[14533] ^ n[14534];
assign t[14535] = t[14534] ^ n[14535];
assign t[14536] = t[14535] ^ n[14536];
assign t[14537] = t[14536] ^ n[14537];
assign t[14538] = t[14537] ^ n[14538];
assign t[14539] = t[14538] ^ n[14539];
assign t[14540] = t[14539] ^ n[14540];
assign t[14541] = t[14540] ^ n[14541];
assign t[14542] = t[14541] ^ n[14542];
assign t[14543] = t[14542] ^ n[14543];
assign t[14544] = t[14543] ^ n[14544];
assign t[14545] = t[14544] ^ n[14545];
assign t[14546] = t[14545] ^ n[14546];
assign t[14547] = t[14546] ^ n[14547];
assign t[14548] = t[14547] ^ n[14548];
assign t[14549] = t[14548] ^ n[14549];
assign t[14550] = t[14549] ^ n[14550];
assign t[14551] = t[14550] ^ n[14551];
assign t[14552] = t[14551] ^ n[14552];
assign t[14553] = t[14552] ^ n[14553];
assign t[14554] = t[14553] ^ n[14554];
assign t[14555] = t[14554] ^ n[14555];
assign t[14556] = t[14555] ^ n[14556];
assign t[14557] = t[14556] ^ n[14557];
assign t[14558] = t[14557] ^ n[14558];
assign t[14559] = t[14558] ^ n[14559];
assign t[14560] = t[14559] ^ n[14560];
assign t[14561] = t[14560] ^ n[14561];
assign t[14562] = t[14561] ^ n[14562];
assign t[14563] = t[14562] ^ n[14563];
assign t[14564] = t[14563] ^ n[14564];
assign t[14565] = t[14564] ^ n[14565];
assign t[14566] = t[14565] ^ n[14566];
assign t[14567] = t[14566] ^ n[14567];
assign t[14568] = t[14567] ^ n[14568];
assign t[14569] = t[14568] ^ n[14569];
assign t[14570] = t[14569] ^ n[14570];
assign t[14571] = t[14570] ^ n[14571];
assign t[14572] = t[14571] ^ n[14572];
assign t[14573] = t[14572] ^ n[14573];
assign t[14574] = t[14573] ^ n[14574];
assign t[14575] = t[14574] ^ n[14575];
assign t[14576] = t[14575] ^ n[14576];
assign t[14577] = t[14576] ^ n[14577];
assign t[14578] = t[14577] ^ n[14578];
assign t[14579] = t[14578] ^ n[14579];
assign t[14580] = t[14579] ^ n[14580];
assign t[14581] = t[14580] ^ n[14581];
assign t[14582] = t[14581] ^ n[14582];
assign t[14583] = t[14582] ^ n[14583];
assign t[14584] = t[14583] ^ n[14584];
assign t[14585] = t[14584] ^ n[14585];
assign t[14586] = t[14585] ^ n[14586];
assign t[14587] = t[14586] ^ n[14587];
assign t[14588] = t[14587] ^ n[14588];
assign t[14589] = t[14588] ^ n[14589];
assign t[14590] = t[14589] ^ n[14590];
assign t[14591] = t[14590] ^ n[14591];
assign t[14592] = t[14591] ^ n[14592];
assign t[14593] = t[14592] ^ n[14593];
assign t[14594] = t[14593] ^ n[14594];
assign t[14595] = t[14594] ^ n[14595];
assign t[14596] = t[14595] ^ n[14596];
assign t[14597] = t[14596] ^ n[14597];
assign t[14598] = t[14597] ^ n[14598];
assign t[14599] = t[14598] ^ n[14599];
assign t[14600] = t[14599] ^ n[14600];
assign t[14601] = t[14600] ^ n[14601];
assign t[14602] = t[14601] ^ n[14602];
assign t[14603] = t[14602] ^ n[14603];
assign t[14604] = t[14603] ^ n[14604];
assign t[14605] = t[14604] ^ n[14605];
assign t[14606] = t[14605] ^ n[14606];
assign t[14607] = t[14606] ^ n[14607];
assign t[14608] = t[14607] ^ n[14608];
assign t[14609] = t[14608] ^ n[14609];
assign t[14610] = t[14609] ^ n[14610];
assign t[14611] = t[14610] ^ n[14611];
assign t[14612] = t[14611] ^ n[14612];
assign t[14613] = t[14612] ^ n[14613];
assign t[14614] = t[14613] ^ n[14614];
assign t[14615] = t[14614] ^ n[14615];
assign t[14616] = t[14615] ^ n[14616];
assign t[14617] = t[14616] ^ n[14617];
assign t[14618] = t[14617] ^ n[14618];
assign t[14619] = t[14618] ^ n[14619];
assign t[14620] = t[14619] ^ n[14620];
assign t[14621] = t[14620] ^ n[14621];
assign t[14622] = t[14621] ^ n[14622];
assign t[14623] = t[14622] ^ n[14623];
assign t[14624] = t[14623] ^ n[14624];
assign t[14625] = t[14624] ^ n[14625];
assign t[14626] = t[14625] ^ n[14626];
assign t[14627] = t[14626] ^ n[14627];
assign t[14628] = t[14627] ^ n[14628];
assign t[14629] = t[14628] ^ n[14629];
assign t[14630] = t[14629] ^ n[14630];
assign t[14631] = t[14630] ^ n[14631];
assign t[14632] = t[14631] ^ n[14632];
assign t[14633] = t[14632] ^ n[14633];
assign t[14634] = t[14633] ^ n[14634];
assign t[14635] = t[14634] ^ n[14635];
assign t[14636] = t[14635] ^ n[14636];
assign t[14637] = t[14636] ^ n[14637];
assign t[14638] = t[14637] ^ n[14638];
assign t[14639] = t[14638] ^ n[14639];
assign t[14640] = t[14639] ^ n[14640];
assign t[14641] = t[14640] ^ n[14641];
assign t[14642] = t[14641] ^ n[14642];
assign t[14643] = t[14642] ^ n[14643];
assign t[14644] = t[14643] ^ n[14644];
assign t[14645] = t[14644] ^ n[14645];
assign t[14646] = t[14645] ^ n[14646];
assign t[14647] = t[14646] ^ n[14647];
assign t[14648] = t[14647] ^ n[14648];
assign t[14649] = t[14648] ^ n[14649];
assign t[14650] = t[14649] ^ n[14650];
assign t[14651] = t[14650] ^ n[14651];
assign t[14652] = t[14651] ^ n[14652];
assign t[14653] = t[14652] ^ n[14653];
assign t[14654] = t[14653] ^ n[14654];
assign t[14655] = t[14654] ^ n[14655];
assign t[14656] = t[14655] ^ n[14656];
assign t[14657] = t[14656] ^ n[14657];
assign t[14658] = t[14657] ^ n[14658];
assign t[14659] = t[14658] ^ n[14659];
assign t[14660] = t[14659] ^ n[14660];
assign t[14661] = t[14660] ^ n[14661];
assign t[14662] = t[14661] ^ n[14662];
assign t[14663] = t[14662] ^ n[14663];
assign t[14664] = t[14663] ^ n[14664];
assign t[14665] = t[14664] ^ n[14665];
assign t[14666] = t[14665] ^ n[14666];
assign t[14667] = t[14666] ^ n[14667];
assign t[14668] = t[14667] ^ n[14668];
assign t[14669] = t[14668] ^ n[14669];
assign t[14670] = t[14669] ^ n[14670];
assign t[14671] = t[14670] ^ n[14671];
assign t[14672] = t[14671] ^ n[14672];
assign t[14673] = t[14672] ^ n[14673];
assign t[14674] = t[14673] ^ n[14674];
assign t[14675] = t[14674] ^ n[14675];
assign t[14676] = t[14675] ^ n[14676];
assign t[14677] = t[14676] ^ n[14677];
assign t[14678] = t[14677] ^ n[14678];
assign t[14679] = t[14678] ^ n[14679];
assign t[14680] = t[14679] ^ n[14680];
assign t[14681] = t[14680] ^ n[14681];
assign t[14682] = t[14681] ^ n[14682];
assign t[14683] = t[14682] ^ n[14683];
assign t[14684] = t[14683] ^ n[14684];
assign t[14685] = t[14684] ^ n[14685];
assign t[14686] = t[14685] ^ n[14686];
assign t[14687] = t[14686] ^ n[14687];
assign t[14688] = t[14687] ^ n[14688];
assign t[14689] = t[14688] ^ n[14689];
assign t[14690] = t[14689] ^ n[14690];
assign t[14691] = t[14690] ^ n[14691];
assign t[14692] = t[14691] ^ n[14692];
assign t[14693] = t[14692] ^ n[14693];
assign t[14694] = t[14693] ^ n[14694];
assign t[14695] = t[14694] ^ n[14695];
assign t[14696] = t[14695] ^ n[14696];
assign t[14697] = t[14696] ^ n[14697];
assign t[14698] = t[14697] ^ n[14698];
assign t[14699] = t[14698] ^ n[14699];
assign t[14700] = t[14699] ^ n[14700];
assign t[14701] = t[14700] ^ n[14701];
assign t[14702] = t[14701] ^ n[14702];
assign t[14703] = t[14702] ^ n[14703];
assign t[14704] = t[14703] ^ n[14704];
assign t[14705] = t[14704] ^ n[14705];
assign t[14706] = t[14705] ^ n[14706];
assign t[14707] = t[14706] ^ n[14707];
assign t[14708] = t[14707] ^ n[14708];
assign t[14709] = t[14708] ^ n[14709];
assign t[14710] = t[14709] ^ n[14710];
assign t[14711] = t[14710] ^ n[14711];
assign t[14712] = t[14711] ^ n[14712];
assign t[14713] = t[14712] ^ n[14713];
assign t[14714] = t[14713] ^ n[14714];
assign t[14715] = t[14714] ^ n[14715];
assign t[14716] = t[14715] ^ n[14716];
assign t[14717] = t[14716] ^ n[14717];
assign t[14718] = t[14717] ^ n[14718];
assign t[14719] = t[14718] ^ n[14719];
assign t[14720] = t[14719] ^ n[14720];
assign t[14721] = t[14720] ^ n[14721];
assign t[14722] = t[14721] ^ n[14722];
assign t[14723] = t[14722] ^ n[14723];
assign t[14724] = t[14723] ^ n[14724];
assign t[14725] = t[14724] ^ n[14725];
assign t[14726] = t[14725] ^ n[14726];
assign t[14727] = t[14726] ^ n[14727];
assign t[14728] = t[14727] ^ n[14728];
assign t[14729] = t[14728] ^ n[14729];
assign t[14730] = t[14729] ^ n[14730];
assign t[14731] = t[14730] ^ n[14731];
assign t[14732] = t[14731] ^ n[14732];
assign t[14733] = t[14732] ^ n[14733];
assign t[14734] = t[14733] ^ n[14734];
assign t[14735] = t[14734] ^ n[14735];
assign t[14736] = t[14735] ^ n[14736];
assign t[14737] = t[14736] ^ n[14737];
assign t[14738] = t[14737] ^ n[14738];
assign t[14739] = t[14738] ^ n[14739];
assign t[14740] = t[14739] ^ n[14740];
assign t[14741] = t[14740] ^ n[14741];
assign t[14742] = t[14741] ^ n[14742];
assign t[14743] = t[14742] ^ n[14743];
assign t[14744] = t[14743] ^ n[14744];
assign t[14745] = t[14744] ^ n[14745];
assign t[14746] = t[14745] ^ n[14746];
assign t[14747] = t[14746] ^ n[14747];
assign t[14748] = t[14747] ^ n[14748];
assign t[14749] = t[14748] ^ n[14749];
assign t[14750] = t[14749] ^ n[14750];
assign t[14751] = t[14750] ^ n[14751];
assign t[14752] = t[14751] ^ n[14752];
assign t[14753] = t[14752] ^ n[14753];
assign t[14754] = t[14753] ^ n[14754];
assign t[14755] = t[14754] ^ n[14755];
assign t[14756] = t[14755] ^ n[14756];
assign t[14757] = t[14756] ^ n[14757];
assign t[14758] = t[14757] ^ n[14758];
assign t[14759] = t[14758] ^ n[14759];
assign t[14760] = t[14759] ^ n[14760];
assign t[14761] = t[14760] ^ n[14761];
assign t[14762] = t[14761] ^ n[14762];
assign t[14763] = t[14762] ^ n[14763];
assign t[14764] = t[14763] ^ n[14764];
assign t[14765] = t[14764] ^ n[14765];
assign t[14766] = t[14765] ^ n[14766];
assign t[14767] = t[14766] ^ n[14767];
assign t[14768] = t[14767] ^ n[14768];
assign t[14769] = t[14768] ^ n[14769];
assign t[14770] = t[14769] ^ n[14770];
assign t[14771] = t[14770] ^ n[14771];
assign t[14772] = t[14771] ^ n[14772];
assign t[14773] = t[14772] ^ n[14773];
assign t[14774] = t[14773] ^ n[14774];
assign t[14775] = t[14774] ^ n[14775];
assign t[14776] = t[14775] ^ n[14776];
assign t[14777] = t[14776] ^ n[14777];
assign t[14778] = t[14777] ^ n[14778];
assign t[14779] = t[14778] ^ n[14779];
assign t[14780] = t[14779] ^ n[14780];
assign t[14781] = t[14780] ^ n[14781];
assign t[14782] = t[14781] ^ n[14782];
assign t[14783] = t[14782] ^ n[14783];
assign t[14784] = t[14783] ^ n[14784];
assign t[14785] = t[14784] ^ n[14785];
assign t[14786] = t[14785] ^ n[14786];
assign t[14787] = t[14786] ^ n[14787];
assign t[14788] = t[14787] ^ n[14788];
assign t[14789] = t[14788] ^ n[14789];
assign t[14790] = t[14789] ^ n[14790];
assign t[14791] = t[14790] ^ n[14791];
assign t[14792] = t[14791] ^ n[14792];
assign t[14793] = t[14792] ^ n[14793];
assign t[14794] = t[14793] ^ n[14794];
assign t[14795] = t[14794] ^ n[14795];
assign t[14796] = t[14795] ^ n[14796];
assign t[14797] = t[14796] ^ n[14797];
assign t[14798] = t[14797] ^ n[14798];
assign t[14799] = t[14798] ^ n[14799];
assign t[14800] = t[14799] ^ n[14800];
assign t[14801] = t[14800] ^ n[14801];
assign t[14802] = t[14801] ^ n[14802];
assign t[14803] = t[14802] ^ n[14803];
assign t[14804] = t[14803] ^ n[14804];
assign t[14805] = t[14804] ^ n[14805];
assign t[14806] = t[14805] ^ n[14806];
assign t[14807] = t[14806] ^ n[14807];
assign t[14808] = t[14807] ^ n[14808];
assign t[14809] = t[14808] ^ n[14809];
assign t[14810] = t[14809] ^ n[14810];
assign t[14811] = t[14810] ^ n[14811];
assign t[14812] = t[14811] ^ n[14812];
assign t[14813] = t[14812] ^ n[14813];
assign t[14814] = t[14813] ^ n[14814];
assign t[14815] = t[14814] ^ n[14815];
assign t[14816] = t[14815] ^ n[14816];
assign t[14817] = t[14816] ^ n[14817];
assign t[14818] = t[14817] ^ n[14818];
assign t[14819] = t[14818] ^ n[14819];
assign t[14820] = t[14819] ^ n[14820];
assign t[14821] = t[14820] ^ n[14821];
assign t[14822] = t[14821] ^ n[14822];
assign t[14823] = t[14822] ^ n[14823];
assign t[14824] = t[14823] ^ n[14824];
assign t[14825] = t[14824] ^ n[14825];
assign t[14826] = t[14825] ^ n[14826];
assign t[14827] = t[14826] ^ n[14827];
assign t[14828] = t[14827] ^ n[14828];
assign t[14829] = t[14828] ^ n[14829];
assign t[14830] = t[14829] ^ n[14830];
assign t[14831] = t[14830] ^ n[14831];
assign t[14832] = t[14831] ^ n[14832];
assign t[14833] = t[14832] ^ n[14833];
assign t[14834] = t[14833] ^ n[14834];
assign t[14835] = t[14834] ^ n[14835];
assign t[14836] = t[14835] ^ n[14836];
assign t[14837] = t[14836] ^ n[14837];
assign t[14838] = t[14837] ^ n[14838];
assign t[14839] = t[14838] ^ n[14839];
assign t[14840] = t[14839] ^ n[14840];
assign t[14841] = t[14840] ^ n[14841];
assign t[14842] = t[14841] ^ n[14842];
assign t[14843] = t[14842] ^ n[14843];
assign t[14844] = t[14843] ^ n[14844];
assign t[14845] = t[14844] ^ n[14845];
assign t[14846] = t[14845] ^ n[14846];
assign t[14847] = t[14846] ^ n[14847];
assign t[14848] = t[14847] ^ n[14848];
assign t[14849] = t[14848] ^ n[14849];
assign t[14850] = t[14849] ^ n[14850];
assign t[14851] = t[14850] ^ n[14851];
assign t[14852] = t[14851] ^ n[14852];
assign t[14853] = t[14852] ^ n[14853];
assign t[14854] = t[14853] ^ n[14854];
assign t[14855] = t[14854] ^ n[14855];
assign t[14856] = t[14855] ^ n[14856];
assign t[14857] = t[14856] ^ n[14857];
assign t[14858] = t[14857] ^ n[14858];
assign t[14859] = t[14858] ^ n[14859];
assign t[14860] = t[14859] ^ n[14860];
assign t[14861] = t[14860] ^ n[14861];
assign t[14862] = t[14861] ^ n[14862];
assign t[14863] = t[14862] ^ n[14863];
assign t[14864] = t[14863] ^ n[14864];
assign t[14865] = t[14864] ^ n[14865];
assign t[14866] = t[14865] ^ n[14866];
assign t[14867] = t[14866] ^ n[14867];
assign t[14868] = t[14867] ^ n[14868];
assign t[14869] = t[14868] ^ n[14869];
assign t[14870] = t[14869] ^ n[14870];
assign t[14871] = t[14870] ^ n[14871];
assign t[14872] = t[14871] ^ n[14872];
assign t[14873] = t[14872] ^ n[14873];
assign t[14874] = t[14873] ^ n[14874];
assign t[14875] = t[14874] ^ n[14875];
assign t[14876] = t[14875] ^ n[14876];
assign t[14877] = t[14876] ^ n[14877];
assign t[14878] = t[14877] ^ n[14878];
assign t[14879] = t[14878] ^ n[14879];
assign t[14880] = t[14879] ^ n[14880];
assign t[14881] = t[14880] ^ n[14881];
assign t[14882] = t[14881] ^ n[14882];
assign t[14883] = t[14882] ^ n[14883];
assign t[14884] = t[14883] ^ n[14884];
assign t[14885] = t[14884] ^ n[14885];
assign t[14886] = t[14885] ^ n[14886];
assign t[14887] = t[14886] ^ n[14887];
assign t[14888] = t[14887] ^ n[14888];
assign t[14889] = t[14888] ^ n[14889];
assign t[14890] = t[14889] ^ n[14890];
assign t[14891] = t[14890] ^ n[14891];
assign t[14892] = t[14891] ^ n[14892];
assign t[14893] = t[14892] ^ n[14893];
assign t[14894] = t[14893] ^ n[14894];
assign t[14895] = t[14894] ^ n[14895];
assign t[14896] = t[14895] ^ n[14896];
assign t[14897] = t[14896] ^ n[14897];
assign t[14898] = t[14897] ^ n[14898];
assign t[14899] = t[14898] ^ n[14899];
assign t[14900] = t[14899] ^ n[14900];
assign t[14901] = t[14900] ^ n[14901];
assign t[14902] = t[14901] ^ n[14902];
assign t[14903] = t[14902] ^ n[14903];
assign t[14904] = t[14903] ^ n[14904];
assign t[14905] = t[14904] ^ n[14905];
assign t[14906] = t[14905] ^ n[14906];
assign t[14907] = t[14906] ^ n[14907];
assign t[14908] = t[14907] ^ n[14908];
assign t[14909] = t[14908] ^ n[14909];
assign t[14910] = t[14909] ^ n[14910];
assign t[14911] = t[14910] ^ n[14911];
assign t[14912] = t[14911] ^ n[14912];
assign t[14913] = t[14912] ^ n[14913];
assign t[14914] = t[14913] ^ n[14914];
assign t[14915] = t[14914] ^ n[14915];
assign t[14916] = t[14915] ^ n[14916];
assign t[14917] = t[14916] ^ n[14917];
assign t[14918] = t[14917] ^ n[14918];
assign t[14919] = t[14918] ^ n[14919];
assign t[14920] = t[14919] ^ n[14920];
assign t[14921] = t[14920] ^ n[14921];
assign t[14922] = t[14921] ^ n[14922];
assign t[14923] = t[14922] ^ n[14923];
assign t[14924] = t[14923] ^ n[14924];
assign t[14925] = t[14924] ^ n[14925];
assign t[14926] = t[14925] ^ n[14926];
assign t[14927] = t[14926] ^ n[14927];
assign t[14928] = t[14927] ^ n[14928];
assign t[14929] = t[14928] ^ n[14929];
assign t[14930] = t[14929] ^ n[14930];
assign t[14931] = t[14930] ^ n[14931];
assign t[14932] = t[14931] ^ n[14932];
assign t[14933] = t[14932] ^ n[14933];
assign t[14934] = t[14933] ^ n[14934];
assign t[14935] = t[14934] ^ n[14935];
assign t[14936] = t[14935] ^ n[14936];
assign t[14937] = t[14936] ^ n[14937];
assign t[14938] = t[14937] ^ n[14938];
assign t[14939] = t[14938] ^ n[14939];
assign t[14940] = t[14939] ^ n[14940];
assign t[14941] = t[14940] ^ n[14941];
assign t[14942] = t[14941] ^ n[14942];
assign t[14943] = t[14942] ^ n[14943];
assign t[14944] = t[14943] ^ n[14944];
assign t[14945] = t[14944] ^ n[14945];
assign t[14946] = t[14945] ^ n[14946];
assign t[14947] = t[14946] ^ n[14947];
assign t[14948] = t[14947] ^ n[14948];
assign t[14949] = t[14948] ^ n[14949];
assign t[14950] = t[14949] ^ n[14950];
assign t[14951] = t[14950] ^ n[14951];
assign t[14952] = t[14951] ^ n[14952];
assign t[14953] = t[14952] ^ n[14953];
assign t[14954] = t[14953] ^ n[14954];
assign t[14955] = t[14954] ^ n[14955];
assign t[14956] = t[14955] ^ n[14956];
assign t[14957] = t[14956] ^ n[14957];
assign t[14958] = t[14957] ^ n[14958];
assign t[14959] = t[14958] ^ n[14959];
assign t[14960] = t[14959] ^ n[14960];
assign t[14961] = t[14960] ^ n[14961];
assign t[14962] = t[14961] ^ n[14962];
assign t[14963] = t[14962] ^ n[14963];
assign t[14964] = t[14963] ^ n[14964];
assign t[14965] = t[14964] ^ n[14965];
assign t[14966] = t[14965] ^ n[14966];
assign t[14967] = t[14966] ^ n[14967];
assign t[14968] = t[14967] ^ n[14968];
assign t[14969] = t[14968] ^ n[14969];
assign t[14970] = t[14969] ^ n[14970];
assign t[14971] = t[14970] ^ n[14971];
assign t[14972] = t[14971] ^ n[14972];
assign t[14973] = t[14972] ^ n[14973];
assign t[14974] = t[14973] ^ n[14974];
assign t[14975] = t[14974] ^ n[14975];
assign t[14976] = t[14975] ^ n[14976];
assign t[14977] = t[14976] ^ n[14977];
assign t[14978] = t[14977] ^ n[14978];
assign t[14979] = t[14978] ^ n[14979];
assign t[14980] = t[14979] ^ n[14980];
assign t[14981] = t[14980] ^ n[14981];
assign t[14982] = t[14981] ^ n[14982];
assign t[14983] = t[14982] ^ n[14983];
assign t[14984] = t[14983] ^ n[14984];
assign t[14985] = t[14984] ^ n[14985];
assign t[14986] = t[14985] ^ n[14986];
assign t[14987] = t[14986] ^ n[14987];
assign t[14988] = t[14987] ^ n[14988];
assign t[14989] = t[14988] ^ n[14989];
assign t[14990] = t[14989] ^ n[14990];
assign t[14991] = t[14990] ^ n[14991];
assign t[14992] = t[14991] ^ n[14992];
assign t[14993] = t[14992] ^ n[14993];
assign t[14994] = t[14993] ^ n[14994];
assign t[14995] = t[14994] ^ n[14995];
assign t[14996] = t[14995] ^ n[14996];
assign t[14997] = t[14996] ^ n[14997];
assign t[14998] = t[14997] ^ n[14998];
assign t[14999] = t[14998] ^ n[14999];
assign t[15000] = t[14999] ^ n[15000];
assign t[15001] = t[15000] ^ n[15001];
assign t[15002] = t[15001] ^ n[15002];
assign t[15003] = t[15002] ^ n[15003];
assign t[15004] = t[15003] ^ n[15004];
assign t[15005] = t[15004] ^ n[15005];
assign t[15006] = t[15005] ^ n[15006];
assign t[15007] = t[15006] ^ n[15007];
assign t[15008] = t[15007] ^ n[15008];
assign t[15009] = t[15008] ^ n[15009];
assign t[15010] = t[15009] ^ n[15010];
assign t[15011] = t[15010] ^ n[15011];
assign t[15012] = t[15011] ^ n[15012];
assign t[15013] = t[15012] ^ n[15013];
assign t[15014] = t[15013] ^ n[15014];
assign t[15015] = t[15014] ^ n[15015];
assign t[15016] = t[15015] ^ n[15016];
assign t[15017] = t[15016] ^ n[15017];
assign t[15018] = t[15017] ^ n[15018];
assign t[15019] = t[15018] ^ n[15019];
assign t[15020] = t[15019] ^ n[15020];
assign t[15021] = t[15020] ^ n[15021];
assign t[15022] = t[15021] ^ n[15022];
assign t[15023] = t[15022] ^ n[15023];
assign t[15024] = t[15023] ^ n[15024];
assign t[15025] = t[15024] ^ n[15025];
assign t[15026] = t[15025] ^ n[15026];
assign t[15027] = t[15026] ^ n[15027];
assign t[15028] = t[15027] ^ n[15028];
assign t[15029] = t[15028] ^ n[15029];
assign t[15030] = t[15029] ^ n[15030];
assign t[15031] = t[15030] ^ n[15031];
assign t[15032] = t[15031] ^ n[15032];
assign t[15033] = t[15032] ^ n[15033];
assign t[15034] = t[15033] ^ n[15034];
assign t[15035] = t[15034] ^ n[15035];
assign t[15036] = t[15035] ^ n[15036];
assign t[15037] = t[15036] ^ n[15037];
assign t[15038] = t[15037] ^ n[15038];
assign t[15039] = t[15038] ^ n[15039];
assign t[15040] = t[15039] ^ n[15040];
assign t[15041] = t[15040] ^ n[15041];
assign t[15042] = t[15041] ^ n[15042];
assign t[15043] = t[15042] ^ n[15043];
assign t[15044] = t[15043] ^ n[15044];
assign t[15045] = t[15044] ^ n[15045];
assign t[15046] = t[15045] ^ n[15046];
assign t[15047] = t[15046] ^ n[15047];
assign t[15048] = t[15047] ^ n[15048];
assign t[15049] = t[15048] ^ n[15049];
assign t[15050] = t[15049] ^ n[15050];
assign t[15051] = t[15050] ^ n[15051];
assign t[15052] = t[15051] ^ n[15052];
assign t[15053] = t[15052] ^ n[15053];
assign t[15054] = t[15053] ^ n[15054];
assign t[15055] = t[15054] ^ n[15055];
assign t[15056] = t[15055] ^ n[15056];
assign t[15057] = t[15056] ^ n[15057];
assign t[15058] = t[15057] ^ n[15058];
assign t[15059] = t[15058] ^ n[15059];
assign t[15060] = t[15059] ^ n[15060];
assign t[15061] = t[15060] ^ n[15061];
assign t[15062] = t[15061] ^ n[15062];
assign t[15063] = t[15062] ^ n[15063];
assign t[15064] = t[15063] ^ n[15064];
assign t[15065] = t[15064] ^ n[15065];
assign t[15066] = t[15065] ^ n[15066];
assign t[15067] = t[15066] ^ n[15067];
assign t[15068] = t[15067] ^ n[15068];
assign t[15069] = t[15068] ^ n[15069];
assign t[15070] = t[15069] ^ n[15070];
assign t[15071] = t[15070] ^ n[15071];
assign t[15072] = t[15071] ^ n[15072];
assign t[15073] = t[15072] ^ n[15073];
assign t[15074] = t[15073] ^ n[15074];
assign t[15075] = t[15074] ^ n[15075];
assign t[15076] = t[15075] ^ n[15076];
assign t[15077] = t[15076] ^ n[15077];
assign t[15078] = t[15077] ^ n[15078];
assign t[15079] = t[15078] ^ n[15079];
assign t[15080] = t[15079] ^ n[15080];
assign t[15081] = t[15080] ^ n[15081];
assign t[15082] = t[15081] ^ n[15082];
assign t[15083] = t[15082] ^ n[15083];
assign t[15084] = t[15083] ^ n[15084];
assign t[15085] = t[15084] ^ n[15085];
assign t[15086] = t[15085] ^ n[15086];
assign t[15087] = t[15086] ^ n[15087];
assign t[15088] = t[15087] ^ n[15088];
assign t[15089] = t[15088] ^ n[15089];
assign t[15090] = t[15089] ^ n[15090];
assign t[15091] = t[15090] ^ n[15091];
assign t[15092] = t[15091] ^ n[15092];
assign t[15093] = t[15092] ^ n[15093];
assign t[15094] = t[15093] ^ n[15094];
assign t[15095] = t[15094] ^ n[15095];
assign t[15096] = t[15095] ^ n[15096];
assign t[15097] = t[15096] ^ n[15097];
assign t[15098] = t[15097] ^ n[15098];
assign t[15099] = t[15098] ^ n[15099];
assign t[15100] = t[15099] ^ n[15100];
assign t[15101] = t[15100] ^ n[15101];
assign t[15102] = t[15101] ^ n[15102];
assign t[15103] = t[15102] ^ n[15103];
assign t[15104] = t[15103] ^ n[15104];
assign t[15105] = t[15104] ^ n[15105];
assign t[15106] = t[15105] ^ n[15106];
assign t[15107] = t[15106] ^ n[15107];
assign t[15108] = t[15107] ^ n[15108];
assign t[15109] = t[15108] ^ n[15109];
assign t[15110] = t[15109] ^ n[15110];
assign t[15111] = t[15110] ^ n[15111];
assign t[15112] = t[15111] ^ n[15112];
assign t[15113] = t[15112] ^ n[15113];
assign t[15114] = t[15113] ^ n[15114];
assign t[15115] = t[15114] ^ n[15115];
assign t[15116] = t[15115] ^ n[15116];
assign t[15117] = t[15116] ^ n[15117];
assign t[15118] = t[15117] ^ n[15118];
assign t[15119] = t[15118] ^ n[15119];
assign t[15120] = t[15119] ^ n[15120];
assign t[15121] = t[15120] ^ n[15121];
assign t[15122] = t[15121] ^ n[15122];
assign t[15123] = t[15122] ^ n[15123];
assign t[15124] = t[15123] ^ n[15124];
assign t[15125] = t[15124] ^ n[15125];
assign t[15126] = t[15125] ^ n[15126];
assign t[15127] = t[15126] ^ n[15127];
assign t[15128] = t[15127] ^ n[15128];
assign t[15129] = t[15128] ^ n[15129];
assign t[15130] = t[15129] ^ n[15130];
assign t[15131] = t[15130] ^ n[15131];
assign t[15132] = t[15131] ^ n[15132];
assign t[15133] = t[15132] ^ n[15133];
assign t[15134] = t[15133] ^ n[15134];
assign t[15135] = t[15134] ^ n[15135];
assign t[15136] = t[15135] ^ n[15136];
assign t[15137] = t[15136] ^ n[15137];
assign t[15138] = t[15137] ^ n[15138];
assign t[15139] = t[15138] ^ n[15139];
assign t[15140] = t[15139] ^ n[15140];
assign t[15141] = t[15140] ^ n[15141];
assign t[15142] = t[15141] ^ n[15142];
assign t[15143] = t[15142] ^ n[15143];
assign t[15144] = t[15143] ^ n[15144];
assign t[15145] = t[15144] ^ n[15145];
assign t[15146] = t[15145] ^ n[15146];
assign t[15147] = t[15146] ^ n[15147];
assign t[15148] = t[15147] ^ n[15148];
assign t[15149] = t[15148] ^ n[15149];
assign t[15150] = t[15149] ^ n[15150];
assign t[15151] = t[15150] ^ n[15151];
assign t[15152] = t[15151] ^ n[15152];
assign t[15153] = t[15152] ^ n[15153];
assign t[15154] = t[15153] ^ n[15154];
assign t[15155] = t[15154] ^ n[15155];
assign t[15156] = t[15155] ^ n[15156];
assign t[15157] = t[15156] ^ n[15157];
assign t[15158] = t[15157] ^ n[15158];
assign t[15159] = t[15158] ^ n[15159];
assign t[15160] = t[15159] ^ n[15160];
assign t[15161] = t[15160] ^ n[15161];
assign t[15162] = t[15161] ^ n[15162];
assign t[15163] = t[15162] ^ n[15163];
assign t[15164] = t[15163] ^ n[15164];
assign t[15165] = t[15164] ^ n[15165];
assign t[15166] = t[15165] ^ n[15166];
assign t[15167] = t[15166] ^ n[15167];
assign t[15168] = t[15167] ^ n[15168];
assign t[15169] = t[15168] ^ n[15169];
assign t[15170] = t[15169] ^ n[15170];
assign t[15171] = t[15170] ^ n[15171];
assign t[15172] = t[15171] ^ n[15172];
assign t[15173] = t[15172] ^ n[15173];
assign t[15174] = t[15173] ^ n[15174];
assign t[15175] = t[15174] ^ n[15175];
assign t[15176] = t[15175] ^ n[15176];
assign t[15177] = t[15176] ^ n[15177];
assign t[15178] = t[15177] ^ n[15178];
assign t[15179] = t[15178] ^ n[15179];
assign t[15180] = t[15179] ^ n[15180];
assign t[15181] = t[15180] ^ n[15181];
assign t[15182] = t[15181] ^ n[15182];
assign t[15183] = t[15182] ^ n[15183];
assign t[15184] = t[15183] ^ n[15184];
assign t[15185] = t[15184] ^ n[15185];
assign t[15186] = t[15185] ^ n[15186];
assign t[15187] = t[15186] ^ n[15187];
assign t[15188] = t[15187] ^ n[15188];
assign t[15189] = t[15188] ^ n[15189];
assign t[15190] = t[15189] ^ n[15190];
assign t[15191] = t[15190] ^ n[15191];
assign t[15192] = t[15191] ^ n[15192];
assign t[15193] = t[15192] ^ n[15193];
assign t[15194] = t[15193] ^ n[15194];
assign t[15195] = t[15194] ^ n[15195];
assign t[15196] = t[15195] ^ n[15196];
assign t[15197] = t[15196] ^ n[15197];
assign t[15198] = t[15197] ^ n[15198];
assign t[15199] = t[15198] ^ n[15199];
assign t[15200] = t[15199] ^ n[15200];
assign t[15201] = t[15200] ^ n[15201];
assign t[15202] = t[15201] ^ n[15202];
assign t[15203] = t[15202] ^ n[15203];
assign t[15204] = t[15203] ^ n[15204];
assign t[15205] = t[15204] ^ n[15205];
assign t[15206] = t[15205] ^ n[15206];
assign t[15207] = t[15206] ^ n[15207];
assign t[15208] = t[15207] ^ n[15208];
assign t[15209] = t[15208] ^ n[15209];
assign t[15210] = t[15209] ^ n[15210];
assign t[15211] = t[15210] ^ n[15211];
assign t[15212] = t[15211] ^ n[15212];
assign t[15213] = t[15212] ^ n[15213];
assign t[15214] = t[15213] ^ n[15214];
assign t[15215] = t[15214] ^ n[15215];
assign t[15216] = t[15215] ^ n[15216];
assign t[15217] = t[15216] ^ n[15217];
assign t[15218] = t[15217] ^ n[15218];
assign t[15219] = t[15218] ^ n[15219];
assign t[15220] = t[15219] ^ n[15220];
assign t[15221] = t[15220] ^ n[15221];
assign t[15222] = t[15221] ^ n[15222];
assign t[15223] = t[15222] ^ n[15223];
assign t[15224] = t[15223] ^ n[15224];
assign t[15225] = t[15224] ^ n[15225];
assign t[15226] = t[15225] ^ n[15226];
assign t[15227] = t[15226] ^ n[15227];
assign t[15228] = t[15227] ^ n[15228];
assign t[15229] = t[15228] ^ n[15229];
assign t[15230] = t[15229] ^ n[15230];
assign t[15231] = t[15230] ^ n[15231];
assign t[15232] = t[15231] ^ n[15232];
assign t[15233] = t[15232] ^ n[15233];
assign t[15234] = t[15233] ^ n[15234];
assign t[15235] = t[15234] ^ n[15235];
assign t[15236] = t[15235] ^ n[15236];
assign t[15237] = t[15236] ^ n[15237];
assign t[15238] = t[15237] ^ n[15238];
assign t[15239] = t[15238] ^ n[15239];
assign t[15240] = t[15239] ^ n[15240];
assign t[15241] = t[15240] ^ n[15241];
assign t[15242] = t[15241] ^ n[15242];
assign t[15243] = t[15242] ^ n[15243];
assign t[15244] = t[15243] ^ n[15244];
assign t[15245] = t[15244] ^ n[15245];
assign t[15246] = t[15245] ^ n[15246];
assign t[15247] = t[15246] ^ n[15247];
assign t[15248] = t[15247] ^ n[15248];
assign t[15249] = t[15248] ^ n[15249];
assign t[15250] = t[15249] ^ n[15250];
assign t[15251] = t[15250] ^ n[15251];
assign t[15252] = t[15251] ^ n[15252];
assign t[15253] = t[15252] ^ n[15253];
assign t[15254] = t[15253] ^ n[15254];
assign t[15255] = t[15254] ^ n[15255];
assign t[15256] = t[15255] ^ n[15256];
assign t[15257] = t[15256] ^ n[15257];
assign t[15258] = t[15257] ^ n[15258];
assign t[15259] = t[15258] ^ n[15259];
assign t[15260] = t[15259] ^ n[15260];
assign t[15261] = t[15260] ^ n[15261];
assign t[15262] = t[15261] ^ n[15262];
assign t[15263] = t[15262] ^ n[15263];
assign t[15264] = t[15263] ^ n[15264];
assign t[15265] = t[15264] ^ n[15265];
assign t[15266] = t[15265] ^ n[15266];
assign t[15267] = t[15266] ^ n[15267];
assign t[15268] = t[15267] ^ n[15268];
assign t[15269] = t[15268] ^ n[15269];
assign t[15270] = t[15269] ^ n[15270];
assign t[15271] = t[15270] ^ n[15271];
assign t[15272] = t[15271] ^ n[15272];
assign t[15273] = t[15272] ^ n[15273];
assign t[15274] = t[15273] ^ n[15274];
assign t[15275] = t[15274] ^ n[15275];
assign t[15276] = t[15275] ^ n[15276];
assign t[15277] = t[15276] ^ n[15277];
assign t[15278] = t[15277] ^ n[15278];
assign t[15279] = t[15278] ^ n[15279];
assign t[15280] = t[15279] ^ n[15280];
assign t[15281] = t[15280] ^ n[15281];
assign t[15282] = t[15281] ^ n[15282];
assign t[15283] = t[15282] ^ n[15283];
assign t[15284] = t[15283] ^ n[15284];
assign t[15285] = t[15284] ^ n[15285];
assign t[15286] = t[15285] ^ n[15286];
assign t[15287] = t[15286] ^ n[15287];
assign t[15288] = t[15287] ^ n[15288];
assign t[15289] = t[15288] ^ n[15289];
assign t[15290] = t[15289] ^ n[15290];
assign t[15291] = t[15290] ^ n[15291];
assign t[15292] = t[15291] ^ n[15292];
assign t[15293] = t[15292] ^ n[15293];
assign t[15294] = t[15293] ^ n[15294];
assign t[15295] = t[15294] ^ n[15295];
assign t[15296] = t[15295] ^ n[15296];
assign t[15297] = t[15296] ^ n[15297];
assign t[15298] = t[15297] ^ n[15298];
assign t[15299] = t[15298] ^ n[15299];
assign t[15300] = t[15299] ^ n[15300];
assign t[15301] = t[15300] ^ n[15301];
assign t[15302] = t[15301] ^ n[15302];
assign t[15303] = t[15302] ^ n[15303];
assign t[15304] = t[15303] ^ n[15304];
assign t[15305] = t[15304] ^ n[15305];
assign t[15306] = t[15305] ^ n[15306];
assign t[15307] = t[15306] ^ n[15307];
assign t[15308] = t[15307] ^ n[15308];
assign t[15309] = t[15308] ^ n[15309];
assign t[15310] = t[15309] ^ n[15310];
assign t[15311] = t[15310] ^ n[15311];
assign t[15312] = t[15311] ^ n[15312];
assign t[15313] = t[15312] ^ n[15313];
assign t[15314] = t[15313] ^ n[15314];
assign t[15315] = t[15314] ^ n[15315];
assign t[15316] = t[15315] ^ n[15316];
assign t[15317] = t[15316] ^ n[15317];
assign t[15318] = t[15317] ^ n[15318];
assign t[15319] = t[15318] ^ n[15319];
assign t[15320] = t[15319] ^ n[15320];
assign t[15321] = t[15320] ^ n[15321];
assign t[15322] = t[15321] ^ n[15322];
assign t[15323] = t[15322] ^ n[15323];
assign t[15324] = t[15323] ^ n[15324];
assign t[15325] = t[15324] ^ n[15325];
assign t[15326] = t[15325] ^ n[15326];
assign t[15327] = t[15326] ^ n[15327];
assign t[15328] = t[15327] ^ n[15328];
assign t[15329] = t[15328] ^ n[15329];
assign t[15330] = t[15329] ^ n[15330];
assign t[15331] = t[15330] ^ n[15331];
assign t[15332] = t[15331] ^ n[15332];
assign t[15333] = t[15332] ^ n[15333];
assign t[15334] = t[15333] ^ n[15334];
assign t[15335] = t[15334] ^ n[15335];
assign t[15336] = t[15335] ^ n[15336];
assign t[15337] = t[15336] ^ n[15337];
assign t[15338] = t[15337] ^ n[15338];
assign t[15339] = t[15338] ^ n[15339];
assign t[15340] = t[15339] ^ n[15340];
assign t[15341] = t[15340] ^ n[15341];
assign t[15342] = t[15341] ^ n[15342];
assign t[15343] = t[15342] ^ n[15343];
assign t[15344] = t[15343] ^ n[15344];
assign t[15345] = t[15344] ^ n[15345];
assign t[15346] = t[15345] ^ n[15346];
assign t[15347] = t[15346] ^ n[15347];
assign t[15348] = t[15347] ^ n[15348];
assign t[15349] = t[15348] ^ n[15349];
assign t[15350] = t[15349] ^ n[15350];
assign t[15351] = t[15350] ^ n[15351];
assign t[15352] = t[15351] ^ n[15352];
assign t[15353] = t[15352] ^ n[15353];
assign t[15354] = t[15353] ^ n[15354];
assign t[15355] = t[15354] ^ n[15355];
assign t[15356] = t[15355] ^ n[15356];
assign t[15357] = t[15356] ^ n[15357];
assign t[15358] = t[15357] ^ n[15358];
assign t[15359] = t[15358] ^ n[15359];
assign t[15360] = t[15359] ^ n[15360];
assign t[15361] = t[15360] ^ n[15361];
assign t[15362] = t[15361] ^ n[15362];
assign t[15363] = t[15362] ^ n[15363];
assign t[15364] = t[15363] ^ n[15364];
assign t[15365] = t[15364] ^ n[15365];
assign t[15366] = t[15365] ^ n[15366];
assign t[15367] = t[15366] ^ n[15367];
assign t[15368] = t[15367] ^ n[15368];
assign t[15369] = t[15368] ^ n[15369];
assign t[15370] = t[15369] ^ n[15370];
assign t[15371] = t[15370] ^ n[15371];
assign t[15372] = t[15371] ^ n[15372];
assign t[15373] = t[15372] ^ n[15373];
assign t[15374] = t[15373] ^ n[15374];
assign t[15375] = t[15374] ^ n[15375];
assign t[15376] = t[15375] ^ n[15376];
assign t[15377] = t[15376] ^ n[15377];
assign t[15378] = t[15377] ^ n[15378];
assign t[15379] = t[15378] ^ n[15379];
assign t[15380] = t[15379] ^ n[15380];
assign t[15381] = t[15380] ^ n[15381];
assign t[15382] = t[15381] ^ n[15382];
assign t[15383] = t[15382] ^ n[15383];
assign t[15384] = t[15383] ^ n[15384];
assign t[15385] = t[15384] ^ n[15385];
assign t[15386] = t[15385] ^ n[15386];
assign t[15387] = t[15386] ^ n[15387];
assign t[15388] = t[15387] ^ n[15388];
assign t[15389] = t[15388] ^ n[15389];
assign t[15390] = t[15389] ^ n[15390];
assign t[15391] = t[15390] ^ n[15391];
assign t[15392] = t[15391] ^ n[15392];
assign t[15393] = t[15392] ^ n[15393];
assign t[15394] = t[15393] ^ n[15394];
assign t[15395] = t[15394] ^ n[15395];
assign t[15396] = t[15395] ^ n[15396];
assign t[15397] = t[15396] ^ n[15397];
assign t[15398] = t[15397] ^ n[15398];
assign t[15399] = t[15398] ^ n[15399];
assign t[15400] = t[15399] ^ n[15400];
assign t[15401] = t[15400] ^ n[15401];
assign t[15402] = t[15401] ^ n[15402];
assign t[15403] = t[15402] ^ n[15403];
assign t[15404] = t[15403] ^ n[15404];
assign t[15405] = t[15404] ^ n[15405];
assign t[15406] = t[15405] ^ n[15406];
assign t[15407] = t[15406] ^ n[15407];
assign t[15408] = t[15407] ^ n[15408];
assign t[15409] = t[15408] ^ n[15409];
assign t[15410] = t[15409] ^ n[15410];
assign t[15411] = t[15410] ^ n[15411];
assign t[15412] = t[15411] ^ n[15412];
assign t[15413] = t[15412] ^ n[15413];
assign t[15414] = t[15413] ^ n[15414];
assign t[15415] = t[15414] ^ n[15415];
assign t[15416] = t[15415] ^ n[15416];
assign t[15417] = t[15416] ^ n[15417];
assign t[15418] = t[15417] ^ n[15418];
assign t[15419] = t[15418] ^ n[15419];
assign t[15420] = t[15419] ^ n[15420];
assign t[15421] = t[15420] ^ n[15421];
assign t[15422] = t[15421] ^ n[15422];
assign t[15423] = t[15422] ^ n[15423];
assign t[15424] = t[15423] ^ n[15424];
assign t[15425] = t[15424] ^ n[15425];
assign t[15426] = t[15425] ^ n[15426];
assign t[15427] = t[15426] ^ n[15427];
assign t[15428] = t[15427] ^ n[15428];
assign t[15429] = t[15428] ^ n[15429];
assign t[15430] = t[15429] ^ n[15430];
assign t[15431] = t[15430] ^ n[15431];
assign t[15432] = t[15431] ^ n[15432];
assign t[15433] = t[15432] ^ n[15433];
assign t[15434] = t[15433] ^ n[15434];
assign t[15435] = t[15434] ^ n[15435];
assign t[15436] = t[15435] ^ n[15436];
assign t[15437] = t[15436] ^ n[15437];
assign t[15438] = t[15437] ^ n[15438];
assign t[15439] = t[15438] ^ n[15439];
assign t[15440] = t[15439] ^ n[15440];
assign t[15441] = t[15440] ^ n[15441];
assign t[15442] = t[15441] ^ n[15442];
assign t[15443] = t[15442] ^ n[15443];
assign t[15444] = t[15443] ^ n[15444];
assign t[15445] = t[15444] ^ n[15445];
assign t[15446] = t[15445] ^ n[15446];
assign t[15447] = t[15446] ^ n[15447];
assign t[15448] = t[15447] ^ n[15448];
assign t[15449] = t[15448] ^ n[15449];
assign t[15450] = t[15449] ^ n[15450];
assign t[15451] = t[15450] ^ n[15451];
assign t[15452] = t[15451] ^ n[15452];
assign t[15453] = t[15452] ^ n[15453];
assign t[15454] = t[15453] ^ n[15454];
assign t[15455] = t[15454] ^ n[15455];
assign t[15456] = t[15455] ^ n[15456];
assign t[15457] = t[15456] ^ n[15457];
assign t[15458] = t[15457] ^ n[15458];
assign t[15459] = t[15458] ^ n[15459];
assign t[15460] = t[15459] ^ n[15460];
assign t[15461] = t[15460] ^ n[15461];
assign t[15462] = t[15461] ^ n[15462];
assign t[15463] = t[15462] ^ n[15463];
assign t[15464] = t[15463] ^ n[15464];
assign t[15465] = t[15464] ^ n[15465];
assign t[15466] = t[15465] ^ n[15466];
assign t[15467] = t[15466] ^ n[15467];
assign t[15468] = t[15467] ^ n[15468];
assign t[15469] = t[15468] ^ n[15469];
assign t[15470] = t[15469] ^ n[15470];
assign t[15471] = t[15470] ^ n[15471];
assign t[15472] = t[15471] ^ n[15472];
assign t[15473] = t[15472] ^ n[15473];
assign t[15474] = t[15473] ^ n[15474];
assign t[15475] = t[15474] ^ n[15475];
assign t[15476] = t[15475] ^ n[15476];
assign t[15477] = t[15476] ^ n[15477];
assign t[15478] = t[15477] ^ n[15478];
assign t[15479] = t[15478] ^ n[15479];
assign t[15480] = t[15479] ^ n[15480];
assign t[15481] = t[15480] ^ n[15481];
assign t[15482] = t[15481] ^ n[15482];
assign t[15483] = t[15482] ^ n[15483];
assign t[15484] = t[15483] ^ n[15484];
assign t[15485] = t[15484] ^ n[15485];
assign t[15486] = t[15485] ^ n[15486];
assign t[15487] = t[15486] ^ n[15487];
assign t[15488] = t[15487] ^ n[15488];
assign t[15489] = t[15488] ^ n[15489];
assign t[15490] = t[15489] ^ n[15490];
assign t[15491] = t[15490] ^ n[15491];
assign t[15492] = t[15491] ^ n[15492];
assign t[15493] = t[15492] ^ n[15493];
assign t[15494] = t[15493] ^ n[15494];
assign t[15495] = t[15494] ^ n[15495];
assign t[15496] = t[15495] ^ n[15496];
assign t[15497] = t[15496] ^ n[15497];
assign t[15498] = t[15497] ^ n[15498];
assign t[15499] = t[15498] ^ n[15499];
assign t[15500] = t[15499] ^ n[15500];
assign t[15501] = t[15500] ^ n[15501];
assign t[15502] = t[15501] ^ n[15502];
assign t[15503] = t[15502] ^ n[15503];
assign t[15504] = t[15503] ^ n[15504];
assign t[15505] = t[15504] ^ n[15505];
assign t[15506] = t[15505] ^ n[15506];
assign t[15507] = t[15506] ^ n[15507];
assign t[15508] = t[15507] ^ n[15508];
assign t[15509] = t[15508] ^ n[15509];
assign t[15510] = t[15509] ^ n[15510];
assign t[15511] = t[15510] ^ n[15511];
assign t[15512] = t[15511] ^ n[15512];
assign t[15513] = t[15512] ^ n[15513];
assign t[15514] = t[15513] ^ n[15514];
assign t[15515] = t[15514] ^ n[15515];
assign t[15516] = t[15515] ^ n[15516];
assign t[15517] = t[15516] ^ n[15517];
assign t[15518] = t[15517] ^ n[15518];
assign t[15519] = t[15518] ^ n[15519];
assign t[15520] = t[15519] ^ n[15520];
assign t[15521] = t[15520] ^ n[15521];
assign t[15522] = t[15521] ^ n[15522];
assign t[15523] = t[15522] ^ n[15523];
assign t[15524] = t[15523] ^ n[15524];
assign t[15525] = t[15524] ^ n[15525];
assign t[15526] = t[15525] ^ n[15526];
assign t[15527] = t[15526] ^ n[15527];
assign t[15528] = t[15527] ^ n[15528];
assign t[15529] = t[15528] ^ n[15529];
assign t[15530] = t[15529] ^ n[15530];
assign t[15531] = t[15530] ^ n[15531];
assign t[15532] = t[15531] ^ n[15532];
assign t[15533] = t[15532] ^ n[15533];
assign t[15534] = t[15533] ^ n[15534];
assign t[15535] = t[15534] ^ n[15535];
assign t[15536] = t[15535] ^ n[15536];
assign t[15537] = t[15536] ^ n[15537];
assign t[15538] = t[15537] ^ n[15538];
assign t[15539] = t[15538] ^ n[15539];
assign t[15540] = t[15539] ^ n[15540];
assign t[15541] = t[15540] ^ n[15541];
assign t[15542] = t[15541] ^ n[15542];
assign t[15543] = t[15542] ^ n[15543];
assign t[15544] = t[15543] ^ n[15544];
assign t[15545] = t[15544] ^ n[15545];
assign t[15546] = t[15545] ^ n[15546];
assign t[15547] = t[15546] ^ n[15547];
assign t[15548] = t[15547] ^ n[15548];
assign t[15549] = t[15548] ^ n[15549];
assign t[15550] = t[15549] ^ n[15550];
assign t[15551] = t[15550] ^ n[15551];
assign t[15552] = t[15551] ^ n[15552];
assign t[15553] = t[15552] ^ n[15553];
assign t[15554] = t[15553] ^ n[15554];
assign t[15555] = t[15554] ^ n[15555];
assign t[15556] = t[15555] ^ n[15556];
assign t[15557] = t[15556] ^ n[15557];
assign t[15558] = t[15557] ^ n[15558];
assign t[15559] = t[15558] ^ n[15559];
assign t[15560] = t[15559] ^ n[15560];
assign t[15561] = t[15560] ^ n[15561];
assign t[15562] = t[15561] ^ n[15562];
assign t[15563] = t[15562] ^ n[15563];
assign t[15564] = t[15563] ^ n[15564];
assign t[15565] = t[15564] ^ n[15565];
assign t[15566] = t[15565] ^ n[15566];
assign t[15567] = t[15566] ^ n[15567];
assign t[15568] = t[15567] ^ n[15568];
assign t[15569] = t[15568] ^ n[15569];
assign t[15570] = t[15569] ^ n[15570];
assign t[15571] = t[15570] ^ n[15571];
assign t[15572] = t[15571] ^ n[15572];
assign t[15573] = t[15572] ^ n[15573];
assign t[15574] = t[15573] ^ n[15574];
assign t[15575] = t[15574] ^ n[15575];
assign t[15576] = t[15575] ^ n[15576];
assign t[15577] = t[15576] ^ n[15577];
assign t[15578] = t[15577] ^ n[15578];
assign t[15579] = t[15578] ^ n[15579];
assign t[15580] = t[15579] ^ n[15580];
assign t[15581] = t[15580] ^ n[15581];
assign t[15582] = t[15581] ^ n[15582];
assign t[15583] = t[15582] ^ n[15583];
assign t[15584] = t[15583] ^ n[15584];
assign t[15585] = t[15584] ^ n[15585];
assign t[15586] = t[15585] ^ n[15586];
assign t[15587] = t[15586] ^ n[15587];
assign t[15588] = t[15587] ^ n[15588];
assign t[15589] = t[15588] ^ n[15589];
assign t[15590] = t[15589] ^ n[15590];
assign t[15591] = t[15590] ^ n[15591];
assign t[15592] = t[15591] ^ n[15592];
assign t[15593] = t[15592] ^ n[15593];
assign t[15594] = t[15593] ^ n[15594];
assign t[15595] = t[15594] ^ n[15595];
assign t[15596] = t[15595] ^ n[15596];
assign t[15597] = t[15596] ^ n[15597];
assign t[15598] = t[15597] ^ n[15598];
assign t[15599] = t[15598] ^ n[15599];
assign t[15600] = t[15599] ^ n[15600];
assign t[15601] = t[15600] ^ n[15601];
assign t[15602] = t[15601] ^ n[15602];
assign t[15603] = t[15602] ^ n[15603];
assign t[15604] = t[15603] ^ n[15604];
assign t[15605] = t[15604] ^ n[15605];
assign t[15606] = t[15605] ^ n[15606];
assign t[15607] = t[15606] ^ n[15607];
assign t[15608] = t[15607] ^ n[15608];
assign t[15609] = t[15608] ^ n[15609];
assign t[15610] = t[15609] ^ n[15610];
assign t[15611] = t[15610] ^ n[15611];
assign t[15612] = t[15611] ^ n[15612];
assign t[15613] = t[15612] ^ n[15613];
assign t[15614] = t[15613] ^ n[15614];
assign t[15615] = t[15614] ^ n[15615];
assign t[15616] = t[15615] ^ n[15616];
assign t[15617] = t[15616] ^ n[15617];
assign t[15618] = t[15617] ^ n[15618];
assign t[15619] = t[15618] ^ n[15619];
assign t[15620] = t[15619] ^ n[15620];
assign t[15621] = t[15620] ^ n[15621];
assign t[15622] = t[15621] ^ n[15622];
assign t[15623] = t[15622] ^ n[15623];
assign t[15624] = t[15623] ^ n[15624];
assign t[15625] = t[15624] ^ n[15625];
assign t[15626] = t[15625] ^ n[15626];
assign t[15627] = t[15626] ^ n[15627];
assign t[15628] = t[15627] ^ n[15628];
assign t[15629] = t[15628] ^ n[15629];
assign t[15630] = t[15629] ^ n[15630];
assign t[15631] = t[15630] ^ n[15631];
assign t[15632] = t[15631] ^ n[15632];
assign t[15633] = t[15632] ^ n[15633];
assign t[15634] = t[15633] ^ n[15634];
assign t[15635] = t[15634] ^ n[15635];
assign t[15636] = t[15635] ^ n[15636];
assign t[15637] = t[15636] ^ n[15637];
assign t[15638] = t[15637] ^ n[15638];
assign t[15639] = t[15638] ^ n[15639];
assign t[15640] = t[15639] ^ n[15640];
assign t[15641] = t[15640] ^ n[15641];
assign t[15642] = t[15641] ^ n[15642];
assign t[15643] = t[15642] ^ n[15643];
assign t[15644] = t[15643] ^ n[15644];
assign t[15645] = t[15644] ^ n[15645];
assign t[15646] = t[15645] ^ n[15646];
assign t[15647] = t[15646] ^ n[15647];
assign t[15648] = t[15647] ^ n[15648];
assign t[15649] = t[15648] ^ n[15649];
assign t[15650] = t[15649] ^ n[15650];
assign t[15651] = t[15650] ^ n[15651];
assign t[15652] = t[15651] ^ n[15652];
assign t[15653] = t[15652] ^ n[15653];
assign t[15654] = t[15653] ^ n[15654];
assign t[15655] = t[15654] ^ n[15655];
assign t[15656] = t[15655] ^ n[15656];
assign t[15657] = t[15656] ^ n[15657];
assign t[15658] = t[15657] ^ n[15658];
assign t[15659] = t[15658] ^ n[15659];
assign t[15660] = t[15659] ^ n[15660];
assign t[15661] = t[15660] ^ n[15661];
assign t[15662] = t[15661] ^ n[15662];
assign t[15663] = t[15662] ^ n[15663];
assign t[15664] = t[15663] ^ n[15664];
assign t[15665] = t[15664] ^ n[15665];
assign t[15666] = t[15665] ^ n[15666];
assign t[15667] = t[15666] ^ n[15667];
assign t[15668] = t[15667] ^ n[15668];
assign t[15669] = t[15668] ^ n[15669];
assign t[15670] = t[15669] ^ n[15670];
assign t[15671] = t[15670] ^ n[15671];
assign t[15672] = t[15671] ^ n[15672];
assign t[15673] = t[15672] ^ n[15673];
assign t[15674] = t[15673] ^ n[15674];
assign t[15675] = t[15674] ^ n[15675];
assign t[15676] = t[15675] ^ n[15676];
assign t[15677] = t[15676] ^ n[15677];
assign t[15678] = t[15677] ^ n[15678];
assign t[15679] = t[15678] ^ n[15679];
assign t[15680] = t[15679] ^ n[15680];
assign t[15681] = t[15680] ^ n[15681];
assign t[15682] = t[15681] ^ n[15682];
assign t[15683] = t[15682] ^ n[15683];
assign t[15684] = t[15683] ^ n[15684];
assign t[15685] = t[15684] ^ n[15685];
assign t[15686] = t[15685] ^ n[15686];
assign t[15687] = t[15686] ^ n[15687];
assign t[15688] = t[15687] ^ n[15688];
assign t[15689] = t[15688] ^ n[15689];
assign t[15690] = t[15689] ^ n[15690];
assign t[15691] = t[15690] ^ n[15691];
assign t[15692] = t[15691] ^ n[15692];
assign t[15693] = t[15692] ^ n[15693];
assign t[15694] = t[15693] ^ n[15694];
assign t[15695] = t[15694] ^ n[15695];
assign t[15696] = t[15695] ^ n[15696];
assign t[15697] = t[15696] ^ n[15697];
assign t[15698] = t[15697] ^ n[15698];
assign t[15699] = t[15698] ^ n[15699];
assign t[15700] = t[15699] ^ n[15700];
assign t[15701] = t[15700] ^ n[15701];
assign t[15702] = t[15701] ^ n[15702];
assign t[15703] = t[15702] ^ n[15703];
assign t[15704] = t[15703] ^ n[15704];
assign t[15705] = t[15704] ^ n[15705];
assign t[15706] = t[15705] ^ n[15706];
assign t[15707] = t[15706] ^ n[15707];
assign t[15708] = t[15707] ^ n[15708];
assign t[15709] = t[15708] ^ n[15709];
assign t[15710] = t[15709] ^ n[15710];
assign t[15711] = t[15710] ^ n[15711];
assign t[15712] = t[15711] ^ n[15712];
assign t[15713] = t[15712] ^ n[15713];
assign t[15714] = t[15713] ^ n[15714];
assign t[15715] = t[15714] ^ n[15715];
assign t[15716] = t[15715] ^ n[15716];
assign t[15717] = t[15716] ^ n[15717];
assign t[15718] = t[15717] ^ n[15718];
assign t[15719] = t[15718] ^ n[15719];
assign t[15720] = t[15719] ^ n[15720];
assign t[15721] = t[15720] ^ n[15721];
assign t[15722] = t[15721] ^ n[15722];
assign t[15723] = t[15722] ^ n[15723];
assign t[15724] = t[15723] ^ n[15724];
assign t[15725] = t[15724] ^ n[15725];
assign t[15726] = t[15725] ^ n[15726];
assign t[15727] = t[15726] ^ n[15727];
assign t[15728] = t[15727] ^ n[15728];
assign t[15729] = t[15728] ^ n[15729];
assign t[15730] = t[15729] ^ n[15730];
assign t[15731] = t[15730] ^ n[15731];
assign t[15732] = t[15731] ^ n[15732];
assign t[15733] = t[15732] ^ n[15733];
assign t[15734] = t[15733] ^ n[15734];
assign t[15735] = t[15734] ^ n[15735];
assign t[15736] = t[15735] ^ n[15736];
assign t[15737] = t[15736] ^ n[15737];
assign t[15738] = t[15737] ^ n[15738];
assign t[15739] = t[15738] ^ n[15739];
assign t[15740] = t[15739] ^ n[15740];
assign t[15741] = t[15740] ^ n[15741];
assign t[15742] = t[15741] ^ n[15742];
assign t[15743] = t[15742] ^ n[15743];
assign t[15744] = t[15743] ^ n[15744];
assign t[15745] = t[15744] ^ n[15745];
assign t[15746] = t[15745] ^ n[15746];
assign t[15747] = t[15746] ^ n[15747];
assign t[15748] = t[15747] ^ n[15748];
assign t[15749] = t[15748] ^ n[15749];
assign t[15750] = t[15749] ^ n[15750];
assign t[15751] = t[15750] ^ n[15751];
assign t[15752] = t[15751] ^ n[15752];
assign t[15753] = t[15752] ^ n[15753];
assign t[15754] = t[15753] ^ n[15754];
assign t[15755] = t[15754] ^ n[15755];
assign t[15756] = t[15755] ^ n[15756];
assign t[15757] = t[15756] ^ n[15757];
assign t[15758] = t[15757] ^ n[15758];
assign t[15759] = t[15758] ^ n[15759];
assign t[15760] = t[15759] ^ n[15760];
assign t[15761] = t[15760] ^ n[15761];
assign t[15762] = t[15761] ^ n[15762];
assign t[15763] = t[15762] ^ n[15763];
assign t[15764] = t[15763] ^ n[15764];
assign t[15765] = t[15764] ^ n[15765];
assign t[15766] = t[15765] ^ n[15766];
assign t[15767] = t[15766] ^ n[15767];
assign t[15768] = t[15767] ^ n[15768];
assign t[15769] = t[15768] ^ n[15769];
assign t[15770] = t[15769] ^ n[15770];
assign t[15771] = t[15770] ^ n[15771];
assign t[15772] = t[15771] ^ n[15772];
assign t[15773] = t[15772] ^ n[15773];
assign t[15774] = t[15773] ^ n[15774];
assign t[15775] = t[15774] ^ n[15775];
assign t[15776] = t[15775] ^ n[15776];
assign t[15777] = t[15776] ^ n[15777];
assign t[15778] = t[15777] ^ n[15778];
assign t[15779] = t[15778] ^ n[15779];
assign t[15780] = t[15779] ^ n[15780];
assign t[15781] = t[15780] ^ n[15781];
assign t[15782] = t[15781] ^ n[15782];
assign t[15783] = t[15782] ^ n[15783];
assign t[15784] = t[15783] ^ n[15784];
assign t[15785] = t[15784] ^ n[15785];
assign t[15786] = t[15785] ^ n[15786];
assign t[15787] = t[15786] ^ n[15787];
assign t[15788] = t[15787] ^ n[15788];
assign t[15789] = t[15788] ^ n[15789];
assign t[15790] = t[15789] ^ n[15790];
assign t[15791] = t[15790] ^ n[15791];
assign t[15792] = t[15791] ^ n[15792];
assign t[15793] = t[15792] ^ n[15793];
assign t[15794] = t[15793] ^ n[15794];
assign t[15795] = t[15794] ^ n[15795];
assign t[15796] = t[15795] ^ n[15796];
assign t[15797] = t[15796] ^ n[15797];
assign t[15798] = t[15797] ^ n[15798];
assign t[15799] = t[15798] ^ n[15799];
assign t[15800] = t[15799] ^ n[15800];
assign t[15801] = t[15800] ^ n[15801];
assign t[15802] = t[15801] ^ n[15802];
assign t[15803] = t[15802] ^ n[15803];
assign t[15804] = t[15803] ^ n[15804];
assign t[15805] = t[15804] ^ n[15805];
assign t[15806] = t[15805] ^ n[15806];
assign t[15807] = t[15806] ^ n[15807];
assign t[15808] = t[15807] ^ n[15808];
assign t[15809] = t[15808] ^ n[15809];
assign t[15810] = t[15809] ^ n[15810];
assign t[15811] = t[15810] ^ n[15811];
assign t[15812] = t[15811] ^ n[15812];
assign t[15813] = t[15812] ^ n[15813];
assign t[15814] = t[15813] ^ n[15814];
assign t[15815] = t[15814] ^ n[15815];
assign t[15816] = t[15815] ^ n[15816];
assign t[15817] = t[15816] ^ n[15817];
assign t[15818] = t[15817] ^ n[15818];
assign t[15819] = t[15818] ^ n[15819];
assign t[15820] = t[15819] ^ n[15820];
assign t[15821] = t[15820] ^ n[15821];
assign t[15822] = t[15821] ^ n[15822];
assign t[15823] = t[15822] ^ n[15823];
assign t[15824] = t[15823] ^ n[15824];
assign t[15825] = t[15824] ^ n[15825];
assign t[15826] = t[15825] ^ n[15826];
assign t[15827] = t[15826] ^ n[15827];
assign t[15828] = t[15827] ^ n[15828];
assign t[15829] = t[15828] ^ n[15829];
assign t[15830] = t[15829] ^ n[15830];
assign t[15831] = t[15830] ^ n[15831];
assign t[15832] = t[15831] ^ n[15832];
assign t[15833] = t[15832] ^ n[15833];
assign t[15834] = t[15833] ^ n[15834];
assign t[15835] = t[15834] ^ n[15835];
assign t[15836] = t[15835] ^ n[15836];
assign t[15837] = t[15836] ^ n[15837];
assign t[15838] = t[15837] ^ n[15838];
assign t[15839] = t[15838] ^ n[15839];
assign t[15840] = t[15839] ^ n[15840];
assign t[15841] = t[15840] ^ n[15841];
assign t[15842] = t[15841] ^ n[15842];
assign t[15843] = t[15842] ^ n[15843];
assign t[15844] = t[15843] ^ n[15844];
assign t[15845] = t[15844] ^ n[15845];
assign t[15846] = t[15845] ^ n[15846];
assign t[15847] = t[15846] ^ n[15847];
assign t[15848] = t[15847] ^ n[15848];
assign t[15849] = t[15848] ^ n[15849];
assign t[15850] = t[15849] ^ n[15850];
assign t[15851] = t[15850] ^ n[15851];
assign t[15852] = t[15851] ^ n[15852];
assign t[15853] = t[15852] ^ n[15853];
assign t[15854] = t[15853] ^ n[15854];
assign t[15855] = t[15854] ^ n[15855];
assign t[15856] = t[15855] ^ n[15856];
assign t[15857] = t[15856] ^ n[15857];
assign t[15858] = t[15857] ^ n[15858];
assign t[15859] = t[15858] ^ n[15859];
assign t[15860] = t[15859] ^ n[15860];
assign t[15861] = t[15860] ^ n[15861];
assign t[15862] = t[15861] ^ n[15862];
assign t[15863] = t[15862] ^ n[15863];
assign t[15864] = t[15863] ^ n[15864];
assign t[15865] = t[15864] ^ n[15865];
assign t[15866] = t[15865] ^ n[15866];
assign t[15867] = t[15866] ^ n[15867];
assign t[15868] = t[15867] ^ n[15868];
assign t[15869] = t[15868] ^ n[15869];
assign t[15870] = t[15869] ^ n[15870];
assign t[15871] = t[15870] ^ n[15871];
assign t[15872] = t[15871] ^ n[15872];
assign t[15873] = t[15872] ^ n[15873];
assign t[15874] = t[15873] ^ n[15874];
assign t[15875] = t[15874] ^ n[15875];
assign t[15876] = t[15875] ^ n[15876];
assign t[15877] = t[15876] ^ n[15877];
assign t[15878] = t[15877] ^ n[15878];
assign t[15879] = t[15878] ^ n[15879];
assign t[15880] = t[15879] ^ n[15880];
assign t[15881] = t[15880] ^ n[15881];
assign t[15882] = t[15881] ^ n[15882];
assign t[15883] = t[15882] ^ n[15883];
assign t[15884] = t[15883] ^ n[15884];
assign t[15885] = t[15884] ^ n[15885];
assign t[15886] = t[15885] ^ n[15886];
assign t[15887] = t[15886] ^ n[15887];
assign t[15888] = t[15887] ^ n[15888];
assign t[15889] = t[15888] ^ n[15889];
assign t[15890] = t[15889] ^ n[15890];
assign t[15891] = t[15890] ^ n[15891];
assign t[15892] = t[15891] ^ n[15892];
assign t[15893] = t[15892] ^ n[15893];
assign t[15894] = t[15893] ^ n[15894];
assign t[15895] = t[15894] ^ n[15895];
assign t[15896] = t[15895] ^ n[15896];
assign t[15897] = t[15896] ^ n[15897];
assign t[15898] = t[15897] ^ n[15898];
assign t[15899] = t[15898] ^ n[15899];
assign t[15900] = t[15899] ^ n[15900];
assign t[15901] = t[15900] ^ n[15901];
assign t[15902] = t[15901] ^ n[15902];
assign t[15903] = t[15902] ^ n[15903];
assign t[15904] = t[15903] ^ n[15904];
assign t[15905] = t[15904] ^ n[15905];
assign t[15906] = t[15905] ^ n[15906];
assign t[15907] = t[15906] ^ n[15907];
assign t[15908] = t[15907] ^ n[15908];
assign t[15909] = t[15908] ^ n[15909];
assign t[15910] = t[15909] ^ n[15910];
assign t[15911] = t[15910] ^ n[15911];
assign t[15912] = t[15911] ^ n[15912];
assign t[15913] = t[15912] ^ n[15913];
assign t[15914] = t[15913] ^ n[15914];
assign t[15915] = t[15914] ^ n[15915];
assign t[15916] = t[15915] ^ n[15916];
assign t[15917] = t[15916] ^ n[15917];
assign t[15918] = t[15917] ^ n[15918];
assign t[15919] = t[15918] ^ n[15919];
assign t[15920] = t[15919] ^ n[15920];
assign t[15921] = t[15920] ^ n[15921];
assign t[15922] = t[15921] ^ n[15922];
assign t[15923] = t[15922] ^ n[15923];
assign t[15924] = t[15923] ^ n[15924];
assign t[15925] = t[15924] ^ n[15925];
assign t[15926] = t[15925] ^ n[15926];
assign t[15927] = t[15926] ^ n[15927];
assign t[15928] = t[15927] ^ n[15928];
assign t[15929] = t[15928] ^ n[15929];
assign t[15930] = t[15929] ^ n[15930];
assign t[15931] = t[15930] ^ n[15931];
assign t[15932] = t[15931] ^ n[15932];
assign t[15933] = t[15932] ^ n[15933];
assign t[15934] = t[15933] ^ n[15934];
assign t[15935] = t[15934] ^ n[15935];
assign t[15936] = t[15935] ^ n[15936];
assign t[15937] = t[15936] ^ n[15937];
assign t[15938] = t[15937] ^ n[15938];
assign t[15939] = t[15938] ^ n[15939];
assign t[15940] = t[15939] ^ n[15940];
assign t[15941] = t[15940] ^ n[15941];
assign t[15942] = t[15941] ^ n[15942];
assign t[15943] = t[15942] ^ n[15943];
assign t[15944] = t[15943] ^ n[15944];
assign t[15945] = t[15944] ^ n[15945];
assign t[15946] = t[15945] ^ n[15946];
assign t[15947] = t[15946] ^ n[15947];
assign t[15948] = t[15947] ^ n[15948];
assign t[15949] = t[15948] ^ n[15949];
assign t[15950] = t[15949] ^ n[15950];
assign t[15951] = t[15950] ^ n[15951];
assign t[15952] = t[15951] ^ n[15952];
assign t[15953] = t[15952] ^ n[15953];
assign t[15954] = t[15953] ^ n[15954];
assign t[15955] = t[15954] ^ n[15955];
assign t[15956] = t[15955] ^ n[15956];
assign t[15957] = t[15956] ^ n[15957];
assign t[15958] = t[15957] ^ n[15958];
assign t[15959] = t[15958] ^ n[15959];
assign t[15960] = t[15959] ^ n[15960];
assign t[15961] = t[15960] ^ n[15961];
assign t[15962] = t[15961] ^ n[15962];
assign t[15963] = t[15962] ^ n[15963];
assign t[15964] = t[15963] ^ n[15964];
assign t[15965] = t[15964] ^ n[15965];
assign t[15966] = t[15965] ^ n[15966];
assign t[15967] = t[15966] ^ n[15967];
assign t[15968] = t[15967] ^ n[15968];
assign t[15969] = t[15968] ^ n[15969];
assign t[15970] = t[15969] ^ n[15970];
assign t[15971] = t[15970] ^ n[15971];
assign t[15972] = t[15971] ^ n[15972];
assign t[15973] = t[15972] ^ n[15973];
assign t[15974] = t[15973] ^ n[15974];
assign t[15975] = t[15974] ^ n[15975];
assign t[15976] = t[15975] ^ n[15976];
assign t[15977] = t[15976] ^ n[15977];
assign t[15978] = t[15977] ^ n[15978];
assign t[15979] = t[15978] ^ n[15979];
assign t[15980] = t[15979] ^ n[15980];
assign t[15981] = t[15980] ^ n[15981];
assign t[15982] = t[15981] ^ n[15982];
assign t[15983] = t[15982] ^ n[15983];
assign t[15984] = t[15983] ^ n[15984];
assign t[15985] = t[15984] ^ n[15985];
assign t[15986] = t[15985] ^ n[15986];
assign t[15987] = t[15986] ^ n[15987];
assign t[15988] = t[15987] ^ n[15988];
assign t[15989] = t[15988] ^ n[15989];
assign t[15990] = t[15989] ^ n[15990];
assign t[15991] = t[15990] ^ n[15991];
assign t[15992] = t[15991] ^ n[15992];
assign t[15993] = t[15992] ^ n[15993];
assign t[15994] = t[15993] ^ n[15994];
assign t[15995] = t[15994] ^ n[15995];
assign t[15996] = t[15995] ^ n[15996];
assign t[15997] = t[15996] ^ n[15997];
assign t[15998] = t[15997] ^ n[15998];
assign t[15999] = t[15998] ^ n[15999];
assign t[16000] = t[15999] ^ n[16000];
assign t[16001] = t[16000] ^ n[16001];
assign t[16002] = t[16001] ^ n[16002];
assign t[16003] = t[16002] ^ n[16003];
assign t[16004] = t[16003] ^ n[16004];
assign t[16005] = t[16004] ^ n[16005];
assign t[16006] = t[16005] ^ n[16006];
assign t[16007] = t[16006] ^ n[16007];
assign t[16008] = t[16007] ^ n[16008];
assign t[16009] = t[16008] ^ n[16009];
assign t[16010] = t[16009] ^ n[16010];
assign t[16011] = t[16010] ^ n[16011];
assign t[16012] = t[16011] ^ n[16012];
assign t[16013] = t[16012] ^ n[16013];
assign t[16014] = t[16013] ^ n[16014];
assign t[16015] = t[16014] ^ n[16015];
assign t[16016] = t[16015] ^ n[16016];
assign t[16017] = t[16016] ^ n[16017];
assign t[16018] = t[16017] ^ n[16018];
assign t[16019] = t[16018] ^ n[16019];
assign t[16020] = t[16019] ^ n[16020];
assign t[16021] = t[16020] ^ n[16021];
assign t[16022] = t[16021] ^ n[16022];
assign t[16023] = t[16022] ^ n[16023];
assign t[16024] = t[16023] ^ n[16024];
assign t[16025] = t[16024] ^ n[16025];
assign t[16026] = t[16025] ^ n[16026];
assign t[16027] = t[16026] ^ n[16027];
assign t[16028] = t[16027] ^ n[16028];
assign t[16029] = t[16028] ^ n[16029];
assign t[16030] = t[16029] ^ n[16030];
assign t[16031] = t[16030] ^ n[16031];
assign t[16032] = t[16031] ^ n[16032];
assign t[16033] = t[16032] ^ n[16033];
assign t[16034] = t[16033] ^ n[16034];
assign t[16035] = t[16034] ^ n[16035];
assign t[16036] = t[16035] ^ n[16036];
assign t[16037] = t[16036] ^ n[16037];
assign t[16038] = t[16037] ^ n[16038];
assign t[16039] = t[16038] ^ n[16039];
assign t[16040] = t[16039] ^ n[16040];
assign t[16041] = t[16040] ^ n[16041];
assign t[16042] = t[16041] ^ n[16042];
assign t[16043] = t[16042] ^ n[16043];
assign t[16044] = t[16043] ^ n[16044];
assign t[16045] = t[16044] ^ n[16045];
assign t[16046] = t[16045] ^ n[16046];
assign t[16047] = t[16046] ^ n[16047];
assign t[16048] = t[16047] ^ n[16048];
assign t[16049] = t[16048] ^ n[16049];
assign t[16050] = t[16049] ^ n[16050];
assign t[16051] = t[16050] ^ n[16051];
assign t[16052] = t[16051] ^ n[16052];
assign t[16053] = t[16052] ^ n[16053];
assign t[16054] = t[16053] ^ n[16054];
assign t[16055] = t[16054] ^ n[16055];
assign t[16056] = t[16055] ^ n[16056];
assign t[16057] = t[16056] ^ n[16057];
assign t[16058] = t[16057] ^ n[16058];
assign t[16059] = t[16058] ^ n[16059];
assign t[16060] = t[16059] ^ n[16060];
assign t[16061] = t[16060] ^ n[16061];
assign t[16062] = t[16061] ^ n[16062];
assign t[16063] = t[16062] ^ n[16063];
assign t[16064] = t[16063] ^ n[16064];
assign t[16065] = t[16064] ^ n[16065];
assign t[16066] = t[16065] ^ n[16066];
assign t[16067] = t[16066] ^ n[16067];
assign t[16068] = t[16067] ^ n[16068];
assign t[16069] = t[16068] ^ n[16069];
assign t[16070] = t[16069] ^ n[16070];
assign t[16071] = t[16070] ^ n[16071];
assign t[16072] = t[16071] ^ n[16072];
assign t[16073] = t[16072] ^ n[16073];
assign t[16074] = t[16073] ^ n[16074];
assign t[16075] = t[16074] ^ n[16075];
assign t[16076] = t[16075] ^ n[16076];
assign t[16077] = t[16076] ^ n[16077];
assign t[16078] = t[16077] ^ n[16078];
assign t[16079] = t[16078] ^ n[16079];
assign t[16080] = t[16079] ^ n[16080];
assign t[16081] = t[16080] ^ n[16081];
assign t[16082] = t[16081] ^ n[16082];
assign t[16083] = t[16082] ^ n[16083];
assign t[16084] = t[16083] ^ n[16084];
assign t[16085] = t[16084] ^ n[16085];
assign t[16086] = t[16085] ^ n[16086];
assign t[16087] = t[16086] ^ n[16087];
assign t[16088] = t[16087] ^ n[16088];
assign t[16089] = t[16088] ^ n[16089];
assign t[16090] = t[16089] ^ n[16090];
assign t[16091] = t[16090] ^ n[16091];
assign t[16092] = t[16091] ^ n[16092];
assign t[16093] = t[16092] ^ n[16093];
assign t[16094] = t[16093] ^ n[16094];
assign t[16095] = t[16094] ^ n[16095];
assign t[16096] = t[16095] ^ n[16096];
assign t[16097] = t[16096] ^ n[16097];
assign t[16098] = t[16097] ^ n[16098];
assign t[16099] = t[16098] ^ n[16099];
assign t[16100] = t[16099] ^ n[16100];
assign t[16101] = t[16100] ^ n[16101];
assign t[16102] = t[16101] ^ n[16102];
assign t[16103] = t[16102] ^ n[16103];
assign t[16104] = t[16103] ^ n[16104];
assign t[16105] = t[16104] ^ n[16105];
assign t[16106] = t[16105] ^ n[16106];
assign t[16107] = t[16106] ^ n[16107];
assign t[16108] = t[16107] ^ n[16108];
assign t[16109] = t[16108] ^ n[16109];
assign t[16110] = t[16109] ^ n[16110];
assign t[16111] = t[16110] ^ n[16111];
assign t[16112] = t[16111] ^ n[16112];
assign t[16113] = t[16112] ^ n[16113];
assign t[16114] = t[16113] ^ n[16114];
assign t[16115] = t[16114] ^ n[16115];
assign t[16116] = t[16115] ^ n[16116];
assign t[16117] = t[16116] ^ n[16117];
assign t[16118] = t[16117] ^ n[16118];
assign t[16119] = t[16118] ^ n[16119];
assign t[16120] = t[16119] ^ n[16120];
assign t[16121] = t[16120] ^ n[16121];
assign t[16122] = t[16121] ^ n[16122];
assign t[16123] = t[16122] ^ n[16123];
assign t[16124] = t[16123] ^ n[16124];
assign t[16125] = t[16124] ^ n[16125];
assign t[16126] = t[16125] ^ n[16126];
assign t[16127] = t[16126] ^ n[16127];
assign t[16128] = t[16127] ^ n[16128];
assign t[16129] = t[16128] ^ n[16129];
assign t[16130] = t[16129] ^ n[16130];
assign t[16131] = t[16130] ^ n[16131];
assign t[16132] = t[16131] ^ n[16132];
assign t[16133] = t[16132] ^ n[16133];
assign t[16134] = t[16133] ^ n[16134];
assign t[16135] = t[16134] ^ n[16135];
assign t[16136] = t[16135] ^ n[16136];
assign t[16137] = t[16136] ^ n[16137];
assign t[16138] = t[16137] ^ n[16138];
assign t[16139] = t[16138] ^ n[16139];
assign t[16140] = t[16139] ^ n[16140];
assign t[16141] = t[16140] ^ n[16141];
assign t[16142] = t[16141] ^ n[16142];
assign t[16143] = t[16142] ^ n[16143];
assign t[16144] = t[16143] ^ n[16144];
assign t[16145] = t[16144] ^ n[16145];
assign t[16146] = t[16145] ^ n[16146];
assign t[16147] = t[16146] ^ n[16147];
assign t[16148] = t[16147] ^ n[16148];
assign t[16149] = t[16148] ^ n[16149];
assign t[16150] = t[16149] ^ n[16150];
assign t[16151] = t[16150] ^ n[16151];
assign t[16152] = t[16151] ^ n[16152];
assign t[16153] = t[16152] ^ n[16153];
assign t[16154] = t[16153] ^ n[16154];
assign t[16155] = t[16154] ^ n[16155];
assign t[16156] = t[16155] ^ n[16156];
assign t[16157] = t[16156] ^ n[16157];
assign t[16158] = t[16157] ^ n[16158];
assign t[16159] = t[16158] ^ n[16159];
assign t[16160] = t[16159] ^ n[16160];
assign t[16161] = t[16160] ^ n[16161];
assign t[16162] = t[16161] ^ n[16162];
assign t[16163] = t[16162] ^ n[16163];
assign t[16164] = t[16163] ^ n[16164];
assign t[16165] = t[16164] ^ n[16165];
assign t[16166] = t[16165] ^ n[16166];
assign t[16167] = t[16166] ^ n[16167];
assign t[16168] = t[16167] ^ n[16168];
assign t[16169] = t[16168] ^ n[16169];
assign t[16170] = t[16169] ^ n[16170];
assign t[16171] = t[16170] ^ n[16171];
assign t[16172] = t[16171] ^ n[16172];
assign t[16173] = t[16172] ^ n[16173];
assign t[16174] = t[16173] ^ n[16174];
assign t[16175] = t[16174] ^ n[16175];
assign t[16176] = t[16175] ^ n[16176];
assign t[16177] = t[16176] ^ n[16177];
assign t[16178] = t[16177] ^ n[16178];
assign t[16179] = t[16178] ^ n[16179];
assign t[16180] = t[16179] ^ n[16180];
assign t[16181] = t[16180] ^ n[16181];
assign t[16182] = t[16181] ^ n[16182];
assign t[16183] = t[16182] ^ n[16183];
assign t[16184] = t[16183] ^ n[16184];
assign t[16185] = t[16184] ^ n[16185];
assign t[16186] = t[16185] ^ n[16186];
assign t[16187] = t[16186] ^ n[16187];
assign t[16188] = t[16187] ^ n[16188];
assign t[16189] = t[16188] ^ n[16189];
assign t[16190] = t[16189] ^ n[16190];
assign t[16191] = t[16190] ^ n[16191];
assign t[16192] = t[16191] ^ n[16192];
assign t[16193] = t[16192] ^ n[16193];
assign t[16194] = t[16193] ^ n[16194];
assign t[16195] = t[16194] ^ n[16195];
assign t[16196] = t[16195] ^ n[16196];
assign t[16197] = t[16196] ^ n[16197];
assign t[16198] = t[16197] ^ n[16198];
assign t[16199] = t[16198] ^ n[16199];
assign t[16200] = t[16199] ^ n[16200];
assign t[16201] = t[16200] ^ n[16201];
assign t[16202] = t[16201] ^ n[16202];
assign t[16203] = t[16202] ^ n[16203];
assign t[16204] = t[16203] ^ n[16204];
assign t[16205] = t[16204] ^ n[16205];
assign t[16206] = t[16205] ^ n[16206];
assign t[16207] = t[16206] ^ n[16207];
assign t[16208] = t[16207] ^ n[16208];
assign t[16209] = t[16208] ^ n[16209];
assign t[16210] = t[16209] ^ n[16210];
assign t[16211] = t[16210] ^ n[16211];
assign t[16212] = t[16211] ^ n[16212];
assign t[16213] = t[16212] ^ n[16213];
assign t[16214] = t[16213] ^ n[16214];
assign t[16215] = t[16214] ^ n[16215];
assign t[16216] = t[16215] ^ n[16216];
assign t[16217] = t[16216] ^ n[16217];
assign t[16218] = t[16217] ^ n[16218];
assign t[16219] = t[16218] ^ n[16219];
assign t[16220] = t[16219] ^ n[16220];
assign t[16221] = t[16220] ^ n[16221];
assign t[16222] = t[16221] ^ n[16222];
assign t[16223] = t[16222] ^ n[16223];
assign t[16224] = t[16223] ^ n[16224];
assign t[16225] = t[16224] ^ n[16225];
assign t[16226] = t[16225] ^ n[16226];
assign t[16227] = t[16226] ^ n[16227];
assign t[16228] = t[16227] ^ n[16228];
assign t[16229] = t[16228] ^ n[16229];
assign t[16230] = t[16229] ^ n[16230];
assign t[16231] = t[16230] ^ n[16231];
assign t[16232] = t[16231] ^ n[16232];
assign t[16233] = t[16232] ^ n[16233];
assign t[16234] = t[16233] ^ n[16234];
assign t[16235] = t[16234] ^ n[16235];
assign t[16236] = t[16235] ^ n[16236];
assign t[16237] = t[16236] ^ n[16237];
assign t[16238] = t[16237] ^ n[16238];
assign t[16239] = t[16238] ^ n[16239];
assign t[16240] = t[16239] ^ n[16240];
assign t[16241] = t[16240] ^ n[16241];
assign t[16242] = t[16241] ^ n[16242];
assign t[16243] = t[16242] ^ n[16243];
assign t[16244] = t[16243] ^ n[16244];
assign t[16245] = t[16244] ^ n[16245];
assign t[16246] = t[16245] ^ n[16246];
assign t[16247] = t[16246] ^ n[16247];
assign t[16248] = t[16247] ^ n[16248];
assign t[16249] = t[16248] ^ n[16249];
assign t[16250] = t[16249] ^ n[16250];
assign t[16251] = t[16250] ^ n[16251];
assign t[16252] = t[16251] ^ n[16252];
assign t[16253] = t[16252] ^ n[16253];
assign t[16254] = t[16253] ^ n[16254];
assign t[16255] = t[16254] ^ n[16255];
assign t[16256] = t[16255] ^ n[16256];
assign t[16257] = t[16256] ^ n[16257];
assign t[16258] = t[16257] ^ n[16258];
assign t[16259] = t[16258] ^ n[16259];
assign t[16260] = t[16259] ^ n[16260];
assign t[16261] = t[16260] ^ n[16261];
assign t[16262] = t[16261] ^ n[16262];
assign t[16263] = t[16262] ^ n[16263];
assign t[16264] = t[16263] ^ n[16264];
assign t[16265] = t[16264] ^ n[16265];
assign t[16266] = t[16265] ^ n[16266];
assign t[16267] = t[16266] ^ n[16267];
assign t[16268] = t[16267] ^ n[16268];
assign t[16269] = t[16268] ^ n[16269];
assign t[16270] = t[16269] ^ n[16270];
assign t[16271] = t[16270] ^ n[16271];
assign t[16272] = t[16271] ^ n[16272];
assign t[16273] = t[16272] ^ n[16273];
assign t[16274] = t[16273] ^ n[16274];
assign t[16275] = t[16274] ^ n[16275];
assign t[16276] = t[16275] ^ n[16276];
assign t[16277] = t[16276] ^ n[16277];
assign t[16278] = t[16277] ^ n[16278];
assign t[16279] = t[16278] ^ n[16279];
assign t[16280] = t[16279] ^ n[16280];
assign t[16281] = t[16280] ^ n[16281];
assign t[16282] = t[16281] ^ n[16282];
assign t[16283] = t[16282] ^ n[16283];
assign t[16284] = t[16283] ^ n[16284];
assign t[16285] = t[16284] ^ n[16285];
assign t[16286] = t[16285] ^ n[16286];
assign t[16287] = t[16286] ^ n[16287];
assign t[16288] = t[16287] ^ n[16288];
assign t[16289] = t[16288] ^ n[16289];
assign t[16290] = t[16289] ^ n[16290];
assign t[16291] = t[16290] ^ n[16291];
assign t[16292] = t[16291] ^ n[16292];
assign t[16293] = t[16292] ^ n[16293];
assign t[16294] = t[16293] ^ n[16294];
assign t[16295] = t[16294] ^ n[16295];
assign t[16296] = t[16295] ^ n[16296];
assign t[16297] = t[16296] ^ n[16297];
assign t[16298] = t[16297] ^ n[16298];
assign t[16299] = t[16298] ^ n[16299];
assign t[16300] = t[16299] ^ n[16300];
assign t[16301] = t[16300] ^ n[16301];
assign t[16302] = t[16301] ^ n[16302];
assign t[16303] = t[16302] ^ n[16303];
assign t[16304] = t[16303] ^ n[16304];
assign t[16305] = t[16304] ^ n[16305];
assign t[16306] = t[16305] ^ n[16306];
assign t[16307] = t[16306] ^ n[16307];
assign t[16308] = t[16307] ^ n[16308];
assign t[16309] = t[16308] ^ n[16309];
assign t[16310] = t[16309] ^ n[16310];
assign t[16311] = t[16310] ^ n[16311];
assign t[16312] = t[16311] ^ n[16312];
assign t[16313] = t[16312] ^ n[16313];
assign t[16314] = t[16313] ^ n[16314];
assign t[16315] = t[16314] ^ n[16315];
assign t[16316] = t[16315] ^ n[16316];
assign t[16317] = t[16316] ^ n[16317];
assign t[16318] = t[16317] ^ n[16318];
assign t[16319] = t[16318] ^ n[16319];
assign t[16320] = t[16319] ^ n[16320];
assign t[16321] = t[16320] ^ n[16321];
assign t[16322] = t[16321] ^ n[16322];
assign t[16323] = t[16322] ^ n[16323];
assign t[16324] = t[16323] ^ n[16324];
assign t[16325] = t[16324] ^ n[16325];
assign t[16326] = t[16325] ^ n[16326];
assign t[16327] = t[16326] ^ n[16327];
assign t[16328] = t[16327] ^ n[16328];
assign t[16329] = t[16328] ^ n[16329];
assign t[16330] = t[16329] ^ n[16330];
assign t[16331] = t[16330] ^ n[16331];
assign t[16332] = t[16331] ^ n[16332];
assign t[16333] = t[16332] ^ n[16333];
assign t[16334] = t[16333] ^ n[16334];
assign t[16335] = t[16334] ^ n[16335];
assign t[16336] = t[16335] ^ n[16336];
assign t[16337] = t[16336] ^ n[16337];
assign t[16338] = t[16337] ^ n[16338];
assign t[16339] = t[16338] ^ n[16339];
assign t[16340] = t[16339] ^ n[16340];
assign t[16341] = t[16340] ^ n[16341];
assign t[16342] = t[16341] ^ n[16342];
assign t[16343] = t[16342] ^ n[16343];
assign t[16344] = t[16343] ^ n[16344];
assign t[16345] = t[16344] ^ n[16345];
assign t[16346] = t[16345] ^ n[16346];
assign t[16347] = t[16346] ^ n[16347];
assign t[16348] = t[16347] ^ n[16348];
assign t[16349] = t[16348] ^ n[16349];
assign t[16350] = t[16349] ^ n[16350];
assign t[16351] = t[16350] ^ n[16351];
assign t[16352] = t[16351] ^ n[16352];
assign t[16353] = t[16352] ^ n[16353];
assign t[16354] = t[16353] ^ n[16354];
assign t[16355] = t[16354] ^ n[16355];
assign t[16356] = t[16355] ^ n[16356];
assign t[16357] = t[16356] ^ n[16357];
assign t[16358] = t[16357] ^ n[16358];
assign t[16359] = t[16358] ^ n[16359];
assign t[16360] = t[16359] ^ n[16360];
assign t[16361] = t[16360] ^ n[16361];
assign t[16362] = t[16361] ^ n[16362];
assign t[16363] = t[16362] ^ n[16363];
assign t[16364] = t[16363] ^ n[16364];
assign t[16365] = t[16364] ^ n[16365];
assign t[16366] = t[16365] ^ n[16366];
assign t[16367] = t[16366] ^ n[16367];
assign t[16368] = t[16367] ^ n[16368];

//asigning bit 13
assign s[13] = ( a[13] ^ b [13] ) ^ t[16368];

assign t[16369] = n[16369];
assign t[16370] = t[16369] ^ n[16370];
assign t[16371] = t[16370] ^ n[16371];
assign t[16372] = t[16371] ^ n[16372];
assign t[16373] = t[16372] ^ n[16373];
assign t[16374] = t[16373] ^ n[16374];
assign t[16375] = t[16374] ^ n[16375];
assign t[16376] = t[16375] ^ n[16376];
assign t[16377] = t[16376] ^ n[16377];
assign t[16378] = t[16377] ^ n[16378];
assign t[16379] = t[16378] ^ n[16379];
assign t[16380] = t[16379] ^ n[16380];
assign t[16381] = t[16380] ^ n[16381];
assign t[16382] = t[16381] ^ n[16382];
assign t[16383] = t[16382] ^ n[16383];
assign t[16384] = t[16383] ^ n[16384];
assign t[16385] = t[16384] ^ n[16385];
assign t[16386] = t[16385] ^ n[16386];
assign t[16387] = t[16386] ^ n[16387];
assign t[16388] = t[16387] ^ n[16388];
assign t[16389] = t[16388] ^ n[16389];
assign t[16390] = t[16389] ^ n[16390];
assign t[16391] = t[16390] ^ n[16391];
assign t[16392] = t[16391] ^ n[16392];
assign t[16393] = t[16392] ^ n[16393];
assign t[16394] = t[16393] ^ n[16394];
assign t[16395] = t[16394] ^ n[16395];
assign t[16396] = t[16395] ^ n[16396];
assign t[16397] = t[16396] ^ n[16397];
assign t[16398] = t[16397] ^ n[16398];
assign t[16399] = t[16398] ^ n[16399];
assign t[16400] = t[16399] ^ n[16400];
assign t[16401] = t[16400] ^ n[16401];
assign t[16402] = t[16401] ^ n[16402];
assign t[16403] = t[16402] ^ n[16403];
assign t[16404] = t[16403] ^ n[16404];
assign t[16405] = t[16404] ^ n[16405];
assign t[16406] = t[16405] ^ n[16406];
assign t[16407] = t[16406] ^ n[16407];
assign t[16408] = t[16407] ^ n[16408];
assign t[16409] = t[16408] ^ n[16409];
assign t[16410] = t[16409] ^ n[16410];
assign t[16411] = t[16410] ^ n[16411];
assign t[16412] = t[16411] ^ n[16412];
assign t[16413] = t[16412] ^ n[16413];
assign t[16414] = t[16413] ^ n[16414];
assign t[16415] = t[16414] ^ n[16415];
assign t[16416] = t[16415] ^ n[16416];
assign t[16417] = t[16416] ^ n[16417];
assign t[16418] = t[16417] ^ n[16418];
assign t[16419] = t[16418] ^ n[16419];
assign t[16420] = t[16419] ^ n[16420];
assign t[16421] = t[16420] ^ n[16421];
assign t[16422] = t[16421] ^ n[16422];
assign t[16423] = t[16422] ^ n[16423];
assign t[16424] = t[16423] ^ n[16424];
assign t[16425] = t[16424] ^ n[16425];
assign t[16426] = t[16425] ^ n[16426];
assign t[16427] = t[16426] ^ n[16427];
assign t[16428] = t[16427] ^ n[16428];
assign t[16429] = t[16428] ^ n[16429];
assign t[16430] = t[16429] ^ n[16430];
assign t[16431] = t[16430] ^ n[16431];
assign t[16432] = t[16431] ^ n[16432];
assign t[16433] = t[16432] ^ n[16433];
assign t[16434] = t[16433] ^ n[16434];
assign t[16435] = t[16434] ^ n[16435];
assign t[16436] = t[16435] ^ n[16436];
assign t[16437] = t[16436] ^ n[16437];
assign t[16438] = t[16437] ^ n[16438];
assign t[16439] = t[16438] ^ n[16439];
assign t[16440] = t[16439] ^ n[16440];
assign t[16441] = t[16440] ^ n[16441];
assign t[16442] = t[16441] ^ n[16442];
assign t[16443] = t[16442] ^ n[16443];
assign t[16444] = t[16443] ^ n[16444];
assign t[16445] = t[16444] ^ n[16445];
assign t[16446] = t[16445] ^ n[16446];
assign t[16447] = t[16446] ^ n[16447];
assign t[16448] = t[16447] ^ n[16448];
assign t[16449] = t[16448] ^ n[16449];
assign t[16450] = t[16449] ^ n[16450];
assign t[16451] = t[16450] ^ n[16451];
assign t[16452] = t[16451] ^ n[16452];
assign t[16453] = t[16452] ^ n[16453];
assign t[16454] = t[16453] ^ n[16454];
assign t[16455] = t[16454] ^ n[16455];
assign t[16456] = t[16455] ^ n[16456];
assign t[16457] = t[16456] ^ n[16457];
assign t[16458] = t[16457] ^ n[16458];
assign t[16459] = t[16458] ^ n[16459];
assign t[16460] = t[16459] ^ n[16460];
assign t[16461] = t[16460] ^ n[16461];
assign t[16462] = t[16461] ^ n[16462];
assign t[16463] = t[16462] ^ n[16463];
assign t[16464] = t[16463] ^ n[16464];
assign t[16465] = t[16464] ^ n[16465];
assign t[16466] = t[16465] ^ n[16466];
assign t[16467] = t[16466] ^ n[16467];
assign t[16468] = t[16467] ^ n[16468];
assign t[16469] = t[16468] ^ n[16469];
assign t[16470] = t[16469] ^ n[16470];
assign t[16471] = t[16470] ^ n[16471];
assign t[16472] = t[16471] ^ n[16472];
assign t[16473] = t[16472] ^ n[16473];
assign t[16474] = t[16473] ^ n[16474];
assign t[16475] = t[16474] ^ n[16475];
assign t[16476] = t[16475] ^ n[16476];
assign t[16477] = t[16476] ^ n[16477];
assign t[16478] = t[16477] ^ n[16478];
assign t[16479] = t[16478] ^ n[16479];
assign t[16480] = t[16479] ^ n[16480];
assign t[16481] = t[16480] ^ n[16481];
assign t[16482] = t[16481] ^ n[16482];
assign t[16483] = t[16482] ^ n[16483];
assign t[16484] = t[16483] ^ n[16484];
assign t[16485] = t[16484] ^ n[16485];
assign t[16486] = t[16485] ^ n[16486];
assign t[16487] = t[16486] ^ n[16487];
assign t[16488] = t[16487] ^ n[16488];
assign t[16489] = t[16488] ^ n[16489];
assign t[16490] = t[16489] ^ n[16490];
assign t[16491] = t[16490] ^ n[16491];
assign t[16492] = t[16491] ^ n[16492];
assign t[16493] = t[16492] ^ n[16493];
assign t[16494] = t[16493] ^ n[16494];
assign t[16495] = t[16494] ^ n[16495];
assign t[16496] = t[16495] ^ n[16496];
assign t[16497] = t[16496] ^ n[16497];
assign t[16498] = t[16497] ^ n[16498];
assign t[16499] = t[16498] ^ n[16499];
assign t[16500] = t[16499] ^ n[16500];
assign t[16501] = t[16500] ^ n[16501];
assign t[16502] = t[16501] ^ n[16502];
assign t[16503] = t[16502] ^ n[16503];
assign t[16504] = t[16503] ^ n[16504];
assign t[16505] = t[16504] ^ n[16505];
assign t[16506] = t[16505] ^ n[16506];
assign t[16507] = t[16506] ^ n[16507];
assign t[16508] = t[16507] ^ n[16508];
assign t[16509] = t[16508] ^ n[16509];
assign t[16510] = t[16509] ^ n[16510];
assign t[16511] = t[16510] ^ n[16511];
assign t[16512] = t[16511] ^ n[16512];
assign t[16513] = t[16512] ^ n[16513];
assign t[16514] = t[16513] ^ n[16514];
assign t[16515] = t[16514] ^ n[16515];
assign t[16516] = t[16515] ^ n[16516];
assign t[16517] = t[16516] ^ n[16517];
assign t[16518] = t[16517] ^ n[16518];
assign t[16519] = t[16518] ^ n[16519];
assign t[16520] = t[16519] ^ n[16520];
assign t[16521] = t[16520] ^ n[16521];
assign t[16522] = t[16521] ^ n[16522];
assign t[16523] = t[16522] ^ n[16523];
assign t[16524] = t[16523] ^ n[16524];
assign t[16525] = t[16524] ^ n[16525];
assign t[16526] = t[16525] ^ n[16526];
assign t[16527] = t[16526] ^ n[16527];
assign t[16528] = t[16527] ^ n[16528];
assign t[16529] = t[16528] ^ n[16529];
assign t[16530] = t[16529] ^ n[16530];
assign t[16531] = t[16530] ^ n[16531];
assign t[16532] = t[16531] ^ n[16532];
assign t[16533] = t[16532] ^ n[16533];
assign t[16534] = t[16533] ^ n[16534];
assign t[16535] = t[16534] ^ n[16535];
assign t[16536] = t[16535] ^ n[16536];
assign t[16537] = t[16536] ^ n[16537];
assign t[16538] = t[16537] ^ n[16538];
assign t[16539] = t[16538] ^ n[16539];
assign t[16540] = t[16539] ^ n[16540];
assign t[16541] = t[16540] ^ n[16541];
assign t[16542] = t[16541] ^ n[16542];
assign t[16543] = t[16542] ^ n[16543];
assign t[16544] = t[16543] ^ n[16544];
assign t[16545] = t[16544] ^ n[16545];
assign t[16546] = t[16545] ^ n[16546];
assign t[16547] = t[16546] ^ n[16547];
assign t[16548] = t[16547] ^ n[16548];
assign t[16549] = t[16548] ^ n[16549];
assign t[16550] = t[16549] ^ n[16550];
assign t[16551] = t[16550] ^ n[16551];
assign t[16552] = t[16551] ^ n[16552];
assign t[16553] = t[16552] ^ n[16553];
assign t[16554] = t[16553] ^ n[16554];
assign t[16555] = t[16554] ^ n[16555];
assign t[16556] = t[16555] ^ n[16556];
assign t[16557] = t[16556] ^ n[16557];
assign t[16558] = t[16557] ^ n[16558];
assign t[16559] = t[16558] ^ n[16559];
assign t[16560] = t[16559] ^ n[16560];
assign t[16561] = t[16560] ^ n[16561];
assign t[16562] = t[16561] ^ n[16562];
assign t[16563] = t[16562] ^ n[16563];
assign t[16564] = t[16563] ^ n[16564];
assign t[16565] = t[16564] ^ n[16565];
assign t[16566] = t[16565] ^ n[16566];
assign t[16567] = t[16566] ^ n[16567];
assign t[16568] = t[16567] ^ n[16568];
assign t[16569] = t[16568] ^ n[16569];
assign t[16570] = t[16569] ^ n[16570];
assign t[16571] = t[16570] ^ n[16571];
assign t[16572] = t[16571] ^ n[16572];
assign t[16573] = t[16572] ^ n[16573];
assign t[16574] = t[16573] ^ n[16574];
assign t[16575] = t[16574] ^ n[16575];
assign t[16576] = t[16575] ^ n[16576];
assign t[16577] = t[16576] ^ n[16577];
assign t[16578] = t[16577] ^ n[16578];
assign t[16579] = t[16578] ^ n[16579];
assign t[16580] = t[16579] ^ n[16580];
assign t[16581] = t[16580] ^ n[16581];
assign t[16582] = t[16581] ^ n[16582];
assign t[16583] = t[16582] ^ n[16583];
assign t[16584] = t[16583] ^ n[16584];
assign t[16585] = t[16584] ^ n[16585];
assign t[16586] = t[16585] ^ n[16586];
assign t[16587] = t[16586] ^ n[16587];
assign t[16588] = t[16587] ^ n[16588];
assign t[16589] = t[16588] ^ n[16589];
assign t[16590] = t[16589] ^ n[16590];
assign t[16591] = t[16590] ^ n[16591];
assign t[16592] = t[16591] ^ n[16592];
assign t[16593] = t[16592] ^ n[16593];
assign t[16594] = t[16593] ^ n[16594];
assign t[16595] = t[16594] ^ n[16595];
assign t[16596] = t[16595] ^ n[16596];
assign t[16597] = t[16596] ^ n[16597];
assign t[16598] = t[16597] ^ n[16598];
assign t[16599] = t[16598] ^ n[16599];
assign t[16600] = t[16599] ^ n[16600];
assign t[16601] = t[16600] ^ n[16601];
assign t[16602] = t[16601] ^ n[16602];
assign t[16603] = t[16602] ^ n[16603];
assign t[16604] = t[16603] ^ n[16604];
assign t[16605] = t[16604] ^ n[16605];
assign t[16606] = t[16605] ^ n[16606];
assign t[16607] = t[16606] ^ n[16607];
assign t[16608] = t[16607] ^ n[16608];
assign t[16609] = t[16608] ^ n[16609];
assign t[16610] = t[16609] ^ n[16610];
assign t[16611] = t[16610] ^ n[16611];
assign t[16612] = t[16611] ^ n[16612];
assign t[16613] = t[16612] ^ n[16613];
assign t[16614] = t[16613] ^ n[16614];
assign t[16615] = t[16614] ^ n[16615];
assign t[16616] = t[16615] ^ n[16616];
assign t[16617] = t[16616] ^ n[16617];
assign t[16618] = t[16617] ^ n[16618];
assign t[16619] = t[16618] ^ n[16619];
assign t[16620] = t[16619] ^ n[16620];
assign t[16621] = t[16620] ^ n[16621];
assign t[16622] = t[16621] ^ n[16622];
assign t[16623] = t[16622] ^ n[16623];
assign t[16624] = t[16623] ^ n[16624];
assign t[16625] = t[16624] ^ n[16625];
assign t[16626] = t[16625] ^ n[16626];
assign t[16627] = t[16626] ^ n[16627];
assign t[16628] = t[16627] ^ n[16628];
assign t[16629] = t[16628] ^ n[16629];
assign t[16630] = t[16629] ^ n[16630];
assign t[16631] = t[16630] ^ n[16631];
assign t[16632] = t[16631] ^ n[16632];
assign t[16633] = t[16632] ^ n[16633];
assign t[16634] = t[16633] ^ n[16634];
assign t[16635] = t[16634] ^ n[16635];
assign t[16636] = t[16635] ^ n[16636];
assign t[16637] = t[16636] ^ n[16637];
assign t[16638] = t[16637] ^ n[16638];
assign t[16639] = t[16638] ^ n[16639];
assign t[16640] = t[16639] ^ n[16640];
assign t[16641] = t[16640] ^ n[16641];
assign t[16642] = t[16641] ^ n[16642];
assign t[16643] = t[16642] ^ n[16643];
assign t[16644] = t[16643] ^ n[16644];
assign t[16645] = t[16644] ^ n[16645];
assign t[16646] = t[16645] ^ n[16646];
assign t[16647] = t[16646] ^ n[16647];
assign t[16648] = t[16647] ^ n[16648];
assign t[16649] = t[16648] ^ n[16649];
assign t[16650] = t[16649] ^ n[16650];
assign t[16651] = t[16650] ^ n[16651];
assign t[16652] = t[16651] ^ n[16652];
assign t[16653] = t[16652] ^ n[16653];
assign t[16654] = t[16653] ^ n[16654];
assign t[16655] = t[16654] ^ n[16655];
assign t[16656] = t[16655] ^ n[16656];
assign t[16657] = t[16656] ^ n[16657];
assign t[16658] = t[16657] ^ n[16658];
assign t[16659] = t[16658] ^ n[16659];
assign t[16660] = t[16659] ^ n[16660];
assign t[16661] = t[16660] ^ n[16661];
assign t[16662] = t[16661] ^ n[16662];
assign t[16663] = t[16662] ^ n[16663];
assign t[16664] = t[16663] ^ n[16664];
assign t[16665] = t[16664] ^ n[16665];
assign t[16666] = t[16665] ^ n[16666];
assign t[16667] = t[16666] ^ n[16667];
assign t[16668] = t[16667] ^ n[16668];
assign t[16669] = t[16668] ^ n[16669];
assign t[16670] = t[16669] ^ n[16670];
assign t[16671] = t[16670] ^ n[16671];
assign t[16672] = t[16671] ^ n[16672];
assign t[16673] = t[16672] ^ n[16673];
assign t[16674] = t[16673] ^ n[16674];
assign t[16675] = t[16674] ^ n[16675];
assign t[16676] = t[16675] ^ n[16676];
assign t[16677] = t[16676] ^ n[16677];
assign t[16678] = t[16677] ^ n[16678];
assign t[16679] = t[16678] ^ n[16679];
assign t[16680] = t[16679] ^ n[16680];
assign t[16681] = t[16680] ^ n[16681];
assign t[16682] = t[16681] ^ n[16682];
assign t[16683] = t[16682] ^ n[16683];
assign t[16684] = t[16683] ^ n[16684];
assign t[16685] = t[16684] ^ n[16685];
assign t[16686] = t[16685] ^ n[16686];
assign t[16687] = t[16686] ^ n[16687];
assign t[16688] = t[16687] ^ n[16688];
assign t[16689] = t[16688] ^ n[16689];
assign t[16690] = t[16689] ^ n[16690];
assign t[16691] = t[16690] ^ n[16691];
assign t[16692] = t[16691] ^ n[16692];
assign t[16693] = t[16692] ^ n[16693];
assign t[16694] = t[16693] ^ n[16694];
assign t[16695] = t[16694] ^ n[16695];
assign t[16696] = t[16695] ^ n[16696];
assign t[16697] = t[16696] ^ n[16697];
assign t[16698] = t[16697] ^ n[16698];
assign t[16699] = t[16698] ^ n[16699];
assign t[16700] = t[16699] ^ n[16700];
assign t[16701] = t[16700] ^ n[16701];
assign t[16702] = t[16701] ^ n[16702];
assign t[16703] = t[16702] ^ n[16703];
assign t[16704] = t[16703] ^ n[16704];
assign t[16705] = t[16704] ^ n[16705];
assign t[16706] = t[16705] ^ n[16706];
assign t[16707] = t[16706] ^ n[16707];
assign t[16708] = t[16707] ^ n[16708];
assign t[16709] = t[16708] ^ n[16709];
assign t[16710] = t[16709] ^ n[16710];
assign t[16711] = t[16710] ^ n[16711];
assign t[16712] = t[16711] ^ n[16712];
assign t[16713] = t[16712] ^ n[16713];
assign t[16714] = t[16713] ^ n[16714];
assign t[16715] = t[16714] ^ n[16715];
assign t[16716] = t[16715] ^ n[16716];
assign t[16717] = t[16716] ^ n[16717];
assign t[16718] = t[16717] ^ n[16718];
assign t[16719] = t[16718] ^ n[16719];
assign t[16720] = t[16719] ^ n[16720];
assign t[16721] = t[16720] ^ n[16721];
assign t[16722] = t[16721] ^ n[16722];
assign t[16723] = t[16722] ^ n[16723];
assign t[16724] = t[16723] ^ n[16724];
assign t[16725] = t[16724] ^ n[16725];
assign t[16726] = t[16725] ^ n[16726];
assign t[16727] = t[16726] ^ n[16727];
assign t[16728] = t[16727] ^ n[16728];
assign t[16729] = t[16728] ^ n[16729];
assign t[16730] = t[16729] ^ n[16730];
assign t[16731] = t[16730] ^ n[16731];
assign t[16732] = t[16731] ^ n[16732];
assign t[16733] = t[16732] ^ n[16733];
assign t[16734] = t[16733] ^ n[16734];
assign t[16735] = t[16734] ^ n[16735];
assign t[16736] = t[16735] ^ n[16736];
assign t[16737] = t[16736] ^ n[16737];
assign t[16738] = t[16737] ^ n[16738];
assign t[16739] = t[16738] ^ n[16739];
assign t[16740] = t[16739] ^ n[16740];
assign t[16741] = t[16740] ^ n[16741];
assign t[16742] = t[16741] ^ n[16742];
assign t[16743] = t[16742] ^ n[16743];
assign t[16744] = t[16743] ^ n[16744];
assign t[16745] = t[16744] ^ n[16745];
assign t[16746] = t[16745] ^ n[16746];
assign t[16747] = t[16746] ^ n[16747];
assign t[16748] = t[16747] ^ n[16748];
assign t[16749] = t[16748] ^ n[16749];
assign t[16750] = t[16749] ^ n[16750];
assign t[16751] = t[16750] ^ n[16751];
assign t[16752] = t[16751] ^ n[16752];
assign t[16753] = t[16752] ^ n[16753];
assign t[16754] = t[16753] ^ n[16754];
assign t[16755] = t[16754] ^ n[16755];
assign t[16756] = t[16755] ^ n[16756];
assign t[16757] = t[16756] ^ n[16757];
assign t[16758] = t[16757] ^ n[16758];
assign t[16759] = t[16758] ^ n[16759];
assign t[16760] = t[16759] ^ n[16760];
assign t[16761] = t[16760] ^ n[16761];
assign t[16762] = t[16761] ^ n[16762];
assign t[16763] = t[16762] ^ n[16763];
assign t[16764] = t[16763] ^ n[16764];
assign t[16765] = t[16764] ^ n[16765];
assign t[16766] = t[16765] ^ n[16766];
assign t[16767] = t[16766] ^ n[16767];
assign t[16768] = t[16767] ^ n[16768];
assign t[16769] = t[16768] ^ n[16769];
assign t[16770] = t[16769] ^ n[16770];
assign t[16771] = t[16770] ^ n[16771];
assign t[16772] = t[16771] ^ n[16772];
assign t[16773] = t[16772] ^ n[16773];
assign t[16774] = t[16773] ^ n[16774];
assign t[16775] = t[16774] ^ n[16775];
assign t[16776] = t[16775] ^ n[16776];
assign t[16777] = t[16776] ^ n[16777];
assign t[16778] = t[16777] ^ n[16778];
assign t[16779] = t[16778] ^ n[16779];
assign t[16780] = t[16779] ^ n[16780];
assign t[16781] = t[16780] ^ n[16781];
assign t[16782] = t[16781] ^ n[16782];
assign t[16783] = t[16782] ^ n[16783];
assign t[16784] = t[16783] ^ n[16784];
assign t[16785] = t[16784] ^ n[16785];
assign t[16786] = t[16785] ^ n[16786];
assign t[16787] = t[16786] ^ n[16787];
assign t[16788] = t[16787] ^ n[16788];
assign t[16789] = t[16788] ^ n[16789];
assign t[16790] = t[16789] ^ n[16790];
assign t[16791] = t[16790] ^ n[16791];
assign t[16792] = t[16791] ^ n[16792];
assign t[16793] = t[16792] ^ n[16793];
assign t[16794] = t[16793] ^ n[16794];
assign t[16795] = t[16794] ^ n[16795];
assign t[16796] = t[16795] ^ n[16796];
assign t[16797] = t[16796] ^ n[16797];
assign t[16798] = t[16797] ^ n[16798];
assign t[16799] = t[16798] ^ n[16799];
assign t[16800] = t[16799] ^ n[16800];
assign t[16801] = t[16800] ^ n[16801];
assign t[16802] = t[16801] ^ n[16802];
assign t[16803] = t[16802] ^ n[16803];
assign t[16804] = t[16803] ^ n[16804];
assign t[16805] = t[16804] ^ n[16805];
assign t[16806] = t[16805] ^ n[16806];
assign t[16807] = t[16806] ^ n[16807];
assign t[16808] = t[16807] ^ n[16808];
assign t[16809] = t[16808] ^ n[16809];
assign t[16810] = t[16809] ^ n[16810];
assign t[16811] = t[16810] ^ n[16811];
assign t[16812] = t[16811] ^ n[16812];
assign t[16813] = t[16812] ^ n[16813];
assign t[16814] = t[16813] ^ n[16814];
assign t[16815] = t[16814] ^ n[16815];
assign t[16816] = t[16815] ^ n[16816];
assign t[16817] = t[16816] ^ n[16817];
assign t[16818] = t[16817] ^ n[16818];
assign t[16819] = t[16818] ^ n[16819];
assign t[16820] = t[16819] ^ n[16820];
assign t[16821] = t[16820] ^ n[16821];
assign t[16822] = t[16821] ^ n[16822];
assign t[16823] = t[16822] ^ n[16823];
assign t[16824] = t[16823] ^ n[16824];
assign t[16825] = t[16824] ^ n[16825];
assign t[16826] = t[16825] ^ n[16826];
assign t[16827] = t[16826] ^ n[16827];
assign t[16828] = t[16827] ^ n[16828];
assign t[16829] = t[16828] ^ n[16829];
assign t[16830] = t[16829] ^ n[16830];
assign t[16831] = t[16830] ^ n[16831];
assign t[16832] = t[16831] ^ n[16832];
assign t[16833] = t[16832] ^ n[16833];
assign t[16834] = t[16833] ^ n[16834];
assign t[16835] = t[16834] ^ n[16835];
assign t[16836] = t[16835] ^ n[16836];
assign t[16837] = t[16836] ^ n[16837];
assign t[16838] = t[16837] ^ n[16838];
assign t[16839] = t[16838] ^ n[16839];
assign t[16840] = t[16839] ^ n[16840];
assign t[16841] = t[16840] ^ n[16841];
assign t[16842] = t[16841] ^ n[16842];
assign t[16843] = t[16842] ^ n[16843];
assign t[16844] = t[16843] ^ n[16844];
assign t[16845] = t[16844] ^ n[16845];
assign t[16846] = t[16845] ^ n[16846];
assign t[16847] = t[16846] ^ n[16847];
assign t[16848] = t[16847] ^ n[16848];
assign t[16849] = t[16848] ^ n[16849];
assign t[16850] = t[16849] ^ n[16850];
assign t[16851] = t[16850] ^ n[16851];
assign t[16852] = t[16851] ^ n[16852];
assign t[16853] = t[16852] ^ n[16853];
assign t[16854] = t[16853] ^ n[16854];
assign t[16855] = t[16854] ^ n[16855];
assign t[16856] = t[16855] ^ n[16856];
assign t[16857] = t[16856] ^ n[16857];
assign t[16858] = t[16857] ^ n[16858];
assign t[16859] = t[16858] ^ n[16859];
assign t[16860] = t[16859] ^ n[16860];
assign t[16861] = t[16860] ^ n[16861];
assign t[16862] = t[16861] ^ n[16862];
assign t[16863] = t[16862] ^ n[16863];
assign t[16864] = t[16863] ^ n[16864];
assign t[16865] = t[16864] ^ n[16865];
assign t[16866] = t[16865] ^ n[16866];
assign t[16867] = t[16866] ^ n[16867];
assign t[16868] = t[16867] ^ n[16868];
assign t[16869] = t[16868] ^ n[16869];
assign t[16870] = t[16869] ^ n[16870];
assign t[16871] = t[16870] ^ n[16871];
assign t[16872] = t[16871] ^ n[16872];
assign t[16873] = t[16872] ^ n[16873];
assign t[16874] = t[16873] ^ n[16874];
assign t[16875] = t[16874] ^ n[16875];
assign t[16876] = t[16875] ^ n[16876];
assign t[16877] = t[16876] ^ n[16877];
assign t[16878] = t[16877] ^ n[16878];
assign t[16879] = t[16878] ^ n[16879];
assign t[16880] = t[16879] ^ n[16880];
assign t[16881] = t[16880] ^ n[16881];
assign t[16882] = t[16881] ^ n[16882];
assign t[16883] = t[16882] ^ n[16883];
assign t[16884] = t[16883] ^ n[16884];
assign t[16885] = t[16884] ^ n[16885];
assign t[16886] = t[16885] ^ n[16886];
assign t[16887] = t[16886] ^ n[16887];
assign t[16888] = t[16887] ^ n[16888];
assign t[16889] = t[16888] ^ n[16889];
assign t[16890] = t[16889] ^ n[16890];
assign t[16891] = t[16890] ^ n[16891];
assign t[16892] = t[16891] ^ n[16892];
assign t[16893] = t[16892] ^ n[16893];
assign t[16894] = t[16893] ^ n[16894];
assign t[16895] = t[16894] ^ n[16895];
assign t[16896] = t[16895] ^ n[16896];
assign t[16897] = t[16896] ^ n[16897];
assign t[16898] = t[16897] ^ n[16898];
assign t[16899] = t[16898] ^ n[16899];
assign t[16900] = t[16899] ^ n[16900];
assign t[16901] = t[16900] ^ n[16901];
assign t[16902] = t[16901] ^ n[16902];
assign t[16903] = t[16902] ^ n[16903];
assign t[16904] = t[16903] ^ n[16904];
assign t[16905] = t[16904] ^ n[16905];
assign t[16906] = t[16905] ^ n[16906];
assign t[16907] = t[16906] ^ n[16907];
assign t[16908] = t[16907] ^ n[16908];
assign t[16909] = t[16908] ^ n[16909];
assign t[16910] = t[16909] ^ n[16910];
assign t[16911] = t[16910] ^ n[16911];
assign t[16912] = t[16911] ^ n[16912];
assign t[16913] = t[16912] ^ n[16913];
assign t[16914] = t[16913] ^ n[16914];
assign t[16915] = t[16914] ^ n[16915];
assign t[16916] = t[16915] ^ n[16916];
assign t[16917] = t[16916] ^ n[16917];
assign t[16918] = t[16917] ^ n[16918];
assign t[16919] = t[16918] ^ n[16919];
assign t[16920] = t[16919] ^ n[16920];
assign t[16921] = t[16920] ^ n[16921];
assign t[16922] = t[16921] ^ n[16922];
assign t[16923] = t[16922] ^ n[16923];
assign t[16924] = t[16923] ^ n[16924];
assign t[16925] = t[16924] ^ n[16925];
assign t[16926] = t[16925] ^ n[16926];
assign t[16927] = t[16926] ^ n[16927];
assign t[16928] = t[16927] ^ n[16928];
assign t[16929] = t[16928] ^ n[16929];
assign t[16930] = t[16929] ^ n[16930];
assign t[16931] = t[16930] ^ n[16931];
assign t[16932] = t[16931] ^ n[16932];
assign t[16933] = t[16932] ^ n[16933];
assign t[16934] = t[16933] ^ n[16934];
assign t[16935] = t[16934] ^ n[16935];
assign t[16936] = t[16935] ^ n[16936];
assign t[16937] = t[16936] ^ n[16937];
assign t[16938] = t[16937] ^ n[16938];
assign t[16939] = t[16938] ^ n[16939];
assign t[16940] = t[16939] ^ n[16940];
assign t[16941] = t[16940] ^ n[16941];
assign t[16942] = t[16941] ^ n[16942];
assign t[16943] = t[16942] ^ n[16943];
assign t[16944] = t[16943] ^ n[16944];
assign t[16945] = t[16944] ^ n[16945];
assign t[16946] = t[16945] ^ n[16946];
assign t[16947] = t[16946] ^ n[16947];
assign t[16948] = t[16947] ^ n[16948];
assign t[16949] = t[16948] ^ n[16949];
assign t[16950] = t[16949] ^ n[16950];
assign t[16951] = t[16950] ^ n[16951];
assign t[16952] = t[16951] ^ n[16952];
assign t[16953] = t[16952] ^ n[16953];
assign t[16954] = t[16953] ^ n[16954];
assign t[16955] = t[16954] ^ n[16955];
assign t[16956] = t[16955] ^ n[16956];
assign t[16957] = t[16956] ^ n[16957];
assign t[16958] = t[16957] ^ n[16958];
assign t[16959] = t[16958] ^ n[16959];
assign t[16960] = t[16959] ^ n[16960];
assign t[16961] = t[16960] ^ n[16961];
assign t[16962] = t[16961] ^ n[16962];
assign t[16963] = t[16962] ^ n[16963];
assign t[16964] = t[16963] ^ n[16964];
assign t[16965] = t[16964] ^ n[16965];
assign t[16966] = t[16965] ^ n[16966];
assign t[16967] = t[16966] ^ n[16967];
assign t[16968] = t[16967] ^ n[16968];
assign t[16969] = t[16968] ^ n[16969];
assign t[16970] = t[16969] ^ n[16970];
assign t[16971] = t[16970] ^ n[16971];
assign t[16972] = t[16971] ^ n[16972];
assign t[16973] = t[16972] ^ n[16973];
assign t[16974] = t[16973] ^ n[16974];
assign t[16975] = t[16974] ^ n[16975];
assign t[16976] = t[16975] ^ n[16976];
assign t[16977] = t[16976] ^ n[16977];
assign t[16978] = t[16977] ^ n[16978];
assign t[16979] = t[16978] ^ n[16979];
assign t[16980] = t[16979] ^ n[16980];
assign t[16981] = t[16980] ^ n[16981];
assign t[16982] = t[16981] ^ n[16982];
assign t[16983] = t[16982] ^ n[16983];
assign t[16984] = t[16983] ^ n[16984];
assign t[16985] = t[16984] ^ n[16985];
assign t[16986] = t[16985] ^ n[16986];
assign t[16987] = t[16986] ^ n[16987];
assign t[16988] = t[16987] ^ n[16988];
assign t[16989] = t[16988] ^ n[16989];
assign t[16990] = t[16989] ^ n[16990];
assign t[16991] = t[16990] ^ n[16991];
assign t[16992] = t[16991] ^ n[16992];
assign t[16993] = t[16992] ^ n[16993];
assign t[16994] = t[16993] ^ n[16994];
assign t[16995] = t[16994] ^ n[16995];
assign t[16996] = t[16995] ^ n[16996];
assign t[16997] = t[16996] ^ n[16997];
assign t[16998] = t[16997] ^ n[16998];
assign t[16999] = t[16998] ^ n[16999];
assign t[17000] = t[16999] ^ n[17000];
assign t[17001] = t[17000] ^ n[17001];
assign t[17002] = t[17001] ^ n[17002];
assign t[17003] = t[17002] ^ n[17003];
assign t[17004] = t[17003] ^ n[17004];
assign t[17005] = t[17004] ^ n[17005];
assign t[17006] = t[17005] ^ n[17006];
assign t[17007] = t[17006] ^ n[17007];
assign t[17008] = t[17007] ^ n[17008];
assign t[17009] = t[17008] ^ n[17009];
assign t[17010] = t[17009] ^ n[17010];
assign t[17011] = t[17010] ^ n[17011];
assign t[17012] = t[17011] ^ n[17012];
assign t[17013] = t[17012] ^ n[17013];
assign t[17014] = t[17013] ^ n[17014];
assign t[17015] = t[17014] ^ n[17015];
assign t[17016] = t[17015] ^ n[17016];
assign t[17017] = t[17016] ^ n[17017];
assign t[17018] = t[17017] ^ n[17018];
assign t[17019] = t[17018] ^ n[17019];
assign t[17020] = t[17019] ^ n[17020];
assign t[17021] = t[17020] ^ n[17021];
assign t[17022] = t[17021] ^ n[17022];
assign t[17023] = t[17022] ^ n[17023];
assign t[17024] = t[17023] ^ n[17024];
assign t[17025] = t[17024] ^ n[17025];
assign t[17026] = t[17025] ^ n[17026];
assign t[17027] = t[17026] ^ n[17027];
assign t[17028] = t[17027] ^ n[17028];
assign t[17029] = t[17028] ^ n[17029];
assign t[17030] = t[17029] ^ n[17030];
assign t[17031] = t[17030] ^ n[17031];
assign t[17032] = t[17031] ^ n[17032];
assign t[17033] = t[17032] ^ n[17033];
assign t[17034] = t[17033] ^ n[17034];
assign t[17035] = t[17034] ^ n[17035];
assign t[17036] = t[17035] ^ n[17036];
assign t[17037] = t[17036] ^ n[17037];
assign t[17038] = t[17037] ^ n[17038];
assign t[17039] = t[17038] ^ n[17039];
assign t[17040] = t[17039] ^ n[17040];
assign t[17041] = t[17040] ^ n[17041];
assign t[17042] = t[17041] ^ n[17042];
assign t[17043] = t[17042] ^ n[17043];
assign t[17044] = t[17043] ^ n[17044];
assign t[17045] = t[17044] ^ n[17045];
assign t[17046] = t[17045] ^ n[17046];
assign t[17047] = t[17046] ^ n[17047];
assign t[17048] = t[17047] ^ n[17048];
assign t[17049] = t[17048] ^ n[17049];
assign t[17050] = t[17049] ^ n[17050];
assign t[17051] = t[17050] ^ n[17051];
assign t[17052] = t[17051] ^ n[17052];
assign t[17053] = t[17052] ^ n[17053];
assign t[17054] = t[17053] ^ n[17054];
assign t[17055] = t[17054] ^ n[17055];
assign t[17056] = t[17055] ^ n[17056];
assign t[17057] = t[17056] ^ n[17057];
assign t[17058] = t[17057] ^ n[17058];
assign t[17059] = t[17058] ^ n[17059];
assign t[17060] = t[17059] ^ n[17060];
assign t[17061] = t[17060] ^ n[17061];
assign t[17062] = t[17061] ^ n[17062];
assign t[17063] = t[17062] ^ n[17063];
assign t[17064] = t[17063] ^ n[17064];
assign t[17065] = t[17064] ^ n[17065];
assign t[17066] = t[17065] ^ n[17066];
assign t[17067] = t[17066] ^ n[17067];
assign t[17068] = t[17067] ^ n[17068];
assign t[17069] = t[17068] ^ n[17069];
assign t[17070] = t[17069] ^ n[17070];
assign t[17071] = t[17070] ^ n[17071];
assign t[17072] = t[17071] ^ n[17072];
assign t[17073] = t[17072] ^ n[17073];
assign t[17074] = t[17073] ^ n[17074];
assign t[17075] = t[17074] ^ n[17075];
assign t[17076] = t[17075] ^ n[17076];
assign t[17077] = t[17076] ^ n[17077];
assign t[17078] = t[17077] ^ n[17078];
assign t[17079] = t[17078] ^ n[17079];
assign t[17080] = t[17079] ^ n[17080];
assign t[17081] = t[17080] ^ n[17081];
assign t[17082] = t[17081] ^ n[17082];
assign t[17083] = t[17082] ^ n[17083];
assign t[17084] = t[17083] ^ n[17084];
assign t[17085] = t[17084] ^ n[17085];
assign t[17086] = t[17085] ^ n[17086];
assign t[17087] = t[17086] ^ n[17087];
assign t[17088] = t[17087] ^ n[17088];
assign t[17089] = t[17088] ^ n[17089];
assign t[17090] = t[17089] ^ n[17090];
assign t[17091] = t[17090] ^ n[17091];
assign t[17092] = t[17091] ^ n[17092];
assign t[17093] = t[17092] ^ n[17093];
assign t[17094] = t[17093] ^ n[17094];
assign t[17095] = t[17094] ^ n[17095];
assign t[17096] = t[17095] ^ n[17096];
assign t[17097] = t[17096] ^ n[17097];
assign t[17098] = t[17097] ^ n[17098];
assign t[17099] = t[17098] ^ n[17099];
assign t[17100] = t[17099] ^ n[17100];
assign t[17101] = t[17100] ^ n[17101];
assign t[17102] = t[17101] ^ n[17102];
assign t[17103] = t[17102] ^ n[17103];
assign t[17104] = t[17103] ^ n[17104];
assign t[17105] = t[17104] ^ n[17105];
assign t[17106] = t[17105] ^ n[17106];
assign t[17107] = t[17106] ^ n[17107];
assign t[17108] = t[17107] ^ n[17108];
assign t[17109] = t[17108] ^ n[17109];
assign t[17110] = t[17109] ^ n[17110];
assign t[17111] = t[17110] ^ n[17111];
assign t[17112] = t[17111] ^ n[17112];
assign t[17113] = t[17112] ^ n[17113];
assign t[17114] = t[17113] ^ n[17114];
assign t[17115] = t[17114] ^ n[17115];
assign t[17116] = t[17115] ^ n[17116];
assign t[17117] = t[17116] ^ n[17117];
assign t[17118] = t[17117] ^ n[17118];
assign t[17119] = t[17118] ^ n[17119];
assign t[17120] = t[17119] ^ n[17120];
assign t[17121] = t[17120] ^ n[17121];
assign t[17122] = t[17121] ^ n[17122];
assign t[17123] = t[17122] ^ n[17123];
assign t[17124] = t[17123] ^ n[17124];
assign t[17125] = t[17124] ^ n[17125];
assign t[17126] = t[17125] ^ n[17126];
assign t[17127] = t[17126] ^ n[17127];
assign t[17128] = t[17127] ^ n[17128];
assign t[17129] = t[17128] ^ n[17129];
assign t[17130] = t[17129] ^ n[17130];
assign t[17131] = t[17130] ^ n[17131];
assign t[17132] = t[17131] ^ n[17132];
assign t[17133] = t[17132] ^ n[17133];
assign t[17134] = t[17133] ^ n[17134];
assign t[17135] = t[17134] ^ n[17135];
assign t[17136] = t[17135] ^ n[17136];
assign t[17137] = t[17136] ^ n[17137];
assign t[17138] = t[17137] ^ n[17138];
assign t[17139] = t[17138] ^ n[17139];
assign t[17140] = t[17139] ^ n[17140];
assign t[17141] = t[17140] ^ n[17141];
assign t[17142] = t[17141] ^ n[17142];
assign t[17143] = t[17142] ^ n[17143];
assign t[17144] = t[17143] ^ n[17144];
assign t[17145] = t[17144] ^ n[17145];
assign t[17146] = t[17145] ^ n[17146];
assign t[17147] = t[17146] ^ n[17147];
assign t[17148] = t[17147] ^ n[17148];
assign t[17149] = t[17148] ^ n[17149];
assign t[17150] = t[17149] ^ n[17150];
assign t[17151] = t[17150] ^ n[17151];
assign t[17152] = t[17151] ^ n[17152];
assign t[17153] = t[17152] ^ n[17153];
assign t[17154] = t[17153] ^ n[17154];
assign t[17155] = t[17154] ^ n[17155];
assign t[17156] = t[17155] ^ n[17156];
assign t[17157] = t[17156] ^ n[17157];
assign t[17158] = t[17157] ^ n[17158];
assign t[17159] = t[17158] ^ n[17159];
assign t[17160] = t[17159] ^ n[17160];
assign t[17161] = t[17160] ^ n[17161];
assign t[17162] = t[17161] ^ n[17162];
assign t[17163] = t[17162] ^ n[17163];
assign t[17164] = t[17163] ^ n[17164];
assign t[17165] = t[17164] ^ n[17165];
assign t[17166] = t[17165] ^ n[17166];
assign t[17167] = t[17166] ^ n[17167];
assign t[17168] = t[17167] ^ n[17168];
assign t[17169] = t[17168] ^ n[17169];
assign t[17170] = t[17169] ^ n[17170];
assign t[17171] = t[17170] ^ n[17171];
assign t[17172] = t[17171] ^ n[17172];
assign t[17173] = t[17172] ^ n[17173];
assign t[17174] = t[17173] ^ n[17174];
assign t[17175] = t[17174] ^ n[17175];
assign t[17176] = t[17175] ^ n[17176];
assign t[17177] = t[17176] ^ n[17177];
assign t[17178] = t[17177] ^ n[17178];
assign t[17179] = t[17178] ^ n[17179];
assign t[17180] = t[17179] ^ n[17180];
assign t[17181] = t[17180] ^ n[17181];
assign t[17182] = t[17181] ^ n[17182];
assign t[17183] = t[17182] ^ n[17183];
assign t[17184] = t[17183] ^ n[17184];
assign t[17185] = t[17184] ^ n[17185];
assign t[17186] = t[17185] ^ n[17186];
assign t[17187] = t[17186] ^ n[17187];
assign t[17188] = t[17187] ^ n[17188];
assign t[17189] = t[17188] ^ n[17189];
assign t[17190] = t[17189] ^ n[17190];
assign t[17191] = t[17190] ^ n[17191];
assign t[17192] = t[17191] ^ n[17192];
assign t[17193] = t[17192] ^ n[17193];
assign t[17194] = t[17193] ^ n[17194];
assign t[17195] = t[17194] ^ n[17195];
assign t[17196] = t[17195] ^ n[17196];
assign t[17197] = t[17196] ^ n[17197];
assign t[17198] = t[17197] ^ n[17198];
assign t[17199] = t[17198] ^ n[17199];
assign t[17200] = t[17199] ^ n[17200];
assign t[17201] = t[17200] ^ n[17201];
assign t[17202] = t[17201] ^ n[17202];
assign t[17203] = t[17202] ^ n[17203];
assign t[17204] = t[17203] ^ n[17204];
assign t[17205] = t[17204] ^ n[17205];
assign t[17206] = t[17205] ^ n[17206];
assign t[17207] = t[17206] ^ n[17207];
assign t[17208] = t[17207] ^ n[17208];
assign t[17209] = t[17208] ^ n[17209];
assign t[17210] = t[17209] ^ n[17210];
assign t[17211] = t[17210] ^ n[17211];
assign t[17212] = t[17211] ^ n[17212];
assign t[17213] = t[17212] ^ n[17213];
assign t[17214] = t[17213] ^ n[17214];
assign t[17215] = t[17214] ^ n[17215];
assign t[17216] = t[17215] ^ n[17216];
assign t[17217] = t[17216] ^ n[17217];
assign t[17218] = t[17217] ^ n[17218];
assign t[17219] = t[17218] ^ n[17219];
assign t[17220] = t[17219] ^ n[17220];
assign t[17221] = t[17220] ^ n[17221];
assign t[17222] = t[17221] ^ n[17222];
assign t[17223] = t[17222] ^ n[17223];
assign t[17224] = t[17223] ^ n[17224];
assign t[17225] = t[17224] ^ n[17225];
assign t[17226] = t[17225] ^ n[17226];
assign t[17227] = t[17226] ^ n[17227];
assign t[17228] = t[17227] ^ n[17228];
assign t[17229] = t[17228] ^ n[17229];
assign t[17230] = t[17229] ^ n[17230];
assign t[17231] = t[17230] ^ n[17231];
assign t[17232] = t[17231] ^ n[17232];
assign t[17233] = t[17232] ^ n[17233];
assign t[17234] = t[17233] ^ n[17234];
assign t[17235] = t[17234] ^ n[17235];
assign t[17236] = t[17235] ^ n[17236];
assign t[17237] = t[17236] ^ n[17237];
assign t[17238] = t[17237] ^ n[17238];
assign t[17239] = t[17238] ^ n[17239];
assign t[17240] = t[17239] ^ n[17240];
assign t[17241] = t[17240] ^ n[17241];
assign t[17242] = t[17241] ^ n[17242];
assign t[17243] = t[17242] ^ n[17243];
assign t[17244] = t[17243] ^ n[17244];
assign t[17245] = t[17244] ^ n[17245];
assign t[17246] = t[17245] ^ n[17246];
assign t[17247] = t[17246] ^ n[17247];
assign t[17248] = t[17247] ^ n[17248];
assign t[17249] = t[17248] ^ n[17249];
assign t[17250] = t[17249] ^ n[17250];
assign t[17251] = t[17250] ^ n[17251];
assign t[17252] = t[17251] ^ n[17252];
assign t[17253] = t[17252] ^ n[17253];
assign t[17254] = t[17253] ^ n[17254];
assign t[17255] = t[17254] ^ n[17255];
assign t[17256] = t[17255] ^ n[17256];
assign t[17257] = t[17256] ^ n[17257];
assign t[17258] = t[17257] ^ n[17258];
assign t[17259] = t[17258] ^ n[17259];
assign t[17260] = t[17259] ^ n[17260];
assign t[17261] = t[17260] ^ n[17261];
assign t[17262] = t[17261] ^ n[17262];
assign t[17263] = t[17262] ^ n[17263];
assign t[17264] = t[17263] ^ n[17264];
assign t[17265] = t[17264] ^ n[17265];
assign t[17266] = t[17265] ^ n[17266];
assign t[17267] = t[17266] ^ n[17267];
assign t[17268] = t[17267] ^ n[17268];
assign t[17269] = t[17268] ^ n[17269];
assign t[17270] = t[17269] ^ n[17270];
assign t[17271] = t[17270] ^ n[17271];
assign t[17272] = t[17271] ^ n[17272];
assign t[17273] = t[17272] ^ n[17273];
assign t[17274] = t[17273] ^ n[17274];
assign t[17275] = t[17274] ^ n[17275];
assign t[17276] = t[17275] ^ n[17276];
assign t[17277] = t[17276] ^ n[17277];
assign t[17278] = t[17277] ^ n[17278];
assign t[17279] = t[17278] ^ n[17279];
assign t[17280] = t[17279] ^ n[17280];
assign t[17281] = t[17280] ^ n[17281];
assign t[17282] = t[17281] ^ n[17282];
assign t[17283] = t[17282] ^ n[17283];
assign t[17284] = t[17283] ^ n[17284];
assign t[17285] = t[17284] ^ n[17285];
assign t[17286] = t[17285] ^ n[17286];
assign t[17287] = t[17286] ^ n[17287];
assign t[17288] = t[17287] ^ n[17288];
assign t[17289] = t[17288] ^ n[17289];
assign t[17290] = t[17289] ^ n[17290];
assign t[17291] = t[17290] ^ n[17291];
assign t[17292] = t[17291] ^ n[17292];
assign t[17293] = t[17292] ^ n[17293];
assign t[17294] = t[17293] ^ n[17294];
assign t[17295] = t[17294] ^ n[17295];
assign t[17296] = t[17295] ^ n[17296];
assign t[17297] = t[17296] ^ n[17297];
assign t[17298] = t[17297] ^ n[17298];
assign t[17299] = t[17298] ^ n[17299];
assign t[17300] = t[17299] ^ n[17300];
assign t[17301] = t[17300] ^ n[17301];
assign t[17302] = t[17301] ^ n[17302];
assign t[17303] = t[17302] ^ n[17303];
assign t[17304] = t[17303] ^ n[17304];
assign t[17305] = t[17304] ^ n[17305];
assign t[17306] = t[17305] ^ n[17306];
assign t[17307] = t[17306] ^ n[17307];
assign t[17308] = t[17307] ^ n[17308];
assign t[17309] = t[17308] ^ n[17309];
assign t[17310] = t[17309] ^ n[17310];
assign t[17311] = t[17310] ^ n[17311];
assign t[17312] = t[17311] ^ n[17312];
assign t[17313] = t[17312] ^ n[17313];
assign t[17314] = t[17313] ^ n[17314];
assign t[17315] = t[17314] ^ n[17315];
assign t[17316] = t[17315] ^ n[17316];
assign t[17317] = t[17316] ^ n[17317];
assign t[17318] = t[17317] ^ n[17318];
assign t[17319] = t[17318] ^ n[17319];
assign t[17320] = t[17319] ^ n[17320];
assign t[17321] = t[17320] ^ n[17321];
assign t[17322] = t[17321] ^ n[17322];
assign t[17323] = t[17322] ^ n[17323];
assign t[17324] = t[17323] ^ n[17324];
assign t[17325] = t[17324] ^ n[17325];
assign t[17326] = t[17325] ^ n[17326];
assign t[17327] = t[17326] ^ n[17327];
assign t[17328] = t[17327] ^ n[17328];
assign t[17329] = t[17328] ^ n[17329];
assign t[17330] = t[17329] ^ n[17330];
assign t[17331] = t[17330] ^ n[17331];
assign t[17332] = t[17331] ^ n[17332];
assign t[17333] = t[17332] ^ n[17333];
assign t[17334] = t[17333] ^ n[17334];
assign t[17335] = t[17334] ^ n[17335];
assign t[17336] = t[17335] ^ n[17336];
assign t[17337] = t[17336] ^ n[17337];
assign t[17338] = t[17337] ^ n[17338];
assign t[17339] = t[17338] ^ n[17339];
assign t[17340] = t[17339] ^ n[17340];
assign t[17341] = t[17340] ^ n[17341];
assign t[17342] = t[17341] ^ n[17342];
assign t[17343] = t[17342] ^ n[17343];
assign t[17344] = t[17343] ^ n[17344];
assign t[17345] = t[17344] ^ n[17345];
assign t[17346] = t[17345] ^ n[17346];
assign t[17347] = t[17346] ^ n[17347];
assign t[17348] = t[17347] ^ n[17348];
assign t[17349] = t[17348] ^ n[17349];
assign t[17350] = t[17349] ^ n[17350];
assign t[17351] = t[17350] ^ n[17351];
assign t[17352] = t[17351] ^ n[17352];
assign t[17353] = t[17352] ^ n[17353];
assign t[17354] = t[17353] ^ n[17354];
assign t[17355] = t[17354] ^ n[17355];
assign t[17356] = t[17355] ^ n[17356];
assign t[17357] = t[17356] ^ n[17357];
assign t[17358] = t[17357] ^ n[17358];
assign t[17359] = t[17358] ^ n[17359];
assign t[17360] = t[17359] ^ n[17360];
assign t[17361] = t[17360] ^ n[17361];
assign t[17362] = t[17361] ^ n[17362];
assign t[17363] = t[17362] ^ n[17363];
assign t[17364] = t[17363] ^ n[17364];
assign t[17365] = t[17364] ^ n[17365];
assign t[17366] = t[17365] ^ n[17366];
assign t[17367] = t[17366] ^ n[17367];
assign t[17368] = t[17367] ^ n[17368];
assign t[17369] = t[17368] ^ n[17369];
assign t[17370] = t[17369] ^ n[17370];
assign t[17371] = t[17370] ^ n[17371];
assign t[17372] = t[17371] ^ n[17372];
assign t[17373] = t[17372] ^ n[17373];
assign t[17374] = t[17373] ^ n[17374];
assign t[17375] = t[17374] ^ n[17375];
assign t[17376] = t[17375] ^ n[17376];
assign t[17377] = t[17376] ^ n[17377];
assign t[17378] = t[17377] ^ n[17378];
assign t[17379] = t[17378] ^ n[17379];
assign t[17380] = t[17379] ^ n[17380];
assign t[17381] = t[17380] ^ n[17381];
assign t[17382] = t[17381] ^ n[17382];
assign t[17383] = t[17382] ^ n[17383];
assign t[17384] = t[17383] ^ n[17384];
assign t[17385] = t[17384] ^ n[17385];
assign t[17386] = t[17385] ^ n[17386];
assign t[17387] = t[17386] ^ n[17387];
assign t[17388] = t[17387] ^ n[17388];
assign t[17389] = t[17388] ^ n[17389];
assign t[17390] = t[17389] ^ n[17390];
assign t[17391] = t[17390] ^ n[17391];
assign t[17392] = t[17391] ^ n[17392];
assign t[17393] = t[17392] ^ n[17393];
assign t[17394] = t[17393] ^ n[17394];
assign t[17395] = t[17394] ^ n[17395];
assign t[17396] = t[17395] ^ n[17396];
assign t[17397] = t[17396] ^ n[17397];
assign t[17398] = t[17397] ^ n[17398];
assign t[17399] = t[17398] ^ n[17399];
assign t[17400] = t[17399] ^ n[17400];
assign t[17401] = t[17400] ^ n[17401];
assign t[17402] = t[17401] ^ n[17402];
assign t[17403] = t[17402] ^ n[17403];
assign t[17404] = t[17403] ^ n[17404];
assign t[17405] = t[17404] ^ n[17405];
assign t[17406] = t[17405] ^ n[17406];
assign t[17407] = t[17406] ^ n[17407];
assign t[17408] = t[17407] ^ n[17408];
assign t[17409] = t[17408] ^ n[17409];
assign t[17410] = t[17409] ^ n[17410];
assign t[17411] = t[17410] ^ n[17411];
assign t[17412] = t[17411] ^ n[17412];
assign t[17413] = t[17412] ^ n[17413];
assign t[17414] = t[17413] ^ n[17414];
assign t[17415] = t[17414] ^ n[17415];
assign t[17416] = t[17415] ^ n[17416];
assign t[17417] = t[17416] ^ n[17417];
assign t[17418] = t[17417] ^ n[17418];
assign t[17419] = t[17418] ^ n[17419];
assign t[17420] = t[17419] ^ n[17420];
assign t[17421] = t[17420] ^ n[17421];
assign t[17422] = t[17421] ^ n[17422];
assign t[17423] = t[17422] ^ n[17423];
assign t[17424] = t[17423] ^ n[17424];
assign t[17425] = t[17424] ^ n[17425];
assign t[17426] = t[17425] ^ n[17426];
assign t[17427] = t[17426] ^ n[17427];
assign t[17428] = t[17427] ^ n[17428];
assign t[17429] = t[17428] ^ n[17429];
assign t[17430] = t[17429] ^ n[17430];
assign t[17431] = t[17430] ^ n[17431];
assign t[17432] = t[17431] ^ n[17432];
assign t[17433] = t[17432] ^ n[17433];
assign t[17434] = t[17433] ^ n[17434];
assign t[17435] = t[17434] ^ n[17435];
assign t[17436] = t[17435] ^ n[17436];
assign t[17437] = t[17436] ^ n[17437];
assign t[17438] = t[17437] ^ n[17438];
assign t[17439] = t[17438] ^ n[17439];
assign t[17440] = t[17439] ^ n[17440];
assign t[17441] = t[17440] ^ n[17441];
assign t[17442] = t[17441] ^ n[17442];
assign t[17443] = t[17442] ^ n[17443];
assign t[17444] = t[17443] ^ n[17444];
assign t[17445] = t[17444] ^ n[17445];
assign t[17446] = t[17445] ^ n[17446];
assign t[17447] = t[17446] ^ n[17447];
assign t[17448] = t[17447] ^ n[17448];
assign t[17449] = t[17448] ^ n[17449];
assign t[17450] = t[17449] ^ n[17450];
assign t[17451] = t[17450] ^ n[17451];
assign t[17452] = t[17451] ^ n[17452];
assign t[17453] = t[17452] ^ n[17453];
assign t[17454] = t[17453] ^ n[17454];
assign t[17455] = t[17454] ^ n[17455];
assign t[17456] = t[17455] ^ n[17456];
assign t[17457] = t[17456] ^ n[17457];
assign t[17458] = t[17457] ^ n[17458];
assign t[17459] = t[17458] ^ n[17459];
assign t[17460] = t[17459] ^ n[17460];
assign t[17461] = t[17460] ^ n[17461];
assign t[17462] = t[17461] ^ n[17462];
assign t[17463] = t[17462] ^ n[17463];
assign t[17464] = t[17463] ^ n[17464];
assign t[17465] = t[17464] ^ n[17465];
assign t[17466] = t[17465] ^ n[17466];
assign t[17467] = t[17466] ^ n[17467];
assign t[17468] = t[17467] ^ n[17468];
assign t[17469] = t[17468] ^ n[17469];
assign t[17470] = t[17469] ^ n[17470];
assign t[17471] = t[17470] ^ n[17471];
assign t[17472] = t[17471] ^ n[17472];
assign t[17473] = t[17472] ^ n[17473];
assign t[17474] = t[17473] ^ n[17474];
assign t[17475] = t[17474] ^ n[17475];
assign t[17476] = t[17475] ^ n[17476];
assign t[17477] = t[17476] ^ n[17477];
assign t[17478] = t[17477] ^ n[17478];
assign t[17479] = t[17478] ^ n[17479];
assign t[17480] = t[17479] ^ n[17480];
assign t[17481] = t[17480] ^ n[17481];
assign t[17482] = t[17481] ^ n[17482];
assign t[17483] = t[17482] ^ n[17483];
assign t[17484] = t[17483] ^ n[17484];
assign t[17485] = t[17484] ^ n[17485];
assign t[17486] = t[17485] ^ n[17486];
assign t[17487] = t[17486] ^ n[17487];
assign t[17488] = t[17487] ^ n[17488];
assign t[17489] = t[17488] ^ n[17489];
assign t[17490] = t[17489] ^ n[17490];
assign t[17491] = t[17490] ^ n[17491];
assign t[17492] = t[17491] ^ n[17492];
assign t[17493] = t[17492] ^ n[17493];
assign t[17494] = t[17493] ^ n[17494];
assign t[17495] = t[17494] ^ n[17495];
assign t[17496] = t[17495] ^ n[17496];
assign t[17497] = t[17496] ^ n[17497];
assign t[17498] = t[17497] ^ n[17498];
assign t[17499] = t[17498] ^ n[17499];
assign t[17500] = t[17499] ^ n[17500];
assign t[17501] = t[17500] ^ n[17501];
assign t[17502] = t[17501] ^ n[17502];
assign t[17503] = t[17502] ^ n[17503];
assign t[17504] = t[17503] ^ n[17504];
assign t[17505] = t[17504] ^ n[17505];
assign t[17506] = t[17505] ^ n[17506];
assign t[17507] = t[17506] ^ n[17507];
assign t[17508] = t[17507] ^ n[17508];
assign t[17509] = t[17508] ^ n[17509];
assign t[17510] = t[17509] ^ n[17510];
assign t[17511] = t[17510] ^ n[17511];
assign t[17512] = t[17511] ^ n[17512];
assign t[17513] = t[17512] ^ n[17513];
assign t[17514] = t[17513] ^ n[17514];
assign t[17515] = t[17514] ^ n[17515];
assign t[17516] = t[17515] ^ n[17516];
assign t[17517] = t[17516] ^ n[17517];
assign t[17518] = t[17517] ^ n[17518];
assign t[17519] = t[17518] ^ n[17519];
assign t[17520] = t[17519] ^ n[17520];
assign t[17521] = t[17520] ^ n[17521];
assign t[17522] = t[17521] ^ n[17522];
assign t[17523] = t[17522] ^ n[17523];
assign t[17524] = t[17523] ^ n[17524];
assign t[17525] = t[17524] ^ n[17525];
assign t[17526] = t[17525] ^ n[17526];
assign t[17527] = t[17526] ^ n[17527];
assign t[17528] = t[17527] ^ n[17528];
assign t[17529] = t[17528] ^ n[17529];
assign t[17530] = t[17529] ^ n[17530];
assign t[17531] = t[17530] ^ n[17531];
assign t[17532] = t[17531] ^ n[17532];
assign t[17533] = t[17532] ^ n[17533];
assign t[17534] = t[17533] ^ n[17534];
assign t[17535] = t[17534] ^ n[17535];
assign t[17536] = t[17535] ^ n[17536];
assign t[17537] = t[17536] ^ n[17537];
assign t[17538] = t[17537] ^ n[17538];
assign t[17539] = t[17538] ^ n[17539];
assign t[17540] = t[17539] ^ n[17540];
assign t[17541] = t[17540] ^ n[17541];
assign t[17542] = t[17541] ^ n[17542];
assign t[17543] = t[17542] ^ n[17543];
assign t[17544] = t[17543] ^ n[17544];
assign t[17545] = t[17544] ^ n[17545];
assign t[17546] = t[17545] ^ n[17546];
assign t[17547] = t[17546] ^ n[17547];
assign t[17548] = t[17547] ^ n[17548];
assign t[17549] = t[17548] ^ n[17549];
assign t[17550] = t[17549] ^ n[17550];
assign t[17551] = t[17550] ^ n[17551];
assign t[17552] = t[17551] ^ n[17552];
assign t[17553] = t[17552] ^ n[17553];
assign t[17554] = t[17553] ^ n[17554];
assign t[17555] = t[17554] ^ n[17555];
assign t[17556] = t[17555] ^ n[17556];
assign t[17557] = t[17556] ^ n[17557];
assign t[17558] = t[17557] ^ n[17558];
assign t[17559] = t[17558] ^ n[17559];
assign t[17560] = t[17559] ^ n[17560];
assign t[17561] = t[17560] ^ n[17561];
assign t[17562] = t[17561] ^ n[17562];
assign t[17563] = t[17562] ^ n[17563];
assign t[17564] = t[17563] ^ n[17564];
assign t[17565] = t[17564] ^ n[17565];
assign t[17566] = t[17565] ^ n[17566];
assign t[17567] = t[17566] ^ n[17567];
assign t[17568] = t[17567] ^ n[17568];
assign t[17569] = t[17568] ^ n[17569];
assign t[17570] = t[17569] ^ n[17570];
assign t[17571] = t[17570] ^ n[17571];
assign t[17572] = t[17571] ^ n[17572];
assign t[17573] = t[17572] ^ n[17573];
assign t[17574] = t[17573] ^ n[17574];
assign t[17575] = t[17574] ^ n[17575];
assign t[17576] = t[17575] ^ n[17576];
assign t[17577] = t[17576] ^ n[17577];
assign t[17578] = t[17577] ^ n[17578];
assign t[17579] = t[17578] ^ n[17579];
assign t[17580] = t[17579] ^ n[17580];
assign t[17581] = t[17580] ^ n[17581];
assign t[17582] = t[17581] ^ n[17582];
assign t[17583] = t[17582] ^ n[17583];
assign t[17584] = t[17583] ^ n[17584];
assign t[17585] = t[17584] ^ n[17585];
assign t[17586] = t[17585] ^ n[17586];
assign t[17587] = t[17586] ^ n[17587];
assign t[17588] = t[17587] ^ n[17588];
assign t[17589] = t[17588] ^ n[17589];
assign t[17590] = t[17589] ^ n[17590];
assign t[17591] = t[17590] ^ n[17591];
assign t[17592] = t[17591] ^ n[17592];
assign t[17593] = t[17592] ^ n[17593];
assign t[17594] = t[17593] ^ n[17594];
assign t[17595] = t[17594] ^ n[17595];
assign t[17596] = t[17595] ^ n[17596];
assign t[17597] = t[17596] ^ n[17597];
assign t[17598] = t[17597] ^ n[17598];
assign t[17599] = t[17598] ^ n[17599];
assign t[17600] = t[17599] ^ n[17600];
assign t[17601] = t[17600] ^ n[17601];
assign t[17602] = t[17601] ^ n[17602];
assign t[17603] = t[17602] ^ n[17603];
assign t[17604] = t[17603] ^ n[17604];
assign t[17605] = t[17604] ^ n[17605];
assign t[17606] = t[17605] ^ n[17606];
assign t[17607] = t[17606] ^ n[17607];
assign t[17608] = t[17607] ^ n[17608];
assign t[17609] = t[17608] ^ n[17609];
assign t[17610] = t[17609] ^ n[17610];
assign t[17611] = t[17610] ^ n[17611];
assign t[17612] = t[17611] ^ n[17612];
assign t[17613] = t[17612] ^ n[17613];
assign t[17614] = t[17613] ^ n[17614];
assign t[17615] = t[17614] ^ n[17615];
assign t[17616] = t[17615] ^ n[17616];
assign t[17617] = t[17616] ^ n[17617];
assign t[17618] = t[17617] ^ n[17618];
assign t[17619] = t[17618] ^ n[17619];
assign t[17620] = t[17619] ^ n[17620];
assign t[17621] = t[17620] ^ n[17621];
assign t[17622] = t[17621] ^ n[17622];
assign t[17623] = t[17622] ^ n[17623];
assign t[17624] = t[17623] ^ n[17624];
assign t[17625] = t[17624] ^ n[17625];
assign t[17626] = t[17625] ^ n[17626];
assign t[17627] = t[17626] ^ n[17627];
assign t[17628] = t[17627] ^ n[17628];
assign t[17629] = t[17628] ^ n[17629];
assign t[17630] = t[17629] ^ n[17630];
assign t[17631] = t[17630] ^ n[17631];
assign t[17632] = t[17631] ^ n[17632];
assign t[17633] = t[17632] ^ n[17633];
assign t[17634] = t[17633] ^ n[17634];
assign t[17635] = t[17634] ^ n[17635];
assign t[17636] = t[17635] ^ n[17636];
assign t[17637] = t[17636] ^ n[17637];
assign t[17638] = t[17637] ^ n[17638];
assign t[17639] = t[17638] ^ n[17639];
assign t[17640] = t[17639] ^ n[17640];
assign t[17641] = t[17640] ^ n[17641];
assign t[17642] = t[17641] ^ n[17642];
assign t[17643] = t[17642] ^ n[17643];
assign t[17644] = t[17643] ^ n[17644];
assign t[17645] = t[17644] ^ n[17645];
assign t[17646] = t[17645] ^ n[17646];
assign t[17647] = t[17646] ^ n[17647];
assign t[17648] = t[17647] ^ n[17648];
assign t[17649] = t[17648] ^ n[17649];
assign t[17650] = t[17649] ^ n[17650];
assign t[17651] = t[17650] ^ n[17651];
assign t[17652] = t[17651] ^ n[17652];
assign t[17653] = t[17652] ^ n[17653];
assign t[17654] = t[17653] ^ n[17654];
assign t[17655] = t[17654] ^ n[17655];
assign t[17656] = t[17655] ^ n[17656];
assign t[17657] = t[17656] ^ n[17657];
assign t[17658] = t[17657] ^ n[17658];
assign t[17659] = t[17658] ^ n[17659];
assign t[17660] = t[17659] ^ n[17660];
assign t[17661] = t[17660] ^ n[17661];
assign t[17662] = t[17661] ^ n[17662];
assign t[17663] = t[17662] ^ n[17663];
assign t[17664] = t[17663] ^ n[17664];
assign t[17665] = t[17664] ^ n[17665];
assign t[17666] = t[17665] ^ n[17666];
assign t[17667] = t[17666] ^ n[17667];
assign t[17668] = t[17667] ^ n[17668];
assign t[17669] = t[17668] ^ n[17669];
assign t[17670] = t[17669] ^ n[17670];
assign t[17671] = t[17670] ^ n[17671];
assign t[17672] = t[17671] ^ n[17672];
assign t[17673] = t[17672] ^ n[17673];
assign t[17674] = t[17673] ^ n[17674];
assign t[17675] = t[17674] ^ n[17675];
assign t[17676] = t[17675] ^ n[17676];
assign t[17677] = t[17676] ^ n[17677];
assign t[17678] = t[17677] ^ n[17678];
assign t[17679] = t[17678] ^ n[17679];
assign t[17680] = t[17679] ^ n[17680];
assign t[17681] = t[17680] ^ n[17681];
assign t[17682] = t[17681] ^ n[17682];
assign t[17683] = t[17682] ^ n[17683];
assign t[17684] = t[17683] ^ n[17684];
assign t[17685] = t[17684] ^ n[17685];
assign t[17686] = t[17685] ^ n[17686];
assign t[17687] = t[17686] ^ n[17687];
assign t[17688] = t[17687] ^ n[17688];
assign t[17689] = t[17688] ^ n[17689];
assign t[17690] = t[17689] ^ n[17690];
assign t[17691] = t[17690] ^ n[17691];
assign t[17692] = t[17691] ^ n[17692];
assign t[17693] = t[17692] ^ n[17693];
assign t[17694] = t[17693] ^ n[17694];
assign t[17695] = t[17694] ^ n[17695];
assign t[17696] = t[17695] ^ n[17696];
assign t[17697] = t[17696] ^ n[17697];
assign t[17698] = t[17697] ^ n[17698];
assign t[17699] = t[17698] ^ n[17699];
assign t[17700] = t[17699] ^ n[17700];
assign t[17701] = t[17700] ^ n[17701];
assign t[17702] = t[17701] ^ n[17702];
assign t[17703] = t[17702] ^ n[17703];
assign t[17704] = t[17703] ^ n[17704];
assign t[17705] = t[17704] ^ n[17705];
assign t[17706] = t[17705] ^ n[17706];
assign t[17707] = t[17706] ^ n[17707];
assign t[17708] = t[17707] ^ n[17708];
assign t[17709] = t[17708] ^ n[17709];
assign t[17710] = t[17709] ^ n[17710];
assign t[17711] = t[17710] ^ n[17711];
assign t[17712] = t[17711] ^ n[17712];
assign t[17713] = t[17712] ^ n[17713];
assign t[17714] = t[17713] ^ n[17714];
assign t[17715] = t[17714] ^ n[17715];
assign t[17716] = t[17715] ^ n[17716];
assign t[17717] = t[17716] ^ n[17717];
assign t[17718] = t[17717] ^ n[17718];
assign t[17719] = t[17718] ^ n[17719];
assign t[17720] = t[17719] ^ n[17720];
assign t[17721] = t[17720] ^ n[17721];
assign t[17722] = t[17721] ^ n[17722];
assign t[17723] = t[17722] ^ n[17723];
assign t[17724] = t[17723] ^ n[17724];
assign t[17725] = t[17724] ^ n[17725];
assign t[17726] = t[17725] ^ n[17726];
assign t[17727] = t[17726] ^ n[17727];
assign t[17728] = t[17727] ^ n[17728];
assign t[17729] = t[17728] ^ n[17729];
assign t[17730] = t[17729] ^ n[17730];
assign t[17731] = t[17730] ^ n[17731];
assign t[17732] = t[17731] ^ n[17732];
assign t[17733] = t[17732] ^ n[17733];
assign t[17734] = t[17733] ^ n[17734];
assign t[17735] = t[17734] ^ n[17735];
assign t[17736] = t[17735] ^ n[17736];
assign t[17737] = t[17736] ^ n[17737];
assign t[17738] = t[17737] ^ n[17738];
assign t[17739] = t[17738] ^ n[17739];
assign t[17740] = t[17739] ^ n[17740];
assign t[17741] = t[17740] ^ n[17741];
assign t[17742] = t[17741] ^ n[17742];
assign t[17743] = t[17742] ^ n[17743];
assign t[17744] = t[17743] ^ n[17744];
assign t[17745] = t[17744] ^ n[17745];
assign t[17746] = t[17745] ^ n[17746];
assign t[17747] = t[17746] ^ n[17747];
assign t[17748] = t[17747] ^ n[17748];
assign t[17749] = t[17748] ^ n[17749];
assign t[17750] = t[17749] ^ n[17750];
assign t[17751] = t[17750] ^ n[17751];
assign t[17752] = t[17751] ^ n[17752];
assign t[17753] = t[17752] ^ n[17753];
assign t[17754] = t[17753] ^ n[17754];
assign t[17755] = t[17754] ^ n[17755];
assign t[17756] = t[17755] ^ n[17756];
assign t[17757] = t[17756] ^ n[17757];
assign t[17758] = t[17757] ^ n[17758];
assign t[17759] = t[17758] ^ n[17759];
assign t[17760] = t[17759] ^ n[17760];
assign t[17761] = t[17760] ^ n[17761];
assign t[17762] = t[17761] ^ n[17762];
assign t[17763] = t[17762] ^ n[17763];
assign t[17764] = t[17763] ^ n[17764];
assign t[17765] = t[17764] ^ n[17765];
assign t[17766] = t[17765] ^ n[17766];
assign t[17767] = t[17766] ^ n[17767];
assign t[17768] = t[17767] ^ n[17768];
assign t[17769] = t[17768] ^ n[17769];
assign t[17770] = t[17769] ^ n[17770];
assign t[17771] = t[17770] ^ n[17771];
assign t[17772] = t[17771] ^ n[17772];
assign t[17773] = t[17772] ^ n[17773];
assign t[17774] = t[17773] ^ n[17774];
assign t[17775] = t[17774] ^ n[17775];
assign t[17776] = t[17775] ^ n[17776];
assign t[17777] = t[17776] ^ n[17777];
assign t[17778] = t[17777] ^ n[17778];
assign t[17779] = t[17778] ^ n[17779];
assign t[17780] = t[17779] ^ n[17780];
assign t[17781] = t[17780] ^ n[17781];
assign t[17782] = t[17781] ^ n[17782];
assign t[17783] = t[17782] ^ n[17783];
assign t[17784] = t[17783] ^ n[17784];
assign t[17785] = t[17784] ^ n[17785];
assign t[17786] = t[17785] ^ n[17786];
assign t[17787] = t[17786] ^ n[17787];
assign t[17788] = t[17787] ^ n[17788];
assign t[17789] = t[17788] ^ n[17789];
assign t[17790] = t[17789] ^ n[17790];
assign t[17791] = t[17790] ^ n[17791];
assign t[17792] = t[17791] ^ n[17792];
assign t[17793] = t[17792] ^ n[17793];
assign t[17794] = t[17793] ^ n[17794];
assign t[17795] = t[17794] ^ n[17795];
assign t[17796] = t[17795] ^ n[17796];
assign t[17797] = t[17796] ^ n[17797];
assign t[17798] = t[17797] ^ n[17798];
assign t[17799] = t[17798] ^ n[17799];
assign t[17800] = t[17799] ^ n[17800];
assign t[17801] = t[17800] ^ n[17801];
assign t[17802] = t[17801] ^ n[17802];
assign t[17803] = t[17802] ^ n[17803];
assign t[17804] = t[17803] ^ n[17804];
assign t[17805] = t[17804] ^ n[17805];
assign t[17806] = t[17805] ^ n[17806];
assign t[17807] = t[17806] ^ n[17807];
assign t[17808] = t[17807] ^ n[17808];
assign t[17809] = t[17808] ^ n[17809];
assign t[17810] = t[17809] ^ n[17810];
assign t[17811] = t[17810] ^ n[17811];
assign t[17812] = t[17811] ^ n[17812];
assign t[17813] = t[17812] ^ n[17813];
assign t[17814] = t[17813] ^ n[17814];
assign t[17815] = t[17814] ^ n[17815];
assign t[17816] = t[17815] ^ n[17816];
assign t[17817] = t[17816] ^ n[17817];
assign t[17818] = t[17817] ^ n[17818];
assign t[17819] = t[17818] ^ n[17819];
assign t[17820] = t[17819] ^ n[17820];
assign t[17821] = t[17820] ^ n[17821];
assign t[17822] = t[17821] ^ n[17822];
assign t[17823] = t[17822] ^ n[17823];
assign t[17824] = t[17823] ^ n[17824];
assign t[17825] = t[17824] ^ n[17825];
assign t[17826] = t[17825] ^ n[17826];
assign t[17827] = t[17826] ^ n[17827];
assign t[17828] = t[17827] ^ n[17828];
assign t[17829] = t[17828] ^ n[17829];
assign t[17830] = t[17829] ^ n[17830];
assign t[17831] = t[17830] ^ n[17831];
assign t[17832] = t[17831] ^ n[17832];
assign t[17833] = t[17832] ^ n[17833];
assign t[17834] = t[17833] ^ n[17834];
assign t[17835] = t[17834] ^ n[17835];
assign t[17836] = t[17835] ^ n[17836];
assign t[17837] = t[17836] ^ n[17837];
assign t[17838] = t[17837] ^ n[17838];
assign t[17839] = t[17838] ^ n[17839];
assign t[17840] = t[17839] ^ n[17840];
assign t[17841] = t[17840] ^ n[17841];
assign t[17842] = t[17841] ^ n[17842];
assign t[17843] = t[17842] ^ n[17843];
assign t[17844] = t[17843] ^ n[17844];
assign t[17845] = t[17844] ^ n[17845];
assign t[17846] = t[17845] ^ n[17846];
assign t[17847] = t[17846] ^ n[17847];
assign t[17848] = t[17847] ^ n[17848];
assign t[17849] = t[17848] ^ n[17849];
assign t[17850] = t[17849] ^ n[17850];
assign t[17851] = t[17850] ^ n[17851];
assign t[17852] = t[17851] ^ n[17852];
assign t[17853] = t[17852] ^ n[17853];
assign t[17854] = t[17853] ^ n[17854];
assign t[17855] = t[17854] ^ n[17855];
assign t[17856] = t[17855] ^ n[17856];
assign t[17857] = t[17856] ^ n[17857];
assign t[17858] = t[17857] ^ n[17858];
assign t[17859] = t[17858] ^ n[17859];
assign t[17860] = t[17859] ^ n[17860];
assign t[17861] = t[17860] ^ n[17861];
assign t[17862] = t[17861] ^ n[17862];
assign t[17863] = t[17862] ^ n[17863];
assign t[17864] = t[17863] ^ n[17864];
assign t[17865] = t[17864] ^ n[17865];
assign t[17866] = t[17865] ^ n[17866];
assign t[17867] = t[17866] ^ n[17867];
assign t[17868] = t[17867] ^ n[17868];
assign t[17869] = t[17868] ^ n[17869];
assign t[17870] = t[17869] ^ n[17870];
assign t[17871] = t[17870] ^ n[17871];
assign t[17872] = t[17871] ^ n[17872];
assign t[17873] = t[17872] ^ n[17873];
assign t[17874] = t[17873] ^ n[17874];
assign t[17875] = t[17874] ^ n[17875];
assign t[17876] = t[17875] ^ n[17876];
assign t[17877] = t[17876] ^ n[17877];
assign t[17878] = t[17877] ^ n[17878];
assign t[17879] = t[17878] ^ n[17879];
assign t[17880] = t[17879] ^ n[17880];
assign t[17881] = t[17880] ^ n[17881];
assign t[17882] = t[17881] ^ n[17882];
assign t[17883] = t[17882] ^ n[17883];
assign t[17884] = t[17883] ^ n[17884];
assign t[17885] = t[17884] ^ n[17885];
assign t[17886] = t[17885] ^ n[17886];
assign t[17887] = t[17886] ^ n[17887];
assign t[17888] = t[17887] ^ n[17888];
assign t[17889] = t[17888] ^ n[17889];
assign t[17890] = t[17889] ^ n[17890];
assign t[17891] = t[17890] ^ n[17891];
assign t[17892] = t[17891] ^ n[17892];
assign t[17893] = t[17892] ^ n[17893];
assign t[17894] = t[17893] ^ n[17894];
assign t[17895] = t[17894] ^ n[17895];
assign t[17896] = t[17895] ^ n[17896];
assign t[17897] = t[17896] ^ n[17897];
assign t[17898] = t[17897] ^ n[17898];
assign t[17899] = t[17898] ^ n[17899];
assign t[17900] = t[17899] ^ n[17900];
assign t[17901] = t[17900] ^ n[17901];
assign t[17902] = t[17901] ^ n[17902];
assign t[17903] = t[17902] ^ n[17903];
assign t[17904] = t[17903] ^ n[17904];
assign t[17905] = t[17904] ^ n[17905];
assign t[17906] = t[17905] ^ n[17906];
assign t[17907] = t[17906] ^ n[17907];
assign t[17908] = t[17907] ^ n[17908];
assign t[17909] = t[17908] ^ n[17909];
assign t[17910] = t[17909] ^ n[17910];
assign t[17911] = t[17910] ^ n[17911];
assign t[17912] = t[17911] ^ n[17912];
assign t[17913] = t[17912] ^ n[17913];
assign t[17914] = t[17913] ^ n[17914];
assign t[17915] = t[17914] ^ n[17915];
assign t[17916] = t[17915] ^ n[17916];
assign t[17917] = t[17916] ^ n[17917];
assign t[17918] = t[17917] ^ n[17918];
assign t[17919] = t[17918] ^ n[17919];
assign t[17920] = t[17919] ^ n[17920];
assign t[17921] = t[17920] ^ n[17921];
assign t[17922] = t[17921] ^ n[17922];
assign t[17923] = t[17922] ^ n[17923];
assign t[17924] = t[17923] ^ n[17924];
assign t[17925] = t[17924] ^ n[17925];
assign t[17926] = t[17925] ^ n[17926];
assign t[17927] = t[17926] ^ n[17927];
assign t[17928] = t[17927] ^ n[17928];
assign t[17929] = t[17928] ^ n[17929];
assign t[17930] = t[17929] ^ n[17930];
assign t[17931] = t[17930] ^ n[17931];
assign t[17932] = t[17931] ^ n[17932];
assign t[17933] = t[17932] ^ n[17933];
assign t[17934] = t[17933] ^ n[17934];
assign t[17935] = t[17934] ^ n[17935];
assign t[17936] = t[17935] ^ n[17936];
assign t[17937] = t[17936] ^ n[17937];
assign t[17938] = t[17937] ^ n[17938];
assign t[17939] = t[17938] ^ n[17939];
assign t[17940] = t[17939] ^ n[17940];
assign t[17941] = t[17940] ^ n[17941];
assign t[17942] = t[17941] ^ n[17942];
assign t[17943] = t[17942] ^ n[17943];
assign t[17944] = t[17943] ^ n[17944];
assign t[17945] = t[17944] ^ n[17945];
assign t[17946] = t[17945] ^ n[17946];
assign t[17947] = t[17946] ^ n[17947];
assign t[17948] = t[17947] ^ n[17948];
assign t[17949] = t[17948] ^ n[17949];
assign t[17950] = t[17949] ^ n[17950];
assign t[17951] = t[17950] ^ n[17951];
assign t[17952] = t[17951] ^ n[17952];
assign t[17953] = t[17952] ^ n[17953];
assign t[17954] = t[17953] ^ n[17954];
assign t[17955] = t[17954] ^ n[17955];
assign t[17956] = t[17955] ^ n[17956];
assign t[17957] = t[17956] ^ n[17957];
assign t[17958] = t[17957] ^ n[17958];
assign t[17959] = t[17958] ^ n[17959];
assign t[17960] = t[17959] ^ n[17960];
assign t[17961] = t[17960] ^ n[17961];
assign t[17962] = t[17961] ^ n[17962];
assign t[17963] = t[17962] ^ n[17963];
assign t[17964] = t[17963] ^ n[17964];
assign t[17965] = t[17964] ^ n[17965];
assign t[17966] = t[17965] ^ n[17966];
assign t[17967] = t[17966] ^ n[17967];
assign t[17968] = t[17967] ^ n[17968];
assign t[17969] = t[17968] ^ n[17969];
assign t[17970] = t[17969] ^ n[17970];
assign t[17971] = t[17970] ^ n[17971];
assign t[17972] = t[17971] ^ n[17972];
assign t[17973] = t[17972] ^ n[17973];
assign t[17974] = t[17973] ^ n[17974];
assign t[17975] = t[17974] ^ n[17975];
assign t[17976] = t[17975] ^ n[17976];
assign t[17977] = t[17976] ^ n[17977];
assign t[17978] = t[17977] ^ n[17978];
assign t[17979] = t[17978] ^ n[17979];
assign t[17980] = t[17979] ^ n[17980];
assign t[17981] = t[17980] ^ n[17981];
assign t[17982] = t[17981] ^ n[17982];
assign t[17983] = t[17982] ^ n[17983];
assign t[17984] = t[17983] ^ n[17984];
assign t[17985] = t[17984] ^ n[17985];
assign t[17986] = t[17985] ^ n[17986];
assign t[17987] = t[17986] ^ n[17987];
assign t[17988] = t[17987] ^ n[17988];
assign t[17989] = t[17988] ^ n[17989];
assign t[17990] = t[17989] ^ n[17990];
assign t[17991] = t[17990] ^ n[17991];
assign t[17992] = t[17991] ^ n[17992];
assign t[17993] = t[17992] ^ n[17993];
assign t[17994] = t[17993] ^ n[17994];
assign t[17995] = t[17994] ^ n[17995];
assign t[17996] = t[17995] ^ n[17996];
assign t[17997] = t[17996] ^ n[17997];
assign t[17998] = t[17997] ^ n[17998];
assign t[17999] = t[17998] ^ n[17999];
assign t[18000] = t[17999] ^ n[18000];
assign t[18001] = t[18000] ^ n[18001];
assign t[18002] = t[18001] ^ n[18002];
assign t[18003] = t[18002] ^ n[18003];
assign t[18004] = t[18003] ^ n[18004];
assign t[18005] = t[18004] ^ n[18005];
assign t[18006] = t[18005] ^ n[18006];
assign t[18007] = t[18006] ^ n[18007];
assign t[18008] = t[18007] ^ n[18008];
assign t[18009] = t[18008] ^ n[18009];
assign t[18010] = t[18009] ^ n[18010];
assign t[18011] = t[18010] ^ n[18011];
assign t[18012] = t[18011] ^ n[18012];
assign t[18013] = t[18012] ^ n[18013];
assign t[18014] = t[18013] ^ n[18014];
assign t[18015] = t[18014] ^ n[18015];
assign t[18016] = t[18015] ^ n[18016];
assign t[18017] = t[18016] ^ n[18017];
assign t[18018] = t[18017] ^ n[18018];
assign t[18019] = t[18018] ^ n[18019];
assign t[18020] = t[18019] ^ n[18020];
assign t[18021] = t[18020] ^ n[18021];
assign t[18022] = t[18021] ^ n[18022];
assign t[18023] = t[18022] ^ n[18023];
assign t[18024] = t[18023] ^ n[18024];
assign t[18025] = t[18024] ^ n[18025];
assign t[18026] = t[18025] ^ n[18026];
assign t[18027] = t[18026] ^ n[18027];
assign t[18028] = t[18027] ^ n[18028];
assign t[18029] = t[18028] ^ n[18029];
assign t[18030] = t[18029] ^ n[18030];
assign t[18031] = t[18030] ^ n[18031];
assign t[18032] = t[18031] ^ n[18032];
assign t[18033] = t[18032] ^ n[18033];
assign t[18034] = t[18033] ^ n[18034];
assign t[18035] = t[18034] ^ n[18035];
assign t[18036] = t[18035] ^ n[18036];
assign t[18037] = t[18036] ^ n[18037];
assign t[18038] = t[18037] ^ n[18038];
assign t[18039] = t[18038] ^ n[18039];
assign t[18040] = t[18039] ^ n[18040];
assign t[18041] = t[18040] ^ n[18041];
assign t[18042] = t[18041] ^ n[18042];
assign t[18043] = t[18042] ^ n[18043];
assign t[18044] = t[18043] ^ n[18044];
assign t[18045] = t[18044] ^ n[18045];
assign t[18046] = t[18045] ^ n[18046];
assign t[18047] = t[18046] ^ n[18047];
assign t[18048] = t[18047] ^ n[18048];
assign t[18049] = t[18048] ^ n[18049];
assign t[18050] = t[18049] ^ n[18050];
assign t[18051] = t[18050] ^ n[18051];
assign t[18052] = t[18051] ^ n[18052];
assign t[18053] = t[18052] ^ n[18053];
assign t[18054] = t[18053] ^ n[18054];
assign t[18055] = t[18054] ^ n[18055];
assign t[18056] = t[18055] ^ n[18056];
assign t[18057] = t[18056] ^ n[18057];
assign t[18058] = t[18057] ^ n[18058];
assign t[18059] = t[18058] ^ n[18059];
assign t[18060] = t[18059] ^ n[18060];
assign t[18061] = t[18060] ^ n[18061];
assign t[18062] = t[18061] ^ n[18062];
assign t[18063] = t[18062] ^ n[18063];
assign t[18064] = t[18063] ^ n[18064];
assign t[18065] = t[18064] ^ n[18065];
assign t[18066] = t[18065] ^ n[18066];
assign t[18067] = t[18066] ^ n[18067];
assign t[18068] = t[18067] ^ n[18068];
assign t[18069] = t[18068] ^ n[18069];
assign t[18070] = t[18069] ^ n[18070];
assign t[18071] = t[18070] ^ n[18071];
assign t[18072] = t[18071] ^ n[18072];
assign t[18073] = t[18072] ^ n[18073];
assign t[18074] = t[18073] ^ n[18074];
assign t[18075] = t[18074] ^ n[18075];
assign t[18076] = t[18075] ^ n[18076];
assign t[18077] = t[18076] ^ n[18077];
assign t[18078] = t[18077] ^ n[18078];
assign t[18079] = t[18078] ^ n[18079];
assign t[18080] = t[18079] ^ n[18080];
assign t[18081] = t[18080] ^ n[18081];
assign t[18082] = t[18081] ^ n[18082];
assign t[18083] = t[18082] ^ n[18083];
assign t[18084] = t[18083] ^ n[18084];
assign t[18085] = t[18084] ^ n[18085];
assign t[18086] = t[18085] ^ n[18086];
assign t[18087] = t[18086] ^ n[18087];
assign t[18088] = t[18087] ^ n[18088];
assign t[18089] = t[18088] ^ n[18089];
assign t[18090] = t[18089] ^ n[18090];
assign t[18091] = t[18090] ^ n[18091];
assign t[18092] = t[18091] ^ n[18092];
assign t[18093] = t[18092] ^ n[18093];
assign t[18094] = t[18093] ^ n[18094];
assign t[18095] = t[18094] ^ n[18095];
assign t[18096] = t[18095] ^ n[18096];
assign t[18097] = t[18096] ^ n[18097];
assign t[18098] = t[18097] ^ n[18098];
assign t[18099] = t[18098] ^ n[18099];
assign t[18100] = t[18099] ^ n[18100];
assign t[18101] = t[18100] ^ n[18101];
assign t[18102] = t[18101] ^ n[18102];
assign t[18103] = t[18102] ^ n[18103];
assign t[18104] = t[18103] ^ n[18104];
assign t[18105] = t[18104] ^ n[18105];
assign t[18106] = t[18105] ^ n[18106];
assign t[18107] = t[18106] ^ n[18107];
assign t[18108] = t[18107] ^ n[18108];
assign t[18109] = t[18108] ^ n[18109];
assign t[18110] = t[18109] ^ n[18110];
assign t[18111] = t[18110] ^ n[18111];
assign t[18112] = t[18111] ^ n[18112];
assign t[18113] = t[18112] ^ n[18113];
assign t[18114] = t[18113] ^ n[18114];
assign t[18115] = t[18114] ^ n[18115];
assign t[18116] = t[18115] ^ n[18116];
assign t[18117] = t[18116] ^ n[18117];
assign t[18118] = t[18117] ^ n[18118];
assign t[18119] = t[18118] ^ n[18119];
assign t[18120] = t[18119] ^ n[18120];
assign t[18121] = t[18120] ^ n[18121];
assign t[18122] = t[18121] ^ n[18122];
assign t[18123] = t[18122] ^ n[18123];
assign t[18124] = t[18123] ^ n[18124];
assign t[18125] = t[18124] ^ n[18125];
assign t[18126] = t[18125] ^ n[18126];
assign t[18127] = t[18126] ^ n[18127];
assign t[18128] = t[18127] ^ n[18128];
assign t[18129] = t[18128] ^ n[18129];
assign t[18130] = t[18129] ^ n[18130];
assign t[18131] = t[18130] ^ n[18131];
assign t[18132] = t[18131] ^ n[18132];
assign t[18133] = t[18132] ^ n[18133];
assign t[18134] = t[18133] ^ n[18134];
assign t[18135] = t[18134] ^ n[18135];
assign t[18136] = t[18135] ^ n[18136];
assign t[18137] = t[18136] ^ n[18137];
assign t[18138] = t[18137] ^ n[18138];
assign t[18139] = t[18138] ^ n[18139];
assign t[18140] = t[18139] ^ n[18140];
assign t[18141] = t[18140] ^ n[18141];
assign t[18142] = t[18141] ^ n[18142];
assign t[18143] = t[18142] ^ n[18143];
assign t[18144] = t[18143] ^ n[18144];
assign t[18145] = t[18144] ^ n[18145];
assign t[18146] = t[18145] ^ n[18146];
assign t[18147] = t[18146] ^ n[18147];
assign t[18148] = t[18147] ^ n[18148];
assign t[18149] = t[18148] ^ n[18149];
assign t[18150] = t[18149] ^ n[18150];
assign t[18151] = t[18150] ^ n[18151];
assign t[18152] = t[18151] ^ n[18152];
assign t[18153] = t[18152] ^ n[18153];
assign t[18154] = t[18153] ^ n[18154];
assign t[18155] = t[18154] ^ n[18155];
assign t[18156] = t[18155] ^ n[18156];
assign t[18157] = t[18156] ^ n[18157];
assign t[18158] = t[18157] ^ n[18158];
assign t[18159] = t[18158] ^ n[18159];
assign t[18160] = t[18159] ^ n[18160];
assign t[18161] = t[18160] ^ n[18161];
assign t[18162] = t[18161] ^ n[18162];
assign t[18163] = t[18162] ^ n[18163];
assign t[18164] = t[18163] ^ n[18164];
assign t[18165] = t[18164] ^ n[18165];
assign t[18166] = t[18165] ^ n[18166];
assign t[18167] = t[18166] ^ n[18167];
assign t[18168] = t[18167] ^ n[18168];
assign t[18169] = t[18168] ^ n[18169];
assign t[18170] = t[18169] ^ n[18170];
assign t[18171] = t[18170] ^ n[18171];
assign t[18172] = t[18171] ^ n[18172];
assign t[18173] = t[18172] ^ n[18173];
assign t[18174] = t[18173] ^ n[18174];
assign t[18175] = t[18174] ^ n[18175];
assign t[18176] = t[18175] ^ n[18176];
assign t[18177] = t[18176] ^ n[18177];
assign t[18178] = t[18177] ^ n[18178];
assign t[18179] = t[18178] ^ n[18179];
assign t[18180] = t[18179] ^ n[18180];
assign t[18181] = t[18180] ^ n[18181];
assign t[18182] = t[18181] ^ n[18182];
assign t[18183] = t[18182] ^ n[18183];
assign t[18184] = t[18183] ^ n[18184];
assign t[18185] = t[18184] ^ n[18185];
assign t[18186] = t[18185] ^ n[18186];
assign t[18187] = t[18186] ^ n[18187];
assign t[18188] = t[18187] ^ n[18188];
assign t[18189] = t[18188] ^ n[18189];
assign t[18190] = t[18189] ^ n[18190];
assign t[18191] = t[18190] ^ n[18191];
assign t[18192] = t[18191] ^ n[18192];
assign t[18193] = t[18192] ^ n[18193];
assign t[18194] = t[18193] ^ n[18194];
assign t[18195] = t[18194] ^ n[18195];
assign t[18196] = t[18195] ^ n[18196];
assign t[18197] = t[18196] ^ n[18197];
assign t[18198] = t[18197] ^ n[18198];
assign t[18199] = t[18198] ^ n[18199];
assign t[18200] = t[18199] ^ n[18200];
assign t[18201] = t[18200] ^ n[18201];
assign t[18202] = t[18201] ^ n[18202];
assign t[18203] = t[18202] ^ n[18203];
assign t[18204] = t[18203] ^ n[18204];
assign t[18205] = t[18204] ^ n[18205];
assign t[18206] = t[18205] ^ n[18206];
assign t[18207] = t[18206] ^ n[18207];
assign t[18208] = t[18207] ^ n[18208];
assign t[18209] = t[18208] ^ n[18209];
assign t[18210] = t[18209] ^ n[18210];
assign t[18211] = t[18210] ^ n[18211];
assign t[18212] = t[18211] ^ n[18212];
assign t[18213] = t[18212] ^ n[18213];
assign t[18214] = t[18213] ^ n[18214];
assign t[18215] = t[18214] ^ n[18215];
assign t[18216] = t[18215] ^ n[18216];
assign t[18217] = t[18216] ^ n[18217];
assign t[18218] = t[18217] ^ n[18218];
assign t[18219] = t[18218] ^ n[18219];
assign t[18220] = t[18219] ^ n[18220];
assign t[18221] = t[18220] ^ n[18221];
assign t[18222] = t[18221] ^ n[18222];
assign t[18223] = t[18222] ^ n[18223];
assign t[18224] = t[18223] ^ n[18224];
assign t[18225] = t[18224] ^ n[18225];
assign t[18226] = t[18225] ^ n[18226];
assign t[18227] = t[18226] ^ n[18227];
assign t[18228] = t[18227] ^ n[18228];
assign t[18229] = t[18228] ^ n[18229];
assign t[18230] = t[18229] ^ n[18230];
assign t[18231] = t[18230] ^ n[18231];
assign t[18232] = t[18231] ^ n[18232];
assign t[18233] = t[18232] ^ n[18233];
assign t[18234] = t[18233] ^ n[18234];
assign t[18235] = t[18234] ^ n[18235];
assign t[18236] = t[18235] ^ n[18236];
assign t[18237] = t[18236] ^ n[18237];
assign t[18238] = t[18237] ^ n[18238];
assign t[18239] = t[18238] ^ n[18239];
assign t[18240] = t[18239] ^ n[18240];
assign t[18241] = t[18240] ^ n[18241];
assign t[18242] = t[18241] ^ n[18242];
assign t[18243] = t[18242] ^ n[18243];
assign t[18244] = t[18243] ^ n[18244];
assign t[18245] = t[18244] ^ n[18245];
assign t[18246] = t[18245] ^ n[18246];
assign t[18247] = t[18246] ^ n[18247];
assign t[18248] = t[18247] ^ n[18248];
assign t[18249] = t[18248] ^ n[18249];
assign t[18250] = t[18249] ^ n[18250];
assign t[18251] = t[18250] ^ n[18251];
assign t[18252] = t[18251] ^ n[18252];
assign t[18253] = t[18252] ^ n[18253];
assign t[18254] = t[18253] ^ n[18254];
assign t[18255] = t[18254] ^ n[18255];
assign t[18256] = t[18255] ^ n[18256];
assign t[18257] = t[18256] ^ n[18257];
assign t[18258] = t[18257] ^ n[18258];
assign t[18259] = t[18258] ^ n[18259];
assign t[18260] = t[18259] ^ n[18260];
assign t[18261] = t[18260] ^ n[18261];
assign t[18262] = t[18261] ^ n[18262];
assign t[18263] = t[18262] ^ n[18263];
assign t[18264] = t[18263] ^ n[18264];
assign t[18265] = t[18264] ^ n[18265];
assign t[18266] = t[18265] ^ n[18266];
assign t[18267] = t[18266] ^ n[18267];
assign t[18268] = t[18267] ^ n[18268];
assign t[18269] = t[18268] ^ n[18269];
assign t[18270] = t[18269] ^ n[18270];
assign t[18271] = t[18270] ^ n[18271];
assign t[18272] = t[18271] ^ n[18272];
assign t[18273] = t[18272] ^ n[18273];
assign t[18274] = t[18273] ^ n[18274];
assign t[18275] = t[18274] ^ n[18275];
assign t[18276] = t[18275] ^ n[18276];
assign t[18277] = t[18276] ^ n[18277];
assign t[18278] = t[18277] ^ n[18278];
assign t[18279] = t[18278] ^ n[18279];
assign t[18280] = t[18279] ^ n[18280];
assign t[18281] = t[18280] ^ n[18281];
assign t[18282] = t[18281] ^ n[18282];
assign t[18283] = t[18282] ^ n[18283];
assign t[18284] = t[18283] ^ n[18284];
assign t[18285] = t[18284] ^ n[18285];
assign t[18286] = t[18285] ^ n[18286];
assign t[18287] = t[18286] ^ n[18287];
assign t[18288] = t[18287] ^ n[18288];
assign t[18289] = t[18288] ^ n[18289];
assign t[18290] = t[18289] ^ n[18290];
assign t[18291] = t[18290] ^ n[18291];
assign t[18292] = t[18291] ^ n[18292];
assign t[18293] = t[18292] ^ n[18293];
assign t[18294] = t[18293] ^ n[18294];
assign t[18295] = t[18294] ^ n[18295];
assign t[18296] = t[18295] ^ n[18296];
assign t[18297] = t[18296] ^ n[18297];
assign t[18298] = t[18297] ^ n[18298];
assign t[18299] = t[18298] ^ n[18299];
assign t[18300] = t[18299] ^ n[18300];
assign t[18301] = t[18300] ^ n[18301];
assign t[18302] = t[18301] ^ n[18302];
assign t[18303] = t[18302] ^ n[18303];
assign t[18304] = t[18303] ^ n[18304];
assign t[18305] = t[18304] ^ n[18305];
assign t[18306] = t[18305] ^ n[18306];
assign t[18307] = t[18306] ^ n[18307];
assign t[18308] = t[18307] ^ n[18308];
assign t[18309] = t[18308] ^ n[18309];
assign t[18310] = t[18309] ^ n[18310];
assign t[18311] = t[18310] ^ n[18311];
assign t[18312] = t[18311] ^ n[18312];
assign t[18313] = t[18312] ^ n[18313];
assign t[18314] = t[18313] ^ n[18314];
assign t[18315] = t[18314] ^ n[18315];
assign t[18316] = t[18315] ^ n[18316];
assign t[18317] = t[18316] ^ n[18317];
assign t[18318] = t[18317] ^ n[18318];
assign t[18319] = t[18318] ^ n[18319];
assign t[18320] = t[18319] ^ n[18320];
assign t[18321] = t[18320] ^ n[18321];
assign t[18322] = t[18321] ^ n[18322];
assign t[18323] = t[18322] ^ n[18323];
assign t[18324] = t[18323] ^ n[18324];
assign t[18325] = t[18324] ^ n[18325];
assign t[18326] = t[18325] ^ n[18326];
assign t[18327] = t[18326] ^ n[18327];
assign t[18328] = t[18327] ^ n[18328];
assign t[18329] = t[18328] ^ n[18329];
assign t[18330] = t[18329] ^ n[18330];
assign t[18331] = t[18330] ^ n[18331];
assign t[18332] = t[18331] ^ n[18332];
assign t[18333] = t[18332] ^ n[18333];
assign t[18334] = t[18333] ^ n[18334];
assign t[18335] = t[18334] ^ n[18335];
assign t[18336] = t[18335] ^ n[18336];
assign t[18337] = t[18336] ^ n[18337];
assign t[18338] = t[18337] ^ n[18338];
assign t[18339] = t[18338] ^ n[18339];
assign t[18340] = t[18339] ^ n[18340];
assign t[18341] = t[18340] ^ n[18341];
assign t[18342] = t[18341] ^ n[18342];
assign t[18343] = t[18342] ^ n[18343];
assign t[18344] = t[18343] ^ n[18344];
assign t[18345] = t[18344] ^ n[18345];
assign t[18346] = t[18345] ^ n[18346];
assign t[18347] = t[18346] ^ n[18347];
assign t[18348] = t[18347] ^ n[18348];
assign t[18349] = t[18348] ^ n[18349];
assign t[18350] = t[18349] ^ n[18350];
assign t[18351] = t[18350] ^ n[18351];
assign t[18352] = t[18351] ^ n[18352];
assign t[18353] = t[18352] ^ n[18353];
assign t[18354] = t[18353] ^ n[18354];
assign t[18355] = t[18354] ^ n[18355];
assign t[18356] = t[18355] ^ n[18356];
assign t[18357] = t[18356] ^ n[18357];
assign t[18358] = t[18357] ^ n[18358];
assign t[18359] = t[18358] ^ n[18359];
assign t[18360] = t[18359] ^ n[18360];
assign t[18361] = t[18360] ^ n[18361];
assign t[18362] = t[18361] ^ n[18362];
assign t[18363] = t[18362] ^ n[18363];
assign t[18364] = t[18363] ^ n[18364];
assign t[18365] = t[18364] ^ n[18365];
assign t[18366] = t[18365] ^ n[18366];
assign t[18367] = t[18366] ^ n[18367];
assign t[18368] = t[18367] ^ n[18368];
assign t[18369] = t[18368] ^ n[18369];
assign t[18370] = t[18369] ^ n[18370];
assign t[18371] = t[18370] ^ n[18371];
assign t[18372] = t[18371] ^ n[18372];
assign t[18373] = t[18372] ^ n[18373];
assign t[18374] = t[18373] ^ n[18374];
assign t[18375] = t[18374] ^ n[18375];
assign t[18376] = t[18375] ^ n[18376];
assign t[18377] = t[18376] ^ n[18377];
assign t[18378] = t[18377] ^ n[18378];
assign t[18379] = t[18378] ^ n[18379];
assign t[18380] = t[18379] ^ n[18380];
assign t[18381] = t[18380] ^ n[18381];
assign t[18382] = t[18381] ^ n[18382];
assign t[18383] = t[18382] ^ n[18383];
assign t[18384] = t[18383] ^ n[18384];
assign t[18385] = t[18384] ^ n[18385];
assign t[18386] = t[18385] ^ n[18386];
assign t[18387] = t[18386] ^ n[18387];
assign t[18388] = t[18387] ^ n[18388];
assign t[18389] = t[18388] ^ n[18389];
assign t[18390] = t[18389] ^ n[18390];
assign t[18391] = t[18390] ^ n[18391];
assign t[18392] = t[18391] ^ n[18392];
assign t[18393] = t[18392] ^ n[18393];
assign t[18394] = t[18393] ^ n[18394];
assign t[18395] = t[18394] ^ n[18395];
assign t[18396] = t[18395] ^ n[18396];
assign t[18397] = t[18396] ^ n[18397];
assign t[18398] = t[18397] ^ n[18398];
assign t[18399] = t[18398] ^ n[18399];
assign t[18400] = t[18399] ^ n[18400];
assign t[18401] = t[18400] ^ n[18401];
assign t[18402] = t[18401] ^ n[18402];
assign t[18403] = t[18402] ^ n[18403];
assign t[18404] = t[18403] ^ n[18404];
assign t[18405] = t[18404] ^ n[18405];
assign t[18406] = t[18405] ^ n[18406];
assign t[18407] = t[18406] ^ n[18407];
assign t[18408] = t[18407] ^ n[18408];
assign t[18409] = t[18408] ^ n[18409];
assign t[18410] = t[18409] ^ n[18410];
assign t[18411] = t[18410] ^ n[18411];
assign t[18412] = t[18411] ^ n[18412];
assign t[18413] = t[18412] ^ n[18413];
assign t[18414] = t[18413] ^ n[18414];
assign t[18415] = t[18414] ^ n[18415];
assign t[18416] = t[18415] ^ n[18416];
assign t[18417] = t[18416] ^ n[18417];
assign t[18418] = t[18417] ^ n[18418];
assign t[18419] = t[18418] ^ n[18419];
assign t[18420] = t[18419] ^ n[18420];
assign t[18421] = t[18420] ^ n[18421];
assign t[18422] = t[18421] ^ n[18422];
assign t[18423] = t[18422] ^ n[18423];
assign t[18424] = t[18423] ^ n[18424];
assign t[18425] = t[18424] ^ n[18425];
assign t[18426] = t[18425] ^ n[18426];
assign t[18427] = t[18426] ^ n[18427];
assign t[18428] = t[18427] ^ n[18428];
assign t[18429] = t[18428] ^ n[18429];
assign t[18430] = t[18429] ^ n[18430];
assign t[18431] = t[18430] ^ n[18431];
assign t[18432] = t[18431] ^ n[18432];
assign t[18433] = t[18432] ^ n[18433];
assign t[18434] = t[18433] ^ n[18434];
assign t[18435] = t[18434] ^ n[18435];
assign t[18436] = t[18435] ^ n[18436];
assign t[18437] = t[18436] ^ n[18437];
assign t[18438] = t[18437] ^ n[18438];
assign t[18439] = t[18438] ^ n[18439];
assign t[18440] = t[18439] ^ n[18440];
assign t[18441] = t[18440] ^ n[18441];
assign t[18442] = t[18441] ^ n[18442];
assign t[18443] = t[18442] ^ n[18443];
assign t[18444] = t[18443] ^ n[18444];
assign t[18445] = t[18444] ^ n[18445];
assign t[18446] = t[18445] ^ n[18446];
assign t[18447] = t[18446] ^ n[18447];
assign t[18448] = t[18447] ^ n[18448];
assign t[18449] = t[18448] ^ n[18449];
assign t[18450] = t[18449] ^ n[18450];
assign t[18451] = t[18450] ^ n[18451];
assign t[18452] = t[18451] ^ n[18452];
assign t[18453] = t[18452] ^ n[18453];
assign t[18454] = t[18453] ^ n[18454];
assign t[18455] = t[18454] ^ n[18455];
assign t[18456] = t[18455] ^ n[18456];
assign t[18457] = t[18456] ^ n[18457];
assign t[18458] = t[18457] ^ n[18458];
assign t[18459] = t[18458] ^ n[18459];
assign t[18460] = t[18459] ^ n[18460];
assign t[18461] = t[18460] ^ n[18461];
assign t[18462] = t[18461] ^ n[18462];
assign t[18463] = t[18462] ^ n[18463];
assign t[18464] = t[18463] ^ n[18464];
assign t[18465] = t[18464] ^ n[18465];
assign t[18466] = t[18465] ^ n[18466];
assign t[18467] = t[18466] ^ n[18467];
assign t[18468] = t[18467] ^ n[18468];
assign t[18469] = t[18468] ^ n[18469];
assign t[18470] = t[18469] ^ n[18470];
assign t[18471] = t[18470] ^ n[18471];
assign t[18472] = t[18471] ^ n[18472];
assign t[18473] = t[18472] ^ n[18473];
assign t[18474] = t[18473] ^ n[18474];
assign t[18475] = t[18474] ^ n[18475];
assign t[18476] = t[18475] ^ n[18476];
assign t[18477] = t[18476] ^ n[18477];
assign t[18478] = t[18477] ^ n[18478];
assign t[18479] = t[18478] ^ n[18479];
assign t[18480] = t[18479] ^ n[18480];
assign t[18481] = t[18480] ^ n[18481];
assign t[18482] = t[18481] ^ n[18482];
assign t[18483] = t[18482] ^ n[18483];
assign t[18484] = t[18483] ^ n[18484];
assign t[18485] = t[18484] ^ n[18485];
assign t[18486] = t[18485] ^ n[18486];
assign t[18487] = t[18486] ^ n[18487];
assign t[18488] = t[18487] ^ n[18488];
assign t[18489] = t[18488] ^ n[18489];
assign t[18490] = t[18489] ^ n[18490];
assign t[18491] = t[18490] ^ n[18491];
assign t[18492] = t[18491] ^ n[18492];
assign t[18493] = t[18492] ^ n[18493];
assign t[18494] = t[18493] ^ n[18494];
assign t[18495] = t[18494] ^ n[18495];
assign t[18496] = t[18495] ^ n[18496];
assign t[18497] = t[18496] ^ n[18497];
assign t[18498] = t[18497] ^ n[18498];
assign t[18499] = t[18498] ^ n[18499];
assign t[18500] = t[18499] ^ n[18500];
assign t[18501] = t[18500] ^ n[18501];
assign t[18502] = t[18501] ^ n[18502];
assign t[18503] = t[18502] ^ n[18503];
assign t[18504] = t[18503] ^ n[18504];
assign t[18505] = t[18504] ^ n[18505];
assign t[18506] = t[18505] ^ n[18506];
assign t[18507] = t[18506] ^ n[18507];
assign t[18508] = t[18507] ^ n[18508];
assign t[18509] = t[18508] ^ n[18509];
assign t[18510] = t[18509] ^ n[18510];
assign t[18511] = t[18510] ^ n[18511];
assign t[18512] = t[18511] ^ n[18512];
assign t[18513] = t[18512] ^ n[18513];
assign t[18514] = t[18513] ^ n[18514];
assign t[18515] = t[18514] ^ n[18515];
assign t[18516] = t[18515] ^ n[18516];
assign t[18517] = t[18516] ^ n[18517];
assign t[18518] = t[18517] ^ n[18518];
assign t[18519] = t[18518] ^ n[18519];
assign t[18520] = t[18519] ^ n[18520];
assign t[18521] = t[18520] ^ n[18521];
assign t[18522] = t[18521] ^ n[18522];
assign t[18523] = t[18522] ^ n[18523];
assign t[18524] = t[18523] ^ n[18524];
assign t[18525] = t[18524] ^ n[18525];
assign t[18526] = t[18525] ^ n[18526];
assign t[18527] = t[18526] ^ n[18527];
assign t[18528] = t[18527] ^ n[18528];
assign t[18529] = t[18528] ^ n[18529];
assign t[18530] = t[18529] ^ n[18530];
assign t[18531] = t[18530] ^ n[18531];
assign t[18532] = t[18531] ^ n[18532];
assign t[18533] = t[18532] ^ n[18533];
assign t[18534] = t[18533] ^ n[18534];
assign t[18535] = t[18534] ^ n[18535];
assign t[18536] = t[18535] ^ n[18536];
assign t[18537] = t[18536] ^ n[18537];
assign t[18538] = t[18537] ^ n[18538];
assign t[18539] = t[18538] ^ n[18539];
assign t[18540] = t[18539] ^ n[18540];
assign t[18541] = t[18540] ^ n[18541];
assign t[18542] = t[18541] ^ n[18542];
assign t[18543] = t[18542] ^ n[18543];
assign t[18544] = t[18543] ^ n[18544];
assign t[18545] = t[18544] ^ n[18545];
assign t[18546] = t[18545] ^ n[18546];
assign t[18547] = t[18546] ^ n[18547];
assign t[18548] = t[18547] ^ n[18548];
assign t[18549] = t[18548] ^ n[18549];
assign t[18550] = t[18549] ^ n[18550];
assign t[18551] = t[18550] ^ n[18551];
assign t[18552] = t[18551] ^ n[18552];
assign t[18553] = t[18552] ^ n[18553];
assign t[18554] = t[18553] ^ n[18554];
assign t[18555] = t[18554] ^ n[18555];
assign t[18556] = t[18555] ^ n[18556];
assign t[18557] = t[18556] ^ n[18557];
assign t[18558] = t[18557] ^ n[18558];
assign t[18559] = t[18558] ^ n[18559];
assign t[18560] = t[18559] ^ n[18560];
assign t[18561] = t[18560] ^ n[18561];
assign t[18562] = t[18561] ^ n[18562];
assign t[18563] = t[18562] ^ n[18563];
assign t[18564] = t[18563] ^ n[18564];
assign t[18565] = t[18564] ^ n[18565];
assign t[18566] = t[18565] ^ n[18566];
assign t[18567] = t[18566] ^ n[18567];
assign t[18568] = t[18567] ^ n[18568];
assign t[18569] = t[18568] ^ n[18569];
assign t[18570] = t[18569] ^ n[18570];
assign t[18571] = t[18570] ^ n[18571];
assign t[18572] = t[18571] ^ n[18572];
assign t[18573] = t[18572] ^ n[18573];
assign t[18574] = t[18573] ^ n[18574];
assign t[18575] = t[18574] ^ n[18575];
assign t[18576] = t[18575] ^ n[18576];
assign t[18577] = t[18576] ^ n[18577];
assign t[18578] = t[18577] ^ n[18578];
assign t[18579] = t[18578] ^ n[18579];
assign t[18580] = t[18579] ^ n[18580];
assign t[18581] = t[18580] ^ n[18581];
assign t[18582] = t[18581] ^ n[18582];
assign t[18583] = t[18582] ^ n[18583];
assign t[18584] = t[18583] ^ n[18584];
assign t[18585] = t[18584] ^ n[18585];
assign t[18586] = t[18585] ^ n[18586];
assign t[18587] = t[18586] ^ n[18587];
assign t[18588] = t[18587] ^ n[18588];
assign t[18589] = t[18588] ^ n[18589];
assign t[18590] = t[18589] ^ n[18590];
assign t[18591] = t[18590] ^ n[18591];
assign t[18592] = t[18591] ^ n[18592];
assign t[18593] = t[18592] ^ n[18593];
assign t[18594] = t[18593] ^ n[18594];
assign t[18595] = t[18594] ^ n[18595];
assign t[18596] = t[18595] ^ n[18596];
assign t[18597] = t[18596] ^ n[18597];
assign t[18598] = t[18597] ^ n[18598];
assign t[18599] = t[18598] ^ n[18599];
assign t[18600] = t[18599] ^ n[18600];
assign t[18601] = t[18600] ^ n[18601];
assign t[18602] = t[18601] ^ n[18602];
assign t[18603] = t[18602] ^ n[18603];
assign t[18604] = t[18603] ^ n[18604];
assign t[18605] = t[18604] ^ n[18605];
assign t[18606] = t[18605] ^ n[18606];
assign t[18607] = t[18606] ^ n[18607];
assign t[18608] = t[18607] ^ n[18608];
assign t[18609] = t[18608] ^ n[18609];
assign t[18610] = t[18609] ^ n[18610];
assign t[18611] = t[18610] ^ n[18611];
assign t[18612] = t[18611] ^ n[18612];
assign t[18613] = t[18612] ^ n[18613];
assign t[18614] = t[18613] ^ n[18614];
assign t[18615] = t[18614] ^ n[18615];
assign t[18616] = t[18615] ^ n[18616];
assign t[18617] = t[18616] ^ n[18617];
assign t[18618] = t[18617] ^ n[18618];
assign t[18619] = t[18618] ^ n[18619];
assign t[18620] = t[18619] ^ n[18620];
assign t[18621] = t[18620] ^ n[18621];
assign t[18622] = t[18621] ^ n[18622];
assign t[18623] = t[18622] ^ n[18623];
assign t[18624] = t[18623] ^ n[18624];
assign t[18625] = t[18624] ^ n[18625];
assign t[18626] = t[18625] ^ n[18626];
assign t[18627] = t[18626] ^ n[18627];
assign t[18628] = t[18627] ^ n[18628];
assign t[18629] = t[18628] ^ n[18629];
assign t[18630] = t[18629] ^ n[18630];
assign t[18631] = t[18630] ^ n[18631];
assign t[18632] = t[18631] ^ n[18632];
assign t[18633] = t[18632] ^ n[18633];
assign t[18634] = t[18633] ^ n[18634];
assign t[18635] = t[18634] ^ n[18635];
assign t[18636] = t[18635] ^ n[18636];
assign t[18637] = t[18636] ^ n[18637];
assign t[18638] = t[18637] ^ n[18638];
assign t[18639] = t[18638] ^ n[18639];
assign t[18640] = t[18639] ^ n[18640];
assign t[18641] = t[18640] ^ n[18641];
assign t[18642] = t[18641] ^ n[18642];
assign t[18643] = t[18642] ^ n[18643];
assign t[18644] = t[18643] ^ n[18644];
assign t[18645] = t[18644] ^ n[18645];
assign t[18646] = t[18645] ^ n[18646];
assign t[18647] = t[18646] ^ n[18647];
assign t[18648] = t[18647] ^ n[18648];
assign t[18649] = t[18648] ^ n[18649];
assign t[18650] = t[18649] ^ n[18650];
assign t[18651] = t[18650] ^ n[18651];
assign t[18652] = t[18651] ^ n[18652];
assign t[18653] = t[18652] ^ n[18653];
assign t[18654] = t[18653] ^ n[18654];
assign t[18655] = t[18654] ^ n[18655];
assign t[18656] = t[18655] ^ n[18656];
assign t[18657] = t[18656] ^ n[18657];
assign t[18658] = t[18657] ^ n[18658];
assign t[18659] = t[18658] ^ n[18659];
assign t[18660] = t[18659] ^ n[18660];
assign t[18661] = t[18660] ^ n[18661];
assign t[18662] = t[18661] ^ n[18662];
assign t[18663] = t[18662] ^ n[18663];
assign t[18664] = t[18663] ^ n[18664];
assign t[18665] = t[18664] ^ n[18665];
assign t[18666] = t[18665] ^ n[18666];
assign t[18667] = t[18666] ^ n[18667];
assign t[18668] = t[18667] ^ n[18668];
assign t[18669] = t[18668] ^ n[18669];
assign t[18670] = t[18669] ^ n[18670];
assign t[18671] = t[18670] ^ n[18671];
assign t[18672] = t[18671] ^ n[18672];
assign t[18673] = t[18672] ^ n[18673];
assign t[18674] = t[18673] ^ n[18674];
assign t[18675] = t[18674] ^ n[18675];
assign t[18676] = t[18675] ^ n[18676];
assign t[18677] = t[18676] ^ n[18677];
assign t[18678] = t[18677] ^ n[18678];
assign t[18679] = t[18678] ^ n[18679];
assign t[18680] = t[18679] ^ n[18680];
assign t[18681] = t[18680] ^ n[18681];
assign t[18682] = t[18681] ^ n[18682];
assign t[18683] = t[18682] ^ n[18683];
assign t[18684] = t[18683] ^ n[18684];
assign t[18685] = t[18684] ^ n[18685];
assign t[18686] = t[18685] ^ n[18686];
assign t[18687] = t[18686] ^ n[18687];
assign t[18688] = t[18687] ^ n[18688];
assign t[18689] = t[18688] ^ n[18689];
assign t[18690] = t[18689] ^ n[18690];
assign t[18691] = t[18690] ^ n[18691];
assign t[18692] = t[18691] ^ n[18692];
assign t[18693] = t[18692] ^ n[18693];
assign t[18694] = t[18693] ^ n[18694];
assign t[18695] = t[18694] ^ n[18695];
assign t[18696] = t[18695] ^ n[18696];
assign t[18697] = t[18696] ^ n[18697];
assign t[18698] = t[18697] ^ n[18698];
assign t[18699] = t[18698] ^ n[18699];
assign t[18700] = t[18699] ^ n[18700];
assign t[18701] = t[18700] ^ n[18701];
assign t[18702] = t[18701] ^ n[18702];
assign t[18703] = t[18702] ^ n[18703];
assign t[18704] = t[18703] ^ n[18704];
assign t[18705] = t[18704] ^ n[18705];
assign t[18706] = t[18705] ^ n[18706];
assign t[18707] = t[18706] ^ n[18707];
assign t[18708] = t[18707] ^ n[18708];
assign t[18709] = t[18708] ^ n[18709];
assign t[18710] = t[18709] ^ n[18710];
assign t[18711] = t[18710] ^ n[18711];
assign t[18712] = t[18711] ^ n[18712];
assign t[18713] = t[18712] ^ n[18713];
assign t[18714] = t[18713] ^ n[18714];
assign t[18715] = t[18714] ^ n[18715];
assign t[18716] = t[18715] ^ n[18716];
assign t[18717] = t[18716] ^ n[18717];
assign t[18718] = t[18717] ^ n[18718];
assign t[18719] = t[18718] ^ n[18719];
assign t[18720] = t[18719] ^ n[18720];
assign t[18721] = t[18720] ^ n[18721];
assign t[18722] = t[18721] ^ n[18722];
assign t[18723] = t[18722] ^ n[18723];
assign t[18724] = t[18723] ^ n[18724];
assign t[18725] = t[18724] ^ n[18725];
assign t[18726] = t[18725] ^ n[18726];
assign t[18727] = t[18726] ^ n[18727];
assign t[18728] = t[18727] ^ n[18728];
assign t[18729] = t[18728] ^ n[18729];
assign t[18730] = t[18729] ^ n[18730];
assign t[18731] = t[18730] ^ n[18731];
assign t[18732] = t[18731] ^ n[18732];
assign t[18733] = t[18732] ^ n[18733];
assign t[18734] = t[18733] ^ n[18734];
assign t[18735] = t[18734] ^ n[18735];
assign t[18736] = t[18735] ^ n[18736];
assign t[18737] = t[18736] ^ n[18737];
assign t[18738] = t[18737] ^ n[18738];
assign t[18739] = t[18738] ^ n[18739];
assign t[18740] = t[18739] ^ n[18740];
assign t[18741] = t[18740] ^ n[18741];
assign t[18742] = t[18741] ^ n[18742];
assign t[18743] = t[18742] ^ n[18743];
assign t[18744] = t[18743] ^ n[18744];
assign t[18745] = t[18744] ^ n[18745];
assign t[18746] = t[18745] ^ n[18746];
assign t[18747] = t[18746] ^ n[18747];
assign t[18748] = t[18747] ^ n[18748];
assign t[18749] = t[18748] ^ n[18749];
assign t[18750] = t[18749] ^ n[18750];
assign t[18751] = t[18750] ^ n[18751];
assign t[18752] = t[18751] ^ n[18752];
assign t[18753] = t[18752] ^ n[18753];
assign t[18754] = t[18753] ^ n[18754];
assign t[18755] = t[18754] ^ n[18755];
assign t[18756] = t[18755] ^ n[18756];
assign t[18757] = t[18756] ^ n[18757];
assign t[18758] = t[18757] ^ n[18758];
assign t[18759] = t[18758] ^ n[18759];
assign t[18760] = t[18759] ^ n[18760];
assign t[18761] = t[18760] ^ n[18761];
assign t[18762] = t[18761] ^ n[18762];
assign t[18763] = t[18762] ^ n[18763];
assign t[18764] = t[18763] ^ n[18764];
assign t[18765] = t[18764] ^ n[18765];
assign t[18766] = t[18765] ^ n[18766];
assign t[18767] = t[18766] ^ n[18767];
assign t[18768] = t[18767] ^ n[18768];
assign t[18769] = t[18768] ^ n[18769];
assign t[18770] = t[18769] ^ n[18770];
assign t[18771] = t[18770] ^ n[18771];
assign t[18772] = t[18771] ^ n[18772];
assign t[18773] = t[18772] ^ n[18773];
assign t[18774] = t[18773] ^ n[18774];
assign t[18775] = t[18774] ^ n[18775];
assign t[18776] = t[18775] ^ n[18776];
assign t[18777] = t[18776] ^ n[18777];
assign t[18778] = t[18777] ^ n[18778];
assign t[18779] = t[18778] ^ n[18779];
assign t[18780] = t[18779] ^ n[18780];
assign t[18781] = t[18780] ^ n[18781];
assign t[18782] = t[18781] ^ n[18782];
assign t[18783] = t[18782] ^ n[18783];
assign t[18784] = t[18783] ^ n[18784];
assign t[18785] = t[18784] ^ n[18785];
assign t[18786] = t[18785] ^ n[18786];
assign t[18787] = t[18786] ^ n[18787];
assign t[18788] = t[18787] ^ n[18788];
assign t[18789] = t[18788] ^ n[18789];
assign t[18790] = t[18789] ^ n[18790];
assign t[18791] = t[18790] ^ n[18791];
assign t[18792] = t[18791] ^ n[18792];
assign t[18793] = t[18792] ^ n[18793];
assign t[18794] = t[18793] ^ n[18794];
assign t[18795] = t[18794] ^ n[18795];
assign t[18796] = t[18795] ^ n[18796];
assign t[18797] = t[18796] ^ n[18797];
assign t[18798] = t[18797] ^ n[18798];
assign t[18799] = t[18798] ^ n[18799];
assign t[18800] = t[18799] ^ n[18800];
assign t[18801] = t[18800] ^ n[18801];
assign t[18802] = t[18801] ^ n[18802];
assign t[18803] = t[18802] ^ n[18803];
assign t[18804] = t[18803] ^ n[18804];
assign t[18805] = t[18804] ^ n[18805];
assign t[18806] = t[18805] ^ n[18806];
assign t[18807] = t[18806] ^ n[18807];
assign t[18808] = t[18807] ^ n[18808];
assign t[18809] = t[18808] ^ n[18809];
assign t[18810] = t[18809] ^ n[18810];
assign t[18811] = t[18810] ^ n[18811];
assign t[18812] = t[18811] ^ n[18812];
assign t[18813] = t[18812] ^ n[18813];
assign t[18814] = t[18813] ^ n[18814];
assign t[18815] = t[18814] ^ n[18815];
assign t[18816] = t[18815] ^ n[18816];
assign t[18817] = t[18816] ^ n[18817];
assign t[18818] = t[18817] ^ n[18818];
assign t[18819] = t[18818] ^ n[18819];
assign t[18820] = t[18819] ^ n[18820];
assign t[18821] = t[18820] ^ n[18821];
assign t[18822] = t[18821] ^ n[18822];
assign t[18823] = t[18822] ^ n[18823];
assign t[18824] = t[18823] ^ n[18824];
assign t[18825] = t[18824] ^ n[18825];
assign t[18826] = t[18825] ^ n[18826];
assign t[18827] = t[18826] ^ n[18827];
assign t[18828] = t[18827] ^ n[18828];
assign t[18829] = t[18828] ^ n[18829];
assign t[18830] = t[18829] ^ n[18830];
assign t[18831] = t[18830] ^ n[18831];
assign t[18832] = t[18831] ^ n[18832];
assign t[18833] = t[18832] ^ n[18833];
assign t[18834] = t[18833] ^ n[18834];
assign t[18835] = t[18834] ^ n[18835];
assign t[18836] = t[18835] ^ n[18836];
assign t[18837] = t[18836] ^ n[18837];
assign t[18838] = t[18837] ^ n[18838];
assign t[18839] = t[18838] ^ n[18839];
assign t[18840] = t[18839] ^ n[18840];
assign t[18841] = t[18840] ^ n[18841];
assign t[18842] = t[18841] ^ n[18842];
assign t[18843] = t[18842] ^ n[18843];
assign t[18844] = t[18843] ^ n[18844];
assign t[18845] = t[18844] ^ n[18845];
assign t[18846] = t[18845] ^ n[18846];
assign t[18847] = t[18846] ^ n[18847];
assign t[18848] = t[18847] ^ n[18848];
assign t[18849] = t[18848] ^ n[18849];
assign t[18850] = t[18849] ^ n[18850];
assign t[18851] = t[18850] ^ n[18851];
assign t[18852] = t[18851] ^ n[18852];
assign t[18853] = t[18852] ^ n[18853];
assign t[18854] = t[18853] ^ n[18854];
assign t[18855] = t[18854] ^ n[18855];
assign t[18856] = t[18855] ^ n[18856];
assign t[18857] = t[18856] ^ n[18857];
assign t[18858] = t[18857] ^ n[18858];
assign t[18859] = t[18858] ^ n[18859];
assign t[18860] = t[18859] ^ n[18860];
assign t[18861] = t[18860] ^ n[18861];
assign t[18862] = t[18861] ^ n[18862];
assign t[18863] = t[18862] ^ n[18863];
assign t[18864] = t[18863] ^ n[18864];
assign t[18865] = t[18864] ^ n[18865];
assign t[18866] = t[18865] ^ n[18866];
assign t[18867] = t[18866] ^ n[18867];
assign t[18868] = t[18867] ^ n[18868];
assign t[18869] = t[18868] ^ n[18869];
assign t[18870] = t[18869] ^ n[18870];
assign t[18871] = t[18870] ^ n[18871];
assign t[18872] = t[18871] ^ n[18872];
assign t[18873] = t[18872] ^ n[18873];
assign t[18874] = t[18873] ^ n[18874];
assign t[18875] = t[18874] ^ n[18875];
assign t[18876] = t[18875] ^ n[18876];
assign t[18877] = t[18876] ^ n[18877];
assign t[18878] = t[18877] ^ n[18878];
assign t[18879] = t[18878] ^ n[18879];
assign t[18880] = t[18879] ^ n[18880];
assign t[18881] = t[18880] ^ n[18881];
assign t[18882] = t[18881] ^ n[18882];
assign t[18883] = t[18882] ^ n[18883];
assign t[18884] = t[18883] ^ n[18884];
assign t[18885] = t[18884] ^ n[18885];
assign t[18886] = t[18885] ^ n[18886];
assign t[18887] = t[18886] ^ n[18887];
assign t[18888] = t[18887] ^ n[18888];
assign t[18889] = t[18888] ^ n[18889];
assign t[18890] = t[18889] ^ n[18890];
assign t[18891] = t[18890] ^ n[18891];
assign t[18892] = t[18891] ^ n[18892];
assign t[18893] = t[18892] ^ n[18893];
assign t[18894] = t[18893] ^ n[18894];
assign t[18895] = t[18894] ^ n[18895];
assign t[18896] = t[18895] ^ n[18896];
assign t[18897] = t[18896] ^ n[18897];
assign t[18898] = t[18897] ^ n[18898];
assign t[18899] = t[18898] ^ n[18899];
assign t[18900] = t[18899] ^ n[18900];
assign t[18901] = t[18900] ^ n[18901];
assign t[18902] = t[18901] ^ n[18902];
assign t[18903] = t[18902] ^ n[18903];
assign t[18904] = t[18903] ^ n[18904];
assign t[18905] = t[18904] ^ n[18905];
assign t[18906] = t[18905] ^ n[18906];
assign t[18907] = t[18906] ^ n[18907];
assign t[18908] = t[18907] ^ n[18908];
assign t[18909] = t[18908] ^ n[18909];
assign t[18910] = t[18909] ^ n[18910];
assign t[18911] = t[18910] ^ n[18911];
assign t[18912] = t[18911] ^ n[18912];
assign t[18913] = t[18912] ^ n[18913];
assign t[18914] = t[18913] ^ n[18914];
assign t[18915] = t[18914] ^ n[18915];
assign t[18916] = t[18915] ^ n[18916];
assign t[18917] = t[18916] ^ n[18917];
assign t[18918] = t[18917] ^ n[18918];
assign t[18919] = t[18918] ^ n[18919];
assign t[18920] = t[18919] ^ n[18920];
assign t[18921] = t[18920] ^ n[18921];
assign t[18922] = t[18921] ^ n[18922];
assign t[18923] = t[18922] ^ n[18923];
assign t[18924] = t[18923] ^ n[18924];
assign t[18925] = t[18924] ^ n[18925];
assign t[18926] = t[18925] ^ n[18926];
assign t[18927] = t[18926] ^ n[18927];
assign t[18928] = t[18927] ^ n[18928];
assign t[18929] = t[18928] ^ n[18929];
assign t[18930] = t[18929] ^ n[18930];
assign t[18931] = t[18930] ^ n[18931];
assign t[18932] = t[18931] ^ n[18932];
assign t[18933] = t[18932] ^ n[18933];
assign t[18934] = t[18933] ^ n[18934];
assign t[18935] = t[18934] ^ n[18935];
assign t[18936] = t[18935] ^ n[18936];
assign t[18937] = t[18936] ^ n[18937];
assign t[18938] = t[18937] ^ n[18938];
assign t[18939] = t[18938] ^ n[18939];
assign t[18940] = t[18939] ^ n[18940];
assign t[18941] = t[18940] ^ n[18941];
assign t[18942] = t[18941] ^ n[18942];
assign t[18943] = t[18942] ^ n[18943];
assign t[18944] = t[18943] ^ n[18944];
assign t[18945] = t[18944] ^ n[18945];
assign t[18946] = t[18945] ^ n[18946];
assign t[18947] = t[18946] ^ n[18947];
assign t[18948] = t[18947] ^ n[18948];
assign t[18949] = t[18948] ^ n[18949];
assign t[18950] = t[18949] ^ n[18950];
assign t[18951] = t[18950] ^ n[18951];
assign t[18952] = t[18951] ^ n[18952];
assign t[18953] = t[18952] ^ n[18953];
assign t[18954] = t[18953] ^ n[18954];
assign t[18955] = t[18954] ^ n[18955];
assign t[18956] = t[18955] ^ n[18956];
assign t[18957] = t[18956] ^ n[18957];
assign t[18958] = t[18957] ^ n[18958];
assign t[18959] = t[18958] ^ n[18959];
assign t[18960] = t[18959] ^ n[18960];
assign t[18961] = t[18960] ^ n[18961];
assign t[18962] = t[18961] ^ n[18962];
assign t[18963] = t[18962] ^ n[18963];
assign t[18964] = t[18963] ^ n[18964];
assign t[18965] = t[18964] ^ n[18965];
assign t[18966] = t[18965] ^ n[18966];
assign t[18967] = t[18966] ^ n[18967];
assign t[18968] = t[18967] ^ n[18968];
assign t[18969] = t[18968] ^ n[18969];
assign t[18970] = t[18969] ^ n[18970];
assign t[18971] = t[18970] ^ n[18971];
assign t[18972] = t[18971] ^ n[18972];
assign t[18973] = t[18972] ^ n[18973];
assign t[18974] = t[18973] ^ n[18974];
assign t[18975] = t[18974] ^ n[18975];
assign t[18976] = t[18975] ^ n[18976];
assign t[18977] = t[18976] ^ n[18977];
assign t[18978] = t[18977] ^ n[18978];
assign t[18979] = t[18978] ^ n[18979];
assign t[18980] = t[18979] ^ n[18980];
assign t[18981] = t[18980] ^ n[18981];
assign t[18982] = t[18981] ^ n[18982];
assign t[18983] = t[18982] ^ n[18983];
assign t[18984] = t[18983] ^ n[18984];
assign t[18985] = t[18984] ^ n[18985];
assign t[18986] = t[18985] ^ n[18986];
assign t[18987] = t[18986] ^ n[18987];
assign t[18988] = t[18987] ^ n[18988];
assign t[18989] = t[18988] ^ n[18989];
assign t[18990] = t[18989] ^ n[18990];
assign t[18991] = t[18990] ^ n[18991];
assign t[18992] = t[18991] ^ n[18992];
assign t[18993] = t[18992] ^ n[18993];
assign t[18994] = t[18993] ^ n[18994];
assign t[18995] = t[18994] ^ n[18995];
assign t[18996] = t[18995] ^ n[18996];
assign t[18997] = t[18996] ^ n[18997];
assign t[18998] = t[18997] ^ n[18998];
assign t[18999] = t[18998] ^ n[18999];
assign t[19000] = t[18999] ^ n[19000];
assign t[19001] = t[19000] ^ n[19001];
assign t[19002] = t[19001] ^ n[19002];
assign t[19003] = t[19002] ^ n[19003];
assign t[19004] = t[19003] ^ n[19004];
assign t[19005] = t[19004] ^ n[19005];
assign t[19006] = t[19005] ^ n[19006];
assign t[19007] = t[19006] ^ n[19007];
assign t[19008] = t[19007] ^ n[19008];
assign t[19009] = t[19008] ^ n[19009];
assign t[19010] = t[19009] ^ n[19010];
assign t[19011] = t[19010] ^ n[19011];
assign t[19012] = t[19011] ^ n[19012];
assign t[19013] = t[19012] ^ n[19013];
assign t[19014] = t[19013] ^ n[19014];
assign t[19015] = t[19014] ^ n[19015];
assign t[19016] = t[19015] ^ n[19016];
assign t[19017] = t[19016] ^ n[19017];
assign t[19018] = t[19017] ^ n[19018];
assign t[19019] = t[19018] ^ n[19019];
assign t[19020] = t[19019] ^ n[19020];
assign t[19021] = t[19020] ^ n[19021];
assign t[19022] = t[19021] ^ n[19022];
assign t[19023] = t[19022] ^ n[19023];
assign t[19024] = t[19023] ^ n[19024];
assign t[19025] = t[19024] ^ n[19025];
assign t[19026] = t[19025] ^ n[19026];
assign t[19027] = t[19026] ^ n[19027];
assign t[19028] = t[19027] ^ n[19028];
assign t[19029] = t[19028] ^ n[19029];
assign t[19030] = t[19029] ^ n[19030];
assign t[19031] = t[19030] ^ n[19031];
assign t[19032] = t[19031] ^ n[19032];
assign t[19033] = t[19032] ^ n[19033];
assign t[19034] = t[19033] ^ n[19034];
assign t[19035] = t[19034] ^ n[19035];
assign t[19036] = t[19035] ^ n[19036];
assign t[19037] = t[19036] ^ n[19037];
assign t[19038] = t[19037] ^ n[19038];
assign t[19039] = t[19038] ^ n[19039];
assign t[19040] = t[19039] ^ n[19040];
assign t[19041] = t[19040] ^ n[19041];
assign t[19042] = t[19041] ^ n[19042];
assign t[19043] = t[19042] ^ n[19043];
assign t[19044] = t[19043] ^ n[19044];
assign t[19045] = t[19044] ^ n[19045];
assign t[19046] = t[19045] ^ n[19046];
assign t[19047] = t[19046] ^ n[19047];
assign t[19048] = t[19047] ^ n[19048];
assign t[19049] = t[19048] ^ n[19049];
assign t[19050] = t[19049] ^ n[19050];
assign t[19051] = t[19050] ^ n[19051];
assign t[19052] = t[19051] ^ n[19052];
assign t[19053] = t[19052] ^ n[19053];
assign t[19054] = t[19053] ^ n[19054];
assign t[19055] = t[19054] ^ n[19055];
assign t[19056] = t[19055] ^ n[19056];
assign t[19057] = t[19056] ^ n[19057];
assign t[19058] = t[19057] ^ n[19058];
assign t[19059] = t[19058] ^ n[19059];
assign t[19060] = t[19059] ^ n[19060];
assign t[19061] = t[19060] ^ n[19061];
assign t[19062] = t[19061] ^ n[19062];
assign t[19063] = t[19062] ^ n[19063];
assign t[19064] = t[19063] ^ n[19064];
assign t[19065] = t[19064] ^ n[19065];
assign t[19066] = t[19065] ^ n[19066];
assign t[19067] = t[19066] ^ n[19067];
assign t[19068] = t[19067] ^ n[19068];
assign t[19069] = t[19068] ^ n[19069];
assign t[19070] = t[19069] ^ n[19070];
assign t[19071] = t[19070] ^ n[19071];
assign t[19072] = t[19071] ^ n[19072];
assign t[19073] = t[19072] ^ n[19073];
assign t[19074] = t[19073] ^ n[19074];
assign t[19075] = t[19074] ^ n[19075];
assign t[19076] = t[19075] ^ n[19076];
assign t[19077] = t[19076] ^ n[19077];
assign t[19078] = t[19077] ^ n[19078];
assign t[19079] = t[19078] ^ n[19079];
assign t[19080] = t[19079] ^ n[19080];
assign t[19081] = t[19080] ^ n[19081];
assign t[19082] = t[19081] ^ n[19082];
assign t[19083] = t[19082] ^ n[19083];
assign t[19084] = t[19083] ^ n[19084];
assign t[19085] = t[19084] ^ n[19085];
assign t[19086] = t[19085] ^ n[19086];
assign t[19087] = t[19086] ^ n[19087];
assign t[19088] = t[19087] ^ n[19088];
assign t[19089] = t[19088] ^ n[19089];
assign t[19090] = t[19089] ^ n[19090];
assign t[19091] = t[19090] ^ n[19091];
assign t[19092] = t[19091] ^ n[19092];
assign t[19093] = t[19092] ^ n[19093];
assign t[19094] = t[19093] ^ n[19094];
assign t[19095] = t[19094] ^ n[19095];
assign t[19096] = t[19095] ^ n[19096];
assign t[19097] = t[19096] ^ n[19097];
assign t[19098] = t[19097] ^ n[19098];
assign t[19099] = t[19098] ^ n[19099];
assign t[19100] = t[19099] ^ n[19100];
assign t[19101] = t[19100] ^ n[19101];
assign t[19102] = t[19101] ^ n[19102];
assign t[19103] = t[19102] ^ n[19103];
assign t[19104] = t[19103] ^ n[19104];
assign t[19105] = t[19104] ^ n[19105];
assign t[19106] = t[19105] ^ n[19106];
assign t[19107] = t[19106] ^ n[19107];
assign t[19108] = t[19107] ^ n[19108];
assign t[19109] = t[19108] ^ n[19109];
assign t[19110] = t[19109] ^ n[19110];
assign t[19111] = t[19110] ^ n[19111];
assign t[19112] = t[19111] ^ n[19112];
assign t[19113] = t[19112] ^ n[19113];
assign t[19114] = t[19113] ^ n[19114];
assign t[19115] = t[19114] ^ n[19115];
assign t[19116] = t[19115] ^ n[19116];
assign t[19117] = t[19116] ^ n[19117];
assign t[19118] = t[19117] ^ n[19118];
assign t[19119] = t[19118] ^ n[19119];
assign t[19120] = t[19119] ^ n[19120];
assign t[19121] = t[19120] ^ n[19121];
assign t[19122] = t[19121] ^ n[19122];
assign t[19123] = t[19122] ^ n[19123];
assign t[19124] = t[19123] ^ n[19124];
assign t[19125] = t[19124] ^ n[19125];
assign t[19126] = t[19125] ^ n[19126];
assign t[19127] = t[19126] ^ n[19127];
assign t[19128] = t[19127] ^ n[19128];
assign t[19129] = t[19128] ^ n[19129];
assign t[19130] = t[19129] ^ n[19130];
assign t[19131] = t[19130] ^ n[19131];
assign t[19132] = t[19131] ^ n[19132];
assign t[19133] = t[19132] ^ n[19133];
assign t[19134] = t[19133] ^ n[19134];
assign t[19135] = t[19134] ^ n[19135];
assign t[19136] = t[19135] ^ n[19136];
assign t[19137] = t[19136] ^ n[19137];
assign t[19138] = t[19137] ^ n[19138];
assign t[19139] = t[19138] ^ n[19139];
assign t[19140] = t[19139] ^ n[19140];
assign t[19141] = t[19140] ^ n[19141];
assign t[19142] = t[19141] ^ n[19142];
assign t[19143] = t[19142] ^ n[19143];
assign t[19144] = t[19143] ^ n[19144];
assign t[19145] = t[19144] ^ n[19145];
assign t[19146] = t[19145] ^ n[19146];
assign t[19147] = t[19146] ^ n[19147];
assign t[19148] = t[19147] ^ n[19148];
assign t[19149] = t[19148] ^ n[19149];
assign t[19150] = t[19149] ^ n[19150];
assign t[19151] = t[19150] ^ n[19151];
assign t[19152] = t[19151] ^ n[19152];
assign t[19153] = t[19152] ^ n[19153];
assign t[19154] = t[19153] ^ n[19154];
assign t[19155] = t[19154] ^ n[19155];
assign t[19156] = t[19155] ^ n[19156];
assign t[19157] = t[19156] ^ n[19157];
assign t[19158] = t[19157] ^ n[19158];
assign t[19159] = t[19158] ^ n[19159];
assign t[19160] = t[19159] ^ n[19160];
assign t[19161] = t[19160] ^ n[19161];
assign t[19162] = t[19161] ^ n[19162];
assign t[19163] = t[19162] ^ n[19163];
assign t[19164] = t[19163] ^ n[19164];
assign t[19165] = t[19164] ^ n[19165];
assign t[19166] = t[19165] ^ n[19166];
assign t[19167] = t[19166] ^ n[19167];
assign t[19168] = t[19167] ^ n[19168];
assign t[19169] = t[19168] ^ n[19169];
assign t[19170] = t[19169] ^ n[19170];
assign t[19171] = t[19170] ^ n[19171];
assign t[19172] = t[19171] ^ n[19172];
assign t[19173] = t[19172] ^ n[19173];
assign t[19174] = t[19173] ^ n[19174];
assign t[19175] = t[19174] ^ n[19175];
assign t[19176] = t[19175] ^ n[19176];
assign t[19177] = t[19176] ^ n[19177];
assign t[19178] = t[19177] ^ n[19178];
assign t[19179] = t[19178] ^ n[19179];
assign t[19180] = t[19179] ^ n[19180];
assign t[19181] = t[19180] ^ n[19181];
assign t[19182] = t[19181] ^ n[19182];
assign t[19183] = t[19182] ^ n[19183];
assign t[19184] = t[19183] ^ n[19184];
assign t[19185] = t[19184] ^ n[19185];
assign t[19186] = t[19185] ^ n[19186];
assign t[19187] = t[19186] ^ n[19187];
assign t[19188] = t[19187] ^ n[19188];
assign t[19189] = t[19188] ^ n[19189];
assign t[19190] = t[19189] ^ n[19190];
assign t[19191] = t[19190] ^ n[19191];
assign t[19192] = t[19191] ^ n[19192];
assign t[19193] = t[19192] ^ n[19193];
assign t[19194] = t[19193] ^ n[19194];
assign t[19195] = t[19194] ^ n[19195];
assign t[19196] = t[19195] ^ n[19196];
assign t[19197] = t[19196] ^ n[19197];
assign t[19198] = t[19197] ^ n[19198];
assign t[19199] = t[19198] ^ n[19199];
assign t[19200] = t[19199] ^ n[19200];
assign t[19201] = t[19200] ^ n[19201];
assign t[19202] = t[19201] ^ n[19202];
assign t[19203] = t[19202] ^ n[19203];
assign t[19204] = t[19203] ^ n[19204];
assign t[19205] = t[19204] ^ n[19205];
assign t[19206] = t[19205] ^ n[19206];
assign t[19207] = t[19206] ^ n[19207];
assign t[19208] = t[19207] ^ n[19208];
assign t[19209] = t[19208] ^ n[19209];
assign t[19210] = t[19209] ^ n[19210];
assign t[19211] = t[19210] ^ n[19211];
assign t[19212] = t[19211] ^ n[19212];
assign t[19213] = t[19212] ^ n[19213];
assign t[19214] = t[19213] ^ n[19214];
assign t[19215] = t[19214] ^ n[19215];
assign t[19216] = t[19215] ^ n[19216];
assign t[19217] = t[19216] ^ n[19217];
assign t[19218] = t[19217] ^ n[19218];
assign t[19219] = t[19218] ^ n[19219];
assign t[19220] = t[19219] ^ n[19220];
assign t[19221] = t[19220] ^ n[19221];
assign t[19222] = t[19221] ^ n[19222];
assign t[19223] = t[19222] ^ n[19223];
assign t[19224] = t[19223] ^ n[19224];
assign t[19225] = t[19224] ^ n[19225];
assign t[19226] = t[19225] ^ n[19226];
assign t[19227] = t[19226] ^ n[19227];
assign t[19228] = t[19227] ^ n[19228];
assign t[19229] = t[19228] ^ n[19229];
assign t[19230] = t[19229] ^ n[19230];
assign t[19231] = t[19230] ^ n[19231];
assign t[19232] = t[19231] ^ n[19232];
assign t[19233] = t[19232] ^ n[19233];
assign t[19234] = t[19233] ^ n[19234];
assign t[19235] = t[19234] ^ n[19235];
assign t[19236] = t[19235] ^ n[19236];
assign t[19237] = t[19236] ^ n[19237];
assign t[19238] = t[19237] ^ n[19238];
assign t[19239] = t[19238] ^ n[19239];
assign t[19240] = t[19239] ^ n[19240];
assign t[19241] = t[19240] ^ n[19241];
assign t[19242] = t[19241] ^ n[19242];
assign t[19243] = t[19242] ^ n[19243];
assign t[19244] = t[19243] ^ n[19244];
assign t[19245] = t[19244] ^ n[19245];
assign t[19246] = t[19245] ^ n[19246];
assign t[19247] = t[19246] ^ n[19247];
assign t[19248] = t[19247] ^ n[19248];
assign t[19249] = t[19248] ^ n[19249];
assign t[19250] = t[19249] ^ n[19250];
assign t[19251] = t[19250] ^ n[19251];
assign t[19252] = t[19251] ^ n[19252];
assign t[19253] = t[19252] ^ n[19253];
assign t[19254] = t[19253] ^ n[19254];
assign t[19255] = t[19254] ^ n[19255];
assign t[19256] = t[19255] ^ n[19256];
assign t[19257] = t[19256] ^ n[19257];
assign t[19258] = t[19257] ^ n[19258];
assign t[19259] = t[19258] ^ n[19259];
assign t[19260] = t[19259] ^ n[19260];
assign t[19261] = t[19260] ^ n[19261];
assign t[19262] = t[19261] ^ n[19262];
assign t[19263] = t[19262] ^ n[19263];
assign t[19264] = t[19263] ^ n[19264];
assign t[19265] = t[19264] ^ n[19265];
assign t[19266] = t[19265] ^ n[19266];
assign t[19267] = t[19266] ^ n[19267];
assign t[19268] = t[19267] ^ n[19268];
assign t[19269] = t[19268] ^ n[19269];
assign t[19270] = t[19269] ^ n[19270];
assign t[19271] = t[19270] ^ n[19271];
assign t[19272] = t[19271] ^ n[19272];
assign t[19273] = t[19272] ^ n[19273];
assign t[19274] = t[19273] ^ n[19274];
assign t[19275] = t[19274] ^ n[19275];
assign t[19276] = t[19275] ^ n[19276];
assign t[19277] = t[19276] ^ n[19277];
assign t[19278] = t[19277] ^ n[19278];
assign t[19279] = t[19278] ^ n[19279];
assign t[19280] = t[19279] ^ n[19280];
assign t[19281] = t[19280] ^ n[19281];
assign t[19282] = t[19281] ^ n[19282];
assign t[19283] = t[19282] ^ n[19283];
assign t[19284] = t[19283] ^ n[19284];
assign t[19285] = t[19284] ^ n[19285];
assign t[19286] = t[19285] ^ n[19286];
assign t[19287] = t[19286] ^ n[19287];
assign t[19288] = t[19287] ^ n[19288];
assign t[19289] = t[19288] ^ n[19289];
assign t[19290] = t[19289] ^ n[19290];
assign t[19291] = t[19290] ^ n[19291];
assign t[19292] = t[19291] ^ n[19292];
assign t[19293] = t[19292] ^ n[19293];
assign t[19294] = t[19293] ^ n[19294];
assign t[19295] = t[19294] ^ n[19295];
assign t[19296] = t[19295] ^ n[19296];
assign t[19297] = t[19296] ^ n[19297];
assign t[19298] = t[19297] ^ n[19298];
assign t[19299] = t[19298] ^ n[19299];
assign t[19300] = t[19299] ^ n[19300];
assign t[19301] = t[19300] ^ n[19301];
assign t[19302] = t[19301] ^ n[19302];
assign t[19303] = t[19302] ^ n[19303];
assign t[19304] = t[19303] ^ n[19304];
assign t[19305] = t[19304] ^ n[19305];
assign t[19306] = t[19305] ^ n[19306];
assign t[19307] = t[19306] ^ n[19307];
assign t[19308] = t[19307] ^ n[19308];
assign t[19309] = t[19308] ^ n[19309];
assign t[19310] = t[19309] ^ n[19310];
assign t[19311] = t[19310] ^ n[19311];
assign t[19312] = t[19311] ^ n[19312];
assign t[19313] = t[19312] ^ n[19313];
assign t[19314] = t[19313] ^ n[19314];
assign t[19315] = t[19314] ^ n[19315];
assign t[19316] = t[19315] ^ n[19316];
assign t[19317] = t[19316] ^ n[19317];
assign t[19318] = t[19317] ^ n[19318];
assign t[19319] = t[19318] ^ n[19319];
assign t[19320] = t[19319] ^ n[19320];
assign t[19321] = t[19320] ^ n[19321];
assign t[19322] = t[19321] ^ n[19322];
assign t[19323] = t[19322] ^ n[19323];
assign t[19324] = t[19323] ^ n[19324];
assign t[19325] = t[19324] ^ n[19325];
assign t[19326] = t[19325] ^ n[19326];
assign t[19327] = t[19326] ^ n[19327];
assign t[19328] = t[19327] ^ n[19328];
assign t[19329] = t[19328] ^ n[19329];
assign t[19330] = t[19329] ^ n[19330];
assign t[19331] = t[19330] ^ n[19331];
assign t[19332] = t[19331] ^ n[19332];
assign t[19333] = t[19332] ^ n[19333];
assign t[19334] = t[19333] ^ n[19334];
assign t[19335] = t[19334] ^ n[19335];
assign t[19336] = t[19335] ^ n[19336];
assign t[19337] = t[19336] ^ n[19337];
assign t[19338] = t[19337] ^ n[19338];
assign t[19339] = t[19338] ^ n[19339];
assign t[19340] = t[19339] ^ n[19340];
assign t[19341] = t[19340] ^ n[19341];
assign t[19342] = t[19341] ^ n[19342];
assign t[19343] = t[19342] ^ n[19343];
assign t[19344] = t[19343] ^ n[19344];
assign t[19345] = t[19344] ^ n[19345];
assign t[19346] = t[19345] ^ n[19346];
assign t[19347] = t[19346] ^ n[19347];
assign t[19348] = t[19347] ^ n[19348];
assign t[19349] = t[19348] ^ n[19349];
assign t[19350] = t[19349] ^ n[19350];
assign t[19351] = t[19350] ^ n[19351];
assign t[19352] = t[19351] ^ n[19352];
assign t[19353] = t[19352] ^ n[19353];
assign t[19354] = t[19353] ^ n[19354];
assign t[19355] = t[19354] ^ n[19355];
assign t[19356] = t[19355] ^ n[19356];
assign t[19357] = t[19356] ^ n[19357];
assign t[19358] = t[19357] ^ n[19358];
assign t[19359] = t[19358] ^ n[19359];
assign t[19360] = t[19359] ^ n[19360];
assign t[19361] = t[19360] ^ n[19361];
assign t[19362] = t[19361] ^ n[19362];
assign t[19363] = t[19362] ^ n[19363];
assign t[19364] = t[19363] ^ n[19364];
assign t[19365] = t[19364] ^ n[19365];
assign t[19366] = t[19365] ^ n[19366];
assign t[19367] = t[19366] ^ n[19367];
assign t[19368] = t[19367] ^ n[19368];
assign t[19369] = t[19368] ^ n[19369];
assign t[19370] = t[19369] ^ n[19370];
assign t[19371] = t[19370] ^ n[19371];
assign t[19372] = t[19371] ^ n[19372];
assign t[19373] = t[19372] ^ n[19373];
assign t[19374] = t[19373] ^ n[19374];
assign t[19375] = t[19374] ^ n[19375];
assign t[19376] = t[19375] ^ n[19376];
assign t[19377] = t[19376] ^ n[19377];
assign t[19378] = t[19377] ^ n[19378];
assign t[19379] = t[19378] ^ n[19379];
assign t[19380] = t[19379] ^ n[19380];
assign t[19381] = t[19380] ^ n[19381];
assign t[19382] = t[19381] ^ n[19382];
assign t[19383] = t[19382] ^ n[19383];
assign t[19384] = t[19383] ^ n[19384];
assign t[19385] = t[19384] ^ n[19385];
assign t[19386] = t[19385] ^ n[19386];
assign t[19387] = t[19386] ^ n[19387];
assign t[19388] = t[19387] ^ n[19388];
assign t[19389] = t[19388] ^ n[19389];
assign t[19390] = t[19389] ^ n[19390];
assign t[19391] = t[19390] ^ n[19391];
assign t[19392] = t[19391] ^ n[19392];
assign t[19393] = t[19392] ^ n[19393];
assign t[19394] = t[19393] ^ n[19394];
assign t[19395] = t[19394] ^ n[19395];
assign t[19396] = t[19395] ^ n[19396];
assign t[19397] = t[19396] ^ n[19397];
assign t[19398] = t[19397] ^ n[19398];
assign t[19399] = t[19398] ^ n[19399];
assign t[19400] = t[19399] ^ n[19400];
assign t[19401] = t[19400] ^ n[19401];
assign t[19402] = t[19401] ^ n[19402];
assign t[19403] = t[19402] ^ n[19403];
assign t[19404] = t[19403] ^ n[19404];
assign t[19405] = t[19404] ^ n[19405];
assign t[19406] = t[19405] ^ n[19406];
assign t[19407] = t[19406] ^ n[19407];
assign t[19408] = t[19407] ^ n[19408];
assign t[19409] = t[19408] ^ n[19409];
assign t[19410] = t[19409] ^ n[19410];
assign t[19411] = t[19410] ^ n[19411];
assign t[19412] = t[19411] ^ n[19412];
assign t[19413] = t[19412] ^ n[19413];
assign t[19414] = t[19413] ^ n[19414];
assign t[19415] = t[19414] ^ n[19415];
assign t[19416] = t[19415] ^ n[19416];
assign t[19417] = t[19416] ^ n[19417];
assign t[19418] = t[19417] ^ n[19418];
assign t[19419] = t[19418] ^ n[19419];
assign t[19420] = t[19419] ^ n[19420];
assign t[19421] = t[19420] ^ n[19421];
assign t[19422] = t[19421] ^ n[19422];
assign t[19423] = t[19422] ^ n[19423];
assign t[19424] = t[19423] ^ n[19424];
assign t[19425] = t[19424] ^ n[19425];
assign t[19426] = t[19425] ^ n[19426];
assign t[19427] = t[19426] ^ n[19427];
assign t[19428] = t[19427] ^ n[19428];
assign t[19429] = t[19428] ^ n[19429];
assign t[19430] = t[19429] ^ n[19430];
assign t[19431] = t[19430] ^ n[19431];
assign t[19432] = t[19431] ^ n[19432];
assign t[19433] = t[19432] ^ n[19433];
assign t[19434] = t[19433] ^ n[19434];
assign t[19435] = t[19434] ^ n[19435];
assign t[19436] = t[19435] ^ n[19436];
assign t[19437] = t[19436] ^ n[19437];
assign t[19438] = t[19437] ^ n[19438];
assign t[19439] = t[19438] ^ n[19439];
assign t[19440] = t[19439] ^ n[19440];
assign t[19441] = t[19440] ^ n[19441];
assign t[19442] = t[19441] ^ n[19442];
assign t[19443] = t[19442] ^ n[19443];
assign t[19444] = t[19443] ^ n[19444];
assign t[19445] = t[19444] ^ n[19445];
assign t[19446] = t[19445] ^ n[19446];
assign t[19447] = t[19446] ^ n[19447];
assign t[19448] = t[19447] ^ n[19448];
assign t[19449] = t[19448] ^ n[19449];
assign t[19450] = t[19449] ^ n[19450];
assign t[19451] = t[19450] ^ n[19451];
assign t[19452] = t[19451] ^ n[19452];
assign t[19453] = t[19452] ^ n[19453];
assign t[19454] = t[19453] ^ n[19454];
assign t[19455] = t[19454] ^ n[19455];
assign t[19456] = t[19455] ^ n[19456];
assign t[19457] = t[19456] ^ n[19457];
assign t[19458] = t[19457] ^ n[19458];
assign t[19459] = t[19458] ^ n[19459];
assign t[19460] = t[19459] ^ n[19460];
assign t[19461] = t[19460] ^ n[19461];
assign t[19462] = t[19461] ^ n[19462];
assign t[19463] = t[19462] ^ n[19463];
assign t[19464] = t[19463] ^ n[19464];
assign t[19465] = t[19464] ^ n[19465];
assign t[19466] = t[19465] ^ n[19466];
assign t[19467] = t[19466] ^ n[19467];
assign t[19468] = t[19467] ^ n[19468];
assign t[19469] = t[19468] ^ n[19469];
assign t[19470] = t[19469] ^ n[19470];
assign t[19471] = t[19470] ^ n[19471];
assign t[19472] = t[19471] ^ n[19472];
assign t[19473] = t[19472] ^ n[19473];
assign t[19474] = t[19473] ^ n[19474];
assign t[19475] = t[19474] ^ n[19475];
assign t[19476] = t[19475] ^ n[19476];
assign t[19477] = t[19476] ^ n[19477];
assign t[19478] = t[19477] ^ n[19478];
assign t[19479] = t[19478] ^ n[19479];
assign t[19480] = t[19479] ^ n[19480];
assign t[19481] = t[19480] ^ n[19481];
assign t[19482] = t[19481] ^ n[19482];
assign t[19483] = t[19482] ^ n[19483];
assign t[19484] = t[19483] ^ n[19484];
assign t[19485] = t[19484] ^ n[19485];
assign t[19486] = t[19485] ^ n[19486];
assign t[19487] = t[19486] ^ n[19487];
assign t[19488] = t[19487] ^ n[19488];
assign t[19489] = t[19488] ^ n[19489];
assign t[19490] = t[19489] ^ n[19490];
assign t[19491] = t[19490] ^ n[19491];
assign t[19492] = t[19491] ^ n[19492];
assign t[19493] = t[19492] ^ n[19493];
assign t[19494] = t[19493] ^ n[19494];
assign t[19495] = t[19494] ^ n[19495];
assign t[19496] = t[19495] ^ n[19496];
assign t[19497] = t[19496] ^ n[19497];
assign t[19498] = t[19497] ^ n[19498];
assign t[19499] = t[19498] ^ n[19499];
assign t[19500] = t[19499] ^ n[19500];
assign t[19501] = t[19500] ^ n[19501];
assign t[19502] = t[19501] ^ n[19502];
assign t[19503] = t[19502] ^ n[19503];
assign t[19504] = t[19503] ^ n[19504];
assign t[19505] = t[19504] ^ n[19505];
assign t[19506] = t[19505] ^ n[19506];
assign t[19507] = t[19506] ^ n[19507];
assign t[19508] = t[19507] ^ n[19508];
assign t[19509] = t[19508] ^ n[19509];
assign t[19510] = t[19509] ^ n[19510];
assign t[19511] = t[19510] ^ n[19511];
assign t[19512] = t[19511] ^ n[19512];
assign t[19513] = t[19512] ^ n[19513];
assign t[19514] = t[19513] ^ n[19514];
assign t[19515] = t[19514] ^ n[19515];
assign t[19516] = t[19515] ^ n[19516];
assign t[19517] = t[19516] ^ n[19517];
assign t[19518] = t[19517] ^ n[19518];
assign t[19519] = t[19518] ^ n[19519];
assign t[19520] = t[19519] ^ n[19520];
assign t[19521] = t[19520] ^ n[19521];
assign t[19522] = t[19521] ^ n[19522];
assign t[19523] = t[19522] ^ n[19523];
assign t[19524] = t[19523] ^ n[19524];
assign t[19525] = t[19524] ^ n[19525];
assign t[19526] = t[19525] ^ n[19526];
assign t[19527] = t[19526] ^ n[19527];
assign t[19528] = t[19527] ^ n[19528];
assign t[19529] = t[19528] ^ n[19529];
assign t[19530] = t[19529] ^ n[19530];
assign t[19531] = t[19530] ^ n[19531];
assign t[19532] = t[19531] ^ n[19532];
assign t[19533] = t[19532] ^ n[19533];
assign t[19534] = t[19533] ^ n[19534];
assign t[19535] = t[19534] ^ n[19535];
assign t[19536] = t[19535] ^ n[19536];
assign t[19537] = t[19536] ^ n[19537];
assign t[19538] = t[19537] ^ n[19538];
assign t[19539] = t[19538] ^ n[19539];
assign t[19540] = t[19539] ^ n[19540];
assign t[19541] = t[19540] ^ n[19541];
assign t[19542] = t[19541] ^ n[19542];
assign t[19543] = t[19542] ^ n[19543];
assign t[19544] = t[19543] ^ n[19544];
assign t[19545] = t[19544] ^ n[19545];
assign t[19546] = t[19545] ^ n[19546];
assign t[19547] = t[19546] ^ n[19547];
assign t[19548] = t[19547] ^ n[19548];
assign t[19549] = t[19548] ^ n[19549];
assign t[19550] = t[19549] ^ n[19550];
assign t[19551] = t[19550] ^ n[19551];
assign t[19552] = t[19551] ^ n[19552];
assign t[19553] = t[19552] ^ n[19553];
assign t[19554] = t[19553] ^ n[19554];
assign t[19555] = t[19554] ^ n[19555];
assign t[19556] = t[19555] ^ n[19556];
assign t[19557] = t[19556] ^ n[19557];
assign t[19558] = t[19557] ^ n[19558];
assign t[19559] = t[19558] ^ n[19559];
assign t[19560] = t[19559] ^ n[19560];
assign t[19561] = t[19560] ^ n[19561];
assign t[19562] = t[19561] ^ n[19562];
assign t[19563] = t[19562] ^ n[19563];
assign t[19564] = t[19563] ^ n[19564];
assign t[19565] = t[19564] ^ n[19565];
assign t[19566] = t[19565] ^ n[19566];
assign t[19567] = t[19566] ^ n[19567];
assign t[19568] = t[19567] ^ n[19568];
assign t[19569] = t[19568] ^ n[19569];
assign t[19570] = t[19569] ^ n[19570];
assign t[19571] = t[19570] ^ n[19571];
assign t[19572] = t[19571] ^ n[19572];
assign t[19573] = t[19572] ^ n[19573];
assign t[19574] = t[19573] ^ n[19574];
assign t[19575] = t[19574] ^ n[19575];
assign t[19576] = t[19575] ^ n[19576];
assign t[19577] = t[19576] ^ n[19577];
assign t[19578] = t[19577] ^ n[19578];
assign t[19579] = t[19578] ^ n[19579];
assign t[19580] = t[19579] ^ n[19580];
assign t[19581] = t[19580] ^ n[19581];
assign t[19582] = t[19581] ^ n[19582];
assign t[19583] = t[19582] ^ n[19583];
assign t[19584] = t[19583] ^ n[19584];
assign t[19585] = t[19584] ^ n[19585];
assign t[19586] = t[19585] ^ n[19586];
assign t[19587] = t[19586] ^ n[19587];
assign t[19588] = t[19587] ^ n[19588];
assign t[19589] = t[19588] ^ n[19589];
assign t[19590] = t[19589] ^ n[19590];
assign t[19591] = t[19590] ^ n[19591];
assign t[19592] = t[19591] ^ n[19592];
assign t[19593] = t[19592] ^ n[19593];
assign t[19594] = t[19593] ^ n[19594];
assign t[19595] = t[19594] ^ n[19595];
assign t[19596] = t[19595] ^ n[19596];
assign t[19597] = t[19596] ^ n[19597];
assign t[19598] = t[19597] ^ n[19598];
assign t[19599] = t[19598] ^ n[19599];
assign t[19600] = t[19599] ^ n[19600];
assign t[19601] = t[19600] ^ n[19601];
assign t[19602] = t[19601] ^ n[19602];
assign t[19603] = t[19602] ^ n[19603];
assign t[19604] = t[19603] ^ n[19604];
assign t[19605] = t[19604] ^ n[19605];
assign t[19606] = t[19605] ^ n[19606];
assign t[19607] = t[19606] ^ n[19607];
assign t[19608] = t[19607] ^ n[19608];
assign t[19609] = t[19608] ^ n[19609];
assign t[19610] = t[19609] ^ n[19610];
assign t[19611] = t[19610] ^ n[19611];
assign t[19612] = t[19611] ^ n[19612];
assign t[19613] = t[19612] ^ n[19613];
assign t[19614] = t[19613] ^ n[19614];
assign t[19615] = t[19614] ^ n[19615];
assign t[19616] = t[19615] ^ n[19616];
assign t[19617] = t[19616] ^ n[19617];
assign t[19618] = t[19617] ^ n[19618];
assign t[19619] = t[19618] ^ n[19619];
assign t[19620] = t[19619] ^ n[19620];
assign t[19621] = t[19620] ^ n[19621];
assign t[19622] = t[19621] ^ n[19622];
assign t[19623] = t[19622] ^ n[19623];
assign t[19624] = t[19623] ^ n[19624];
assign t[19625] = t[19624] ^ n[19625];
assign t[19626] = t[19625] ^ n[19626];
assign t[19627] = t[19626] ^ n[19627];
assign t[19628] = t[19627] ^ n[19628];
assign t[19629] = t[19628] ^ n[19629];
assign t[19630] = t[19629] ^ n[19630];
assign t[19631] = t[19630] ^ n[19631];
assign t[19632] = t[19631] ^ n[19632];
assign t[19633] = t[19632] ^ n[19633];
assign t[19634] = t[19633] ^ n[19634];
assign t[19635] = t[19634] ^ n[19635];
assign t[19636] = t[19635] ^ n[19636];
assign t[19637] = t[19636] ^ n[19637];
assign t[19638] = t[19637] ^ n[19638];
assign t[19639] = t[19638] ^ n[19639];
assign t[19640] = t[19639] ^ n[19640];
assign t[19641] = t[19640] ^ n[19641];
assign t[19642] = t[19641] ^ n[19642];
assign t[19643] = t[19642] ^ n[19643];
assign t[19644] = t[19643] ^ n[19644];
assign t[19645] = t[19644] ^ n[19645];
assign t[19646] = t[19645] ^ n[19646];
assign t[19647] = t[19646] ^ n[19647];
assign t[19648] = t[19647] ^ n[19648];
assign t[19649] = t[19648] ^ n[19649];
assign t[19650] = t[19649] ^ n[19650];
assign t[19651] = t[19650] ^ n[19651];
assign t[19652] = t[19651] ^ n[19652];
assign t[19653] = t[19652] ^ n[19653];
assign t[19654] = t[19653] ^ n[19654];
assign t[19655] = t[19654] ^ n[19655];
assign t[19656] = t[19655] ^ n[19656];
assign t[19657] = t[19656] ^ n[19657];
assign t[19658] = t[19657] ^ n[19658];
assign t[19659] = t[19658] ^ n[19659];
assign t[19660] = t[19659] ^ n[19660];
assign t[19661] = t[19660] ^ n[19661];
assign t[19662] = t[19661] ^ n[19662];
assign t[19663] = t[19662] ^ n[19663];
assign t[19664] = t[19663] ^ n[19664];
assign t[19665] = t[19664] ^ n[19665];
assign t[19666] = t[19665] ^ n[19666];
assign t[19667] = t[19666] ^ n[19667];
assign t[19668] = t[19667] ^ n[19668];
assign t[19669] = t[19668] ^ n[19669];
assign t[19670] = t[19669] ^ n[19670];
assign t[19671] = t[19670] ^ n[19671];
assign t[19672] = t[19671] ^ n[19672];
assign t[19673] = t[19672] ^ n[19673];
assign t[19674] = t[19673] ^ n[19674];
assign t[19675] = t[19674] ^ n[19675];
assign t[19676] = t[19675] ^ n[19676];
assign t[19677] = t[19676] ^ n[19677];
assign t[19678] = t[19677] ^ n[19678];
assign t[19679] = t[19678] ^ n[19679];
assign t[19680] = t[19679] ^ n[19680];
assign t[19681] = t[19680] ^ n[19681];
assign t[19682] = t[19681] ^ n[19682];
assign t[19683] = t[19682] ^ n[19683];
assign t[19684] = t[19683] ^ n[19684];
assign t[19685] = t[19684] ^ n[19685];
assign t[19686] = t[19685] ^ n[19686];
assign t[19687] = t[19686] ^ n[19687];
assign t[19688] = t[19687] ^ n[19688];
assign t[19689] = t[19688] ^ n[19689];
assign t[19690] = t[19689] ^ n[19690];
assign t[19691] = t[19690] ^ n[19691];
assign t[19692] = t[19691] ^ n[19692];
assign t[19693] = t[19692] ^ n[19693];
assign t[19694] = t[19693] ^ n[19694];
assign t[19695] = t[19694] ^ n[19695];
assign t[19696] = t[19695] ^ n[19696];
assign t[19697] = t[19696] ^ n[19697];
assign t[19698] = t[19697] ^ n[19698];
assign t[19699] = t[19698] ^ n[19699];
assign t[19700] = t[19699] ^ n[19700];
assign t[19701] = t[19700] ^ n[19701];
assign t[19702] = t[19701] ^ n[19702];
assign t[19703] = t[19702] ^ n[19703];
assign t[19704] = t[19703] ^ n[19704];
assign t[19705] = t[19704] ^ n[19705];
assign t[19706] = t[19705] ^ n[19706];
assign t[19707] = t[19706] ^ n[19707];
assign t[19708] = t[19707] ^ n[19708];
assign t[19709] = t[19708] ^ n[19709];
assign t[19710] = t[19709] ^ n[19710];
assign t[19711] = t[19710] ^ n[19711];
assign t[19712] = t[19711] ^ n[19712];
assign t[19713] = t[19712] ^ n[19713];
assign t[19714] = t[19713] ^ n[19714];
assign t[19715] = t[19714] ^ n[19715];
assign t[19716] = t[19715] ^ n[19716];
assign t[19717] = t[19716] ^ n[19717];
assign t[19718] = t[19717] ^ n[19718];
assign t[19719] = t[19718] ^ n[19719];
assign t[19720] = t[19719] ^ n[19720];
assign t[19721] = t[19720] ^ n[19721];
assign t[19722] = t[19721] ^ n[19722];
assign t[19723] = t[19722] ^ n[19723];
assign t[19724] = t[19723] ^ n[19724];
assign t[19725] = t[19724] ^ n[19725];
assign t[19726] = t[19725] ^ n[19726];
assign t[19727] = t[19726] ^ n[19727];
assign t[19728] = t[19727] ^ n[19728];
assign t[19729] = t[19728] ^ n[19729];
assign t[19730] = t[19729] ^ n[19730];
assign t[19731] = t[19730] ^ n[19731];
assign t[19732] = t[19731] ^ n[19732];
assign t[19733] = t[19732] ^ n[19733];
assign t[19734] = t[19733] ^ n[19734];
assign t[19735] = t[19734] ^ n[19735];
assign t[19736] = t[19735] ^ n[19736];
assign t[19737] = t[19736] ^ n[19737];
assign t[19738] = t[19737] ^ n[19738];
assign t[19739] = t[19738] ^ n[19739];
assign t[19740] = t[19739] ^ n[19740];
assign t[19741] = t[19740] ^ n[19741];
assign t[19742] = t[19741] ^ n[19742];
assign t[19743] = t[19742] ^ n[19743];
assign t[19744] = t[19743] ^ n[19744];
assign t[19745] = t[19744] ^ n[19745];
assign t[19746] = t[19745] ^ n[19746];
assign t[19747] = t[19746] ^ n[19747];
assign t[19748] = t[19747] ^ n[19748];
assign t[19749] = t[19748] ^ n[19749];
assign t[19750] = t[19749] ^ n[19750];
assign t[19751] = t[19750] ^ n[19751];
assign t[19752] = t[19751] ^ n[19752];
assign t[19753] = t[19752] ^ n[19753];
assign t[19754] = t[19753] ^ n[19754];
assign t[19755] = t[19754] ^ n[19755];
assign t[19756] = t[19755] ^ n[19756];
assign t[19757] = t[19756] ^ n[19757];
assign t[19758] = t[19757] ^ n[19758];
assign t[19759] = t[19758] ^ n[19759];
assign t[19760] = t[19759] ^ n[19760];
assign t[19761] = t[19760] ^ n[19761];
assign t[19762] = t[19761] ^ n[19762];
assign t[19763] = t[19762] ^ n[19763];
assign t[19764] = t[19763] ^ n[19764];
assign t[19765] = t[19764] ^ n[19765];
assign t[19766] = t[19765] ^ n[19766];
assign t[19767] = t[19766] ^ n[19767];
assign t[19768] = t[19767] ^ n[19768];
assign t[19769] = t[19768] ^ n[19769];
assign t[19770] = t[19769] ^ n[19770];
assign t[19771] = t[19770] ^ n[19771];
assign t[19772] = t[19771] ^ n[19772];
assign t[19773] = t[19772] ^ n[19773];
assign t[19774] = t[19773] ^ n[19774];
assign t[19775] = t[19774] ^ n[19775];
assign t[19776] = t[19775] ^ n[19776];
assign t[19777] = t[19776] ^ n[19777];
assign t[19778] = t[19777] ^ n[19778];
assign t[19779] = t[19778] ^ n[19779];
assign t[19780] = t[19779] ^ n[19780];
assign t[19781] = t[19780] ^ n[19781];
assign t[19782] = t[19781] ^ n[19782];
assign t[19783] = t[19782] ^ n[19783];
assign t[19784] = t[19783] ^ n[19784];
assign t[19785] = t[19784] ^ n[19785];
assign t[19786] = t[19785] ^ n[19786];
assign t[19787] = t[19786] ^ n[19787];
assign t[19788] = t[19787] ^ n[19788];
assign t[19789] = t[19788] ^ n[19789];
assign t[19790] = t[19789] ^ n[19790];
assign t[19791] = t[19790] ^ n[19791];
assign t[19792] = t[19791] ^ n[19792];
assign t[19793] = t[19792] ^ n[19793];
assign t[19794] = t[19793] ^ n[19794];
assign t[19795] = t[19794] ^ n[19795];
assign t[19796] = t[19795] ^ n[19796];
assign t[19797] = t[19796] ^ n[19797];
assign t[19798] = t[19797] ^ n[19798];
assign t[19799] = t[19798] ^ n[19799];
assign t[19800] = t[19799] ^ n[19800];
assign t[19801] = t[19800] ^ n[19801];
assign t[19802] = t[19801] ^ n[19802];
assign t[19803] = t[19802] ^ n[19803];
assign t[19804] = t[19803] ^ n[19804];
assign t[19805] = t[19804] ^ n[19805];
assign t[19806] = t[19805] ^ n[19806];
assign t[19807] = t[19806] ^ n[19807];
assign t[19808] = t[19807] ^ n[19808];
assign t[19809] = t[19808] ^ n[19809];
assign t[19810] = t[19809] ^ n[19810];
assign t[19811] = t[19810] ^ n[19811];
assign t[19812] = t[19811] ^ n[19812];
assign t[19813] = t[19812] ^ n[19813];
assign t[19814] = t[19813] ^ n[19814];
assign t[19815] = t[19814] ^ n[19815];
assign t[19816] = t[19815] ^ n[19816];
assign t[19817] = t[19816] ^ n[19817];
assign t[19818] = t[19817] ^ n[19818];
assign t[19819] = t[19818] ^ n[19819];
assign t[19820] = t[19819] ^ n[19820];
assign t[19821] = t[19820] ^ n[19821];
assign t[19822] = t[19821] ^ n[19822];
assign t[19823] = t[19822] ^ n[19823];
assign t[19824] = t[19823] ^ n[19824];
assign t[19825] = t[19824] ^ n[19825];
assign t[19826] = t[19825] ^ n[19826];
assign t[19827] = t[19826] ^ n[19827];
assign t[19828] = t[19827] ^ n[19828];
assign t[19829] = t[19828] ^ n[19829];
assign t[19830] = t[19829] ^ n[19830];
assign t[19831] = t[19830] ^ n[19831];
assign t[19832] = t[19831] ^ n[19832];
assign t[19833] = t[19832] ^ n[19833];
assign t[19834] = t[19833] ^ n[19834];
assign t[19835] = t[19834] ^ n[19835];
assign t[19836] = t[19835] ^ n[19836];
assign t[19837] = t[19836] ^ n[19837];
assign t[19838] = t[19837] ^ n[19838];
assign t[19839] = t[19838] ^ n[19839];
assign t[19840] = t[19839] ^ n[19840];
assign t[19841] = t[19840] ^ n[19841];
assign t[19842] = t[19841] ^ n[19842];
assign t[19843] = t[19842] ^ n[19843];
assign t[19844] = t[19843] ^ n[19844];
assign t[19845] = t[19844] ^ n[19845];
assign t[19846] = t[19845] ^ n[19846];
assign t[19847] = t[19846] ^ n[19847];
assign t[19848] = t[19847] ^ n[19848];
assign t[19849] = t[19848] ^ n[19849];
assign t[19850] = t[19849] ^ n[19850];
assign t[19851] = t[19850] ^ n[19851];
assign t[19852] = t[19851] ^ n[19852];
assign t[19853] = t[19852] ^ n[19853];
assign t[19854] = t[19853] ^ n[19854];
assign t[19855] = t[19854] ^ n[19855];
assign t[19856] = t[19855] ^ n[19856];
assign t[19857] = t[19856] ^ n[19857];
assign t[19858] = t[19857] ^ n[19858];
assign t[19859] = t[19858] ^ n[19859];
assign t[19860] = t[19859] ^ n[19860];
assign t[19861] = t[19860] ^ n[19861];
assign t[19862] = t[19861] ^ n[19862];
assign t[19863] = t[19862] ^ n[19863];
assign t[19864] = t[19863] ^ n[19864];
assign t[19865] = t[19864] ^ n[19865];
assign t[19866] = t[19865] ^ n[19866];
assign t[19867] = t[19866] ^ n[19867];
assign t[19868] = t[19867] ^ n[19868];
assign t[19869] = t[19868] ^ n[19869];
assign t[19870] = t[19869] ^ n[19870];
assign t[19871] = t[19870] ^ n[19871];
assign t[19872] = t[19871] ^ n[19872];
assign t[19873] = t[19872] ^ n[19873];
assign t[19874] = t[19873] ^ n[19874];
assign t[19875] = t[19874] ^ n[19875];
assign t[19876] = t[19875] ^ n[19876];
assign t[19877] = t[19876] ^ n[19877];
assign t[19878] = t[19877] ^ n[19878];
assign t[19879] = t[19878] ^ n[19879];
assign t[19880] = t[19879] ^ n[19880];
assign t[19881] = t[19880] ^ n[19881];
assign t[19882] = t[19881] ^ n[19882];
assign t[19883] = t[19882] ^ n[19883];
assign t[19884] = t[19883] ^ n[19884];
assign t[19885] = t[19884] ^ n[19885];
assign t[19886] = t[19885] ^ n[19886];
assign t[19887] = t[19886] ^ n[19887];
assign t[19888] = t[19887] ^ n[19888];
assign t[19889] = t[19888] ^ n[19889];
assign t[19890] = t[19889] ^ n[19890];
assign t[19891] = t[19890] ^ n[19891];
assign t[19892] = t[19891] ^ n[19892];
assign t[19893] = t[19892] ^ n[19893];
assign t[19894] = t[19893] ^ n[19894];
assign t[19895] = t[19894] ^ n[19895];
assign t[19896] = t[19895] ^ n[19896];
assign t[19897] = t[19896] ^ n[19897];
assign t[19898] = t[19897] ^ n[19898];
assign t[19899] = t[19898] ^ n[19899];
assign t[19900] = t[19899] ^ n[19900];
assign t[19901] = t[19900] ^ n[19901];
assign t[19902] = t[19901] ^ n[19902];
assign t[19903] = t[19902] ^ n[19903];
assign t[19904] = t[19903] ^ n[19904];
assign t[19905] = t[19904] ^ n[19905];
assign t[19906] = t[19905] ^ n[19906];
assign t[19907] = t[19906] ^ n[19907];
assign t[19908] = t[19907] ^ n[19908];
assign t[19909] = t[19908] ^ n[19909];
assign t[19910] = t[19909] ^ n[19910];
assign t[19911] = t[19910] ^ n[19911];
assign t[19912] = t[19911] ^ n[19912];
assign t[19913] = t[19912] ^ n[19913];
assign t[19914] = t[19913] ^ n[19914];
assign t[19915] = t[19914] ^ n[19915];
assign t[19916] = t[19915] ^ n[19916];
assign t[19917] = t[19916] ^ n[19917];
assign t[19918] = t[19917] ^ n[19918];
assign t[19919] = t[19918] ^ n[19919];
assign t[19920] = t[19919] ^ n[19920];
assign t[19921] = t[19920] ^ n[19921];
assign t[19922] = t[19921] ^ n[19922];
assign t[19923] = t[19922] ^ n[19923];
assign t[19924] = t[19923] ^ n[19924];
assign t[19925] = t[19924] ^ n[19925];
assign t[19926] = t[19925] ^ n[19926];
assign t[19927] = t[19926] ^ n[19927];
assign t[19928] = t[19927] ^ n[19928];
assign t[19929] = t[19928] ^ n[19929];
assign t[19930] = t[19929] ^ n[19930];
assign t[19931] = t[19930] ^ n[19931];
assign t[19932] = t[19931] ^ n[19932];
assign t[19933] = t[19932] ^ n[19933];
assign t[19934] = t[19933] ^ n[19934];
assign t[19935] = t[19934] ^ n[19935];
assign t[19936] = t[19935] ^ n[19936];
assign t[19937] = t[19936] ^ n[19937];
assign t[19938] = t[19937] ^ n[19938];
assign t[19939] = t[19938] ^ n[19939];
assign t[19940] = t[19939] ^ n[19940];
assign t[19941] = t[19940] ^ n[19941];
assign t[19942] = t[19941] ^ n[19942];
assign t[19943] = t[19942] ^ n[19943];
assign t[19944] = t[19943] ^ n[19944];
assign t[19945] = t[19944] ^ n[19945];
assign t[19946] = t[19945] ^ n[19946];
assign t[19947] = t[19946] ^ n[19947];
assign t[19948] = t[19947] ^ n[19948];
assign t[19949] = t[19948] ^ n[19949];
assign t[19950] = t[19949] ^ n[19950];
assign t[19951] = t[19950] ^ n[19951];
assign t[19952] = t[19951] ^ n[19952];
assign t[19953] = t[19952] ^ n[19953];
assign t[19954] = t[19953] ^ n[19954];
assign t[19955] = t[19954] ^ n[19955];
assign t[19956] = t[19955] ^ n[19956];
assign t[19957] = t[19956] ^ n[19957];
assign t[19958] = t[19957] ^ n[19958];
assign t[19959] = t[19958] ^ n[19959];
assign t[19960] = t[19959] ^ n[19960];
assign t[19961] = t[19960] ^ n[19961];
assign t[19962] = t[19961] ^ n[19962];
assign t[19963] = t[19962] ^ n[19963];
assign t[19964] = t[19963] ^ n[19964];
assign t[19965] = t[19964] ^ n[19965];
assign t[19966] = t[19965] ^ n[19966];
assign t[19967] = t[19966] ^ n[19967];
assign t[19968] = t[19967] ^ n[19968];
assign t[19969] = t[19968] ^ n[19969];
assign t[19970] = t[19969] ^ n[19970];
assign t[19971] = t[19970] ^ n[19971];
assign t[19972] = t[19971] ^ n[19972];
assign t[19973] = t[19972] ^ n[19973];
assign t[19974] = t[19973] ^ n[19974];
assign t[19975] = t[19974] ^ n[19975];
assign t[19976] = t[19975] ^ n[19976];
assign t[19977] = t[19976] ^ n[19977];
assign t[19978] = t[19977] ^ n[19978];
assign t[19979] = t[19978] ^ n[19979];
assign t[19980] = t[19979] ^ n[19980];
assign t[19981] = t[19980] ^ n[19981];
assign t[19982] = t[19981] ^ n[19982];
assign t[19983] = t[19982] ^ n[19983];
assign t[19984] = t[19983] ^ n[19984];
assign t[19985] = t[19984] ^ n[19985];
assign t[19986] = t[19985] ^ n[19986];
assign t[19987] = t[19986] ^ n[19987];
assign t[19988] = t[19987] ^ n[19988];
assign t[19989] = t[19988] ^ n[19989];
assign t[19990] = t[19989] ^ n[19990];
assign t[19991] = t[19990] ^ n[19991];
assign t[19992] = t[19991] ^ n[19992];
assign t[19993] = t[19992] ^ n[19993];
assign t[19994] = t[19993] ^ n[19994];
assign t[19995] = t[19994] ^ n[19995];
assign t[19996] = t[19995] ^ n[19996];
assign t[19997] = t[19996] ^ n[19997];
assign t[19998] = t[19997] ^ n[19998];
assign t[19999] = t[19998] ^ n[19999];
assign t[20000] = t[19999] ^ n[20000];
assign t[20001] = t[20000] ^ n[20001];
assign t[20002] = t[20001] ^ n[20002];
assign t[20003] = t[20002] ^ n[20003];
assign t[20004] = t[20003] ^ n[20004];
assign t[20005] = t[20004] ^ n[20005];
assign t[20006] = t[20005] ^ n[20006];
assign t[20007] = t[20006] ^ n[20007];
assign t[20008] = t[20007] ^ n[20008];
assign t[20009] = t[20008] ^ n[20009];
assign t[20010] = t[20009] ^ n[20010];
assign t[20011] = t[20010] ^ n[20011];
assign t[20012] = t[20011] ^ n[20012];
assign t[20013] = t[20012] ^ n[20013];
assign t[20014] = t[20013] ^ n[20014];
assign t[20015] = t[20014] ^ n[20015];
assign t[20016] = t[20015] ^ n[20016];
assign t[20017] = t[20016] ^ n[20017];
assign t[20018] = t[20017] ^ n[20018];
assign t[20019] = t[20018] ^ n[20019];
assign t[20020] = t[20019] ^ n[20020];
assign t[20021] = t[20020] ^ n[20021];
assign t[20022] = t[20021] ^ n[20022];
assign t[20023] = t[20022] ^ n[20023];
assign t[20024] = t[20023] ^ n[20024];
assign t[20025] = t[20024] ^ n[20025];
assign t[20026] = t[20025] ^ n[20026];
assign t[20027] = t[20026] ^ n[20027];
assign t[20028] = t[20027] ^ n[20028];
assign t[20029] = t[20028] ^ n[20029];
assign t[20030] = t[20029] ^ n[20030];
assign t[20031] = t[20030] ^ n[20031];
assign t[20032] = t[20031] ^ n[20032];
assign t[20033] = t[20032] ^ n[20033];
assign t[20034] = t[20033] ^ n[20034];
assign t[20035] = t[20034] ^ n[20035];
assign t[20036] = t[20035] ^ n[20036];
assign t[20037] = t[20036] ^ n[20037];
assign t[20038] = t[20037] ^ n[20038];
assign t[20039] = t[20038] ^ n[20039];
assign t[20040] = t[20039] ^ n[20040];
assign t[20041] = t[20040] ^ n[20041];
assign t[20042] = t[20041] ^ n[20042];
assign t[20043] = t[20042] ^ n[20043];
assign t[20044] = t[20043] ^ n[20044];
assign t[20045] = t[20044] ^ n[20045];
assign t[20046] = t[20045] ^ n[20046];
assign t[20047] = t[20046] ^ n[20047];
assign t[20048] = t[20047] ^ n[20048];
assign t[20049] = t[20048] ^ n[20049];
assign t[20050] = t[20049] ^ n[20050];
assign t[20051] = t[20050] ^ n[20051];
assign t[20052] = t[20051] ^ n[20052];
assign t[20053] = t[20052] ^ n[20053];
assign t[20054] = t[20053] ^ n[20054];
assign t[20055] = t[20054] ^ n[20055];
assign t[20056] = t[20055] ^ n[20056];
assign t[20057] = t[20056] ^ n[20057];
assign t[20058] = t[20057] ^ n[20058];
assign t[20059] = t[20058] ^ n[20059];
assign t[20060] = t[20059] ^ n[20060];
assign t[20061] = t[20060] ^ n[20061];
assign t[20062] = t[20061] ^ n[20062];
assign t[20063] = t[20062] ^ n[20063];
assign t[20064] = t[20063] ^ n[20064];
assign t[20065] = t[20064] ^ n[20065];
assign t[20066] = t[20065] ^ n[20066];
assign t[20067] = t[20066] ^ n[20067];
assign t[20068] = t[20067] ^ n[20068];
assign t[20069] = t[20068] ^ n[20069];
assign t[20070] = t[20069] ^ n[20070];
assign t[20071] = t[20070] ^ n[20071];
assign t[20072] = t[20071] ^ n[20072];
assign t[20073] = t[20072] ^ n[20073];
assign t[20074] = t[20073] ^ n[20074];
assign t[20075] = t[20074] ^ n[20075];
assign t[20076] = t[20075] ^ n[20076];
assign t[20077] = t[20076] ^ n[20077];
assign t[20078] = t[20077] ^ n[20078];
assign t[20079] = t[20078] ^ n[20079];
assign t[20080] = t[20079] ^ n[20080];
assign t[20081] = t[20080] ^ n[20081];
assign t[20082] = t[20081] ^ n[20082];
assign t[20083] = t[20082] ^ n[20083];
assign t[20084] = t[20083] ^ n[20084];
assign t[20085] = t[20084] ^ n[20085];
assign t[20086] = t[20085] ^ n[20086];
assign t[20087] = t[20086] ^ n[20087];
assign t[20088] = t[20087] ^ n[20088];
assign t[20089] = t[20088] ^ n[20089];
assign t[20090] = t[20089] ^ n[20090];
assign t[20091] = t[20090] ^ n[20091];
assign t[20092] = t[20091] ^ n[20092];
assign t[20093] = t[20092] ^ n[20093];
assign t[20094] = t[20093] ^ n[20094];
assign t[20095] = t[20094] ^ n[20095];
assign t[20096] = t[20095] ^ n[20096];
assign t[20097] = t[20096] ^ n[20097];
assign t[20098] = t[20097] ^ n[20098];
assign t[20099] = t[20098] ^ n[20099];
assign t[20100] = t[20099] ^ n[20100];
assign t[20101] = t[20100] ^ n[20101];
assign t[20102] = t[20101] ^ n[20102];
assign t[20103] = t[20102] ^ n[20103];
assign t[20104] = t[20103] ^ n[20104];
assign t[20105] = t[20104] ^ n[20105];
assign t[20106] = t[20105] ^ n[20106];
assign t[20107] = t[20106] ^ n[20107];
assign t[20108] = t[20107] ^ n[20108];
assign t[20109] = t[20108] ^ n[20109];
assign t[20110] = t[20109] ^ n[20110];
assign t[20111] = t[20110] ^ n[20111];
assign t[20112] = t[20111] ^ n[20112];
assign t[20113] = t[20112] ^ n[20113];
assign t[20114] = t[20113] ^ n[20114];
assign t[20115] = t[20114] ^ n[20115];
assign t[20116] = t[20115] ^ n[20116];
assign t[20117] = t[20116] ^ n[20117];
assign t[20118] = t[20117] ^ n[20118];
assign t[20119] = t[20118] ^ n[20119];
assign t[20120] = t[20119] ^ n[20120];
assign t[20121] = t[20120] ^ n[20121];
assign t[20122] = t[20121] ^ n[20122];
assign t[20123] = t[20122] ^ n[20123];
assign t[20124] = t[20123] ^ n[20124];
assign t[20125] = t[20124] ^ n[20125];
assign t[20126] = t[20125] ^ n[20126];
assign t[20127] = t[20126] ^ n[20127];
assign t[20128] = t[20127] ^ n[20128];
assign t[20129] = t[20128] ^ n[20129];
assign t[20130] = t[20129] ^ n[20130];
assign t[20131] = t[20130] ^ n[20131];
assign t[20132] = t[20131] ^ n[20132];
assign t[20133] = t[20132] ^ n[20133];
assign t[20134] = t[20133] ^ n[20134];
assign t[20135] = t[20134] ^ n[20135];
assign t[20136] = t[20135] ^ n[20136];
assign t[20137] = t[20136] ^ n[20137];
assign t[20138] = t[20137] ^ n[20138];
assign t[20139] = t[20138] ^ n[20139];
assign t[20140] = t[20139] ^ n[20140];
assign t[20141] = t[20140] ^ n[20141];
assign t[20142] = t[20141] ^ n[20142];
assign t[20143] = t[20142] ^ n[20143];
assign t[20144] = t[20143] ^ n[20144];
assign t[20145] = t[20144] ^ n[20145];
assign t[20146] = t[20145] ^ n[20146];
assign t[20147] = t[20146] ^ n[20147];
assign t[20148] = t[20147] ^ n[20148];
assign t[20149] = t[20148] ^ n[20149];
assign t[20150] = t[20149] ^ n[20150];
assign t[20151] = t[20150] ^ n[20151];
assign t[20152] = t[20151] ^ n[20152];
assign t[20153] = t[20152] ^ n[20153];
assign t[20154] = t[20153] ^ n[20154];
assign t[20155] = t[20154] ^ n[20155];
assign t[20156] = t[20155] ^ n[20156];
assign t[20157] = t[20156] ^ n[20157];
assign t[20158] = t[20157] ^ n[20158];
assign t[20159] = t[20158] ^ n[20159];
assign t[20160] = t[20159] ^ n[20160];
assign t[20161] = t[20160] ^ n[20161];
assign t[20162] = t[20161] ^ n[20162];
assign t[20163] = t[20162] ^ n[20163];
assign t[20164] = t[20163] ^ n[20164];
assign t[20165] = t[20164] ^ n[20165];
assign t[20166] = t[20165] ^ n[20166];
assign t[20167] = t[20166] ^ n[20167];
assign t[20168] = t[20167] ^ n[20168];
assign t[20169] = t[20168] ^ n[20169];
assign t[20170] = t[20169] ^ n[20170];
assign t[20171] = t[20170] ^ n[20171];
assign t[20172] = t[20171] ^ n[20172];
assign t[20173] = t[20172] ^ n[20173];
assign t[20174] = t[20173] ^ n[20174];
assign t[20175] = t[20174] ^ n[20175];
assign t[20176] = t[20175] ^ n[20176];
assign t[20177] = t[20176] ^ n[20177];
assign t[20178] = t[20177] ^ n[20178];
assign t[20179] = t[20178] ^ n[20179];
assign t[20180] = t[20179] ^ n[20180];
assign t[20181] = t[20180] ^ n[20181];
assign t[20182] = t[20181] ^ n[20182];
assign t[20183] = t[20182] ^ n[20183];
assign t[20184] = t[20183] ^ n[20184];
assign t[20185] = t[20184] ^ n[20185];
assign t[20186] = t[20185] ^ n[20186];
assign t[20187] = t[20186] ^ n[20187];
assign t[20188] = t[20187] ^ n[20188];
assign t[20189] = t[20188] ^ n[20189];
assign t[20190] = t[20189] ^ n[20190];
assign t[20191] = t[20190] ^ n[20191];
assign t[20192] = t[20191] ^ n[20192];
assign t[20193] = t[20192] ^ n[20193];
assign t[20194] = t[20193] ^ n[20194];
assign t[20195] = t[20194] ^ n[20195];
assign t[20196] = t[20195] ^ n[20196];
assign t[20197] = t[20196] ^ n[20197];
assign t[20198] = t[20197] ^ n[20198];
assign t[20199] = t[20198] ^ n[20199];
assign t[20200] = t[20199] ^ n[20200];
assign t[20201] = t[20200] ^ n[20201];
assign t[20202] = t[20201] ^ n[20202];
assign t[20203] = t[20202] ^ n[20203];
assign t[20204] = t[20203] ^ n[20204];
assign t[20205] = t[20204] ^ n[20205];
assign t[20206] = t[20205] ^ n[20206];
assign t[20207] = t[20206] ^ n[20207];
assign t[20208] = t[20207] ^ n[20208];
assign t[20209] = t[20208] ^ n[20209];
assign t[20210] = t[20209] ^ n[20210];
assign t[20211] = t[20210] ^ n[20211];
assign t[20212] = t[20211] ^ n[20212];
assign t[20213] = t[20212] ^ n[20213];
assign t[20214] = t[20213] ^ n[20214];
assign t[20215] = t[20214] ^ n[20215];
assign t[20216] = t[20215] ^ n[20216];
assign t[20217] = t[20216] ^ n[20217];
assign t[20218] = t[20217] ^ n[20218];
assign t[20219] = t[20218] ^ n[20219];
assign t[20220] = t[20219] ^ n[20220];
assign t[20221] = t[20220] ^ n[20221];
assign t[20222] = t[20221] ^ n[20222];
assign t[20223] = t[20222] ^ n[20223];
assign t[20224] = t[20223] ^ n[20224];
assign t[20225] = t[20224] ^ n[20225];
assign t[20226] = t[20225] ^ n[20226];
assign t[20227] = t[20226] ^ n[20227];
assign t[20228] = t[20227] ^ n[20228];
assign t[20229] = t[20228] ^ n[20229];
assign t[20230] = t[20229] ^ n[20230];
assign t[20231] = t[20230] ^ n[20231];
assign t[20232] = t[20231] ^ n[20232];
assign t[20233] = t[20232] ^ n[20233];
assign t[20234] = t[20233] ^ n[20234];
assign t[20235] = t[20234] ^ n[20235];
assign t[20236] = t[20235] ^ n[20236];
assign t[20237] = t[20236] ^ n[20237];
assign t[20238] = t[20237] ^ n[20238];
assign t[20239] = t[20238] ^ n[20239];
assign t[20240] = t[20239] ^ n[20240];
assign t[20241] = t[20240] ^ n[20241];
assign t[20242] = t[20241] ^ n[20242];
assign t[20243] = t[20242] ^ n[20243];
assign t[20244] = t[20243] ^ n[20244];
assign t[20245] = t[20244] ^ n[20245];
assign t[20246] = t[20245] ^ n[20246];
assign t[20247] = t[20246] ^ n[20247];
assign t[20248] = t[20247] ^ n[20248];
assign t[20249] = t[20248] ^ n[20249];
assign t[20250] = t[20249] ^ n[20250];
assign t[20251] = t[20250] ^ n[20251];
assign t[20252] = t[20251] ^ n[20252];
assign t[20253] = t[20252] ^ n[20253];
assign t[20254] = t[20253] ^ n[20254];
assign t[20255] = t[20254] ^ n[20255];
assign t[20256] = t[20255] ^ n[20256];
assign t[20257] = t[20256] ^ n[20257];
assign t[20258] = t[20257] ^ n[20258];
assign t[20259] = t[20258] ^ n[20259];
assign t[20260] = t[20259] ^ n[20260];
assign t[20261] = t[20260] ^ n[20261];
assign t[20262] = t[20261] ^ n[20262];
assign t[20263] = t[20262] ^ n[20263];
assign t[20264] = t[20263] ^ n[20264];
assign t[20265] = t[20264] ^ n[20265];
assign t[20266] = t[20265] ^ n[20266];
assign t[20267] = t[20266] ^ n[20267];
assign t[20268] = t[20267] ^ n[20268];
assign t[20269] = t[20268] ^ n[20269];
assign t[20270] = t[20269] ^ n[20270];
assign t[20271] = t[20270] ^ n[20271];
assign t[20272] = t[20271] ^ n[20272];
assign t[20273] = t[20272] ^ n[20273];
assign t[20274] = t[20273] ^ n[20274];
assign t[20275] = t[20274] ^ n[20275];
assign t[20276] = t[20275] ^ n[20276];
assign t[20277] = t[20276] ^ n[20277];
assign t[20278] = t[20277] ^ n[20278];
assign t[20279] = t[20278] ^ n[20279];
assign t[20280] = t[20279] ^ n[20280];
assign t[20281] = t[20280] ^ n[20281];
assign t[20282] = t[20281] ^ n[20282];
assign t[20283] = t[20282] ^ n[20283];
assign t[20284] = t[20283] ^ n[20284];
assign t[20285] = t[20284] ^ n[20285];
assign t[20286] = t[20285] ^ n[20286];
assign t[20287] = t[20286] ^ n[20287];
assign t[20288] = t[20287] ^ n[20288];
assign t[20289] = t[20288] ^ n[20289];
assign t[20290] = t[20289] ^ n[20290];
assign t[20291] = t[20290] ^ n[20291];
assign t[20292] = t[20291] ^ n[20292];
assign t[20293] = t[20292] ^ n[20293];
assign t[20294] = t[20293] ^ n[20294];
assign t[20295] = t[20294] ^ n[20295];
assign t[20296] = t[20295] ^ n[20296];
assign t[20297] = t[20296] ^ n[20297];
assign t[20298] = t[20297] ^ n[20298];
assign t[20299] = t[20298] ^ n[20299];
assign t[20300] = t[20299] ^ n[20300];
assign t[20301] = t[20300] ^ n[20301];
assign t[20302] = t[20301] ^ n[20302];
assign t[20303] = t[20302] ^ n[20303];
assign t[20304] = t[20303] ^ n[20304];
assign t[20305] = t[20304] ^ n[20305];
assign t[20306] = t[20305] ^ n[20306];
assign t[20307] = t[20306] ^ n[20307];
assign t[20308] = t[20307] ^ n[20308];
assign t[20309] = t[20308] ^ n[20309];
assign t[20310] = t[20309] ^ n[20310];
assign t[20311] = t[20310] ^ n[20311];
assign t[20312] = t[20311] ^ n[20312];
assign t[20313] = t[20312] ^ n[20313];
assign t[20314] = t[20313] ^ n[20314];
assign t[20315] = t[20314] ^ n[20315];
assign t[20316] = t[20315] ^ n[20316];
assign t[20317] = t[20316] ^ n[20317];
assign t[20318] = t[20317] ^ n[20318];
assign t[20319] = t[20318] ^ n[20319];
assign t[20320] = t[20319] ^ n[20320];
assign t[20321] = t[20320] ^ n[20321];
assign t[20322] = t[20321] ^ n[20322];
assign t[20323] = t[20322] ^ n[20323];
assign t[20324] = t[20323] ^ n[20324];
assign t[20325] = t[20324] ^ n[20325];
assign t[20326] = t[20325] ^ n[20326];
assign t[20327] = t[20326] ^ n[20327];
assign t[20328] = t[20327] ^ n[20328];
assign t[20329] = t[20328] ^ n[20329];
assign t[20330] = t[20329] ^ n[20330];
assign t[20331] = t[20330] ^ n[20331];
assign t[20332] = t[20331] ^ n[20332];
assign t[20333] = t[20332] ^ n[20333];
assign t[20334] = t[20333] ^ n[20334];
assign t[20335] = t[20334] ^ n[20335];
assign t[20336] = t[20335] ^ n[20336];
assign t[20337] = t[20336] ^ n[20337];
assign t[20338] = t[20337] ^ n[20338];
assign t[20339] = t[20338] ^ n[20339];
assign t[20340] = t[20339] ^ n[20340];
assign t[20341] = t[20340] ^ n[20341];
assign t[20342] = t[20341] ^ n[20342];
assign t[20343] = t[20342] ^ n[20343];
assign t[20344] = t[20343] ^ n[20344];
assign t[20345] = t[20344] ^ n[20345];
assign t[20346] = t[20345] ^ n[20346];
assign t[20347] = t[20346] ^ n[20347];
assign t[20348] = t[20347] ^ n[20348];
assign t[20349] = t[20348] ^ n[20349];
assign t[20350] = t[20349] ^ n[20350];
assign t[20351] = t[20350] ^ n[20351];
assign t[20352] = t[20351] ^ n[20352];
assign t[20353] = t[20352] ^ n[20353];
assign t[20354] = t[20353] ^ n[20354];
assign t[20355] = t[20354] ^ n[20355];
assign t[20356] = t[20355] ^ n[20356];
assign t[20357] = t[20356] ^ n[20357];
assign t[20358] = t[20357] ^ n[20358];
assign t[20359] = t[20358] ^ n[20359];
assign t[20360] = t[20359] ^ n[20360];
assign t[20361] = t[20360] ^ n[20361];
assign t[20362] = t[20361] ^ n[20362];
assign t[20363] = t[20362] ^ n[20363];
assign t[20364] = t[20363] ^ n[20364];
assign t[20365] = t[20364] ^ n[20365];
assign t[20366] = t[20365] ^ n[20366];
assign t[20367] = t[20366] ^ n[20367];
assign t[20368] = t[20367] ^ n[20368];
assign t[20369] = t[20368] ^ n[20369];
assign t[20370] = t[20369] ^ n[20370];
assign t[20371] = t[20370] ^ n[20371];
assign t[20372] = t[20371] ^ n[20372];
assign t[20373] = t[20372] ^ n[20373];
assign t[20374] = t[20373] ^ n[20374];
assign t[20375] = t[20374] ^ n[20375];
assign t[20376] = t[20375] ^ n[20376];
assign t[20377] = t[20376] ^ n[20377];
assign t[20378] = t[20377] ^ n[20378];
assign t[20379] = t[20378] ^ n[20379];
assign t[20380] = t[20379] ^ n[20380];
assign t[20381] = t[20380] ^ n[20381];
assign t[20382] = t[20381] ^ n[20382];
assign t[20383] = t[20382] ^ n[20383];
assign t[20384] = t[20383] ^ n[20384];
assign t[20385] = t[20384] ^ n[20385];
assign t[20386] = t[20385] ^ n[20386];
assign t[20387] = t[20386] ^ n[20387];
assign t[20388] = t[20387] ^ n[20388];
assign t[20389] = t[20388] ^ n[20389];
assign t[20390] = t[20389] ^ n[20390];
assign t[20391] = t[20390] ^ n[20391];
assign t[20392] = t[20391] ^ n[20392];
assign t[20393] = t[20392] ^ n[20393];
assign t[20394] = t[20393] ^ n[20394];
assign t[20395] = t[20394] ^ n[20395];
assign t[20396] = t[20395] ^ n[20396];
assign t[20397] = t[20396] ^ n[20397];
assign t[20398] = t[20397] ^ n[20398];
assign t[20399] = t[20398] ^ n[20399];
assign t[20400] = t[20399] ^ n[20400];
assign t[20401] = t[20400] ^ n[20401];
assign t[20402] = t[20401] ^ n[20402];
assign t[20403] = t[20402] ^ n[20403];
assign t[20404] = t[20403] ^ n[20404];
assign t[20405] = t[20404] ^ n[20405];
assign t[20406] = t[20405] ^ n[20406];
assign t[20407] = t[20406] ^ n[20407];
assign t[20408] = t[20407] ^ n[20408];
assign t[20409] = t[20408] ^ n[20409];
assign t[20410] = t[20409] ^ n[20410];
assign t[20411] = t[20410] ^ n[20411];
assign t[20412] = t[20411] ^ n[20412];
assign t[20413] = t[20412] ^ n[20413];
assign t[20414] = t[20413] ^ n[20414];
assign t[20415] = t[20414] ^ n[20415];
assign t[20416] = t[20415] ^ n[20416];
assign t[20417] = t[20416] ^ n[20417];
assign t[20418] = t[20417] ^ n[20418];
assign t[20419] = t[20418] ^ n[20419];
assign t[20420] = t[20419] ^ n[20420];
assign t[20421] = t[20420] ^ n[20421];
assign t[20422] = t[20421] ^ n[20422];
assign t[20423] = t[20422] ^ n[20423];
assign t[20424] = t[20423] ^ n[20424];
assign t[20425] = t[20424] ^ n[20425];
assign t[20426] = t[20425] ^ n[20426];
assign t[20427] = t[20426] ^ n[20427];
assign t[20428] = t[20427] ^ n[20428];
assign t[20429] = t[20428] ^ n[20429];
assign t[20430] = t[20429] ^ n[20430];
assign t[20431] = t[20430] ^ n[20431];
assign t[20432] = t[20431] ^ n[20432];
assign t[20433] = t[20432] ^ n[20433];
assign t[20434] = t[20433] ^ n[20434];
assign t[20435] = t[20434] ^ n[20435];
assign t[20436] = t[20435] ^ n[20436];
assign t[20437] = t[20436] ^ n[20437];
assign t[20438] = t[20437] ^ n[20438];
assign t[20439] = t[20438] ^ n[20439];
assign t[20440] = t[20439] ^ n[20440];
assign t[20441] = t[20440] ^ n[20441];
assign t[20442] = t[20441] ^ n[20442];
assign t[20443] = t[20442] ^ n[20443];
assign t[20444] = t[20443] ^ n[20444];
assign t[20445] = t[20444] ^ n[20445];
assign t[20446] = t[20445] ^ n[20446];
assign t[20447] = t[20446] ^ n[20447];
assign t[20448] = t[20447] ^ n[20448];
assign t[20449] = t[20448] ^ n[20449];
assign t[20450] = t[20449] ^ n[20450];
assign t[20451] = t[20450] ^ n[20451];
assign t[20452] = t[20451] ^ n[20452];
assign t[20453] = t[20452] ^ n[20453];
assign t[20454] = t[20453] ^ n[20454];
assign t[20455] = t[20454] ^ n[20455];
assign t[20456] = t[20455] ^ n[20456];
assign t[20457] = t[20456] ^ n[20457];
assign t[20458] = t[20457] ^ n[20458];
assign t[20459] = t[20458] ^ n[20459];
assign t[20460] = t[20459] ^ n[20460];
assign t[20461] = t[20460] ^ n[20461];
assign t[20462] = t[20461] ^ n[20462];
assign t[20463] = t[20462] ^ n[20463];
assign t[20464] = t[20463] ^ n[20464];
assign t[20465] = t[20464] ^ n[20465];
assign t[20466] = t[20465] ^ n[20466];
assign t[20467] = t[20466] ^ n[20467];
assign t[20468] = t[20467] ^ n[20468];
assign t[20469] = t[20468] ^ n[20469];
assign t[20470] = t[20469] ^ n[20470];
assign t[20471] = t[20470] ^ n[20471];
assign t[20472] = t[20471] ^ n[20472];
assign t[20473] = t[20472] ^ n[20473];
assign t[20474] = t[20473] ^ n[20474];
assign t[20475] = t[20474] ^ n[20475];
assign t[20476] = t[20475] ^ n[20476];
assign t[20477] = t[20476] ^ n[20477];
assign t[20478] = t[20477] ^ n[20478];
assign t[20479] = t[20478] ^ n[20479];
assign t[20480] = t[20479] ^ n[20480];
assign t[20481] = t[20480] ^ n[20481];
assign t[20482] = t[20481] ^ n[20482];
assign t[20483] = t[20482] ^ n[20483];
assign t[20484] = t[20483] ^ n[20484];
assign t[20485] = t[20484] ^ n[20485];
assign t[20486] = t[20485] ^ n[20486];
assign t[20487] = t[20486] ^ n[20487];
assign t[20488] = t[20487] ^ n[20488];
assign t[20489] = t[20488] ^ n[20489];
assign t[20490] = t[20489] ^ n[20490];
assign t[20491] = t[20490] ^ n[20491];
assign t[20492] = t[20491] ^ n[20492];
assign t[20493] = t[20492] ^ n[20493];
assign t[20494] = t[20493] ^ n[20494];
assign t[20495] = t[20494] ^ n[20495];
assign t[20496] = t[20495] ^ n[20496];
assign t[20497] = t[20496] ^ n[20497];
assign t[20498] = t[20497] ^ n[20498];
assign t[20499] = t[20498] ^ n[20499];
assign t[20500] = t[20499] ^ n[20500];
assign t[20501] = t[20500] ^ n[20501];
assign t[20502] = t[20501] ^ n[20502];
assign t[20503] = t[20502] ^ n[20503];
assign t[20504] = t[20503] ^ n[20504];
assign t[20505] = t[20504] ^ n[20505];
assign t[20506] = t[20505] ^ n[20506];
assign t[20507] = t[20506] ^ n[20507];
assign t[20508] = t[20507] ^ n[20508];
assign t[20509] = t[20508] ^ n[20509];
assign t[20510] = t[20509] ^ n[20510];
assign t[20511] = t[20510] ^ n[20511];
assign t[20512] = t[20511] ^ n[20512];
assign t[20513] = t[20512] ^ n[20513];
assign t[20514] = t[20513] ^ n[20514];
assign t[20515] = t[20514] ^ n[20515];
assign t[20516] = t[20515] ^ n[20516];
assign t[20517] = t[20516] ^ n[20517];
assign t[20518] = t[20517] ^ n[20518];
assign t[20519] = t[20518] ^ n[20519];
assign t[20520] = t[20519] ^ n[20520];
assign t[20521] = t[20520] ^ n[20521];
assign t[20522] = t[20521] ^ n[20522];
assign t[20523] = t[20522] ^ n[20523];
assign t[20524] = t[20523] ^ n[20524];
assign t[20525] = t[20524] ^ n[20525];
assign t[20526] = t[20525] ^ n[20526];
assign t[20527] = t[20526] ^ n[20527];
assign t[20528] = t[20527] ^ n[20528];
assign t[20529] = t[20528] ^ n[20529];
assign t[20530] = t[20529] ^ n[20530];
assign t[20531] = t[20530] ^ n[20531];
assign t[20532] = t[20531] ^ n[20532];
assign t[20533] = t[20532] ^ n[20533];
assign t[20534] = t[20533] ^ n[20534];
assign t[20535] = t[20534] ^ n[20535];
assign t[20536] = t[20535] ^ n[20536];
assign t[20537] = t[20536] ^ n[20537];
assign t[20538] = t[20537] ^ n[20538];
assign t[20539] = t[20538] ^ n[20539];
assign t[20540] = t[20539] ^ n[20540];
assign t[20541] = t[20540] ^ n[20541];
assign t[20542] = t[20541] ^ n[20542];
assign t[20543] = t[20542] ^ n[20543];
assign t[20544] = t[20543] ^ n[20544];
assign t[20545] = t[20544] ^ n[20545];
assign t[20546] = t[20545] ^ n[20546];
assign t[20547] = t[20546] ^ n[20547];
assign t[20548] = t[20547] ^ n[20548];
assign t[20549] = t[20548] ^ n[20549];
assign t[20550] = t[20549] ^ n[20550];
assign t[20551] = t[20550] ^ n[20551];
assign t[20552] = t[20551] ^ n[20552];
assign t[20553] = t[20552] ^ n[20553];
assign t[20554] = t[20553] ^ n[20554];
assign t[20555] = t[20554] ^ n[20555];
assign t[20556] = t[20555] ^ n[20556];
assign t[20557] = t[20556] ^ n[20557];
assign t[20558] = t[20557] ^ n[20558];
assign t[20559] = t[20558] ^ n[20559];
assign t[20560] = t[20559] ^ n[20560];
assign t[20561] = t[20560] ^ n[20561];
assign t[20562] = t[20561] ^ n[20562];
assign t[20563] = t[20562] ^ n[20563];
assign t[20564] = t[20563] ^ n[20564];
assign t[20565] = t[20564] ^ n[20565];
assign t[20566] = t[20565] ^ n[20566];
assign t[20567] = t[20566] ^ n[20567];
assign t[20568] = t[20567] ^ n[20568];
assign t[20569] = t[20568] ^ n[20569];
assign t[20570] = t[20569] ^ n[20570];
assign t[20571] = t[20570] ^ n[20571];
assign t[20572] = t[20571] ^ n[20572];
assign t[20573] = t[20572] ^ n[20573];
assign t[20574] = t[20573] ^ n[20574];
assign t[20575] = t[20574] ^ n[20575];
assign t[20576] = t[20575] ^ n[20576];
assign t[20577] = t[20576] ^ n[20577];
assign t[20578] = t[20577] ^ n[20578];
assign t[20579] = t[20578] ^ n[20579];
assign t[20580] = t[20579] ^ n[20580];
assign t[20581] = t[20580] ^ n[20581];
assign t[20582] = t[20581] ^ n[20582];
assign t[20583] = t[20582] ^ n[20583];
assign t[20584] = t[20583] ^ n[20584];
assign t[20585] = t[20584] ^ n[20585];
assign t[20586] = t[20585] ^ n[20586];
assign t[20587] = t[20586] ^ n[20587];
assign t[20588] = t[20587] ^ n[20588];
assign t[20589] = t[20588] ^ n[20589];
assign t[20590] = t[20589] ^ n[20590];
assign t[20591] = t[20590] ^ n[20591];
assign t[20592] = t[20591] ^ n[20592];
assign t[20593] = t[20592] ^ n[20593];
assign t[20594] = t[20593] ^ n[20594];
assign t[20595] = t[20594] ^ n[20595];
assign t[20596] = t[20595] ^ n[20596];
assign t[20597] = t[20596] ^ n[20597];
assign t[20598] = t[20597] ^ n[20598];
assign t[20599] = t[20598] ^ n[20599];
assign t[20600] = t[20599] ^ n[20600];
assign t[20601] = t[20600] ^ n[20601];
assign t[20602] = t[20601] ^ n[20602];
assign t[20603] = t[20602] ^ n[20603];
assign t[20604] = t[20603] ^ n[20604];
assign t[20605] = t[20604] ^ n[20605];
assign t[20606] = t[20605] ^ n[20606];
assign t[20607] = t[20606] ^ n[20607];
assign t[20608] = t[20607] ^ n[20608];
assign t[20609] = t[20608] ^ n[20609];
assign t[20610] = t[20609] ^ n[20610];
assign t[20611] = t[20610] ^ n[20611];
assign t[20612] = t[20611] ^ n[20612];
assign t[20613] = t[20612] ^ n[20613];
assign t[20614] = t[20613] ^ n[20614];
assign t[20615] = t[20614] ^ n[20615];
assign t[20616] = t[20615] ^ n[20616];
assign t[20617] = t[20616] ^ n[20617];
assign t[20618] = t[20617] ^ n[20618];
assign t[20619] = t[20618] ^ n[20619];
assign t[20620] = t[20619] ^ n[20620];
assign t[20621] = t[20620] ^ n[20621];
assign t[20622] = t[20621] ^ n[20622];
assign t[20623] = t[20622] ^ n[20623];
assign t[20624] = t[20623] ^ n[20624];
assign t[20625] = t[20624] ^ n[20625];
assign t[20626] = t[20625] ^ n[20626];
assign t[20627] = t[20626] ^ n[20627];
assign t[20628] = t[20627] ^ n[20628];
assign t[20629] = t[20628] ^ n[20629];
assign t[20630] = t[20629] ^ n[20630];
assign t[20631] = t[20630] ^ n[20631];
assign t[20632] = t[20631] ^ n[20632];
assign t[20633] = t[20632] ^ n[20633];
assign t[20634] = t[20633] ^ n[20634];
assign t[20635] = t[20634] ^ n[20635];
assign t[20636] = t[20635] ^ n[20636];
assign t[20637] = t[20636] ^ n[20637];
assign t[20638] = t[20637] ^ n[20638];
assign t[20639] = t[20638] ^ n[20639];
assign t[20640] = t[20639] ^ n[20640];
assign t[20641] = t[20640] ^ n[20641];
assign t[20642] = t[20641] ^ n[20642];
assign t[20643] = t[20642] ^ n[20643];
assign t[20644] = t[20643] ^ n[20644];
assign t[20645] = t[20644] ^ n[20645];
assign t[20646] = t[20645] ^ n[20646];
assign t[20647] = t[20646] ^ n[20647];
assign t[20648] = t[20647] ^ n[20648];
assign t[20649] = t[20648] ^ n[20649];
assign t[20650] = t[20649] ^ n[20650];
assign t[20651] = t[20650] ^ n[20651];
assign t[20652] = t[20651] ^ n[20652];
assign t[20653] = t[20652] ^ n[20653];
assign t[20654] = t[20653] ^ n[20654];
assign t[20655] = t[20654] ^ n[20655];
assign t[20656] = t[20655] ^ n[20656];
assign t[20657] = t[20656] ^ n[20657];
assign t[20658] = t[20657] ^ n[20658];
assign t[20659] = t[20658] ^ n[20659];
assign t[20660] = t[20659] ^ n[20660];
assign t[20661] = t[20660] ^ n[20661];
assign t[20662] = t[20661] ^ n[20662];
assign t[20663] = t[20662] ^ n[20663];
assign t[20664] = t[20663] ^ n[20664];
assign t[20665] = t[20664] ^ n[20665];
assign t[20666] = t[20665] ^ n[20666];
assign t[20667] = t[20666] ^ n[20667];
assign t[20668] = t[20667] ^ n[20668];
assign t[20669] = t[20668] ^ n[20669];
assign t[20670] = t[20669] ^ n[20670];
assign t[20671] = t[20670] ^ n[20671];
assign t[20672] = t[20671] ^ n[20672];
assign t[20673] = t[20672] ^ n[20673];
assign t[20674] = t[20673] ^ n[20674];
assign t[20675] = t[20674] ^ n[20675];
assign t[20676] = t[20675] ^ n[20676];
assign t[20677] = t[20676] ^ n[20677];
assign t[20678] = t[20677] ^ n[20678];
assign t[20679] = t[20678] ^ n[20679];
assign t[20680] = t[20679] ^ n[20680];
assign t[20681] = t[20680] ^ n[20681];
assign t[20682] = t[20681] ^ n[20682];
assign t[20683] = t[20682] ^ n[20683];
assign t[20684] = t[20683] ^ n[20684];
assign t[20685] = t[20684] ^ n[20685];
assign t[20686] = t[20685] ^ n[20686];
assign t[20687] = t[20686] ^ n[20687];
assign t[20688] = t[20687] ^ n[20688];
assign t[20689] = t[20688] ^ n[20689];
assign t[20690] = t[20689] ^ n[20690];
assign t[20691] = t[20690] ^ n[20691];
assign t[20692] = t[20691] ^ n[20692];
assign t[20693] = t[20692] ^ n[20693];
assign t[20694] = t[20693] ^ n[20694];
assign t[20695] = t[20694] ^ n[20695];
assign t[20696] = t[20695] ^ n[20696];
assign t[20697] = t[20696] ^ n[20697];
assign t[20698] = t[20697] ^ n[20698];
assign t[20699] = t[20698] ^ n[20699];
assign t[20700] = t[20699] ^ n[20700];
assign t[20701] = t[20700] ^ n[20701];
assign t[20702] = t[20701] ^ n[20702];
assign t[20703] = t[20702] ^ n[20703];
assign t[20704] = t[20703] ^ n[20704];
assign t[20705] = t[20704] ^ n[20705];
assign t[20706] = t[20705] ^ n[20706];
assign t[20707] = t[20706] ^ n[20707];
assign t[20708] = t[20707] ^ n[20708];
assign t[20709] = t[20708] ^ n[20709];
assign t[20710] = t[20709] ^ n[20710];
assign t[20711] = t[20710] ^ n[20711];
assign t[20712] = t[20711] ^ n[20712];
assign t[20713] = t[20712] ^ n[20713];
assign t[20714] = t[20713] ^ n[20714];
assign t[20715] = t[20714] ^ n[20715];
assign t[20716] = t[20715] ^ n[20716];
assign t[20717] = t[20716] ^ n[20717];
assign t[20718] = t[20717] ^ n[20718];
assign t[20719] = t[20718] ^ n[20719];
assign t[20720] = t[20719] ^ n[20720];
assign t[20721] = t[20720] ^ n[20721];
assign t[20722] = t[20721] ^ n[20722];
assign t[20723] = t[20722] ^ n[20723];
assign t[20724] = t[20723] ^ n[20724];
assign t[20725] = t[20724] ^ n[20725];
assign t[20726] = t[20725] ^ n[20726];
assign t[20727] = t[20726] ^ n[20727];
assign t[20728] = t[20727] ^ n[20728];
assign t[20729] = t[20728] ^ n[20729];
assign t[20730] = t[20729] ^ n[20730];
assign t[20731] = t[20730] ^ n[20731];
assign t[20732] = t[20731] ^ n[20732];
assign t[20733] = t[20732] ^ n[20733];
assign t[20734] = t[20733] ^ n[20734];
assign t[20735] = t[20734] ^ n[20735];
assign t[20736] = t[20735] ^ n[20736];
assign t[20737] = t[20736] ^ n[20737];
assign t[20738] = t[20737] ^ n[20738];
assign t[20739] = t[20738] ^ n[20739];
assign t[20740] = t[20739] ^ n[20740];
assign t[20741] = t[20740] ^ n[20741];
assign t[20742] = t[20741] ^ n[20742];
assign t[20743] = t[20742] ^ n[20743];
assign t[20744] = t[20743] ^ n[20744];
assign t[20745] = t[20744] ^ n[20745];
assign t[20746] = t[20745] ^ n[20746];
assign t[20747] = t[20746] ^ n[20747];
assign t[20748] = t[20747] ^ n[20748];
assign t[20749] = t[20748] ^ n[20749];
assign t[20750] = t[20749] ^ n[20750];
assign t[20751] = t[20750] ^ n[20751];
assign t[20752] = t[20751] ^ n[20752];
assign t[20753] = t[20752] ^ n[20753];
assign t[20754] = t[20753] ^ n[20754];
assign t[20755] = t[20754] ^ n[20755];
assign t[20756] = t[20755] ^ n[20756];
assign t[20757] = t[20756] ^ n[20757];
assign t[20758] = t[20757] ^ n[20758];
assign t[20759] = t[20758] ^ n[20759];
assign t[20760] = t[20759] ^ n[20760];
assign t[20761] = t[20760] ^ n[20761];
assign t[20762] = t[20761] ^ n[20762];
assign t[20763] = t[20762] ^ n[20763];
assign t[20764] = t[20763] ^ n[20764];
assign t[20765] = t[20764] ^ n[20765];
assign t[20766] = t[20765] ^ n[20766];
assign t[20767] = t[20766] ^ n[20767];
assign t[20768] = t[20767] ^ n[20768];
assign t[20769] = t[20768] ^ n[20769];
assign t[20770] = t[20769] ^ n[20770];
assign t[20771] = t[20770] ^ n[20771];
assign t[20772] = t[20771] ^ n[20772];
assign t[20773] = t[20772] ^ n[20773];
assign t[20774] = t[20773] ^ n[20774];
assign t[20775] = t[20774] ^ n[20775];
assign t[20776] = t[20775] ^ n[20776];
assign t[20777] = t[20776] ^ n[20777];
assign t[20778] = t[20777] ^ n[20778];
assign t[20779] = t[20778] ^ n[20779];
assign t[20780] = t[20779] ^ n[20780];
assign t[20781] = t[20780] ^ n[20781];
assign t[20782] = t[20781] ^ n[20782];
assign t[20783] = t[20782] ^ n[20783];
assign t[20784] = t[20783] ^ n[20784];
assign t[20785] = t[20784] ^ n[20785];
assign t[20786] = t[20785] ^ n[20786];
assign t[20787] = t[20786] ^ n[20787];
assign t[20788] = t[20787] ^ n[20788];
assign t[20789] = t[20788] ^ n[20789];
assign t[20790] = t[20789] ^ n[20790];
assign t[20791] = t[20790] ^ n[20791];
assign t[20792] = t[20791] ^ n[20792];
assign t[20793] = t[20792] ^ n[20793];
assign t[20794] = t[20793] ^ n[20794];
assign t[20795] = t[20794] ^ n[20795];
assign t[20796] = t[20795] ^ n[20796];
assign t[20797] = t[20796] ^ n[20797];
assign t[20798] = t[20797] ^ n[20798];
assign t[20799] = t[20798] ^ n[20799];
assign t[20800] = t[20799] ^ n[20800];
assign t[20801] = t[20800] ^ n[20801];
assign t[20802] = t[20801] ^ n[20802];
assign t[20803] = t[20802] ^ n[20803];
assign t[20804] = t[20803] ^ n[20804];
assign t[20805] = t[20804] ^ n[20805];
assign t[20806] = t[20805] ^ n[20806];
assign t[20807] = t[20806] ^ n[20807];
assign t[20808] = t[20807] ^ n[20808];
assign t[20809] = t[20808] ^ n[20809];
assign t[20810] = t[20809] ^ n[20810];
assign t[20811] = t[20810] ^ n[20811];
assign t[20812] = t[20811] ^ n[20812];
assign t[20813] = t[20812] ^ n[20813];
assign t[20814] = t[20813] ^ n[20814];
assign t[20815] = t[20814] ^ n[20815];
assign t[20816] = t[20815] ^ n[20816];
assign t[20817] = t[20816] ^ n[20817];
assign t[20818] = t[20817] ^ n[20818];
assign t[20819] = t[20818] ^ n[20819];
assign t[20820] = t[20819] ^ n[20820];
assign t[20821] = t[20820] ^ n[20821];
assign t[20822] = t[20821] ^ n[20822];
assign t[20823] = t[20822] ^ n[20823];
assign t[20824] = t[20823] ^ n[20824];
assign t[20825] = t[20824] ^ n[20825];
assign t[20826] = t[20825] ^ n[20826];
assign t[20827] = t[20826] ^ n[20827];
assign t[20828] = t[20827] ^ n[20828];
assign t[20829] = t[20828] ^ n[20829];
assign t[20830] = t[20829] ^ n[20830];
assign t[20831] = t[20830] ^ n[20831];
assign t[20832] = t[20831] ^ n[20832];
assign t[20833] = t[20832] ^ n[20833];
assign t[20834] = t[20833] ^ n[20834];
assign t[20835] = t[20834] ^ n[20835];
assign t[20836] = t[20835] ^ n[20836];
assign t[20837] = t[20836] ^ n[20837];
assign t[20838] = t[20837] ^ n[20838];
assign t[20839] = t[20838] ^ n[20839];
assign t[20840] = t[20839] ^ n[20840];
assign t[20841] = t[20840] ^ n[20841];
assign t[20842] = t[20841] ^ n[20842];
assign t[20843] = t[20842] ^ n[20843];
assign t[20844] = t[20843] ^ n[20844];
assign t[20845] = t[20844] ^ n[20845];
assign t[20846] = t[20845] ^ n[20846];
assign t[20847] = t[20846] ^ n[20847];
assign t[20848] = t[20847] ^ n[20848];
assign t[20849] = t[20848] ^ n[20849];
assign t[20850] = t[20849] ^ n[20850];
assign t[20851] = t[20850] ^ n[20851];
assign t[20852] = t[20851] ^ n[20852];
assign t[20853] = t[20852] ^ n[20853];
assign t[20854] = t[20853] ^ n[20854];
assign t[20855] = t[20854] ^ n[20855];
assign t[20856] = t[20855] ^ n[20856];
assign t[20857] = t[20856] ^ n[20857];
assign t[20858] = t[20857] ^ n[20858];
assign t[20859] = t[20858] ^ n[20859];
assign t[20860] = t[20859] ^ n[20860];
assign t[20861] = t[20860] ^ n[20861];
assign t[20862] = t[20861] ^ n[20862];
assign t[20863] = t[20862] ^ n[20863];
assign t[20864] = t[20863] ^ n[20864];
assign t[20865] = t[20864] ^ n[20865];
assign t[20866] = t[20865] ^ n[20866];
assign t[20867] = t[20866] ^ n[20867];
assign t[20868] = t[20867] ^ n[20868];
assign t[20869] = t[20868] ^ n[20869];
assign t[20870] = t[20869] ^ n[20870];
assign t[20871] = t[20870] ^ n[20871];
assign t[20872] = t[20871] ^ n[20872];
assign t[20873] = t[20872] ^ n[20873];
assign t[20874] = t[20873] ^ n[20874];
assign t[20875] = t[20874] ^ n[20875];
assign t[20876] = t[20875] ^ n[20876];
assign t[20877] = t[20876] ^ n[20877];
assign t[20878] = t[20877] ^ n[20878];
assign t[20879] = t[20878] ^ n[20879];
assign t[20880] = t[20879] ^ n[20880];
assign t[20881] = t[20880] ^ n[20881];
assign t[20882] = t[20881] ^ n[20882];
assign t[20883] = t[20882] ^ n[20883];
assign t[20884] = t[20883] ^ n[20884];
assign t[20885] = t[20884] ^ n[20885];
assign t[20886] = t[20885] ^ n[20886];
assign t[20887] = t[20886] ^ n[20887];
assign t[20888] = t[20887] ^ n[20888];
assign t[20889] = t[20888] ^ n[20889];
assign t[20890] = t[20889] ^ n[20890];
assign t[20891] = t[20890] ^ n[20891];
assign t[20892] = t[20891] ^ n[20892];
assign t[20893] = t[20892] ^ n[20893];
assign t[20894] = t[20893] ^ n[20894];
assign t[20895] = t[20894] ^ n[20895];
assign t[20896] = t[20895] ^ n[20896];
assign t[20897] = t[20896] ^ n[20897];
assign t[20898] = t[20897] ^ n[20898];
assign t[20899] = t[20898] ^ n[20899];
assign t[20900] = t[20899] ^ n[20900];
assign t[20901] = t[20900] ^ n[20901];
assign t[20902] = t[20901] ^ n[20902];
assign t[20903] = t[20902] ^ n[20903];
assign t[20904] = t[20903] ^ n[20904];
assign t[20905] = t[20904] ^ n[20905];
assign t[20906] = t[20905] ^ n[20906];
assign t[20907] = t[20906] ^ n[20907];
assign t[20908] = t[20907] ^ n[20908];
assign t[20909] = t[20908] ^ n[20909];
assign t[20910] = t[20909] ^ n[20910];
assign t[20911] = t[20910] ^ n[20911];
assign t[20912] = t[20911] ^ n[20912];
assign t[20913] = t[20912] ^ n[20913];
assign t[20914] = t[20913] ^ n[20914];
assign t[20915] = t[20914] ^ n[20915];
assign t[20916] = t[20915] ^ n[20916];
assign t[20917] = t[20916] ^ n[20917];
assign t[20918] = t[20917] ^ n[20918];
assign t[20919] = t[20918] ^ n[20919];
assign t[20920] = t[20919] ^ n[20920];
assign t[20921] = t[20920] ^ n[20921];
assign t[20922] = t[20921] ^ n[20922];
assign t[20923] = t[20922] ^ n[20923];
assign t[20924] = t[20923] ^ n[20924];
assign t[20925] = t[20924] ^ n[20925];
assign t[20926] = t[20925] ^ n[20926];
assign t[20927] = t[20926] ^ n[20927];
assign t[20928] = t[20927] ^ n[20928];
assign t[20929] = t[20928] ^ n[20929];
assign t[20930] = t[20929] ^ n[20930];
assign t[20931] = t[20930] ^ n[20931];
assign t[20932] = t[20931] ^ n[20932];
assign t[20933] = t[20932] ^ n[20933];
assign t[20934] = t[20933] ^ n[20934];
assign t[20935] = t[20934] ^ n[20935];
assign t[20936] = t[20935] ^ n[20936];
assign t[20937] = t[20936] ^ n[20937];
assign t[20938] = t[20937] ^ n[20938];
assign t[20939] = t[20938] ^ n[20939];
assign t[20940] = t[20939] ^ n[20940];
assign t[20941] = t[20940] ^ n[20941];
assign t[20942] = t[20941] ^ n[20942];
assign t[20943] = t[20942] ^ n[20943];
assign t[20944] = t[20943] ^ n[20944];
assign t[20945] = t[20944] ^ n[20945];
assign t[20946] = t[20945] ^ n[20946];
assign t[20947] = t[20946] ^ n[20947];
assign t[20948] = t[20947] ^ n[20948];
assign t[20949] = t[20948] ^ n[20949];
assign t[20950] = t[20949] ^ n[20950];
assign t[20951] = t[20950] ^ n[20951];
assign t[20952] = t[20951] ^ n[20952];
assign t[20953] = t[20952] ^ n[20953];
assign t[20954] = t[20953] ^ n[20954];
assign t[20955] = t[20954] ^ n[20955];
assign t[20956] = t[20955] ^ n[20956];
assign t[20957] = t[20956] ^ n[20957];
assign t[20958] = t[20957] ^ n[20958];
assign t[20959] = t[20958] ^ n[20959];
assign t[20960] = t[20959] ^ n[20960];
assign t[20961] = t[20960] ^ n[20961];
assign t[20962] = t[20961] ^ n[20962];
assign t[20963] = t[20962] ^ n[20963];
assign t[20964] = t[20963] ^ n[20964];
assign t[20965] = t[20964] ^ n[20965];
assign t[20966] = t[20965] ^ n[20966];
assign t[20967] = t[20966] ^ n[20967];
assign t[20968] = t[20967] ^ n[20968];
assign t[20969] = t[20968] ^ n[20969];
assign t[20970] = t[20969] ^ n[20970];
assign t[20971] = t[20970] ^ n[20971];
assign t[20972] = t[20971] ^ n[20972];
assign t[20973] = t[20972] ^ n[20973];
assign t[20974] = t[20973] ^ n[20974];
assign t[20975] = t[20974] ^ n[20975];
assign t[20976] = t[20975] ^ n[20976];
assign t[20977] = t[20976] ^ n[20977];
assign t[20978] = t[20977] ^ n[20978];
assign t[20979] = t[20978] ^ n[20979];
assign t[20980] = t[20979] ^ n[20980];
assign t[20981] = t[20980] ^ n[20981];
assign t[20982] = t[20981] ^ n[20982];
assign t[20983] = t[20982] ^ n[20983];
assign t[20984] = t[20983] ^ n[20984];
assign t[20985] = t[20984] ^ n[20985];
assign t[20986] = t[20985] ^ n[20986];
assign t[20987] = t[20986] ^ n[20987];
assign t[20988] = t[20987] ^ n[20988];
assign t[20989] = t[20988] ^ n[20989];
assign t[20990] = t[20989] ^ n[20990];
assign t[20991] = t[20990] ^ n[20991];
assign t[20992] = t[20991] ^ n[20992];
assign t[20993] = t[20992] ^ n[20993];
assign t[20994] = t[20993] ^ n[20994];
assign t[20995] = t[20994] ^ n[20995];
assign t[20996] = t[20995] ^ n[20996];
assign t[20997] = t[20996] ^ n[20997];
assign t[20998] = t[20997] ^ n[20998];
assign t[20999] = t[20998] ^ n[20999];
assign t[21000] = t[20999] ^ n[21000];
assign t[21001] = t[21000] ^ n[21001];
assign t[21002] = t[21001] ^ n[21002];
assign t[21003] = t[21002] ^ n[21003];
assign t[21004] = t[21003] ^ n[21004];
assign t[21005] = t[21004] ^ n[21005];
assign t[21006] = t[21005] ^ n[21006];
assign t[21007] = t[21006] ^ n[21007];
assign t[21008] = t[21007] ^ n[21008];
assign t[21009] = t[21008] ^ n[21009];
assign t[21010] = t[21009] ^ n[21010];
assign t[21011] = t[21010] ^ n[21011];
assign t[21012] = t[21011] ^ n[21012];
assign t[21013] = t[21012] ^ n[21013];
assign t[21014] = t[21013] ^ n[21014];
assign t[21015] = t[21014] ^ n[21015];
assign t[21016] = t[21015] ^ n[21016];
assign t[21017] = t[21016] ^ n[21017];
assign t[21018] = t[21017] ^ n[21018];
assign t[21019] = t[21018] ^ n[21019];
assign t[21020] = t[21019] ^ n[21020];
assign t[21021] = t[21020] ^ n[21021];
assign t[21022] = t[21021] ^ n[21022];
assign t[21023] = t[21022] ^ n[21023];
assign t[21024] = t[21023] ^ n[21024];
assign t[21025] = t[21024] ^ n[21025];
assign t[21026] = t[21025] ^ n[21026];
assign t[21027] = t[21026] ^ n[21027];
assign t[21028] = t[21027] ^ n[21028];
assign t[21029] = t[21028] ^ n[21029];
assign t[21030] = t[21029] ^ n[21030];
assign t[21031] = t[21030] ^ n[21031];
assign t[21032] = t[21031] ^ n[21032];
assign t[21033] = t[21032] ^ n[21033];
assign t[21034] = t[21033] ^ n[21034];
assign t[21035] = t[21034] ^ n[21035];
assign t[21036] = t[21035] ^ n[21036];
assign t[21037] = t[21036] ^ n[21037];
assign t[21038] = t[21037] ^ n[21038];
assign t[21039] = t[21038] ^ n[21039];
assign t[21040] = t[21039] ^ n[21040];
assign t[21041] = t[21040] ^ n[21041];
assign t[21042] = t[21041] ^ n[21042];
assign t[21043] = t[21042] ^ n[21043];
assign t[21044] = t[21043] ^ n[21044];
assign t[21045] = t[21044] ^ n[21045];
assign t[21046] = t[21045] ^ n[21046];
assign t[21047] = t[21046] ^ n[21047];
assign t[21048] = t[21047] ^ n[21048];
assign t[21049] = t[21048] ^ n[21049];
assign t[21050] = t[21049] ^ n[21050];
assign t[21051] = t[21050] ^ n[21051];
assign t[21052] = t[21051] ^ n[21052];
assign t[21053] = t[21052] ^ n[21053];
assign t[21054] = t[21053] ^ n[21054];
assign t[21055] = t[21054] ^ n[21055];
assign t[21056] = t[21055] ^ n[21056];
assign t[21057] = t[21056] ^ n[21057];
assign t[21058] = t[21057] ^ n[21058];
assign t[21059] = t[21058] ^ n[21059];
assign t[21060] = t[21059] ^ n[21060];
assign t[21061] = t[21060] ^ n[21061];
assign t[21062] = t[21061] ^ n[21062];
assign t[21063] = t[21062] ^ n[21063];
assign t[21064] = t[21063] ^ n[21064];
assign t[21065] = t[21064] ^ n[21065];
assign t[21066] = t[21065] ^ n[21066];
assign t[21067] = t[21066] ^ n[21067];
assign t[21068] = t[21067] ^ n[21068];
assign t[21069] = t[21068] ^ n[21069];
assign t[21070] = t[21069] ^ n[21070];
assign t[21071] = t[21070] ^ n[21071];
assign t[21072] = t[21071] ^ n[21072];
assign t[21073] = t[21072] ^ n[21073];
assign t[21074] = t[21073] ^ n[21074];
assign t[21075] = t[21074] ^ n[21075];
assign t[21076] = t[21075] ^ n[21076];
assign t[21077] = t[21076] ^ n[21077];
assign t[21078] = t[21077] ^ n[21078];
assign t[21079] = t[21078] ^ n[21079];
assign t[21080] = t[21079] ^ n[21080];
assign t[21081] = t[21080] ^ n[21081];
assign t[21082] = t[21081] ^ n[21082];
assign t[21083] = t[21082] ^ n[21083];
assign t[21084] = t[21083] ^ n[21084];
assign t[21085] = t[21084] ^ n[21085];
assign t[21086] = t[21085] ^ n[21086];
assign t[21087] = t[21086] ^ n[21087];
assign t[21088] = t[21087] ^ n[21088];
assign t[21089] = t[21088] ^ n[21089];
assign t[21090] = t[21089] ^ n[21090];
assign t[21091] = t[21090] ^ n[21091];
assign t[21092] = t[21091] ^ n[21092];
assign t[21093] = t[21092] ^ n[21093];
assign t[21094] = t[21093] ^ n[21094];
assign t[21095] = t[21094] ^ n[21095];
assign t[21096] = t[21095] ^ n[21096];
assign t[21097] = t[21096] ^ n[21097];
assign t[21098] = t[21097] ^ n[21098];
assign t[21099] = t[21098] ^ n[21099];
assign t[21100] = t[21099] ^ n[21100];
assign t[21101] = t[21100] ^ n[21101];
assign t[21102] = t[21101] ^ n[21102];
assign t[21103] = t[21102] ^ n[21103];
assign t[21104] = t[21103] ^ n[21104];
assign t[21105] = t[21104] ^ n[21105];
assign t[21106] = t[21105] ^ n[21106];
assign t[21107] = t[21106] ^ n[21107];
assign t[21108] = t[21107] ^ n[21108];
assign t[21109] = t[21108] ^ n[21109];
assign t[21110] = t[21109] ^ n[21110];
assign t[21111] = t[21110] ^ n[21111];
assign t[21112] = t[21111] ^ n[21112];
assign t[21113] = t[21112] ^ n[21113];
assign t[21114] = t[21113] ^ n[21114];
assign t[21115] = t[21114] ^ n[21115];
assign t[21116] = t[21115] ^ n[21116];
assign t[21117] = t[21116] ^ n[21117];
assign t[21118] = t[21117] ^ n[21118];
assign t[21119] = t[21118] ^ n[21119];
assign t[21120] = t[21119] ^ n[21120];
assign t[21121] = t[21120] ^ n[21121];
assign t[21122] = t[21121] ^ n[21122];
assign t[21123] = t[21122] ^ n[21123];
assign t[21124] = t[21123] ^ n[21124];
assign t[21125] = t[21124] ^ n[21125];
assign t[21126] = t[21125] ^ n[21126];
assign t[21127] = t[21126] ^ n[21127];
assign t[21128] = t[21127] ^ n[21128];
assign t[21129] = t[21128] ^ n[21129];
assign t[21130] = t[21129] ^ n[21130];
assign t[21131] = t[21130] ^ n[21131];
assign t[21132] = t[21131] ^ n[21132];
assign t[21133] = t[21132] ^ n[21133];
assign t[21134] = t[21133] ^ n[21134];
assign t[21135] = t[21134] ^ n[21135];
assign t[21136] = t[21135] ^ n[21136];
assign t[21137] = t[21136] ^ n[21137];
assign t[21138] = t[21137] ^ n[21138];
assign t[21139] = t[21138] ^ n[21139];
assign t[21140] = t[21139] ^ n[21140];
assign t[21141] = t[21140] ^ n[21141];
assign t[21142] = t[21141] ^ n[21142];
assign t[21143] = t[21142] ^ n[21143];
assign t[21144] = t[21143] ^ n[21144];
assign t[21145] = t[21144] ^ n[21145];
assign t[21146] = t[21145] ^ n[21146];
assign t[21147] = t[21146] ^ n[21147];
assign t[21148] = t[21147] ^ n[21148];
assign t[21149] = t[21148] ^ n[21149];
assign t[21150] = t[21149] ^ n[21150];
assign t[21151] = t[21150] ^ n[21151];
assign t[21152] = t[21151] ^ n[21152];
assign t[21153] = t[21152] ^ n[21153];
assign t[21154] = t[21153] ^ n[21154];
assign t[21155] = t[21154] ^ n[21155];
assign t[21156] = t[21155] ^ n[21156];
assign t[21157] = t[21156] ^ n[21157];
assign t[21158] = t[21157] ^ n[21158];
assign t[21159] = t[21158] ^ n[21159];
assign t[21160] = t[21159] ^ n[21160];
assign t[21161] = t[21160] ^ n[21161];
assign t[21162] = t[21161] ^ n[21162];
assign t[21163] = t[21162] ^ n[21163];
assign t[21164] = t[21163] ^ n[21164];
assign t[21165] = t[21164] ^ n[21165];
assign t[21166] = t[21165] ^ n[21166];
assign t[21167] = t[21166] ^ n[21167];
assign t[21168] = t[21167] ^ n[21168];
assign t[21169] = t[21168] ^ n[21169];
assign t[21170] = t[21169] ^ n[21170];
assign t[21171] = t[21170] ^ n[21171];
assign t[21172] = t[21171] ^ n[21172];
assign t[21173] = t[21172] ^ n[21173];
assign t[21174] = t[21173] ^ n[21174];
assign t[21175] = t[21174] ^ n[21175];
assign t[21176] = t[21175] ^ n[21176];
assign t[21177] = t[21176] ^ n[21177];
assign t[21178] = t[21177] ^ n[21178];
assign t[21179] = t[21178] ^ n[21179];
assign t[21180] = t[21179] ^ n[21180];
assign t[21181] = t[21180] ^ n[21181];
assign t[21182] = t[21181] ^ n[21182];
assign t[21183] = t[21182] ^ n[21183];
assign t[21184] = t[21183] ^ n[21184];
assign t[21185] = t[21184] ^ n[21185];
assign t[21186] = t[21185] ^ n[21186];
assign t[21187] = t[21186] ^ n[21187];
assign t[21188] = t[21187] ^ n[21188];
assign t[21189] = t[21188] ^ n[21189];
assign t[21190] = t[21189] ^ n[21190];
assign t[21191] = t[21190] ^ n[21191];
assign t[21192] = t[21191] ^ n[21192];
assign t[21193] = t[21192] ^ n[21193];
assign t[21194] = t[21193] ^ n[21194];
assign t[21195] = t[21194] ^ n[21195];
assign t[21196] = t[21195] ^ n[21196];
assign t[21197] = t[21196] ^ n[21197];
assign t[21198] = t[21197] ^ n[21198];
assign t[21199] = t[21198] ^ n[21199];
assign t[21200] = t[21199] ^ n[21200];
assign t[21201] = t[21200] ^ n[21201];
assign t[21202] = t[21201] ^ n[21202];
assign t[21203] = t[21202] ^ n[21203];
assign t[21204] = t[21203] ^ n[21204];
assign t[21205] = t[21204] ^ n[21205];
assign t[21206] = t[21205] ^ n[21206];
assign t[21207] = t[21206] ^ n[21207];
assign t[21208] = t[21207] ^ n[21208];
assign t[21209] = t[21208] ^ n[21209];
assign t[21210] = t[21209] ^ n[21210];
assign t[21211] = t[21210] ^ n[21211];
assign t[21212] = t[21211] ^ n[21212];
assign t[21213] = t[21212] ^ n[21213];
assign t[21214] = t[21213] ^ n[21214];
assign t[21215] = t[21214] ^ n[21215];
assign t[21216] = t[21215] ^ n[21216];
assign t[21217] = t[21216] ^ n[21217];
assign t[21218] = t[21217] ^ n[21218];
assign t[21219] = t[21218] ^ n[21219];
assign t[21220] = t[21219] ^ n[21220];
assign t[21221] = t[21220] ^ n[21221];
assign t[21222] = t[21221] ^ n[21222];
assign t[21223] = t[21222] ^ n[21223];
assign t[21224] = t[21223] ^ n[21224];
assign t[21225] = t[21224] ^ n[21225];
assign t[21226] = t[21225] ^ n[21226];
assign t[21227] = t[21226] ^ n[21227];
assign t[21228] = t[21227] ^ n[21228];
assign t[21229] = t[21228] ^ n[21229];
assign t[21230] = t[21229] ^ n[21230];
assign t[21231] = t[21230] ^ n[21231];
assign t[21232] = t[21231] ^ n[21232];
assign t[21233] = t[21232] ^ n[21233];
assign t[21234] = t[21233] ^ n[21234];
assign t[21235] = t[21234] ^ n[21235];
assign t[21236] = t[21235] ^ n[21236];
assign t[21237] = t[21236] ^ n[21237];
assign t[21238] = t[21237] ^ n[21238];
assign t[21239] = t[21238] ^ n[21239];
assign t[21240] = t[21239] ^ n[21240];
assign t[21241] = t[21240] ^ n[21241];
assign t[21242] = t[21241] ^ n[21242];
assign t[21243] = t[21242] ^ n[21243];
assign t[21244] = t[21243] ^ n[21244];
assign t[21245] = t[21244] ^ n[21245];
assign t[21246] = t[21245] ^ n[21246];
assign t[21247] = t[21246] ^ n[21247];
assign t[21248] = t[21247] ^ n[21248];
assign t[21249] = t[21248] ^ n[21249];
assign t[21250] = t[21249] ^ n[21250];
assign t[21251] = t[21250] ^ n[21251];
assign t[21252] = t[21251] ^ n[21252];
assign t[21253] = t[21252] ^ n[21253];
assign t[21254] = t[21253] ^ n[21254];
assign t[21255] = t[21254] ^ n[21255];
assign t[21256] = t[21255] ^ n[21256];
assign t[21257] = t[21256] ^ n[21257];
assign t[21258] = t[21257] ^ n[21258];
assign t[21259] = t[21258] ^ n[21259];
assign t[21260] = t[21259] ^ n[21260];
assign t[21261] = t[21260] ^ n[21261];
assign t[21262] = t[21261] ^ n[21262];
assign t[21263] = t[21262] ^ n[21263];
assign t[21264] = t[21263] ^ n[21264];
assign t[21265] = t[21264] ^ n[21265];
assign t[21266] = t[21265] ^ n[21266];
assign t[21267] = t[21266] ^ n[21267];
assign t[21268] = t[21267] ^ n[21268];
assign t[21269] = t[21268] ^ n[21269];
assign t[21270] = t[21269] ^ n[21270];
assign t[21271] = t[21270] ^ n[21271];
assign t[21272] = t[21271] ^ n[21272];
assign t[21273] = t[21272] ^ n[21273];
assign t[21274] = t[21273] ^ n[21274];
assign t[21275] = t[21274] ^ n[21275];
assign t[21276] = t[21275] ^ n[21276];
assign t[21277] = t[21276] ^ n[21277];
assign t[21278] = t[21277] ^ n[21278];
assign t[21279] = t[21278] ^ n[21279];
assign t[21280] = t[21279] ^ n[21280];
assign t[21281] = t[21280] ^ n[21281];
assign t[21282] = t[21281] ^ n[21282];
assign t[21283] = t[21282] ^ n[21283];
assign t[21284] = t[21283] ^ n[21284];
assign t[21285] = t[21284] ^ n[21285];
assign t[21286] = t[21285] ^ n[21286];
assign t[21287] = t[21286] ^ n[21287];
assign t[21288] = t[21287] ^ n[21288];
assign t[21289] = t[21288] ^ n[21289];
assign t[21290] = t[21289] ^ n[21290];
assign t[21291] = t[21290] ^ n[21291];
assign t[21292] = t[21291] ^ n[21292];
assign t[21293] = t[21292] ^ n[21293];
assign t[21294] = t[21293] ^ n[21294];
assign t[21295] = t[21294] ^ n[21295];
assign t[21296] = t[21295] ^ n[21296];
assign t[21297] = t[21296] ^ n[21297];
assign t[21298] = t[21297] ^ n[21298];
assign t[21299] = t[21298] ^ n[21299];
assign t[21300] = t[21299] ^ n[21300];
assign t[21301] = t[21300] ^ n[21301];
assign t[21302] = t[21301] ^ n[21302];
assign t[21303] = t[21302] ^ n[21303];
assign t[21304] = t[21303] ^ n[21304];
assign t[21305] = t[21304] ^ n[21305];
assign t[21306] = t[21305] ^ n[21306];
assign t[21307] = t[21306] ^ n[21307];
assign t[21308] = t[21307] ^ n[21308];
assign t[21309] = t[21308] ^ n[21309];
assign t[21310] = t[21309] ^ n[21310];
assign t[21311] = t[21310] ^ n[21311];
assign t[21312] = t[21311] ^ n[21312];
assign t[21313] = t[21312] ^ n[21313];
assign t[21314] = t[21313] ^ n[21314];
assign t[21315] = t[21314] ^ n[21315];
assign t[21316] = t[21315] ^ n[21316];
assign t[21317] = t[21316] ^ n[21317];
assign t[21318] = t[21317] ^ n[21318];
assign t[21319] = t[21318] ^ n[21319];
assign t[21320] = t[21319] ^ n[21320];
assign t[21321] = t[21320] ^ n[21321];
assign t[21322] = t[21321] ^ n[21322];
assign t[21323] = t[21322] ^ n[21323];
assign t[21324] = t[21323] ^ n[21324];
assign t[21325] = t[21324] ^ n[21325];
assign t[21326] = t[21325] ^ n[21326];
assign t[21327] = t[21326] ^ n[21327];
assign t[21328] = t[21327] ^ n[21328];
assign t[21329] = t[21328] ^ n[21329];
assign t[21330] = t[21329] ^ n[21330];
assign t[21331] = t[21330] ^ n[21331];
assign t[21332] = t[21331] ^ n[21332];
assign t[21333] = t[21332] ^ n[21333];
assign t[21334] = t[21333] ^ n[21334];
assign t[21335] = t[21334] ^ n[21335];
assign t[21336] = t[21335] ^ n[21336];
assign t[21337] = t[21336] ^ n[21337];
assign t[21338] = t[21337] ^ n[21338];
assign t[21339] = t[21338] ^ n[21339];
assign t[21340] = t[21339] ^ n[21340];
assign t[21341] = t[21340] ^ n[21341];
assign t[21342] = t[21341] ^ n[21342];
assign t[21343] = t[21342] ^ n[21343];
assign t[21344] = t[21343] ^ n[21344];
assign t[21345] = t[21344] ^ n[21345];
assign t[21346] = t[21345] ^ n[21346];
assign t[21347] = t[21346] ^ n[21347];
assign t[21348] = t[21347] ^ n[21348];
assign t[21349] = t[21348] ^ n[21349];
assign t[21350] = t[21349] ^ n[21350];
assign t[21351] = t[21350] ^ n[21351];
assign t[21352] = t[21351] ^ n[21352];
assign t[21353] = t[21352] ^ n[21353];
assign t[21354] = t[21353] ^ n[21354];
assign t[21355] = t[21354] ^ n[21355];
assign t[21356] = t[21355] ^ n[21356];
assign t[21357] = t[21356] ^ n[21357];
assign t[21358] = t[21357] ^ n[21358];
assign t[21359] = t[21358] ^ n[21359];
assign t[21360] = t[21359] ^ n[21360];
assign t[21361] = t[21360] ^ n[21361];
assign t[21362] = t[21361] ^ n[21362];
assign t[21363] = t[21362] ^ n[21363];
assign t[21364] = t[21363] ^ n[21364];
assign t[21365] = t[21364] ^ n[21365];
assign t[21366] = t[21365] ^ n[21366];
assign t[21367] = t[21366] ^ n[21367];
assign t[21368] = t[21367] ^ n[21368];
assign t[21369] = t[21368] ^ n[21369];
assign t[21370] = t[21369] ^ n[21370];
assign t[21371] = t[21370] ^ n[21371];
assign t[21372] = t[21371] ^ n[21372];
assign t[21373] = t[21372] ^ n[21373];
assign t[21374] = t[21373] ^ n[21374];
assign t[21375] = t[21374] ^ n[21375];
assign t[21376] = t[21375] ^ n[21376];
assign t[21377] = t[21376] ^ n[21377];
assign t[21378] = t[21377] ^ n[21378];
assign t[21379] = t[21378] ^ n[21379];
assign t[21380] = t[21379] ^ n[21380];
assign t[21381] = t[21380] ^ n[21381];
assign t[21382] = t[21381] ^ n[21382];
assign t[21383] = t[21382] ^ n[21383];
assign t[21384] = t[21383] ^ n[21384];
assign t[21385] = t[21384] ^ n[21385];
assign t[21386] = t[21385] ^ n[21386];
assign t[21387] = t[21386] ^ n[21387];
assign t[21388] = t[21387] ^ n[21388];
assign t[21389] = t[21388] ^ n[21389];
assign t[21390] = t[21389] ^ n[21390];
assign t[21391] = t[21390] ^ n[21391];
assign t[21392] = t[21391] ^ n[21392];
assign t[21393] = t[21392] ^ n[21393];
assign t[21394] = t[21393] ^ n[21394];
assign t[21395] = t[21394] ^ n[21395];
assign t[21396] = t[21395] ^ n[21396];
assign t[21397] = t[21396] ^ n[21397];
assign t[21398] = t[21397] ^ n[21398];
assign t[21399] = t[21398] ^ n[21399];
assign t[21400] = t[21399] ^ n[21400];
assign t[21401] = t[21400] ^ n[21401];
assign t[21402] = t[21401] ^ n[21402];
assign t[21403] = t[21402] ^ n[21403];
assign t[21404] = t[21403] ^ n[21404];
assign t[21405] = t[21404] ^ n[21405];
assign t[21406] = t[21405] ^ n[21406];
assign t[21407] = t[21406] ^ n[21407];
assign t[21408] = t[21407] ^ n[21408];
assign t[21409] = t[21408] ^ n[21409];
assign t[21410] = t[21409] ^ n[21410];
assign t[21411] = t[21410] ^ n[21411];
assign t[21412] = t[21411] ^ n[21412];
assign t[21413] = t[21412] ^ n[21413];
assign t[21414] = t[21413] ^ n[21414];
assign t[21415] = t[21414] ^ n[21415];
assign t[21416] = t[21415] ^ n[21416];
assign t[21417] = t[21416] ^ n[21417];
assign t[21418] = t[21417] ^ n[21418];
assign t[21419] = t[21418] ^ n[21419];
assign t[21420] = t[21419] ^ n[21420];
assign t[21421] = t[21420] ^ n[21421];
assign t[21422] = t[21421] ^ n[21422];
assign t[21423] = t[21422] ^ n[21423];
assign t[21424] = t[21423] ^ n[21424];
assign t[21425] = t[21424] ^ n[21425];
assign t[21426] = t[21425] ^ n[21426];
assign t[21427] = t[21426] ^ n[21427];
assign t[21428] = t[21427] ^ n[21428];
assign t[21429] = t[21428] ^ n[21429];
assign t[21430] = t[21429] ^ n[21430];
assign t[21431] = t[21430] ^ n[21431];
assign t[21432] = t[21431] ^ n[21432];
assign t[21433] = t[21432] ^ n[21433];
assign t[21434] = t[21433] ^ n[21434];
assign t[21435] = t[21434] ^ n[21435];
assign t[21436] = t[21435] ^ n[21436];
assign t[21437] = t[21436] ^ n[21437];
assign t[21438] = t[21437] ^ n[21438];
assign t[21439] = t[21438] ^ n[21439];
assign t[21440] = t[21439] ^ n[21440];
assign t[21441] = t[21440] ^ n[21441];
assign t[21442] = t[21441] ^ n[21442];
assign t[21443] = t[21442] ^ n[21443];
assign t[21444] = t[21443] ^ n[21444];
assign t[21445] = t[21444] ^ n[21445];
assign t[21446] = t[21445] ^ n[21446];
assign t[21447] = t[21446] ^ n[21447];
assign t[21448] = t[21447] ^ n[21448];
assign t[21449] = t[21448] ^ n[21449];
assign t[21450] = t[21449] ^ n[21450];
assign t[21451] = t[21450] ^ n[21451];
assign t[21452] = t[21451] ^ n[21452];
assign t[21453] = t[21452] ^ n[21453];
assign t[21454] = t[21453] ^ n[21454];
assign t[21455] = t[21454] ^ n[21455];
assign t[21456] = t[21455] ^ n[21456];
assign t[21457] = t[21456] ^ n[21457];
assign t[21458] = t[21457] ^ n[21458];
assign t[21459] = t[21458] ^ n[21459];
assign t[21460] = t[21459] ^ n[21460];
assign t[21461] = t[21460] ^ n[21461];
assign t[21462] = t[21461] ^ n[21462];
assign t[21463] = t[21462] ^ n[21463];
assign t[21464] = t[21463] ^ n[21464];
assign t[21465] = t[21464] ^ n[21465];
assign t[21466] = t[21465] ^ n[21466];
assign t[21467] = t[21466] ^ n[21467];
assign t[21468] = t[21467] ^ n[21468];
assign t[21469] = t[21468] ^ n[21469];
assign t[21470] = t[21469] ^ n[21470];
assign t[21471] = t[21470] ^ n[21471];
assign t[21472] = t[21471] ^ n[21472];
assign t[21473] = t[21472] ^ n[21473];
assign t[21474] = t[21473] ^ n[21474];
assign t[21475] = t[21474] ^ n[21475];
assign t[21476] = t[21475] ^ n[21476];
assign t[21477] = t[21476] ^ n[21477];
assign t[21478] = t[21477] ^ n[21478];
assign t[21479] = t[21478] ^ n[21479];
assign t[21480] = t[21479] ^ n[21480];
assign t[21481] = t[21480] ^ n[21481];
assign t[21482] = t[21481] ^ n[21482];
assign t[21483] = t[21482] ^ n[21483];
assign t[21484] = t[21483] ^ n[21484];
assign t[21485] = t[21484] ^ n[21485];
assign t[21486] = t[21485] ^ n[21486];
assign t[21487] = t[21486] ^ n[21487];
assign t[21488] = t[21487] ^ n[21488];
assign t[21489] = t[21488] ^ n[21489];
assign t[21490] = t[21489] ^ n[21490];
assign t[21491] = t[21490] ^ n[21491];
assign t[21492] = t[21491] ^ n[21492];
assign t[21493] = t[21492] ^ n[21493];
assign t[21494] = t[21493] ^ n[21494];
assign t[21495] = t[21494] ^ n[21495];
assign t[21496] = t[21495] ^ n[21496];
assign t[21497] = t[21496] ^ n[21497];
assign t[21498] = t[21497] ^ n[21498];
assign t[21499] = t[21498] ^ n[21499];
assign t[21500] = t[21499] ^ n[21500];
assign t[21501] = t[21500] ^ n[21501];
assign t[21502] = t[21501] ^ n[21502];
assign t[21503] = t[21502] ^ n[21503];
assign t[21504] = t[21503] ^ n[21504];
assign t[21505] = t[21504] ^ n[21505];
assign t[21506] = t[21505] ^ n[21506];
assign t[21507] = t[21506] ^ n[21507];
assign t[21508] = t[21507] ^ n[21508];
assign t[21509] = t[21508] ^ n[21509];
assign t[21510] = t[21509] ^ n[21510];
assign t[21511] = t[21510] ^ n[21511];
assign t[21512] = t[21511] ^ n[21512];
assign t[21513] = t[21512] ^ n[21513];
assign t[21514] = t[21513] ^ n[21514];
assign t[21515] = t[21514] ^ n[21515];
assign t[21516] = t[21515] ^ n[21516];
assign t[21517] = t[21516] ^ n[21517];
assign t[21518] = t[21517] ^ n[21518];
assign t[21519] = t[21518] ^ n[21519];
assign t[21520] = t[21519] ^ n[21520];
assign t[21521] = t[21520] ^ n[21521];
assign t[21522] = t[21521] ^ n[21522];
assign t[21523] = t[21522] ^ n[21523];
assign t[21524] = t[21523] ^ n[21524];
assign t[21525] = t[21524] ^ n[21525];
assign t[21526] = t[21525] ^ n[21526];
assign t[21527] = t[21526] ^ n[21527];
assign t[21528] = t[21527] ^ n[21528];
assign t[21529] = t[21528] ^ n[21529];
assign t[21530] = t[21529] ^ n[21530];
assign t[21531] = t[21530] ^ n[21531];
assign t[21532] = t[21531] ^ n[21532];
assign t[21533] = t[21532] ^ n[21533];
assign t[21534] = t[21533] ^ n[21534];
assign t[21535] = t[21534] ^ n[21535];
assign t[21536] = t[21535] ^ n[21536];
assign t[21537] = t[21536] ^ n[21537];
assign t[21538] = t[21537] ^ n[21538];
assign t[21539] = t[21538] ^ n[21539];
assign t[21540] = t[21539] ^ n[21540];
assign t[21541] = t[21540] ^ n[21541];
assign t[21542] = t[21541] ^ n[21542];
assign t[21543] = t[21542] ^ n[21543];
assign t[21544] = t[21543] ^ n[21544];
assign t[21545] = t[21544] ^ n[21545];
assign t[21546] = t[21545] ^ n[21546];
assign t[21547] = t[21546] ^ n[21547];
assign t[21548] = t[21547] ^ n[21548];
assign t[21549] = t[21548] ^ n[21549];
assign t[21550] = t[21549] ^ n[21550];
assign t[21551] = t[21550] ^ n[21551];
assign t[21552] = t[21551] ^ n[21552];
assign t[21553] = t[21552] ^ n[21553];
assign t[21554] = t[21553] ^ n[21554];
assign t[21555] = t[21554] ^ n[21555];
assign t[21556] = t[21555] ^ n[21556];
assign t[21557] = t[21556] ^ n[21557];
assign t[21558] = t[21557] ^ n[21558];
assign t[21559] = t[21558] ^ n[21559];
assign t[21560] = t[21559] ^ n[21560];
assign t[21561] = t[21560] ^ n[21561];
assign t[21562] = t[21561] ^ n[21562];
assign t[21563] = t[21562] ^ n[21563];
assign t[21564] = t[21563] ^ n[21564];
assign t[21565] = t[21564] ^ n[21565];
assign t[21566] = t[21565] ^ n[21566];
assign t[21567] = t[21566] ^ n[21567];
assign t[21568] = t[21567] ^ n[21568];
assign t[21569] = t[21568] ^ n[21569];
assign t[21570] = t[21569] ^ n[21570];
assign t[21571] = t[21570] ^ n[21571];
assign t[21572] = t[21571] ^ n[21572];
assign t[21573] = t[21572] ^ n[21573];
assign t[21574] = t[21573] ^ n[21574];
assign t[21575] = t[21574] ^ n[21575];
assign t[21576] = t[21575] ^ n[21576];
assign t[21577] = t[21576] ^ n[21577];
assign t[21578] = t[21577] ^ n[21578];
assign t[21579] = t[21578] ^ n[21579];
assign t[21580] = t[21579] ^ n[21580];
assign t[21581] = t[21580] ^ n[21581];
assign t[21582] = t[21581] ^ n[21582];
assign t[21583] = t[21582] ^ n[21583];
assign t[21584] = t[21583] ^ n[21584];
assign t[21585] = t[21584] ^ n[21585];
assign t[21586] = t[21585] ^ n[21586];
assign t[21587] = t[21586] ^ n[21587];
assign t[21588] = t[21587] ^ n[21588];
assign t[21589] = t[21588] ^ n[21589];
assign t[21590] = t[21589] ^ n[21590];
assign t[21591] = t[21590] ^ n[21591];
assign t[21592] = t[21591] ^ n[21592];
assign t[21593] = t[21592] ^ n[21593];
assign t[21594] = t[21593] ^ n[21594];
assign t[21595] = t[21594] ^ n[21595];
assign t[21596] = t[21595] ^ n[21596];
assign t[21597] = t[21596] ^ n[21597];
assign t[21598] = t[21597] ^ n[21598];
assign t[21599] = t[21598] ^ n[21599];
assign t[21600] = t[21599] ^ n[21600];
assign t[21601] = t[21600] ^ n[21601];
assign t[21602] = t[21601] ^ n[21602];
assign t[21603] = t[21602] ^ n[21603];
assign t[21604] = t[21603] ^ n[21604];
assign t[21605] = t[21604] ^ n[21605];
assign t[21606] = t[21605] ^ n[21606];
assign t[21607] = t[21606] ^ n[21607];
assign t[21608] = t[21607] ^ n[21608];
assign t[21609] = t[21608] ^ n[21609];
assign t[21610] = t[21609] ^ n[21610];
assign t[21611] = t[21610] ^ n[21611];
assign t[21612] = t[21611] ^ n[21612];
assign t[21613] = t[21612] ^ n[21613];
assign t[21614] = t[21613] ^ n[21614];
assign t[21615] = t[21614] ^ n[21615];
assign t[21616] = t[21615] ^ n[21616];
assign t[21617] = t[21616] ^ n[21617];
assign t[21618] = t[21617] ^ n[21618];
assign t[21619] = t[21618] ^ n[21619];
assign t[21620] = t[21619] ^ n[21620];
assign t[21621] = t[21620] ^ n[21621];
assign t[21622] = t[21621] ^ n[21622];
assign t[21623] = t[21622] ^ n[21623];
assign t[21624] = t[21623] ^ n[21624];
assign t[21625] = t[21624] ^ n[21625];
assign t[21626] = t[21625] ^ n[21626];
assign t[21627] = t[21626] ^ n[21627];
assign t[21628] = t[21627] ^ n[21628];
assign t[21629] = t[21628] ^ n[21629];
assign t[21630] = t[21629] ^ n[21630];
assign t[21631] = t[21630] ^ n[21631];
assign t[21632] = t[21631] ^ n[21632];
assign t[21633] = t[21632] ^ n[21633];
assign t[21634] = t[21633] ^ n[21634];
assign t[21635] = t[21634] ^ n[21635];
assign t[21636] = t[21635] ^ n[21636];
assign t[21637] = t[21636] ^ n[21637];
assign t[21638] = t[21637] ^ n[21638];
assign t[21639] = t[21638] ^ n[21639];
assign t[21640] = t[21639] ^ n[21640];
assign t[21641] = t[21640] ^ n[21641];
assign t[21642] = t[21641] ^ n[21642];
assign t[21643] = t[21642] ^ n[21643];
assign t[21644] = t[21643] ^ n[21644];
assign t[21645] = t[21644] ^ n[21645];
assign t[21646] = t[21645] ^ n[21646];
assign t[21647] = t[21646] ^ n[21647];
assign t[21648] = t[21647] ^ n[21648];
assign t[21649] = t[21648] ^ n[21649];
assign t[21650] = t[21649] ^ n[21650];
assign t[21651] = t[21650] ^ n[21651];
assign t[21652] = t[21651] ^ n[21652];
assign t[21653] = t[21652] ^ n[21653];
assign t[21654] = t[21653] ^ n[21654];
assign t[21655] = t[21654] ^ n[21655];
assign t[21656] = t[21655] ^ n[21656];
assign t[21657] = t[21656] ^ n[21657];
assign t[21658] = t[21657] ^ n[21658];
assign t[21659] = t[21658] ^ n[21659];
assign t[21660] = t[21659] ^ n[21660];
assign t[21661] = t[21660] ^ n[21661];
assign t[21662] = t[21661] ^ n[21662];
assign t[21663] = t[21662] ^ n[21663];
assign t[21664] = t[21663] ^ n[21664];
assign t[21665] = t[21664] ^ n[21665];
assign t[21666] = t[21665] ^ n[21666];
assign t[21667] = t[21666] ^ n[21667];
assign t[21668] = t[21667] ^ n[21668];
assign t[21669] = t[21668] ^ n[21669];
assign t[21670] = t[21669] ^ n[21670];
assign t[21671] = t[21670] ^ n[21671];
assign t[21672] = t[21671] ^ n[21672];
assign t[21673] = t[21672] ^ n[21673];
assign t[21674] = t[21673] ^ n[21674];
assign t[21675] = t[21674] ^ n[21675];
assign t[21676] = t[21675] ^ n[21676];
assign t[21677] = t[21676] ^ n[21677];
assign t[21678] = t[21677] ^ n[21678];
assign t[21679] = t[21678] ^ n[21679];
assign t[21680] = t[21679] ^ n[21680];
assign t[21681] = t[21680] ^ n[21681];
assign t[21682] = t[21681] ^ n[21682];
assign t[21683] = t[21682] ^ n[21683];
assign t[21684] = t[21683] ^ n[21684];
assign t[21685] = t[21684] ^ n[21685];
assign t[21686] = t[21685] ^ n[21686];
assign t[21687] = t[21686] ^ n[21687];
assign t[21688] = t[21687] ^ n[21688];
assign t[21689] = t[21688] ^ n[21689];
assign t[21690] = t[21689] ^ n[21690];
assign t[21691] = t[21690] ^ n[21691];
assign t[21692] = t[21691] ^ n[21692];
assign t[21693] = t[21692] ^ n[21693];
assign t[21694] = t[21693] ^ n[21694];
assign t[21695] = t[21694] ^ n[21695];
assign t[21696] = t[21695] ^ n[21696];
assign t[21697] = t[21696] ^ n[21697];
assign t[21698] = t[21697] ^ n[21698];
assign t[21699] = t[21698] ^ n[21699];
assign t[21700] = t[21699] ^ n[21700];
assign t[21701] = t[21700] ^ n[21701];
assign t[21702] = t[21701] ^ n[21702];
assign t[21703] = t[21702] ^ n[21703];
assign t[21704] = t[21703] ^ n[21704];
assign t[21705] = t[21704] ^ n[21705];
assign t[21706] = t[21705] ^ n[21706];
assign t[21707] = t[21706] ^ n[21707];
assign t[21708] = t[21707] ^ n[21708];
assign t[21709] = t[21708] ^ n[21709];
assign t[21710] = t[21709] ^ n[21710];
assign t[21711] = t[21710] ^ n[21711];
assign t[21712] = t[21711] ^ n[21712];
assign t[21713] = t[21712] ^ n[21713];
assign t[21714] = t[21713] ^ n[21714];
assign t[21715] = t[21714] ^ n[21715];
assign t[21716] = t[21715] ^ n[21716];
assign t[21717] = t[21716] ^ n[21717];
assign t[21718] = t[21717] ^ n[21718];
assign t[21719] = t[21718] ^ n[21719];
assign t[21720] = t[21719] ^ n[21720];
assign t[21721] = t[21720] ^ n[21721];
assign t[21722] = t[21721] ^ n[21722];
assign t[21723] = t[21722] ^ n[21723];
assign t[21724] = t[21723] ^ n[21724];
assign t[21725] = t[21724] ^ n[21725];
assign t[21726] = t[21725] ^ n[21726];
assign t[21727] = t[21726] ^ n[21727];
assign t[21728] = t[21727] ^ n[21728];
assign t[21729] = t[21728] ^ n[21729];
assign t[21730] = t[21729] ^ n[21730];
assign t[21731] = t[21730] ^ n[21731];
assign t[21732] = t[21731] ^ n[21732];
assign t[21733] = t[21732] ^ n[21733];
assign t[21734] = t[21733] ^ n[21734];
assign t[21735] = t[21734] ^ n[21735];
assign t[21736] = t[21735] ^ n[21736];
assign t[21737] = t[21736] ^ n[21737];
assign t[21738] = t[21737] ^ n[21738];
assign t[21739] = t[21738] ^ n[21739];
assign t[21740] = t[21739] ^ n[21740];
assign t[21741] = t[21740] ^ n[21741];
assign t[21742] = t[21741] ^ n[21742];
assign t[21743] = t[21742] ^ n[21743];
assign t[21744] = t[21743] ^ n[21744];
assign t[21745] = t[21744] ^ n[21745];
assign t[21746] = t[21745] ^ n[21746];
assign t[21747] = t[21746] ^ n[21747];
assign t[21748] = t[21747] ^ n[21748];
assign t[21749] = t[21748] ^ n[21749];
assign t[21750] = t[21749] ^ n[21750];
assign t[21751] = t[21750] ^ n[21751];
assign t[21752] = t[21751] ^ n[21752];
assign t[21753] = t[21752] ^ n[21753];
assign t[21754] = t[21753] ^ n[21754];
assign t[21755] = t[21754] ^ n[21755];
assign t[21756] = t[21755] ^ n[21756];
assign t[21757] = t[21756] ^ n[21757];
assign t[21758] = t[21757] ^ n[21758];
assign t[21759] = t[21758] ^ n[21759];
assign t[21760] = t[21759] ^ n[21760];
assign t[21761] = t[21760] ^ n[21761];
assign t[21762] = t[21761] ^ n[21762];
assign t[21763] = t[21762] ^ n[21763];
assign t[21764] = t[21763] ^ n[21764];
assign t[21765] = t[21764] ^ n[21765];
assign t[21766] = t[21765] ^ n[21766];
assign t[21767] = t[21766] ^ n[21767];
assign t[21768] = t[21767] ^ n[21768];
assign t[21769] = t[21768] ^ n[21769];
assign t[21770] = t[21769] ^ n[21770];
assign t[21771] = t[21770] ^ n[21771];
assign t[21772] = t[21771] ^ n[21772];
assign t[21773] = t[21772] ^ n[21773];
assign t[21774] = t[21773] ^ n[21774];
assign t[21775] = t[21774] ^ n[21775];
assign t[21776] = t[21775] ^ n[21776];
assign t[21777] = t[21776] ^ n[21777];
assign t[21778] = t[21777] ^ n[21778];
assign t[21779] = t[21778] ^ n[21779];
assign t[21780] = t[21779] ^ n[21780];
assign t[21781] = t[21780] ^ n[21781];
assign t[21782] = t[21781] ^ n[21782];
assign t[21783] = t[21782] ^ n[21783];
assign t[21784] = t[21783] ^ n[21784];
assign t[21785] = t[21784] ^ n[21785];
assign t[21786] = t[21785] ^ n[21786];
assign t[21787] = t[21786] ^ n[21787];
assign t[21788] = t[21787] ^ n[21788];
assign t[21789] = t[21788] ^ n[21789];
assign t[21790] = t[21789] ^ n[21790];
assign t[21791] = t[21790] ^ n[21791];
assign t[21792] = t[21791] ^ n[21792];
assign t[21793] = t[21792] ^ n[21793];
assign t[21794] = t[21793] ^ n[21794];
assign t[21795] = t[21794] ^ n[21795];
assign t[21796] = t[21795] ^ n[21796];
assign t[21797] = t[21796] ^ n[21797];
assign t[21798] = t[21797] ^ n[21798];
assign t[21799] = t[21798] ^ n[21799];
assign t[21800] = t[21799] ^ n[21800];
assign t[21801] = t[21800] ^ n[21801];
assign t[21802] = t[21801] ^ n[21802];
assign t[21803] = t[21802] ^ n[21803];
assign t[21804] = t[21803] ^ n[21804];
assign t[21805] = t[21804] ^ n[21805];
assign t[21806] = t[21805] ^ n[21806];
assign t[21807] = t[21806] ^ n[21807];
assign t[21808] = t[21807] ^ n[21808];
assign t[21809] = t[21808] ^ n[21809];
assign t[21810] = t[21809] ^ n[21810];
assign t[21811] = t[21810] ^ n[21811];
assign t[21812] = t[21811] ^ n[21812];
assign t[21813] = t[21812] ^ n[21813];
assign t[21814] = t[21813] ^ n[21814];
assign t[21815] = t[21814] ^ n[21815];
assign t[21816] = t[21815] ^ n[21816];
assign t[21817] = t[21816] ^ n[21817];
assign t[21818] = t[21817] ^ n[21818];
assign t[21819] = t[21818] ^ n[21819];
assign t[21820] = t[21819] ^ n[21820];
assign t[21821] = t[21820] ^ n[21821];
assign t[21822] = t[21821] ^ n[21822];
assign t[21823] = t[21822] ^ n[21823];
assign t[21824] = t[21823] ^ n[21824];
assign t[21825] = t[21824] ^ n[21825];
assign t[21826] = t[21825] ^ n[21826];
assign t[21827] = t[21826] ^ n[21827];
assign t[21828] = t[21827] ^ n[21828];
assign t[21829] = t[21828] ^ n[21829];
assign t[21830] = t[21829] ^ n[21830];
assign t[21831] = t[21830] ^ n[21831];
assign t[21832] = t[21831] ^ n[21832];
assign t[21833] = t[21832] ^ n[21833];
assign t[21834] = t[21833] ^ n[21834];
assign t[21835] = t[21834] ^ n[21835];
assign t[21836] = t[21835] ^ n[21836];
assign t[21837] = t[21836] ^ n[21837];
assign t[21838] = t[21837] ^ n[21838];
assign t[21839] = t[21838] ^ n[21839];
assign t[21840] = t[21839] ^ n[21840];
assign t[21841] = t[21840] ^ n[21841];
assign t[21842] = t[21841] ^ n[21842];
assign t[21843] = t[21842] ^ n[21843];
assign t[21844] = t[21843] ^ n[21844];
assign t[21845] = t[21844] ^ n[21845];
assign t[21846] = t[21845] ^ n[21846];
assign t[21847] = t[21846] ^ n[21847];
assign t[21848] = t[21847] ^ n[21848];
assign t[21849] = t[21848] ^ n[21849];
assign t[21850] = t[21849] ^ n[21850];
assign t[21851] = t[21850] ^ n[21851];
assign t[21852] = t[21851] ^ n[21852];
assign t[21853] = t[21852] ^ n[21853];
assign t[21854] = t[21853] ^ n[21854];
assign t[21855] = t[21854] ^ n[21855];
assign t[21856] = t[21855] ^ n[21856];
assign t[21857] = t[21856] ^ n[21857];
assign t[21858] = t[21857] ^ n[21858];
assign t[21859] = t[21858] ^ n[21859];
assign t[21860] = t[21859] ^ n[21860];
assign t[21861] = t[21860] ^ n[21861];
assign t[21862] = t[21861] ^ n[21862];
assign t[21863] = t[21862] ^ n[21863];
assign t[21864] = t[21863] ^ n[21864];
assign t[21865] = t[21864] ^ n[21865];
assign t[21866] = t[21865] ^ n[21866];
assign t[21867] = t[21866] ^ n[21867];
assign t[21868] = t[21867] ^ n[21868];
assign t[21869] = t[21868] ^ n[21869];
assign t[21870] = t[21869] ^ n[21870];
assign t[21871] = t[21870] ^ n[21871];
assign t[21872] = t[21871] ^ n[21872];
assign t[21873] = t[21872] ^ n[21873];
assign t[21874] = t[21873] ^ n[21874];
assign t[21875] = t[21874] ^ n[21875];
assign t[21876] = t[21875] ^ n[21876];
assign t[21877] = t[21876] ^ n[21877];
assign t[21878] = t[21877] ^ n[21878];
assign t[21879] = t[21878] ^ n[21879];
assign t[21880] = t[21879] ^ n[21880];
assign t[21881] = t[21880] ^ n[21881];
assign t[21882] = t[21881] ^ n[21882];
assign t[21883] = t[21882] ^ n[21883];
assign t[21884] = t[21883] ^ n[21884];
assign t[21885] = t[21884] ^ n[21885];
assign t[21886] = t[21885] ^ n[21886];
assign t[21887] = t[21886] ^ n[21887];
assign t[21888] = t[21887] ^ n[21888];
assign t[21889] = t[21888] ^ n[21889];
assign t[21890] = t[21889] ^ n[21890];
assign t[21891] = t[21890] ^ n[21891];
assign t[21892] = t[21891] ^ n[21892];
assign t[21893] = t[21892] ^ n[21893];
assign t[21894] = t[21893] ^ n[21894];
assign t[21895] = t[21894] ^ n[21895];
assign t[21896] = t[21895] ^ n[21896];
assign t[21897] = t[21896] ^ n[21897];
assign t[21898] = t[21897] ^ n[21898];
assign t[21899] = t[21898] ^ n[21899];
assign t[21900] = t[21899] ^ n[21900];
assign t[21901] = t[21900] ^ n[21901];
assign t[21902] = t[21901] ^ n[21902];
assign t[21903] = t[21902] ^ n[21903];
assign t[21904] = t[21903] ^ n[21904];
assign t[21905] = t[21904] ^ n[21905];
assign t[21906] = t[21905] ^ n[21906];
assign t[21907] = t[21906] ^ n[21907];
assign t[21908] = t[21907] ^ n[21908];
assign t[21909] = t[21908] ^ n[21909];
assign t[21910] = t[21909] ^ n[21910];
assign t[21911] = t[21910] ^ n[21911];
assign t[21912] = t[21911] ^ n[21912];
assign t[21913] = t[21912] ^ n[21913];
assign t[21914] = t[21913] ^ n[21914];
assign t[21915] = t[21914] ^ n[21915];
assign t[21916] = t[21915] ^ n[21916];
assign t[21917] = t[21916] ^ n[21917];
assign t[21918] = t[21917] ^ n[21918];
assign t[21919] = t[21918] ^ n[21919];
assign t[21920] = t[21919] ^ n[21920];
assign t[21921] = t[21920] ^ n[21921];
assign t[21922] = t[21921] ^ n[21922];
assign t[21923] = t[21922] ^ n[21923];
assign t[21924] = t[21923] ^ n[21924];
assign t[21925] = t[21924] ^ n[21925];
assign t[21926] = t[21925] ^ n[21926];
assign t[21927] = t[21926] ^ n[21927];
assign t[21928] = t[21927] ^ n[21928];
assign t[21929] = t[21928] ^ n[21929];
assign t[21930] = t[21929] ^ n[21930];
assign t[21931] = t[21930] ^ n[21931];
assign t[21932] = t[21931] ^ n[21932];
assign t[21933] = t[21932] ^ n[21933];
assign t[21934] = t[21933] ^ n[21934];
assign t[21935] = t[21934] ^ n[21935];
assign t[21936] = t[21935] ^ n[21936];
assign t[21937] = t[21936] ^ n[21937];
assign t[21938] = t[21937] ^ n[21938];
assign t[21939] = t[21938] ^ n[21939];
assign t[21940] = t[21939] ^ n[21940];
assign t[21941] = t[21940] ^ n[21941];
assign t[21942] = t[21941] ^ n[21942];
assign t[21943] = t[21942] ^ n[21943];
assign t[21944] = t[21943] ^ n[21944];
assign t[21945] = t[21944] ^ n[21945];
assign t[21946] = t[21945] ^ n[21946];
assign t[21947] = t[21946] ^ n[21947];
assign t[21948] = t[21947] ^ n[21948];
assign t[21949] = t[21948] ^ n[21949];
assign t[21950] = t[21949] ^ n[21950];
assign t[21951] = t[21950] ^ n[21951];
assign t[21952] = t[21951] ^ n[21952];
assign t[21953] = t[21952] ^ n[21953];
assign t[21954] = t[21953] ^ n[21954];
assign t[21955] = t[21954] ^ n[21955];
assign t[21956] = t[21955] ^ n[21956];
assign t[21957] = t[21956] ^ n[21957];
assign t[21958] = t[21957] ^ n[21958];
assign t[21959] = t[21958] ^ n[21959];
assign t[21960] = t[21959] ^ n[21960];
assign t[21961] = t[21960] ^ n[21961];
assign t[21962] = t[21961] ^ n[21962];
assign t[21963] = t[21962] ^ n[21963];
assign t[21964] = t[21963] ^ n[21964];
assign t[21965] = t[21964] ^ n[21965];
assign t[21966] = t[21965] ^ n[21966];
assign t[21967] = t[21966] ^ n[21967];
assign t[21968] = t[21967] ^ n[21968];
assign t[21969] = t[21968] ^ n[21969];
assign t[21970] = t[21969] ^ n[21970];
assign t[21971] = t[21970] ^ n[21971];
assign t[21972] = t[21971] ^ n[21972];
assign t[21973] = t[21972] ^ n[21973];
assign t[21974] = t[21973] ^ n[21974];
assign t[21975] = t[21974] ^ n[21975];
assign t[21976] = t[21975] ^ n[21976];
assign t[21977] = t[21976] ^ n[21977];
assign t[21978] = t[21977] ^ n[21978];
assign t[21979] = t[21978] ^ n[21979];
assign t[21980] = t[21979] ^ n[21980];
assign t[21981] = t[21980] ^ n[21981];
assign t[21982] = t[21981] ^ n[21982];
assign t[21983] = t[21982] ^ n[21983];
assign t[21984] = t[21983] ^ n[21984];
assign t[21985] = t[21984] ^ n[21985];
assign t[21986] = t[21985] ^ n[21986];
assign t[21987] = t[21986] ^ n[21987];
assign t[21988] = t[21987] ^ n[21988];
assign t[21989] = t[21988] ^ n[21989];
assign t[21990] = t[21989] ^ n[21990];
assign t[21991] = t[21990] ^ n[21991];
assign t[21992] = t[21991] ^ n[21992];
assign t[21993] = t[21992] ^ n[21993];
assign t[21994] = t[21993] ^ n[21994];
assign t[21995] = t[21994] ^ n[21995];
assign t[21996] = t[21995] ^ n[21996];
assign t[21997] = t[21996] ^ n[21997];
assign t[21998] = t[21997] ^ n[21998];
assign t[21999] = t[21998] ^ n[21999];
assign t[22000] = t[21999] ^ n[22000];
assign t[22001] = t[22000] ^ n[22001];
assign t[22002] = t[22001] ^ n[22002];
assign t[22003] = t[22002] ^ n[22003];
assign t[22004] = t[22003] ^ n[22004];
assign t[22005] = t[22004] ^ n[22005];
assign t[22006] = t[22005] ^ n[22006];
assign t[22007] = t[22006] ^ n[22007];
assign t[22008] = t[22007] ^ n[22008];
assign t[22009] = t[22008] ^ n[22009];
assign t[22010] = t[22009] ^ n[22010];
assign t[22011] = t[22010] ^ n[22011];
assign t[22012] = t[22011] ^ n[22012];
assign t[22013] = t[22012] ^ n[22013];
assign t[22014] = t[22013] ^ n[22014];
assign t[22015] = t[22014] ^ n[22015];
assign t[22016] = t[22015] ^ n[22016];
assign t[22017] = t[22016] ^ n[22017];
assign t[22018] = t[22017] ^ n[22018];
assign t[22019] = t[22018] ^ n[22019];
assign t[22020] = t[22019] ^ n[22020];
assign t[22021] = t[22020] ^ n[22021];
assign t[22022] = t[22021] ^ n[22022];
assign t[22023] = t[22022] ^ n[22023];
assign t[22024] = t[22023] ^ n[22024];
assign t[22025] = t[22024] ^ n[22025];
assign t[22026] = t[22025] ^ n[22026];
assign t[22027] = t[22026] ^ n[22027];
assign t[22028] = t[22027] ^ n[22028];
assign t[22029] = t[22028] ^ n[22029];
assign t[22030] = t[22029] ^ n[22030];
assign t[22031] = t[22030] ^ n[22031];
assign t[22032] = t[22031] ^ n[22032];
assign t[22033] = t[22032] ^ n[22033];
assign t[22034] = t[22033] ^ n[22034];
assign t[22035] = t[22034] ^ n[22035];
assign t[22036] = t[22035] ^ n[22036];
assign t[22037] = t[22036] ^ n[22037];
assign t[22038] = t[22037] ^ n[22038];
assign t[22039] = t[22038] ^ n[22039];
assign t[22040] = t[22039] ^ n[22040];
assign t[22041] = t[22040] ^ n[22041];
assign t[22042] = t[22041] ^ n[22042];
assign t[22043] = t[22042] ^ n[22043];
assign t[22044] = t[22043] ^ n[22044];
assign t[22045] = t[22044] ^ n[22045];
assign t[22046] = t[22045] ^ n[22046];
assign t[22047] = t[22046] ^ n[22047];
assign t[22048] = t[22047] ^ n[22048];
assign t[22049] = t[22048] ^ n[22049];
assign t[22050] = t[22049] ^ n[22050];
assign t[22051] = t[22050] ^ n[22051];
assign t[22052] = t[22051] ^ n[22052];
assign t[22053] = t[22052] ^ n[22053];
assign t[22054] = t[22053] ^ n[22054];
assign t[22055] = t[22054] ^ n[22055];
assign t[22056] = t[22055] ^ n[22056];
assign t[22057] = t[22056] ^ n[22057];
assign t[22058] = t[22057] ^ n[22058];
assign t[22059] = t[22058] ^ n[22059];
assign t[22060] = t[22059] ^ n[22060];
assign t[22061] = t[22060] ^ n[22061];
assign t[22062] = t[22061] ^ n[22062];
assign t[22063] = t[22062] ^ n[22063];
assign t[22064] = t[22063] ^ n[22064];
assign t[22065] = t[22064] ^ n[22065];
assign t[22066] = t[22065] ^ n[22066];
assign t[22067] = t[22066] ^ n[22067];
assign t[22068] = t[22067] ^ n[22068];
assign t[22069] = t[22068] ^ n[22069];
assign t[22070] = t[22069] ^ n[22070];
assign t[22071] = t[22070] ^ n[22071];
assign t[22072] = t[22071] ^ n[22072];
assign t[22073] = t[22072] ^ n[22073];
assign t[22074] = t[22073] ^ n[22074];
assign t[22075] = t[22074] ^ n[22075];
assign t[22076] = t[22075] ^ n[22076];
assign t[22077] = t[22076] ^ n[22077];
assign t[22078] = t[22077] ^ n[22078];
assign t[22079] = t[22078] ^ n[22079];
assign t[22080] = t[22079] ^ n[22080];
assign t[22081] = t[22080] ^ n[22081];
assign t[22082] = t[22081] ^ n[22082];
assign t[22083] = t[22082] ^ n[22083];
assign t[22084] = t[22083] ^ n[22084];
assign t[22085] = t[22084] ^ n[22085];
assign t[22086] = t[22085] ^ n[22086];
assign t[22087] = t[22086] ^ n[22087];
assign t[22088] = t[22087] ^ n[22088];
assign t[22089] = t[22088] ^ n[22089];
assign t[22090] = t[22089] ^ n[22090];
assign t[22091] = t[22090] ^ n[22091];
assign t[22092] = t[22091] ^ n[22092];
assign t[22093] = t[22092] ^ n[22093];
assign t[22094] = t[22093] ^ n[22094];
assign t[22095] = t[22094] ^ n[22095];
assign t[22096] = t[22095] ^ n[22096];
assign t[22097] = t[22096] ^ n[22097];
assign t[22098] = t[22097] ^ n[22098];
assign t[22099] = t[22098] ^ n[22099];
assign t[22100] = t[22099] ^ n[22100];
assign t[22101] = t[22100] ^ n[22101];
assign t[22102] = t[22101] ^ n[22102];
assign t[22103] = t[22102] ^ n[22103];
assign t[22104] = t[22103] ^ n[22104];
assign t[22105] = t[22104] ^ n[22105];
assign t[22106] = t[22105] ^ n[22106];
assign t[22107] = t[22106] ^ n[22107];
assign t[22108] = t[22107] ^ n[22108];
assign t[22109] = t[22108] ^ n[22109];
assign t[22110] = t[22109] ^ n[22110];
assign t[22111] = t[22110] ^ n[22111];
assign t[22112] = t[22111] ^ n[22112];
assign t[22113] = t[22112] ^ n[22113];
assign t[22114] = t[22113] ^ n[22114];
assign t[22115] = t[22114] ^ n[22115];
assign t[22116] = t[22115] ^ n[22116];
assign t[22117] = t[22116] ^ n[22117];
assign t[22118] = t[22117] ^ n[22118];
assign t[22119] = t[22118] ^ n[22119];
assign t[22120] = t[22119] ^ n[22120];
assign t[22121] = t[22120] ^ n[22121];
assign t[22122] = t[22121] ^ n[22122];
assign t[22123] = t[22122] ^ n[22123];
assign t[22124] = t[22123] ^ n[22124];
assign t[22125] = t[22124] ^ n[22125];
assign t[22126] = t[22125] ^ n[22126];
assign t[22127] = t[22126] ^ n[22127];
assign t[22128] = t[22127] ^ n[22128];
assign t[22129] = t[22128] ^ n[22129];
assign t[22130] = t[22129] ^ n[22130];
assign t[22131] = t[22130] ^ n[22131];
assign t[22132] = t[22131] ^ n[22132];
assign t[22133] = t[22132] ^ n[22133];
assign t[22134] = t[22133] ^ n[22134];
assign t[22135] = t[22134] ^ n[22135];
assign t[22136] = t[22135] ^ n[22136];
assign t[22137] = t[22136] ^ n[22137];
assign t[22138] = t[22137] ^ n[22138];
assign t[22139] = t[22138] ^ n[22139];
assign t[22140] = t[22139] ^ n[22140];
assign t[22141] = t[22140] ^ n[22141];
assign t[22142] = t[22141] ^ n[22142];
assign t[22143] = t[22142] ^ n[22143];
assign t[22144] = t[22143] ^ n[22144];
assign t[22145] = t[22144] ^ n[22145];
assign t[22146] = t[22145] ^ n[22146];
assign t[22147] = t[22146] ^ n[22147];
assign t[22148] = t[22147] ^ n[22148];
assign t[22149] = t[22148] ^ n[22149];
assign t[22150] = t[22149] ^ n[22150];
assign t[22151] = t[22150] ^ n[22151];
assign t[22152] = t[22151] ^ n[22152];
assign t[22153] = t[22152] ^ n[22153];
assign t[22154] = t[22153] ^ n[22154];
assign t[22155] = t[22154] ^ n[22155];
assign t[22156] = t[22155] ^ n[22156];
assign t[22157] = t[22156] ^ n[22157];
assign t[22158] = t[22157] ^ n[22158];
assign t[22159] = t[22158] ^ n[22159];
assign t[22160] = t[22159] ^ n[22160];
assign t[22161] = t[22160] ^ n[22161];
assign t[22162] = t[22161] ^ n[22162];
assign t[22163] = t[22162] ^ n[22163];
assign t[22164] = t[22163] ^ n[22164];
assign t[22165] = t[22164] ^ n[22165];
assign t[22166] = t[22165] ^ n[22166];
assign t[22167] = t[22166] ^ n[22167];
assign t[22168] = t[22167] ^ n[22168];
assign t[22169] = t[22168] ^ n[22169];
assign t[22170] = t[22169] ^ n[22170];
assign t[22171] = t[22170] ^ n[22171];
assign t[22172] = t[22171] ^ n[22172];
assign t[22173] = t[22172] ^ n[22173];
assign t[22174] = t[22173] ^ n[22174];
assign t[22175] = t[22174] ^ n[22175];
assign t[22176] = t[22175] ^ n[22176];
assign t[22177] = t[22176] ^ n[22177];
assign t[22178] = t[22177] ^ n[22178];
assign t[22179] = t[22178] ^ n[22179];
assign t[22180] = t[22179] ^ n[22180];
assign t[22181] = t[22180] ^ n[22181];
assign t[22182] = t[22181] ^ n[22182];
assign t[22183] = t[22182] ^ n[22183];
assign t[22184] = t[22183] ^ n[22184];
assign t[22185] = t[22184] ^ n[22185];
assign t[22186] = t[22185] ^ n[22186];
assign t[22187] = t[22186] ^ n[22187];
assign t[22188] = t[22187] ^ n[22188];
assign t[22189] = t[22188] ^ n[22189];
assign t[22190] = t[22189] ^ n[22190];
assign t[22191] = t[22190] ^ n[22191];
assign t[22192] = t[22191] ^ n[22192];
assign t[22193] = t[22192] ^ n[22193];
assign t[22194] = t[22193] ^ n[22194];
assign t[22195] = t[22194] ^ n[22195];
assign t[22196] = t[22195] ^ n[22196];
assign t[22197] = t[22196] ^ n[22197];
assign t[22198] = t[22197] ^ n[22198];
assign t[22199] = t[22198] ^ n[22199];
assign t[22200] = t[22199] ^ n[22200];
assign t[22201] = t[22200] ^ n[22201];
assign t[22202] = t[22201] ^ n[22202];
assign t[22203] = t[22202] ^ n[22203];
assign t[22204] = t[22203] ^ n[22204];
assign t[22205] = t[22204] ^ n[22205];
assign t[22206] = t[22205] ^ n[22206];
assign t[22207] = t[22206] ^ n[22207];
assign t[22208] = t[22207] ^ n[22208];
assign t[22209] = t[22208] ^ n[22209];
assign t[22210] = t[22209] ^ n[22210];
assign t[22211] = t[22210] ^ n[22211];
assign t[22212] = t[22211] ^ n[22212];
assign t[22213] = t[22212] ^ n[22213];
assign t[22214] = t[22213] ^ n[22214];
assign t[22215] = t[22214] ^ n[22215];
assign t[22216] = t[22215] ^ n[22216];
assign t[22217] = t[22216] ^ n[22217];
assign t[22218] = t[22217] ^ n[22218];
assign t[22219] = t[22218] ^ n[22219];
assign t[22220] = t[22219] ^ n[22220];
assign t[22221] = t[22220] ^ n[22221];
assign t[22222] = t[22221] ^ n[22222];
assign t[22223] = t[22222] ^ n[22223];
assign t[22224] = t[22223] ^ n[22224];
assign t[22225] = t[22224] ^ n[22225];
assign t[22226] = t[22225] ^ n[22226];
assign t[22227] = t[22226] ^ n[22227];
assign t[22228] = t[22227] ^ n[22228];
assign t[22229] = t[22228] ^ n[22229];
assign t[22230] = t[22229] ^ n[22230];
assign t[22231] = t[22230] ^ n[22231];
assign t[22232] = t[22231] ^ n[22232];
assign t[22233] = t[22232] ^ n[22233];
assign t[22234] = t[22233] ^ n[22234];
assign t[22235] = t[22234] ^ n[22235];
assign t[22236] = t[22235] ^ n[22236];
assign t[22237] = t[22236] ^ n[22237];
assign t[22238] = t[22237] ^ n[22238];
assign t[22239] = t[22238] ^ n[22239];
assign t[22240] = t[22239] ^ n[22240];
assign t[22241] = t[22240] ^ n[22241];
assign t[22242] = t[22241] ^ n[22242];
assign t[22243] = t[22242] ^ n[22243];
assign t[22244] = t[22243] ^ n[22244];
assign t[22245] = t[22244] ^ n[22245];
assign t[22246] = t[22245] ^ n[22246];
assign t[22247] = t[22246] ^ n[22247];
assign t[22248] = t[22247] ^ n[22248];
assign t[22249] = t[22248] ^ n[22249];
assign t[22250] = t[22249] ^ n[22250];
assign t[22251] = t[22250] ^ n[22251];
assign t[22252] = t[22251] ^ n[22252];
assign t[22253] = t[22252] ^ n[22253];
assign t[22254] = t[22253] ^ n[22254];
assign t[22255] = t[22254] ^ n[22255];
assign t[22256] = t[22255] ^ n[22256];
assign t[22257] = t[22256] ^ n[22257];
assign t[22258] = t[22257] ^ n[22258];
assign t[22259] = t[22258] ^ n[22259];
assign t[22260] = t[22259] ^ n[22260];
assign t[22261] = t[22260] ^ n[22261];
assign t[22262] = t[22261] ^ n[22262];
assign t[22263] = t[22262] ^ n[22263];
assign t[22264] = t[22263] ^ n[22264];
assign t[22265] = t[22264] ^ n[22265];
assign t[22266] = t[22265] ^ n[22266];
assign t[22267] = t[22266] ^ n[22267];
assign t[22268] = t[22267] ^ n[22268];
assign t[22269] = t[22268] ^ n[22269];
assign t[22270] = t[22269] ^ n[22270];
assign t[22271] = t[22270] ^ n[22271];
assign t[22272] = t[22271] ^ n[22272];
assign t[22273] = t[22272] ^ n[22273];
assign t[22274] = t[22273] ^ n[22274];
assign t[22275] = t[22274] ^ n[22275];
assign t[22276] = t[22275] ^ n[22276];
assign t[22277] = t[22276] ^ n[22277];
assign t[22278] = t[22277] ^ n[22278];
assign t[22279] = t[22278] ^ n[22279];
assign t[22280] = t[22279] ^ n[22280];
assign t[22281] = t[22280] ^ n[22281];
assign t[22282] = t[22281] ^ n[22282];
assign t[22283] = t[22282] ^ n[22283];
assign t[22284] = t[22283] ^ n[22284];
assign t[22285] = t[22284] ^ n[22285];
assign t[22286] = t[22285] ^ n[22286];
assign t[22287] = t[22286] ^ n[22287];
assign t[22288] = t[22287] ^ n[22288];
assign t[22289] = t[22288] ^ n[22289];
assign t[22290] = t[22289] ^ n[22290];
assign t[22291] = t[22290] ^ n[22291];
assign t[22292] = t[22291] ^ n[22292];
assign t[22293] = t[22292] ^ n[22293];
assign t[22294] = t[22293] ^ n[22294];
assign t[22295] = t[22294] ^ n[22295];
assign t[22296] = t[22295] ^ n[22296];
assign t[22297] = t[22296] ^ n[22297];
assign t[22298] = t[22297] ^ n[22298];
assign t[22299] = t[22298] ^ n[22299];
assign t[22300] = t[22299] ^ n[22300];
assign t[22301] = t[22300] ^ n[22301];
assign t[22302] = t[22301] ^ n[22302];
assign t[22303] = t[22302] ^ n[22303];
assign t[22304] = t[22303] ^ n[22304];
assign t[22305] = t[22304] ^ n[22305];
assign t[22306] = t[22305] ^ n[22306];
assign t[22307] = t[22306] ^ n[22307];
assign t[22308] = t[22307] ^ n[22308];
assign t[22309] = t[22308] ^ n[22309];
assign t[22310] = t[22309] ^ n[22310];
assign t[22311] = t[22310] ^ n[22311];
assign t[22312] = t[22311] ^ n[22312];
assign t[22313] = t[22312] ^ n[22313];
assign t[22314] = t[22313] ^ n[22314];
assign t[22315] = t[22314] ^ n[22315];
assign t[22316] = t[22315] ^ n[22316];
assign t[22317] = t[22316] ^ n[22317];
assign t[22318] = t[22317] ^ n[22318];
assign t[22319] = t[22318] ^ n[22319];
assign t[22320] = t[22319] ^ n[22320];
assign t[22321] = t[22320] ^ n[22321];
assign t[22322] = t[22321] ^ n[22322];
assign t[22323] = t[22322] ^ n[22323];
assign t[22324] = t[22323] ^ n[22324];
assign t[22325] = t[22324] ^ n[22325];
assign t[22326] = t[22325] ^ n[22326];
assign t[22327] = t[22326] ^ n[22327];
assign t[22328] = t[22327] ^ n[22328];
assign t[22329] = t[22328] ^ n[22329];
assign t[22330] = t[22329] ^ n[22330];
assign t[22331] = t[22330] ^ n[22331];
assign t[22332] = t[22331] ^ n[22332];
assign t[22333] = t[22332] ^ n[22333];
assign t[22334] = t[22333] ^ n[22334];
assign t[22335] = t[22334] ^ n[22335];
assign t[22336] = t[22335] ^ n[22336];
assign t[22337] = t[22336] ^ n[22337];
assign t[22338] = t[22337] ^ n[22338];
assign t[22339] = t[22338] ^ n[22339];
assign t[22340] = t[22339] ^ n[22340];
assign t[22341] = t[22340] ^ n[22341];
assign t[22342] = t[22341] ^ n[22342];
assign t[22343] = t[22342] ^ n[22343];
assign t[22344] = t[22343] ^ n[22344];
assign t[22345] = t[22344] ^ n[22345];
assign t[22346] = t[22345] ^ n[22346];
assign t[22347] = t[22346] ^ n[22347];
assign t[22348] = t[22347] ^ n[22348];
assign t[22349] = t[22348] ^ n[22349];
assign t[22350] = t[22349] ^ n[22350];
assign t[22351] = t[22350] ^ n[22351];
assign t[22352] = t[22351] ^ n[22352];
assign t[22353] = t[22352] ^ n[22353];
assign t[22354] = t[22353] ^ n[22354];
assign t[22355] = t[22354] ^ n[22355];
assign t[22356] = t[22355] ^ n[22356];
assign t[22357] = t[22356] ^ n[22357];
assign t[22358] = t[22357] ^ n[22358];
assign t[22359] = t[22358] ^ n[22359];
assign t[22360] = t[22359] ^ n[22360];
assign t[22361] = t[22360] ^ n[22361];
assign t[22362] = t[22361] ^ n[22362];
assign t[22363] = t[22362] ^ n[22363];
assign t[22364] = t[22363] ^ n[22364];
assign t[22365] = t[22364] ^ n[22365];
assign t[22366] = t[22365] ^ n[22366];
assign t[22367] = t[22366] ^ n[22367];
assign t[22368] = t[22367] ^ n[22368];
assign t[22369] = t[22368] ^ n[22369];
assign t[22370] = t[22369] ^ n[22370];
assign t[22371] = t[22370] ^ n[22371];
assign t[22372] = t[22371] ^ n[22372];
assign t[22373] = t[22372] ^ n[22373];
assign t[22374] = t[22373] ^ n[22374];
assign t[22375] = t[22374] ^ n[22375];
assign t[22376] = t[22375] ^ n[22376];
assign t[22377] = t[22376] ^ n[22377];
assign t[22378] = t[22377] ^ n[22378];
assign t[22379] = t[22378] ^ n[22379];
assign t[22380] = t[22379] ^ n[22380];
assign t[22381] = t[22380] ^ n[22381];
assign t[22382] = t[22381] ^ n[22382];
assign t[22383] = t[22382] ^ n[22383];
assign t[22384] = t[22383] ^ n[22384];
assign t[22385] = t[22384] ^ n[22385];
assign t[22386] = t[22385] ^ n[22386];
assign t[22387] = t[22386] ^ n[22387];
assign t[22388] = t[22387] ^ n[22388];
assign t[22389] = t[22388] ^ n[22389];
assign t[22390] = t[22389] ^ n[22390];
assign t[22391] = t[22390] ^ n[22391];
assign t[22392] = t[22391] ^ n[22392];
assign t[22393] = t[22392] ^ n[22393];
assign t[22394] = t[22393] ^ n[22394];
assign t[22395] = t[22394] ^ n[22395];
assign t[22396] = t[22395] ^ n[22396];
assign t[22397] = t[22396] ^ n[22397];
assign t[22398] = t[22397] ^ n[22398];
assign t[22399] = t[22398] ^ n[22399];
assign t[22400] = t[22399] ^ n[22400];
assign t[22401] = t[22400] ^ n[22401];
assign t[22402] = t[22401] ^ n[22402];
assign t[22403] = t[22402] ^ n[22403];
assign t[22404] = t[22403] ^ n[22404];
assign t[22405] = t[22404] ^ n[22405];
assign t[22406] = t[22405] ^ n[22406];
assign t[22407] = t[22406] ^ n[22407];
assign t[22408] = t[22407] ^ n[22408];
assign t[22409] = t[22408] ^ n[22409];
assign t[22410] = t[22409] ^ n[22410];
assign t[22411] = t[22410] ^ n[22411];
assign t[22412] = t[22411] ^ n[22412];
assign t[22413] = t[22412] ^ n[22413];
assign t[22414] = t[22413] ^ n[22414];
assign t[22415] = t[22414] ^ n[22415];
assign t[22416] = t[22415] ^ n[22416];
assign t[22417] = t[22416] ^ n[22417];
assign t[22418] = t[22417] ^ n[22418];
assign t[22419] = t[22418] ^ n[22419];
assign t[22420] = t[22419] ^ n[22420];
assign t[22421] = t[22420] ^ n[22421];
assign t[22422] = t[22421] ^ n[22422];
assign t[22423] = t[22422] ^ n[22423];
assign t[22424] = t[22423] ^ n[22424];
assign t[22425] = t[22424] ^ n[22425];
assign t[22426] = t[22425] ^ n[22426];
assign t[22427] = t[22426] ^ n[22427];
assign t[22428] = t[22427] ^ n[22428];
assign t[22429] = t[22428] ^ n[22429];
assign t[22430] = t[22429] ^ n[22430];
assign t[22431] = t[22430] ^ n[22431];
assign t[22432] = t[22431] ^ n[22432];
assign t[22433] = t[22432] ^ n[22433];
assign t[22434] = t[22433] ^ n[22434];
assign t[22435] = t[22434] ^ n[22435];
assign t[22436] = t[22435] ^ n[22436];
assign t[22437] = t[22436] ^ n[22437];
assign t[22438] = t[22437] ^ n[22438];
assign t[22439] = t[22438] ^ n[22439];
assign t[22440] = t[22439] ^ n[22440];
assign t[22441] = t[22440] ^ n[22441];
assign t[22442] = t[22441] ^ n[22442];
assign t[22443] = t[22442] ^ n[22443];
assign t[22444] = t[22443] ^ n[22444];
assign t[22445] = t[22444] ^ n[22445];
assign t[22446] = t[22445] ^ n[22446];
assign t[22447] = t[22446] ^ n[22447];
assign t[22448] = t[22447] ^ n[22448];
assign t[22449] = t[22448] ^ n[22449];
assign t[22450] = t[22449] ^ n[22450];
assign t[22451] = t[22450] ^ n[22451];
assign t[22452] = t[22451] ^ n[22452];
assign t[22453] = t[22452] ^ n[22453];
assign t[22454] = t[22453] ^ n[22454];
assign t[22455] = t[22454] ^ n[22455];
assign t[22456] = t[22455] ^ n[22456];
assign t[22457] = t[22456] ^ n[22457];
assign t[22458] = t[22457] ^ n[22458];
assign t[22459] = t[22458] ^ n[22459];
assign t[22460] = t[22459] ^ n[22460];
assign t[22461] = t[22460] ^ n[22461];
assign t[22462] = t[22461] ^ n[22462];
assign t[22463] = t[22462] ^ n[22463];
assign t[22464] = t[22463] ^ n[22464];
assign t[22465] = t[22464] ^ n[22465];
assign t[22466] = t[22465] ^ n[22466];
assign t[22467] = t[22466] ^ n[22467];
assign t[22468] = t[22467] ^ n[22468];
assign t[22469] = t[22468] ^ n[22469];
assign t[22470] = t[22469] ^ n[22470];
assign t[22471] = t[22470] ^ n[22471];
assign t[22472] = t[22471] ^ n[22472];
assign t[22473] = t[22472] ^ n[22473];
assign t[22474] = t[22473] ^ n[22474];
assign t[22475] = t[22474] ^ n[22475];
assign t[22476] = t[22475] ^ n[22476];
assign t[22477] = t[22476] ^ n[22477];
assign t[22478] = t[22477] ^ n[22478];
assign t[22479] = t[22478] ^ n[22479];
assign t[22480] = t[22479] ^ n[22480];
assign t[22481] = t[22480] ^ n[22481];
assign t[22482] = t[22481] ^ n[22482];
assign t[22483] = t[22482] ^ n[22483];
assign t[22484] = t[22483] ^ n[22484];
assign t[22485] = t[22484] ^ n[22485];
assign t[22486] = t[22485] ^ n[22486];
assign t[22487] = t[22486] ^ n[22487];
assign t[22488] = t[22487] ^ n[22488];
assign t[22489] = t[22488] ^ n[22489];
assign t[22490] = t[22489] ^ n[22490];
assign t[22491] = t[22490] ^ n[22491];
assign t[22492] = t[22491] ^ n[22492];
assign t[22493] = t[22492] ^ n[22493];
assign t[22494] = t[22493] ^ n[22494];
assign t[22495] = t[22494] ^ n[22495];
assign t[22496] = t[22495] ^ n[22496];
assign t[22497] = t[22496] ^ n[22497];
assign t[22498] = t[22497] ^ n[22498];
assign t[22499] = t[22498] ^ n[22499];
assign t[22500] = t[22499] ^ n[22500];
assign t[22501] = t[22500] ^ n[22501];
assign t[22502] = t[22501] ^ n[22502];
assign t[22503] = t[22502] ^ n[22503];
assign t[22504] = t[22503] ^ n[22504];
assign t[22505] = t[22504] ^ n[22505];
assign t[22506] = t[22505] ^ n[22506];
assign t[22507] = t[22506] ^ n[22507];
assign t[22508] = t[22507] ^ n[22508];
assign t[22509] = t[22508] ^ n[22509];
assign t[22510] = t[22509] ^ n[22510];
assign t[22511] = t[22510] ^ n[22511];
assign t[22512] = t[22511] ^ n[22512];
assign t[22513] = t[22512] ^ n[22513];
assign t[22514] = t[22513] ^ n[22514];
assign t[22515] = t[22514] ^ n[22515];
assign t[22516] = t[22515] ^ n[22516];
assign t[22517] = t[22516] ^ n[22517];
assign t[22518] = t[22517] ^ n[22518];
assign t[22519] = t[22518] ^ n[22519];
assign t[22520] = t[22519] ^ n[22520];
assign t[22521] = t[22520] ^ n[22521];
assign t[22522] = t[22521] ^ n[22522];
assign t[22523] = t[22522] ^ n[22523];
assign t[22524] = t[22523] ^ n[22524];
assign t[22525] = t[22524] ^ n[22525];
assign t[22526] = t[22525] ^ n[22526];
assign t[22527] = t[22526] ^ n[22527];
assign t[22528] = t[22527] ^ n[22528];
assign t[22529] = t[22528] ^ n[22529];
assign t[22530] = t[22529] ^ n[22530];
assign t[22531] = t[22530] ^ n[22531];
assign t[22532] = t[22531] ^ n[22532];
assign t[22533] = t[22532] ^ n[22533];
assign t[22534] = t[22533] ^ n[22534];
assign t[22535] = t[22534] ^ n[22535];
assign t[22536] = t[22535] ^ n[22536];
assign t[22537] = t[22536] ^ n[22537];
assign t[22538] = t[22537] ^ n[22538];
assign t[22539] = t[22538] ^ n[22539];
assign t[22540] = t[22539] ^ n[22540];
assign t[22541] = t[22540] ^ n[22541];
assign t[22542] = t[22541] ^ n[22542];
assign t[22543] = t[22542] ^ n[22543];
assign t[22544] = t[22543] ^ n[22544];
assign t[22545] = t[22544] ^ n[22545];
assign t[22546] = t[22545] ^ n[22546];
assign t[22547] = t[22546] ^ n[22547];
assign t[22548] = t[22547] ^ n[22548];
assign t[22549] = t[22548] ^ n[22549];
assign t[22550] = t[22549] ^ n[22550];
assign t[22551] = t[22550] ^ n[22551];
assign t[22552] = t[22551] ^ n[22552];
assign t[22553] = t[22552] ^ n[22553];
assign t[22554] = t[22553] ^ n[22554];
assign t[22555] = t[22554] ^ n[22555];
assign t[22556] = t[22555] ^ n[22556];
assign t[22557] = t[22556] ^ n[22557];
assign t[22558] = t[22557] ^ n[22558];
assign t[22559] = t[22558] ^ n[22559];
assign t[22560] = t[22559] ^ n[22560];
assign t[22561] = t[22560] ^ n[22561];
assign t[22562] = t[22561] ^ n[22562];
assign t[22563] = t[22562] ^ n[22563];
assign t[22564] = t[22563] ^ n[22564];
assign t[22565] = t[22564] ^ n[22565];
assign t[22566] = t[22565] ^ n[22566];
assign t[22567] = t[22566] ^ n[22567];
assign t[22568] = t[22567] ^ n[22568];
assign t[22569] = t[22568] ^ n[22569];
assign t[22570] = t[22569] ^ n[22570];
assign t[22571] = t[22570] ^ n[22571];
assign t[22572] = t[22571] ^ n[22572];
assign t[22573] = t[22572] ^ n[22573];
assign t[22574] = t[22573] ^ n[22574];
assign t[22575] = t[22574] ^ n[22575];
assign t[22576] = t[22575] ^ n[22576];
assign t[22577] = t[22576] ^ n[22577];
assign t[22578] = t[22577] ^ n[22578];
assign t[22579] = t[22578] ^ n[22579];
assign t[22580] = t[22579] ^ n[22580];
assign t[22581] = t[22580] ^ n[22581];
assign t[22582] = t[22581] ^ n[22582];
assign t[22583] = t[22582] ^ n[22583];
assign t[22584] = t[22583] ^ n[22584];
assign t[22585] = t[22584] ^ n[22585];
assign t[22586] = t[22585] ^ n[22586];
assign t[22587] = t[22586] ^ n[22587];
assign t[22588] = t[22587] ^ n[22588];
assign t[22589] = t[22588] ^ n[22589];
assign t[22590] = t[22589] ^ n[22590];
assign t[22591] = t[22590] ^ n[22591];
assign t[22592] = t[22591] ^ n[22592];
assign t[22593] = t[22592] ^ n[22593];
assign t[22594] = t[22593] ^ n[22594];
assign t[22595] = t[22594] ^ n[22595];
assign t[22596] = t[22595] ^ n[22596];
assign t[22597] = t[22596] ^ n[22597];
assign t[22598] = t[22597] ^ n[22598];
assign t[22599] = t[22598] ^ n[22599];
assign t[22600] = t[22599] ^ n[22600];
assign t[22601] = t[22600] ^ n[22601];
assign t[22602] = t[22601] ^ n[22602];
assign t[22603] = t[22602] ^ n[22603];
assign t[22604] = t[22603] ^ n[22604];
assign t[22605] = t[22604] ^ n[22605];
assign t[22606] = t[22605] ^ n[22606];
assign t[22607] = t[22606] ^ n[22607];
assign t[22608] = t[22607] ^ n[22608];
assign t[22609] = t[22608] ^ n[22609];
assign t[22610] = t[22609] ^ n[22610];
assign t[22611] = t[22610] ^ n[22611];
assign t[22612] = t[22611] ^ n[22612];
assign t[22613] = t[22612] ^ n[22613];
assign t[22614] = t[22613] ^ n[22614];
assign t[22615] = t[22614] ^ n[22615];
assign t[22616] = t[22615] ^ n[22616];
assign t[22617] = t[22616] ^ n[22617];
assign t[22618] = t[22617] ^ n[22618];
assign t[22619] = t[22618] ^ n[22619];
assign t[22620] = t[22619] ^ n[22620];
assign t[22621] = t[22620] ^ n[22621];
assign t[22622] = t[22621] ^ n[22622];
assign t[22623] = t[22622] ^ n[22623];
assign t[22624] = t[22623] ^ n[22624];
assign t[22625] = t[22624] ^ n[22625];
assign t[22626] = t[22625] ^ n[22626];
assign t[22627] = t[22626] ^ n[22627];
assign t[22628] = t[22627] ^ n[22628];
assign t[22629] = t[22628] ^ n[22629];
assign t[22630] = t[22629] ^ n[22630];
assign t[22631] = t[22630] ^ n[22631];
assign t[22632] = t[22631] ^ n[22632];
assign t[22633] = t[22632] ^ n[22633];
assign t[22634] = t[22633] ^ n[22634];
assign t[22635] = t[22634] ^ n[22635];
assign t[22636] = t[22635] ^ n[22636];
assign t[22637] = t[22636] ^ n[22637];
assign t[22638] = t[22637] ^ n[22638];
assign t[22639] = t[22638] ^ n[22639];
assign t[22640] = t[22639] ^ n[22640];
assign t[22641] = t[22640] ^ n[22641];
assign t[22642] = t[22641] ^ n[22642];
assign t[22643] = t[22642] ^ n[22643];
assign t[22644] = t[22643] ^ n[22644];
assign t[22645] = t[22644] ^ n[22645];
assign t[22646] = t[22645] ^ n[22646];
assign t[22647] = t[22646] ^ n[22647];
assign t[22648] = t[22647] ^ n[22648];
assign t[22649] = t[22648] ^ n[22649];
assign t[22650] = t[22649] ^ n[22650];
assign t[22651] = t[22650] ^ n[22651];
assign t[22652] = t[22651] ^ n[22652];
assign t[22653] = t[22652] ^ n[22653];
assign t[22654] = t[22653] ^ n[22654];
assign t[22655] = t[22654] ^ n[22655];
assign t[22656] = t[22655] ^ n[22656];
assign t[22657] = t[22656] ^ n[22657];
assign t[22658] = t[22657] ^ n[22658];
assign t[22659] = t[22658] ^ n[22659];
assign t[22660] = t[22659] ^ n[22660];
assign t[22661] = t[22660] ^ n[22661];
assign t[22662] = t[22661] ^ n[22662];
assign t[22663] = t[22662] ^ n[22663];
assign t[22664] = t[22663] ^ n[22664];
assign t[22665] = t[22664] ^ n[22665];
assign t[22666] = t[22665] ^ n[22666];
assign t[22667] = t[22666] ^ n[22667];
assign t[22668] = t[22667] ^ n[22668];
assign t[22669] = t[22668] ^ n[22669];
assign t[22670] = t[22669] ^ n[22670];
assign t[22671] = t[22670] ^ n[22671];
assign t[22672] = t[22671] ^ n[22672];
assign t[22673] = t[22672] ^ n[22673];
assign t[22674] = t[22673] ^ n[22674];
assign t[22675] = t[22674] ^ n[22675];
assign t[22676] = t[22675] ^ n[22676];
assign t[22677] = t[22676] ^ n[22677];
assign t[22678] = t[22677] ^ n[22678];
assign t[22679] = t[22678] ^ n[22679];
assign t[22680] = t[22679] ^ n[22680];
assign t[22681] = t[22680] ^ n[22681];
assign t[22682] = t[22681] ^ n[22682];
assign t[22683] = t[22682] ^ n[22683];
assign t[22684] = t[22683] ^ n[22684];
assign t[22685] = t[22684] ^ n[22685];
assign t[22686] = t[22685] ^ n[22686];
assign t[22687] = t[22686] ^ n[22687];
assign t[22688] = t[22687] ^ n[22688];
assign t[22689] = t[22688] ^ n[22689];
assign t[22690] = t[22689] ^ n[22690];
assign t[22691] = t[22690] ^ n[22691];
assign t[22692] = t[22691] ^ n[22692];
assign t[22693] = t[22692] ^ n[22693];
assign t[22694] = t[22693] ^ n[22694];
assign t[22695] = t[22694] ^ n[22695];
assign t[22696] = t[22695] ^ n[22696];
assign t[22697] = t[22696] ^ n[22697];
assign t[22698] = t[22697] ^ n[22698];
assign t[22699] = t[22698] ^ n[22699];
assign t[22700] = t[22699] ^ n[22700];
assign t[22701] = t[22700] ^ n[22701];
assign t[22702] = t[22701] ^ n[22702];
assign t[22703] = t[22702] ^ n[22703];
assign t[22704] = t[22703] ^ n[22704];
assign t[22705] = t[22704] ^ n[22705];
assign t[22706] = t[22705] ^ n[22706];
assign t[22707] = t[22706] ^ n[22707];
assign t[22708] = t[22707] ^ n[22708];
assign t[22709] = t[22708] ^ n[22709];
assign t[22710] = t[22709] ^ n[22710];
assign t[22711] = t[22710] ^ n[22711];
assign t[22712] = t[22711] ^ n[22712];
assign t[22713] = t[22712] ^ n[22713];
assign t[22714] = t[22713] ^ n[22714];
assign t[22715] = t[22714] ^ n[22715];
assign t[22716] = t[22715] ^ n[22716];
assign t[22717] = t[22716] ^ n[22717];
assign t[22718] = t[22717] ^ n[22718];
assign t[22719] = t[22718] ^ n[22719];
assign t[22720] = t[22719] ^ n[22720];
assign t[22721] = t[22720] ^ n[22721];
assign t[22722] = t[22721] ^ n[22722];
assign t[22723] = t[22722] ^ n[22723];
assign t[22724] = t[22723] ^ n[22724];
assign t[22725] = t[22724] ^ n[22725];
assign t[22726] = t[22725] ^ n[22726];
assign t[22727] = t[22726] ^ n[22727];
assign t[22728] = t[22727] ^ n[22728];
assign t[22729] = t[22728] ^ n[22729];
assign t[22730] = t[22729] ^ n[22730];
assign t[22731] = t[22730] ^ n[22731];
assign t[22732] = t[22731] ^ n[22732];
assign t[22733] = t[22732] ^ n[22733];
assign t[22734] = t[22733] ^ n[22734];
assign t[22735] = t[22734] ^ n[22735];
assign t[22736] = t[22735] ^ n[22736];
assign t[22737] = t[22736] ^ n[22737];
assign t[22738] = t[22737] ^ n[22738];
assign t[22739] = t[22738] ^ n[22739];
assign t[22740] = t[22739] ^ n[22740];
assign t[22741] = t[22740] ^ n[22741];
assign t[22742] = t[22741] ^ n[22742];
assign t[22743] = t[22742] ^ n[22743];
assign t[22744] = t[22743] ^ n[22744];
assign t[22745] = t[22744] ^ n[22745];
assign t[22746] = t[22745] ^ n[22746];
assign t[22747] = t[22746] ^ n[22747];
assign t[22748] = t[22747] ^ n[22748];
assign t[22749] = t[22748] ^ n[22749];
assign t[22750] = t[22749] ^ n[22750];
assign t[22751] = t[22750] ^ n[22751];
assign t[22752] = t[22751] ^ n[22752];
assign t[22753] = t[22752] ^ n[22753];
assign t[22754] = t[22753] ^ n[22754];
assign t[22755] = t[22754] ^ n[22755];
assign t[22756] = t[22755] ^ n[22756];
assign t[22757] = t[22756] ^ n[22757];
assign t[22758] = t[22757] ^ n[22758];
assign t[22759] = t[22758] ^ n[22759];
assign t[22760] = t[22759] ^ n[22760];
assign t[22761] = t[22760] ^ n[22761];
assign t[22762] = t[22761] ^ n[22762];
assign t[22763] = t[22762] ^ n[22763];
assign t[22764] = t[22763] ^ n[22764];
assign t[22765] = t[22764] ^ n[22765];
assign t[22766] = t[22765] ^ n[22766];
assign t[22767] = t[22766] ^ n[22767];
assign t[22768] = t[22767] ^ n[22768];
assign t[22769] = t[22768] ^ n[22769];
assign t[22770] = t[22769] ^ n[22770];
assign t[22771] = t[22770] ^ n[22771];
assign t[22772] = t[22771] ^ n[22772];
assign t[22773] = t[22772] ^ n[22773];
assign t[22774] = t[22773] ^ n[22774];
assign t[22775] = t[22774] ^ n[22775];
assign t[22776] = t[22775] ^ n[22776];
assign t[22777] = t[22776] ^ n[22777];
assign t[22778] = t[22777] ^ n[22778];
assign t[22779] = t[22778] ^ n[22779];
assign t[22780] = t[22779] ^ n[22780];
assign t[22781] = t[22780] ^ n[22781];
assign t[22782] = t[22781] ^ n[22782];
assign t[22783] = t[22782] ^ n[22783];
assign t[22784] = t[22783] ^ n[22784];
assign t[22785] = t[22784] ^ n[22785];
assign t[22786] = t[22785] ^ n[22786];
assign t[22787] = t[22786] ^ n[22787];
assign t[22788] = t[22787] ^ n[22788];
assign t[22789] = t[22788] ^ n[22789];
assign t[22790] = t[22789] ^ n[22790];
assign t[22791] = t[22790] ^ n[22791];
assign t[22792] = t[22791] ^ n[22792];
assign t[22793] = t[22792] ^ n[22793];
assign t[22794] = t[22793] ^ n[22794];
assign t[22795] = t[22794] ^ n[22795];
assign t[22796] = t[22795] ^ n[22796];
assign t[22797] = t[22796] ^ n[22797];
assign t[22798] = t[22797] ^ n[22798];
assign t[22799] = t[22798] ^ n[22799];
assign t[22800] = t[22799] ^ n[22800];
assign t[22801] = t[22800] ^ n[22801];
assign t[22802] = t[22801] ^ n[22802];
assign t[22803] = t[22802] ^ n[22803];
assign t[22804] = t[22803] ^ n[22804];
assign t[22805] = t[22804] ^ n[22805];
assign t[22806] = t[22805] ^ n[22806];
assign t[22807] = t[22806] ^ n[22807];
assign t[22808] = t[22807] ^ n[22808];
assign t[22809] = t[22808] ^ n[22809];
assign t[22810] = t[22809] ^ n[22810];
assign t[22811] = t[22810] ^ n[22811];
assign t[22812] = t[22811] ^ n[22812];
assign t[22813] = t[22812] ^ n[22813];
assign t[22814] = t[22813] ^ n[22814];
assign t[22815] = t[22814] ^ n[22815];
assign t[22816] = t[22815] ^ n[22816];
assign t[22817] = t[22816] ^ n[22817];
assign t[22818] = t[22817] ^ n[22818];
assign t[22819] = t[22818] ^ n[22819];
assign t[22820] = t[22819] ^ n[22820];
assign t[22821] = t[22820] ^ n[22821];
assign t[22822] = t[22821] ^ n[22822];
assign t[22823] = t[22822] ^ n[22823];
assign t[22824] = t[22823] ^ n[22824];
assign t[22825] = t[22824] ^ n[22825];
assign t[22826] = t[22825] ^ n[22826];
assign t[22827] = t[22826] ^ n[22827];
assign t[22828] = t[22827] ^ n[22828];
assign t[22829] = t[22828] ^ n[22829];
assign t[22830] = t[22829] ^ n[22830];
assign t[22831] = t[22830] ^ n[22831];
assign t[22832] = t[22831] ^ n[22832];
assign t[22833] = t[22832] ^ n[22833];
assign t[22834] = t[22833] ^ n[22834];
assign t[22835] = t[22834] ^ n[22835];
assign t[22836] = t[22835] ^ n[22836];
assign t[22837] = t[22836] ^ n[22837];
assign t[22838] = t[22837] ^ n[22838];
assign t[22839] = t[22838] ^ n[22839];
assign t[22840] = t[22839] ^ n[22840];
assign t[22841] = t[22840] ^ n[22841];
assign t[22842] = t[22841] ^ n[22842];
assign t[22843] = t[22842] ^ n[22843];
assign t[22844] = t[22843] ^ n[22844];
assign t[22845] = t[22844] ^ n[22845];
assign t[22846] = t[22845] ^ n[22846];
assign t[22847] = t[22846] ^ n[22847];
assign t[22848] = t[22847] ^ n[22848];
assign t[22849] = t[22848] ^ n[22849];
assign t[22850] = t[22849] ^ n[22850];
assign t[22851] = t[22850] ^ n[22851];
assign t[22852] = t[22851] ^ n[22852];
assign t[22853] = t[22852] ^ n[22853];
assign t[22854] = t[22853] ^ n[22854];
assign t[22855] = t[22854] ^ n[22855];
assign t[22856] = t[22855] ^ n[22856];
assign t[22857] = t[22856] ^ n[22857];
assign t[22858] = t[22857] ^ n[22858];
assign t[22859] = t[22858] ^ n[22859];
assign t[22860] = t[22859] ^ n[22860];
assign t[22861] = t[22860] ^ n[22861];
assign t[22862] = t[22861] ^ n[22862];
assign t[22863] = t[22862] ^ n[22863];
assign t[22864] = t[22863] ^ n[22864];
assign t[22865] = t[22864] ^ n[22865];
assign t[22866] = t[22865] ^ n[22866];
assign t[22867] = t[22866] ^ n[22867];
assign t[22868] = t[22867] ^ n[22868];
assign t[22869] = t[22868] ^ n[22869];
assign t[22870] = t[22869] ^ n[22870];
assign t[22871] = t[22870] ^ n[22871];
assign t[22872] = t[22871] ^ n[22872];
assign t[22873] = t[22872] ^ n[22873];
assign t[22874] = t[22873] ^ n[22874];
assign t[22875] = t[22874] ^ n[22875];
assign t[22876] = t[22875] ^ n[22876];
assign t[22877] = t[22876] ^ n[22877];
assign t[22878] = t[22877] ^ n[22878];
assign t[22879] = t[22878] ^ n[22879];
assign t[22880] = t[22879] ^ n[22880];
assign t[22881] = t[22880] ^ n[22881];
assign t[22882] = t[22881] ^ n[22882];
assign t[22883] = t[22882] ^ n[22883];
assign t[22884] = t[22883] ^ n[22884];
assign t[22885] = t[22884] ^ n[22885];
assign t[22886] = t[22885] ^ n[22886];
assign t[22887] = t[22886] ^ n[22887];
assign t[22888] = t[22887] ^ n[22888];
assign t[22889] = t[22888] ^ n[22889];
assign t[22890] = t[22889] ^ n[22890];
assign t[22891] = t[22890] ^ n[22891];
assign t[22892] = t[22891] ^ n[22892];
assign t[22893] = t[22892] ^ n[22893];
assign t[22894] = t[22893] ^ n[22894];
assign t[22895] = t[22894] ^ n[22895];
assign t[22896] = t[22895] ^ n[22896];
assign t[22897] = t[22896] ^ n[22897];
assign t[22898] = t[22897] ^ n[22898];
assign t[22899] = t[22898] ^ n[22899];
assign t[22900] = t[22899] ^ n[22900];
assign t[22901] = t[22900] ^ n[22901];
assign t[22902] = t[22901] ^ n[22902];
assign t[22903] = t[22902] ^ n[22903];
assign t[22904] = t[22903] ^ n[22904];
assign t[22905] = t[22904] ^ n[22905];
assign t[22906] = t[22905] ^ n[22906];
assign t[22907] = t[22906] ^ n[22907];
assign t[22908] = t[22907] ^ n[22908];
assign t[22909] = t[22908] ^ n[22909];
assign t[22910] = t[22909] ^ n[22910];
assign t[22911] = t[22910] ^ n[22911];
assign t[22912] = t[22911] ^ n[22912];
assign t[22913] = t[22912] ^ n[22913];
assign t[22914] = t[22913] ^ n[22914];
assign t[22915] = t[22914] ^ n[22915];
assign t[22916] = t[22915] ^ n[22916];
assign t[22917] = t[22916] ^ n[22917];
assign t[22918] = t[22917] ^ n[22918];
assign t[22919] = t[22918] ^ n[22919];
assign t[22920] = t[22919] ^ n[22920];
assign t[22921] = t[22920] ^ n[22921];
assign t[22922] = t[22921] ^ n[22922];
assign t[22923] = t[22922] ^ n[22923];
assign t[22924] = t[22923] ^ n[22924];
assign t[22925] = t[22924] ^ n[22925];
assign t[22926] = t[22925] ^ n[22926];
assign t[22927] = t[22926] ^ n[22927];
assign t[22928] = t[22927] ^ n[22928];
assign t[22929] = t[22928] ^ n[22929];
assign t[22930] = t[22929] ^ n[22930];
assign t[22931] = t[22930] ^ n[22931];
assign t[22932] = t[22931] ^ n[22932];
assign t[22933] = t[22932] ^ n[22933];
assign t[22934] = t[22933] ^ n[22934];
assign t[22935] = t[22934] ^ n[22935];
assign t[22936] = t[22935] ^ n[22936];
assign t[22937] = t[22936] ^ n[22937];
assign t[22938] = t[22937] ^ n[22938];
assign t[22939] = t[22938] ^ n[22939];
assign t[22940] = t[22939] ^ n[22940];
assign t[22941] = t[22940] ^ n[22941];
assign t[22942] = t[22941] ^ n[22942];
assign t[22943] = t[22942] ^ n[22943];
assign t[22944] = t[22943] ^ n[22944];
assign t[22945] = t[22944] ^ n[22945];
assign t[22946] = t[22945] ^ n[22946];
assign t[22947] = t[22946] ^ n[22947];
assign t[22948] = t[22947] ^ n[22948];
assign t[22949] = t[22948] ^ n[22949];
assign t[22950] = t[22949] ^ n[22950];
assign t[22951] = t[22950] ^ n[22951];
assign t[22952] = t[22951] ^ n[22952];
assign t[22953] = t[22952] ^ n[22953];
assign t[22954] = t[22953] ^ n[22954];
assign t[22955] = t[22954] ^ n[22955];
assign t[22956] = t[22955] ^ n[22956];
assign t[22957] = t[22956] ^ n[22957];
assign t[22958] = t[22957] ^ n[22958];
assign t[22959] = t[22958] ^ n[22959];
assign t[22960] = t[22959] ^ n[22960];
assign t[22961] = t[22960] ^ n[22961];
assign t[22962] = t[22961] ^ n[22962];
assign t[22963] = t[22962] ^ n[22963];
assign t[22964] = t[22963] ^ n[22964];
assign t[22965] = t[22964] ^ n[22965];
assign t[22966] = t[22965] ^ n[22966];
assign t[22967] = t[22966] ^ n[22967];
assign t[22968] = t[22967] ^ n[22968];
assign t[22969] = t[22968] ^ n[22969];
assign t[22970] = t[22969] ^ n[22970];
assign t[22971] = t[22970] ^ n[22971];
assign t[22972] = t[22971] ^ n[22972];
assign t[22973] = t[22972] ^ n[22973];
assign t[22974] = t[22973] ^ n[22974];
assign t[22975] = t[22974] ^ n[22975];
assign t[22976] = t[22975] ^ n[22976];
assign t[22977] = t[22976] ^ n[22977];
assign t[22978] = t[22977] ^ n[22978];
assign t[22979] = t[22978] ^ n[22979];
assign t[22980] = t[22979] ^ n[22980];
assign t[22981] = t[22980] ^ n[22981];
assign t[22982] = t[22981] ^ n[22982];
assign t[22983] = t[22982] ^ n[22983];
assign t[22984] = t[22983] ^ n[22984];
assign t[22985] = t[22984] ^ n[22985];
assign t[22986] = t[22985] ^ n[22986];
assign t[22987] = t[22986] ^ n[22987];
assign t[22988] = t[22987] ^ n[22988];
assign t[22989] = t[22988] ^ n[22989];
assign t[22990] = t[22989] ^ n[22990];
assign t[22991] = t[22990] ^ n[22991];
assign t[22992] = t[22991] ^ n[22992];
assign t[22993] = t[22992] ^ n[22993];
assign t[22994] = t[22993] ^ n[22994];
assign t[22995] = t[22994] ^ n[22995];
assign t[22996] = t[22995] ^ n[22996];
assign t[22997] = t[22996] ^ n[22997];
assign t[22998] = t[22997] ^ n[22998];
assign t[22999] = t[22998] ^ n[22999];
assign t[23000] = t[22999] ^ n[23000];
assign t[23001] = t[23000] ^ n[23001];
assign t[23002] = t[23001] ^ n[23002];
assign t[23003] = t[23002] ^ n[23003];
assign t[23004] = t[23003] ^ n[23004];
assign t[23005] = t[23004] ^ n[23005];
assign t[23006] = t[23005] ^ n[23006];
assign t[23007] = t[23006] ^ n[23007];
assign t[23008] = t[23007] ^ n[23008];
assign t[23009] = t[23008] ^ n[23009];
assign t[23010] = t[23009] ^ n[23010];
assign t[23011] = t[23010] ^ n[23011];
assign t[23012] = t[23011] ^ n[23012];
assign t[23013] = t[23012] ^ n[23013];
assign t[23014] = t[23013] ^ n[23014];
assign t[23015] = t[23014] ^ n[23015];
assign t[23016] = t[23015] ^ n[23016];
assign t[23017] = t[23016] ^ n[23017];
assign t[23018] = t[23017] ^ n[23018];
assign t[23019] = t[23018] ^ n[23019];
assign t[23020] = t[23019] ^ n[23020];
assign t[23021] = t[23020] ^ n[23021];
assign t[23022] = t[23021] ^ n[23022];
assign t[23023] = t[23022] ^ n[23023];
assign t[23024] = t[23023] ^ n[23024];
assign t[23025] = t[23024] ^ n[23025];
assign t[23026] = t[23025] ^ n[23026];
assign t[23027] = t[23026] ^ n[23027];
assign t[23028] = t[23027] ^ n[23028];
assign t[23029] = t[23028] ^ n[23029];
assign t[23030] = t[23029] ^ n[23030];
assign t[23031] = t[23030] ^ n[23031];
assign t[23032] = t[23031] ^ n[23032];
assign t[23033] = t[23032] ^ n[23033];
assign t[23034] = t[23033] ^ n[23034];
assign t[23035] = t[23034] ^ n[23035];
assign t[23036] = t[23035] ^ n[23036];
assign t[23037] = t[23036] ^ n[23037];
assign t[23038] = t[23037] ^ n[23038];
assign t[23039] = t[23038] ^ n[23039];
assign t[23040] = t[23039] ^ n[23040];
assign t[23041] = t[23040] ^ n[23041];
assign t[23042] = t[23041] ^ n[23042];
assign t[23043] = t[23042] ^ n[23043];
assign t[23044] = t[23043] ^ n[23044];
assign t[23045] = t[23044] ^ n[23045];
assign t[23046] = t[23045] ^ n[23046];
assign t[23047] = t[23046] ^ n[23047];
assign t[23048] = t[23047] ^ n[23048];
assign t[23049] = t[23048] ^ n[23049];
assign t[23050] = t[23049] ^ n[23050];
assign t[23051] = t[23050] ^ n[23051];
assign t[23052] = t[23051] ^ n[23052];
assign t[23053] = t[23052] ^ n[23053];
assign t[23054] = t[23053] ^ n[23054];
assign t[23055] = t[23054] ^ n[23055];
assign t[23056] = t[23055] ^ n[23056];
assign t[23057] = t[23056] ^ n[23057];
assign t[23058] = t[23057] ^ n[23058];
assign t[23059] = t[23058] ^ n[23059];
assign t[23060] = t[23059] ^ n[23060];
assign t[23061] = t[23060] ^ n[23061];
assign t[23062] = t[23061] ^ n[23062];
assign t[23063] = t[23062] ^ n[23063];
assign t[23064] = t[23063] ^ n[23064];
assign t[23065] = t[23064] ^ n[23065];
assign t[23066] = t[23065] ^ n[23066];
assign t[23067] = t[23066] ^ n[23067];
assign t[23068] = t[23067] ^ n[23068];
assign t[23069] = t[23068] ^ n[23069];
assign t[23070] = t[23069] ^ n[23070];
assign t[23071] = t[23070] ^ n[23071];
assign t[23072] = t[23071] ^ n[23072];
assign t[23073] = t[23072] ^ n[23073];
assign t[23074] = t[23073] ^ n[23074];
assign t[23075] = t[23074] ^ n[23075];
assign t[23076] = t[23075] ^ n[23076];
assign t[23077] = t[23076] ^ n[23077];
assign t[23078] = t[23077] ^ n[23078];
assign t[23079] = t[23078] ^ n[23079];
assign t[23080] = t[23079] ^ n[23080];
assign t[23081] = t[23080] ^ n[23081];
assign t[23082] = t[23081] ^ n[23082];
assign t[23083] = t[23082] ^ n[23083];
assign t[23084] = t[23083] ^ n[23084];
assign t[23085] = t[23084] ^ n[23085];
assign t[23086] = t[23085] ^ n[23086];
assign t[23087] = t[23086] ^ n[23087];
assign t[23088] = t[23087] ^ n[23088];
assign t[23089] = t[23088] ^ n[23089];
assign t[23090] = t[23089] ^ n[23090];
assign t[23091] = t[23090] ^ n[23091];
assign t[23092] = t[23091] ^ n[23092];
assign t[23093] = t[23092] ^ n[23093];
assign t[23094] = t[23093] ^ n[23094];
assign t[23095] = t[23094] ^ n[23095];
assign t[23096] = t[23095] ^ n[23096];
assign t[23097] = t[23096] ^ n[23097];
assign t[23098] = t[23097] ^ n[23098];
assign t[23099] = t[23098] ^ n[23099];
assign t[23100] = t[23099] ^ n[23100];
assign t[23101] = t[23100] ^ n[23101];
assign t[23102] = t[23101] ^ n[23102];
assign t[23103] = t[23102] ^ n[23103];
assign t[23104] = t[23103] ^ n[23104];
assign t[23105] = t[23104] ^ n[23105];
assign t[23106] = t[23105] ^ n[23106];
assign t[23107] = t[23106] ^ n[23107];
assign t[23108] = t[23107] ^ n[23108];
assign t[23109] = t[23108] ^ n[23109];
assign t[23110] = t[23109] ^ n[23110];
assign t[23111] = t[23110] ^ n[23111];
assign t[23112] = t[23111] ^ n[23112];
assign t[23113] = t[23112] ^ n[23113];
assign t[23114] = t[23113] ^ n[23114];
assign t[23115] = t[23114] ^ n[23115];
assign t[23116] = t[23115] ^ n[23116];
assign t[23117] = t[23116] ^ n[23117];
assign t[23118] = t[23117] ^ n[23118];
assign t[23119] = t[23118] ^ n[23119];
assign t[23120] = t[23119] ^ n[23120];
assign t[23121] = t[23120] ^ n[23121];
assign t[23122] = t[23121] ^ n[23122];
assign t[23123] = t[23122] ^ n[23123];
assign t[23124] = t[23123] ^ n[23124];
assign t[23125] = t[23124] ^ n[23125];
assign t[23126] = t[23125] ^ n[23126];
assign t[23127] = t[23126] ^ n[23127];
assign t[23128] = t[23127] ^ n[23128];
assign t[23129] = t[23128] ^ n[23129];
assign t[23130] = t[23129] ^ n[23130];
assign t[23131] = t[23130] ^ n[23131];
assign t[23132] = t[23131] ^ n[23132];
assign t[23133] = t[23132] ^ n[23133];
assign t[23134] = t[23133] ^ n[23134];
assign t[23135] = t[23134] ^ n[23135];
assign t[23136] = t[23135] ^ n[23136];
assign t[23137] = t[23136] ^ n[23137];
assign t[23138] = t[23137] ^ n[23138];
assign t[23139] = t[23138] ^ n[23139];
assign t[23140] = t[23139] ^ n[23140];
assign t[23141] = t[23140] ^ n[23141];
assign t[23142] = t[23141] ^ n[23142];
assign t[23143] = t[23142] ^ n[23143];
assign t[23144] = t[23143] ^ n[23144];
assign t[23145] = t[23144] ^ n[23145];
assign t[23146] = t[23145] ^ n[23146];
assign t[23147] = t[23146] ^ n[23147];
assign t[23148] = t[23147] ^ n[23148];
assign t[23149] = t[23148] ^ n[23149];
assign t[23150] = t[23149] ^ n[23150];
assign t[23151] = t[23150] ^ n[23151];
assign t[23152] = t[23151] ^ n[23152];
assign t[23153] = t[23152] ^ n[23153];
assign t[23154] = t[23153] ^ n[23154];
assign t[23155] = t[23154] ^ n[23155];
assign t[23156] = t[23155] ^ n[23156];
assign t[23157] = t[23156] ^ n[23157];
assign t[23158] = t[23157] ^ n[23158];
assign t[23159] = t[23158] ^ n[23159];
assign t[23160] = t[23159] ^ n[23160];
assign t[23161] = t[23160] ^ n[23161];
assign t[23162] = t[23161] ^ n[23162];
assign t[23163] = t[23162] ^ n[23163];
assign t[23164] = t[23163] ^ n[23164];
assign t[23165] = t[23164] ^ n[23165];
assign t[23166] = t[23165] ^ n[23166];
assign t[23167] = t[23166] ^ n[23167];
assign t[23168] = t[23167] ^ n[23168];
assign t[23169] = t[23168] ^ n[23169];
assign t[23170] = t[23169] ^ n[23170];
assign t[23171] = t[23170] ^ n[23171];
assign t[23172] = t[23171] ^ n[23172];
assign t[23173] = t[23172] ^ n[23173];
assign t[23174] = t[23173] ^ n[23174];
assign t[23175] = t[23174] ^ n[23175];
assign t[23176] = t[23175] ^ n[23176];
assign t[23177] = t[23176] ^ n[23177];
assign t[23178] = t[23177] ^ n[23178];
assign t[23179] = t[23178] ^ n[23179];
assign t[23180] = t[23179] ^ n[23180];
assign t[23181] = t[23180] ^ n[23181];
assign t[23182] = t[23181] ^ n[23182];
assign t[23183] = t[23182] ^ n[23183];
assign t[23184] = t[23183] ^ n[23184];
assign t[23185] = t[23184] ^ n[23185];
assign t[23186] = t[23185] ^ n[23186];
assign t[23187] = t[23186] ^ n[23187];
assign t[23188] = t[23187] ^ n[23188];
assign t[23189] = t[23188] ^ n[23189];
assign t[23190] = t[23189] ^ n[23190];
assign t[23191] = t[23190] ^ n[23191];
assign t[23192] = t[23191] ^ n[23192];
assign t[23193] = t[23192] ^ n[23193];
assign t[23194] = t[23193] ^ n[23194];
assign t[23195] = t[23194] ^ n[23195];
assign t[23196] = t[23195] ^ n[23196];
assign t[23197] = t[23196] ^ n[23197];
assign t[23198] = t[23197] ^ n[23198];
assign t[23199] = t[23198] ^ n[23199];
assign t[23200] = t[23199] ^ n[23200];
assign t[23201] = t[23200] ^ n[23201];
assign t[23202] = t[23201] ^ n[23202];
assign t[23203] = t[23202] ^ n[23203];
assign t[23204] = t[23203] ^ n[23204];
assign t[23205] = t[23204] ^ n[23205];
assign t[23206] = t[23205] ^ n[23206];
assign t[23207] = t[23206] ^ n[23207];
assign t[23208] = t[23207] ^ n[23208];
assign t[23209] = t[23208] ^ n[23209];
assign t[23210] = t[23209] ^ n[23210];
assign t[23211] = t[23210] ^ n[23211];
assign t[23212] = t[23211] ^ n[23212];
assign t[23213] = t[23212] ^ n[23213];
assign t[23214] = t[23213] ^ n[23214];
assign t[23215] = t[23214] ^ n[23215];
assign t[23216] = t[23215] ^ n[23216];
assign t[23217] = t[23216] ^ n[23217];
assign t[23218] = t[23217] ^ n[23218];
assign t[23219] = t[23218] ^ n[23219];
assign t[23220] = t[23219] ^ n[23220];
assign t[23221] = t[23220] ^ n[23221];
assign t[23222] = t[23221] ^ n[23222];
assign t[23223] = t[23222] ^ n[23223];
assign t[23224] = t[23223] ^ n[23224];
assign t[23225] = t[23224] ^ n[23225];
assign t[23226] = t[23225] ^ n[23226];
assign t[23227] = t[23226] ^ n[23227];
assign t[23228] = t[23227] ^ n[23228];
assign t[23229] = t[23228] ^ n[23229];
assign t[23230] = t[23229] ^ n[23230];
assign t[23231] = t[23230] ^ n[23231];
assign t[23232] = t[23231] ^ n[23232];
assign t[23233] = t[23232] ^ n[23233];
assign t[23234] = t[23233] ^ n[23234];
assign t[23235] = t[23234] ^ n[23235];
assign t[23236] = t[23235] ^ n[23236];
assign t[23237] = t[23236] ^ n[23237];
assign t[23238] = t[23237] ^ n[23238];
assign t[23239] = t[23238] ^ n[23239];
assign t[23240] = t[23239] ^ n[23240];
assign t[23241] = t[23240] ^ n[23241];
assign t[23242] = t[23241] ^ n[23242];
assign t[23243] = t[23242] ^ n[23243];
assign t[23244] = t[23243] ^ n[23244];
assign t[23245] = t[23244] ^ n[23245];
assign t[23246] = t[23245] ^ n[23246];
assign t[23247] = t[23246] ^ n[23247];
assign t[23248] = t[23247] ^ n[23248];
assign t[23249] = t[23248] ^ n[23249];
assign t[23250] = t[23249] ^ n[23250];
assign t[23251] = t[23250] ^ n[23251];
assign t[23252] = t[23251] ^ n[23252];
assign t[23253] = t[23252] ^ n[23253];
assign t[23254] = t[23253] ^ n[23254];
assign t[23255] = t[23254] ^ n[23255];
assign t[23256] = t[23255] ^ n[23256];
assign t[23257] = t[23256] ^ n[23257];
assign t[23258] = t[23257] ^ n[23258];
assign t[23259] = t[23258] ^ n[23259];
assign t[23260] = t[23259] ^ n[23260];
assign t[23261] = t[23260] ^ n[23261];
assign t[23262] = t[23261] ^ n[23262];
assign t[23263] = t[23262] ^ n[23263];
assign t[23264] = t[23263] ^ n[23264];
assign t[23265] = t[23264] ^ n[23265];
assign t[23266] = t[23265] ^ n[23266];
assign t[23267] = t[23266] ^ n[23267];
assign t[23268] = t[23267] ^ n[23268];
assign t[23269] = t[23268] ^ n[23269];
assign t[23270] = t[23269] ^ n[23270];
assign t[23271] = t[23270] ^ n[23271];
assign t[23272] = t[23271] ^ n[23272];
assign t[23273] = t[23272] ^ n[23273];
assign t[23274] = t[23273] ^ n[23274];
assign t[23275] = t[23274] ^ n[23275];
assign t[23276] = t[23275] ^ n[23276];
assign t[23277] = t[23276] ^ n[23277];
assign t[23278] = t[23277] ^ n[23278];
assign t[23279] = t[23278] ^ n[23279];
assign t[23280] = t[23279] ^ n[23280];
assign t[23281] = t[23280] ^ n[23281];
assign t[23282] = t[23281] ^ n[23282];
assign t[23283] = t[23282] ^ n[23283];
assign t[23284] = t[23283] ^ n[23284];
assign t[23285] = t[23284] ^ n[23285];
assign t[23286] = t[23285] ^ n[23286];
assign t[23287] = t[23286] ^ n[23287];
assign t[23288] = t[23287] ^ n[23288];
assign t[23289] = t[23288] ^ n[23289];
assign t[23290] = t[23289] ^ n[23290];
assign t[23291] = t[23290] ^ n[23291];
assign t[23292] = t[23291] ^ n[23292];
assign t[23293] = t[23292] ^ n[23293];
assign t[23294] = t[23293] ^ n[23294];
assign t[23295] = t[23294] ^ n[23295];
assign t[23296] = t[23295] ^ n[23296];
assign t[23297] = t[23296] ^ n[23297];
assign t[23298] = t[23297] ^ n[23298];
assign t[23299] = t[23298] ^ n[23299];
assign t[23300] = t[23299] ^ n[23300];
assign t[23301] = t[23300] ^ n[23301];
assign t[23302] = t[23301] ^ n[23302];
assign t[23303] = t[23302] ^ n[23303];
assign t[23304] = t[23303] ^ n[23304];
assign t[23305] = t[23304] ^ n[23305];
assign t[23306] = t[23305] ^ n[23306];
assign t[23307] = t[23306] ^ n[23307];
assign t[23308] = t[23307] ^ n[23308];
assign t[23309] = t[23308] ^ n[23309];
assign t[23310] = t[23309] ^ n[23310];
assign t[23311] = t[23310] ^ n[23311];
assign t[23312] = t[23311] ^ n[23312];
assign t[23313] = t[23312] ^ n[23313];
assign t[23314] = t[23313] ^ n[23314];
assign t[23315] = t[23314] ^ n[23315];
assign t[23316] = t[23315] ^ n[23316];
assign t[23317] = t[23316] ^ n[23317];
assign t[23318] = t[23317] ^ n[23318];
assign t[23319] = t[23318] ^ n[23319];
assign t[23320] = t[23319] ^ n[23320];
assign t[23321] = t[23320] ^ n[23321];
assign t[23322] = t[23321] ^ n[23322];
assign t[23323] = t[23322] ^ n[23323];
assign t[23324] = t[23323] ^ n[23324];
assign t[23325] = t[23324] ^ n[23325];
assign t[23326] = t[23325] ^ n[23326];
assign t[23327] = t[23326] ^ n[23327];
assign t[23328] = t[23327] ^ n[23328];
assign t[23329] = t[23328] ^ n[23329];
assign t[23330] = t[23329] ^ n[23330];
assign t[23331] = t[23330] ^ n[23331];
assign t[23332] = t[23331] ^ n[23332];
assign t[23333] = t[23332] ^ n[23333];
assign t[23334] = t[23333] ^ n[23334];
assign t[23335] = t[23334] ^ n[23335];
assign t[23336] = t[23335] ^ n[23336];
assign t[23337] = t[23336] ^ n[23337];
assign t[23338] = t[23337] ^ n[23338];
assign t[23339] = t[23338] ^ n[23339];
assign t[23340] = t[23339] ^ n[23340];
assign t[23341] = t[23340] ^ n[23341];
assign t[23342] = t[23341] ^ n[23342];
assign t[23343] = t[23342] ^ n[23343];
assign t[23344] = t[23343] ^ n[23344];
assign t[23345] = t[23344] ^ n[23345];
assign t[23346] = t[23345] ^ n[23346];
assign t[23347] = t[23346] ^ n[23347];
assign t[23348] = t[23347] ^ n[23348];
assign t[23349] = t[23348] ^ n[23349];
assign t[23350] = t[23349] ^ n[23350];
assign t[23351] = t[23350] ^ n[23351];
assign t[23352] = t[23351] ^ n[23352];
assign t[23353] = t[23352] ^ n[23353];
assign t[23354] = t[23353] ^ n[23354];
assign t[23355] = t[23354] ^ n[23355];
assign t[23356] = t[23355] ^ n[23356];
assign t[23357] = t[23356] ^ n[23357];
assign t[23358] = t[23357] ^ n[23358];
assign t[23359] = t[23358] ^ n[23359];
assign t[23360] = t[23359] ^ n[23360];
assign t[23361] = t[23360] ^ n[23361];
assign t[23362] = t[23361] ^ n[23362];
assign t[23363] = t[23362] ^ n[23363];
assign t[23364] = t[23363] ^ n[23364];
assign t[23365] = t[23364] ^ n[23365];
assign t[23366] = t[23365] ^ n[23366];
assign t[23367] = t[23366] ^ n[23367];
assign t[23368] = t[23367] ^ n[23368];
assign t[23369] = t[23368] ^ n[23369];
assign t[23370] = t[23369] ^ n[23370];
assign t[23371] = t[23370] ^ n[23371];
assign t[23372] = t[23371] ^ n[23372];
assign t[23373] = t[23372] ^ n[23373];
assign t[23374] = t[23373] ^ n[23374];
assign t[23375] = t[23374] ^ n[23375];
assign t[23376] = t[23375] ^ n[23376];
assign t[23377] = t[23376] ^ n[23377];
assign t[23378] = t[23377] ^ n[23378];
assign t[23379] = t[23378] ^ n[23379];
assign t[23380] = t[23379] ^ n[23380];
assign t[23381] = t[23380] ^ n[23381];
assign t[23382] = t[23381] ^ n[23382];
assign t[23383] = t[23382] ^ n[23383];
assign t[23384] = t[23383] ^ n[23384];
assign t[23385] = t[23384] ^ n[23385];
assign t[23386] = t[23385] ^ n[23386];
assign t[23387] = t[23386] ^ n[23387];
assign t[23388] = t[23387] ^ n[23388];
assign t[23389] = t[23388] ^ n[23389];
assign t[23390] = t[23389] ^ n[23390];
assign t[23391] = t[23390] ^ n[23391];
assign t[23392] = t[23391] ^ n[23392];
assign t[23393] = t[23392] ^ n[23393];
assign t[23394] = t[23393] ^ n[23394];
assign t[23395] = t[23394] ^ n[23395];
assign t[23396] = t[23395] ^ n[23396];
assign t[23397] = t[23396] ^ n[23397];
assign t[23398] = t[23397] ^ n[23398];
assign t[23399] = t[23398] ^ n[23399];
assign t[23400] = t[23399] ^ n[23400];
assign t[23401] = t[23400] ^ n[23401];
assign t[23402] = t[23401] ^ n[23402];
assign t[23403] = t[23402] ^ n[23403];
assign t[23404] = t[23403] ^ n[23404];
assign t[23405] = t[23404] ^ n[23405];
assign t[23406] = t[23405] ^ n[23406];
assign t[23407] = t[23406] ^ n[23407];
assign t[23408] = t[23407] ^ n[23408];
assign t[23409] = t[23408] ^ n[23409];
assign t[23410] = t[23409] ^ n[23410];
assign t[23411] = t[23410] ^ n[23411];
assign t[23412] = t[23411] ^ n[23412];
assign t[23413] = t[23412] ^ n[23413];
assign t[23414] = t[23413] ^ n[23414];
assign t[23415] = t[23414] ^ n[23415];
assign t[23416] = t[23415] ^ n[23416];
assign t[23417] = t[23416] ^ n[23417];
assign t[23418] = t[23417] ^ n[23418];
assign t[23419] = t[23418] ^ n[23419];
assign t[23420] = t[23419] ^ n[23420];
assign t[23421] = t[23420] ^ n[23421];
assign t[23422] = t[23421] ^ n[23422];
assign t[23423] = t[23422] ^ n[23423];
assign t[23424] = t[23423] ^ n[23424];
assign t[23425] = t[23424] ^ n[23425];
assign t[23426] = t[23425] ^ n[23426];
assign t[23427] = t[23426] ^ n[23427];
assign t[23428] = t[23427] ^ n[23428];
assign t[23429] = t[23428] ^ n[23429];
assign t[23430] = t[23429] ^ n[23430];
assign t[23431] = t[23430] ^ n[23431];
assign t[23432] = t[23431] ^ n[23432];
assign t[23433] = t[23432] ^ n[23433];
assign t[23434] = t[23433] ^ n[23434];
assign t[23435] = t[23434] ^ n[23435];
assign t[23436] = t[23435] ^ n[23436];
assign t[23437] = t[23436] ^ n[23437];
assign t[23438] = t[23437] ^ n[23438];
assign t[23439] = t[23438] ^ n[23439];
assign t[23440] = t[23439] ^ n[23440];
assign t[23441] = t[23440] ^ n[23441];
assign t[23442] = t[23441] ^ n[23442];
assign t[23443] = t[23442] ^ n[23443];
assign t[23444] = t[23443] ^ n[23444];
assign t[23445] = t[23444] ^ n[23445];
assign t[23446] = t[23445] ^ n[23446];
assign t[23447] = t[23446] ^ n[23447];
assign t[23448] = t[23447] ^ n[23448];
assign t[23449] = t[23448] ^ n[23449];
assign t[23450] = t[23449] ^ n[23450];
assign t[23451] = t[23450] ^ n[23451];
assign t[23452] = t[23451] ^ n[23452];
assign t[23453] = t[23452] ^ n[23453];
assign t[23454] = t[23453] ^ n[23454];
assign t[23455] = t[23454] ^ n[23455];
assign t[23456] = t[23455] ^ n[23456];
assign t[23457] = t[23456] ^ n[23457];
assign t[23458] = t[23457] ^ n[23458];
assign t[23459] = t[23458] ^ n[23459];
assign t[23460] = t[23459] ^ n[23460];
assign t[23461] = t[23460] ^ n[23461];
assign t[23462] = t[23461] ^ n[23462];
assign t[23463] = t[23462] ^ n[23463];
assign t[23464] = t[23463] ^ n[23464];
assign t[23465] = t[23464] ^ n[23465];
assign t[23466] = t[23465] ^ n[23466];
assign t[23467] = t[23466] ^ n[23467];
assign t[23468] = t[23467] ^ n[23468];
assign t[23469] = t[23468] ^ n[23469];
assign t[23470] = t[23469] ^ n[23470];
assign t[23471] = t[23470] ^ n[23471];
assign t[23472] = t[23471] ^ n[23472];
assign t[23473] = t[23472] ^ n[23473];
assign t[23474] = t[23473] ^ n[23474];
assign t[23475] = t[23474] ^ n[23475];
assign t[23476] = t[23475] ^ n[23476];
assign t[23477] = t[23476] ^ n[23477];
assign t[23478] = t[23477] ^ n[23478];
assign t[23479] = t[23478] ^ n[23479];
assign t[23480] = t[23479] ^ n[23480];
assign t[23481] = t[23480] ^ n[23481];
assign t[23482] = t[23481] ^ n[23482];
assign t[23483] = t[23482] ^ n[23483];
assign t[23484] = t[23483] ^ n[23484];
assign t[23485] = t[23484] ^ n[23485];
assign t[23486] = t[23485] ^ n[23486];
assign t[23487] = t[23486] ^ n[23487];
assign t[23488] = t[23487] ^ n[23488];
assign t[23489] = t[23488] ^ n[23489];
assign t[23490] = t[23489] ^ n[23490];
assign t[23491] = t[23490] ^ n[23491];
assign t[23492] = t[23491] ^ n[23492];
assign t[23493] = t[23492] ^ n[23493];
assign t[23494] = t[23493] ^ n[23494];
assign t[23495] = t[23494] ^ n[23495];
assign t[23496] = t[23495] ^ n[23496];
assign t[23497] = t[23496] ^ n[23497];
assign t[23498] = t[23497] ^ n[23498];
assign t[23499] = t[23498] ^ n[23499];
assign t[23500] = t[23499] ^ n[23500];
assign t[23501] = t[23500] ^ n[23501];
assign t[23502] = t[23501] ^ n[23502];
assign t[23503] = t[23502] ^ n[23503];
assign t[23504] = t[23503] ^ n[23504];
assign t[23505] = t[23504] ^ n[23505];
assign t[23506] = t[23505] ^ n[23506];
assign t[23507] = t[23506] ^ n[23507];
assign t[23508] = t[23507] ^ n[23508];
assign t[23509] = t[23508] ^ n[23509];
assign t[23510] = t[23509] ^ n[23510];
assign t[23511] = t[23510] ^ n[23511];
assign t[23512] = t[23511] ^ n[23512];
assign t[23513] = t[23512] ^ n[23513];
assign t[23514] = t[23513] ^ n[23514];
assign t[23515] = t[23514] ^ n[23515];
assign t[23516] = t[23515] ^ n[23516];
assign t[23517] = t[23516] ^ n[23517];
assign t[23518] = t[23517] ^ n[23518];
assign t[23519] = t[23518] ^ n[23519];
assign t[23520] = t[23519] ^ n[23520];
assign t[23521] = t[23520] ^ n[23521];
assign t[23522] = t[23521] ^ n[23522];
assign t[23523] = t[23522] ^ n[23523];
assign t[23524] = t[23523] ^ n[23524];
assign t[23525] = t[23524] ^ n[23525];
assign t[23526] = t[23525] ^ n[23526];
assign t[23527] = t[23526] ^ n[23527];
assign t[23528] = t[23527] ^ n[23528];
assign t[23529] = t[23528] ^ n[23529];
assign t[23530] = t[23529] ^ n[23530];
assign t[23531] = t[23530] ^ n[23531];
assign t[23532] = t[23531] ^ n[23532];
assign t[23533] = t[23532] ^ n[23533];
assign t[23534] = t[23533] ^ n[23534];
assign t[23535] = t[23534] ^ n[23535];
assign t[23536] = t[23535] ^ n[23536];
assign t[23537] = t[23536] ^ n[23537];
assign t[23538] = t[23537] ^ n[23538];
assign t[23539] = t[23538] ^ n[23539];
assign t[23540] = t[23539] ^ n[23540];
assign t[23541] = t[23540] ^ n[23541];
assign t[23542] = t[23541] ^ n[23542];
assign t[23543] = t[23542] ^ n[23543];
assign t[23544] = t[23543] ^ n[23544];
assign t[23545] = t[23544] ^ n[23545];
assign t[23546] = t[23545] ^ n[23546];
assign t[23547] = t[23546] ^ n[23547];
assign t[23548] = t[23547] ^ n[23548];
assign t[23549] = t[23548] ^ n[23549];
assign t[23550] = t[23549] ^ n[23550];
assign t[23551] = t[23550] ^ n[23551];
assign t[23552] = t[23551] ^ n[23552];
assign t[23553] = t[23552] ^ n[23553];
assign t[23554] = t[23553] ^ n[23554];
assign t[23555] = t[23554] ^ n[23555];
assign t[23556] = t[23555] ^ n[23556];
assign t[23557] = t[23556] ^ n[23557];
assign t[23558] = t[23557] ^ n[23558];
assign t[23559] = t[23558] ^ n[23559];
assign t[23560] = t[23559] ^ n[23560];
assign t[23561] = t[23560] ^ n[23561];
assign t[23562] = t[23561] ^ n[23562];
assign t[23563] = t[23562] ^ n[23563];
assign t[23564] = t[23563] ^ n[23564];
assign t[23565] = t[23564] ^ n[23565];
assign t[23566] = t[23565] ^ n[23566];
assign t[23567] = t[23566] ^ n[23567];
assign t[23568] = t[23567] ^ n[23568];
assign t[23569] = t[23568] ^ n[23569];
assign t[23570] = t[23569] ^ n[23570];
assign t[23571] = t[23570] ^ n[23571];
assign t[23572] = t[23571] ^ n[23572];
assign t[23573] = t[23572] ^ n[23573];
assign t[23574] = t[23573] ^ n[23574];
assign t[23575] = t[23574] ^ n[23575];
assign t[23576] = t[23575] ^ n[23576];
assign t[23577] = t[23576] ^ n[23577];
assign t[23578] = t[23577] ^ n[23578];
assign t[23579] = t[23578] ^ n[23579];
assign t[23580] = t[23579] ^ n[23580];
assign t[23581] = t[23580] ^ n[23581];
assign t[23582] = t[23581] ^ n[23582];
assign t[23583] = t[23582] ^ n[23583];
assign t[23584] = t[23583] ^ n[23584];
assign t[23585] = t[23584] ^ n[23585];
assign t[23586] = t[23585] ^ n[23586];
assign t[23587] = t[23586] ^ n[23587];
assign t[23588] = t[23587] ^ n[23588];
assign t[23589] = t[23588] ^ n[23589];
assign t[23590] = t[23589] ^ n[23590];
assign t[23591] = t[23590] ^ n[23591];
assign t[23592] = t[23591] ^ n[23592];
assign t[23593] = t[23592] ^ n[23593];
assign t[23594] = t[23593] ^ n[23594];
assign t[23595] = t[23594] ^ n[23595];
assign t[23596] = t[23595] ^ n[23596];
assign t[23597] = t[23596] ^ n[23597];
assign t[23598] = t[23597] ^ n[23598];
assign t[23599] = t[23598] ^ n[23599];
assign t[23600] = t[23599] ^ n[23600];
assign t[23601] = t[23600] ^ n[23601];
assign t[23602] = t[23601] ^ n[23602];
assign t[23603] = t[23602] ^ n[23603];
assign t[23604] = t[23603] ^ n[23604];
assign t[23605] = t[23604] ^ n[23605];
assign t[23606] = t[23605] ^ n[23606];
assign t[23607] = t[23606] ^ n[23607];
assign t[23608] = t[23607] ^ n[23608];
assign t[23609] = t[23608] ^ n[23609];
assign t[23610] = t[23609] ^ n[23610];
assign t[23611] = t[23610] ^ n[23611];
assign t[23612] = t[23611] ^ n[23612];
assign t[23613] = t[23612] ^ n[23613];
assign t[23614] = t[23613] ^ n[23614];
assign t[23615] = t[23614] ^ n[23615];
assign t[23616] = t[23615] ^ n[23616];
assign t[23617] = t[23616] ^ n[23617];
assign t[23618] = t[23617] ^ n[23618];
assign t[23619] = t[23618] ^ n[23619];
assign t[23620] = t[23619] ^ n[23620];
assign t[23621] = t[23620] ^ n[23621];
assign t[23622] = t[23621] ^ n[23622];
assign t[23623] = t[23622] ^ n[23623];
assign t[23624] = t[23623] ^ n[23624];
assign t[23625] = t[23624] ^ n[23625];
assign t[23626] = t[23625] ^ n[23626];
assign t[23627] = t[23626] ^ n[23627];
assign t[23628] = t[23627] ^ n[23628];
assign t[23629] = t[23628] ^ n[23629];
assign t[23630] = t[23629] ^ n[23630];
assign t[23631] = t[23630] ^ n[23631];
assign t[23632] = t[23631] ^ n[23632];
assign t[23633] = t[23632] ^ n[23633];
assign t[23634] = t[23633] ^ n[23634];
assign t[23635] = t[23634] ^ n[23635];
assign t[23636] = t[23635] ^ n[23636];
assign t[23637] = t[23636] ^ n[23637];
assign t[23638] = t[23637] ^ n[23638];
assign t[23639] = t[23638] ^ n[23639];
assign t[23640] = t[23639] ^ n[23640];
assign t[23641] = t[23640] ^ n[23641];
assign t[23642] = t[23641] ^ n[23642];
assign t[23643] = t[23642] ^ n[23643];
assign t[23644] = t[23643] ^ n[23644];
assign t[23645] = t[23644] ^ n[23645];
assign t[23646] = t[23645] ^ n[23646];
assign t[23647] = t[23646] ^ n[23647];
assign t[23648] = t[23647] ^ n[23648];
assign t[23649] = t[23648] ^ n[23649];
assign t[23650] = t[23649] ^ n[23650];
assign t[23651] = t[23650] ^ n[23651];
assign t[23652] = t[23651] ^ n[23652];
assign t[23653] = t[23652] ^ n[23653];
assign t[23654] = t[23653] ^ n[23654];
assign t[23655] = t[23654] ^ n[23655];
assign t[23656] = t[23655] ^ n[23656];
assign t[23657] = t[23656] ^ n[23657];
assign t[23658] = t[23657] ^ n[23658];
assign t[23659] = t[23658] ^ n[23659];
assign t[23660] = t[23659] ^ n[23660];
assign t[23661] = t[23660] ^ n[23661];
assign t[23662] = t[23661] ^ n[23662];
assign t[23663] = t[23662] ^ n[23663];
assign t[23664] = t[23663] ^ n[23664];
assign t[23665] = t[23664] ^ n[23665];
assign t[23666] = t[23665] ^ n[23666];
assign t[23667] = t[23666] ^ n[23667];
assign t[23668] = t[23667] ^ n[23668];
assign t[23669] = t[23668] ^ n[23669];
assign t[23670] = t[23669] ^ n[23670];
assign t[23671] = t[23670] ^ n[23671];
assign t[23672] = t[23671] ^ n[23672];
assign t[23673] = t[23672] ^ n[23673];
assign t[23674] = t[23673] ^ n[23674];
assign t[23675] = t[23674] ^ n[23675];
assign t[23676] = t[23675] ^ n[23676];
assign t[23677] = t[23676] ^ n[23677];
assign t[23678] = t[23677] ^ n[23678];
assign t[23679] = t[23678] ^ n[23679];
assign t[23680] = t[23679] ^ n[23680];
assign t[23681] = t[23680] ^ n[23681];
assign t[23682] = t[23681] ^ n[23682];
assign t[23683] = t[23682] ^ n[23683];
assign t[23684] = t[23683] ^ n[23684];
assign t[23685] = t[23684] ^ n[23685];
assign t[23686] = t[23685] ^ n[23686];
assign t[23687] = t[23686] ^ n[23687];
assign t[23688] = t[23687] ^ n[23688];
assign t[23689] = t[23688] ^ n[23689];
assign t[23690] = t[23689] ^ n[23690];
assign t[23691] = t[23690] ^ n[23691];
assign t[23692] = t[23691] ^ n[23692];
assign t[23693] = t[23692] ^ n[23693];
assign t[23694] = t[23693] ^ n[23694];
assign t[23695] = t[23694] ^ n[23695];
assign t[23696] = t[23695] ^ n[23696];
assign t[23697] = t[23696] ^ n[23697];
assign t[23698] = t[23697] ^ n[23698];
assign t[23699] = t[23698] ^ n[23699];
assign t[23700] = t[23699] ^ n[23700];
assign t[23701] = t[23700] ^ n[23701];
assign t[23702] = t[23701] ^ n[23702];
assign t[23703] = t[23702] ^ n[23703];
assign t[23704] = t[23703] ^ n[23704];
assign t[23705] = t[23704] ^ n[23705];
assign t[23706] = t[23705] ^ n[23706];
assign t[23707] = t[23706] ^ n[23707];
assign t[23708] = t[23707] ^ n[23708];
assign t[23709] = t[23708] ^ n[23709];
assign t[23710] = t[23709] ^ n[23710];
assign t[23711] = t[23710] ^ n[23711];
assign t[23712] = t[23711] ^ n[23712];
assign t[23713] = t[23712] ^ n[23713];
assign t[23714] = t[23713] ^ n[23714];
assign t[23715] = t[23714] ^ n[23715];
assign t[23716] = t[23715] ^ n[23716];
assign t[23717] = t[23716] ^ n[23717];
assign t[23718] = t[23717] ^ n[23718];
assign t[23719] = t[23718] ^ n[23719];
assign t[23720] = t[23719] ^ n[23720];
assign t[23721] = t[23720] ^ n[23721];
assign t[23722] = t[23721] ^ n[23722];
assign t[23723] = t[23722] ^ n[23723];
assign t[23724] = t[23723] ^ n[23724];
assign t[23725] = t[23724] ^ n[23725];
assign t[23726] = t[23725] ^ n[23726];
assign t[23727] = t[23726] ^ n[23727];
assign t[23728] = t[23727] ^ n[23728];
assign t[23729] = t[23728] ^ n[23729];
assign t[23730] = t[23729] ^ n[23730];
assign t[23731] = t[23730] ^ n[23731];
assign t[23732] = t[23731] ^ n[23732];
assign t[23733] = t[23732] ^ n[23733];
assign t[23734] = t[23733] ^ n[23734];
assign t[23735] = t[23734] ^ n[23735];
assign t[23736] = t[23735] ^ n[23736];
assign t[23737] = t[23736] ^ n[23737];
assign t[23738] = t[23737] ^ n[23738];
assign t[23739] = t[23738] ^ n[23739];
assign t[23740] = t[23739] ^ n[23740];
assign t[23741] = t[23740] ^ n[23741];
assign t[23742] = t[23741] ^ n[23742];
assign t[23743] = t[23742] ^ n[23743];
assign t[23744] = t[23743] ^ n[23744];
assign t[23745] = t[23744] ^ n[23745];
assign t[23746] = t[23745] ^ n[23746];
assign t[23747] = t[23746] ^ n[23747];
assign t[23748] = t[23747] ^ n[23748];
assign t[23749] = t[23748] ^ n[23749];
assign t[23750] = t[23749] ^ n[23750];
assign t[23751] = t[23750] ^ n[23751];
assign t[23752] = t[23751] ^ n[23752];
assign t[23753] = t[23752] ^ n[23753];
assign t[23754] = t[23753] ^ n[23754];
assign t[23755] = t[23754] ^ n[23755];
assign t[23756] = t[23755] ^ n[23756];
assign t[23757] = t[23756] ^ n[23757];
assign t[23758] = t[23757] ^ n[23758];
assign t[23759] = t[23758] ^ n[23759];
assign t[23760] = t[23759] ^ n[23760];
assign t[23761] = t[23760] ^ n[23761];
assign t[23762] = t[23761] ^ n[23762];
assign t[23763] = t[23762] ^ n[23763];
assign t[23764] = t[23763] ^ n[23764];
assign t[23765] = t[23764] ^ n[23765];
assign t[23766] = t[23765] ^ n[23766];
assign t[23767] = t[23766] ^ n[23767];
assign t[23768] = t[23767] ^ n[23768];
assign t[23769] = t[23768] ^ n[23769];
assign t[23770] = t[23769] ^ n[23770];
assign t[23771] = t[23770] ^ n[23771];
assign t[23772] = t[23771] ^ n[23772];
assign t[23773] = t[23772] ^ n[23773];
assign t[23774] = t[23773] ^ n[23774];
assign t[23775] = t[23774] ^ n[23775];
assign t[23776] = t[23775] ^ n[23776];
assign t[23777] = t[23776] ^ n[23777];
assign t[23778] = t[23777] ^ n[23778];
assign t[23779] = t[23778] ^ n[23779];
assign t[23780] = t[23779] ^ n[23780];
assign t[23781] = t[23780] ^ n[23781];
assign t[23782] = t[23781] ^ n[23782];
assign t[23783] = t[23782] ^ n[23783];
assign t[23784] = t[23783] ^ n[23784];
assign t[23785] = t[23784] ^ n[23785];
assign t[23786] = t[23785] ^ n[23786];
assign t[23787] = t[23786] ^ n[23787];
assign t[23788] = t[23787] ^ n[23788];
assign t[23789] = t[23788] ^ n[23789];
assign t[23790] = t[23789] ^ n[23790];
assign t[23791] = t[23790] ^ n[23791];
assign t[23792] = t[23791] ^ n[23792];
assign t[23793] = t[23792] ^ n[23793];
assign t[23794] = t[23793] ^ n[23794];
assign t[23795] = t[23794] ^ n[23795];
assign t[23796] = t[23795] ^ n[23796];
assign t[23797] = t[23796] ^ n[23797];
assign t[23798] = t[23797] ^ n[23798];
assign t[23799] = t[23798] ^ n[23799];
assign t[23800] = t[23799] ^ n[23800];
assign t[23801] = t[23800] ^ n[23801];
assign t[23802] = t[23801] ^ n[23802];
assign t[23803] = t[23802] ^ n[23803];
assign t[23804] = t[23803] ^ n[23804];
assign t[23805] = t[23804] ^ n[23805];
assign t[23806] = t[23805] ^ n[23806];
assign t[23807] = t[23806] ^ n[23807];
assign t[23808] = t[23807] ^ n[23808];
assign t[23809] = t[23808] ^ n[23809];
assign t[23810] = t[23809] ^ n[23810];
assign t[23811] = t[23810] ^ n[23811];
assign t[23812] = t[23811] ^ n[23812];
assign t[23813] = t[23812] ^ n[23813];
assign t[23814] = t[23813] ^ n[23814];
assign t[23815] = t[23814] ^ n[23815];
assign t[23816] = t[23815] ^ n[23816];
assign t[23817] = t[23816] ^ n[23817];
assign t[23818] = t[23817] ^ n[23818];
assign t[23819] = t[23818] ^ n[23819];
assign t[23820] = t[23819] ^ n[23820];
assign t[23821] = t[23820] ^ n[23821];
assign t[23822] = t[23821] ^ n[23822];
assign t[23823] = t[23822] ^ n[23823];
assign t[23824] = t[23823] ^ n[23824];
assign t[23825] = t[23824] ^ n[23825];
assign t[23826] = t[23825] ^ n[23826];
assign t[23827] = t[23826] ^ n[23827];
assign t[23828] = t[23827] ^ n[23828];
assign t[23829] = t[23828] ^ n[23829];
assign t[23830] = t[23829] ^ n[23830];
assign t[23831] = t[23830] ^ n[23831];
assign t[23832] = t[23831] ^ n[23832];
assign t[23833] = t[23832] ^ n[23833];
assign t[23834] = t[23833] ^ n[23834];
assign t[23835] = t[23834] ^ n[23835];
assign t[23836] = t[23835] ^ n[23836];
assign t[23837] = t[23836] ^ n[23837];
assign t[23838] = t[23837] ^ n[23838];
assign t[23839] = t[23838] ^ n[23839];
assign t[23840] = t[23839] ^ n[23840];
assign t[23841] = t[23840] ^ n[23841];
assign t[23842] = t[23841] ^ n[23842];
assign t[23843] = t[23842] ^ n[23843];
assign t[23844] = t[23843] ^ n[23844];
assign t[23845] = t[23844] ^ n[23845];
assign t[23846] = t[23845] ^ n[23846];
assign t[23847] = t[23846] ^ n[23847];
assign t[23848] = t[23847] ^ n[23848];
assign t[23849] = t[23848] ^ n[23849];
assign t[23850] = t[23849] ^ n[23850];
assign t[23851] = t[23850] ^ n[23851];
assign t[23852] = t[23851] ^ n[23852];
assign t[23853] = t[23852] ^ n[23853];
assign t[23854] = t[23853] ^ n[23854];
assign t[23855] = t[23854] ^ n[23855];
assign t[23856] = t[23855] ^ n[23856];
assign t[23857] = t[23856] ^ n[23857];
assign t[23858] = t[23857] ^ n[23858];
assign t[23859] = t[23858] ^ n[23859];
assign t[23860] = t[23859] ^ n[23860];
assign t[23861] = t[23860] ^ n[23861];
assign t[23862] = t[23861] ^ n[23862];
assign t[23863] = t[23862] ^ n[23863];
assign t[23864] = t[23863] ^ n[23864];
assign t[23865] = t[23864] ^ n[23865];
assign t[23866] = t[23865] ^ n[23866];
assign t[23867] = t[23866] ^ n[23867];
assign t[23868] = t[23867] ^ n[23868];
assign t[23869] = t[23868] ^ n[23869];
assign t[23870] = t[23869] ^ n[23870];
assign t[23871] = t[23870] ^ n[23871];
assign t[23872] = t[23871] ^ n[23872];
assign t[23873] = t[23872] ^ n[23873];
assign t[23874] = t[23873] ^ n[23874];
assign t[23875] = t[23874] ^ n[23875];
assign t[23876] = t[23875] ^ n[23876];
assign t[23877] = t[23876] ^ n[23877];
assign t[23878] = t[23877] ^ n[23878];
assign t[23879] = t[23878] ^ n[23879];
assign t[23880] = t[23879] ^ n[23880];
assign t[23881] = t[23880] ^ n[23881];
assign t[23882] = t[23881] ^ n[23882];
assign t[23883] = t[23882] ^ n[23883];
assign t[23884] = t[23883] ^ n[23884];
assign t[23885] = t[23884] ^ n[23885];
assign t[23886] = t[23885] ^ n[23886];
assign t[23887] = t[23886] ^ n[23887];
assign t[23888] = t[23887] ^ n[23888];
assign t[23889] = t[23888] ^ n[23889];
assign t[23890] = t[23889] ^ n[23890];
assign t[23891] = t[23890] ^ n[23891];
assign t[23892] = t[23891] ^ n[23892];
assign t[23893] = t[23892] ^ n[23893];
assign t[23894] = t[23893] ^ n[23894];
assign t[23895] = t[23894] ^ n[23895];
assign t[23896] = t[23895] ^ n[23896];
assign t[23897] = t[23896] ^ n[23897];
assign t[23898] = t[23897] ^ n[23898];
assign t[23899] = t[23898] ^ n[23899];
assign t[23900] = t[23899] ^ n[23900];
assign t[23901] = t[23900] ^ n[23901];
assign t[23902] = t[23901] ^ n[23902];
assign t[23903] = t[23902] ^ n[23903];
assign t[23904] = t[23903] ^ n[23904];
assign t[23905] = t[23904] ^ n[23905];
assign t[23906] = t[23905] ^ n[23906];
assign t[23907] = t[23906] ^ n[23907];
assign t[23908] = t[23907] ^ n[23908];
assign t[23909] = t[23908] ^ n[23909];
assign t[23910] = t[23909] ^ n[23910];
assign t[23911] = t[23910] ^ n[23911];
assign t[23912] = t[23911] ^ n[23912];
assign t[23913] = t[23912] ^ n[23913];
assign t[23914] = t[23913] ^ n[23914];
assign t[23915] = t[23914] ^ n[23915];
assign t[23916] = t[23915] ^ n[23916];
assign t[23917] = t[23916] ^ n[23917];
assign t[23918] = t[23917] ^ n[23918];
assign t[23919] = t[23918] ^ n[23919];
assign t[23920] = t[23919] ^ n[23920];
assign t[23921] = t[23920] ^ n[23921];
assign t[23922] = t[23921] ^ n[23922];
assign t[23923] = t[23922] ^ n[23923];
assign t[23924] = t[23923] ^ n[23924];
assign t[23925] = t[23924] ^ n[23925];
assign t[23926] = t[23925] ^ n[23926];
assign t[23927] = t[23926] ^ n[23927];
assign t[23928] = t[23927] ^ n[23928];
assign t[23929] = t[23928] ^ n[23929];
assign t[23930] = t[23929] ^ n[23930];
assign t[23931] = t[23930] ^ n[23931];
assign t[23932] = t[23931] ^ n[23932];
assign t[23933] = t[23932] ^ n[23933];
assign t[23934] = t[23933] ^ n[23934];
assign t[23935] = t[23934] ^ n[23935];
assign t[23936] = t[23935] ^ n[23936];
assign t[23937] = t[23936] ^ n[23937];
assign t[23938] = t[23937] ^ n[23938];
assign t[23939] = t[23938] ^ n[23939];
assign t[23940] = t[23939] ^ n[23940];
assign t[23941] = t[23940] ^ n[23941];
assign t[23942] = t[23941] ^ n[23942];
assign t[23943] = t[23942] ^ n[23943];
assign t[23944] = t[23943] ^ n[23944];
assign t[23945] = t[23944] ^ n[23945];
assign t[23946] = t[23945] ^ n[23946];
assign t[23947] = t[23946] ^ n[23947];
assign t[23948] = t[23947] ^ n[23948];
assign t[23949] = t[23948] ^ n[23949];
assign t[23950] = t[23949] ^ n[23950];
assign t[23951] = t[23950] ^ n[23951];
assign t[23952] = t[23951] ^ n[23952];
assign t[23953] = t[23952] ^ n[23953];
assign t[23954] = t[23953] ^ n[23954];
assign t[23955] = t[23954] ^ n[23955];
assign t[23956] = t[23955] ^ n[23956];
assign t[23957] = t[23956] ^ n[23957];
assign t[23958] = t[23957] ^ n[23958];
assign t[23959] = t[23958] ^ n[23959];
assign t[23960] = t[23959] ^ n[23960];
assign t[23961] = t[23960] ^ n[23961];
assign t[23962] = t[23961] ^ n[23962];
assign t[23963] = t[23962] ^ n[23963];
assign t[23964] = t[23963] ^ n[23964];
assign t[23965] = t[23964] ^ n[23965];
assign t[23966] = t[23965] ^ n[23966];
assign t[23967] = t[23966] ^ n[23967];
assign t[23968] = t[23967] ^ n[23968];
assign t[23969] = t[23968] ^ n[23969];
assign t[23970] = t[23969] ^ n[23970];
assign t[23971] = t[23970] ^ n[23971];
assign t[23972] = t[23971] ^ n[23972];
assign t[23973] = t[23972] ^ n[23973];
assign t[23974] = t[23973] ^ n[23974];
assign t[23975] = t[23974] ^ n[23975];
assign t[23976] = t[23975] ^ n[23976];
assign t[23977] = t[23976] ^ n[23977];
assign t[23978] = t[23977] ^ n[23978];
assign t[23979] = t[23978] ^ n[23979];
assign t[23980] = t[23979] ^ n[23980];
assign t[23981] = t[23980] ^ n[23981];
assign t[23982] = t[23981] ^ n[23982];
assign t[23983] = t[23982] ^ n[23983];
assign t[23984] = t[23983] ^ n[23984];
assign t[23985] = t[23984] ^ n[23985];
assign t[23986] = t[23985] ^ n[23986];
assign t[23987] = t[23986] ^ n[23987];
assign t[23988] = t[23987] ^ n[23988];
assign t[23989] = t[23988] ^ n[23989];
assign t[23990] = t[23989] ^ n[23990];
assign t[23991] = t[23990] ^ n[23991];
assign t[23992] = t[23991] ^ n[23992];
assign t[23993] = t[23992] ^ n[23993];
assign t[23994] = t[23993] ^ n[23994];
assign t[23995] = t[23994] ^ n[23995];
assign t[23996] = t[23995] ^ n[23996];
assign t[23997] = t[23996] ^ n[23997];
assign t[23998] = t[23997] ^ n[23998];
assign t[23999] = t[23998] ^ n[23999];
assign t[24000] = t[23999] ^ n[24000];
assign t[24001] = t[24000] ^ n[24001];
assign t[24002] = t[24001] ^ n[24002];
assign t[24003] = t[24002] ^ n[24003];
assign t[24004] = t[24003] ^ n[24004];
assign t[24005] = t[24004] ^ n[24005];
assign t[24006] = t[24005] ^ n[24006];
assign t[24007] = t[24006] ^ n[24007];
assign t[24008] = t[24007] ^ n[24008];
assign t[24009] = t[24008] ^ n[24009];
assign t[24010] = t[24009] ^ n[24010];
assign t[24011] = t[24010] ^ n[24011];
assign t[24012] = t[24011] ^ n[24012];
assign t[24013] = t[24012] ^ n[24013];
assign t[24014] = t[24013] ^ n[24014];
assign t[24015] = t[24014] ^ n[24015];
assign t[24016] = t[24015] ^ n[24016];
assign t[24017] = t[24016] ^ n[24017];
assign t[24018] = t[24017] ^ n[24018];
assign t[24019] = t[24018] ^ n[24019];
assign t[24020] = t[24019] ^ n[24020];
assign t[24021] = t[24020] ^ n[24021];
assign t[24022] = t[24021] ^ n[24022];
assign t[24023] = t[24022] ^ n[24023];
assign t[24024] = t[24023] ^ n[24024];
assign t[24025] = t[24024] ^ n[24025];
assign t[24026] = t[24025] ^ n[24026];
assign t[24027] = t[24026] ^ n[24027];
assign t[24028] = t[24027] ^ n[24028];
assign t[24029] = t[24028] ^ n[24029];
assign t[24030] = t[24029] ^ n[24030];
assign t[24031] = t[24030] ^ n[24031];
assign t[24032] = t[24031] ^ n[24032];
assign t[24033] = t[24032] ^ n[24033];
assign t[24034] = t[24033] ^ n[24034];
assign t[24035] = t[24034] ^ n[24035];
assign t[24036] = t[24035] ^ n[24036];
assign t[24037] = t[24036] ^ n[24037];
assign t[24038] = t[24037] ^ n[24038];
assign t[24039] = t[24038] ^ n[24039];
assign t[24040] = t[24039] ^ n[24040];
assign t[24041] = t[24040] ^ n[24041];
assign t[24042] = t[24041] ^ n[24042];
assign t[24043] = t[24042] ^ n[24043];
assign t[24044] = t[24043] ^ n[24044];
assign t[24045] = t[24044] ^ n[24045];
assign t[24046] = t[24045] ^ n[24046];
assign t[24047] = t[24046] ^ n[24047];
assign t[24048] = t[24047] ^ n[24048];
assign t[24049] = t[24048] ^ n[24049];
assign t[24050] = t[24049] ^ n[24050];
assign t[24051] = t[24050] ^ n[24051];
assign t[24052] = t[24051] ^ n[24052];
assign t[24053] = t[24052] ^ n[24053];
assign t[24054] = t[24053] ^ n[24054];
assign t[24055] = t[24054] ^ n[24055];
assign t[24056] = t[24055] ^ n[24056];
assign t[24057] = t[24056] ^ n[24057];
assign t[24058] = t[24057] ^ n[24058];
assign t[24059] = t[24058] ^ n[24059];
assign t[24060] = t[24059] ^ n[24060];
assign t[24061] = t[24060] ^ n[24061];
assign t[24062] = t[24061] ^ n[24062];
assign t[24063] = t[24062] ^ n[24063];
assign t[24064] = t[24063] ^ n[24064];
assign t[24065] = t[24064] ^ n[24065];
assign t[24066] = t[24065] ^ n[24066];
assign t[24067] = t[24066] ^ n[24067];
assign t[24068] = t[24067] ^ n[24068];
assign t[24069] = t[24068] ^ n[24069];
assign t[24070] = t[24069] ^ n[24070];
assign t[24071] = t[24070] ^ n[24071];
assign t[24072] = t[24071] ^ n[24072];
assign t[24073] = t[24072] ^ n[24073];
assign t[24074] = t[24073] ^ n[24074];
assign t[24075] = t[24074] ^ n[24075];
assign t[24076] = t[24075] ^ n[24076];
assign t[24077] = t[24076] ^ n[24077];
assign t[24078] = t[24077] ^ n[24078];
assign t[24079] = t[24078] ^ n[24079];
assign t[24080] = t[24079] ^ n[24080];
assign t[24081] = t[24080] ^ n[24081];
assign t[24082] = t[24081] ^ n[24082];
assign t[24083] = t[24082] ^ n[24083];
assign t[24084] = t[24083] ^ n[24084];
assign t[24085] = t[24084] ^ n[24085];
assign t[24086] = t[24085] ^ n[24086];
assign t[24087] = t[24086] ^ n[24087];
assign t[24088] = t[24087] ^ n[24088];
assign t[24089] = t[24088] ^ n[24089];
assign t[24090] = t[24089] ^ n[24090];
assign t[24091] = t[24090] ^ n[24091];
assign t[24092] = t[24091] ^ n[24092];
assign t[24093] = t[24092] ^ n[24093];
assign t[24094] = t[24093] ^ n[24094];
assign t[24095] = t[24094] ^ n[24095];
assign t[24096] = t[24095] ^ n[24096];
assign t[24097] = t[24096] ^ n[24097];
assign t[24098] = t[24097] ^ n[24098];
assign t[24099] = t[24098] ^ n[24099];
assign t[24100] = t[24099] ^ n[24100];
assign t[24101] = t[24100] ^ n[24101];
assign t[24102] = t[24101] ^ n[24102];
assign t[24103] = t[24102] ^ n[24103];
assign t[24104] = t[24103] ^ n[24104];
assign t[24105] = t[24104] ^ n[24105];
assign t[24106] = t[24105] ^ n[24106];
assign t[24107] = t[24106] ^ n[24107];
assign t[24108] = t[24107] ^ n[24108];
assign t[24109] = t[24108] ^ n[24109];
assign t[24110] = t[24109] ^ n[24110];
assign t[24111] = t[24110] ^ n[24111];
assign t[24112] = t[24111] ^ n[24112];
assign t[24113] = t[24112] ^ n[24113];
assign t[24114] = t[24113] ^ n[24114];
assign t[24115] = t[24114] ^ n[24115];
assign t[24116] = t[24115] ^ n[24116];
assign t[24117] = t[24116] ^ n[24117];
assign t[24118] = t[24117] ^ n[24118];
assign t[24119] = t[24118] ^ n[24119];
assign t[24120] = t[24119] ^ n[24120];
assign t[24121] = t[24120] ^ n[24121];
assign t[24122] = t[24121] ^ n[24122];
assign t[24123] = t[24122] ^ n[24123];
assign t[24124] = t[24123] ^ n[24124];
assign t[24125] = t[24124] ^ n[24125];
assign t[24126] = t[24125] ^ n[24126];
assign t[24127] = t[24126] ^ n[24127];
assign t[24128] = t[24127] ^ n[24128];
assign t[24129] = t[24128] ^ n[24129];
assign t[24130] = t[24129] ^ n[24130];
assign t[24131] = t[24130] ^ n[24131];
assign t[24132] = t[24131] ^ n[24132];
assign t[24133] = t[24132] ^ n[24133];
assign t[24134] = t[24133] ^ n[24134];
assign t[24135] = t[24134] ^ n[24135];
assign t[24136] = t[24135] ^ n[24136];
assign t[24137] = t[24136] ^ n[24137];
assign t[24138] = t[24137] ^ n[24138];
assign t[24139] = t[24138] ^ n[24139];
assign t[24140] = t[24139] ^ n[24140];
assign t[24141] = t[24140] ^ n[24141];
assign t[24142] = t[24141] ^ n[24142];
assign t[24143] = t[24142] ^ n[24143];
assign t[24144] = t[24143] ^ n[24144];
assign t[24145] = t[24144] ^ n[24145];
assign t[24146] = t[24145] ^ n[24146];
assign t[24147] = t[24146] ^ n[24147];
assign t[24148] = t[24147] ^ n[24148];
assign t[24149] = t[24148] ^ n[24149];
assign t[24150] = t[24149] ^ n[24150];
assign t[24151] = t[24150] ^ n[24151];
assign t[24152] = t[24151] ^ n[24152];
assign t[24153] = t[24152] ^ n[24153];
assign t[24154] = t[24153] ^ n[24154];
assign t[24155] = t[24154] ^ n[24155];
assign t[24156] = t[24155] ^ n[24156];
assign t[24157] = t[24156] ^ n[24157];
assign t[24158] = t[24157] ^ n[24158];
assign t[24159] = t[24158] ^ n[24159];
assign t[24160] = t[24159] ^ n[24160];
assign t[24161] = t[24160] ^ n[24161];
assign t[24162] = t[24161] ^ n[24162];
assign t[24163] = t[24162] ^ n[24163];
assign t[24164] = t[24163] ^ n[24164];
assign t[24165] = t[24164] ^ n[24165];
assign t[24166] = t[24165] ^ n[24166];
assign t[24167] = t[24166] ^ n[24167];
assign t[24168] = t[24167] ^ n[24168];
assign t[24169] = t[24168] ^ n[24169];
assign t[24170] = t[24169] ^ n[24170];
assign t[24171] = t[24170] ^ n[24171];
assign t[24172] = t[24171] ^ n[24172];
assign t[24173] = t[24172] ^ n[24173];
assign t[24174] = t[24173] ^ n[24174];
assign t[24175] = t[24174] ^ n[24175];
assign t[24176] = t[24175] ^ n[24176];
assign t[24177] = t[24176] ^ n[24177];
assign t[24178] = t[24177] ^ n[24178];
assign t[24179] = t[24178] ^ n[24179];
assign t[24180] = t[24179] ^ n[24180];
assign t[24181] = t[24180] ^ n[24181];
assign t[24182] = t[24181] ^ n[24182];
assign t[24183] = t[24182] ^ n[24183];
assign t[24184] = t[24183] ^ n[24184];
assign t[24185] = t[24184] ^ n[24185];
assign t[24186] = t[24185] ^ n[24186];
assign t[24187] = t[24186] ^ n[24187];
assign t[24188] = t[24187] ^ n[24188];
assign t[24189] = t[24188] ^ n[24189];
assign t[24190] = t[24189] ^ n[24190];
assign t[24191] = t[24190] ^ n[24191];
assign t[24192] = t[24191] ^ n[24192];
assign t[24193] = t[24192] ^ n[24193];
assign t[24194] = t[24193] ^ n[24194];
assign t[24195] = t[24194] ^ n[24195];
assign t[24196] = t[24195] ^ n[24196];
assign t[24197] = t[24196] ^ n[24197];
assign t[24198] = t[24197] ^ n[24198];
assign t[24199] = t[24198] ^ n[24199];
assign t[24200] = t[24199] ^ n[24200];
assign t[24201] = t[24200] ^ n[24201];
assign t[24202] = t[24201] ^ n[24202];
assign t[24203] = t[24202] ^ n[24203];
assign t[24204] = t[24203] ^ n[24204];
assign t[24205] = t[24204] ^ n[24205];
assign t[24206] = t[24205] ^ n[24206];
assign t[24207] = t[24206] ^ n[24207];
assign t[24208] = t[24207] ^ n[24208];
assign t[24209] = t[24208] ^ n[24209];
assign t[24210] = t[24209] ^ n[24210];
assign t[24211] = t[24210] ^ n[24211];
assign t[24212] = t[24211] ^ n[24212];
assign t[24213] = t[24212] ^ n[24213];
assign t[24214] = t[24213] ^ n[24214];
assign t[24215] = t[24214] ^ n[24215];
assign t[24216] = t[24215] ^ n[24216];
assign t[24217] = t[24216] ^ n[24217];
assign t[24218] = t[24217] ^ n[24218];
assign t[24219] = t[24218] ^ n[24219];
assign t[24220] = t[24219] ^ n[24220];
assign t[24221] = t[24220] ^ n[24221];
assign t[24222] = t[24221] ^ n[24222];
assign t[24223] = t[24222] ^ n[24223];
assign t[24224] = t[24223] ^ n[24224];
assign t[24225] = t[24224] ^ n[24225];
assign t[24226] = t[24225] ^ n[24226];
assign t[24227] = t[24226] ^ n[24227];
assign t[24228] = t[24227] ^ n[24228];
assign t[24229] = t[24228] ^ n[24229];
assign t[24230] = t[24229] ^ n[24230];
assign t[24231] = t[24230] ^ n[24231];
assign t[24232] = t[24231] ^ n[24232];
assign t[24233] = t[24232] ^ n[24233];
assign t[24234] = t[24233] ^ n[24234];
assign t[24235] = t[24234] ^ n[24235];
assign t[24236] = t[24235] ^ n[24236];
assign t[24237] = t[24236] ^ n[24237];
assign t[24238] = t[24237] ^ n[24238];
assign t[24239] = t[24238] ^ n[24239];
assign t[24240] = t[24239] ^ n[24240];
assign t[24241] = t[24240] ^ n[24241];
assign t[24242] = t[24241] ^ n[24242];
assign t[24243] = t[24242] ^ n[24243];
assign t[24244] = t[24243] ^ n[24244];
assign t[24245] = t[24244] ^ n[24245];
assign t[24246] = t[24245] ^ n[24246];
assign t[24247] = t[24246] ^ n[24247];
assign t[24248] = t[24247] ^ n[24248];
assign t[24249] = t[24248] ^ n[24249];
assign t[24250] = t[24249] ^ n[24250];
assign t[24251] = t[24250] ^ n[24251];
assign t[24252] = t[24251] ^ n[24252];
assign t[24253] = t[24252] ^ n[24253];
assign t[24254] = t[24253] ^ n[24254];
assign t[24255] = t[24254] ^ n[24255];
assign t[24256] = t[24255] ^ n[24256];
assign t[24257] = t[24256] ^ n[24257];
assign t[24258] = t[24257] ^ n[24258];
assign t[24259] = t[24258] ^ n[24259];
assign t[24260] = t[24259] ^ n[24260];
assign t[24261] = t[24260] ^ n[24261];
assign t[24262] = t[24261] ^ n[24262];
assign t[24263] = t[24262] ^ n[24263];
assign t[24264] = t[24263] ^ n[24264];
assign t[24265] = t[24264] ^ n[24265];
assign t[24266] = t[24265] ^ n[24266];
assign t[24267] = t[24266] ^ n[24267];
assign t[24268] = t[24267] ^ n[24268];
assign t[24269] = t[24268] ^ n[24269];
assign t[24270] = t[24269] ^ n[24270];
assign t[24271] = t[24270] ^ n[24271];
assign t[24272] = t[24271] ^ n[24272];
assign t[24273] = t[24272] ^ n[24273];
assign t[24274] = t[24273] ^ n[24274];
assign t[24275] = t[24274] ^ n[24275];
assign t[24276] = t[24275] ^ n[24276];
assign t[24277] = t[24276] ^ n[24277];
assign t[24278] = t[24277] ^ n[24278];
assign t[24279] = t[24278] ^ n[24279];
assign t[24280] = t[24279] ^ n[24280];
assign t[24281] = t[24280] ^ n[24281];
assign t[24282] = t[24281] ^ n[24282];
assign t[24283] = t[24282] ^ n[24283];
assign t[24284] = t[24283] ^ n[24284];
assign t[24285] = t[24284] ^ n[24285];
assign t[24286] = t[24285] ^ n[24286];
assign t[24287] = t[24286] ^ n[24287];
assign t[24288] = t[24287] ^ n[24288];
assign t[24289] = t[24288] ^ n[24289];
assign t[24290] = t[24289] ^ n[24290];
assign t[24291] = t[24290] ^ n[24291];
assign t[24292] = t[24291] ^ n[24292];
assign t[24293] = t[24292] ^ n[24293];
assign t[24294] = t[24293] ^ n[24294];
assign t[24295] = t[24294] ^ n[24295];
assign t[24296] = t[24295] ^ n[24296];
assign t[24297] = t[24296] ^ n[24297];
assign t[24298] = t[24297] ^ n[24298];
assign t[24299] = t[24298] ^ n[24299];
assign t[24300] = t[24299] ^ n[24300];
assign t[24301] = t[24300] ^ n[24301];
assign t[24302] = t[24301] ^ n[24302];
assign t[24303] = t[24302] ^ n[24303];
assign t[24304] = t[24303] ^ n[24304];
assign t[24305] = t[24304] ^ n[24305];
assign t[24306] = t[24305] ^ n[24306];
assign t[24307] = t[24306] ^ n[24307];
assign t[24308] = t[24307] ^ n[24308];
assign t[24309] = t[24308] ^ n[24309];
assign t[24310] = t[24309] ^ n[24310];
assign t[24311] = t[24310] ^ n[24311];
assign t[24312] = t[24311] ^ n[24312];
assign t[24313] = t[24312] ^ n[24313];
assign t[24314] = t[24313] ^ n[24314];
assign t[24315] = t[24314] ^ n[24315];
assign t[24316] = t[24315] ^ n[24316];
assign t[24317] = t[24316] ^ n[24317];
assign t[24318] = t[24317] ^ n[24318];
assign t[24319] = t[24318] ^ n[24319];
assign t[24320] = t[24319] ^ n[24320];
assign t[24321] = t[24320] ^ n[24321];
assign t[24322] = t[24321] ^ n[24322];
assign t[24323] = t[24322] ^ n[24323];
assign t[24324] = t[24323] ^ n[24324];
assign t[24325] = t[24324] ^ n[24325];
assign t[24326] = t[24325] ^ n[24326];
assign t[24327] = t[24326] ^ n[24327];
assign t[24328] = t[24327] ^ n[24328];
assign t[24329] = t[24328] ^ n[24329];
assign t[24330] = t[24329] ^ n[24330];
assign t[24331] = t[24330] ^ n[24331];
assign t[24332] = t[24331] ^ n[24332];
assign t[24333] = t[24332] ^ n[24333];
assign t[24334] = t[24333] ^ n[24334];
assign t[24335] = t[24334] ^ n[24335];
assign t[24336] = t[24335] ^ n[24336];
assign t[24337] = t[24336] ^ n[24337];
assign t[24338] = t[24337] ^ n[24338];
assign t[24339] = t[24338] ^ n[24339];
assign t[24340] = t[24339] ^ n[24340];
assign t[24341] = t[24340] ^ n[24341];
assign t[24342] = t[24341] ^ n[24342];
assign t[24343] = t[24342] ^ n[24343];
assign t[24344] = t[24343] ^ n[24344];
assign t[24345] = t[24344] ^ n[24345];
assign t[24346] = t[24345] ^ n[24346];
assign t[24347] = t[24346] ^ n[24347];
assign t[24348] = t[24347] ^ n[24348];
assign t[24349] = t[24348] ^ n[24349];
assign t[24350] = t[24349] ^ n[24350];
assign t[24351] = t[24350] ^ n[24351];
assign t[24352] = t[24351] ^ n[24352];
assign t[24353] = t[24352] ^ n[24353];
assign t[24354] = t[24353] ^ n[24354];
assign t[24355] = t[24354] ^ n[24355];
assign t[24356] = t[24355] ^ n[24356];
assign t[24357] = t[24356] ^ n[24357];
assign t[24358] = t[24357] ^ n[24358];
assign t[24359] = t[24358] ^ n[24359];
assign t[24360] = t[24359] ^ n[24360];
assign t[24361] = t[24360] ^ n[24361];
assign t[24362] = t[24361] ^ n[24362];
assign t[24363] = t[24362] ^ n[24363];
assign t[24364] = t[24363] ^ n[24364];
assign t[24365] = t[24364] ^ n[24365];
assign t[24366] = t[24365] ^ n[24366];
assign t[24367] = t[24366] ^ n[24367];
assign t[24368] = t[24367] ^ n[24368];
assign t[24369] = t[24368] ^ n[24369];
assign t[24370] = t[24369] ^ n[24370];
assign t[24371] = t[24370] ^ n[24371];
assign t[24372] = t[24371] ^ n[24372];
assign t[24373] = t[24372] ^ n[24373];
assign t[24374] = t[24373] ^ n[24374];
assign t[24375] = t[24374] ^ n[24375];
assign t[24376] = t[24375] ^ n[24376];
assign t[24377] = t[24376] ^ n[24377];
assign t[24378] = t[24377] ^ n[24378];
assign t[24379] = t[24378] ^ n[24379];
assign t[24380] = t[24379] ^ n[24380];
assign t[24381] = t[24380] ^ n[24381];
assign t[24382] = t[24381] ^ n[24382];
assign t[24383] = t[24382] ^ n[24383];
assign t[24384] = t[24383] ^ n[24384];
assign t[24385] = t[24384] ^ n[24385];
assign t[24386] = t[24385] ^ n[24386];
assign t[24387] = t[24386] ^ n[24387];
assign t[24388] = t[24387] ^ n[24388];
assign t[24389] = t[24388] ^ n[24389];
assign t[24390] = t[24389] ^ n[24390];
assign t[24391] = t[24390] ^ n[24391];
assign t[24392] = t[24391] ^ n[24392];
assign t[24393] = t[24392] ^ n[24393];
assign t[24394] = t[24393] ^ n[24394];
assign t[24395] = t[24394] ^ n[24395];
assign t[24396] = t[24395] ^ n[24396];
assign t[24397] = t[24396] ^ n[24397];
assign t[24398] = t[24397] ^ n[24398];
assign t[24399] = t[24398] ^ n[24399];
assign t[24400] = t[24399] ^ n[24400];
assign t[24401] = t[24400] ^ n[24401];
assign t[24402] = t[24401] ^ n[24402];
assign t[24403] = t[24402] ^ n[24403];
assign t[24404] = t[24403] ^ n[24404];
assign t[24405] = t[24404] ^ n[24405];
assign t[24406] = t[24405] ^ n[24406];
assign t[24407] = t[24406] ^ n[24407];
assign t[24408] = t[24407] ^ n[24408];
assign t[24409] = t[24408] ^ n[24409];
assign t[24410] = t[24409] ^ n[24410];
assign t[24411] = t[24410] ^ n[24411];
assign t[24412] = t[24411] ^ n[24412];
assign t[24413] = t[24412] ^ n[24413];
assign t[24414] = t[24413] ^ n[24414];
assign t[24415] = t[24414] ^ n[24415];
assign t[24416] = t[24415] ^ n[24416];
assign t[24417] = t[24416] ^ n[24417];
assign t[24418] = t[24417] ^ n[24418];
assign t[24419] = t[24418] ^ n[24419];
assign t[24420] = t[24419] ^ n[24420];
assign t[24421] = t[24420] ^ n[24421];
assign t[24422] = t[24421] ^ n[24422];
assign t[24423] = t[24422] ^ n[24423];
assign t[24424] = t[24423] ^ n[24424];
assign t[24425] = t[24424] ^ n[24425];
assign t[24426] = t[24425] ^ n[24426];
assign t[24427] = t[24426] ^ n[24427];
assign t[24428] = t[24427] ^ n[24428];
assign t[24429] = t[24428] ^ n[24429];
assign t[24430] = t[24429] ^ n[24430];
assign t[24431] = t[24430] ^ n[24431];
assign t[24432] = t[24431] ^ n[24432];
assign t[24433] = t[24432] ^ n[24433];
assign t[24434] = t[24433] ^ n[24434];
assign t[24435] = t[24434] ^ n[24435];
assign t[24436] = t[24435] ^ n[24436];
assign t[24437] = t[24436] ^ n[24437];
assign t[24438] = t[24437] ^ n[24438];
assign t[24439] = t[24438] ^ n[24439];
assign t[24440] = t[24439] ^ n[24440];
assign t[24441] = t[24440] ^ n[24441];
assign t[24442] = t[24441] ^ n[24442];
assign t[24443] = t[24442] ^ n[24443];
assign t[24444] = t[24443] ^ n[24444];
assign t[24445] = t[24444] ^ n[24445];
assign t[24446] = t[24445] ^ n[24446];
assign t[24447] = t[24446] ^ n[24447];
assign t[24448] = t[24447] ^ n[24448];
assign t[24449] = t[24448] ^ n[24449];
assign t[24450] = t[24449] ^ n[24450];
assign t[24451] = t[24450] ^ n[24451];
assign t[24452] = t[24451] ^ n[24452];
assign t[24453] = t[24452] ^ n[24453];
assign t[24454] = t[24453] ^ n[24454];
assign t[24455] = t[24454] ^ n[24455];
assign t[24456] = t[24455] ^ n[24456];
assign t[24457] = t[24456] ^ n[24457];
assign t[24458] = t[24457] ^ n[24458];
assign t[24459] = t[24458] ^ n[24459];
assign t[24460] = t[24459] ^ n[24460];
assign t[24461] = t[24460] ^ n[24461];
assign t[24462] = t[24461] ^ n[24462];
assign t[24463] = t[24462] ^ n[24463];
assign t[24464] = t[24463] ^ n[24464];
assign t[24465] = t[24464] ^ n[24465];
assign t[24466] = t[24465] ^ n[24466];
assign t[24467] = t[24466] ^ n[24467];
assign t[24468] = t[24467] ^ n[24468];
assign t[24469] = t[24468] ^ n[24469];
assign t[24470] = t[24469] ^ n[24470];
assign t[24471] = t[24470] ^ n[24471];
assign t[24472] = t[24471] ^ n[24472];
assign t[24473] = t[24472] ^ n[24473];
assign t[24474] = t[24473] ^ n[24474];
assign t[24475] = t[24474] ^ n[24475];
assign t[24476] = t[24475] ^ n[24476];
assign t[24477] = t[24476] ^ n[24477];
assign t[24478] = t[24477] ^ n[24478];
assign t[24479] = t[24478] ^ n[24479];
assign t[24480] = t[24479] ^ n[24480];
assign t[24481] = t[24480] ^ n[24481];
assign t[24482] = t[24481] ^ n[24482];
assign t[24483] = t[24482] ^ n[24483];
assign t[24484] = t[24483] ^ n[24484];
assign t[24485] = t[24484] ^ n[24485];
assign t[24486] = t[24485] ^ n[24486];
assign t[24487] = t[24486] ^ n[24487];
assign t[24488] = t[24487] ^ n[24488];
assign t[24489] = t[24488] ^ n[24489];
assign t[24490] = t[24489] ^ n[24490];
assign t[24491] = t[24490] ^ n[24491];
assign t[24492] = t[24491] ^ n[24492];
assign t[24493] = t[24492] ^ n[24493];
assign t[24494] = t[24493] ^ n[24494];
assign t[24495] = t[24494] ^ n[24495];
assign t[24496] = t[24495] ^ n[24496];
assign t[24497] = t[24496] ^ n[24497];
assign t[24498] = t[24497] ^ n[24498];
assign t[24499] = t[24498] ^ n[24499];
assign t[24500] = t[24499] ^ n[24500];
assign t[24501] = t[24500] ^ n[24501];
assign t[24502] = t[24501] ^ n[24502];
assign t[24503] = t[24502] ^ n[24503];
assign t[24504] = t[24503] ^ n[24504];
assign t[24505] = t[24504] ^ n[24505];
assign t[24506] = t[24505] ^ n[24506];
assign t[24507] = t[24506] ^ n[24507];
assign t[24508] = t[24507] ^ n[24508];
assign t[24509] = t[24508] ^ n[24509];
assign t[24510] = t[24509] ^ n[24510];
assign t[24511] = t[24510] ^ n[24511];
assign t[24512] = t[24511] ^ n[24512];
assign t[24513] = t[24512] ^ n[24513];
assign t[24514] = t[24513] ^ n[24514];
assign t[24515] = t[24514] ^ n[24515];
assign t[24516] = t[24515] ^ n[24516];
assign t[24517] = t[24516] ^ n[24517];
assign t[24518] = t[24517] ^ n[24518];
assign t[24519] = t[24518] ^ n[24519];
assign t[24520] = t[24519] ^ n[24520];
assign t[24521] = t[24520] ^ n[24521];
assign t[24522] = t[24521] ^ n[24522];
assign t[24523] = t[24522] ^ n[24523];
assign t[24524] = t[24523] ^ n[24524];
assign t[24525] = t[24524] ^ n[24525];
assign t[24526] = t[24525] ^ n[24526];
assign t[24527] = t[24526] ^ n[24527];
assign t[24528] = t[24527] ^ n[24528];
assign t[24529] = t[24528] ^ n[24529];
assign t[24530] = t[24529] ^ n[24530];
assign t[24531] = t[24530] ^ n[24531];
assign t[24532] = t[24531] ^ n[24532];
assign t[24533] = t[24532] ^ n[24533];
assign t[24534] = t[24533] ^ n[24534];
assign t[24535] = t[24534] ^ n[24535];
assign t[24536] = t[24535] ^ n[24536];
assign t[24537] = t[24536] ^ n[24537];
assign t[24538] = t[24537] ^ n[24538];
assign t[24539] = t[24538] ^ n[24539];
assign t[24540] = t[24539] ^ n[24540];
assign t[24541] = t[24540] ^ n[24541];
assign t[24542] = t[24541] ^ n[24542];
assign t[24543] = t[24542] ^ n[24543];
assign t[24544] = t[24543] ^ n[24544];
assign t[24545] = t[24544] ^ n[24545];
assign t[24546] = t[24545] ^ n[24546];
assign t[24547] = t[24546] ^ n[24547];
assign t[24548] = t[24547] ^ n[24548];
assign t[24549] = t[24548] ^ n[24549];
assign t[24550] = t[24549] ^ n[24550];
assign t[24551] = t[24550] ^ n[24551];
assign t[24552] = t[24551] ^ n[24552];
assign t[24553] = t[24552] ^ n[24553];
assign t[24554] = t[24553] ^ n[24554];
assign t[24555] = t[24554] ^ n[24555];
assign t[24556] = t[24555] ^ n[24556];
assign t[24557] = t[24556] ^ n[24557];
assign t[24558] = t[24557] ^ n[24558];
assign t[24559] = t[24558] ^ n[24559];
assign t[24560] = t[24559] ^ n[24560];
assign t[24561] = t[24560] ^ n[24561];
assign t[24562] = t[24561] ^ n[24562];
assign t[24563] = t[24562] ^ n[24563];
assign t[24564] = t[24563] ^ n[24564];
assign t[24565] = t[24564] ^ n[24565];
assign t[24566] = t[24565] ^ n[24566];
assign t[24567] = t[24566] ^ n[24567];
assign t[24568] = t[24567] ^ n[24568];
assign t[24569] = t[24568] ^ n[24569];
assign t[24570] = t[24569] ^ n[24570];
assign t[24571] = t[24570] ^ n[24571];
assign t[24572] = t[24571] ^ n[24572];
assign t[24573] = t[24572] ^ n[24573];
assign t[24574] = t[24573] ^ n[24574];
assign t[24575] = t[24574] ^ n[24575];
assign t[24576] = t[24575] ^ n[24576];
assign t[24577] = t[24576] ^ n[24577];
assign t[24578] = t[24577] ^ n[24578];
assign t[24579] = t[24578] ^ n[24579];
assign t[24580] = t[24579] ^ n[24580];
assign t[24581] = t[24580] ^ n[24581];
assign t[24582] = t[24581] ^ n[24582];
assign t[24583] = t[24582] ^ n[24583];
assign t[24584] = t[24583] ^ n[24584];
assign t[24585] = t[24584] ^ n[24585];
assign t[24586] = t[24585] ^ n[24586];
assign t[24587] = t[24586] ^ n[24587];
assign t[24588] = t[24587] ^ n[24588];
assign t[24589] = t[24588] ^ n[24589];
assign t[24590] = t[24589] ^ n[24590];
assign t[24591] = t[24590] ^ n[24591];
assign t[24592] = t[24591] ^ n[24592];
assign t[24593] = t[24592] ^ n[24593];
assign t[24594] = t[24593] ^ n[24594];
assign t[24595] = t[24594] ^ n[24595];
assign t[24596] = t[24595] ^ n[24596];
assign t[24597] = t[24596] ^ n[24597];
assign t[24598] = t[24597] ^ n[24598];
assign t[24599] = t[24598] ^ n[24599];
assign t[24600] = t[24599] ^ n[24600];
assign t[24601] = t[24600] ^ n[24601];
assign t[24602] = t[24601] ^ n[24602];
assign t[24603] = t[24602] ^ n[24603];
assign t[24604] = t[24603] ^ n[24604];
assign t[24605] = t[24604] ^ n[24605];
assign t[24606] = t[24605] ^ n[24606];
assign t[24607] = t[24606] ^ n[24607];
assign t[24608] = t[24607] ^ n[24608];
assign t[24609] = t[24608] ^ n[24609];
assign t[24610] = t[24609] ^ n[24610];
assign t[24611] = t[24610] ^ n[24611];
assign t[24612] = t[24611] ^ n[24612];
assign t[24613] = t[24612] ^ n[24613];
assign t[24614] = t[24613] ^ n[24614];
assign t[24615] = t[24614] ^ n[24615];
assign t[24616] = t[24615] ^ n[24616];
assign t[24617] = t[24616] ^ n[24617];
assign t[24618] = t[24617] ^ n[24618];
assign t[24619] = t[24618] ^ n[24619];
assign t[24620] = t[24619] ^ n[24620];
assign t[24621] = t[24620] ^ n[24621];
assign t[24622] = t[24621] ^ n[24622];
assign t[24623] = t[24622] ^ n[24623];
assign t[24624] = t[24623] ^ n[24624];
assign t[24625] = t[24624] ^ n[24625];
assign t[24626] = t[24625] ^ n[24626];
assign t[24627] = t[24626] ^ n[24627];
assign t[24628] = t[24627] ^ n[24628];
assign t[24629] = t[24628] ^ n[24629];
assign t[24630] = t[24629] ^ n[24630];
assign t[24631] = t[24630] ^ n[24631];
assign t[24632] = t[24631] ^ n[24632];
assign t[24633] = t[24632] ^ n[24633];
assign t[24634] = t[24633] ^ n[24634];
assign t[24635] = t[24634] ^ n[24635];
assign t[24636] = t[24635] ^ n[24636];
assign t[24637] = t[24636] ^ n[24637];
assign t[24638] = t[24637] ^ n[24638];
assign t[24639] = t[24638] ^ n[24639];
assign t[24640] = t[24639] ^ n[24640];
assign t[24641] = t[24640] ^ n[24641];
assign t[24642] = t[24641] ^ n[24642];
assign t[24643] = t[24642] ^ n[24643];
assign t[24644] = t[24643] ^ n[24644];
assign t[24645] = t[24644] ^ n[24645];
assign t[24646] = t[24645] ^ n[24646];
assign t[24647] = t[24646] ^ n[24647];
assign t[24648] = t[24647] ^ n[24648];
assign t[24649] = t[24648] ^ n[24649];
assign t[24650] = t[24649] ^ n[24650];
assign t[24651] = t[24650] ^ n[24651];
assign t[24652] = t[24651] ^ n[24652];
assign t[24653] = t[24652] ^ n[24653];
assign t[24654] = t[24653] ^ n[24654];
assign t[24655] = t[24654] ^ n[24655];
assign t[24656] = t[24655] ^ n[24656];
assign t[24657] = t[24656] ^ n[24657];
assign t[24658] = t[24657] ^ n[24658];
assign t[24659] = t[24658] ^ n[24659];
assign t[24660] = t[24659] ^ n[24660];
assign t[24661] = t[24660] ^ n[24661];
assign t[24662] = t[24661] ^ n[24662];
assign t[24663] = t[24662] ^ n[24663];
assign t[24664] = t[24663] ^ n[24664];
assign t[24665] = t[24664] ^ n[24665];
assign t[24666] = t[24665] ^ n[24666];
assign t[24667] = t[24666] ^ n[24667];
assign t[24668] = t[24667] ^ n[24668];
assign t[24669] = t[24668] ^ n[24669];
assign t[24670] = t[24669] ^ n[24670];
assign t[24671] = t[24670] ^ n[24671];
assign t[24672] = t[24671] ^ n[24672];
assign t[24673] = t[24672] ^ n[24673];
assign t[24674] = t[24673] ^ n[24674];
assign t[24675] = t[24674] ^ n[24675];
assign t[24676] = t[24675] ^ n[24676];
assign t[24677] = t[24676] ^ n[24677];
assign t[24678] = t[24677] ^ n[24678];
assign t[24679] = t[24678] ^ n[24679];
assign t[24680] = t[24679] ^ n[24680];
assign t[24681] = t[24680] ^ n[24681];
assign t[24682] = t[24681] ^ n[24682];
assign t[24683] = t[24682] ^ n[24683];
assign t[24684] = t[24683] ^ n[24684];
assign t[24685] = t[24684] ^ n[24685];
assign t[24686] = t[24685] ^ n[24686];
assign t[24687] = t[24686] ^ n[24687];
assign t[24688] = t[24687] ^ n[24688];
assign t[24689] = t[24688] ^ n[24689];
assign t[24690] = t[24689] ^ n[24690];
assign t[24691] = t[24690] ^ n[24691];
assign t[24692] = t[24691] ^ n[24692];
assign t[24693] = t[24692] ^ n[24693];
assign t[24694] = t[24693] ^ n[24694];
assign t[24695] = t[24694] ^ n[24695];
assign t[24696] = t[24695] ^ n[24696];
assign t[24697] = t[24696] ^ n[24697];
assign t[24698] = t[24697] ^ n[24698];
assign t[24699] = t[24698] ^ n[24699];
assign t[24700] = t[24699] ^ n[24700];
assign t[24701] = t[24700] ^ n[24701];
assign t[24702] = t[24701] ^ n[24702];
assign t[24703] = t[24702] ^ n[24703];
assign t[24704] = t[24703] ^ n[24704];
assign t[24705] = t[24704] ^ n[24705];
assign t[24706] = t[24705] ^ n[24706];
assign t[24707] = t[24706] ^ n[24707];
assign t[24708] = t[24707] ^ n[24708];
assign t[24709] = t[24708] ^ n[24709];
assign t[24710] = t[24709] ^ n[24710];
assign t[24711] = t[24710] ^ n[24711];
assign t[24712] = t[24711] ^ n[24712];
assign t[24713] = t[24712] ^ n[24713];
assign t[24714] = t[24713] ^ n[24714];
assign t[24715] = t[24714] ^ n[24715];
assign t[24716] = t[24715] ^ n[24716];
assign t[24717] = t[24716] ^ n[24717];
assign t[24718] = t[24717] ^ n[24718];
assign t[24719] = t[24718] ^ n[24719];
assign t[24720] = t[24719] ^ n[24720];
assign t[24721] = t[24720] ^ n[24721];
assign t[24722] = t[24721] ^ n[24722];
assign t[24723] = t[24722] ^ n[24723];
assign t[24724] = t[24723] ^ n[24724];
assign t[24725] = t[24724] ^ n[24725];
assign t[24726] = t[24725] ^ n[24726];
assign t[24727] = t[24726] ^ n[24727];
assign t[24728] = t[24727] ^ n[24728];
assign t[24729] = t[24728] ^ n[24729];
assign t[24730] = t[24729] ^ n[24730];
assign t[24731] = t[24730] ^ n[24731];
assign t[24732] = t[24731] ^ n[24732];
assign t[24733] = t[24732] ^ n[24733];
assign t[24734] = t[24733] ^ n[24734];
assign t[24735] = t[24734] ^ n[24735];
assign t[24736] = t[24735] ^ n[24736];
assign t[24737] = t[24736] ^ n[24737];
assign t[24738] = t[24737] ^ n[24738];
assign t[24739] = t[24738] ^ n[24739];
assign t[24740] = t[24739] ^ n[24740];
assign t[24741] = t[24740] ^ n[24741];
assign t[24742] = t[24741] ^ n[24742];
assign t[24743] = t[24742] ^ n[24743];
assign t[24744] = t[24743] ^ n[24744];
assign t[24745] = t[24744] ^ n[24745];
assign t[24746] = t[24745] ^ n[24746];
assign t[24747] = t[24746] ^ n[24747];
assign t[24748] = t[24747] ^ n[24748];
assign t[24749] = t[24748] ^ n[24749];
assign t[24750] = t[24749] ^ n[24750];
assign t[24751] = t[24750] ^ n[24751];
assign t[24752] = t[24751] ^ n[24752];
assign t[24753] = t[24752] ^ n[24753];
assign t[24754] = t[24753] ^ n[24754];
assign t[24755] = t[24754] ^ n[24755];
assign t[24756] = t[24755] ^ n[24756];
assign t[24757] = t[24756] ^ n[24757];
assign t[24758] = t[24757] ^ n[24758];
assign t[24759] = t[24758] ^ n[24759];
assign t[24760] = t[24759] ^ n[24760];
assign t[24761] = t[24760] ^ n[24761];
assign t[24762] = t[24761] ^ n[24762];
assign t[24763] = t[24762] ^ n[24763];
assign t[24764] = t[24763] ^ n[24764];
assign t[24765] = t[24764] ^ n[24765];
assign t[24766] = t[24765] ^ n[24766];
assign t[24767] = t[24766] ^ n[24767];
assign t[24768] = t[24767] ^ n[24768];
assign t[24769] = t[24768] ^ n[24769];
assign t[24770] = t[24769] ^ n[24770];
assign t[24771] = t[24770] ^ n[24771];
assign t[24772] = t[24771] ^ n[24772];
assign t[24773] = t[24772] ^ n[24773];
assign t[24774] = t[24773] ^ n[24774];
assign t[24775] = t[24774] ^ n[24775];
assign t[24776] = t[24775] ^ n[24776];
assign t[24777] = t[24776] ^ n[24777];
assign t[24778] = t[24777] ^ n[24778];
assign t[24779] = t[24778] ^ n[24779];
assign t[24780] = t[24779] ^ n[24780];
assign t[24781] = t[24780] ^ n[24781];
assign t[24782] = t[24781] ^ n[24782];
assign t[24783] = t[24782] ^ n[24783];
assign t[24784] = t[24783] ^ n[24784];
assign t[24785] = t[24784] ^ n[24785];
assign t[24786] = t[24785] ^ n[24786];
assign t[24787] = t[24786] ^ n[24787];
assign t[24788] = t[24787] ^ n[24788];
assign t[24789] = t[24788] ^ n[24789];
assign t[24790] = t[24789] ^ n[24790];
assign t[24791] = t[24790] ^ n[24791];
assign t[24792] = t[24791] ^ n[24792];
assign t[24793] = t[24792] ^ n[24793];
assign t[24794] = t[24793] ^ n[24794];
assign t[24795] = t[24794] ^ n[24795];
assign t[24796] = t[24795] ^ n[24796];
assign t[24797] = t[24796] ^ n[24797];
assign t[24798] = t[24797] ^ n[24798];
assign t[24799] = t[24798] ^ n[24799];
assign t[24800] = t[24799] ^ n[24800];
assign t[24801] = t[24800] ^ n[24801];
assign t[24802] = t[24801] ^ n[24802];
assign t[24803] = t[24802] ^ n[24803];
assign t[24804] = t[24803] ^ n[24804];
assign t[24805] = t[24804] ^ n[24805];
assign t[24806] = t[24805] ^ n[24806];
assign t[24807] = t[24806] ^ n[24807];
assign t[24808] = t[24807] ^ n[24808];
assign t[24809] = t[24808] ^ n[24809];
assign t[24810] = t[24809] ^ n[24810];
assign t[24811] = t[24810] ^ n[24811];
assign t[24812] = t[24811] ^ n[24812];
assign t[24813] = t[24812] ^ n[24813];
assign t[24814] = t[24813] ^ n[24814];
assign t[24815] = t[24814] ^ n[24815];
assign t[24816] = t[24815] ^ n[24816];
assign t[24817] = t[24816] ^ n[24817];
assign t[24818] = t[24817] ^ n[24818];
assign t[24819] = t[24818] ^ n[24819];
assign t[24820] = t[24819] ^ n[24820];
assign t[24821] = t[24820] ^ n[24821];
assign t[24822] = t[24821] ^ n[24822];
assign t[24823] = t[24822] ^ n[24823];
assign t[24824] = t[24823] ^ n[24824];
assign t[24825] = t[24824] ^ n[24825];
assign t[24826] = t[24825] ^ n[24826];
assign t[24827] = t[24826] ^ n[24827];
assign t[24828] = t[24827] ^ n[24828];
assign t[24829] = t[24828] ^ n[24829];
assign t[24830] = t[24829] ^ n[24830];
assign t[24831] = t[24830] ^ n[24831];
assign t[24832] = t[24831] ^ n[24832];
assign t[24833] = t[24832] ^ n[24833];
assign t[24834] = t[24833] ^ n[24834];
assign t[24835] = t[24834] ^ n[24835];
assign t[24836] = t[24835] ^ n[24836];
assign t[24837] = t[24836] ^ n[24837];
assign t[24838] = t[24837] ^ n[24838];
assign t[24839] = t[24838] ^ n[24839];
assign t[24840] = t[24839] ^ n[24840];
assign t[24841] = t[24840] ^ n[24841];
assign t[24842] = t[24841] ^ n[24842];
assign t[24843] = t[24842] ^ n[24843];
assign t[24844] = t[24843] ^ n[24844];
assign t[24845] = t[24844] ^ n[24845];
assign t[24846] = t[24845] ^ n[24846];
assign t[24847] = t[24846] ^ n[24847];
assign t[24848] = t[24847] ^ n[24848];
assign t[24849] = t[24848] ^ n[24849];
assign t[24850] = t[24849] ^ n[24850];
assign t[24851] = t[24850] ^ n[24851];
assign t[24852] = t[24851] ^ n[24852];
assign t[24853] = t[24852] ^ n[24853];
assign t[24854] = t[24853] ^ n[24854];
assign t[24855] = t[24854] ^ n[24855];
assign t[24856] = t[24855] ^ n[24856];
assign t[24857] = t[24856] ^ n[24857];
assign t[24858] = t[24857] ^ n[24858];
assign t[24859] = t[24858] ^ n[24859];
assign t[24860] = t[24859] ^ n[24860];
assign t[24861] = t[24860] ^ n[24861];
assign t[24862] = t[24861] ^ n[24862];
assign t[24863] = t[24862] ^ n[24863];
assign t[24864] = t[24863] ^ n[24864];
assign t[24865] = t[24864] ^ n[24865];
assign t[24866] = t[24865] ^ n[24866];
assign t[24867] = t[24866] ^ n[24867];
assign t[24868] = t[24867] ^ n[24868];
assign t[24869] = t[24868] ^ n[24869];
assign t[24870] = t[24869] ^ n[24870];
assign t[24871] = t[24870] ^ n[24871];
assign t[24872] = t[24871] ^ n[24872];
assign t[24873] = t[24872] ^ n[24873];
assign t[24874] = t[24873] ^ n[24874];
assign t[24875] = t[24874] ^ n[24875];
assign t[24876] = t[24875] ^ n[24876];
assign t[24877] = t[24876] ^ n[24877];
assign t[24878] = t[24877] ^ n[24878];
assign t[24879] = t[24878] ^ n[24879];
assign t[24880] = t[24879] ^ n[24880];
assign t[24881] = t[24880] ^ n[24881];
assign t[24882] = t[24881] ^ n[24882];
assign t[24883] = t[24882] ^ n[24883];
assign t[24884] = t[24883] ^ n[24884];
assign t[24885] = t[24884] ^ n[24885];
assign t[24886] = t[24885] ^ n[24886];
assign t[24887] = t[24886] ^ n[24887];
assign t[24888] = t[24887] ^ n[24888];
assign t[24889] = t[24888] ^ n[24889];
assign t[24890] = t[24889] ^ n[24890];
assign t[24891] = t[24890] ^ n[24891];
assign t[24892] = t[24891] ^ n[24892];
assign t[24893] = t[24892] ^ n[24893];
assign t[24894] = t[24893] ^ n[24894];
assign t[24895] = t[24894] ^ n[24895];
assign t[24896] = t[24895] ^ n[24896];
assign t[24897] = t[24896] ^ n[24897];
assign t[24898] = t[24897] ^ n[24898];
assign t[24899] = t[24898] ^ n[24899];
assign t[24900] = t[24899] ^ n[24900];
assign t[24901] = t[24900] ^ n[24901];
assign t[24902] = t[24901] ^ n[24902];
assign t[24903] = t[24902] ^ n[24903];
assign t[24904] = t[24903] ^ n[24904];
assign t[24905] = t[24904] ^ n[24905];
assign t[24906] = t[24905] ^ n[24906];
assign t[24907] = t[24906] ^ n[24907];
assign t[24908] = t[24907] ^ n[24908];
assign t[24909] = t[24908] ^ n[24909];
assign t[24910] = t[24909] ^ n[24910];
assign t[24911] = t[24910] ^ n[24911];
assign t[24912] = t[24911] ^ n[24912];
assign t[24913] = t[24912] ^ n[24913];
assign t[24914] = t[24913] ^ n[24914];
assign t[24915] = t[24914] ^ n[24915];
assign t[24916] = t[24915] ^ n[24916];
assign t[24917] = t[24916] ^ n[24917];
assign t[24918] = t[24917] ^ n[24918];
assign t[24919] = t[24918] ^ n[24919];
assign t[24920] = t[24919] ^ n[24920];
assign t[24921] = t[24920] ^ n[24921];
assign t[24922] = t[24921] ^ n[24922];
assign t[24923] = t[24922] ^ n[24923];
assign t[24924] = t[24923] ^ n[24924];
assign t[24925] = t[24924] ^ n[24925];
assign t[24926] = t[24925] ^ n[24926];
assign t[24927] = t[24926] ^ n[24927];
assign t[24928] = t[24927] ^ n[24928];
assign t[24929] = t[24928] ^ n[24929];
assign t[24930] = t[24929] ^ n[24930];
assign t[24931] = t[24930] ^ n[24931];
assign t[24932] = t[24931] ^ n[24932];
assign t[24933] = t[24932] ^ n[24933];
assign t[24934] = t[24933] ^ n[24934];
assign t[24935] = t[24934] ^ n[24935];
assign t[24936] = t[24935] ^ n[24936];
assign t[24937] = t[24936] ^ n[24937];
assign t[24938] = t[24937] ^ n[24938];
assign t[24939] = t[24938] ^ n[24939];
assign t[24940] = t[24939] ^ n[24940];
assign t[24941] = t[24940] ^ n[24941];
assign t[24942] = t[24941] ^ n[24942];
assign t[24943] = t[24942] ^ n[24943];
assign t[24944] = t[24943] ^ n[24944];
assign t[24945] = t[24944] ^ n[24945];
assign t[24946] = t[24945] ^ n[24946];
assign t[24947] = t[24946] ^ n[24947];
assign t[24948] = t[24947] ^ n[24948];
assign t[24949] = t[24948] ^ n[24949];
assign t[24950] = t[24949] ^ n[24950];
assign t[24951] = t[24950] ^ n[24951];
assign t[24952] = t[24951] ^ n[24952];
assign t[24953] = t[24952] ^ n[24953];
assign t[24954] = t[24953] ^ n[24954];
assign t[24955] = t[24954] ^ n[24955];
assign t[24956] = t[24955] ^ n[24956];
assign t[24957] = t[24956] ^ n[24957];
assign t[24958] = t[24957] ^ n[24958];
assign t[24959] = t[24958] ^ n[24959];
assign t[24960] = t[24959] ^ n[24960];
assign t[24961] = t[24960] ^ n[24961];
assign t[24962] = t[24961] ^ n[24962];
assign t[24963] = t[24962] ^ n[24963];
assign t[24964] = t[24963] ^ n[24964];
assign t[24965] = t[24964] ^ n[24965];
assign t[24966] = t[24965] ^ n[24966];
assign t[24967] = t[24966] ^ n[24967];
assign t[24968] = t[24967] ^ n[24968];
assign t[24969] = t[24968] ^ n[24969];
assign t[24970] = t[24969] ^ n[24970];
assign t[24971] = t[24970] ^ n[24971];
assign t[24972] = t[24971] ^ n[24972];
assign t[24973] = t[24972] ^ n[24973];
assign t[24974] = t[24973] ^ n[24974];
assign t[24975] = t[24974] ^ n[24975];
assign t[24976] = t[24975] ^ n[24976];
assign t[24977] = t[24976] ^ n[24977];
assign t[24978] = t[24977] ^ n[24978];
assign t[24979] = t[24978] ^ n[24979];
assign t[24980] = t[24979] ^ n[24980];
assign t[24981] = t[24980] ^ n[24981];
assign t[24982] = t[24981] ^ n[24982];
assign t[24983] = t[24982] ^ n[24983];
assign t[24984] = t[24983] ^ n[24984];
assign t[24985] = t[24984] ^ n[24985];
assign t[24986] = t[24985] ^ n[24986];
assign t[24987] = t[24986] ^ n[24987];
assign t[24988] = t[24987] ^ n[24988];
assign t[24989] = t[24988] ^ n[24989];
assign t[24990] = t[24989] ^ n[24990];
assign t[24991] = t[24990] ^ n[24991];
assign t[24992] = t[24991] ^ n[24992];
assign t[24993] = t[24992] ^ n[24993];
assign t[24994] = t[24993] ^ n[24994];
assign t[24995] = t[24994] ^ n[24995];
assign t[24996] = t[24995] ^ n[24996];
assign t[24997] = t[24996] ^ n[24997];
assign t[24998] = t[24997] ^ n[24998];
assign t[24999] = t[24998] ^ n[24999];
assign t[25000] = t[24999] ^ n[25000];
assign t[25001] = t[25000] ^ n[25001];
assign t[25002] = t[25001] ^ n[25002];
assign t[25003] = t[25002] ^ n[25003];
assign t[25004] = t[25003] ^ n[25004];
assign t[25005] = t[25004] ^ n[25005];
assign t[25006] = t[25005] ^ n[25006];
assign t[25007] = t[25006] ^ n[25007];
assign t[25008] = t[25007] ^ n[25008];
assign t[25009] = t[25008] ^ n[25009];
assign t[25010] = t[25009] ^ n[25010];
assign t[25011] = t[25010] ^ n[25011];
assign t[25012] = t[25011] ^ n[25012];
assign t[25013] = t[25012] ^ n[25013];
assign t[25014] = t[25013] ^ n[25014];
assign t[25015] = t[25014] ^ n[25015];
assign t[25016] = t[25015] ^ n[25016];
assign t[25017] = t[25016] ^ n[25017];
assign t[25018] = t[25017] ^ n[25018];
assign t[25019] = t[25018] ^ n[25019];
assign t[25020] = t[25019] ^ n[25020];
assign t[25021] = t[25020] ^ n[25021];
assign t[25022] = t[25021] ^ n[25022];
assign t[25023] = t[25022] ^ n[25023];
assign t[25024] = t[25023] ^ n[25024];
assign t[25025] = t[25024] ^ n[25025];
assign t[25026] = t[25025] ^ n[25026];
assign t[25027] = t[25026] ^ n[25027];
assign t[25028] = t[25027] ^ n[25028];
assign t[25029] = t[25028] ^ n[25029];
assign t[25030] = t[25029] ^ n[25030];
assign t[25031] = t[25030] ^ n[25031];
assign t[25032] = t[25031] ^ n[25032];
assign t[25033] = t[25032] ^ n[25033];
assign t[25034] = t[25033] ^ n[25034];
assign t[25035] = t[25034] ^ n[25035];
assign t[25036] = t[25035] ^ n[25036];
assign t[25037] = t[25036] ^ n[25037];
assign t[25038] = t[25037] ^ n[25038];
assign t[25039] = t[25038] ^ n[25039];
assign t[25040] = t[25039] ^ n[25040];
assign t[25041] = t[25040] ^ n[25041];
assign t[25042] = t[25041] ^ n[25042];
assign t[25043] = t[25042] ^ n[25043];
assign t[25044] = t[25043] ^ n[25044];
assign t[25045] = t[25044] ^ n[25045];
assign t[25046] = t[25045] ^ n[25046];
assign t[25047] = t[25046] ^ n[25047];
assign t[25048] = t[25047] ^ n[25048];
assign t[25049] = t[25048] ^ n[25049];
assign t[25050] = t[25049] ^ n[25050];
assign t[25051] = t[25050] ^ n[25051];
assign t[25052] = t[25051] ^ n[25052];
assign t[25053] = t[25052] ^ n[25053];
assign t[25054] = t[25053] ^ n[25054];
assign t[25055] = t[25054] ^ n[25055];
assign t[25056] = t[25055] ^ n[25056];
assign t[25057] = t[25056] ^ n[25057];
assign t[25058] = t[25057] ^ n[25058];
assign t[25059] = t[25058] ^ n[25059];
assign t[25060] = t[25059] ^ n[25060];
assign t[25061] = t[25060] ^ n[25061];
assign t[25062] = t[25061] ^ n[25062];
assign t[25063] = t[25062] ^ n[25063];
assign t[25064] = t[25063] ^ n[25064];
assign t[25065] = t[25064] ^ n[25065];
assign t[25066] = t[25065] ^ n[25066];
assign t[25067] = t[25066] ^ n[25067];
assign t[25068] = t[25067] ^ n[25068];
assign t[25069] = t[25068] ^ n[25069];
assign t[25070] = t[25069] ^ n[25070];
assign t[25071] = t[25070] ^ n[25071];
assign t[25072] = t[25071] ^ n[25072];
assign t[25073] = t[25072] ^ n[25073];
assign t[25074] = t[25073] ^ n[25074];
assign t[25075] = t[25074] ^ n[25075];
assign t[25076] = t[25075] ^ n[25076];
assign t[25077] = t[25076] ^ n[25077];
assign t[25078] = t[25077] ^ n[25078];
assign t[25079] = t[25078] ^ n[25079];
assign t[25080] = t[25079] ^ n[25080];
assign t[25081] = t[25080] ^ n[25081];
assign t[25082] = t[25081] ^ n[25082];
assign t[25083] = t[25082] ^ n[25083];
assign t[25084] = t[25083] ^ n[25084];
assign t[25085] = t[25084] ^ n[25085];
assign t[25086] = t[25085] ^ n[25086];
assign t[25087] = t[25086] ^ n[25087];
assign t[25088] = t[25087] ^ n[25088];
assign t[25089] = t[25088] ^ n[25089];
assign t[25090] = t[25089] ^ n[25090];
assign t[25091] = t[25090] ^ n[25091];
assign t[25092] = t[25091] ^ n[25092];
assign t[25093] = t[25092] ^ n[25093];
assign t[25094] = t[25093] ^ n[25094];
assign t[25095] = t[25094] ^ n[25095];
assign t[25096] = t[25095] ^ n[25096];
assign t[25097] = t[25096] ^ n[25097];
assign t[25098] = t[25097] ^ n[25098];
assign t[25099] = t[25098] ^ n[25099];
assign t[25100] = t[25099] ^ n[25100];
assign t[25101] = t[25100] ^ n[25101];
assign t[25102] = t[25101] ^ n[25102];
assign t[25103] = t[25102] ^ n[25103];
assign t[25104] = t[25103] ^ n[25104];
assign t[25105] = t[25104] ^ n[25105];
assign t[25106] = t[25105] ^ n[25106];
assign t[25107] = t[25106] ^ n[25107];
assign t[25108] = t[25107] ^ n[25108];
assign t[25109] = t[25108] ^ n[25109];
assign t[25110] = t[25109] ^ n[25110];
assign t[25111] = t[25110] ^ n[25111];
assign t[25112] = t[25111] ^ n[25112];
assign t[25113] = t[25112] ^ n[25113];
assign t[25114] = t[25113] ^ n[25114];
assign t[25115] = t[25114] ^ n[25115];
assign t[25116] = t[25115] ^ n[25116];
assign t[25117] = t[25116] ^ n[25117];
assign t[25118] = t[25117] ^ n[25118];
assign t[25119] = t[25118] ^ n[25119];
assign t[25120] = t[25119] ^ n[25120];
assign t[25121] = t[25120] ^ n[25121];
assign t[25122] = t[25121] ^ n[25122];
assign t[25123] = t[25122] ^ n[25123];
assign t[25124] = t[25123] ^ n[25124];
assign t[25125] = t[25124] ^ n[25125];
assign t[25126] = t[25125] ^ n[25126];
assign t[25127] = t[25126] ^ n[25127];
assign t[25128] = t[25127] ^ n[25128];
assign t[25129] = t[25128] ^ n[25129];
assign t[25130] = t[25129] ^ n[25130];
assign t[25131] = t[25130] ^ n[25131];
assign t[25132] = t[25131] ^ n[25132];
assign t[25133] = t[25132] ^ n[25133];
assign t[25134] = t[25133] ^ n[25134];
assign t[25135] = t[25134] ^ n[25135];
assign t[25136] = t[25135] ^ n[25136];
assign t[25137] = t[25136] ^ n[25137];
assign t[25138] = t[25137] ^ n[25138];
assign t[25139] = t[25138] ^ n[25139];
assign t[25140] = t[25139] ^ n[25140];
assign t[25141] = t[25140] ^ n[25141];
assign t[25142] = t[25141] ^ n[25142];
assign t[25143] = t[25142] ^ n[25143];
assign t[25144] = t[25143] ^ n[25144];
assign t[25145] = t[25144] ^ n[25145];
assign t[25146] = t[25145] ^ n[25146];
assign t[25147] = t[25146] ^ n[25147];
assign t[25148] = t[25147] ^ n[25148];
assign t[25149] = t[25148] ^ n[25149];
assign t[25150] = t[25149] ^ n[25150];
assign t[25151] = t[25150] ^ n[25151];
assign t[25152] = t[25151] ^ n[25152];
assign t[25153] = t[25152] ^ n[25153];
assign t[25154] = t[25153] ^ n[25154];
assign t[25155] = t[25154] ^ n[25155];
assign t[25156] = t[25155] ^ n[25156];
assign t[25157] = t[25156] ^ n[25157];
assign t[25158] = t[25157] ^ n[25158];
assign t[25159] = t[25158] ^ n[25159];
assign t[25160] = t[25159] ^ n[25160];
assign t[25161] = t[25160] ^ n[25161];
assign t[25162] = t[25161] ^ n[25162];
assign t[25163] = t[25162] ^ n[25163];
assign t[25164] = t[25163] ^ n[25164];
assign t[25165] = t[25164] ^ n[25165];
assign t[25166] = t[25165] ^ n[25166];
assign t[25167] = t[25166] ^ n[25167];
assign t[25168] = t[25167] ^ n[25168];
assign t[25169] = t[25168] ^ n[25169];
assign t[25170] = t[25169] ^ n[25170];
assign t[25171] = t[25170] ^ n[25171];
assign t[25172] = t[25171] ^ n[25172];
assign t[25173] = t[25172] ^ n[25173];
assign t[25174] = t[25173] ^ n[25174];
assign t[25175] = t[25174] ^ n[25175];
assign t[25176] = t[25175] ^ n[25176];
assign t[25177] = t[25176] ^ n[25177];
assign t[25178] = t[25177] ^ n[25178];
assign t[25179] = t[25178] ^ n[25179];
assign t[25180] = t[25179] ^ n[25180];
assign t[25181] = t[25180] ^ n[25181];
assign t[25182] = t[25181] ^ n[25182];
assign t[25183] = t[25182] ^ n[25183];
assign t[25184] = t[25183] ^ n[25184];
assign t[25185] = t[25184] ^ n[25185];
assign t[25186] = t[25185] ^ n[25186];
assign t[25187] = t[25186] ^ n[25187];
assign t[25188] = t[25187] ^ n[25188];
assign t[25189] = t[25188] ^ n[25189];
assign t[25190] = t[25189] ^ n[25190];
assign t[25191] = t[25190] ^ n[25191];
assign t[25192] = t[25191] ^ n[25192];
assign t[25193] = t[25192] ^ n[25193];
assign t[25194] = t[25193] ^ n[25194];
assign t[25195] = t[25194] ^ n[25195];
assign t[25196] = t[25195] ^ n[25196];
assign t[25197] = t[25196] ^ n[25197];
assign t[25198] = t[25197] ^ n[25198];
assign t[25199] = t[25198] ^ n[25199];
assign t[25200] = t[25199] ^ n[25200];
assign t[25201] = t[25200] ^ n[25201];
assign t[25202] = t[25201] ^ n[25202];
assign t[25203] = t[25202] ^ n[25203];
assign t[25204] = t[25203] ^ n[25204];
assign t[25205] = t[25204] ^ n[25205];
assign t[25206] = t[25205] ^ n[25206];
assign t[25207] = t[25206] ^ n[25207];
assign t[25208] = t[25207] ^ n[25208];
assign t[25209] = t[25208] ^ n[25209];
assign t[25210] = t[25209] ^ n[25210];
assign t[25211] = t[25210] ^ n[25211];
assign t[25212] = t[25211] ^ n[25212];
assign t[25213] = t[25212] ^ n[25213];
assign t[25214] = t[25213] ^ n[25214];
assign t[25215] = t[25214] ^ n[25215];
assign t[25216] = t[25215] ^ n[25216];
assign t[25217] = t[25216] ^ n[25217];
assign t[25218] = t[25217] ^ n[25218];
assign t[25219] = t[25218] ^ n[25219];
assign t[25220] = t[25219] ^ n[25220];
assign t[25221] = t[25220] ^ n[25221];
assign t[25222] = t[25221] ^ n[25222];
assign t[25223] = t[25222] ^ n[25223];
assign t[25224] = t[25223] ^ n[25224];
assign t[25225] = t[25224] ^ n[25225];
assign t[25226] = t[25225] ^ n[25226];
assign t[25227] = t[25226] ^ n[25227];
assign t[25228] = t[25227] ^ n[25228];
assign t[25229] = t[25228] ^ n[25229];
assign t[25230] = t[25229] ^ n[25230];
assign t[25231] = t[25230] ^ n[25231];
assign t[25232] = t[25231] ^ n[25232];
assign t[25233] = t[25232] ^ n[25233];
assign t[25234] = t[25233] ^ n[25234];
assign t[25235] = t[25234] ^ n[25235];
assign t[25236] = t[25235] ^ n[25236];
assign t[25237] = t[25236] ^ n[25237];
assign t[25238] = t[25237] ^ n[25238];
assign t[25239] = t[25238] ^ n[25239];
assign t[25240] = t[25239] ^ n[25240];
assign t[25241] = t[25240] ^ n[25241];
assign t[25242] = t[25241] ^ n[25242];
assign t[25243] = t[25242] ^ n[25243];
assign t[25244] = t[25243] ^ n[25244];
assign t[25245] = t[25244] ^ n[25245];
assign t[25246] = t[25245] ^ n[25246];
assign t[25247] = t[25246] ^ n[25247];
assign t[25248] = t[25247] ^ n[25248];
assign t[25249] = t[25248] ^ n[25249];
assign t[25250] = t[25249] ^ n[25250];
assign t[25251] = t[25250] ^ n[25251];
assign t[25252] = t[25251] ^ n[25252];
assign t[25253] = t[25252] ^ n[25253];
assign t[25254] = t[25253] ^ n[25254];
assign t[25255] = t[25254] ^ n[25255];
assign t[25256] = t[25255] ^ n[25256];
assign t[25257] = t[25256] ^ n[25257];
assign t[25258] = t[25257] ^ n[25258];
assign t[25259] = t[25258] ^ n[25259];
assign t[25260] = t[25259] ^ n[25260];
assign t[25261] = t[25260] ^ n[25261];
assign t[25262] = t[25261] ^ n[25262];
assign t[25263] = t[25262] ^ n[25263];
assign t[25264] = t[25263] ^ n[25264];
assign t[25265] = t[25264] ^ n[25265];
assign t[25266] = t[25265] ^ n[25266];
assign t[25267] = t[25266] ^ n[25267];
assign t[25268] = t[25267] ^ n[25268];
assign t[25269] = t[25268] ^ n[25269];
assign t[25270] = t[25269] ^ n[25270];
assign t[25271] = t[25270] ^ n[25271];
assign t[25272] = t[25271] ^ n[25272];
assign t[25273] = t[25272] ^ n[25273];
assign t[25274] = t[25273] ^ n[25274];
assign t[25275] = t[25274] ^ n[25275];
assign t[25276] = t[25275] ^ n[25276];
assign t[25277] = t[25276] ^ n[25277];
assign t[25278] = t[25277] ^ n[25278];
assign t[25279] = t[25278] ^ n[25279];
assign t[25280] = t[25279] ^ n[25280];
assign t[25281] = t[25280] ^ n[25281];
assign t[25282] = t[25281] ^ n[25282];
assign t[25283] = t[25282] ^ n[25283];
assign t[25284] = t[25283] ^ n[25284];
assign t[25285] = t[25284] ^ n[25285];
assign t[25286] = t[25285] ^ n[25286];
assign t[25287] = t[25286] ^ n[25287];
assign t[25288] = t[25287] ^ n[25288];
assign t[25289] = t[25288] ^ n[25289];
assign t[25290] = t[25289] ^ n[25290];
assign t[25291] = t[25290] ^ n[25291];
assign t[25292] = t[25291] ^ n[25292];
assign t[25293] = t[25292] ^ n[25293];
assign t[25294] = t[25293] ^ n[25294];
assign t[25295] = t[25294] ^ n[25295];
assign t[25296] = t[25295] ^ n[25296];
assign t[25297] = t[25296] ^ n[25297];
assign t[25298] = t[25297] ^ n[25298];
assign t[25299] = t[25298] ^ n[25299];
assign t[25300] = t[25299] ^ n[25300];
assign t[25301] = t[25300] ^ n[25301];
assign t[25302] = t[25301] ^ n[25302];
assign t[25303] = t[25302] ^ n[25303];
assign t[25304] = t[25303] ^ n[25304];
assign t[25305] = t[25304] ^ n[25305];
assign t[25306] = t[25305] ^ n[25306];
assign t[25307] = t[25306] ^ n[25307];
assign t[25308] = t[25307] ^ n[25308];
assign t[25309] = t[25308] ^ n[25309];
assign t[25310] = t[25309] ^ n[25310];
assign t[25311] = t[25310] ^ n[25311];
assign t[25312] = t[25311] ^ n[25312];
assign t[25313] = t[25312] ^ n[25313];
assign t[25314] = t[25313] ^ n[25314];
assign t[25315] = t[25314] ^ n[25315];
assign t[25316] = t[25315] ^ n[25316];
assign t[25317] = t[25316] ^ n[25317];
assign t[25318] = t[25317] ^ n[25318];
assign t[25319] = t[25318] ^ n[25319];
assign t[25320] = t[25319] ^ n[25320];
assign t[25321] = t[25320] ^ n[25321];
assign t[25322] = t[25321] ^ n[25322];
assign t[25323] = t[25322] ^ n[25323];
assign t[25324] = t[25323] ^ n[25324];
assign t[25325] = t[25324] ^ n[25325];
assign t[25326] = t[25325] ^ n[25326];
assign t[25327] = t[25326] ^ n[25327];
assign t[25328] = t[25327] ^ n[25328];
assign t[25329] = t[25328] ^ n[25329];
assign t[25330] = t[25329] ^ n[25330];
assign t[25331] = t[25330] ^ n[25331];
assign t[25332] = t[25331] ^ n[25332];
assign t[25333] = t[25332] ^ n[25333];
assign t[25334] = t[25333] ^ n[25334];
assign t[25335] = t[25334] ^ n[25335];
assign t[25336] = t[25335] ^ n[25336];
assign t[25337] = t[25336] ^ n[25337];
assign t[25338] = t[25337] ^ n[25338];
assign t[25339] = t[25338] ^ n[25339];
assign t[25340] = t[25339] ^ n[25340];
assign t[25341] = t[25340] ^ n[25341];
assign t[25342] = t[25341] ^ n[25342];
assign t[25343] = t[25342] ^ n[25343];
assign t[25344] = t[25343] ^ n[25344];
assign t[25345] = t[25344] ^ n[25345];
assign t[25346] = t[25345] ^ n[25346];
assign t[25347] = t[25346] ^ n[25347];
assign t[25348] = t[25347] ^ n[25348];
assign t[25349] = t[25348] ^ n[25349];
assign t[25350] = t[25349] ^ n[25350];
assign t[25351] = t[25350] ^ n[25351];
assign t[25352] = t[25351] ^ n[25352];
assign t[25353] = t[25352] ^ n[25353];
assign t[25354] = t[25353] ^ n[25354];
assign t[25355] = t[25354] ^ n[25355];
assign t[25356] = t[25355] ^ n[25356];
assign t[25357] = t[25356] ^ n[25357];
assign t[25358] = t[25357] ^ n[25358];
assign t[25359] = t[25358] ^ n[25359];
assign t[25360] = t[25359] ^ n[25360];
assign t[25361] = t[25360] ^ n[25361];
assign t[25362] = t[25361] ^ n[25362];
assign t[25363] = t[25362] ^ n[25363];
assign t[25364] = t[25363] ^ n[25364];
assign t[25365] = t[25364] ^ n[25365];
assign t[25366] = t[25365] ^ n[25366];
assign t[25367] = t[25366] ^ n[25367];
assign t[25368] = t[25367] ^ n[25368];
assign t[25369] = t[25368] ^ n[25369];
assign t[25370] = t[25369] ^ n[25370];
assign t[25371] = t[25370] ^ n[25371];
assign t[25372] = t[25371] ^ n[25372];
assign t[25373] = t[25372] ^ n[25373];
assign t[25374] = t[25373] ^ n[25374];
assign t[25375] = t[25374] ^ n[25375];
assign t[25376] = t[25375] ^ n[25376];
assign t[25377] = t[25376] ^ n[25377];
assign t[25378] = t[25377] ^ n[25378];
assign t[25379] = t[25378] ^ n[25379];
assign t[25380] = t[25379] ^ n[25380];
assign t[25381] = t[25380] ^ n[25381];
assign t[25382] = t[25381] ^ n[25382];
assign t[25383] = t[25382] ^ n[25383];
assign t[25384] = t[25383] ^ n[25384];
assign t[25385] = t[25384] ^ n[25385];
assign t[25386] = t[25385] ^ n[25386];
assign t[25387] = t[25386] ^ n[25387];
assign t[25388] = t[25387] ^ n[25388];
assign t[25389] = t[25388] ^ n[25389];
assign t[25390] = t[25389] ^ n[25390];
assign t[25391] = t[25390] ^ n[25391];
assign t[25392] = t[25391] ^ n[25392];
assign t[25393] = t[25392] ^ n[25393];
assign t[25394] = t[25393] ^ n[25394];
assign t[25395] = t[25394] ^ n[25395];
assign t[25396] = t[25395] ^ n[25396];
assign t[25397] = t[25396] ^ n[25397];
assign t[25398] = t[25397] ^ n[25398];
assign t[25399] = t[25398] ^ n[25399];
assign t[25400] = t[25399] ^ n[25400];
assign t[25401] = t[25400] ^ n[25401];
assign t[25402] = t[25401] ^ n[25402];
assign t[25403] = t[25402] ^ n[25403];
assign t[25404] = t[25403] ^ n[25404];
assign t[25405] = t[25404] ^ n[25405];
assign t[25406] = t[25405] ^ n[25406];
assign t[25407] = t[25406] ^ n[25407];
assign t[25408] = t[25407] ^ n[25408];
assign t[25409] = t[25408] ^ n[25409];
assign t[25410] = t[25409] ^ n[25410];
assign t[25411] = t[25410] ^ n[25411];
assign t[25412] = t[25411] ^ n[25412];
assign t[25413] = t[25412] ^ n[25413];
assign t[25414] = t[25413] ^ n[25414];
assign t[25415] = t[25414] ^ n[25415];
assign t[25416] = t[25415] ^ n[25416];
assign t[25417] = t[25416] ^ n[25417];
assign t[25418] = t[25417] ^ n[25418];
assign t[25419] = t[25418] ^ n[25419];
assign t[25420] = t[25419] ^ n[25420];
assign t[25421] = t[25420] ^ n[25421];
assign t[25422] = t[25421] ^ n[25422];
assign t[25423] = t[25422] ^ n[25423];
assign t[25424] = t[25423] ^ n[25424];
assign t[25425] = t[25424] ^ n[25425];
assign t[25426] = t[25425] ^ n[25426];
assign t[25427] = t[25426] ^ n[25427];
assign t[25428] = t[25427] ^ n[25428];
assign t[25429] = t[25428] ^ n[25429];
assign t[25430] = t[25429] ^ n[25430];
assign t[25431] = t[25430] ^ n[25431];
assign t[25432] = t[25431] ^ n[25432];
assign t[25433] = t[25432] ^ n[25433];
assign t[25434] = t[25433] ^ n[25434];
assign t[25435] = t[25434] ^ n[25435];
assign t[25436] = t[25435] ^ n[25436];
assign t[25437] = t[25436] ^ n[25437];
assign t[25438] = t[25437] ^ n[25438];
assign t[25439] = t[25438] ^ n[25439];
assign t[25440] = t[25439] ^ n[25440];
assign t[25441] = t[25440] ^ n[25441];
assign t[25442] = t[25441] ^ n[25442];
assign t[25443] = t[25442] ^ n[25443];
assign t[25444] = t[25443] ^ n[25444];
assign t[25445] = t[25444] ^ n[25445];
assign t[25446] = t[25445] ^ n[25446];
assign t[25447] = t[25446] ^ n[25447];
assign t[25448] = t[25447] ^ n[25448];
assign t[25449] = t[25448] ^ n[25449];
assign t[25450] = t[25449] ^ n[25450];
assign t[25451] = t[25450] ^ n[25451];
assign t[25452] = t[25451] ^ n[25452];
assign t[25453] = t[25452] ^ n[25453];
assign t[25454] = t[25453] ^ n[25454];
assign t[25455] = t[25454] ^ n[25455];
assign t[25456] = t[25455] ^ n[25456];
assign t[25457] = t[25456] ^ n[25457];
assign t[25458] = t[25457] ^ n[25458];
assign t[25459] = t[25458] ^ n[25459];
assign t[25460] = t[25459] ^ n[25460];
assign t[25461] = t[25460] ^ n[25461];
assign t[25462] = t[25461] ^ n[25462];
assign t[25463] = t[25462] ^ n[25463];
assign t[25464] = t[25463] ^ n[25464];
assign t[25465] = t[25464] ^ n[25465];
assign t[25466] = t[25465] ^ n[25466];
assign t[25467] = t[25466] ^ n[25467];
assign t[25468] = t[25467] ^ n[25468];
assign t[25469] = t[25468] ^ n[25469];
assign t[25470] = t[25469] ^ n[25470];
assign t[25471] = t[25470] ^ n[25471];
assign t[25472] = t[25471] ^ n[25472];
assign t[25473] = t[25472] ^ n[25473];
assign t[25474] = t[25473] ^ n[25474];
assign t[25475] = t[25474] ^ n[25475];
assign t[25476] = t[25475] ^ n[25476];
assign t[25477] = t[25476] ^ n[25477];
assign t[25478] = t[25477] ^ n[25478];
assign t[25479] = t[25478] ^ n[25479];
assign t[25480] = t[25479] ^ n[25480];
assign t[25481] = t[25480] ^ n[25481];
assign t[25482] = t[25481] ^ n[25482];
assign t[25483] = t[25482] ^ n[25483];
assign t[25484] = t[25483] ^ n[25484];
assign t[25485] = t[25484] ^ n[25485];
assign t[25486] = t[25485] ^ n[25486];
assign t[25487] = t[25486] ^ n[25487];
assign t[25488] = t[25487] ^ n[25488];
assign t[25489] = t[25488] ^ n[25489];
assign t[25490] = t[25489] ^ n[25490];
assign t[25491] = t[25490] ^ n[25491];
assign t[25492] = t[25491] ^ n[25492];
assign t[25493] = t[25492] ^ n[25493];
assign t[25494] = t[25493] ^ n[25494];
assign t[25495] = t[25494] ^ n[25495];
assign t[25496] = t[25495] ^ n[25496];
assign t[25497] = t[25496] ^ n[25497];
assign t[25498] = t[25497] ^ n[25498];
assign t[25499] = t[25498] ^ n[25499];
assign t[25500] = t[25499] ^ n[25500];
assign t[25501] = t[25500] ^ n[25501];
assign t[25502] = t[25501] ^ n[25502];
assign t[25503] = t[25502] ^ n[25503];
assign t[25504] = t[25503] ^ n[25504];
assign t[25505] = t[25504] ^ n[25505];
assign t[25506] = t[25505] ^ n[25506];
assign t[25507] = t[25506] ^ n[25507];
assign t[25508] = t[25507] ^ n[25508];
assign t[25509] = t[25508] ^ n[25509];
assign t[25510] = t[25509] ^ n[25510];
assign t[25511] = t[25510] ^ n[25511];
assign t[25512] = t[25511] ^ n[25512];
assign t[25513] = t[25512] ^ n[25513];
assign t[25514] = t[25513] ^ n[25514];
assign t[25515] = t[25514] ^ n[25515];
assign t[25516] = t[25515] ^ n[25516];
assign t[25517] = t[25516] ^ n[25517];
assign t[25518] = t[25517] ^ n[25518];
assign t[25519] = t[25518] ^ n[25519];
assign t[25520] = t[25519] ^ n[25520];
assign t[25521] = t[25520] ^ n[25521];
assign t[25522] = t[25521] ^ n[25522];
assign t[25523] = t[25522] ^ n[25523];
assign t[25524] = t[25523] ^ n[25524];
assign t[25525] = t[25524] ^ n[25525];
assign t[25526] = t[25525] ^ n[25526];
assign t[25527] = t[25526] ^ n[25527];
assign t[25528] = t[25527] ^ n[25528];
assign t[25529] = t[25528] ^ n[25529];
assign t[25530] = t[25529] ^ n[25530];
assign t[25531] = t[25530] ^ n[25531];
assign t[25532] = t[25531] ^ n[25532];
assign t[25533] = t[25532] ^ n[25533];
assign t[25534] = t[25533] ^ n[25534];
assign t[25535] = t[25534] ^ n[25535];
assign t[25536] = t[25535] ^ n[25536];
assign t[25537] = t[25536] ^ n[25537];
assign t[25538] = t[25537] ^ n[25538];
assign t[25539] = t[25538] ^ n[25539];
assign t[25540] = t[25539] ^ n[25540];
assign t[25541] = t[25540] ^ n[25541];
assign t[25542] = t[25541] ^ n[25542];
assign t[25543] = t[25542] ^ n[25543];
assign t[25544] = t[25543] ^ n[25544];
assign t[25545] = t[25544] ^ n[25545];
assign t[25546] = t[25545] ^ n[25546];
assign t[25547] = t[25546] ^ n[25547];
assign t[25548] = t[25547] ^ n[25548];
assign t[25549] = t[25548] ^ n[25549];
assign t[25550] = t[25549] ^ n[25550];
assign t[25551] = t[25550] ^ n[25551];
assign t[25552] = t[25551] ^ n[25552];
assign t[25553] = t[25552] ^ n[25553];
assign t[25554] = t[25553] ^ n[25554];
assign t[25555] = t[25554] ^ n[25555];
assign t[25556] = t[25555] ^ n[25556];
assign t[25557] = t[25556] ^ n[25557];
assign t[25558] = t[25557] ^ n[25558];
assign t[25559] = t[25558] ^ n[25559];
assign t[25560] = t[25559] ^ n[25560];
assign t[25561] = t[25560] ^ n[25561];
assign t[25562] = t[25561] ^ n[25562];
assign t[25563] = t[25562] ^ n[25563];
assign t[25564] = t[25563] ^ n[25564];
assign t[25565] = t[25564] ^ n[25565];
assign t[25566] = t[25565] ^ n[25566];
assign t[25567] = t[25566] ^ n[25567];
assign t[25568] = t[25567] ^ n[25568];
assign t[25569] = t[25568] ^ n[25569];
assign t[25570] = t[25569] ^ n[25570];
assign t[25571] = t[25570] ^ n[25571];
assign t[25572] = t[25571] ^ n[25572];
assign t[25573] = t[25572] ^ n[25573];
assign t[25574] = t[25573] ^ n[25574];
assign t[25575] = t[25574] ^ n[25575];
assign t[25576] = t[25575] ^ n[25576];
assign t[25577] = t[25576] ^ n[25577];
assign t[25578] = t[25577] ^ n[25578];
assign t[25579] = t[25578] ^ n[25579];
assign t[25580] = t[25579] ^ n[25580];
assign t[25581] = t[25580] ^ n[25581];
assign t[25582] = t[25581] ^ n[25582];
assign t[25583] = t[25582] ^ n[25583];
assign t[25584] = t[25583] ^ n[25584];
assign t[25585] = t[25584] ^ n[25585];
assign t[25586] = t[25585] ^ n[25586];
assign t[25587] = t[25586] ^ n[25587];
assign t[25588] = t[25587] ^ n[25588];
assign t[25589] = t[25588] ^ n[25589];
assign t[25590] = t[25589] ^ n[25590];
assign t[25591] = t[25590] ^ n[25591];
assign t[25592] = t[25591] ^ n[25592];
assign t[25593] = t[25592] ^ n[25593];
assign t[25594] = t[25593] ^ n[25594];
assign t[25595] = t[25594] ^ n[25595];
assign t[25596] = t[25595] ^ n[25596];
assign t[25597] = t[25596] ^ n[25597];
assign t[25598] = t[25597] ^ n[25598];
assign t[25599] = t[25598] ^ n[25599];
assign t[25600] = t[25599] ^ n[25600];
assign t[25601] = t[25600] ^ n[25601];
assign t[25602] = t[25601] ^ n[25602];
assign t[25603] = t[25602] ^ n[25603];
assign t[25604] = t[25603] ^ n[25604];
assign t[25605] = t[25604] ^ n[25605];
assign t[25606] = t[25605] ^ n[25606];
assign t[25607] = t[25606] ^ n[25607];
assign t[25608] = t[25607] ^ n[25608];
assign t[25609] = t[25608] ^ n[25609];
assign t[25610] = t[25609] ^ n[25610];
assign t[25611] = t[25610] ^ n[25611];
assign t[25612] = t[25611] ^ n[25612];
assign t[25613] = t[25612] ^ n[25613];
assign t[25614] = t[25613] ^ n[25614];
assign t[25615] = t[25614] ^ n[25615];
assign t[25616] = t[25615] ^ n[25616];
assign t[25617] = t[25616] ^ n[25617];
assign t[25618] = t[25617] ^ n[25618];
assign t[25619] = t[25618] ^ n[25619];
assign t[25620] = t[25619] ^ n[25620];
assign t[25621] = t[25620] ^ n[25621];
assign t[25622] = t[25621] ^ n[25622];
assign t[25623] = t[25622] ^ n[25623];
assign t[25624] = t[25623] ^ n[25624];
assign t[25625] = t[25624] ^ n[25625];
assign t[25626] = t[25625] ^ n[25626];
assign t[25627] = t[25626] ^ n[25627];
assign t[25628] = t[25627] ^ n[25628];
assign t[25629] = t[25628] ^ n[25629];
assign t[25630] = t[25629] ^ n[25630];
assign t[25631] = t[25630] ^ n[25631];
assign t[25632] = t[25631] ^ n[25632];
assign t[25633] = t[25632] ^ n[25633];
assign t[25634] = t[25633] ^ n[25634];
assign t[25635] = t[25634] ^ n[25635];
assign t[25636] = t[25635] ^ n[25636];
assign t[25637] = t[25636] ^ n[25637];
assign t[25638] = t[25637] ^ n[25638];
assign t[25639] = t[25638] ^ n[25639];
assign t[25640] = t[25639] ^ n[25640];
assign t[25641] = t[25640] ^ n[25641];
assign t[25642] = t[25641] ^ n[25642];
assign t[25643] = t[25642] ^ n[25643];
assign t[25644] = t[25643] ^ n[25644];
assign t[25645] = t[25644] ^ n[25645];
assign t[25646] = t[25645] ^ n[25646];
assign t[25647] = t[25646] ^ n[25647];
assign t[25648] = t[25647] ^ n[25648];
assign t[25649] = t[25648] ^ n[25649];
assign t[25650] = t[25649] ^ n[25650];
assign t[25651] = t[25650] ^ n[25651];
assign t[25652] = t[25651] ^ n[25652];
assign t[25653] = t[25652] ^ n[25653];
assign t[25654] = t[25653] ^ n[25654];
assign t[25655] = t[25654] ^ n[25655];
assign t[25656] = t[25655] ^ n[25656];
assign t[25657] = t[25656] ^ n[25657];
assign t[25658] = t[25657] ^ n[25658];
assign t[25659] = t[25658] ^ n[25659];
assign t[25660] = t[25659] ^ n[25660];
assign t[25661] = t[25660] ^ n[25661];
assign t[25662] = t[25661] ^ n[25662];
assign t[25663] = t[25662] ^ n[25663];
assign t[25664] = t[25663] ^ n[25664];
assign t[25665] = t[25664] ^ n[25665];
assign t[25666] = t[25665] ^ n[25666];
assign t[25667] = t[25666] ^ n[25667];
assign t[25668] = t[25667] ^ n[25668];
assign t[25669] = t[25668] ^ n[25669];
assign t[25670] = t[25669] ^ n[25670];
assign t[25671] = t[25670] ^ n[25671];
assign t[25672] = t[25671] ^ n[25672];
assign t[25673] = t[25672] ^ n[25673];
assign t[25674] = t[25673] ^ n[25674];
assign t[25675] = t[25674] ^ n[25675];
assign t[25676] = t[25675] ^ n[25676];
assign t[25677] = t[25676] ^ n[25677];
assign t[25678] = t[25677] ^ n[25678];
assign t[25679] = t[25678] ^ n[25679];
assign t[25680] = t[25679] ^ n[25680];
assign t[25681] = t[25680] ^ n[25681];
assign t[25682] = t[25681] ^ n[25682];
assign t[25683] = t[25682] ^ n[25683];
assign t[25684] = t[25683] ^ n[25684];
assign t[25685] = t[25684] ^ n[25685];
assign t[25686] = t[25685] ^ n[25686];
assign t[25687] = t[25686] ^ n[25687];
assign t[25688] = t[25687] ^ n[25688];
assign t[25689] = t[25688] ^ n[25689];
assign t[25690] = t[25689] ^ n[25690];
assign t[25691] = t[25690] ^ n[25691];
assign t[25692] = t[25691] ^ n[25692];
assign t[25693] = t[25692] ^ n[25693];
assign t[25694] = t[25693] ^ n[25694];
assign t[25695] = t[25694] ^ n[25695];
assign t[25696] = t[25695] ^ n[25696];
assign t[25697] = t[25696] ^ n[25697];
assign t[25698] = t[25697] ^ n[25698];
assign t[25699] = t[25698] ^ n[25699];
assign t[25700] = t[25699] ^ n[25700];
assign t[25701] = t[25700] ^ n[25701];
assign t[25702] = t[25701] ^ n[25702];
assign t[25703] = t[25702] ^ n[25703];
assign t[25704] = t[25703] ^ n[25704];
assign t[25705] = t[25704] ^ n[25705];
assign t[25706] = t[25705] ^ n[25706];
assign t[25707] = t[25706] ^ n[25707];
assign t[25708] = t[25707] ^ n[25708];
assign t[25709] = t[25708] ^ n[25709];
assign t[25710] = t[25709] ^ n[25710];
assign t[25711] = t[25710] ^ n[25711];
assign t[25712] = t[25711] ^ n[25712];
assign t[25713] = t[25712] ^ n[25713];
assign t[25714] = t[25713] ^ n[25714];
assign t[25715] = t[25714] ^ n[25715];
assign t[25716] = t[25715] ^ n[25716];
assign t[25717] = t[25716] ^ n[25717];
assign t[25718] = t[25717] ^ n[25718];
assign t[25719] = t[25718] ^ n[25719];
assign t[25720] = t[25719] ^ n[25720];
assign t[25721] = t[25720] ^ n[25721];
assign t[25722] = t[25721] ^ n[25722];
assign t[25723] = t[25722] ^ n[25723];
assign t[25724] = t[25723] ^ n[25724];
assign t[25725] = t[25724] ^ n[25725];
assign t[25726] = t[25725] ^ n[25726];
assign t[25727] = t[25726] ^ n[25727];
assign t[25728] = t[25727] ^ n[25728];
assign t[25729] = t[25728] ^ n[25729];
assign t[25730] = t[25729] ^ n[25730];
assign t[25731] = t[25730] ^ n[25731];
assign t[25732] = t[25731] ^ n[25732];
assign t[25733] = t[25732] ^ n[25733];
assign t[25734] = t[25733] ^ n[25734];
assign t[25735] = t[25734] ^ n[25735];
assign t[25736] = t[25735] ^ n[25736];
assign t[25737] = t[25736] ^ n[25737];
assign t[25738] = t[25737] ^ n[25738];
assign t[25739] = t[25738] ^ n[25739];
assign t[25740] = t[25739] ^ n[25740];
assign t[25741] = t[25740] ^ n[25741];
assign t[25742] = t[25741] ^ n[25742];
assign t[25743] = t[25742] ^ n[25743];
assign t[25744] = t[25743] ^ n[25744];
assign t[25745] = t[25744] ^ n[25745];
assign t[25746] = t[25745] ^ n[25746];
assign t[25747] = t[25746] ^ n[25747];
assign t[25748] = t[25747] ^ n[25748];
assign t[25749] = t[25748] ^ n[25749];
assign t[25750] = t[25749] ^ n[25750];
assign t[25751] = t[25750] ^ n[25751];
assign t[25752] = t[25751] ^ n[25752];
assign t[25753] = t[25752] ^ n[25753];
assign t[25754] = t[25753] ^ n[25754];
assign t[25755] = t[25754] ^ n[25755];
assign t[25756] = t[25755] ^ n[25756];
assign t[25757] = t[25756] ^ n[25757];
assign t[25758] = t[25757] ^ n[25758];
assign t[25759] = t[25758] ^ n[25759];
assign t[25760] = t[25759] ^ n[25760];
assign t[25761] = t[25760] ^ n[25761];
assign t[25762] = t[25761] ^ n[25762];
assign t[25763] = t[25762] ^ n[25763];
assign t[25764] = t[25763] ^ n[25764];
assign t[25765] = t[25764] ^ n[25765];
assign t[25766] = t[25765] ^ n[25766];
assign t[25767] = t[25766] ^ n[25767];
assign t[25768] = t[25767] ^ n[25768];
assign t[25769] = t[25768] ^ n[25769];
assign t[25770] = t[25769] ^ n[25770];
assign t[25771] = t[25770] ^ n[25771];
assign t[25772] = t[25771] ^ n[25772];
assign t[25773] = t[25772] ^ n[25773];
assign t[25774] = t[25773] ^ n[25774];
assign t[25775] = t[25774] ^ n[25775];
assign t[25776] = t[25775] ^ n[25776];
assign t[25777] = t[25776] ^ n[25777];
assign t[25778] = t[25777] ^ n[25778];
assign t[25779] = t[25778] ^ n[25779];
assign t[25780] = t[25779] ^ n[25780];
assign t[25781] = t[25780] ^ n[25781];
assign t[25782] = t[25781] ^ n[25782];
assign t[25783] = t[25782] ^ n[25783];
assign t[25784] = t[25783] ^ n[25784];
assign t[25785] = t[25784] ^ n[25785];
assign t[25786] = t[25785] ^ n[25786];
assign t[25787] = t[25786] ^ n[25787];
assign t[25788] = t[25787] ^ n[25788];
assign t[25789] = t[25788] ^ n[25789];
assign t[25790] = t[25789] ^ n[25790];
assign t[25791] = t[25790] ^ n[25791];
assign t[25792] = t[25791] ^ n[25792];
assign t[25793] = t[25792] ^ n[25793];
assign t[25794] = t[25793] ^ n[25794];
assign t[25795] = t[25794] ^ n[25795];
assign t[25796] = t[25795] ^ n[25796];
assign t[25797] = t[25796] ^ n[25797];
assign t[25798] = t[25797] ^ n[25798];
assign t[25799] = t[25798] ^ n[25799];
assign t[25800] = t[25799] ^ n[25800];
assign t[25801] = t[25800] ^ n[25801];
assign t[25802] = t[25801] ^ n[25802];
assign t[25803] = t[25802] ^ n[25803];
assign t[25804] = t[25803] ^ n[25804];
assign t[25805] = t[25804] ^ n[25805];
assign t[25806] = t[25805] ^ n[25806];
assign t[25807] = t[25806] ^ n[25807];
assign t[25808] = t[25807] ^ n[25808];
assign t[25809] = t[25808] ^ n[25809];
assign t[25810] = t[25809] ^ n[25810];
assign t[25811] = t[25810] ^ n[25811];
assign t[25812] = t[25811] ^ n[25812];
assign t[25813] = t[25812] ^ n[25813];
assign t[25814] = t[25813] ^ n[25814];
assign t[25815] = t[25814] ^ n[25815];
assign t[25816] = t[25815] ^ n[25816];
assign t[25817] = t[25816] ^ n[25817];
assign t[25818] = t[25817] ^ n[25818];
assign t[25819] = t[25818] ^ n[25819];
assign t[25820] = t[25819] ^ n[25820];
assign t[25821] = t[25820] ^ n[25821];
assign t[25822] = t[25821] ^ n[25822];
assign t[25823] = t[25822] ^ n[25823];
assign t[25824] = t[25823] ^ n[25824];
assign t[25825] = t[25824] ^ n[25825];
assign t[25826] = t[25825] ^ n[25826];
assign t[25827] = t[25826] ^ n[25827];
assign t[25828] = t[25827] ^ n[25828];
assign t[25829] = t[25828] ^ n[25829];
assign t[25830] = t[25829] ^ n[25830];
assign t[25831] = t[25830] ^ n[25831];
assign t[25832] = t[25831] ^ n[25832];
assign t[25833] = t[25832] ^ n[25833];
assign t[25834] = t[25833] ^ n[25834];
assign t[25835] = t[25834] ^ n[25835];
assign t[25836] = t[25835] ^ n[25836];
assign t[25837] = t[25836] ^ n[25837];
assign t[25838] = t[25837] ^ n[25838];
assign t[25839] = t[25838] ^ n[25839];
assign t[25840] = t[25839] ^ n[25840];
assign t[25841] = t[25840] ^ n[25841];
assign t[25842] = t[25841] ^ n[25842];
assign t[25843] = t[25842] ^ n[25843];
assign t[25844] = t[25843] ^ n[25844];
assign t[25845] = t[25844] ^ n[25845];
assign t[25846] = t[25845] ^ n[25846];
assign t[25847] = t[25846] ^ n[25847];
assign t[25848] = t[25847] ^ n[25848];
assign t[25849] = t[25848] ^ n[25849];
assign t[25850] = t[25849] ^ n[25850];
assign t[25851] = t[25850] ^ n[25851];
assign t[25852] = t[25851] ^ n[25852];
assign t[25853] = t[25852] ^ n[25853];
assign t[25854] = t[25853] ^ n[25854];
assign t[25855] = t[25854] ^ n[25855];
assign t[25856] = t[25855] ^ n[25856];
assign t[25857] = t[25856] ^ n[25857];
assign t[25858] = t[25857] ^ n[25858];
assign t[25859] = t[25858] ^ n[25859];
assign t[25860] = t[25859] ^ n[25860];
assign t[25861] = t[25860] ^ n[25861];
assign t[25862] = t[25861] ^ n[25862];
assign t[25863] = t[25862] ^ n[25863];
assign t[25864] = t[25863] ^ n[25864];
assign t[25865] = t[25864] ^ n[25865];
assign t[25866] = t[25865] ^ n[25866];
assign t[25867] = t[25866] ^ n[25867];
assign t[25868] = t[25867] ^ n[25868];
assign t[25869] = t[25868] ^ n[25869];
assign t[25870] = t[25869] ^ n[25870];
assign t[25871] = t[25870] ^ n[25871];
assign t[25872] = t[25871] ^ n[25872];
assign t[25873] = t[25872] ^ n[25873];
assign t[25874] = t[25873] ^ n[25874];
assign t[25875] = t[25874] ^ n[25875];
assign t[25876] = t[25875] ^ n[25876];
assign t[25877] = t[25876] ^ n[25877];
assign t[25878] = t[25877] ^ n[25878];
assign t[25879] = t[25878] ^ n[25879];
assign t[25880] = t[25879] ^ n[25880];
assign t[25881] = t[25880] ^ n[25881];
assign t[25882] = t[25881] ^ n[25882];
assign t[25883] = t[25882] ^ n[25883];
assign t[25884] = t[25883] ^ n[25884];
assign t[25885] = t[25884] ^ n[25885];
assign t[25886] = t[25885] ^ n[25886];
assign t[25887] = t[25886] ^ n[25887];
assign t[25888] = t[25887] ^ n[25888];
assign t[25889] = t[25888] ^ n[25889];
assign t[25890] = t[25889] ^ n[25890];
assign t[25891] = t[25890] ^ n[25891];
assign t[25892] = t[25891] ^ n[25892];
assign t[25893] = t[25892] ^ n[25893];
assign t[25894] = t[25893] ^ n[25894];
assign t[25895] = t[25894] ^ n[25895];
assign t[25896] = t[25895] ^ n[25896];
assign t[25897] = t[25896] ^ n[25897];
assign t[25898] = t[25897] ^ n[25898];
assign t[25899] = t[25898] ^ n[25899];
assign t[25900] = t[25899] ^ n[25900];
assign t[25901] = t[25900] ^ n[25901];
assign t[25902] = t[25901] ^ n[25902];
assign t[25903] = t[25902] ^ n[25903];
assign t[25904] = t[25903] ^ n[25904];
assign t[25905] = t[25904] ^ n[25905];
assign t[25906] = t[25905] ^ n[25906];
assign t[25907] = t[25906] ^ n[25907];
assign t[25908] = t[25907] ^ n[25908];
assign t[25909] = t[25908] ^ n[25909];
assign t[25910] = t[25909] ^ n[25910];
assign t[25911] = t[25910] ^ n[25911];
assign t[25912] = t[25911] ^ n[25912];
assign t[25913] = t[25912] ^ n[25913];
assign t[25914] = t[25913] ^ n[25914];
assign t[25915] = t[25914] ^ n[25915];
assign t[25916] = t[25915] ^ n[25916];
assign t[25917] = t[25916] ^ n[25917];
assign t[25918] = t[25917] ^ n[25918];
assign t[25919] = t[25918] ^ n[25919];
assign t[25920] = t[25919] ^ n[25920];
assign t[25921] = t[25920] ^ n[25921];
assign t[25922] = t[25921] ^ n[25922];
assign t[25923] = t[25922] ^ n[25923];
assign t[25924] = t[25923] ^ n[25924];
assign t[25925] = t[25924] ^ n[25925];
assign t[25926] = t[25925] ^ n[25926];
assign t[25927] = t[25926] ^ n[25927];
assign t[25928] = t[25927] ^ n[25928];
assign t[25929] = t[25928] ^ n[25929];
assign t[25930] = t[25929] ^ n[25930];
assign t[25931] = t[25930] ^ n[25931];
assign t[25932] = t[25931] ^ n[25932];
assign t[25933] = t[25932] ^ n[25933];
assign t[25934] = t[25933] ^ n[25934];
assign t[25935] = t[25934] ^ n[25935];
assign t[25936] = t[25935] ^ n[25936];
assign t[25937] = t[25936] ^ n[25937];
assign t[25938] = t[25937] ^ n[25938];
assign t[25939] = t[25938] ^ n[25939];
assign t[25940] = t[25939] ^ n[25940];
assign t[25941] = t[25940] ^ n[25941];
assign t[25942] = t[25941] ^ n[25942];
assign t[25943] = t[25942] ^ n[25943];
assign t[25944] = t[25943] ^ n[25944];
assign t[25945] = t[25944] ^ n[25945];
assign t[25946] = t[25945] ^ n[25946];
assign t[25947] = t[25946] ^ n[25947];
assign t[25948] = t[25947] ^ n[25948];
assign t[25949] = t[25948] ^ n[25949];
assign t[25950] = t[25949] ^ n[25950];
assign t[25951] = t[25950] ^ n[25951];
assign t[25952] = t[25951] ^ n[25952];
assign t[25953] = t[25952] ^ n[25953];
assign t[25954] = t[25953] ^ n[25954];
assign t[25955] = t[25954] ^ n[25955];
assign t[25956] = t[25955] ^ n[25956];
assign t[25957] = t[25956] ^ n[25957];
assign t[25958] = t[25957] ^ n[25958];
assign t[25959] = t[25958] ^ n[25959];
assign t[25960] = t[25959] ^ n[25960];
assign t[25961] = t[25960] ^ n[25961];
assign t[25962] = t[25961] ^ n[25962];
assign t[25963] = t[25962] ^ n[25963];
assign t[25964] = t[25963] ^ n[25964];
assign t[25965] = t[25964] ^ n[25965];
assign t[25966] = t[25965] ^ n[25966];
assign t[25967] = t[25966] ^ n[25967];
assign t[25968] = t[25967] ^ n[25968];
assign t[25969] = t[25968] ^ n[25969];
assign t[25970] = t[25969] ^ n[25970];
assign t[25971] = t[25970] ^ n[25971];
assign t[25972] = t[25971] ^ n[25972];
assign t[25973] = t[25972] ^ n[25973];
assign t[25974] = t[25973] ^ n[25974];
assign t[25975] = t[25974] ^ n[25975];
assign t[25976] = t[25975] ^ n[25976];
assign t[25977] = t[25976] ^ n[25977];
assign t[25978] = t[25977] ^ n[25978];
assign t[25979] = t[25978] ^ n[25979];
assign t[25980] = t[25979] ^ n[25980];
assign t[25981] = t[25980] ^ n[25981];
assign t[25982] = t[25981] ^ n[25982];
assign t[25983] = t[25982] ^ n[25983];
assign t[25984] = t[25983] ^ n[25984];
assign t[25985] = t[25984] ^ n[25985];
assign t[25986] = t[25985] ^ n[25986];
assign t[25987] = t[25986] ^ n[25987];
assign t[25988] = t[25987] ^ n[25988];
assign t[25989] = t[25988] ^ n[25989];
assign t[25990] = t[25989] ^ n[25990];
assign t[25991] = t[25990] ^ n[25991];
assign t[25992] = t[25991] ^ n[25992];
assign t[25993] = t[25992] ^ n[25993];
assign t[25994] = t[25993] ^ n[25994];
assign t[25995] = t[25994] ^ n[25995];
assign t[25996] = t[25995] ^ n[25996];
assign t[25997] = t[25996] ^ n[25997];
assign t[25998] = t[25997] ^ n[25998];
assign t[25999] = t[25998] ^ n[25999];
assign t[26000] = t[25999] ^ n[26000];
assign t[26001] = t[26000] ^ n[26001];
assign t[26002] = t[26001] ^ n[26002];
assign t[26003] = t[26002] ^ n[26003];
assign t[26004] = t[26003] ^ n[26004];
assign t[26005] = t[26004] ^ n[26005];
assign t[26006] = t[26005] ^ n[26006];
assign t[26007] = t[26006] ^ n[26007];
assign t[26008] = t[26007] ^ n[26008];
assign t[26009] = t[26008] ^ n[26009];
assign t[26010] = t[26009] ^ n[26010];
assign t[26011] = t[26010] ^ n[26011];
assign t[26012] = t[26011] ^ n[26012];
assign t[26013] = t[26012] ^ n[26013];
assign t[26014] = t[26013] ^ n[26014];
assign t[26015] = t[26014] ^ n[26015];
assign t[26016] = t[26015] ^ n[26016];
assign t[26017] = t[26016] ^ n[26017];
assign t[26018] = t[26017] ^ n[26018];
assign t[26019] = t[26018] ^ n[26019];
assign t[26020] = t[26019] ^ n[26020];
assign t[26021] = t[26020] ^ n[26021];
assign t[26022] = t[26021] ^ n[26022];
assign t[26023] = t[26022] ^ n[26023];
assign t[26024] = t[26023] ^ n[26024];
assign t[26025] = t[26024] ^ n[26025];
assign t[26026] = t[26025] ^ n[26026];
assign t[26027] = t[26026] ^ n[26027];
assign t[26028] = t[26027] ^ n[26028];
assign t[26029] = t[26028] ^ n[26029];
assign t[26030] = t[26029] ^ n[26030];
assign t[26031] = t[26030] ^ n[26031];
assign t[26032] = t[26031] ^ n[26032];
assign t[26033] = t[26032] ^ n[26033];
assign t[26034] = t[26033] ^ n[26034];
assign t[26035] = t[26034] ^ n[26035];
assign t[26036] = t[26035] ^ n[26036];
assign t[26037] = t[26036] ^ n[26037];
assign t[26038] = t[26037] ^ n[26038];
assign t[26039] = t[26038] ^ n[26039];
assign t[26040] = t[26039] ^ n[26040];
assign t[26041] = t[26040] ^ n[26041];
assign t[26042] = t[26041] ^ n[26042];
assign t[26043] = t[26042] ^ n[26043];
assign t[26044] = t[26043] ^ n[26044];
assign t[26045] = t[26044] ^ n[26045];
assign t[26046] = t[26045] ^ n[26046];
assign t[26047] = t[26046] ^ n[26047];
assign t[26048] = t[26047] ^ n[26048];
assign t[26049] = t[26048] ^ n[26049];
assign t[26050] = t[26049] ^ n[26050];
assign t[26051] = t[26050] ^ n[26051];
assign t[26052] = t[26051] ^ n[26052];
assign t[26053] = t[26052] ^ n[26053];
assign t[26054] = t[26053] ^ n[26054];
assign t[26055] = t[26054] ^ n[26055];
assign t[26056] = t[26055] ^ n[26056];
assign t[26057] = t[26056] ^ n[26057];
assign t[26058] = t[26057] ^ n[26058];
assign t[26059] = t[26058] ^ n[26059];
assign t[26060] = t[26059] ^ n[26060];
assign t[26061] = t[26060] ^ n[26061];
assign t[26062] = t[26061] ^ n[26062];
assign t[26063] = t[26062] ^ n[26063];
assign t[26064] = t[26063] ^ n[26064];
assign t[26065] = t[26064] ^ n[26065];
assign t[26066] = t[26065] ^ n[26066];
assign t[26067] = t[26066] ^ n[26067];
assign t[26068] = t[26067] ^ n[26068];
assign t[26069] = t[26068] ^ n[26069];
assign t[26070] = t[26069] ^ n[26070];
assign t[26071] = t[26070] ^ n[26071];
assign t[26072] = t[26071] ^ n[26072];
assign t[26073] = t[26072] ^ n[26073];
assign t[26074] = t[26073] ^ n[26074];
assign t[26075] = t[26074] ^ n[26075];
assign t[26076] = t[26075] ^ n[26076];
assign t[26077] = t[26076] ^ n[26077];
assign t[26078] = t[26077] ^ n[26078];
assign t[26079] = t[26078] ^ n[26079];
assign t[26080] = t[26079] ^ n[26080];
assign t[26081] = t[26080] ^ n[26081];
assign t[26082] = t[26081] ^ n[26082];
assign t[26083] = t[26082] ^ n[26083];
assign t[26084] = t[26083] ^ n[26084];
assign t[26085] = t[26084] ^ n[26085];
assign t[26086] = t[26085] ^ n[26086];
assign t[26087] = t[26086] ^ n[26087];
assign t[26088] = t[26087] ^ n[26088];
assign t[26089] = t[26088] ^ n[26089];
assign t[26090] = t[26089] ^ n[26090];
assign t[26091] = t[26090] ^ n[26091];
assign t[26092] = t[26091] ^ n[26092];
assign t[26093] = t[26092] ^ n[26093];
assign t[26094] = t[26093] ^ n[26094];
assign t[26095] = t[26094] ^ n[26095];
assign t[26096] = t[26095] ^ n[26096];
assign t[26097] = t[26096] ^ n[26097];
assign t[26098] = t[26097] ^ n[26098];
assign t[26099] = t[26098] ^ n[26099];
assign t[26100] = t[26099] ^ n[26100];
assign t[26101] = t[26100] ^ n[26101];
assign t[26102] = t[26101] ^ n[26102];
assign t[26103] = t[26102] ^ n[26103];
assign t[26104] = t[26103] ^ n[26104];
assign t[26105] = t[26104] ^ n[26105];
assign t[26106] = t[26105] ^ n[26106];
assign t[26107] = t[26106] ^ n[26107];
assign t[26108] = t[26107] ^ n[26108];
assign t[26109] = t[26108] ^ n[26109];
assign t[26110] = t[26109] ^ n[26110];
assign t[26111] = t[26110] ^ n[26111];
assign t[26112] = t[26111] ^ n[26112];
assign t[26113] = t[26112] ^ n[26113];
assign t[26114] = t[26113] ^ n[26114];
assign t[26115] = t[26114] ^ n[26115];
assign t[26116] = t[26115] ^ n[26116];
assign t[26117] = t[26116] ^ n[26117];
assign t[26118] = t[26117] ^ n[26118];
assign t[26119] = t[26118] ^ n[26119];
assign t[26120] = t[26119] ^ n[26120];
assign t[26121] = t[26120] ^ n[26121];
assign t[26122] = t[26121] ^ n[26122];
assign t[26123] = t[26122] ^ n[26123];
assign t[26124] = t[26123] ^ n[26124];
assign t[26125] = t[26124] ^ n[26125];
assign t[26126] = t[26125] ^ n[26126];
assign t[26127] = t[26126] ^ n[26127];
assign t[26128] = t[26127] ^ n[26128];
assign t[26129] = t[26128] ^ n[26129];
assign t[26130] = t[26129] ^ n[26130];
assign t[26131] = t[26130] ^ n[26131];
assign t[26132] = t[26131] ^ n[26132];
assign t[26133] = t[26132] ^ n[26133];
assign t[26134] = t[26133] ^ n[26134];
assign t[26135] = t[26134] ^ n[26135];
assign t[26136] = t[26135] ^ n[26136];
assign t[26137] = t[26136] ^ n[26137];
assign t[26138] = t[26137] ^ n[26138];
assign t[26139] = t[26138] ^ n[26139];
assign t[26140] = t[26139] ^ n[26140];
assign t[26141] = t[26140] ^ n[26141];
assign t[26142] = t[26141] ^ n[26142];
assign t[26143] = t[26142] ^ n[26143];
assign t[26144] = t[26143] ^ n[26144];
assign t[26145] = t[26144] ^ n[26145];
assign t[26146] = t[26145] ^ n[26146];
assign t[26147] = t[26146] ^ n[26147];
assign t[26148] = t[26147] ^ n[26148];
assign t[26149] = t[26148] ^ n[26149];
assign t[26150] = t[26149] ^ n[26150];
assign t[26151] = t[26150] ^ n[26151];
assign t[26152] = t[26151] ^ n[26152];
assign t[26153] = t[26152] ^ n[26153];
assign t[26154] = t[26153] ^ n[26154];
assign t[26155] = t[26154] ^ n[26155];
assign t[26156] = t[26155] ^ n[26156];
assign t[26157] = t[26156] ^ n[26157];
assign t[26158] = t[26157] ^ n[26158];
assign t[26159] = t[26158] ^ n[26159];
assign t[26160] = t[26159] ^ n[26160];
assign t[26161] = t[26160] ^ n[26161];
assign t[26162] = t[26161] ^ n[26162];
assign t[26163] = t[26162] ^ n[26163];
assign t[26164] = t[26163] ^ n[26164];
assign t[26165] = t[26164] ^ n[26165];
assign t[26166] = t[26165] ^ n[26166];
assign t[26167] = t[26166] ^ n[26167];
assign t[26168] = t[26167] ^ n[26168];
assign t[26169] = t[26168] ^ n[26169];
assign t[26170] = t[26169] ^ n[26170];
assign t[26171] = t[26170] ^ n[26171];
assign t[26172] = t[26171] ^ n[26172];
assign t[26173] = t[26172] ^ n[26173];
assign t[26174] = t[26173] ^ n[26174];
assign t[26175] = t[26174] ^ n[26175];
assign t[26176] = t[26175] ^ n[26176];
assign t[26177] = t[26176] ^ n[26177];
assign t[26178] = t[26177] ^ n[26178];
assign t[26179] = t[26178] ^ n[26179];
assign t[26180] = t[26179] ^ n[26180];
assign t[26181] = t[26180] ^ n[26181];
assign t[26182] = t[26181] ^ n[26182];
assign t[26183] = t[26182] ^ n[26183];
assign t[26184] = t[26183] ^ n[26184];
assign t[26185] = t[26184] ^ n[26185];
assign t[26186] = t[26185] ^ n[26186];
assign t[26187] = t[26186] ^ n[26187];
assign t[26188] = t[26187] ^ n[26188];
assign t[26189] = t[26188] ^ n[26189];
assign t[26190] = t[26189] ^ n[26190];
assign t[26191] = t[26190] ^ n[26191];
assign t[26192] = t[26191] ^ n[26192];
assign t[26193] = t[26192] ^ n[26193];
assign t[26194] = t[26193] ^ n[26194];
assign t[26195] = t[26194] ^ n[26195];
assign t[26196] = t[26195] ^ n[26196];
assign t[26197] = t[26196] ^ n[26197];
assign t[26198] = t[26197] ^ n[26198];
assign t[26199] = t[26198] ^ n[26199];
assign t[26200] = t[26199] ^ n[26200];
assign t[26201] = t[26200] ^ n[26201];
assign t[26202] = t[26201] ^ n[26202];
assign t[26203] = t[26202] ^ n[26203];
assign t[26204] = t[26203] ^ n[26204];
assign t[26205] = t[26204] ^ n[26205];
assign t[26206] = t[26205] ^ n[26206];
assign t[26207] = t[26206] ^ n[26207];
assign t[26208] = t[26207] ^ n[26208];
assign t[26209] = t[26208] ^ n[26209];
assign t[26210] = t[26209] ^ n[26210];
assign t[26211] = t[26210] ^ n[26211];
assign t[26212] = t[26211] ^ n[26212];
assign t[26213] = t[26212] ^ n[26213];
assign t[26214] = t[26213] ^ n[26214];
assign t[26215] = t[26214] ^ n[26215];
assign t[26216] = t[26215] ^ n[26216];
assign t[26217] = t[26216] ^ n[26217];
assign t[26218] = t[26217] ^ n[26218];
assign t[26219] = t[26218] ^ n[26219];
assign t[26220] = t[26219] ^ n[26220];
assign t[26221] = t[26220] ^ n[26221];
assign t[26222] = t[26221] ^ n[26222];
assign t[26223] = t[26222] ^ n[26223];
assign t[26224] = t[26223] ^ n[26224];
assign t[26225] = t[26224] ^ n[26225];
assign t[26226] = t[26225] ^ n[26226];
assign t[26227] = t[26226] ^ n[26227];
assign t[26228] = t[26227] ^ n[26228];
assign t[26229] = t[26228] ^ n[26229];
assign t[26230] = t[26229] ^ n[26230];
assign t[26231] = t[26230] ^ n[26231];
assign t[26232] = t[26231] ^ n[26232];
assign t[26233] = t[26232] ^ n[26233];
assign t[26234] = t[26233] ^ n[26234];
assign t[26235] = t[26234] ^ n[26235];
assign t[26236] = t[26235] ^ n[26236];
assign t[26237] = t[26236] ^ n[26237];
assign t[26238] = t[26237] ^ n[26238];
assign t[26239] = t[26238] ^ n[26239];
assign t[26240] = t[26239] ^ n[26240];
assign t[26241] = t[26240] ^ n[26241];
assign t[26242] = t[26241] ^ n[26242];
assign t[26243] = t[26242] ^ n[26243];
assign t[26244] = t[26243] ^ n[26244];
assign t[26245] = t[26244] ^ n[26245];
assign t[26246] = t[26245] ^ n[26246];
assign t[26247] = t[26246] ^ n[26247];
assign t[26248] = t[26247] ^ n[26248];
assign t[26249] = t[26248] ^ n[26249];
assign t[26250] = t[26249] ^ n[26250];
assign t[26251] = t[26250] ^ n[26251];
assign t[26252] = t[26251] ^ n[26252];
assign t[26253] = t[26252] ^ n[26253];
assign t[26254] = t[26253] ^ n[26254];
assign t[26255] = t[26254] ^ n[26255];
assign t[26256] = t[26255] ^ n[26256];
assign t[26257] = t[26256] ^ n[26257];
assign t[26258] = t[26257] ^ n[26258];
assign t[26259] = t[26258] ^ n[26259];
assign t[26260] = t[26259] ^ n[26260];
assign t[26261] = t[26260] ^ n[26261];
assign t[26262] = t[26261] ^ n[26262];
assign t[26263] = t[26262] ^ n[26263];
assign t[26264] = t[26263] ^ n[26264];
assign t[26265] = t[26264] ^ n[26265];
assign t[26266] = t[26265] ^ n[26266];
assign t[26267] = t[26266] ^ n[26267];
assign t[26268] = t[26267] ^ n[26268];
assign t[26269] = t[26268] ^ n[26269];
assign t[26270] = t[26269] ^ n[26270];
assign t[26271] = t[26270] ^ n[26271];
assign t[26272] = t[26271] ^ n[26272];
assign t[26273] = t[26272] ^ n[26273];
assign t[26274] = t[26273] ^ n[26274];
assign t[26275] = t[26274] ^ n[26275];
assign t[26276] = t[26275] ^ n[26276];
assign t[26277] = t[26276] ^ n[26277];
assign t[26278] = t[26277] ^ n[26278];
assign t[26279] = t[26278] ^ n[26279];
assign t[26280] = t[26279] ^ n[26280];
assign t[26281] = t[26280] ^ n[26281];
assign t[26282] = t[26281] ^ n[26282];
assign t[26283] = t[26282] ^ n[26283];
assign t[26284] = t[26283] ^ n[26284];
assign t[26285] = t[26284] ^ n[26285];
assign t[26286] = t[26285] ^ n[26286];
assign t[26287] = t[26286] ^ n[26287];
assign t[26288] = t[26287] ^ n[26288];
assign t[26289] = t[26288] ^ n[26289];
assign t[26290] = t[26289] ^ n[26290];
assign t[26291] = t[26290] ^ n[26291];
assign t[26292] = t[26291] ^ n[26292];
assign t[26293] = t[26292] ^ n[26293];
assign t[26294] = t[26293] ^ n[26294];
assign t[26295] = t[26294] ^ n[26295];
assign t[26296] = t[26295] ^ n[26296];
assign t[26297] = t[26296] ^ n[26297];
assign t[26298] = t[26297] ^ n[26298];
assign t[26299] = t[26298] ^ n[26299];
assign t[26300] = t[26299] ^ n[26300];
assign t[26301] = t[26300] ^ n[26301];
assign t[26302] = t[26301] ^ n[26302];
assign t[26303] = t[26302] ^ n[26303];
assign t[26304] = t[26303] ^ n[26304];
assign t[26305] = t[26304] ^ n[26305];
assign t[26306] = t[26305] ^ n[26306];
assign t[26307] = t[26306] ^ n[26307];
assign t[26308] = t[26307] ^ n[26308];
assign t[26309] = t[26308] ^ n[26309];
assign t[26310] = t[26309] ^ n[26310];
assign t[26311] = t[26310] ^ n[26311];
assign t[26312] = t[26311] ^ n[26312];
assign t[26313] = t[26312] ^ n[26313];
assign t[26314] = t[26313] ^ n[26314];
assign t[26315] = t[26314] ^ n[26315];
assign t[26316] = t[26315] ^ n[26316];
assign t[26317] = t[26316] ^ n[26317];
assign t[26318] = t[26317] ^ n[26318];
assign t[26319] = t[26318] ^ n[26319];
assign t[26320] = t[26319] ^ n[26320];
assign t[26321] = t[26320] ^ n[26321];
assign t[26322] = t[26321] ^ n[26322];
assign t[26323] = t[26322] ^ n[26323];
assign t[26324] = t[26323] ^ n[26324];
assign t[26325] = t[26324] ^ n[26325];
assign t[26326] = t[26325] ^ n[26326];
assign t[26327] = t[26326] ^ n[26327];
assign t[26328] = t[26327] ^ n[26328];
assign t[26329] = t[26328] ^ n[26329];
assign t[26330] = t[26329] ^ n[26330];
assign t[26331] = t[26330] ^ n[26331];
assign t[26332] = t[26331] ^ n[26332];
assign t[26333] = t[26332] ^ n[26333];
assign t[26334] = t[26333] ^ n[26334];
assign t[26335] = t[26334] ^ n[26335];
assign t[26336] = t[26335] ^ n[26336];
assign t[26337] = t[26336] ^ n[26337];
assign t[26338] = t[26337] ^ n[26338];
assign t[26339] = t[26338] ^ n[26339];
assign t[26340] = t[26339] ^ n[26340];
assign t[26341] = t[26340] ^ n[26341];
assign t[26342] = t[26341] ^ n[26342];
assign t[26343] = t[26342] ^ n[26343];
assign t[26344] = t[26343] ^ n[26344];
assign t[26345] = t[26344] ^ n[26345];
assign t[26346] = t[26345] ^ n[26346];
assign t[26347] = t[26346] ^ n[26347];
assign t[26348] = t[26347] ^ n[26348];
assign t[26349] = t[26348] ^ n[26349];
assign t[26350] = t[26349] ^ n[26350];
assign t[26351] = t[26350] ^ n[26351];
assign t[26352] = t[26351] ^ n[26352];
assign t[26353] = t[26352] ^ n[26353];
assign t[26354] = t[26353] ^ n[26354];
assign t[26355] = t[26354] ^ n[26355];
assign t[26356] = t[26355] ^ n[26356];
assign t[26357] = t[26356] ^ n[26357];
assign t[26358] = t[26357] ^ n[26358];
assign t[26359] = t[26358] ^ n[26359];
assign t[26360] = t[26359] ^ n[26360];
assign t[26361] = t[26360] ^ n[26361];
assign t[26362] = t[26361] ^ n[26362];
assign t[26363] = t[26362] ^ n[26363];
assign t[26364] = t[26363] ^ n[26364];
assign t[26365] = t[26364] ^ n[26365];
assign t[26366] = t[26365] ^ n[26366];
assign t[26367] = t[26366] ^ n[26367];
assign t[26368] = t[26367] ^ n[26368];
assign t[26369] = t[26368] ^ n[26369];
assign t[26370] = t[26369] ^ n[26370];
assign t[26371] = t[26370] ^ n[26371];
assign t[26372] = t[26371] ^ n[26372];
assign t[26373] = t[26372] ^ n[26373];
assign t[26374] = t[26373] ^ n[26374];
assign t[26375] = t[26374] ^ n[26375];
assign t[26376] = t[26375] ^ n[26376];
assign t[26377] = t[26376] ^ n[26377];
assign t[26378] = t[26377] ^ n[26378];
assign t[26379] = t[26378] ^ n[26379];
assign t[26380] = t[26379] ^ n[26380];
assign t[26381] = t[26380] ^ n[26381];
assign t[26382] = t[26381] ^ n[26382];
assign t[26383] = t[26382] ^ n[26383];
assign t[26384] = t[26383] ^ n[26384];
assign t[26385] = t[26384] ^ n[26385];
assign t[26386] = t[26385] ^ n[26386];
assign t[26387] = t[26386] ^ n[26387];
assign t[26388] = t[26387] ^ n[26388];
assign t[26389] = t[26388] ^ n[26389];
assign t[26390] = t[26389] ^ n[26390];
assign t[26391] = t[26390] ^ n[26391];
assign t[26392] = t[26391] ^ n[26392];
assign t[26393] = t[26392] ^ n[26393];
assign t[26394] = t[26393] ^ n[26394];
assign t[26395] = t[26394] ^ n[26395];
assign t[26396] = t[26395] ^ n[26396];
assign t[26397] = t[26396] ^ n[26397];
assign t[26398] = t[26397] ^ n[26398];
assign t[26399] = t[26398] ^ n[26399];
assign t[26400] = t[26399] ^ n[26400];
assign t[26401] = t[26400] ^ n[26401];
assign t[26402] = t[26401] ^ n[26402];
assign t[26403] = t[26402] ^ n[26403];
assign t[26404] = t[26403] ^ n[26404];
assign t[26405] = t[26404] ^ n[26405];
assign t[26406] = t[26405] ^ n[26406];
assign t[26407] = t[26406] ^ n[26407];
assign t[26408] = t[26407] ^ n[26408];
assign t[26409] = t[26408] ^ n[26409];
assign t[26410] = t[26409] ^ n[26410];
assign t[26411] = t[26410] ^ n[26411];
assign t[26412] = t[26411] ^ n[26412];
assign t[26413] = t[26412] ^ n[26413];
assign t[26414] = t[26413] ^ n[26414];
assign t[26415] = t[26414] ^ n[26415];
assign t[26416] = t[26415] ^ n[26416];
assign t[26417] = t[26416] ^ n[26417];
assign t[26418] = t[26417] ^ n[26418];
assign t[26419] = t[26418] ^ n[26419];
assign t[26420] = t[26419] ^ n[26420];
assign t[26421] = t[26420] ^ n[26421];
assign t[26422] = t[26421] ^ n[26422];
assign t[26423] = t[26422] ^ n[26423];
assign t[26424] = t[26423] ^ n[26424];
assign t[26425] = t[26424] ^ n[26425];
assign t[26426] = t[26425] ^ n[26426];
assign t[26427] = t[26426] ^ n[26427];
assign t[26428] = t[26427] ^ n[26428];
assign t[26429] = t[26428] ^ n[26429];
assign t[26430] = t[26429] ^ n[26430];
assign t[26431] = t[26430] ^ n[26431];
assign t[26432] = t[26431] ^ n[26432];
assign t[26433] = t[26432] ^ n[26433];
assign t[26434] = t[26433] ^ n[26434];
assign t[26435] = t[26434] ^ n[26435];
assign t[26436] = t[26435] ^ n[26436];
assign t[26437] = t[26436] ^ n[26437];
assign t[26438] = t[26437] ^ n[26438];
assign t[26439] = t[26438] ^ n[26439];
assign t[26440] = t[26439] ^ n[26440];
assign t[26441] = t[26440] ^ n[26441];
assign t[26442] = t[26441] ^ n[26442];
assign t[26443] = t[26442] ^ n[26443];
assign t[26444] = t[26443] ^ n[26444];
assign t[26445] = t[26444] ^ n[26445];
assign t[26446] = t[26445] ^ n[26446];
assign t[26447] = t[26446] ^ n[26447];
assign t[26448] = t[26447] ^ n[26448];
assign t[26449] = t[26448] ^ n[26449];
assign t[26450] = t[26449] ^ n[26450];
assign t[26451] = t[26450] ^ n[26451];
assign t[26452] = t[26451] ^ n[26452];
assign t[26453] = t[26452] ^ n[26453];
assign t[26454] = t[26453] ^ n[26454];
assign t[26455] = t[26454] ^ n[26455];
assign t[26456] = t[26455] ^ n[26456];
assign t[26457] = t[26456] ^ n[26457];
assign t[26458] = t[26457] ^ n[26458];
assign t[26459] = t[26458] ^ n[26459];
assign t[26460] = t[26459] ^ n[26460];
assign t[26461] = t[26460] ^ n[26461];
assign t[26462] = t[26461] ^ n[26462];
assign t[26463] = t[26462] ^ n[26463];
assign t[26464] = t[26463] ^ n[26464];
assign t[26465] = t[26464] ^ n[26465];
assign t[26466] = t[26465] ^ n[26466];
assign t[26467] = t[26466] ^ n[26467];
assign t[26468] = t[26467] ^ n[26468];
assign t[26469] = t[26468] ^ n[26469];
assign t[26470] = t[26469] ^ n[26470];
assign t[26471] = t[26470] ^ n[26471];
assign t[26472] = t[26471] ^ n[26472];
assign t[26473] = t[26472] ^ n[26473];
assign t[26474] = t[26473] ^ n[26474];
assign t[26475] = t[26474] ^ n[26475];
assign t[26476] = t[26475] ^ n[26476];
assign t[26477] = t[26476] ^ n[26477];
assign t[26478] = t[26477] ^ n[26478];
assign t[26479] = t[26478] ^ n[26479];
assign t[26480] = t[26479] ^ n[26480];
assign t[26481] = t[26480] ^ n[26481];
assign t[26482] = t[26481] ^ n[26482];
assign t[26483] = t[26482] ^ n[26483];
assign t[26484] = t[26483] ^ n[26484];
assign t[26485] = t[26484] ^ n[26485];
assign t[26486] = t[26485] ^ n[26486];
assign t[26487] = t[26486] ^ n[26487];
assign t[26488] = t[26487] ^ n[26488];
assign t[26489] = t[26488] ^ n[26489];
assign t[26490] = t[26489] ^ n[26490];
assign t[26491] = t[26490] ^ n[26491];
assign t[26492] = t[26491] ^ n[26492];
assign t[26493] = t[26492] ^ n[26493];
assign t[26494] = t[26493] ^ n[26494];
assign t[26495] = t[26494] ^ n[26495];
assign t[26496] = t[26495] ^ n[26496];
assign t[26497] = t[26496] ^ n[26497];
assign t[26498] = t[26497] ^ n[26498];
assign t[26499] = t[26498] ^ n[26499];
assign t[26500] = t[26499] ^ n[26500];
assign t[26501] = t[26500] ^ n[26501];
assign t[26502] = t[26501] ^ n[26502];
assign t[26503] = t[26502] ^ n[26503];
assign t[26504] = t[26503] ^ n[26504];
assign t[26505] = t[26504] ^ n[26505];
assign t[26506] = t[26505] ^ n[26506];
assign t[26507] = t[26506] ^ n[26507];
assign t[26508] = t[26507] ^ n[26508];
assign t[26509] = t[26508] ^ n[26509];
assign t[26510] = t[26509] ^ n[26510];
assign t[26511] = t[26510] ^ n[26511];
assign t[26512] = t[26511] ^ n[26512];
assign t[26513] = t[26512] ^ n[26513];
assign t[26514] = t[26513] ^ n[26514];
assign t[26515] = t[26514] ^ n[26515];
assign t[26516] = t[26515] ^ n[26516];
assign t[26517] = t[26516] ^ n[26517];
assign t[26518] = t[26517] ^ n[26518];
assign t[26519] = t[26518] ^ n[26519];
assign t[26520] = t[26519] ^ n[26520];
assign t[26521] = t[26520] ^ n[26521];
assign t[26522] = t[26521] ^ n[26522];
assign t[26523] = t[26522] ^ n[26523];
assign t[26524] = t[26523] ^ n[26524];
assign t[26525] = t[26524] ^ n[26525];
assign t[26526] = t[26525] ^ n[26526];
assign t[26527] = t[26526] ^ n[26527];
assign t[26528] = t[26527] ^ n[26528];
assign t[26529] = t[26528] ^ n[26529];
assign t[26530] = t[26529] ^ n[26530];
assign t[26531] = t[26530] ^ n[26531];
assign t[26532] = t[26531] ^ n[26532];
assign t[26533] = t[26532] ^ n[26533];
assign t[26534] = t[26533] ^ n[26534];
assign t[26535] = t[26534] ^ n[26535];
assign t[26536] = t[26535] ^ n[26536];
assign t[26537] = t[26536] ^ n[26537];
assign t[26538] = t[26537] ^ n[26538];
assign t[26539] = t[26538] ^ n[26539];
assign t[26540] = t[26539] ^ n[26540];
assign t[26541] = t[26540] ^ n[26541];
assign t[26542] = t[26541] ^ n[26542];
assign t[26543] = t[26542] ^ n[26543];
assign t[26544] = t[26543] ^ n[26544];
assign t[26545] = t[26544] ^ n[26545];
assign t[26546] = t[26545] ^ n[26546];
assign t[26547] = t[26546] ^ n[26547];
assign t[26548] = t[26547] ^ n[26548];
assign t[26549] = t[26548] ^ n[26549];
assign t[26550] = t[26549] ^ n[26550];
assign t[26551] = t[26550] ^ n[26551];
assign t[26552] = t[26551] ^ n[26552];
assign t[26553] = t[26552] ^ n[26553];
assign t[26554] = t[26553] ^ n[26554];
assign t[26555] = t[26554] ^ n[26555];
assign t[26556] = t[26555] ^ n[26556];
assign t[26557] = t[26556] ^ n[26557];
assign t[26558] = t[26557] ^ n[26558];
assign t[26559] = t[26558] ^ n[26559];
assign t[26560] = t[26559] ^ n[26560];
assign t[26561] = t[26560] ^ n[26561];
assign t[26562] = t[26561] ^ n[26562];
assign t[26563] = t[26562] ^ n[26563];
assign t[26564] = t[26563] ^ n[26564];
assign t[26565] = t[26564] ^ n[26565];
assign t[26566] = t[26565] ^ n[26566];
assign t[26567] = t[26566] ^ n[26567];
assign t[26568] = t[26567] ^ n[26568];
assign t[26569] = t[26568] ^ n[26569];
assign t[26570] = t[26569] ^ n[26570];
assign t[26571] = t[26570] ^ n[26571];
assign t[26572] = t[26571] ^ n[26572];
assign t[26573] = t[26572] ^ n[26573];
assign t[26574] = t[26573] ^ n[26574];
assign t[26575] = t[26574] ^ n[26575];
assign t[26576] = t[26575] ^ n[26576];
assign t[26577] = t[26576] ^ n[26577];
assign t[26578] = t[26577] ^ n[26578];
assign t[26579] = t[26578] ^ n[26579];
assign t[26580] = t[26579] ^ n[26580];
assign t[26581] = t[26580] ^ n[26581];
assign t[26582] = t[26581] ^ n[26582];
assign t[26583] = t[26582] ^ n[26583];
assign t[26584] = t[26583] ^ n[26584];
assign t[26585] = t[26584] ^ n[26585];
assign t[26586] = t[26585] ^ n[26586];
assign t[26587] = t[26586] ^ n[26587];
assign t[26588] = t[26587] ^ n[26588];
assign t[26589] = t[26588] ^ n[26589];
assign t[26590] = t[26589] ^ n[26590];
assign t[26591] = t[26590] ^ n[26591];
assign t[26592] = t[26591] ^ n[26592];
assign t[26593] = t[26592] ^ n[26593];
assign t[26594] = t[26593] ^ n[26594];
assign t[26595] = t[26594] ^ n[26595];
assign t[26596] = t[26595] ^ n[26596];
assign t[26597] = t[26596] ^ n[26597];
assign t[26598] = t[26597] ^ n[26598];
assign t[26599] = t[26598] ^ n[26599];
assign t[26600] = t[26599] ^ n[26600];
assign t[26601] = t[26600] ^ n[26601];
assign t[26602] = t[26601] ^ n[26602];
assign t[26603] = t[26602] ^ n[26603];
assign t[26604] = t[26603] ^ n[26604];
assign t[26605] = t[26604] ^ n[26605];
assign t[26606] = t[26605] ^ n[26606];
assign t[26607] = t[26606] ^ n[26607];
assign t[26608] = t[26607] ^ n[26608];
assign t[26609] = t[26608] ^ n[26609];
assign t[26610] = t[26609] ^ n[26610];
assign t[26611] = t[26610] ^ n[26611];
assign t[26612] = t[26611] ^ n[26612];
assign t[26613] = t[26612] ^ n[26613];
assign t[26614] = t[26613] ^ n[26614];
assign t[26615] = t[26614] ^ n[26615];
assign t[26616] = t[26615] ^ n[26616];
assign t[26617] = t[26616] ^ n[26617];
assign t[26618] = t[26617] ^ n[26618];
assign t[26619] = t[26618] ^ n[26619];
assign t[26620] = t[26619] ^ n[26620];
assign t[26621] = t[26620] ^ n[26621];
assign t[26622] = t[26621] ^ n[26622];
assign t[26623] = t[26622] ^ n[26623];
assign t[26624] = t[26623] ^ n[26624];
assign t[26625] = t[26624] ^ n[26625];
assign t[26626] = t[26625] ^ n[26626];
assign t[26627] = t[26626] ^ n[26627];
assign t[26628] = t[26627] ^ n[26628];
assign t[26629] = t[26628] ^ n[26629];
assign t[26630] = t[26629] ^ n[26630];
assign t[26631] = t[26630] ^ n[26631];
assign t[26632] = t[26631] ^ n[26632];
assign t[26633] = t[26632] ^ n[26633];
assign t[26634] = t[26633] ^ n[26634];
assign t[26635] = t[26634] ^ n[26635];
assign t[26636] = t[26635] ^ n[26636];
assign t[26637] = t[26636] ^ n[26637];
assign t[26638] = t[26637] ^ n[26638];
assign t[26639] = t[26638] ^ n[26639];
assign t[26640] = t[26639] ^ n[26640];
assign t[26641] = t[26640] ^ n[26641];
assign t[26642] = t[26641] ^ n[26642];
assign t[26643] = t[26642] ^ n[26643];
assign t[26644] = t[26643] ^ n[26644];
assign t[26645] = t[26644] ^ n[26645];
assign t[26646] = t[26645] ^ n[26646];
assign t[26647] = t[26646] ^ n[26647];
assign t[26648] = t[26647] ^ n[26648];
assign t[26649] = t[26648] ^ n[26649];
assign t[26650] = t[26649] ^ n[26650];
assign t[26651] = t[26650] ^ n[26651];
assign t[26652] = t[26651] ^ n[26652];
assign t[26653] = t[26652] ^ n[26653];
assign t[26654] = t[26653] ^ n[26654];
assign t[26655] = t[26654] ^ n[26655];
assign t[26656] = t[26655] ^ n[26656];
assign t[26657] = t[26656] ^ n[26657];
assign t[26658] = t[26657] ^ n[26658];
assign t[26659] = t[26658] ^ n[26659];
assign t[26660] = t[26659] ^ n[26660];
assign t[26661] = t[26660] ^ n[26661];
assign t[26662] = t[26661] ^ n[26662];
assign t[26663] = t[26662] ^ n[26663];
assign t[26664] = t[26663] ^ n[26664];
assign t[26665] = t[26664] ^ n[26665];
assign t[26666] = t[26665] ^ n[26666];
assign t[26667] = t[26666] ^ n[26667];
assign t[26668] = t[26667] ^ n[26668];
assign t[26669] = t[26668] ^ n[26669];
assign t[26670] = t[26669] ^ n[26670];
assign t[26671] = t[26670] ^ n[26671];
assign t[26672] = t[26671] ^ n[26672];
assign t[26673] = t[26672] ^ n[26673];
assign t[26674] = t[26673] ^ n[26674];
assign t[26675] = t[26674] ^ n[26675];
assign t[26676] = t[26675] ^ n[26676];
assign t[26677] = t[26676] ^ n[26677];
assign t[26678] = t[26677] ^ n[26678];
assign t[26679] = t[26678] ^ n[26679];
assign t[26680] = t[26679] ^ n[26680];
assign t[26681] = t[26680] ^ n[26681];
assign t[26682] = t[26681] ^ n[26682];
assign t[26683] = t[26682] ^ n[26683];
assign t[26684] = t[26683] ^ n[26684];
assign t[26685] = t[26684] ^ n[26685];
assign t[26686] = t[26685] ^ n[26686];
assign t[26687] = t[26686] ^ n[26687];
assign t[26688] = t[26687] ^ n[26688];
assign t[26689] = t[26688] ^ n[26689];
assign t[26690] = t[26689] ^ n[26690];
assign t[26691] = t[26690] ^ n[26691];
assign t[26692] = t[26691] ^ n[26692];
assign t[26693] = t[26692] ^ n[26693];
assign t[26694] = t[26693] ^ n[26694];
assign t[26695] = t[26694] ^ n[26695];
assign t[26696] = t[26695] ^ n[26696];
assign t[26697] = t[26696] ^ n[26697];
assign t[26698] = t[26697] ^ n[26698];
assign t[26699] = t[26698] ^ n[26699];
assign t[26700] = t[26699] ^ n[26700];
assign t[26701] = t[26700] ^ n[26701];
assign t[26702] = t[26701] ^ n[26702];
assign t[26703] = t[26702] ^ n[26703];
assign t[26704] = t[26703] ^ n[26704];
assign t[26705] = t[26704] ^ n[26705];
assign t[26706] = t[26705] ^ n[26706];
assign t[26707] = t[26706] ^ n[26707];
assign t[26708] = t[26707] ^ n[26708];
assign t[26709] = t[26708] ^ n[26709];
assign t[26710] = t[26709] ^ n[26710];
assign t[26711] = t[26710] ^ n[26711];
assign t[26712] = t[26711] ^ n[26712];
assign t[26713] = t[26712] ^ n[26713];
assign t[26714] = t[26713] ^ n[26714];
assign t[26715] = t[26714] ^ n[26715];
assign t[26716] = t[26715] ^ n[26716];
assign t[26717] = t[26716] ^ n[26717];
assign t[26718] = t[26717] ^ n[26718];
assign t[26719] = t[26718] ^ n[26719];
assign t[26720] = t[26719] ^ n[26720];
assign t[26721] = t[26720] ^ n[26721];
assign t[26722] = t[26721] ^ n[26722];
assign t[26723] = t[26722] ^ n[26723];
assign t[26724] = t[26723] ^ n[26724];
assign t[26725] = t[26724] ^ n[26725];
assign t[26726] = t[26725] ^ n[26726];
assign t[26727] = t[26726] ^ n[26727];
assign t[26728] = t[26727] ^ n[26728];
assign t[26729] = t[26728] ^ n[26729];
assign t[26730] = t[26729] ^ n[26730];
assign t[26731] = t[26730] ^ n[26731];
assign t[26732] = t[26731] ^ n[26732];
assign t[26733] = t[26732] ^ n[26733];
assign t[26734] = t[26733] ^ n[26734];
assign t[26735] = t[26734] ^ n[26735];
assign t[26736] = t[26735] ^ n[26736];
assign t[26737] = t[26736] ^ n[26737];
assign t[26738] = t[26737] ^ n[26738];
assign t[26739] = t[26738] ^ n[26739];
assign t[26740] = t[26739] ^ n[26740];
assign t[26741] = t[26740] ^ n[26741];
assign t[26742] = t[26741] ^ n[26742];
assign t[26743] = t[26742] ^ n[26743];
assign t[26744] = t[26743] ^ n[26744];
assign t[26745] = t[26744] ^ n[26745];
assign t[26746] = t[26745] ^ n[26746];
assign t[26747] = t[26746] ^ n[26747];
assign t[26748] = t[26747] ^ n[26748];
assign t[26749] = t[26748] ^ n[26749];
assign t[26750] = t[26749] ^ n[26750];
assign t[26751] = t[26750] ^ n[26751];
assign t[26752] = t[26751] ^ n[26752];
assign t[26753] = t[26752] ^ n[26753];
assign t[26754] = t[26753] ^ n[26754];
assign t[26755] = t[26754] ^ n[26755];
assign t[26756] = t[26755] ^ n[26756];
assign t[26757] = t[26756] ^ n[26757];
assign t[26758] = t[26757] ^ n[26758];
assign t[26759] = t[26758] ^ n[26759];
assign t[26760] = t[26759] ^ n[26760];
assign t[26761] = t[26760] ^ n[26761];
assign t[26762] = t[26761] ^ n[26762];
assign t[26763] = t[26762] ^ n[26763];
assign t[26764] = t[26763] ^ n[26764];
assign t[26765] = t[26764] ^ n[26765];
assign t[26766] = t[26765] ^ n[26766];
assign t[26767] = t[26766] ^ n[26767];
assign t[26768] = t[26767] ^ n[26768];
assign t[26769] = t[26768] ^ n[26769];
assign t[26770] = t[26769] ^ n[26770];
assign t[26771] = t[26770] ^ n[26771];
assign t[26772] = t[26771] ^ n[26772];
assign t[26773] = t[26772] ^ n[26773];
assign t[26774] = t[26773] ^ n[26774];
assign t[26775] = t[26774] ^ n[26775];
assign t[26776] = t[26775] ^ n[26776];
assign t[26777] = t[26776] ^ n[26777];
assign t[26778] = t[26777] ^ n[26778];
assign t[26779] = t[26778] ^ n[26779];
assign t[26780] = t[26779] ^ n[26780];
assign t[26781] = t[26780] ^ n[26781];
assign t[26782] = t[26781] ^ n[26782];
assign t[26783] = t[26782] ^ n[26783];
assign t[26784] = t[26783] ^ n[26784];
assign t[26785] = t[26784] ^ n[26785];
assign t[26786] = t[26785] ^ n[26786];
assign t[26787] = t[26786] ^ n[26787];
assign t[26788] = t[26787] ^ n[26788];
assign t[26789] = t[26788] ^ n[26789];
assign t[26790] = t[26789] ^ n[26790];
assign t[26791] = t[26790] ^ n[26791];
assign t[26792] = t[26791] ^ n[26792];
assign t[26793] = t[26792] ^ n[26793];
assign t[26794] = t[26793] ^ n[26794];
assign t[26795] = t[26794] ^ n[26795];
assign t[26796] = t[26795] ^ n[26796];
assign t[26797] = t[26796] ^ n[26797];
assign t[26798] = t[26797] ^ n[26798];
assign t[26799] = t[26798] ^ n[26799];
assign t[26800] = t[26799] ^ n[26800];
assign t[26801] = t[26800] ^ n[26801];
assign t[26802] = t[26801] ^ n[26802];
assign t[26803] = t[26802] ^ n[26803];
assign t[26804] = t[26803] ^ n[26804];
assign t[26805] = t[26804] ^ n[26805];
assign t[26806] = t[26805] ^ n[26806];
assign t[26807] = t[26806] ^ n[26807];
assign t[26808] = t[26807] ^ n[26808];
assign t[26809] = t[26808] ^ n[26809];
assign t[26810] = t[26809] ^ n[26810];
assign t[26811] = t[26810] ^ n[26811];
assign t[26812] = t[26811] ^ n[26812];
assign t[26813] = t[26812] ^ n[26813];
assign t[26814] = t[26813] ^ n[26814];
assign t[26815] = t[26814] ^ n[26815];
assign t[26816] = t[26815] ^ n[26816];
assign t[26817] = t[26816] ^ n[26817];
assign t[26818] = t[26817] ^ n[26818];
assign t[26819] = t[26818] ^ n[26819];
assign t[26820] = t[26819] ^ n[26820];
assign t[26821] = t[26820] ^ n[26821];
assign t[26822] = t[26821] ^ n[26822];
assign t[26823] = t[26822] ^ n[26823];
assign t[26824] = t[26823] ^ n[26824];
assign t[26825] = t[26824] ^ n[26825];
assign t[26826] = t[26825] ^ n[26826];
assign t[26827] = t[26826] ^ n[26827];
assign t[26828] = t[26827] ^ n[26828];
assign t[26829] = t[26828] ^ n[26829];
assign t[26830] = t[26829] ^ n[26830];
assign t[26831] = t[26830] ^ n[26831];
assign t[26832] = t[26831] ^ n[26832];
assign t[26833] = t[26832] ^ n[26833];
assign t[26834] = t[26833] ^ n[26834];
assign t[26835] = t[26834] ^ n[26835];
assign t[26836] = t[26835] ^ n[26836];
assign t[26837] = t[26836] ^ n[26837];
assign t[26838] = t[26837] ^ n[26838];
assign t[26839] = t[26838] ^ n[26839];
assign t[26840] = t[26839] ^ n[26840];
assign t[26841] = t[26840] ^ n[26841];
assign t[26842] = t[26841] ^ n[26842];
assign t[26843] = t[26842] ^ n[26843];
assign t[26844] = t[26843] ^ n[26844];
assign t[26845] = t[26844] ^ n[26845];
assign t[26846] = t[26845] ^ n[26846];
assign t[26847] = t[26846] ^ n[26847];
assign t[26848] = t[26847] ^ n[26848];
assign t[26849] = t[26848] ^ n[26849];
assign t[26850] = t[26849] ^ n[26850];
assign t[26851] = t[26850] ^ n[26851];
assign t[26852] = t[26851] ^ n[26852];
assign t[26853] = t[26852] ^ n[26853];
assign t[26854] = t[26853] ^ n[26854];
assign t[26855] = t[26854] ^ n[26855];
assign t[26856] = t[26855] ^ n[26856];
assign t[26857] = t[26856] ^ n[26857];
assign t[26858] = t[26857] ^ n[26858];
assign t[26859] = t[26858] ^ n[26859];
assign t[26860] = t[26859] ^ n[26860];
assign t[26861] = t[26860] ^ n[26861];
assign t[26862] = t[26861] ^ n[26862];
assign t[26863] = t[26862] ^ n[26863];
assign t[26864] = t[26863] ^ n[26864];
assign t[26865] = t[26864] ^ n[26865];
assign t[26866] = t[26865] ^ n[26866];
assign t[26867] = t[26866] ^ n[26867];
assign t[26868] = t[26867] ^ n[26868];
assign t[26869] = t[26868] ^ n[26869];
assign t[26870] = t[26869] ^ n[26870];
assign t[26871] = t[26870] ^ n[26871];
assign t[26872] = t[26871] ^ n[26872];
assign t[26873] = t[26872] ^ n[26873];
assign t[26874] = t[26873] ^ n[26874];
assign t[26875] = t[26874] ^ n[26875];
assign t[26876] = t[26875] ^ n[26876];
assign t[26877] = t[26876] ^ n[26877];
assign t[26878] = t[26877] ^ n[26878];
assign t[26879] = t[26878] ^ n[26879];
assign t[26880] = t[26879] ^ n[26880];
assign t[26881] = t[26880] ^ n[26881];
assign t[26882] = t[26881] ^ n[26882];
assign t[26883] = t[26882] ^ n[26883];
assign t[26884] = t[26883] ^ n[26884];
assign t[26885] = t[26884] ^ n[26885];
assign t[26886] = t[26885] ^ n[26886];
assign t[26887] = t[26886] ^ n[26887];
assign t[26888] = t[26887] ^ n[26888];
assign t[26889] = t[26888] ^ n[26889];
assign t[26890] = t[26889] ^ n[26890];
assign t[26891] = t[26890] ^ n[26891];
assign t[26892] = t[26891] ^ n[26892];
assign t[26893] = t[26892] ^ n[26893];
assign t[26894] = t[26893] ^ n[26894];
assign t[26895] = t[26894] ^ n[26895];
assign t[26896] = t[26895] ^ n[26896];
assign t[26897] = t[26896] ^ n[26897];
assign t[26898] = t[26897] ^ n[26898];
assign t[26899] = t[26898] ^ n[26899];
assign t[26900] = t[26899] ^ n[26900];
assign t[26901] = t[26900] ^ n[26901];
assign t[26902] = t[26901] ^ n[26902];
assign t[26903] = t[26902] ^ n[26903];
assign t[26904] = t[26903] ^ n[26904];
assign t[26905] = t[26904] ^ n[26905];
assign t[26906] = t[26905] ^ n[26906];
assign t[26907] = t[26906] ^ n[26907];
assign t[26908] = t[26907] ^ n[26908];
assign t[26909] = t[26908] ^ n[26909];
assign t[26910] = t[26909] ^ n[26910];
assign t[26911] = t[26910] ^ n[26911];
assign t[26912] = t[26911] ^ n[26912];
assign t[26913] = t[26912] ^ n[26913];
assign t[26914] = t[26913] ^ n[26914];
assign t[26915] = t[26914] ^ n[26915];
assign t[26916] = t[26915] ^ n[26916];
assign t[26917] = t[26916] ^ n[26917];
assign t[26918] = t[26917] ^ n[26918];
assign t[26919] = t[26918] ^ n[26919];
assign t[26920] = t[26919] ^ n[26920];
assign t[26921] = t[26920] ^ n[26921];
assign t[26922] = t[26921] ^ n[26922];
assign t[26923] = t[26922] ^ n[26923];
assign t[26924] = t[26923] ^ n[26924];
assign t[26925] = t[26924] ^ n[26925];
assign t[26926] = t[26925] ^ n[26926];
assign t[26927] = t[26926] ^ n[26927];
assign t[26928] = t[26927] ^ n[26928];
assign t[26929] = t[26928] ^ n[26929];
assign t[26930] = t[26929] ^ n[26930];
assign t[26931] = t[26930] ^ n[26931];
assign t[26932] = t[26931] ^ n[26932];
assign t[26933] = t[26932] ^ n[26933];
assign t[26934] = t[26933] ^ n[26934];
assign t[26935] = t[26934] ^ n[26935];
assign t[26936] = t[26935] ^ n[26936];
assign t[26937] = t[26936] ^ n[26937];
assign t[26938] = t[26937] ^ n[26938];
assign t[26939] = t[26938] ^ n[26939];
assign t[26940] = t[26939] ^ n[26940];
assign t[26941] = t[26940] ^ n[26941];
assign t[26942] = t[26941] ^ n[26942];
assign t[26943] = t[26942] ^ n[26943];
assign t[26944] = t[26943] ^ n[26944];
assign t[26945] = t[26944] ^ n[26945];
assign t[26946] = t[26945] ^ n[26946];
assign t[26947] = t[26946] ^ n[26947];
assign t[26948] = t[26947] ^ n[26948];
assign t[26949] = t[26948] ^ n[26949];
assign t[26950] = t[26949] ^ n[26950];
assign t[26951] = t[26950] ^ n[26951];
assign t[26952] = t[26951] ^ n[26952];
assign t[26953] = t[26952] ^ n[26953];
assign t[26954] = t[26953] ^ n[26954];
assign t[26955] = t[26954] ^ n[26955];
assign t[26956] = t[26955] ^ n[26956];
assign t[26957] = t[26956] ^ n[26957];
assign t[26958] = t[26957] ^ n[26958];
assign t[26959] = t[26958] ^ n[26959];
assign t[26960] = t[26959] ^ n[26960];
assign t[26961] = t[26960] ^ n[26961];
assign t[26962] = t[26961] ^ n[26962];
assign t[26963] = t[26962] ^ n[26963];
assign t[26964] = t[26963] ^ n[26964];
assign t[26965] = t[26964] ^ n[26965];
assign t[26966] = t[26965] ^ n[26966];
assign t[26967] = t[26966] ^ n[26967];
assign t[26968] = t[26967] ^ n[26968];
assign t[26969] = t[26968] ^ n[26969];
assign t[26970] = t[26969] ^ n[26970];
assign t[26971] = t[26970] ^ n[26971];
assign t[26972] = t[26971] ^ n[26972];
assign t[26973] = t[26972] ^ n[26973];
assign t[26974] = t[26973] ^ n[26974];
assign t[26975] = t[26974] ^ n[26975];
assign t[26976] = t[26975] ^ n[26976];
assign t[26977] = t[26976] ^ n[26977];
assign t[26978] = t[26977] ^ n[26978];
assign t[26979] = t[26978] ^ n[26979];
assign t[26980] = t[26979] ^ n[26980];
assign t[26981] = t[26980] ^ n[26981];
assign t[26982] = t[26981] ^ n[26982];
assign t[26983] = t[26982] ^ n[26983];
assign t[26984] = t[26983] ^ n[26984];
assign t[26985] = t[26984] ^ n[26985];
assign t[26986] = t[26985] ^ n[26986];
assign t[26987] = t[26986] ^ n[26987];
assign t[26988] = t[26987] ^ n[26988];
assign t[26989] = t[26988] ^ n[26989];
assign t[26990] = t[26989] ^ n[26990];
assign t[26991] = t[26990] ^ n[26991];
assign t[26992] = t[26991] ^ n[26992];
assign t[26993] = t[26992] ^ n[26993];
assign t[26994] = t[26993] ^ n[26994];
assign t[26995] = t[26994] ^ n[26995];
assign t[26996] = t[26995] ^ n[26996];
assign t[26997] = t[26996] ^ n[26997];
assign t[26998] = t[26997] ^ n[26998];
assign t[26999] = t[26998] ^ n[26999];
assign t[27000] = t[26999] ^ n[27000];
assign t[27001] = t[27000] ^ n[27001];
assign t[27002] = t[27001] ^ n[27002];
assign t[27003] = t[27002] ^ n[27003];
assign t[27004] = t[27003] ^ n[27004];
assign t[27005] = t[27004] ^ n[27005];
assign t[27006] = t[27005] ^ n[27006];
assign t[27007] = t[27006] ^ n[27007];
assign t[27008] = t[27007] ^ n[27008];
assign t[27009] = t[27008] ^ n[27009];
assign t[27010] = t[27009] ^ n[27010];
assign t[27011] = t[27010] ^ n[27011];
assign t[27012] = t[27011] ^ n[27012];
assign t[27013] = t[27012] ^ n[27013];
assign t[27014] = t[27013] ^ n[27014];
assign t[27015] = t[27014] ^ n[27015];
assign t[27016] = t[27015] ^ n[27016];
assign t[27017] = t[27016] ^ n[27017];
assign t[27018] = t[27017] ^ n[27018];
assign t[27019] = t[27018] ^ n[27019];
assign t[27020] = t[27019] ^ n[27020];
assign t[27021] = t[27020] ^ n[27021];
assign t[27022] = t[27021] ^ n[27022];
assign t[27023] = t[27022] ^ n[27023];
assign t[27024] = t[27023] ^ n[27024];
assign t[27025] = t[27024] ^ n[27025];
assign t[27026] = t[27025] ^ n[27026];
assign t[27027] = t[27026] ^ n[27027];
assign t[27028] = t[27027] ^ n[27028];
assign t[27029] = t[27028] ^ n[27029];
assign t[27030] = t[27029] ^ n[27030];
assign t[27031] = t[27030] ^ n[27031];
assign t[27032] = t[27031] ^ n[27032];
assign t[27033] = t[27032] ^ n[27033];
assign t[27034] = t[27033] ^ n[27034];
assign t[27035] = t[27034] ^ n[27035];
assign t[27036] = t[27035] ^ n[27036];
assign t[27037] = t[27036] ^ n[27037];
assign t[27038] = t[27037] ^ n[27038];
assign t[27039] = t[27038] ^ n[27039];
assign t[27040] = t[27039] ^ n[27040];
assign t[27041] = t[27040] ^ n[27041];
assign t[27042] = t[27041] ^ n[27042];
assign t[27043] = t[27042] ^ n[27043];
assign t[27044] = t[27043] ^ n[27044];
assign t[27045] = t[27044] ^ n[27045];
assign t[27046] = t[27045] ^ n[27046];
assign t[27047] = t[27046] ^ n[27047];
assign t[27048] = t[27047] ^ n[27048];
assign t[27049] = t[27048] ^ n[27049];
assign t[27050] = t[27049] ^ n[27050];
assign t[27051] = t[27050] ^ n[27051];
assign t[27052] = t[27051] ^ n[27052];
assign t[27053] = t[27052] ^ n[27053];
assign t[27054] = t[27053] ^ n[27054];
assign t[27055] = t[27054] ^ n[27055];
assign t[27056] = t[27055] ^ n[27056];
assign t[27057] = t[27056] ^ n[27057];
assign t[27058] = t[27057] ^ n[27058];
assign t[27059] = t[27058] ^ n[27059];
assign t[27060] = t[27059] ^ n[27060];
assign t[27061] = t[27060] ^ n[27061];
assign t[27062] = t[27061] ^ n[27062];
assign t[27063] = t[27062] ^ n[27063];
assign t[27064] = t[27063] ^ n[27064];
assign t[27065] = t[27064] ^ n[27065];
assign t[27066] = t[27065] ^ n[27066];
assign t[27067] = t[27066] ^ n[27067];
assign t[27068] = t[27067] ^ n[27068];
assign t[27069] = t[27068] ^ n[27069];
assign t[27070] = t[27069] ^ n[27070];
assign t[27071] = t[27070] ^ n[27071];
assign t[27072] = t[27071] ^ n[27072];
assign t[27073] = t[27072] ^ n[27073];
assign t[27074] = t[27073] ^ n[27074];
assign t[27075] = t[27074] ^ n[27075];
assign t[27076] = t[27075] ^ n[27076];
assign t[27077] = t[27076] ^ n[27077];
assign t[27078] = t[27077] ^ n[27078];
assign t[27079] = t[27078] ^ n[27079];
assign t[27080] = t[27079] ^ n[27080];
assign t[27081] = t[27080] ^ n[27081];
assign t[27082] = t[27081] ^ n[27082];
assign t[27083] = t[27082] ^ n[27083];
assign t[27084] = t[27083] ^ n[27084];
assign t[27085] = t[27084] ^ n[27085];
assign t[27086] = t[27085] ^ n[27086];
assign t[27087] = t[27086] ^ n[27087];
assign t[27088] = t[27087] ^ n[27088];
assign t[27089] = t[27088] ^ n[27089];
assign t[27090] = t[27089] ^ n[27090];
assign t[27091] = t[27090] ^ n[27091];
assign t[27092] = t[27091] ^ n[27092];
assign t[27093] = t[27092] ^ n[27093];
assign t[27094] = t[27093] ^ n[27094];
assign t[27095] = t[27094] ^ n[27095];
assign t[27096] = t[27095] ^ n[27096];
assign t[27097] = t[27096] ^ n[27097];
assign t[27098] = t[27097] ^ n[27098];
assign t[27099] = t[27098] ^ n[27099];
assign t[27100] = t[27099] ^ n[27100];
assign t[27101] = t[27100] ^ n[27101];
assign t[27102] = t[27101] ^ n[27102];
assign t[27103] = t[27102] ^ n[27103];
assign t[27104] = t[27103] ^ n[27104];
assign t[27105] = t[27104] ^ n[27105];
assign t[27106] = t[27105] ^ n[27106];
assign t[27107] = t[27106] ^ n[27107];
assign t[27108] = t[27107] ^ n[27108];
assign t[27109] = t[27108] ^ n[27109];
assign t[27110] = t[27109] ^ n[27110];
assign t[27111] = t[27110] ^ n[27111];
assign t[27112] = t[27111] ^ n[27112];
assign t[27113] = t[27112] ^ n[27113];
assign t[27114] = t[27113] ^ n[27114];
assign t[27115] = t[27114] ^ n[27115];
assign t[27116] = t[27115] ^ n[27116];
assign t[27117] = t[27116] ^ n[27117];
assign t[27118] = t[27117] ^ n[27118];
assign t[27119] = t[27118] ^ n[27119];
assign t[27120] = t[27119] ^ n[27120];
assign t[27121] = t[27120] ^ n[27121];
assign t[27122] = t[27121] ^ n[27122];
assign t[27123] = t[27122] ^ n[27123];
assign t[27124] = t[27123] ^ n[27124];
assign t[27125] = t[27124] ^ n[27125];
assign t[27126] = t[27125] ^ n[27126];
assign t[27127] = t[27126] ^ n[27127];
assign t[27128] = t[27127] ^ n[27128];
assign t[27129] = t[27128] ^ n[27129];
assign t[27130] = t[27129] ^ n[27130];
assign t[27131] = t[27130] ^ n[27131];
assign t[27132] = t[27131] ^ n[27132];
assign t[27133] = t[27132] ^ n[27133];
assign t[27134] = t[27133] ^ n[27134];
assign t[27135] = t[27134] ^ n[27135];
assign t[27136] = t[27135] ^ n[27136];
assign t[27137] = t[27136] ^ n[27137];
assign t[27138] = t[27137] ^ n[27138];
assign t[27139] = t[27138] ^ n[27139];
assign t[27140] = t[27139] ^ n[27140];
assign t[27141] = t[27140] ^ n[27141];
assign t[27142] = t[27141] ^ n[27142];
assign t[27143] = t[27142] ^ n[27143];
assign t[27144] = t[27143] ^ n[27144];
assign t[27145] = t[27144] ^ n[27145];
assign t[27146] = t[27145] ^ n[27146];
assign t[27147] = t[27146] ^ n[27147];
assign t[27148] = t[27147] ^ n[27148];
assign t[27149] = t[27148] ^ n[27149];
assign t[27150] = t[27149] ^ n[27150];
assign t[27151] = t[27150] ^ n[27151];
assign t[27152] = t[27151] ^ n[27152];
assign t[27153] = t[27152] ^ n[27153];
assign t[27154] = t[27153] ^ n[27154];
assign t[27155] = t[27154] ^ n[27155];
assign t[27156] = t[27155] ^ n[27156];
assign t[27157] = t[27156] ^ n[27157];
assign t[27158] = t[27157] ^ n[27158];
assign t[27159] = t[27158] ^ n[27159];
assign t[27160] = t[27159] ^ n[27160];
assign t[27161] = t[27160] ^ n[27161];
assign t[27162] = t[27161] ^ n[27162];
assign t[27163] = t[27162] ^ n[27163];
assign t[27164] = t[27163] ^ n[27164];
assign t[27165] = t[27164] ^ n[27165];
assign t[27166] = t[27165] ^ n[27166];
assign t[27167] = t[27166] ^ n[27167];
assign t[27168] = t[27167] ^ n[27168];
assign t[27169] = t[27168] ^ n[27169];
assign t[27170] = t[27169] ^ n[27170];
assign t[27171] = t[27170] ^ n[27171];
assign t[27172] = t[27171] ^ n[27172];
assign t[27173] = t[27172] ^ n[27173];
assign t[27174] = t[27173] ^ n[27174];
assign t[27175] = t[27174] ^ n[27175];
assign t[27176] = t[27175] ^ n[27176];
assign t[27177] = t[27176] ^ n[27177];
assign t[27178] = t[27177] ^ n[27178];
assign t[27179] = t[27178] ^ n[27179];
assign t[27180] = t[27179] ^ n[27180];
assign t[27181] = t[27180] ^ n[27181];
assign t[27182] = t[27181] ^ n[27182];
assign t[27183] = t[27182] ^ n[27183];
assign t[27184] = t[27183] ^ n[27184];
assign t[27185] = t[27184] ^ n[27185];
assign t[27186] = t[27185] ^ n[27186];
assign t[27187] = t[27186] ^ n[27187];
assign t[27188] = t[27187] ^ n[27188];
assign t[27189] = t[27188] ^ n[27189];
assign t[27190] = t[27189] ^ n[27190];
assign t[27191] = t[27190] ^ n[27191];
assign t[27192] = t[27191] ^ n[27192];
assign t[27193] = t[27192] ^ n[27193];
assign t[27194] = t[27193] ^ n[27194];
assign t[27195] = t[27194] ^ n[27195];
assign t[27196] = t[27195] ^ n[27196];
assign t[27197] = t[27196] ^ n[27197];
assign t[27198] = t[27197] ^ n[27198];
assign t[27199] = t[27198] ^ n[27199];
assign t[27200] = t[27199] ^ n[27200];
assign t[27201] = t[27200] ^ n[27201];
assign t[27202] = t[27201] ^ n[27202];
assign t[27203] = t[27202] ^ n[27203];
assign t[27204] = t[27203] ^ n[27204];
assign t[27205] = t[27204] ^ n[27205];
assign t[27206] = t[27205] ^ n[27206];
assign t[27207] = t[27206] ^ n[27207];
assign t[27208] = t[27207] ^ n[27208];
assign t[27209] = t[27208] ^ n[27209];
assign t[27210] = t[27209] ^ n[27210];
assign t[27211] = t[27210] ^ n[27211];
assign t[27212] = t[27211] ^ n[27212];
assign t[27213] = t[27212] ^ n[27213];
assign t[27214] = t[27213] ^ n[27214];
assign t[27215] = t[27214] ^ n[27215];
assign t[27216] = t[27215] ^ n[27216];
assign t[27217] = t[27216] ^ n[27217];
assign t[27218] = t[27217] ^ n[27218];
assign t[27219] = t[27218] ^ n[27219];
assign t[27220] = t[27219] ^ n[27220];
assign t[27221] = t[27220] ^ n[27221];
assign t[27222] = t[27221] ^ n[27222];
assign t[27223] = t[27222] ^ n[27223];
assign t[27224] = t[27223] ^ n[27224];
assign t[27225] = t[27224] ^ n[27225];
assign t[27226] = t[27225] ^ n[27226];
assign t[27227] = t[27226] ^ n[27227];
assign t[27228] = t[27227] ^ n[27228];
assign t[27229] = t[27228] ^ n[27229];
assign t[27230] = t[27229] ^ n[27230];
assign t[27231] = t[27230] ^ n[27231];
assign t[27232] = t[27231] ^ n[27232];
assign t[27233] = t[27232] ^ n[27233];
assign t[27234] = t[27233] ^ n[27234];
assign t[27235] = t[27234] ^ n[27235];
assign t[27236] = t[27235] ^ n[27236];
assign t[27237] = t[27236] ^ n[27237];
assign t[27238] = t[27237] ^ n[27238];
assign t[27239] = t[27238] ^ n[27239];
assign t[27240] = t[27239] ^ n[27240];
assign t[27241] = t[27240] ^ n[27241];
assign t[27242] = t[27241] ^ n[27242];
assign t[27243] = t[27242] ^ n[27243];
assign t[27244] = t[27243] ^ n[27244];
assign t[27245] = t[27244] ^ n[27245];
assign t[27246] = t[27245] ^ n[27246];
assign t[27247] = t[27246] ^ n[27247];
assign t[27248] = t[27247] ^ n[27248];
assign t[27249] = t[27248] ^ n[27249];
assign t[27250] = t[27249] ^ n[27250];
assign t[27251] = t[27250] ^ n[27251];
assign t[27252] = t[27251] ^ n[27252];
assign t[27253] = t[27252] ^ n[27253];
assign t[27254] = t[27253] ^ n[27254];
assign t[27255] = t[27254] ^ n[27255];
assign t[27256] = t[27255] ^ n[27256];
assign t[27257] = t[27256] ^ n[27257];
assign t[27258] = t[27257] ^ n[27258];
assign t[27259] = t[27258] ^ n[27259];
assign t[27260] = t[27259] ^ n[27260];
assign t[27261] = t[27260] ^ n[27261];
assign t[27262] = t[27261] ^ n[27262];
assign t[27263] = t[27262] ^ n[27263];
assign t[27264] = t[27263] ^ n[27264];
assign t[27265] = t[27264] ^ n[27265];
assign t[27266] = t[27265] ^ n[27266];
assign t[27267] = t[27266] ^ n[27267];
assign t[27268] = t[27267] ^ n[27268];
assign t[27269] = t[27268] ^ n[27269];
assign t[27270] = t[27269] ^ n[27270];
assign t[27271] = t[27270] ^ n[27271];
assign t[27272] = t[27271] ^ n[27272];
assign t[27273] = t[27272] ^ n[27273];
assign t[27274] = t[27273] ^ n[27274];
assign t[27275] = t[27274] ^ n[27275];
assign t[27276] = t[27275] ^ n[27276];
assign t[27277] = t[27276] ^ n[27277];
assign t[27278] = t[27277] ^ n[27278];
assign t[27279] = t[27278] ^ n[27279];
assign t[27280] = t[27279] ^ n[27280];
assign t[27281] = t[27280] ^ n[27281];
assign t[27282] = t[27281] ^ n[27282];
assign t[27283] = t[27282] ^ n[27283];
assign t[27284] = t[27283] ^ n[27284];
assign t[27285] = t[27284] ^ n[27285];
assign t[27286] = t[27285] ^ n[27286];
assign t[27287] = t[27286] ^ n[27287];
assign t[27288] = t[27287] ^ n[27288];
assign t[27289] = t[27288] ^ n[27289];
assign t[27290] = t[27289] ^ n[27290];
assign t[27291] = t[27290] ^ n[27291];
assign t[27292] = t[27291] ^ n[27292];
assign t[27293] = t[27292] ^ n[27293];
assign t[27294] = t[27293] ^ n[27294];
assign t[27295] = t[27294] ^ n[27295];
assign t[27296] = t[27295] ^ n[27296];
assign t[27297] = t[27296] ^ n[27297];
assign t[27298] = t[27297] ^ n[27298];
assign t[27299] = t[27298] ^ n[27299];
assign t[27300] = t[27299] ^ n[27300];
assign t[27301] = t[27300] ^ n[27301];
assign t[27302] = t[27301] ^ n[27302];
assign t[27303] = t[27302] ^ n[27303];
assign t[27304] = t[27303] ^ n[27304];
assign t[27305] = t[27304] ^ n[27305];
assign t[27306] = t[27305] ^ n[27306];
assign t[27307] = t[27306] ^ n[27307];
assign t[27308] = t[27307] ^ n[27308];
assign t[27309] = t[27308] ^ n[27309];
assign t[27310] = t[27309] ^ n[27310];
assign t[27311] = t[27310] ^ n[27311];
assign t[27312] = t[27311] ^ n[27312];
assign t[27313] = t[27312] ^ n[27313];
assign t[27314] = t[27313] ^ n[27314];
assign t[27315] = t[27314] ^ n[27315];
assign t[27316] = t[27315] ^ n[27316];
assign t[27317] = t[27316] ^ n[27317];
assign t[27318] = t[27317] ^ n[27318];
assign t[27319] = t[27318] ^ n[27319];
assign t[27320] = t[27319] ^ n[27320];
assign t[27321] = t[27320] ^ n[27321];
assign t[27322] = t[27321] ^ n[27322];
assign t[27323] = t[27322] ^ n[27323];
assign t[27324] = t[27323] ^ n[27324];
assign t[27325] = t[27324] ^ n[27325];
assign t[27326] = t[27325] ^ n[27326];
assign t[27327] = t[27326] ^ n[27327];
assign t[27328] = t[27327] ^ n[27328];
assign t[27329] = t[27328] ^ n[27329];
assign t[27330] = t[27329] ^ n[27330];
assign t[27331] = t[27330] ^ n[27331];
assign t[27332] = t[27331] ^ n[27332];
assign t[27333] = t[27332] ^ n[27333];
assign t[27334] = t[27333] ^ n[27334];
assign t[27335] = t[27334] ^ n[27335];
assign t[27336] = t[27335] ^ n[27336];
assign t[27337] = t[27336] ^ n[27337];
assign t[27338] = t[27337] ^ n[27338];
assign t[27339] = t[27338] ^ n[27339];
assign t[27340] = t[27339] ^ n[27340];
assign t[27341] = t[27340] ^ n[27341];
assign t[27342] = t[27341] ^ n[27342];
assign t[27343] = t[27342] ^ n[27343];
assign t[27344] = t[27343] ^ n[27344];
assign t[27345] = t[27344] ^ n[27345];
assign t[27346] = t[27345] ^ n[27346];
assign t[27347] = t[27346] ^ n[27347];
assign t[27348] = t[27347] ^ n[27348];
assign t[27349] = t[27348] ^ n[27349];
assign t[27350] = t[27349] ^ n[27350];
assign t[27351] = t[27350] ^ n[27351];
assign t[27352] = t[27351] ^ n[27352];
assign t[27353] = t[27352] ^ n[27353];
assign t[27354] = t[27353] ^ n[27354];
assign t[27355] = t[27354] ^ n[27355];
assign t[27356] = t[27355] ^ n[27356];
assign t[27357] = t[27356] ^ n[27357];
assign t[27358] = t[27357] ^ n[27358];
assign t[27359] = t[27358] ^ n[27359];
assign t[27360] = t[27359] ^ n[27360];
assign t[27361] = t[27360] ^ n[27361];
assign t[27362] = t[27361] ^ n[27362];
assign t[27363] = t[27362] ^ n[27363];
assign t[27364] = t[27363] ^ n[27364];
assign t[27365] = t[27364] ^ n[27365];
assign t[27366] = t[27365] ^ n[27366];
assign t[27367] = t[27366] ^ n[27367];
assign t[27368] = t[27367] ^ n[27368];
assign t[27369] = t[27368] ^ n[27369];
assign t[27370] = t[27369] ^ n[27370];
assign t[27371] = t[27370] ^ n[27371];
assign t[27372] = t[27371] ^ n[27372];
assign t[27373] = t[27372] ^ n[27373];
assign t[27374] = t[27373] ^ n[27374];
assign t[27375] = t[27374] ^ n[27375];
assign t[27376] = t[27375] ^ n[27376];
assign t[27377] = t[27376] ^ n[27377];
assign t[27378] = t[27377] ^ n[27378];
assign t[27379] = t[27378] ^ n[27379];
assign t[27380] = t[27379] ^ n[27380];
assign t[27381] = t[27380] ^ n[27381];
assign t[27382] = t[27381] ^ n[27382];
assign t[27383] = t[27382] ^ n[27383];
assign t[27384] = t[27383] ^ n[27384];
assign t[27385] = t[27384] ^ n[27385];
assign t[27386] = t[27385] ^ n[27386];
assign t[27387] = t[27386] ^ n[27387];
assign t[27388] = t[27387] ^ n[27388];
assign t[27389] = t[27388] ^ n[27389];
assign t[27390] = t[27389] ^ n[27390];
assign t[27391] = t[27390] ^ n[27391];
assign t[27392] = t[27391] ^ n[27392];
assign t[27393] = t[27392] ^ n[27393];
assign t[27394] = t[27393] ^ n[27394];
assign t[27395] = t[27394] ^ n[27395];
assign t[27396] = t[27395] ^ n[27396];
assign t[27397] = t[27396] ^ n[27397];
assign t[27398] = t[27397] ^ n[27398];
assign t[27399] = t[27398] ^ n[27399];
assign t[27400] = t[27399] ^ n[27400];
assign t[27401] = t[27400] ^ n[27401];
assign t[27402] = t[27401] ^ n[27402];
assign t[27403] = t[27402] ^ n[27403];
assign t[27404] = t[27403] ^ n[27404];
assign t[27405] = t[27404] ^ n[27405];
assign t[27406] = t[27405] ^ n[27406];
assign t[27407] = t[27406] ^ n[27407];
assign t[27408] = t[27407] ^ n[27408];
assign t[27409] = t[27408] ^ n[27409];
assign t[27410] = t[27409] ^ n[27410];
assign t[27411] = t[27410] ^ n[27411];
assign t[27412] = t[27411] ^ n[27412];
assign t[27413] = t[27412] ^ n[27413];
assign t[27414] = t[27413] ^ n[27414];
assign t[27415] = t[27414] ^ n[27415];
assign t[27416] = t[27415] ^ n[27416];
assign t[27417] = t[27416] ^ n[27417];
assign t[27418] = t[27417] ^ n[27418];
assign t[27419] = t[27418] ^ n[27419];
assign t[27420] = t[27419] ^ n[27420];
assign t[27421] = t[27420] ^ n[27421];
assign t[27422] = t[27421] ^ n[27422];
assign t[27423] = t[27422] ^ n[27423];
assign t[27424] = t[27423] ^ n[27424];
assign t[27425] = t[27424] ^ n[27425];
assign t[27426] = t[27425] ^ n[27426];
assign t[27427] = t[27426] ^ n[27427];
assign t[27428] = t[27427] ^ n[27428];
assign t[27429] = t[27428] ^ n[27429];
assign t[27430] = t[27429] ^ n[27430];
assign t[27431] = t[27430] ^ n[27431];
assign t[27432] = t[27431] ^ n[27432];
assign t[27433] = t[27432] ^ n[27433];
assign t[27434] = t[27433] ^ n[27434];
assign t[27435] = t[27434] ^ n[27435];
assign t[27436] = t[27435] ^ n[27436];
assign t[27437] = t[27436] ^ n[27437];
assign t[27438] = t[27437] ^ n[27438];
assign t[27439] = t[27438] ^ n[27439];
assign t[27440] = t[27439] ^ n[27440];
assign t[27441] = t[27440] ^ n[27441];
assign t[27442] = t[27441] ^ n[27442];
assign t[27443] = t[27442] ^ n[27443];
assign t[27444] = t[27443] ^ n[27444];
assign t[27445] = t[27444] ^ n[27445];
assign t[27446] = t[27445] ^ n[27446];
assign t[27447] = t[27446] ^ n[27447];
assign t[27448] = t[27447] ^ n[27448];
assign t[27449] = t[27448] ^ n[27449];
assign t[27450] = t[27449] ^ n[27450];
assign t[27451] = t[27450] ^ n[27451];
assign t[27452] = t[27451] ^ n[27452];
assign t[27453] = t[27452] ^ n[27453];
assign t[27454] = t[27453] ^ n[27454];
assign t[27455] = t[27454] ^ n[27455];
assign t[27456] = t[27455] ^ n[27456];
assign t[27457] = t[27456] ^ n[27457];
assign t[27458] = t[27457] ^ n[27458];
assign t[27459] = t[27458] ^ n[27459];
assign t[27460] = t[27459] ^ n[27460];
assign t[27461] = t[27460] ^ n[27461];
assign t[27462] = t[27461] ^ n[27462];
assign t[27463] = t[27462] ^ n[27463];
assign t[27464] = t[27463] ^ n[27464];
assign t[27465] = t[27464] ^ n[27465];
assign t[27466] = t[27465] ^ n[27466];
assign t[27467] = t[27466] ^ n[27467];
assign t[27468] = t[27467] ^ n[27468];
assign t[27469] = t[27468] ^ n[27469];
assign t[27470] = t[27469] ^ n[27470];
assign t[27471] = t[27470] ^ n[27471];
assign t[27472] = t[27471] ^ n[27472];
assign t[27473] = t[27472] ^ n[27473];
assign t[27474] = t[27473] ^ n[27474];
assign t[27475] = t[27474] ^ n[27475];
assign t[27476] = t[27475] ^ n[27476];
assign t[27477] = t[27476] ^ n[27477];
assign t[27478] = t[27477] ^ n[27478];
assign t[27479] = t[27478] ^ n[27479];
assign t[27480] = t[27479] ^ n[27480];
assign t[27481] = t[27480] ^ n[27481];
assign t[27482] = t[27481] ^ n[27482];
assign t[27483] = t[27482] ^ n[27483];
assign t[27484] = t[27483] ^ n[27484];
assign t[27485] = t[27484] ^ n[27485];
assign t[27486] = t[27485] ^ n[27486];
assign t[27487] = t[27486] ^ n[27487];
assign t[27488] = t[27487] ^ n[27488];
assign t[27489] = t[27488] ^ n[27489];
assign t[27490] = t[27489] ^ n[27490];
assign t[27491] = t[27490] ^ n[27491];
assign t[27492] = t[27491] ^ n[27492];
assign t[27493] = t[27492] ^ n[27493];
assign t[27494] = t[27493] ^ n[27494];
assign t[27495] = t[27494] ^ n[27495];
assign t[27496] = t[27495] ^ n[27496];
assign t[27497] = t[27496] ^ n[27497];
assign t[27498] = t[27497] ^ n[27498];
assign t[27499] = t[27498] ^ n[27499];
assign t[27500] = t[27499] ^ n[27500];
assign t[27501] = t[27500] ^ n[27501];
assign t[27502] = t[27501] ^ n[27502];
assign t[27503] = t[27502] ^ n[27503];
assign t[27504] = t[27503] ^ n[27504];
assign t[27505] = t[27504] ^ n[27505];
assign t[27506] = t[27505] ^ n[27506];
assign t[27507] = t[27506] ^ n[27507];
assign t[27508] = t[27507] ^ n[27508];
assign t[27509] = t[27508] ^ n[27509];
assign t[27510] = t[27509] ^ n[27510];
assign t[27511] = t[27510] ^ n[27511];
assign t[27512] = t[27511] ^ n[27512];
assign t[27513] = t[27512] ^ n[27513];
assign t[27514] = t[27513] ^ n[27514];
assign t[27515] = t[27514] ^ n[27515];
assign t[27516] = t[27515] ^ n[27516];
assign t[27517] = t[27516] ^ n[27517];
assign t[27518] = t[27517] ^ n[27518];
assign t[27519] = t[27518] ^ n[27519];
assign t[27520] = t[27519] ^ n[27520];
assign t[27521] = t[27520] ^ n[27521];
assign t[27522] = t[27521] ^ n[27522];
assign t[27523] = t[27522] ^ n[27523];
assign t[27524] = t[27523] ^ n[27524];
assign t[27525] = t[27524] ^ n[27525];
assign t[27526] = t[27525] ^ n[27526];
assign t[27527] = t[27526] ^ n[27527];
assign t[27528] = t[27527] ^ n[27528];
assign t[27529] = t[27528] ^ n[27529];
assign t[27530] = t[27529] ^ n[27530];
assign t[27531] = t[27530] ^ n[27531];
assign t[27532] = t[27531] ^ n[27532];
assign t[27533] = t[27532] ^ n[27533];
assign t[27534] = t[27533] ^ n[27534];
assign t[27535] = t[27534] ^ n[27535];
assign t[27536] = t[27535] ^ n[27536];
assign t[27537] = t[27536] ^ n[27537];
assign t[27538] = t[27537] ^ n[27538];
assign t[27539] = t[27538] ^ n[27539];
assign t[27540] = t[27539] ^ n[27540];
assign t[27541] = t[27540] ^ n[27541];
assign t[27542] = t[27541] ^ n[27542];
assign t[27543] = t[27542] ^ n[27543];
assign t[27544] = t[27543] ^ n[27544];
assign t[27545] = t[27544] ^ n[27545];
assign t[27546] = t[27545] ^ n[27546];
assign t[27547] = t[27546] ^ n[27547];
assign t[27548] = t[27547] ^ n[27548];
assign t[27549] = t[27548] ^ n[27549];
assign t[27550] = t[27549] ^ n[27550];
assign t[27551] = t[27550] ^ n[27551];
assign t[27552] = t[27551] ^ n[27552];
assign t[27553] = t[27552] ^ n[27553];
assign t[27554] = t[27553] ^ n[27554];
assign t[27555] = t[27554] ^ n[27555];
assign t[27556] = t[27555] ^ n[27556];
assign t[27557] = t[27556] ^ n[27557];
assign t[27558] = t[27557] ^ n[27558];
assign t[27559] = t[27558] ^ n[27559];
assign t[27560] = t[27559] ^ n[27560];
assign t[27561] = t[27560] ^ n[27561];
assign t[27562] = t[27561] ^ n[27562];
assign t[27563] = t[27562] ^ n[27563];
assign t[27564] = t[27563] ^ n[27564];
assign t[27565] = t[27564] ^ n[27565];
assign t[27566] = t[27565] ^ n[27566];
assign t[27567] = t[27566] ^ n[27567];
assign t[27568] = t[27567] ^ n[27568];
assign t[27569] = t[27568] ^ n[27569];
assign t[27570] = t[27569] ^ n[27570];
assign t[27571] = t[27570] ^ n[27571];
assign t[27572] = t[27571] ^ n[27572];
assign t[27573] = t[27572] ^ n[27573];
assign t[27574] = t[27573] ^ n[27574];
assign t[27575] = t[27574] ^ n[27575];
assign t[27576] = t[27575] ^ n[27576];
assign t[27577] = t[27576] ^ n[27577];
assign t[27578] = t[27577] ^ n[27578];
assign t[27579] = t[27578] ^ n[27579];
assign t[27580] = t[27579] ^ n[27580];
assign t[27581] = t[27580] ^ n[27581];
assign t[27582] = t[27581] ^ n[27582];
assign t[27583] = t[27582] ^ n[27583];
assign t[27584] = t[27583] ^ n[27584];
assign t[27585] = t[27584] ^ n[27585];
assign t[27586] = t[27585] ^ n[27586];
assign t[27587] = t[27586] ^ n[27587];
assign t[27588] = t[27587] ^ n[27588];
assign t[27589] = t[27588] ^ n[27589];
assign t[27590] = t[27589] ^ n[27590];
assign t[27591] = t[27590] ^ n[27591];
assign t[27592] = t[27591] ^ n[27592];
assign t[27593] = t[27592] ^ n[27593];
assign t[27594] = t[27593] ^ n[27594];
assign t[27595] = t[27594] ^ n[27595];
assign t[27596] = t[27595] ^ n[27596];
assign t[27597] = t[27596] ^ n[27597];
assign t[27598] = t[27597] ^ n[27598];
assign t[27599] = t[27598] ^ n[27599];
assign t[27600] = t[27599] ^ n[27600];
assign t[27601] = t[27600] ^ n[27601];
assign t[27602] = t[27601] ^ n[27602];
assign t[27603] = t[27602] ^ n[27603];
assign t[27604] = t[27603] ^ n[27604];
assign t[27605] = t[27604] ^ n[27605];
assign t[27606] = t[27605] ^ n[27606];
assign t[27607] = t[27606] ^ n[27607];
assign t[27608] = t[27607] ^ n[27608];
assign t[27609] = t[27608] ^ n[27609];
assign t[27610] = t[27609] ^ n[27610];
assign t[27611] = t[27610] ^ n[27611];
assign t[27612] = t[27611] ^ n[27612];
assign t[27613] = t[27612] ^ n[27613];
assign t[27614] = t[27613] ^ n[27614];
assign t[27615] = t[27614] ^ n[27615];
assign t[27616] = t[27615] ^ n[27616];
assign t[27617] = t[27616] ^ n[27617];
assign t[27618] = t[27617] ^ n[27618];
assign t[27619] = t[27618] ^ n[27619];
assign t[27620] = t[27619] ^ n[27620];
assign t[27621] = t[27620] ^ n[27621];
assign t[27622] = t[27621] ^ n[27622];
assign t[27623] = t[27622] ^ n[27623];
assign t[27624] = t[27623] ^ n[27624];
assign t[27625] = t[27624] ^ n[27625];
assign t[27626] = t[27625] ^ n[27626];
assign t[27627] = t[27626] ^ n[27627];
assign t[27628] = t[27627] ^ n[27628];
assign t[27629] = t[27628] ^ n[27629];
assign t[27630] = t[27629] ^ n[27630];
assign t[27631] = t[27630] ^ n[27631];
assign t[27632] = t[27631] ^ n[27632];
assign t[27633] = t[27632] ^ n[27633];
assign t[27634] = t[27633] ^ n[27634];
assign t[27635] = t[27634] ^ n[27635];
assign t[27636] = t[27635] ^ n[27636];
assign t[27637] = t[27636] ^ n[27637];
assign t[27638] = t[27637] ^ n[27638];
assign t[27639] = t[27638] ^ n[27639];
assign t[27640] = t[27639] ^ n[27640];
assign t[27641] = t[27640] ^ n[27641];
assign t[27642] = t[27641] ^ n[27642];
assign t[27643] = t[27642] ^ n[27643];
assign t[27644] = t[27643] ^ n[27644];
assign t[27645] = t[27644] ^ n[27645];
assign t[27646] = t[27645] ^ n[27646];
assign t[27647] = t[27646] ^ n[27647];
assign t[27648] = t[27647] ^ n[27648];
assign t[27649] = t[27648] ^ n[27649];
assign t[27650] = t[27649] ^ n[27650];
assign t[27651] = t[27650] ^ n[27651];
assign t[27652] = t[27651] ^ n[27652];
assign t[27653] = t[27652] ^ n[27653];
assign t[27654] = t[27653] ^ n[27654];
assign t[27655] = t[27654] ^ n[27655];
assign t[27656] = t[27655] ^ n[27656];
assign t[27657] = t[27656] ^ n[27657];
assign t[27658] = t[27657] ^ n[27658];
assign t[27659] = t[27658] ^ n[27659];
assign t[27660] = t[27659] ^ n[27660];
assign t[27661] = t[27660] ^ n[27661];
assign t[27662] = t[27661] ^ n[27662];
assign t[27663] = t[27662] ^ n[27663];
assign t[27664] = t[27663] ^ n[27664];
assign t[27665] = t[27664] ^ n[27665];
assign t[27666] = t[27665] ^ n[27666];
assign t[27667] = t[27666] ^ n[27667];
assign t[27668] = t[27667] ^ n[27668];
assign t[27669] = t[27668] ^ n[27669];
assign t[27670] = t[27669] ^ n[27670];
assign t[27671] = t[27670] ^ n[27671];
assign t[27672] = t[27671] ^ n[27672];
assign t[27673] = t[27672] ^ n[27673];
assign t[27674] = t[27673] ^ n[27674];
assign t[27675] = t[27674] ^ n[27675];
assign t[27676] = t[27675] ^ n[27676];
assign t[27677] = t[27676] ^ n[27677];
assign t[27678] = t[27677] ^ n[27678];
assign t[27679] = t[27678] ^ n[27679];
assign t[27680] = t[27679] ^ n[27680];
assign t[27681] = t[27680] ^ n[27681];
assign t[27682] = t[27681] ^ n[27682];
assign t[27683] = t[27682] ^ n[27683];
assign t[27684] = t[27683] ^ n[27684];
assign t[27685] = t[27684] ^ n[27685];
assign t[27686] = t[27685] ^ n[27686];
assign t[27687] = t[27686] ^ n[27687];
assign t[27688] = t[27687] ^ n[27688];
assign t[27689] = t[27688] ^ n[27689];
assign t[27690] = t[27689] ^ n[27690];
assign t[27691] = t[27690] ^ n[27691];
assign t[27692] = t[27691] ^ n[27692];
assign t[27693] = t[27692] ^ n[27693];
assign t[27694] = t[27693] ^ n[27694];
assign t[27695] = t[27694] ^ n[27695];
assign t[27696] = t[27695] ^ n[27696];
assign t[27697] = t[27696] ^ n[27697];
assign t[27698] = t[27697] ^ n[27698];
assign t[27699] = t[27698] ^ n[27699];
assign t[27700] = t[27699] ^ n[27700];
assign t[27701] = t[27700] ^ n[27701];
assign t[27702] = t[27701] ^ n[27702];
assign t[27703] = t[27702] ^ n[27703];
assign t[27704] = t[27703] ^ n[27704];
assign t[27705] = t[27704] ^ n[27705];
assign t[27706] = t[27705] ^ n[27706];
assign t[27707] = t[27706] ^ n[27707];
assign t[27708] = t[27707] ^ n[27708];
assign t[27709] = t[27708] ^ n[27709];
assign t[27710] = t[27709] ^ n[27710];
assign t[27711] = t[27710] ^ n[27711];
assign t[27712] = t[27711] ^ n[27712];
assign t[27713] = t[27712] ^ n[27713];
assign t[27714] = t[27713] ^ n[27714];
assign t[27715] = t[27714] ^ n[27715];
assign t[27716] = t[27715] ^ n[27716];
assign t[27717] = t[27716] ^ n[27717];
assign t[27718] = t[27717] ^ n[27718];
assign t[27719] = t[27718] ^ n[27719];
assign t[27720] = t[27719] ^ n[27720];
assign t[27721] = t[27720] ^ n[27721];
assign t[27722] = t[27721] ^ n[27722];
assign t[27723] = t[27722] ^ n[27723];
assign t[27724] = t[27723] ^ n[27724];
assign t[27725] = t[27724] ^ n[27725];
assign t[27726] = t[27725] ^ n[27726];
assign t[27727] = t[27726] ^ n[27727];
assign t[27728] = t[27727] ^ n[27728];
assign t[27729] = t[27728] ^ n[27729];
assign t[27730] = t[27729] ^ n[27730];
assign t[27731] = t[27730] ^ n[27731];
assign t[27732] = t[27731] ^ n[27732];
assign t[27733] = t[27732] ^ n[27733];
assign t[27734] = t[27733] ^ n[27734];
assign t[27735] = t[27734] ^ n[27735];
assign t[27736] = t[27735] ^ n[27736];
assign t[27737] = t[27736] ^ n[27737];
assign t[27738] = t[27737] ^ n[27738];
assign t[27739] = t[27738] ^ n[27739];
assign t[27740] = t[27739] ^ n[27740];
assign t[27741] = t[27740] ^ n[27741];
assign t[27742] = t[27741] ^ n[27742];
assign t[27743] = t[27742] ^ n[27743];
assign t[27744] = t[27743] ^ n[27744];
assign t[27745] = t[27744] ^ n[27745];
assign t[27746] = t[27745] ^ n[27746];
assign t[27747] = t[27746] ^ n[27747];
assign t[27748] = t[27747] ^ n[27748];
assign t[27749] = t[27748] ^ n[27749];
assign t[27750] = t[27749] ^ n[27750];
assign t[27751] = t[27750] ^ n[27751];
assign t[27752] = t[27751] ^ n[27752];
assign t[27753] = t[27752] ^ n[27753];
assign t[27754] = t[27753] ^ n[27754];
assign t[27755] = t[27754] ^ n[27755];
assign t[27756] = t[27755] ^ n[27756];
assign t[27757] = t[27756] ^ n[27757];
assign t[27758] = t[27757] ^ n[27758];
assign t[27759] = t[27758] ^ n[27759];
assign t[27760] = t[27759] ^ n[27760];
assign t[27761] = t[27760] ^ n[27761];
assign t[27762] = t[27761] ^ n[27762];
assign t[27763] = t[27762] ^ n[27763];
assign t[27764] = t[27763] ^ n[27764];
assign t[27765] = t[27764] ^ n[27765];
assign t[27766] = t[27765] ^ n[27766];
assign t[27767] = t[27766] ^ n[27767];
assign t[27768] = t[27767] ^ n[27768];
assign t[27769] = t[27768] ^ n[27769];
assign t[27770] = t[27769] ^ n[27770];
assign t[27771] = t[27770] ^ n[27771];
assign t[27772] = t[27771] ^ n[27772];
assign t[27773] = t[27772] ^ n[27773];
assign t[27774] = t[27773] ^ n[27774];
assign t[27775] = t[27774] ^ n[27775];
assign t[27776] = t[27775] ^ n[27776];
assign t[27777] = t[27776] ^ n[27777];
assign t[27778] = t[27777] ^ n[27778];
assign t[27779] = t[27778] ^ n[27779];
assign t[27780] = t[27779] ^ n[27780];
assign t[27781] = t[27780] ^ n[27781];
assign t[27782] = t[27781] ^ n[27782];
assign t[27783] = t[27782] ^ n[27783];
assign t[27784] = t[27783] ^ n[27784];
assign t[27785] = t[27784] ^ n[27785];
assign t[27786] = t[27785] ^ n[27786];
assign t[27787] = t[27786] ^ n[27787];
assign t[27788] = t[27787] ^ n[27788];
assign t[27789] = t[27788] ^ n[27789];
assign t[27790] = t[27789] ^ n[27790];
assign t[27791] = t[27790] ^ n[27791];
assign t[27792] = t[27791] ^ n[27792];
assign t[27793] = t[27792] ^ n[27793];
assign t[27794] = t[27793] ^ n[27794];
assign t[27795] = t[27794] ^ n[27795];
assign t[27796] = t[27795] ^ n[27796];
assign t[27797] = t[27796] ^ n[27797];
assign t[27798] = t[27797] ^ n[27798];
assign t[27799] = t[27798] ^ n[27799];
assign t[27800] = t[27799] ^ n[27800];
assign t[27801] = t[27800] ^ n[27801];
assign t[27802] = t[27801] ^ n[27802];
assign t[27803] = t[27802] ^ n[27803];
assign t[27804] = t[27803] ^ n[27804];
assign t[27805] = t[27804] ^ n[27805];
assign t[27806] = t[27805] ^ n[27806];
assign t[27807] = t[27806] ^ n[27807];
assign t[27808] = t[27807] ^ n[27808];
assign t[27809] = t[27808] ^ n[27809];
assign t[27810] = t[27809] ^ n[27810];
assign t[27811] = t[27810] ^ n[27811];
assign t[27812] = t[27811] ^ n[27812];
assign t[27813] = t[27812] ^ n[27813];
assign t[27814] = t[27813] ^ n[27814];
assign t[27815] = t[27814] ^ n[27815];
assign t[27816] = t[27815] ^ n[27816];
assign t[27817] = t[27816] ^ n[27817];
assign t[27818] = t[27817] ^ n[27818];
assign t[27819] = t[27818] ^ n[27819];
assign t[27820] = t[27819] ^ n[27820];
assign t[27821] = t[27820] ^ n[27821];
assign t[27822] = t[27821] ^ n[27822];
assign t[27823] = t[27822] ^ n[27823];
assign t[27824] = t[27823] ^ n[27824];
assign t[27825] = t[27824] ^ n[27825];
assign t[27826] = t[27825] ^ n[27826];
assign t[27827] = t[27826] ^ n[27827];
assign t[27828] = t[27827] ^ n[27828];
assign t[27829] = t[27828] ^ n[27829];
assign t[27830] = t[27829] ^ n[27830];
assign t[27831] = t[27830] ^ n[27831];
assign t[27832] = t[27831] ^ n[27832];
assign t[27833] = t[27832] ^ n[27833];
assign t[27834] = t[27833] ^ n[27834];
assign t[27835] = t[27834] ^ n[27835];
assign t[27836] = t[27835] ^ n[27836];
assign t[27837] = t[27836] ^ n[27837];
assign t[27838] = t[27837] ^ n[27838];
assign t[27839] = t[27838] ^ n[27839];
assign t[27840] = t[27839] ^ n[27840];
assign t[27841] = t[27840] ^ n[27841];
assign t[27842] = t[27841] ^ n[27842];
assign t[27843] = t[27842] ^ n[27843];
assign t[27844] = t[27843] ^ n[27844];
assign t[27845] = t[27844] ^ n[27845];
assign t[27846] = t[27845] ^ n[27846];
assign t[27847] = t[27846] ^ n[27847];
assign t[27848] = t[27847] ^ n[27848];
assign t[27849] = t[27848] ^ n[27849];
assign t[27850] = t[27849] ^ n[27850];
assign t[27851] = t[27850] ^ n[27851];
assign t[27852] = t[27851] ^ n[27852];
assign t[27853] = t[27852] ^ n[27853];
assign t[27854] = t[27853] ^ n[27854];
assign t[27855] = t[27854] ^ n[27855];
assign t[27856] = t[27855] ^ n[27856];
assign t[27857] = t[27856] ^ n[27857];
assign t[27858] = t[27857] ^ n[27858];
assign t[27859] = t[27858] ^ n[27859];
assign t[27860] = t[27859] ^ n[27860];
assign t[27861] = t[27860] ^ n[27861];
assign t[27862] = t[27861] ^ n[27862];
assign t[27863] = t[27862] ^ n[27863];
assign t[27864] = t[27863] ^ n[27864];
assign t[27865] = t[27864] ^ n[27865];
assign t[27866] = t[27865] ^ n[27866];
assign t[27867] = t[27866] ^ n[27867];
assign t[27868] = t[27867] ^ n[27868];
assign t[27869] = t[27868] ^ n[27869];
assign t[27870] = t[27869] ^ n[27870];
assign t[27871] = t[27870] ^ n[27871];
assign t[27872] = t[27871] ^ n[27872];
assign t[27873] = t[27872] ^ n[27873];
assign t[27874] = t[27873] ^ n[27874];
assign t[27875] = t[27874] ^ n[27875];
assign t[27876] = t[27875] ^ n[27876];
assign t[27877] = t[27876] ^ n[27877];
assign t[27878] = t[27877] ^ n[27878];
assign t[27879] = t[27878] ^ n[27879];
assign t[27880] = t[27879] ^ n[27880];
assign t[27881] = t[27880] ^ n[27881];
assign t[27882] = t[27881] ^ n[27882];
assign t[27883] = t[27882] ^ n[27883];
assign t[27884] = t[27883] ^ n[27884];
assign t[27885] = t[27884] ^ n[27885];
assign t[27886] = t[27885] ^ n[27886];
assign t[27887] = t[27886] ^ n[27887];
assign t[27888] = t[27887] ^ n[27888];
assign t[27889] = t[27888] ^ n[27889];
assign t[27890] = t[27889] ^ n[27890];
assign t[27891] = t[27890] ^ n[27891];
assign t[27892] = t[27891] ^ n[27892];
assign t[27893] = t[27892] ^ n[27893];
assign t[27894] = t[27893] ^ n[27894];
assign t[27895] = t[27894] ^ n[27895];
assign t[27896] = t[27895] ^ n[27896];
assign t[27897] = t[27896] ^ n[27897];
assign t[27898] = t[27897] ^ n[27898];
assign t[27899] = t[27898] ^ n[27899];
assign t[27900] = t[27899] ^ n[27900];
assign t[27901] = t[27900] ^ n[27901];
assign t[27902] = t[27901] ^ n[27902];
assign t[27903] = t[27902] ^ n[27903];
assign t[27904] = t[27903] ^ n[27904];
assign t[27905] = t[27904] ^ n[27905];
assign t[27906] = t[27905] ^ n[27906];
assign t[27907] = t[27906] ^ n[27907];
assign t[27908] = t[27907] ^ n[27908];
assign t[27909] = t[27908] ^ n[27909];
assign t[27910] = t[27909] ^ n[27910];
assign t[27911] = t[27910] ^ n[27911];
assign t[27912] = t[27911] ^ n[27912];
assign t[27913] = t[27912] ^ n[27913];
assign t[27914] = t[27913] ^ n[27914];
assign t[27915] = t[27914] ^ n[27915];
assign t[27916] = t[27915] ^ n[27916];
assign t[27917] = t[27916] ^ n[27917];
assign t[27918] = t[27917] ^ n[27918];
assign t[27919] = t[27918] ^ n[27919];
assign t[27920] = t[27919] ^ n[27920];
assign t[27921] = t[27920] ^ n[27921];
assign t[27922] = t[27921] ^ n[27922];
assign t[27923] = t[27922] ^ n[27923];
assign t[27924] = t[27923] ^ n[27924];
assign t[27925] = t[27924] ^ n[27925];
assign t[27926] = t[27925] ^ n[27926];
assign t[27927] = t[27926] ^ n[27927];
assign t[27928] = t[27927] ^ n[27928];
assign t[27929] = t[27928] ^ n[27929];
assign t[27930] = t[27929] ^ n[27930];
assign t[27931] = t[27930] ^ n[27931];
assign t[27932] = t[27931] ^ n[27932];
assign t[27933] = t[27932] ^ n[27933];
assign t[27934] = t[27933] ^ n[27934];
assign t[27935] = t[27934] ^ n[27935];
assign t[27936] = t[27935] ^ n[27936];
assign t[27937] = t[27936] ^ n[27937];
assign t[27938] = t[27937] ^ n[27938];
assign t[27939] = t[27938] ^ n[27939];
assign t[27940] = t[27939] ^ n[27940];
assign t[27941] = t[27940] ^ n[27941];
assign t[27942] = t[27941] ^ n[27942];
assign t[27943] = t[27942] ^ n[27943];
assign t[27944] = t[27943] ^ n[27944];
assign t[27945] = t[27944] ^ n[27945];
assign t[27946] = t[27945] ^ n[27946];
assign t[27947] = t[27946] ^ n[27947];
assign t[27948] = t[27947] ^ n[27948];
assign t[27949] = t[27948] ^ n[27949];
assign t[27950] = t[27949] ^ n[27950];
assign t[27951] = t[27950] ^ n[27951];
assign t[27952] = t[27951] ^ n[27952];
assign t[27953] = t[27952] ^ n[27953];
assign t[27954] = t[27953] ^ n[27954];
assign t[27955] = t[27954] ^ n[27955];
assign t[27956] = t[27955] ^ n[27956];
assign t[27957] = t[27956] ^ n[27957];
assign t[27958] = t[27957] ^ n[27958];
assign t[27959] = t[27958] ^ n[27959];
assign t[27960] = t[27959] ^ n[27960];
assign t[27961] = t[27960] ^ n[27961];
assign t[27962] = t[27961] ^ n[27962];
assign t[27963] = t[27962] ^ n[27963];
assign t[27964] = t[27963] ^ n[27964];
assign t[27965] = t[27964] ^ n[27965];
assign t[27966] = t[27965] ^ n[27966];
assign t[27967] = t[27966] ^ n[27967];
assign t[27968] = t[27967] ^ n[27968];
assign t[27969] = t[27968] ^ n[27969];
assign t[27970] = t[27969] ^ n[27970];
assign t[27971] = t[27970] ^ n[27971];
assign t[27972] = t[27971] ^ n[27972];
assign t[27973] = t[27972] ^ n[27973];
assign t[27974] = t[27973] ^ n[27974];
assign t[27975] = t[27974] ^ n[27975];
assign t[27976] = t[27975] ^ n[27976];
assign t[27977] = t[27976] ^ n[27977];
assign t[27978] = t[27977] ^ n[27978];
assign t[27979] = t[27978] ^ n[27979];
assign t[27980] = t[27979] ^ n[27980];
assign t[27981] = t[27980] ^ n[27981];
assign t[27982] = t[27981] ^ n[27982];
assign t[27983] = t[27982] ^ n[27983];
assign t[27984] = t[27983] ^ n[27984];
assign t[27985] = t[27984] ^ n[27985];
assign t[27986] = t[27985] ^ n[27986];
assign t[27987] = t[27986] ^ n[27987];
assign t[27988] = t[27987] ^ n[27988];
assign t[27989] = t[27988] ^ n[27989];
assign t[27990] = t[27989] ^ n[27990];
assign t[27991] = t[27990] ^ n[27991];
assign t[27992] = t[27991] ^ n[27992];
assign t[27993] = t[27992] ^ n[27993];
assign t[27994] = t[27993] ^ n[27994];
assign t[27995] = t[27994] ^ n[27995];
assign t[27996] = t[27995] ^ n[27996];
assign t[27997] = t[27996] ^ n[27997];
assign t[27998] = t[27997] ^ n[27998];
assign t[27999] = t[27998] ^ n[27999];
assign t[28000] = t[27999] ^ n[28000];
assign t[28001] = t[28000] ^ n[28001];
assign t[28002] = t[28001] ^ n[28002];
assign t[28003] = t[28002] ^ n[28003];
assign t[28004] = t[28003] ^ n[28004];
assign t[28005] = t[28004] ^ n[28005];
assign t[28006] = t[28005] ^ n[28006];
assign t[28007] = t[28006] ^ n[28007];
assign t[28008] = t[28007] ^ n[28008];
assign t[28009] = t[28008] ^ n[28009];
assign t[28010] = t[28009] ^ n[28010];
assign t[28011] = t[28010] ^ n[28011];
assign t[28012] = t[28011] ^ n[28012];
assign t[28013] = t[28012] ^ n[28013];
assign t[28014] = t[28013] ^ n[28014];
assign t[28015] = t[28014] ^ n[28015];
assign t[28016] = t[28015] ^ n[28016];
assign t[28017] = t[28016] ^ n[28017];
assign t[28018] = t[28017] ^ n[28018];
assign t[28019] = t[28018] ^ n[28019];
assign t[28020] = t[28019] ^ n[28020];
assign t[28021] = t[28020] ^ n[28021];
assign t[28022] = t[28021] ^ n[28022];
assign t[28023] = t[28022] ^ n[28023];
assign t[28024] = t[28023] ^ n[28024];
assign t[28025] = t[28024] ^ n[28025];
assign t[28026] = t[28025] ^ n[28026];
assign t[28027] = t[28026] ^ n[28027];
assign t[28028] = t[28027] ^ n[28028];
assign t[28029] = t[28028] ^ n[28029];
assign t[28030] = t[28029] ^ n[28030];
assign t[28031] = t[28030] ^ n[28031];
assign t[28032] = t[28031] ^ n[28032];
assign t[28033] = t[28032] ^ n[28033];
assign t[28034] = t[28033] ^ n[28034];
assign t[28035] = t[28034] ^ n[28035];
assign t[28036] = t[28035] ^ n[28036];
assign t[28037] = t[28036] ^ n[28037];
assign t[28038] = t[28037] ^ n[28038];
assign t[28039] = t[28038] ^ n[28039];
assign t[28040] = t[28039] ^ n[28040];
assign t[28041] = t[28040] ^ n[28041];
assign t[28042] = t[28041] ^ n[28042];
assign t[28043] = t[28042] ^ n[28043];
assign t[28044] = t[28043] ^ n[28044];
assign t[28045] = t[28044] ^ n[28045];
assign t[28046] = t[28045] ^ n[28046];
assign t[28047] = t[28046] ^ n[28047];
assign t[28048] = t[28047] ^ n[28048];
assign t[28049] = t[28048] ^ n[28049];
assign t[28050] = t[28049] ^ n[28050];
assign t[28051] = t[28050] ^ n[28051];
assign t[28052] = t[28051] ^ n[28052];
assign t[28053] = t[28052] ^ n[28053];
assign t[28054] = t[28053] ^ n[28054];
assign t[28055] = t[28054] ^ n[28055];
assign t[28056] = t[28055] ^ n[28056];
assign t[28057] = t[28056] ^ n[28057];
assign t[28058] = t[28057] ^ n[28058];
assign t[28059] = t[28058] ^ n[28059];
assign t[28060] = t[28059] ^ n[28060];
assign t[28061] = t[28060] ^ n[28061];
assign t[28062] = t[28061] ^ n[28062];
assign t[28063] = t[28062] ^ n[28063];
assign t[28064] = t[28063] ^ n[28064];
assign t[28065] = t[28064] ^ n[28065];
assign t[28066] = t[28065] ^ n[28066];
assign t[28067] = t[28066] ^ n[28067];
assign t[28068] = t[28067] ^ n[28068];
assign t[28069] = t[28068] ^ n[28069];
assign t[28070] = t[28069] ^ n[28070];
assign t[28071] = t[28070] ^ n[28071];
assign t[28072] = t[28071] ^ n[28072];
assign t[28073] = t[28072] ^ n[28073];
assign t[28074] = t[28073] ^ n[28074];
assign t[28075] = t[28074] ^ n[28075];
assign t[28076] = t[28075] ^ n[28076];
assign t[28077] = t[28076] ^ n[28077];
assign t[28078] = t[28077] ^ n[28078];
assign t[28079] = t[28078] ^ n[28079];
assign t[28080] = t[28079] ^ n[28080];
assign t[28081] = t[28080] ^ n[28081];
assign t[28082] = t[28081] ^ n[28082];
assign t[28083] = t[28082] ^ n[28083];
assign t[28084] = t[28083] ^ n[28084];
assign t[28085] = t[28084] ^ n[28085];
assign t[28086] = t[28085] ^ n[28086];
assign t[28087] = t[28086] ^ n[28087];
assign t[28088] = t[28087] ^ n[28088];
assign t[28089] = t[28088] ^ n[28089];
assign t[28090] = t[28089] ^ n[28090];
assign t[28091] = t[28090] ^ n[28091];
assign t[28092] = t[28091] ^ n[28092];
assign t[28093] = t[28092] ^ n[28093];
assign t[28094] = t[28093] ^ n[28094];
assign t[28095] = t[28094] ^ n[28095];
assign t[28096] = t[28095] ^ n[28096];
assign t[28097] = t[28096] ^ n[28097];
assign t[28098] = t[28097] ^ n[28098];
assign t[28099] = t[28098] ^ n[28099];
assign t[28100] = t[28099] ^ n[28100];
assign t[28101] = t[28100] ^ n[28101];
assign t[28102] = t[28101] ^ n[28102];
assign t[28103] = t[28102] ^ n[28103];
assign t[28104] = t[28103] ^ n[28104];
assign t[28105] = t[28104] ^ n[28105];
assign t[28106] = t[28105] ^ n[28106];
assign t[28107] = t[28106] ^ n[28107];
assign t[28108] = t[28107] ^ n[28108];
assign t[28109] = t[28108] ^ n[28109];
assign t[28110] = t[28109] ^ n[28110];
assign t[28111] = t[28110] ^ n[28111];
assign t[28112] = t[28111] ^ n[28112];
assign t[28113] = t[28112] ^ n[28113];
assign t[28114] = t[28113] ^ n[28114];
assign t[28115] = t[28114] ^ n[28115];
assign t[28116] = t[28115] ^ n[28116];
assign t[28117] = t[28116] ^ n[28117];
assign t[28118] = t[28117] ^ n[28118];
assign t[28119] = t[28118] ^ n[28119];
assign t[28120] = t[28119] ^ n[28120];
assign t[28121] = t[28120] ^ n[28121];
assign t[28122] = t[28121] ^ n[28122];
assign t[28123] = t[28122] ^ n[28123];
assign t[28124] = t[28123] ^ n[28124];
assign t[28125] = t[28124] ^ n[28125];
assign t[28126] = t[28125] ^ n[28126];
assign t[28127] = t[28126] ^ n[28127];
assign t[28128] = t[28127] ^ n[28128];
assign t[28129] = t[28128] ^ n[28129];
assign t[28130] = t[28129] ^ n[28130];
assign t[28131] = t[28130] ^ n[28131];
assign t[28132] = t[28131] ^ n[28132];
assign t[28133] = t[28132] ^ n[28133];
assign t[28134] = t[28133] ^ n[28134];
assign t[28135] = t[28134] ^ n[28135];
assign t[28136] = t[28135] ^ n[28136];
assign t[28137] = t[28136] ^ n[28137];
assign t[28138] = t[28137] ^ n[28138];
assign t[28139] = t[28138] ^ n[28139];
assign t[28140] = t[28139] ^ n[28140];
assign t[28141] = t[28140] ^ n[28141];
assign t[28142] = t[28141] ^ n[28142];
assign t[28143] = t[28142] ^ n[28143];
assign t[28144] = t[28143] ^ n[28144];
assign t[28145] = t[28144] ^ n[28145];
assign t[28146] = t[28145] ^ n[28146];
assign t[28147] = t[28146] ^ n[28147];
assign t[28148] = t[28147] ^ n[28148];
assign t[28149] = t[28148] ^ n[28149];
assign t[28150] = t[28149] ^ n[28150];
assign t[28151] = t[28150] ^ n[28151];
assign t[28152] = t[28151] ^ n[28152];
assign t[28153] = t[28152] ^ n[28153];
assign t[28154] = t[28153] ^ n[28154];
assign t[28155] = t[28154] ^ n[28155];
assign t[28156] = t[28155] ^ n[28156];
assign t[28157] = t[28156] ^ n[28157];
assign t[28158] = t[28157] ^ n[28158];
assign t[28159] = t[28158] ^ n[28159];
assign t[28160] = t[28159] ^ n[28160];
assign t[28161] = t[28160] ^ n[28161];
assign t[28162] = t[28161] ^ n[28162];
assign t[28163] = t[28162] ^ n[28163];
assign t[28164] = t[28163] ^ n[28164];
assign t[28165] = t[28164] ^ n[28165];
assign t[28166] = t[28165] ^ n[28166];
assign t[28167] = t[28166] ^ n[28167];
assign t[28168] = t[28167] ^ n[28168];
assign t[28169] = t[28168] ^ n[28169];
assign t[28170] = t[28169] ^ n[28170];
assign t[28171] = t[28170] ^ n[28171];
assign t[28172] = t[28171] ^ n[28172];
assign t[28173] = t[28172] ^ n[28173];
assign t[28174] = t[28173] ^ n[28174];
assign t[28175] = t[28174] ^ n[28175];
assign t[28176] = t[28175] ^ n[28176];
assign t[28177] = t[28176] ^ n[28177];
assign t[28178] = t[28177] ^ n[28178];
assign t[28179] = t[28178] ^ n[28179];
assign t[28180] = t[28179] ^ n[28180];
assign t[28181] = t[28180] ^ n[28181];
assign t[28182] = t[28181] ^ n[28182];
assign t[28183] = t[28182] ^ n[28183];
assign t[28184] = t[28183] ^ n[28184];
assign t[28185] = t[28184] ^ n[28185];
assign t[28186] = t[28185] ^ n[28186];
assign t[28187] = t[28186] ^ n[28187];
assign t[28188] = t[28187] ^ n[28188];
assign t[28189] = t[28188] ^ n[28189];
assign t[28190] = t[28189] ^ n[28190];
assign t[28191] = t[28190] ^ n[28191];
assign t[28192] = t[28191] ^ n[28192];
assign t[28193] = t[28192] ^ n[28193];
assign t[28194] = t[28193] ^ n[28194];
assign t[28195] = t[28194] ^ n[28195];
assign t[28196] = t[28195] ^ n[28196];
assign t[28197] = t[28196] ^ n[28197];
assign t[28198] = t[28197] ^ n[28198];
assign t[28199] = t[28198] ^ n[28199];
assign t[28200] = t[28199] ^ n[28200];
assign t[28201] = t[28200] ^ n[28201];
assign t[28202] = t[28201] ^ n[28202];
assign t[28203] = t[28202] ^ n[28203];
assign t[28204] = t[28203] ^ n[28204];
assign t[28205] = t[28204] ^ n[28205];
assign t[28206] = t[28205] ^ n[28206];
assign t[28207] = t[28206] ^ n[28207];
assign t[28208] = t[28207] ^ n[28208];
assign t[28209] = t[28208] ^ n[28209];
assign t[28210] = t[28209] ^ n[28210];
assign t[28211] = t[28210] ^ n[28211];
assign t[28212] = t[28211] ^ n[28212];
assign t[28213] = t[28212] ^ n[28213];
assign t[28214] = t[28213] ^ n[28214];
assign t[28215] = t[28214] ^ n[28215];
assign t[28216] = t[28215] ^ n[28216];
assign t[28217] = t[28216] ^ n[28217];
assign t[28218] = t[28217] ^ n[28218];
assign t[28219] = t[28218] ^ n[28219];
assign t[28220] = t[28219] ^ n[28220];
assign t[28221] = t[28220] ^ n[28221];
assign t[28222] = t[28221] ^ n[28222];
assign t[28223] = t[28222] ^ n[28223];
assign t[28224] = t[28223] ^ n[28224];
assign t[28225] = t[28224] ^ n[28225];
assign t[28226] = t[28225] ^ n[28226];
assign t[28227] = t[28226] ^ n[28227];
assign t[28228] = t[28227] ^ n[28228];
assign t[28229] = t[28228] ^ n[28229];
assign t[28230] = t[28229] ^ n[28230];
assign t[28231] = t[28230] ^ n[28231];
assign t[28232] = t[28231] ^ n[28232];
assign t[28233] = t[28232] ^ n[28233];
assign t[28234] = t[28233] ^ n[28234];
assign t[28235] = t[28234] ^ n[28235];
assign t[28236] = t[28235] ^ n[28236];
assign t[28237] = t[28236] ^ n[28237];
assign t[28238] = t[28237] ^ n[28238];
assign t[28239] = t[28238] ^ n[28239];
assign t[28240] = t[28239] ^ n[28240];
assign t[28241] = t[28240] ^ n[28241];
assign t[28242] = t[28241] ^ n[28242];
assign t[28243] = t[28242] ^ n[28243];
assign t[28244] = t[28243] ^ n[28244];
assign t[28245] = t[28244] ^ n[28245];
assign t[28246] = t[28245] ^ n[28246];
assign t[28247] = t[28246] ^ n[28247];
assign t[28248] = t[28247] ^ n[28248];
assign t[28249] = t[28248] ^ n[28249];
assign t[28250] = t[28249] ^ n[28250];
assign t[28251] = t[28250] ^ n[28251];
assign t[28252] = t[28251] ^ n[28252];
assign t[28253] = t[28252] ^ n[28253];
assign t[28254] = t[28253] ^ n[28254];
assign t[28255] = t[28254] ^ n[28255];
assign t[28256] = t[28255] ^ n[28256];
assign t[28257] = t[28256] ^ n[28257];
assign t[28258] = t[28257] ^ n[28258];
assign t[28259] = t[28258] ^ n[28259];
assign t[28260] = t[28259] ^ n[28260];
assign t[28261] = t[28260] ^ n[28261];
assign t[28262] = t[28261] ^ n[28262];
assign t[28263] = t[28262] ^ n[28263];
assign t[28264] = t[28263] ^ n[28264];
assign t[28265] = t[28264] ^ n[28265];
assign t[28266] = t[28265] ^ n[28266];
assign t[28267] = t[28266] ^ n[28267];
assign t[28268] = t[28267] ^ n[28268];
assign t[28269] = t[28268] ^ n[28269];
assign t[28270] = t[28269] ^ n[28270];
assign t[28271] = t[28270] ^ n[28271];
assign t[28272] = t[28271] ^ n[28272];
assign t[28273] = t[28272] ^ n[28273];
assign t[28274] = t[28273] ^ n[28274];
assign t[28275] = t[28274] ^ n[28275];
assign t[28276] = t[28275] ^ n[28276];
assign t[28277] = t[28276] ^ n[28277];
assign t[28278] = t[28277] ^ n[28278];
assign t[28279] = t[28278] ^ n[28279];
assign t[28280] = t[28279] ^ n[28280];
assign t[28281] = t[28280] ^ n[28281];
assign t[28282] = t[28281] ^ n[28282];
assign t[28283] = t[28282] ^ n[28283];
assign t[28284] = t[28283] ^ n[28284];
assign t[28285] = t[28284] ^ n[28285];
assign t[28286] = t[28285] ^ n[28286];
assign t[28287] = t[28286] ^ n[28287];
assign t[28288] = t[28287] ^ n[28288];
assign t[28289] = t[28288] ^ n[28289];
assign t[28290] = t[28289] ^ n[28290];
assign t[28291] = t[28290] ^ n[28291];
assign t[28292] = t[28291] ^ n[28292];
assign t[28293] = t[28292] ^ n[28293];
assign t[28294] = t[28293] ^ n[28294];
assign t[28295] = t[28294] ^ n[28295];
assign t[28296] = t[28295] ^ n[28296];
assign t[28297] = t[28296] ^ n[28297];
assign t[28298] = t[28297] ^ n[28298];
assign t[28299] = t[28298] ^ n[28299];
assign t[28300] = t[28299] ^ n[28300];
assign t[28301] = t[28300] ^ n[28301];
assign t[28302] = t[28301] ^ n[28302];
assign t[28303] = t[28302] ^ n[28303];
assign t[28304] = t[28303] ^ n[28304];
assign t[28305] = t[28304] ^ n[28305];
assign t[28306] = t[28305] ^ n[28306];
assign t[28307] = t[28306] ^ n[28307];
assign t[28308] = t[28307] ^ n[28308];
assign t[28309] = t[28308] ^ n[28309];
assign t[28310] = t[28309] ^ n[28310];
assign t[28311] = t[28310] ^ n[28311];
assign t[28312] = t[28311] ^ n[28312];
assign t[28313] = t[28312] ^ n[28313];
assign t[28314] = t[28313] ^ n[28314];
assign t[28315] = t[28314] ^ n[28315];
assign t[28316] = t[28315] ^ n[28316];
assign t[28317] = t[28316] ^ n[28317];
assign t[28318] = t[28317] ^ n[28318];
assign t[28319] = t[28318] ^ n[28319];
assign t[28320] = t[28319] ^ n[28320];
assign t[28321] = t[28320] ^ n[28321];
assign t[28322] = t[28321] ^ n[28322];
assign t[28323] = t[28322] ^ n[28323];
assign t[28324] = t[28323] ^ n[28324];
assign t[28325] = t[28324] ^ n[28325];
assign t[28326] = t[28325] ^ n[28326];
assign t[28327] = t[28326] ^ n[28327];
assign t[28328] = t[28327] ^ n[28328];
assign t[28329] = t[28328] ^ n[28329];
assign t[28330] = t[28329] ^ n[28330];
assign t[28331] = t[28330] ^ n[28331];
assign t[28332] = t[28331] ^ n[28332];
assign t[28333] = t[28332] ^ n[28333];
assign t[28334] = t[28333] ^ n[28334];
assign t[28335] = t[28334] ^ n[28335];
assign t[28336] = t[28335] ^ n[28336];
assign t[28337] = t[28336] ^ n[28337];
assign t[28338] = t[28337] ^ n[28338];
assign t[28339] = t[28338] ^ n[28339];
assign t[28340] = t[28339] ^ n[28340];
assign t[28341] = t[28340] ^ n[28341];
assign t[28342] = t[28341] ^ n[28342];
assign t[28343] = t[28342] ^ n[28343];
assign t[28344] = t[28343] ^ n[28344];
assign t[28345] = t[28344] ^ n[28345];
assign t[28346] = t[28345] ^ n[28346];
assign t[28347] = t[28346] ^ n[28347];
assign t[28348] = t[28347] ^ n[28348];
assign t[28349] = t[28348] ^ n[28349];
assign t[28350] = t[28349] ^ n[28350];
assign t[28351] = t[28350] ^ n[28351];
assign t[28352] = t[28351] ^ n[28352];
assign t[28353] = t[28352] ^ n[28353];
assign t[28354] = t[28353] ^ n[28354];
assign t[28355] = t[28354] ^ n[28355];
assign t[28356] = t[28355] ^ n[28356];
assign t[28357] = t[28356] ^ n[28357];
assign t[28358] = t[28357] ^ n[28358];
assign t[28359] = t[28358] ^ n[28359];
assign t[28360] = t[28359] ^ n[28360];
assign t[28361] = t[28360] ^ n[28361];
assign t[28362] = t[28361] ^ n[28362];
assign t[28363] = t[28362] ^ n[28363];
assign t[28364] = t[28363] ^ n[28364];
assign t[28365] = t[28364] ^ n[28365];
assign t[28366] = t[28365] ^ n[28366];
assign t[28367] = t[28366] ^ n[28367];
assign t[28368] = t[28367] ^ n[28368];
assign t[28369] = t[28368] ^ n[28369];
assign t[28370] = t[28369] ^ n[28370];
assign t[28371] = t[28370] ^ n[28371];
assign t[28372] = t[28371] ^ n[28372];
assign t[28373] = t[28372] ^ n[28373];
assign t[28374] = t[28373] ^ n[28374];
assign t[28375] = t[28374] ^ n[28375];
assign t[28376] = t[28375] ^ n[28376];
assign t[28377] = t[28376] ^ n[28377];
assign t[28378] = t[28377] ^ n[28378];
assign t[28379] = t[28378] ^ n[28379];
assign t[28380] = t[28379] ^ n[28380];
assign t[28381] = t[28380] ^ n[28381];
assign t[28382] = t[28381] ^ n[28382];
assign t[28383] = t[28382] ^ n[28383];
assign t[28384] = t[28383] ^ n[28384];
assign t[28385] = t[28384] ^ n[28385];
assign t[28386] = t[28385] ^ n[28386];
assign t[28387] = t[28386] ^ n[28387];
assign t[28388] = t[28387] ^ n[28388];
assign t[28389] = t[28388] ^ n[28389];
assign t[28390] = t[28389] ^ n[28390];
assign t[28391] = t[28390] ^ n[28391];
assign t[28392] = t[28391] ^ n[28392];
assign t[28393] = t[28392] ^ n[28393];
assign t[28394] = t[28393] ^ n[28394];
assign t[28395] = t[28394] ^ n[28395];
assign t[28396] = t[28395] ^ n[28396];
assign t[28397] = t[28396] ^ n[28397];
assign t[28398] = t[28397] ^ n[28398];
assign t[28399] = t[28398] ^ n[28399];
assign t[28400] = t[28399] ^ n[28400];
assign t[28401] = t[28400] ^ n[28401];
assign t[28402] = t[28401] ^ n[28402];
assign t[28403] = t[28402] ^ n[28403];
assign t[28404] = t[28403] ^ n[28404];
assign t[28405] = t[28404] ^ n[28405];
assign t[28406] = t[28405] ^ n[28406];
assign t[28407] = t[28406] ^ n[28407];
assign t[28408] = t[28407] ^ n[28408];
assign t[28409] = t[28408] ^ n[28409];
assign t[28410] = t[28409] ^ n[28410];
assign t[28411] = t[28410] ^ n[28411];
assign t[28412] = t[28411] ^ n[28412];
assign t[28413] = t[28412] ^ n[28413];
assign t[28414] = t[28413] ^ n[28414];
assign t[28415] = t[28414] ^ n[28415];
assign t[28416] = t[28415] ^ n[28416];
assign t[28417] = t[28416] ^ n[28417];
assign t[28418] = t[28417] ^ n[28418];
assign t[28419] = t[28418] ^ n[28419];
assign t[28420] = t[28419] ^ n[28420];
assign t[28421] = t[28420] ^ n[28421];
assign t[28422] = t[28421] ^ n[28422];
assign t[28423] = t[28422] ^ n[28423];
assign t[28424] = t[28423] ^ n[28424];
assign t[28425] = t[28424] ^ n[28425];
assign t[28426] = t[28425] ^ n[28426];
assign t[28427] = t[28426] ^ n[28427];
assign t[28428] = t[28427] ^ n[28428];
assign t[28429] = t[28428] ^ n[28429];
assign t[28430] = t[28429] ^ n[28430];
assign t[28431] = t[28430] ^ n[28431];
assign t[28432] = t[28431] ^ n[28432];
assign t[28433] = t[28432] ^ n[28433];
assign t[28434] = t[28433] ^ n[28434];
assign t[28435] = t[28434] ^ n[28435];
assign t[28436] = t[28435] ^ n[28436];
assign t[28437] = t[28436] ^ n[28437];
assign t[28438] = t[28437] ^ n[28438];
assign t[28439] = t[28438] ^ n[28439];
assign t[28440] = t[28439] ^ n[28440];
assign t[28441] = t[28440] ^ n[28441];
assign t[28442] = t[28441] ^ n[28442];
assign t[28443] = t[28442] ^ n[28443];
assign t[28444] = t[28443] ^ n[28444];
assign t[28445] = t[28444] ^ n[28445];
assign t[28446] = t[28445] ^ n[28446];
assign t[28447] = t[28446] ^ n[28447];
assign t[28448] = t[28447] ^ n[28448];
assign t[28449] = t[28448] ^ n[28449];
assign t[28450] = t[28449] ^ n[28450];
assign t[28451] = t[28450] ^ n[28451];
assign t[28452] = t[28451] ^ n[28452];
assign t[28453] = t[28452] ^ n[28453];
assign t[28454] = t[28453] ^ n[28454];
assign t[28455] = t[28454] ^ n[28455];
assign t[28456] = t[28455] ^ n[28456];
assign t[28457] = t[28456] ^ n[28457];
assign t[28458] = t[28457] ^ n[28458];
assign t[28459] = t[28458] ^ n[28459];
assign t[28460] = t[28459] ^ n[28460];
assign t[28461] = t[28460] ^ n[28461];
assign t[28462] = t[28461] ^ n[28462];
assign t[28463] = t[28462] ^ n[28463];
assign t[28464] = t[28463] ^ n[28464];
assign t[28465] = t[28464] ^ n[28465];
assign t[28466] = t[28465] ^ n[28466];
assign t[28467] = t[28466] ^ n[28467];
assign t[28468] = t[28467] ^ n[28468];
assign t[28469] = t[28468] ^ n[28469];
assign t[28470] = t[28469] ^ n[28470];
assign t[28471] = t[28470] ^ n[28471];
assign t[28472] = t[28471] ^ n[28472];
assign t[28473] = t[28472] ^ n[28473];
assign t[28474] = t[28473] ^ n[28474];
assign t[28475] = t[28474] ^ n[28475];
assign t[28476] = t[28475] ^ n[28476];
assign t[28477] = t[28476] ^ n[28477];
assign t[28478] = t[28477] ^ n[28478];
assign t[28479] = t[28478] ^ n[28479];
assign t[28480] = t[28479] ^ n[28480];
assign t[28481] = t[28480] ^ n[28481];
assign t[28482] = t[28481] ^ n[28482];
assign t[28483] = t[28482] ^ n[28483];
assign t[28484] = t[28483] ^ n[28484];
assign t[28485] = t[28484] ^ n[28485];
assign t[28486] = t[28485] ^ n[28486];
assign t[28487] = t[28486] ^ n[28487];
assign t[28488] = t[28487] ^ n[28488];
assign t[28489] = t[28488] ^ n[28489];
assign t[28490] = t[28489] ^ n[28490];
assign t[28491] = t[28490] ^ n[28491];
assign t[28492] = t[28491] ^ n[28492];
assign t[28493] = t[28492] ^ n[28493];
assign t[28494] = t[28493] ^ n[28494];
assign t[28495] = t[28494] ^ n[28495];
assign t[28496] = t[28495] ^ n[28496];
assign t[28497] = t[28496] ^ n[28497];
assign t[28498] = t[28497] ^ n[28498];
assign t[28499] = t[28498] ^ n[28499];
assign t[28500] = t[28499] ^ n[28500];
assign t[28501] = t[28500] ^ n[28501];
assign t[28502] = t[28501] ^ n[28502];
assign t[28503] = t[28502] ^ n[28503];
assign t[28504] = t[28503] ^ n[28504];
assign t[28505] = t[28504] ^ n[28505];
assign t[28506] = t[28505] ^ n[28506];
assign t[28507] = t[28506] ^ n[28507];
assign t[28508] = t[28507] ^ n[28508];
assign t[28509] = t[28508] ^ n[28509];
assign t[28510] = t[28509] ^ n[28510];
assign t[28511] = t[28510] ^ n[28511];
assign t[28512] = t[28511] ^ n[28512];
assign t[28513] = t[28512] ^ n[28513];
assign t[28514] = t[28513] ^ n[28514];
assign t[28515] = t[28514] ^ n[28515];
assign t[28516] = t[28515] ^ n[28516];
assign t[28517] = t[28516] ^ n[28517];
assign t[28518] = t[28517] ^ n[28518];
assign t[28519] = t[28518] ^ n[28519];
assign t[28520] = t[28519] ^ n[28520];
assign t[28521] = t[28520] ^ n[28521];
assign t[28522] = t[28521] ^ n[28522];
assign t[28523] = t[28522] ^ n[28523];
assign t[28524] = t[28523] ^ n[28524];
assign t[28525] = t[28524] ^ n[28525];
assign t[28526] = t[28525] ^ n[28526];
assign t[28527] = t[28526] ^ n[28527];
assign t[28528] = t[28527] ^ n[28528];
assign t[28529] = t[28528] ^ n[28529];
assign t[28530] = t[28529] ^ n[28530];
assign t[28531] = t[28530] ^ n[28531];
assign t[28532] = t[28531] ^ n[28532];
assign t[28533] = t[28532] ^ n[28533];
assign t[28534] = t[28533] ^ n[28534];
assign t[28535] = t[28534] ^ n[28535];
assign t[28536] = t[28535] ^ n[28536];
assign t[28537] = t[28536] ^ n[28537];
assign t[28538] = t[28537] ^ n[28538];
assign t[28539] = t[28538] ^ n[28539];
assign t[28540] = t[28539] ^ n[28540];
assign t[28541] = t[28540] ^ n[28541];
assign t[28542] = t[28541] ^ n[28542];
assign t[28543] = t[28542] ^ n[28543];
assign t[28544] = t[28543] ^ n[28544];
assign t[28545] = t[28544] ^ n[28545];
assign t[28546] = t[28545] ^ n[28546];
assign t[28547] = t[28546] ^ n[28547];
assign t[28548] = t[28547] ^ n[28548];
assign t[28549] = t[28548] ^ n[28549];
assign t[28550] = t[28549] ^ n[28550];
assign t[28551] = t[28550] ^ n[28551];
assign t[28552] = t[28551] ^ n[28552];
assign t[28553] = t[28552] ^ n[28553];
assign t[28554] = t[28553] ^ n[28554];
assign t[28555] = t[28554] ^ n[28555];
assign t[28556] = t[28555] ^ n[28556];
assign t[28557] = t[28556] ^ n[28557];
assign t[28558] = t[28557] ^ n[28558];
assign t[28559] = t[28558] ^ n[28559];
assign t[28560] = t[28559] ^ n[28560];
assign t[28561] = t[28560] ^ n[28561];
assign t[28562] = t[28561] ^ n[28562];
assign t[28563] = t[28562] ^ n[28563];
assign t[28564] = t[28563] ^ n[28564];
assign t[28565] = t[28564] ^ n[28565];
assign t[28566] = t[28565] ^ n[28566];
assign t[28567] = t[28566] ^ n[28567];
assign t[28568] = t[28567] ^ n[28568];
assign t[28569] = t[28568] ^ n[28569];
assign t[28570] = t[28569] ^ n[28570];
assign t[28571] = t[28570] ^ n[28571];
assign t[28572] = t[28571] ^ n[28572];
assign t[28573] = t[28572] ^ n[28573];
assign t[28574] = t[28573] ^ n[28574];
assign t[28575] = t[28574] ^ n[28575];
assign t[28576] = t[28575] ^ n[28576];
assign t[28577] = t[28576] ^ n[28577];
assign t[28578] = t[28577] ^ n[28578];
assign t[28579] = t[28578] ^ n[28579];
assign t[28580] = t[28579] ^ n[28580];
assign t[28581] = t[28580] ^ n[28581];
assign t[28582] = t[28581] ^ n[28582];
assign t[28583] = t[28582] ^ n[28583];
assign t[28584] = t[28583] ^ n[28584];
assign t[28585] = t[28584] ^ n[28585];
assign t[28586] = t[28585] ^ n[28586];
assign t[28587] = t[28586] ^ n[28587];
assign t[28588] = t[28587] ^ n[28588];
assign t[28589] = t[28588] ^ n[28589];
assign t[28590] = t[28589] ^ n[28590];
assign t[28591] = t[28590] ^ n[28591];
assign t[28592] = t[28591] ^ n[28592];
assign t[28593] = t[28592] ^ n[28593];
assign t[28594] = t[28593] ^ n[28594];
assign t[28595] = t[28594] ^ n[28595];
assign t[28596] = t[28595] ^ n[28596];
assign t[28597] = t[28596] ^ n[28597];
assign t[28598] = t[28597] ^ n[28598];
assign t[28599] = t[28598] ^ n[28599];
assign t[28600] = t[28599] ^ n[28600];
assign t[28601] = t[28600] ^ n[28601];
assign t[28602] = t[28601] ^ n[28602];
assign t[28603] = t[28602] ^ n[28603];
assign t[28604] = t[28603] ^ n[28604];
assign t[28605] = t[28604] ^ n[28605];
assign t[28606] = t[28605] ^ n[28606];
assign t[28607] = t[28606] ^ n[28607];
assign t[28608] = t[28607] ^ n[28608];
assign t[28609] = t[28608] ^ n[28609];
assign t[28610] = t[28609] ^ n[28610];
assign t[28611] = t[28610] ^ n[28611];
assign t[28612] = t[28611] ^ n[28612];
assign t[28613] = t[28612] ^ n[28613];
assign t[28614] = t[28613] ^ n[28614];
assign t[28615] = t[28614] ^ n[28615];
assign t[28616] = t[28615] ^ n[28616];
assign t[28617] = t[28616] ^ n[28617];
assign t[28618] = t[28617] ^ n[28618];
assign t[28619] = t[28618] ^ n[28619];
assign t[28620] = t[28619] ^ n[28620];
assign t[28621] = t[28620] ^ n[28621];
assign t[28622] = t[28621] ^ n[28622];
assign t[28623] = t[28622] ^ n[28623];
assign t[28624] = t[28623] ^ n[28624];
assign t[28625] = t[28624] ^ n[28625];
assign t[28626] = t[28625] ^ n[28626];
assign t[28627] = t[28626] ^ n[28627];
assign t[28628] = t[28627] ^ n[28628];
assign t[28629] = t[28628] ^ n[28629];
assign t[28630] = t[28629] ^ n[28630];
assign t[28631] = t[28630] ^ n[28631];
assign t[28632] = t[28631] ^ n[28632];
assign t[28633] = t[28632] ^ n[28633];
assign t[28634] = t[28633] ^ n[28634];
assign t[28635] = t[28634] ^ n[28635];
assign t[28636] = t[28635] ^ n[28636];
assign t[28637] = t[28636] ^ n[28637];
assign t[28638] = t[28637] ^ n[28638];
assign t[28639] = t[28638] ^ n[28639];
assign t[28640] = t[28639] ^ n[28640];
assign t[28641] = t[28640] ^ n[28641];
assign t[28642] = t[28641] ^ n[28642];
assign t[28643] = t[28642] ^ n[28643];
assign t[28644] = t[28643] ^ n[28644];
assign t[28645] = t[28644] ^ n[28645];
assign t[28646] = t[28645] ^ n[28646];
assign t[28647] = t[28646] ^ n[28647];
assign t[28648] = t[28647] ^ n[28648];
assign t[28649] = t[28648] ^ n[28649];
assign t[28650] = t[28649] ^ n[28650];
assign t[28651] = t[28650] ^ n[28651];
assign t[28652] = t[28651] ^ n[28652];
assign t[28653] = t[28652] ^ n[28653];
assign t[28654] = t[28653] ^ n[28654];
assign t[28655] = t[28654] ^ n[28655];
assign t[28656] = t[28655] ^ n[28656];
assign t[28657] = t[28656] ^ n[28657];
assign t[28658] = t[28657] ^ n[28658];
assign t[28659] = t[28658] ^ n[28659];
assign t[28660] = t[28659] ^ n[28660];
assign t[28661] = t[28660] ^ n[28661];
assign t[28662] = t[28661] ^ n[28662];
assign t[28663] = t[28662] ^ n[28663];
assign t[28664] = t[28663] ^ n[28664];
assign t[28665] = t[28664] ^ n[28665];
assign t[28666] = t[28665] ^ n[28666];
assign t[28667] = t[28666] ^ n[28667];
assign t[28668] = t[28667] ^ n[28668];
assign t[28669] = t[28668] ^ n[28669];
assign t[28670] = t[28669] ^ n[28670];
assign t[28671] = t[28670] ^ n[28671];
assign t[28672] = t[28671] ^ n[28672];
assign t[28673] = t[28672] ^ n[28673];
assign t[28674] = t[28673] ^ n[28674];
assign t[28675] = t[28674] ^ n[28675];
assign t[28676] = t[28675] ^ n[28676];
assign t[28677] = t[28676] ^ n[28677];
assign t[28678] = t[28677] ^ n[28678];
assign t[28679] = t[28678] ^ n[28679];
assign t[28680] = t[28679] ^ n[28680];
assign t[28681] = t[28680] ^ n[28681];
assign t[28682] = t[28681] ^ n[28682];
assign t[28683] = t[28682] ^ n[28683];
assign t[28684] = t[28683] ^ n[28684];
assign t[28685] = t[28684] ^ n[28685];
assign t[28686] = t[28685] ^ n[28686];
assign t[28687] = t[28686] ^ n[28687];
assign t[28688] = t[28687] ^ n[28688];
assign t[28689] = t[28688] ^ n[28689];
assign t[28690] = t[28689] ^ n[28690];
assign t[28691] = t[28690] ^ n[28691];
assign t[28692] = t[28691] ^ n[28692];
assign t[28693] = t[28692] ^ n[28693];
assign t[28694] = t[28693] ^ n[28694];
assign t[28695] = t[28694] ^ n[28695];
assign t[28696] = t[28695] ^ n[28696];
assign t[28697] = t[28696] ^ n[28697];
assign t[28698] = t[28697] ^ n[28698];
assign t[28699] = t[28698] ^ n[28699];
assign t[28700] = t[28699] ^ n[28700];
assign t[28701] = t[28700] ^ n[28701];
assign t[28702] = t[28701] ^ n[28702];
assign t[28703] = t[28702] ^ n[28703];
assign t[28704] = t[28703] ^ n[28704];
assign t[28705] = t[28704] ^ n[28705];
assign t[28706] = t[28705] ^ n[28706];
assign t[28707] = t[28706] ^ n[28707];
assign t[28708] = t[28707] ^ n[28708];
assign t[28709] = t[28708] ^ n[28709];
assign t[28710] = t[28709] ^ n[28710];
assign t[28711] = t[28710] ^ n[28711];
assign t[28712] = t[28711] ^ n[28712];
assign t[28713] = t[28712] ^ n[28713];
assign t[28714] = t[28713] ^ n[28714];
assign t[28715] = t[28714] ^ n[28715];
assign t[28716] = t[28715] ^ n[28716];
assign t[28717] = t[28716] ^ n[28717];
assign t[28718] = t[28717] ^ n[28718];
assign t[28719] = t[28718] ^ n[28719];
assign t[28720] = t[28719] ^ n[28720];
assign t[28721] = t[28720] ^ n[28721];
assign t[28722] = t[28721] ^ n[28722];
assign t[28723] = t[28722] ^ n[28723];
assign t[28724] = t[28723] ^ n[28724];
assign t[28725] = t[28724] ^ n[28725];
assign t[28726] = t[28725] ^ n[28726];
assign t[28727] = t[28726] ^ n[28727];
assign t[28728] = t[28727] ^ n[28728];
assign t[28729] = t[28728] ^ n[28729];
assign t[28730] = t[28729] ^ n[28730];
assign t[28731] = t[28730] ^ n[28731];
assign t[28732] = t[28731] ^ n[28732];
assign t[28733] = t[28732] ^ n[28733];
assign t[28734] = t[28733] ^ n[28734];
assign t[28735] = t[28734] ^ n[28735];
assign t[28736] = t[28735] ^ n[28736];
assign t[28737] = t[28736] ^ n[28737];
assign t[28738] = t[28737] ^ n[28738];
assign t[28739] = t[28738] ^ n[28739];
assign t[28740] = t[28739] ^ n[28740];
assign t[28741] = t[28740] ^ n[28741];
assign t[28742] = t[28741] ^ n[28742];
assign t[28743] = t[28742] ^ n[28743];
assign t[28744] = t[28743] ^ n[28744];
assign t[28745] = t[28744] ^ n[28745];
assign t[28746] = t[28745] ^ n[28746];
assign t[28747] = t[28746] ^ n[28747];
assign t[28748] = t[28747] ^ n[28748];
assign t[28749] = t[28748] ^ n[28749];
assign t[28750] = t[28749] ^ n[28750];
assign t[28751] = t[28750] ^ n[28751];
assign t[28752] = t[28751] ^ n[28752];
assign t[28753] = t[28752] ^ n[28753];
assign t[28754] = t[28753] ^ n[28754];
assign t[28755] = t[28754] ^ n[28755];
assign t[28756] = t[28755] ^ n[28756];
assign t[28757] = t[28756] ^ n[28757];
assign t[28758] = t[28757] ^ n[28758];
assign t[28759] = t[28758] ^ n[28759];
assign t[28760] = t[28759] ^ n[28760];
assign t[28761] = t[28760] ^ n[28761];
assign t[28762] = t[28761] ^ n[28762];
assign t[28763] = t[28762] ^ n[28763];
assign t[28764] = t[28763] ^ n[28764];
assign t[28765] = t[28764] ^ n[28765];
assign t[28766] = t[28765] ^ n[28766];
assign t[28767] = t[28766] ^ n[28767];
assign t[28768] = t[28767] ^ n[28768];
assign t[28769] = t[28768] ^ n[28769];
assign t[28770] = t[28769] ^ n[28770];
assign t[28771] = t[28770] ^ n[28771];
assign t[28772] = t[28771] ^ n[28772];
assign t[28773] = t[28772] ^ n[28773];
assign t[28774] = t[28773] ^ n[28774];
assign t[28775] = t[28774] ^ n[28775];
assign t[28776] = t[28775] ^ n[28776];
assign t[28777] = t[28776] ^ n[28777];
assign t[28778] = t[28777] ^ n[28778];
assign t[28779] = t[28778] ^ n[28779];
assign t[28780] = t[28779] ^ n[28780];
assign t[28781] = t[28780] ^ n[28781];
assign t[28782] = t[28781] ^ n[28782];
assign t[28783] = t[28782] ^ n[28783];
assign t[28784] = t[28783] ^ n[28784];
assign t[28785] = t[28784] ^ n[28785];
assign t[28786] = t[28785] ^ n[28786];
assign t[28787] = t[28786] ^ n[28787];
assign t[28788] = t[28787] ^ n[28788];
assign t[28789] = t[28788] ^ n[28789];
assign t[28790] = t[28789] ^ n[28790];
assign t[28791] = t[28790] ^ n[28791];
assign t[28792] = t[28791] ^ n[28792];
assign t[28793] = t[28792] ^ n[28793];
assign t[28794] = t[28793] ^ n[28794];
assign t[28795] = t[28794] ^ n[28795];
assign t[28796] = t[28795] ^ n[28796];
assign t[28797] = t[28796] ^ n[28797];
assign t[28798] = t[28797] ^ n[28798];
assign t[28799] = t[28798] ^ n[28799];
assign t[28800] = t[28799] ^ n[28800];
assign t[28801] = t[28800] ^ n[28801];
assign t[28802] = t[28801] ^ n[28802];
assign t[28803] = t[28802] ^ n[28803];
assign t[28804] = t[28803] ^ n[28804];
assign t[28805] = t[28804] ^ n[28805];
assign t[28806] = t[28805] ^ n[28806];
assign t[28807] = t[28806] ^ n[28807];
assign t[28808] = t[28807] ^ n[28808];
assign t[28809] = t[28808] ^ n[28809];
assign t[28810] = t[28809] ^ n[28810];
assign t[28811] = t[28810] ^ n[28811];
assign t[28812] = t[28811] ^ n[28812];
assign t[28813] = t[28812] ^ n[28813];
assign t[28814] = t[28813] ^ n[28814];
assign t[28815] = t[28814] ^ n[28815];
assign t[28816] = t[28815] ^ n[28816];
assign t[28817] = t[28816] ^ n[28817];
assign t[28818] = t[28817] ^ n[28818];
assign t[28819] = t[28818] ^ n[28819];
assign t[28820] = t[28819] ^ n[28820];
assign t[28821] = t[28820] ^ n[28821];
assign t[28822] = t[28821] ^ n[28822];
assign t[28823] = t[28822] ^ n[28823];
assign t[28824] = t[28823] ^ n[28824];
assign t[28825] = t[28824] ^ n[28825];
assign t[28826] = t[28825] ^ n[28826];
assign t[28827] = t[28826] ^ n[28827];
assign t[28828] = t[28827] ^ n[28828];
assign t[28829] = t[28828] ^ n[28829];
assign t[28830] = t[28829] ^ n[28830];
assign t[28831] = t[28830] ^ n[28831];
assign t[28832] = t[28831] ^ n[28832];
assign t[28833] = t[28832] ^ n[28833];
assign t[28834] = t[28833] ^ n[28834];
assign t[28835] = t[28834] ^ n[28835];
assign t[28836] = t[28835] ^ n[28836];
assign t[28837] = t[28836] ^ n[28837];
assign t[28838] = t[28837] ^ n[28838];
assign t[28839] = t[28838] ^ n[28839];
assign t[28840] = t[28839] ^ n[28840];
assign t[28841] = t[28840] ^ n[28841];
assign t[28842] = t[28841] ^ n[28842];
assign t[28843] = t[28842] ^ n[28843];
assign t[28844] = t[28843] ^ n[28844];
assign t[28845] = t[28844] ^ n[28845];
assign t[28846] = t[28845] ^ n[28846];
assign t[28847] = t[28846] ^ n[28847];
assign t[28848] = t[28847] ^ n[28848];
assign t[28849] = t[28848] ^ n[28849];
assign t[28850] = t[28849] ^ n[28850];
assign t[28851] = t[28850] ^ n[28851];
assign t[28852] = t[28851] ^ n[28852];
assign t[28853] = t[28852] ^ n[28853];
assign t[28854] = t[28853] ^ n[28854];
assign t[28855] = t[28854] ^ n[28855];
assign t[28856] = t[28855] ^ n[28856];
assign t[28857] = t[28856] ^ n[28857];
assign t[28858] = t[28857] ^ n[28858];
assign t[28859] = t[28858] ^ n[28859];
assign t[28860] = t[28859] ^ n[28860];
assign t[28861] = t[28860] ^ n[28861];
assign t[28862] = t[28861] ^ n[28862];
assign t[28863] = t[28862] ^ n[28863];
assign t[28864] = t[28863] ^ n[28864];
assign t[28865] = t[28864] ^ n[28865];
assign t[28866] = t[28865] ^ n[28866];
assign t[28867] = t[28866] ^ n[28867];
assign t[28868] = t[28867] ^ n[28868];
assign t[28869] = t[28868] ^ n[28869];
assign t[28870] = t[28869] ^ n[28870];
assign t[28871] = t[28870] ^ n[28871];
assign t[28872] = t[28871] ^ n[28872];
assign t[28873] = t[28872] ^ n[28873];
assign t[28874] = t[28873] ^ n[28874];
assign t[28875] = t[28874] ^ n[28875];
assign t[28876] = t[28875] ^ n[28876];
assign t[28877] = t[28876] ^ n[28877];
assign t[28878] = t[28877] ^ n[28878];
assign t[28879] = t[28878] ^ n[28879];
assign t[28880] = t[28879] ^ n[28880];
assign t[28881] = t[28880] ^ n[28881];
assign t[28882] = t[28881] ^ n[28882];
assign t[28883] = t[28882] ^ n[28883];
assign t[28884] = t[28883] ^ n[28884];
assign t[28885] = t[28884] ^ n[28885];
assign t[28886] = t[28885] ^ n[28886];
assign t[28887] = t[28886] ^ n[28887];
assign t[28888] = t[28887] ^ n[28888];
assign t[28889] = t[28888] ^ n[28889];
assign t[28890] = t[28889] ^ n[28890];
assign t[28891] = t[28890] ^ n[28891];
assign t[28892] = t[28891] ^ n[28892];
assign t[28893] = t[28892] ^ n[28893];
assign t[28894] = t[28893] ^ n[28894];
assign t[28895] = t[28894] ^ n[28895];
assign t[28896] = t[28895] ^ n[28896];
assign t[28897] = t[28896] ^ n[28897];
assign t[28898] = t[28897] ^ n[28898];
assign t[28899] = t[28898] ^ n[28899];
assign t[28900] = t[28899] ^ n[28900];
assign t[28901] = t[28900] ^ n[28901];
assign t[28902] = t[28901] ^ n[28902];
assign t[28903] = t[28902] ^ n[28903];
assign t[28904] = t[28903] ^ n[28904];
assign t[28905] = t[28904] ^ n[28905];
assign t[28906] = t[28905] ^ n[28906];
assign t[28907] = t[28906] ^ n[28907];
assign t[28908] = t[28907] ^ n[28908];
assign t[28909] = t[28908] ^ n[28909];
assign t[28910] = t[28909] ^ n[28910];
assign t[28911] = t[28910] ^ n[28911];
assign t[28912] = t[28911] ^ n[28912];
assign t[28913] = t[28912] ^ n[28913];
assign t[28914] = t[28913] ^ n[28914];
assign t[28915] = t[28914] ^ n[28915];
assign t[28916] = t[28915] ^ n[28916];
assign t[28917] = t[28916] ^ n[28917];
assign t[28918] = t[28917] ^ n[28918];
assign t[28919] = t[28918] ^ n[28919];
assign t[28920] = t[28919] ^ n[28920];
assign t[28921] = t[28920] ^ n[28921];
assign t[28922] = t[28921] ^ n[28922];
assign t[28923] = t[28922] ^ n[28923];
assign t[28924] = t[28923] ^ n[28924];
assign t[28925] = t[28924] ^ n[28925];
assign t[28926] = t[28925] ^ n[28926];
assign t[28927] = t[28926] ^ n[28927];
assign t[28928] = t[28927] ^ n[28928];
assign t[28929] = t[28928] ^ n[28929];
assign t[28930] = t[28929] ^ n[28930];
assign t[28931] = t[28930] ^ n[28931];
assign t[28932] = t[28931] ^ n[28932];
assign t[28933] = t[28932] ^ n[28933];
assign t[28934] = t[28933] ^ n[28934];
assign t[28935] = t[28934] ^ n[28935];
assign t[28936] = t[28935] ^ n[28936];
assign t[28937] = t[28936] ^ n[28937];
assign t[28938] = t[28937] ^ n[28938];
assign t[28939] = t[28938] ^ n[28939];
assign t[28940] = t[28939] ^ n[28940];
assign t[28941] = t[28940] ^ n[28941];
assign t[28942] = t[28941] ^ n[28942];
assign t[28943] = t[28942] ^ n[28943];
assign t[28944] = t[28943] ^ n[28944];
assign t[28945] = t[28944] ^ n[28945];
assign t[28946] = t[28945] ^ n[28946];
assign t[28947] = t[28946] ^ n[28947];
assign t[28948] = t[28947] ^ n[28948];
assign t[28949] = t[28948] ^ n[28949];
assign t[28950] = t[28949] ^ n[28950];
assign t[28951] = t[28950] ^ n[28951];
assign t[28952] = t[28951] ^ n[28952];
assign t[28953] = t[28952] ^ n[28953];
assign t[28954] = t[28953] ^ n[28954];
assign t[28955] = t[28954] ^ n[28955];
assign t[28956] = t[28955] ^ n[28956];
assign t[28957] = t[28956] ^ n[28957];
assign t[28958] = t[28957] ^ n[28958];
assign t[28959] = t[28958] ^ n[28959];
assign t[28960] = t[28959] ^ n[28960];
assign t[28961] = t[28960] ^ n[28961];
assign t[28962] = t[28961] ^ n[28962];
assign t[28963] = t[28962] ^ n[28963];
assign t[28964] = t[28963] ^ n[28964];
assign t[28965] = t[28964] ^ n[28965];
assign t[28966] = t[28965] ^ n[28966];
assign t[28967] = t[28966] ^ n[28967];
assign t[28968] = t[28967] ^ n[28968];
assign t[28969] = t[28968] ^ n[28969];
assign t[28970] = t[28969] ^ n[28970];
assign t[28971] = t[28970] ^ n[28971];
assign t[28972] = t[28971] ^ n[28972];
assign t[28973] = t[28972] ^ n[28973];
assign t[28974] = t[28973] ^ n[28974];
assign t[28975] = t[28974] ^ n[28975];
assign t[28976] = t[28975] ^ n[28976];
assign t[28977] = t[28976] ^ n[28977];
assign t[28978] = t[28977] ^ n[28978];
assign t[28979] = t[28978] ^ n[28979];
assign t[28980] = t[28979] ^ n[28980];
assign t[28981] = t[28980] ^ n[28981];
assign t[28982] = t[28981] ^ n[28982];
assign t[28983] = t[28982] ^ n[28983];
assign t[28984] = t[28983] ^ n[28984];
assign t[28985] = t[28984] ^ n[28985];
assign t[28986] = t[28985] ^ n[28986];
assign t[28987] = t[28986] ^ n[28987];
assign t[28988] = t[28987] ^ n[28988];
assign t[28989] = t[28988] ^ n[28989];
assign t[28990] = t[28989] ^ n[28990];
assign t[28991] = t[28990] ^ n[28991];
assign t[28992] = t[28991] ^ n[28992];
assign t[28993] = t[28992] ^ n[28993];
assign t[28994] = t[28993] ^ n[28994];
assign t[28995] = t[28994] ^ n[28995];
assign t[28996] = t[28995] ^ n[28996];
assign t[28997] = t[28996] ^ n[28997];
assign t[28998] = t[28997] ^ n[28998];
assign t[28999] = t[28998] ^ n[28999];
assign t[29000] = t[28999] ^ n[29000];
assign t[29001] = t[29000] ^ n[29001];
assign t[29002] = t[29001] ^ n[29002];
assign t[29003] = t[29002] ^ n[29003];
assign t[29004] = t[29003] ^ n[29004];
assign t[29005] = t[29004] ^ n[29005];
assign t[29006] = t[29005] ^ n[29006];
assign t[29007] = t[29006] ^ n[29007];
assign t[29008] = t[29007] ^ n[29008];
assign t[29009] = t[29008] ^ n[29009];
assign t[29010] = t[29009] ^ n[29010];
assign t[29011] = t[29010] ^ n[29011];
assign t[29012] = t[29011] ^ n[29012];
assign t[29013] = t[29012] ^ n[29013];
assign t[29014] = t[29013] ^ n[29014];
assign t[29015] = t[29014] ^ n[29015];
assign t[29016] = t[29015] ^ n[29016];
assign t[29017] = t[29016] ^ n[29017];
assign t[29018] = t[29017] ^ n[29018];
assign t[29019] = t[29018] ^ n[29019];
assign t[29020] = t[29019] ^ n[29020];
assign t[29021] = t[29020] ^ n[29021];
assign t[29022] = t[29021] ^ n[29022];
assign t[29023] = t[29022] ^ n[29023];
assign t[29024] = t[29023] ^ n[29024];
assign t[29025] = t[29024] ^ n[29025];
assign t[29026] = t[29025] ^ n[29026];
assign t[29027] = t[29026] ^ n[29027];
assign t[29028] = t[29027] ^ n[29028];
assign t[29029] = t[29028] ^ n[29029];
assign t[29030] = t[29029] ^ n[29030];
assign t[29031] = t[29030] ^ n[29031];
assign t[29032] = t[29031] ^ n[29032];
assign t[29033] = t[29032] ^ n[29033];
assign t[29034] = t[29033] ^ n[29034];
assign t[29035] = t[29034] ^ n[29035];
assign t[29036] = t[29035] ^ n[29036];
assign t[29037] = t[29036] ^ n[29037];
assign t[29038] = t[29037] ^ n[29038];
assign t[29039] = t[29038] ^ n[29039];
assign t[29040] = t[29039] ^ n[29040];
assign t[29041] = t[29040] ^ n[29041];
assign t[29042] = t[29041] ^ n[29042];
assign t[29043] = t[29042] ^ n[29043];
assign t[29044] = t[29043] ^ n[29044];
assign t[29045] = t[29044] ^ n[29045];
assign t[29046] = t[29045] ^ n[29046];
assign t[29047] = t[29046] ^ n[29047];
assign t[29048] = t[29047] ^ n[29048];
assign t[29049] = t[29048] ^ n[29049];
assign t[29050] = t[29049] ^ n[29050];
assign t[29051] = t[29050] ^ n[29051];
assign t[29052] = t[29051] ^ n[29052];
assign t[29053] = t[29052] ^ n[29053];
assign t[29054] = t[29053] ^ n[29054];
assign t[29055] = t[29054] ^ n[29055];
assign t[29056] = t[29055] ^ n[29056];
assign t[29057] = t[29056] ^ n[29057];
assign t[29058] = t[29057] ^ n[29058];
assign t[29059] = t[29058] ^ n[29059];
assign t[29060] = t[29059] ^ n[29060];
assign t[29061] = t[29060] ^ n[29061];
assign t[29062] = t[29061] ^ n[29062];
assign t[29063] = t[29062] ^ n[29063];
assign t[29064] = t[29063] ^ n[29064];
assign t[29065] = t[29064] ^ n[29065];
assign t[29066] = t[29065] ^ n[29066];
assign t[29067] = t[29066] ^ n[29067];
assign t[29068] = t[29067] ^ n[29068];
assign t[29069] = t[29068] ^ n[29069];
assign t[29070] = t[29069] ^ n[29070];
assign t[29071] = t[29070] ^ n[29071];
assign t[29072] = t[29071] ^ n[29072];
assign t[29073] = t[29072] ^ n[29073];
assign t[29074] = t[29073] ^ n[29074];
assign t[29075] = t[29074] ^ n[29075];
assign t[29076] = t[29075] ^ n[29076];
assign t[29077] = t[29076] ^ n[29077];
assign t[29078] = t[29077] ^ n[29078];
assign t[29079] = t[29078] ^ n[29079];
assign t[29080] = t[29079] ^ n[29080];
assign t[29081] = t[29080] ^ n[29081];
assign t[29082] = t[29081] ^ n[29082];
assign t[29083] = t[29082] ^ n[29083];
assign t[29084] = t[29083] ^ n[29084];
assign t[29085] = t[29084] ^ n[29085];
assign t[29086] = t[29085] ^ n[29086];
assign t[29087] = t[29086] ^ n[29087];
assign t[29088] = t[29087] ^ n[29088];
assign t[29089] = t[29088] ^ n[29089];
assign t[29090] = t[29089] ^ n[29090];
assign t[29091] = t[29090] ^ n[29091];
assign t[29092] = t[29091] ^ n[29092];
assign t[29093] = t[29092] ^ n[29093];
assign t[29094] = t[29093] ^ n[29094];
assign t[29095] = t[29094] ^ n[29095];
assign t[29096] = t[29095] ^ n[29096];
assign t[29097] = t[29096] ^ n[29097];
assign t[29098] = t[29097] ^ n[29098];
assign t[29099] = t[29098] ^ n[29099];
assign t[29100] = t[29099] ^ n[29100];
assign t[29101] = t[29100] ^ n[29101];
assign t[29102] = t[29101] ^ n[29102];
assign t[29103] = t[29102] ^ n[29103];
assign t[29104] = t[29103] ^ n[29104];
assign t[29105] = t[29104] ^ n[29105];
assign t[29106] = t[29105] ^ n[29106];
assign t[29107] = t[29106] ^ n[29107];
assign t[29108] = t[29107] ^ n[29108];
assign t[29109] = t[29108] ^ n[29109];
assign t[29110] = t[29109] ^ n[29110];
assign t[29111] = t[29110] ^ n[29111];
assign t[29112] = t[29111] ^ n[29112];
assign t[29113] = t[29112] ^ n[29113];
assign t[29114] = t[29113] ^ n[29114];
assign t[29115] = t[29114] ^ n[29115];
assign t[29116] = t[29115] ^ n[29116];
assign t[29117] = t[29116] ^ n[29117];
assign t[29118] = t[29117] ^ n[29118];
assign t[29119] = t[29118] ^ n[29119];
assign t[29120] = t[29119] ^ n[29120];
assign t[29121] = t[29120] ^ n[29121];
assign t[29122] = t[29121] ^ n[29122];
assign t[29123] = t[29122] ^ n[29123];
assign t[29124] = t[29123] ^ n[29124];
assign t[29125] = t[29124] ^ n[29125];
assign t[29126] = t[29125] ^ n[29126];
assign t[29127] = t[29126] ^ n[29127];
assign t[29128] = t[29127] ^ n[29128];
assign t[29129] = t[29128] ^ n[29129];
assign t[29130] = t[29129] ^ n[29130];
assign t[29131] = t[29130] ^ n[29131];
assign t[29132] = t[29131] ^ n[29132];
assign t[29133] = t[29132] ^ n[29133];
assign t[29134] = t[29133] ^ n[29134];
assign t[29135] = t[29134] ^ n[29135];
assign t[29136] = t[29135] ^ n[29136];
assign t[29137] = t[29136] ^ n[29137];
assign t[29138] = t[29137] ^ n[29138];
assign t[29139] = t[29138] ^ n[29139];
assign t[29140] = t[29139] ^ n[29140];
assign t[29141] = t[29140] ^ n[29141];
assign t[29142] = t[29141] ^ n[29142];
assign t[29143] = t[29142] ^ n[29143];
assign t[29144] = t[29143] ^ n[29144];
assign t[29145] = t[29144] ^ n[29145];
assign t[29146] = t[29145] ^ n[29146];
assign t[29147] = t[29146] ^ n[29147];
assign t[29148] = t[29147] ^ n[29148];
assign t[29149] = t[29148] ^ n[29149];
assign t[29150] = t[29149] ^ n[29150];
assign t[29151] = t[29150] ^ n[29151];
assign t[29152] = t[29151] ^ n[29152];
assign t[29153] = t[29152] ^ n[29153];
assign t[29154] = t[29153] ^ n[29154];
assign t[29155] = t[29154] ^ n[29155];
assign t[29156] = t[29155] ^ n[29156];
assign t[29157] = t[29156] ^ n[29157];
assign t[29158] = t[29157] ^ n[29158];
assign t[29159] = t[29158] ^ n[29159];
assign t[29160] = t[29159] ^ n[29160];
assign t[29161] = t[29160] ^ n[29161];
assign t[29162] = t[29161] ^ n[29162];
assign t[29163] = t[29162] ^ n[29163];
assign t[29164] = t[29163] ^ n[29164];
assign t[29165] = t[29164] ^ n[29165];
assign t[29166] = t[29165] ^ n[29166];
assign t[29167] = t[29166] ^ n[29167];
assign t[29168] = t[29167] ^ n[29168];
assign t[29169] = t[29168] ^ n[29169];
assign t[29170] = t[29169] ^ n[29170];
assign t[29171] = t[29170] ^ n[29171];
assign t[29172] = t[29171] ^ n[29172];
assign t[29173] = t[29172] ^ n[29173];
assign t[29174] = t[29173] ^ n[29174];
assign t[29175] = t[29174] ^ n[29175];
assign t[29176] = t[29175] ^ n[29176];
assign t[29177] = t[29176] ^ n[29177];
assign t[29178] = t[29177] ^ n[29178];
assign t[29179] = t[29178] ^ n[29179];
assign t[29180] = t[29179] ^ n[29180];
assign t[29181] = t[29180] ^ n[29181];
assign t[29182] = t[29181] ^ n[29182];
assign t[29183] = t[29182] ^ n[29183];
assign t[29184] = t[29183] ^ n[29184];
assign t[29185] = t[29184] ^ n[29185];
assign t[29186] = t[29185] ^ n[29186];
assign t[29187] = t[29186] ^ n[29187];
assign t[29188] = t[29187] ^ n[29188];
assign t[29189] = t[29188] ^ n[29189];
assign t[29190] = t[29189] ^ n[29190];
assign t[29191] = t[29190] ^ n[29191];
assign t[29192] = t[29191] ^ n[29192];
assign t[29193] = t[29192] ^ n[29193];
assign t[29194] = t[29193] ^ n[29194];
assign t[29195] = t[29194] ^ n[29195];
assign t[29196] = t[29195] ^ n[29196];
assign t[29197] = t[29196] ^ n[29197];
assign t[29198] = t[29197] ^ n[29198];
assign t[29199] = t[29198] ^ n[29199];
assign t[29200] = t[29199] ^ n[29200];
assign t[29201] = t[29200] ^ n[29201];
assign t[29202] = t[29201] ^ n[29202];
assign t[29203] = t[29202] ^ n[29203];
assign t[29204] = t[29203] ^ n[29204];
assign t[29205] = t[29204] ^ n[29205];
assign t[29206] = t[29205] ^ n[29206];
assign t[29207] = t[29206] ^ n[29207];
assign t[29208] = t[29207] ^ n[29208];
assign t[29209] = t[29208] ^ n[29209];
assign t[29210] = t[29209] ^ n[29210];
assign t[29211] = t[29210] ^ n[29211];
assign t[29212] = t[29211] ^ n[29212];
assign t[29213] = t[29212] ^ n[29213];
assign t[29214] = t[29213] ^ n[29214];
assign t[29215] = t[29214] ^ n[29215];
assign t[29216] = t[29215] ^ n[29216];
assign t[29217] = t[29216] ^ n[29217];
assign t[29218] = t[29217] ^ n[29218];
assign t[29219] = t[29218] ^ n[29219];
assign t[29220] = t[29219] ^ n[29220];
assign t[29221] = t[29220] ^ n[29221];
assign t[29222] = t[29221] ^ n[29222];
assign t[29223] = t[29222] ^ n[29223];
assign t[29224] = t[29223] ^ n[29224];
assign t[29225] = t[29224] ^ n[29225];
assign t[29226] = t[29225] ^ n[29226];
assign t[29227] = t[29226] ^ n[29227];
assign t[29228] = t[29227] ^ n[29228];
assign t[29229] = t[29228] ^ n[29229];
assign t[29230] = t[29229] ^ n[29230];
assign t[29231] = t[29230] ^ n[29231];
assign t[29232] = t[29231] ^ n[29232];
assign t[29233] = t[29232] ^ n[29233];
assign t[29234] = t[29233] ^ n[29234];
assign t[29235] = t[29234] ^ n[29235];
assign t[29236] = t[29235] ^ n[29236];
assign t[29237] = t[29236] ^ n[29237];
assign t[29238] = t[29237] ^ n[29238];
assign t[29239] = t[29238] ^ n[29239];
assign t[29240] = t[29239] ^ n[29240];
assign t[29241] = t[29240] ^ n[29241];
assign t[29242] = t[29241] ^ n[29242];
assign t[29243] = t[29242] ^ n[29243];
assign t[29244] = t[29243] ^ n[29244];
assign t[29245] = t[29244] ^ n[29245];
assign t[29246] = t[29245] ^ n[29246];
assign t[29247] = t[29246] ^ n[29247];
assign t[29248] = t[29247] ^ n[29248];
assign t[29249] = t[29248] ^ n[29249];
assign t[29250] = t[29249] ^ n[29250];
assign t[29251] = t[29250] ^ n[29251];
assign t[29252] = t[29251] ^ n[29252];
assign t[29253] = t[29252] ^ n[29253];
assign t[29254] = t[29253] ^ n[29254];
assign t[29255] = t[29254] ^ n[29255];
assign t[29256] = t[29255] ^ n[29256];
assign t[29257] = t[29256] ^ n[29257];
assign t[29258] = t[29257] ^ n[29258];
assign t[29259] = t[29258] ^ n[29259];
assign t[29260] = t[29259] ^ n[29260];
assign t[29261] = t[29260] ^ n[29261];
assign t[29262] = t[29261] ^ n[29262];
assign t[29263] = t[29262] ^ n[29263];
assign t[29264] = t[29263] ^ n[29264];
assign t[29265] = t[29264] ^ n[29265];
assign t[29266] = t[29265] ^ n[29266];
assign t[29267] = t[29266] ^ n[29267];
assign t[29268] = t[29267] ^ n[29268];
assign t[29269] = t[29268] ^ n[29269];
assign t[29270] = t[29269] ^ n[29270];
assign t[29271] = t[29270] ^ n[29271];
assign t[29272] = t[29271] ^ n[29272];
assign t[29273] = t[29272] ^ n[29273];
assign t[29274] = t[29273] ^ n[29274];
assign t[29275] = t[29274] ^ n[29275];
assign t[29276] = t[29275] ^ n[29276];
assign t[29277] = t[29276] ^ n[29277];
assign t[29278] = t[29277] ^ n[29278];
assign t[29279] = t[29278] ^ n[29279];
assign t[29280] = t[29279] ^ n[29280];
assign t[29281] = t[29280] ^ n[29281];
assign t[29282] = t[29281] ^ n[29282];
assign t[29283] = t[29282] ^ n[29283];
assign t[29284] = t[29283] ^ n[29284];
assign t[29285] = t[29284] ^ n[29285];
assign t[29286] = t[29285] ^ n[29286];
assign t[29287] = t[29286] ^ n[29287];
assign t[29288] = t[29287] ^ n[29288];
assign t[29289] = t[29288] ^ n[29289];
assign t[29290] = t[29289] ^ n[29290];
assign t[29291] = t[29290] ^ n[29291];
assign t[29292] = t[29291] ^ n[29292];
assign t[29293] = t[29292] ^ n[29293];
assign t[29294] = t[29293] ^ n[29294];
assign t[29295] = t[29294] ^ n[29295];
assign t[29296] = t[29295] ^ n[29296];
assign t[29297] = t[29296] ^ n[29297];
assign t[29298] = t[29297] ^ n[29298];
assign t[29299] = t[29298] ^ n[29299];
assign t[29300] = t[29299] ^ n[29300];
assign t[29301] = t[29300] ^ n[29301];
assign t[29302] = t[29301] ^ n[29302];
assign t[29303] = t[29302] ^ n[29303];
assign t[29304] = t[29303] ^ n[29304];
assign t[29305] = t[29304] ^ n[29305];
assign t[29306] = t[29305] ^ n[29306];
assign t[29307] = t[29306] ^ n[29307];
assign t[29308] = t[29307] ^ n[29308];
assign t[29309] = t[29308] ^ n[29309];
assign t[29310] = t[29309] ^ n[29310];
assign t[29311] = t[29310] ^ n[29311];
assign t[29312] = t[29311] ^ n[29312];
assign t[29313] = t[29312] ^ n[29313];
assign t[29314] = t[29313] ^ n[29314];
assign t[29315] = t[29314] ^ n[29315];
assign t[29316] = t[29315] ^ n[29316];
assign t[29317] = t[29316] ^ n[29317];
assign t[29318] = t[29317] ^ n[29318];
assign t[29319] = t[29318] ^ n[29319];
assign t[29320] = t[29319] ^ n[29320];
assign t[29321] = t[29320] ^ n[29321];
assign t[29322] = t[29321] ^ n[29322];
assign t[29323] = t[29322] ^ n[29323];
assign t[29324] = t[29323] ^ n[29324];
assign t[29325] = t[29324] ^ n[29325];
assign t[29326] = t[29325] ^ n[29326];
assign t[29327] = t[29326] ^ n[29327];
assign t[29328] = t[29327] ^ n[29328];
assign t[29329] = t[29328] ^ n[29329];
assign t[29330] = t[29329] ^ n[29330];
assign t[29331] = t[29330] ^ n[29331];
assign t[29332] = t[29331] ^ n[29332];
assign t[29333] = t[29332] ^ n[29333];
assign t[29334] = t[29333] ^ n[29334];
assign t[29335] = t[29334] ^ n[29335];
assign t[29336] = t[29335] ^ n[29336];
assign t[29337] = t[29336] ^ n[29337];
assign t[29338] = t[29337] ^ n[29338];
assign t[29339] = t[29338] ^ n[29339];
assign t[29340] = t[29339] ^ n[29340];
assign t[29341] = t[29340] ^ n[29341];
assign t[29342] = t[29341] ^ n[29342];
assign t[29343] = t[29342] ^ n[29343];
assign t[29344] = t[29343] ^ n[29344];
assign t[29345] = t[29344] ^ n[29345];
assign t[29346] = t[29345] ^ n[29346];
assign t[29347] = t[29346] ^ n[29347];
assign t[29348] = t[29347] ^ n[29348];
assign t[29349] = t[29348] ^ n[29349];
assign t[29350] = t[29349] ^ n[29350];
assign t[29351] = t[29350] ^ n[29351];
assign t[29352] = t[29351] ^ n[29352];
assign t[29353] = t[29352] ^ n[29353];
assign t[29354] = t[29353] ^ n[29354];
assign t[29355] = t[29354] ^ n[29355];
assign t[29356] = t[29355] ^ n[29356];
assign t[29357] = t[29356] ^ n[29357];
assign t[29358] = t[29357] ^ n[29358];
assign t[29359] = t[29358] ^ n[29359];
assign t[29360] = t[29359] ^ n[29360];
assign t[29361] = t[29360] ^ n[29361];
assign t[29362] = t[29361] ^ n[29362];
assign t[29363] = t[29362] ^ n[29363];
assign t[29364] = t[29363] ^ n[29364];
assign t[29365] = t[29364] ^ n[29365];
assign t[29366] = t[29365] ^ n[29366];
assign t[29367] = t[29366] ^ n[29367];
assign t[29368] = t[29367] ^ n[29368];
assign t[29369] = t[29368] ^ n[29369];
assign t[29370] = t[29369] ^ n[29370];
assign t[29371] = t[29370] ^ n[29371];
assign t[29372] = t[29371] ^ n[29372];
assign t[29373] = t[29372] ^ n[29373];
assign t[29374] = t[29373] ^ n[29374];
assign t[29375] = t[29374] ^ n[29375];
assign t[29376] = t[29375] ^ n[29376];
assign t[29377] = t[29376] ^ n[29377];
assign t[29378] = t[29377] ^ n[29378];
assign t[29379] = t[29378] ^ n[29379];
assign t[29380] = t[29379] ^ n[29380];
assign t[29381] = t[29380] ^ n[29381];
assign t[29382] = t[29381] ^ n[29382];
assign t[29383] = t[29382] ^ n[29383];
assign t[29384] = t[29383] ^ n[29384];
assign t[29385] = t[29384] ^ n[29385];
assign t[29386] = t[29385] ^ n[29386];
assign t[29387] = t[29386] ^ n[29387];
assign t[29388] = t[29387] ^ n[29388];
assign t[29389] = t[29388] ^ n[29389];
assign t[29390] = t[29389] ^ n[29390];
assign t[29391] = t[29390] ^ n[29391];
assign t[29392] = t[29391] ^ n[29392];
assign t[29393] = t[29392] ^ n[29393];
assign t[29394] = t[29393] ^ n[29394];
assign t[29395] = t[29394] ^ n[29395];
assign t[29396] = t[29395] ^ n[29396];
assign t[29397] = t[29396] ^ n[29397];
assign t[29398] = t[29397] ^ n[29398];
assign t[29399] = t[29398] ^ n[29399];
assign t[29400] = t[29399] ^ n[29400];
assign t[29401] = t[29400] ^ n[29401];
assign t[29402] = t[29401] ^ n[29402];
assign t[29403] = t[29402] ^ n[29403];
assign t[29404] = t[29403] ^ n[29404];
assign t[29405] = t[29404] ^ n[29405];
assign t[29406] = t[29405] ^ n[29406];
assign t[29407] = t[29406] ^ n[29407];
assign t[29408] = t[29407] ^ n[29408];
assign t[29409] = t[29408] ^ n[29409];
assign t[29410] = t[29409] ^ n[29410];
assign t[29411] = t[29410] ^ n[29411];
assign t[29412] = t[29411] ^ n[29412];
assign t[29413] = t[29412] ^ n[29413];
assign t[29414] = t[29413] ^ n[29414];
assign t[29415] = t[29414] ^ n[29415];
assign t[29416] = t[29415] ^ n[29416];
assign t[29417] = t[29416] ^ n[29417];
assign t[29418] = t[29417] ^ n[29418];
assign t[29419] = t[29418] ^ n[29419];
assign t[29420] = t[29419] ^ n[29420];
assign t[29421] = t[29420] ^ n[29421];
assign t[29422] = t[29421] ^ n[29422];
assign t[29423] = t[29422] ^ n[29423];
assign t[29424] = t[29423] ^ n[29424];
assign t[29425] = t[29424] ^ n[29425];
assign t[29426] = t[29425] ^ n[29426];
assign t[29427] = t[29426] ^ n[29427];
assign t[29428] = t[29427] ^ n[29428];
assign t[29429] = t[29428] ^ n[29429];
assign t[29430] = t[29429] ^ n[29430];
assign t[29431] = t[29430] ^ n[29431];
assign t[29432] = t[29431] ^ n[29432];
assign t[29433] = t[29432] ^ n[29433];
assign t[29434] = t[29433] ^ n[29434];
assign t[29435] = t[29434] ^ n[29435];
assign t[29436] = t[29435] ^ n[29436];
assign t[29437] = t[29436] ^ n[29437];
assign t[29438] = t[29437] ^ n[29438];
assign t[29439] = t[29438] ^ n[29439];
assign t[29440] = t[29439] ^ n[29440];
assign t[29441] = t[29440] ^ n[29441];
assign t[29442] = t[29441] ^ n[29442];
assign t[29443] = t[29442] ^ n[29443];
assign t[29444] = t[29443] ^ n[29444];
assign t[29445] = t[29444] ^ n[29445];
assign t[29446] = t[29445] ^ n[29446];
assign t[29447] = t[29446] ^ n[29447];
assign t[29448] = t[29447] ^ n[29448];
assign t[29449] = t[29448] ^ n[29449];
assign t[29450] = t[29449] ^ n[29450];
assign t[29451] = t[29450] ^ n[29451];
assign t[29452] = t[29451] ^ n[29452];
assign t[29453] = t[29452] ^ n[29453];
assign t[29454] = t[29453] ^ n[29454];
assign t[29455] = t[29454] ^ n[29455];
assign t[29456] = t[29455] ^ n[29456];
assign t[29457] = t[29456] ^ n[29457];
assign t[29458] = t[29457] ^ n[29458];
assign t[29459] = t[29458] ^ n[29459];
assign t[29460] = t[29459] ^ n[29460];
assign t[29461] = t[29460] ^ n[29461];
assign t[29462] = t[29461] ^ n[29462];
assign t[29463] = t[29462] ^ n[29463];
assign t[29464] = t[29463] ^ n[29464];
assign t[29465] = t[29464] ^ n[29465];
assign t[29466] = t[29465] ^ n[29466];
assign t[29467] = t[29466] ^ n[29467];
assign t[29468] = t[29467] ^ n[29468];
assign t[29469] = t[29468] ^ n[29469];
assign t[29470] = t[29469] ^ n[29470];
assign t[29471] = t[29470] ^ n[29471];
assign t[29472] = t[29471] ^ n[29472];
assign t[29473] = t[29472] ^ n[29473];
assign t[29474] = t[29473] ^ n[29474];
assign t[29475] = t[29474] ^ n[29475];
assign t[29476] = t[29475] ^ n[29476];
assign t[29477] = t[29476] ^ n[29477];
assign t[29478] = t[29477] ^ n[29478];
assign t[29479] = t[29478] ^ n[29479];
assign t[29480] = t[29479] ^ n[29480];
assign t[29481] = t[29480] ^ n[29481];
assign t[29482] = t[29481] ^ n[29482];
assign t[29483] = t[29482] ^ n[29483];
assign t[29484] = t[29483] ^ n[29484];
assign t[29485] = t[29484] ^ n[29485];
assign t[29486] = t[29485] ^ n[29486];
assign t[29487] = t[29486] ^ n[29487];
assign t[29488] = t[29487] ^ n[29488];
assign t[29489] = t[29488] ^ n[29489];
assign t[29490] = t[29489] ^ n[29490];
assign t[29491] = t[29490] ^ n[29491];
assign t[29492] = t[29491] ^ n[29492];
assign t[29493] = t[29492] ^ n[29493];
assign t[29494] = t[29493] ^ n[29494];
assign t[29495] = t[29494] ^ n[29495];
assign t[29496] = t[29495] ^ n[29496];
assign t[29497] = t[29496] ^ n[29497];
assign t[29498] = t[29497] ^ n[29498];
assign t[29499] = t[29498] ^ n[29499];
assign t[29500] = t[29499] ^ n[29500];
assign t[29501] = t[29500] ^ n[29501];
assign t[29502] = t[29501] ^ n[29502];
assign t[29503] = t[29502] ^ n[29503];
assign t[29504] = t[29503] ^ n[29504];
assign t[29505] = t[29504] ^ n[29505];
assign t[29506] = t[29505] ^ n[29506];
assign t[29507] = t[29506] ^ n[29507];
assign t[29508] = t[29507] ^ n[29508];
assign t[29509] = t[29508] ^ n[29509];
assign t[29510] = t[29509] ^ n[29510];
assign t[29511] = t[29510] ^ n[29511];
assign t[29512] = t[29511] ^ n[29512];
assign t[29513] = t[29512] ^ n[29513];
assign t[29514] = t[29513] ^ n[29514];
assign t[29515] = t[29514] ^ n[29515];
assign t[29516] = t[29515] ^ n[29516];
assign t[29517] = t[29516] ^ n[29517];
assign t[29518] = t[29517] ^ n[29518];
assign t[29519] = t[29518] ^ n[29519];
assign t[29520] = t[29519] ^ n[29520];
assign t[29521] = t[29520] ^ n[29521];
assign t[29522] = t[29521] ^ n[29522];
assign t[29523] = t[29522] ^ n[29523];
assign t[29524] = t[29523] ^ n[29524];
assign t[29525] = t[29524] ^ n[29525];
assign t[29526] = t[29525] ^ n[29526];
assign t[29527] = t[29526] ^ n[29527];
assign t[29528] = t[29527] ^ n[29528];
assign t[29529] = t[29528] ^ n[29529];
assign t[29530] = t[29529] ^ n[29530];
assign t[29531] = t[29530] ^ n[29531];
assign t[29532] = t[29531] ^ n[29532];
assign t[29533] = t[29532] ^ n[29533];
assign t[29534] = t[29533] ^ n[29534];
assign t[29535] = t[29534] ^ n[29535];
assign t[29536] = t[29535] ^ n[29536];
assign t[29537] = t[29536] ^ n[29537];
assign t[29538] = t[29537] ^ n[29538];
assign t[29539] = t[29538] ^ n[29539];
assign t[29540] = t[29539] ^ n[29540];
assign t[29541] = t[29540] ^ n[29541];
assign t[29542] = t[29541] ^ n[29542];
assign t[29543] = t[29542] ^ n[29543];
assign t[29544] = t[29543] ^ n[29544];
assign t[29545] = t[29544] ^ n[29545];
assign t[29546] = t[29545] ^ n[29546];
assign t[29547] = t[29546] ^ n[29547];
assign t[29548] = t[29547] ^ n[29548];
assign t[29549] = t[29548] ^ n[29549];
assign t[29550] = t[29549] ^ n[29550];
assign t[29551] = t[29550] ^ n[29551];
assign t[29552] = t[29551] ^ n[29552];
assign t[29553] = t[29552] ^ n[29553];
assign t[29554] = t[29553] ^ n[29554];
assign t[29555] = t[29554] ^ n[29555];
assign t[29556] = t[29555] ^ n[29556];
assign t[29557] = t[29556] ^ n[29557];
assign t[29558] = t[29557] ^ n[29558];
assign t[29559] = t[29558] ^ n[29559];
assign t[29560] = t[29559] ^ n[29560];
assign t[29561] = t[29560] ^ n[29561];
assign t[29562] = t[29561] ^ n[29562];
assign t[29563] = t[29562] ^ n[29563];
assign t[29564] = t[29563] ^ n[29564];
assign t[29565] = t[29564] ^ n[29565];
assign t[29566] = t[29565] ^ n[29566];
assign t[29567] = t[29566] ^ n[29567];
assign t[29568] = t[29567] ^ n[29568];
assign t[29569] = t[29568] ^ n[29569];
assign t[29570] = t[29569] ^ n[29570];
assign t[29571] = t[29570] ^ n[29571];
assign t[29572] = t[29571] ^ n[29572];
assign t[29573] = t[29572] ^ n[29573];
assign t[29574] = t[29573] ^ n[29574];
assign t[29575] = t[29574] ^ n[29575];
assign t[29576] = t[29575] ^ n[29576];
assign t[29577] = t[29576] ^ n[29577];
assign t[29578] = t[29577] ^ n[29578];
assign t[29579] = t[29578] ^ n[29579];
assign t[29580] = t[29579] ^ n[29580];
assign t[29581] = t[29580] ^ n[29581];
assign t[29582] = t[29581] ^ n[29582];
assign t[29583] = t[29582] ^ n[29583];
assign t[29584] = t[29583] ^ n[29584];
assign t[29585] = t[29584] ^ n[29585];
assign t[29586] = t[29585] ^ n[29586];
assign t[29587] = t[29586] ^ n[29587];
assign t[29588] = t[29587] ^ n[29588];
assign t[29589] = t[29588] ^ n[29589];
assign t[29590] = t[29589] ^ n[29590];
assign t[29591] = t[29590] ^ n[29591];
assign t[29592] = t[29591] ^ n[29592];
assign t[29593] = t[29592] ^ n[29593];
assign t[29594] = t[29593] ^ n[29594];
assign t[29595] = t[29594] ^ n[29595];
assign t[29596] = t[29595] ^ n[29596];
assign t[29597] = t[29596] ^ n[29597];
assign t[29598] = t[29597] ^ n[29598];
assign t[29599] = t[29598] ^ n[29599];
assign t[29600] = t[29599] ^ n[29600];
assign t[29601] = t[29600] ^ n[29601];
assign t[29602] = t[29601] ^ n[29602];
assign t[29603] = t[29602] ^ n[29603];
assign t[29604] = t[29603] ^ n[29604];
assign t[29605] = t[29604] ^ n[29605];
assign t[29606] = t[29605] ^ n[29606];
assign t[29607] = t[29606] ^ n[29607];
assign t[29608] = t[29607] ^ n[29608];
assign t[29609] = t[29608] ^ n[29609];
assign t[29610] = t[29609] ^ n[29610];
assign t[29611] = t[29610] ^ n[29611];
assign t[29612] = t[29611] ^ n[29612];
assign t[29613] = t[29612] ^ n[29613];
assign t[29614] = t[29613] ^ n[29614];
assign t[29615] = t[29614] ^ n[29615];
assign t[29616] = t[29615] ^ n[29616];
assign t[29617] = t[29616] ^ n[29617];
assign t[29618] = t[29617] ^ n[29618];
assign t[29619] = t[29618] ^ n[29619];
assign t[29620] = t[29619] ^ n[29620];
assign t[29621] = t[29620] ^ n[29621];
assign t[29622] = t[29621] ^ n[29622];
assign t[29623] = t[29622] ^ n[29623];
assign t[29624] = t[29623] ^ n[29624];
assign t[29625] = t[29624] ^ n[29625];
assign t[29626] = t[29625] ^ n[29626];
assign t[29627] = t[29626] ^ n[29627];
assign t[29628] = t[29627] ^ n[29628];
assign t[29629] = t[29628] ^ n[29629];
assign t[29630] = t[29629] ^ n[29630];
assign t[29631] = t[29630] ^ n[29631];
assign t[29632] = t[29631] ^ n[29632];
assign t[29633] = t[29632] ^ n[29633];
assign t[29634] = t[29633] ^ n[29634];
assign t[29635] = t[29634] ^ n[29635];
assign t[29636] = t[29635] ^ n[29636];
assign t[29637] = t[29636] ^ n[29637];
assign t[29638] = t[29637] ^ n[29638];
assign t[29639] = t[29638] ^ n[29639];
assign t[29640] = t[29639] ^ n[29640];
assign t[29641] = t[29640] ^ n[29641];
assign t[29642] = t[29641] ^ n[29642];
assign t[29643] = t[29642] ^ n[29643];
assign t[29644] = t[29643] ^ n[29644];
assign t[29645] = t[29644] ^ n[29645];
assign t[29646] = t[29645] ^ n[29646];
assign t[29647] = t[29646] ^ n[29647];
assign t[29648] = t[29647] ^ n[29648];
assign t[29649] = t[29648] ^ n[29649];
assign t[29650] = t[29649] ^ n[29650];
assign t[29651] = t[29650] ^ n[29651];
assign t[29652] = t[29651] ^ n[29652];
assign t[29653] = t[29652] ^ n[29653];
assign t[29654] = t[29653] ^ n[29654];
assign t[29655] = t[29654] ^ n[29655];
assign t[29656] = t[29655] ^ n[29656];
assign t[29657] = t[29656] ^ n[29657];
assign t[29658] = t[29657] ^ n[29658];
assign t[29659] = t[29658] ^ n[29659];
assign t[29660] = t[29659] ^ n[29660];
assign t[29661] = t[29660] ^ n[29661];
assign t[29662] = t[29661] ^ n[29662];
assign t[29663] = t[29662] ^ n[29663];
assign t[29664] = t[29663] ^ n[29664];
assign t[29665] = t[29664] ^ n[29665];
assign t[29666] = t[29665] ^ n[29666];
assign t[29667] = t[29666] ^ n[29667];
assign t[29668] = t[29667] ^ n[29668];
assign t[29669] = t[29668] ^ n[29669];
assign t[29670] = t[29669] ^ n[29670];
assign t[29671] = t[29670] ^ n[29671];
assign t[29672] = t[29671] ^ n[29672];
assign t[29673] = t[29672] ^ n[29673];
assign t[29674] = t[29673] ^ n[29674];
assign t[29675] = t[29674] ^ n[29675];
assign t[29676] = t[29675] ^ n[29676];
assign t[29677] = t[29676] ^ n[29677];
assign t[29678] = t[29677] ^ n[29678];
assign t[29679] = t[29678] ^ n[29679];
assign t[29680] = t[29679] ^ n[29680];
assign t[29681] = t[29680] ^ n[29681];
assign t[29682] = t[29681] ^ n[29682];
assign t[29683] = t[29682] ^ n[29683];
assign t[29684] = t[29683] ^ n[29684];
assign t[29685] = t[29684] ^ n[29685];
assign t[29686] = t[29685] ^ n[29686];
assign t[29687] = t[29686] ^ n[29687];
assign t[29688] = t[29687] ^ n[29688];
assign t[29689] = t[29688] ^ n[29689];
assign t[29690] = t[29689] ^ n[29690];
assign t[29691] = t[29690] ^ n[29691];
assign t[29692] = t[29691] ^ n[29692];
assign t[29693] = t[29692] ^ n[29693];
assign t[29694] = t[29693] ^ n[29694];
assign t[29695] = t[29694] ^ n[29695];
assign t[29696] = t[29695] ^ n[29696];
assign t[29697] = t[29696] ^ n[29697];
assign t[29698] = t[29697] ^ n[29698];
assign t[29699] = t[29698] ^ n[29699];
assign t[29700] = t[29699] ^ n[29700];
assign t[29701] = t[29700] ^ n[29701];
assign t[29702] = t[29701] ^ n[29702];
assign t[29703] = t[29702] ^ n[29703];
assign t[29704] = t[29703] ^ n[29704];
assign t[29705] = t[29704] ^ n[29705];
assign t[29706] = t[29705] ^ n[29706];
assign t[29707] = t[29706] ^ n[29707];
assign t[29708] = t[29707] ^ n[29708];
assign t[29709] = t[29708] ^ n[29709];
assign t[29710] = t[29709] ^ n[29710];
assign t[29711] = t[29710] ^ n[29711];
assign t[29712] = t[29711] ^ n[29712];
assign t[29713] = t[29712] ^ n[29713];
assign t[29714] = t[29713] ^ n[29714];
assign t[29715] = t[29714] ^ n[29715];
assign t[29716] = t[29715] ^ n[29716];
assign t[29717] = t[29716] ^ n[29717];
assign t[29718] = t[29717] ^ n[29718];
assign t[29719] = t[29718] ^ n[29719];
assign t[29720] = t[29719] ^ n[29720];
assign t[29721] = t[29720] ^ n[29721];
assign t[29722] = t[29721] ^ n[29722];
assign t[29723] = t[29722] ^ n[29723];
assign t[29724] = t[29723] ^ n[29724];
assign t[29725] = t[29724] ^ n[29725];
assign t[29726] = t[29725] ^ n[29726];
assign t[29727] = t[29726] ^ n[29727];
assign t[29728] = t[29727] ^ n[29728];
assign t[29729] = t[29728] ^ n[29729];
assign t[29730] = t[29729] ^ n[29730];
assign t[29731] = t[29730] ^ n[29731];
assign t[29732] = t[29731] ^ n[29732];
assign t[29733] = t[29732] ^ n[29733];
assign t[29734] = t[29733] ^ n[29734];
assign t[29735] = t[29734] ^ n[29735];
assign t[29736] = t[29735] ^ n[29736];
assign t[29737] = t[29736] ^ n[29737];
assign t[29738] = t[29737] ^ n[29738];
assign t[29739] = t[29738] ^ n[29739];
assign t[29740] = t[29739] ^ n[29740];
assign t[29741] = t[29740] ^ n[29741];
assign t[29742] = t[29741] ^ n[29742];
assign t[29743] = t[29742] ^ n[29743];
assign t[29744] = t[29743] ^ n[29744];
assign t[29745] = t[29744] ^ n[29745];
assign t[29746] = t[29745] ^ n[29746];
assign t[29747] = t[29746] ^ n[29747];
assign t[29748] = t[29747] ^ n[29748];
assign t[29749] = t[29748] ^ n[29749];
assign t[29750] = t[29749] ^ n[29750];
assign t[29751] = t[29750] ^ n[29751];
assign t[29752] = t[29751] ^ n[29752];
assign t[29753] = t[29752] ^ n[29753];
assign t[29754] = t[29753] ^ n[29754];
assign t[29755] = t[29754] ^ n[29755];
assign t[29756] = t[29755] ^ n[29756];
assign t[29757] = t[29756] ^ n[29757];
assign t[29758] = t[29757] ^ n[29758];
assign t[29759] = t[29758] ^ n[29759];
assign t[29760] = t[29759] ^ n[29760];
assign t[29761] = t[29760] ^ n[29761];
assign t[29762] = t[29761] ^ n[29762];
assign t[29763] = t[29762] ^ n[29763];
assign t[29764] = t[29763] ^ n[29764];
assign t[29765] = t[29764] ^ n[29765];
assign t[29766] = t[29765] ^ n[29766];
assign t[29767] = t[29766] ^ n[29767];
assign t[29768] = t[29767] ^ n[29768];
assign t[29769] = t[29768] ^ n[29769];
assign t[29770] = t[29769] ^ n[29770];
assign t[29771] = t[29770] ^ n[29771];
assign t[29772] = t[29771] ^ n[29772];
assign t[29773] = t[29772] ^ n[29773];
assign t[29774] = t[29773] ^ n[29774];
assign t[29775] = t[29774] ^ n[29775];
assign t[29776] = t[29775] ^ n[29776];
assign t[29777] = t[29776] ^ n[29777];
assign t[29778] = t[29777] ^ n[29778];
assign t[29779] = t[29778] ^ n[29779];
assign t[29780] = t[29779] ^ n[29780];
assign t[29781] = t[29780] ^ n[29781];
assign t[29782] = t[29781] ^ n[29782];
assign t[29783] = t[29782] ^ n[29783];
assign t[29784] = t[29783] ^ n[29784];
assign t[29785] = t[29784] ^ n[29785];
assign t[29786] = t[29785] ^ n[29786];
assign t[29787] = t[29786] ^ n[29787];
assign t[29788] = t[29787] ^ n[29788];
assign t[29789] = t[29788] ^ n[29789];
assign t[29790] = t[29789] ^ n[29790];
assign t[29791] = t[29790] ^ n[29791];
assign t[29792] = t[29791] ^ n[29792];
assign t[29793] = t[29792] ^ n[29793];
assign t[29794] = t[29793] ^ n[29794];
assign t[29795] = t[29794] ^ n[29795];
assign t[29796] = t[29795] ^ n[29796];
assign t[29797] = t[29796] ^ n[29797];
assign t[29798] = t[29797] ^ n[29798];
assign t[29799] = t[29798] ^ n[29799];
assign t[29800] = t[29799] ^ n[29800];
assign t[29801] = t[29800] ^ n[29801];
assign t[29802] = t[29801] ^ n[29802];
assign t[29803] = t[29802] ^ n[29803];
assign t[29804] = t[29803] ^ n[29804];
assign t[29805] = t[29804] ^ n[29805];
assign t[29806] = t[29805] ^ n[29806];
assign t[29807] = t[29806] ^ n[29807];
assign t[29808] = t[29807] ^ n[29808];
assign t[29809] = t[29808] ^ n[29809];
assign t[29810] = t[29809] ^ n[29810];
assign t[29811] = t[29810] ^ n[29811];
assign t[29812] = t[29811] ^ n[29812];
assign t[29813] = t[29812] ^ n[29813];
assign t[29814] = t[29813] ^ n[29814];
assign t[29815] = t[29814] ^ n[29815];
assign t[29816] = t[29815] ^ n[29816];
assign t[29817] = t[29816] ^ n[29817];
assign t[29818] = t[29817] ^ n[29818];
assign t[29819] = t[29818] ^ n[29819];
assign t[29820] = t[29819] ^ n[29820];
assign t[29821] = t[29820] ^ n[29821];
assign t[29822] = t[29821] ^ n[29822];
assign t[29823] = t[29822] ^ n[29823];
assign t[29824] = t[29823] ^ n[29824];
assign t[29825] = t[29824] ^ n[29825];
assign t[29826] = t[29825] ^ n[29826];
assign t[29827] = t[29826] ^ n[29827];
assign t[29828] = t[29827] ^ n[29828];
assign t[29829] = t[29828] ^ n[29829];
assign t[29830] = t[29829] ^ n[29830];
assign t[29831] = t[29830] ^ n[29831];
assign t[29832] = t[29831] ^ n[29832];
assign t[29833] = t[29832] ^ n[29833];
assign t[29834] = t[29833] ^ n[29834];
assign t[29835] = t[29834] ^ n[29835];
assign t[29836] = t[29835] ^ n[29836];
assign t[29837] = t[29836] ^ n[29837];
assign t[29838] = t[29837] ^ n[29838];
assign t[29839] = t[29838] ^ n[29839];
assign t[29840] = t[29839] ^ n[29840];
assign t[29841] = t[29840] ^ n[29841];
assign t[29842] = t[29841] ^ n[29842];
assign t[29843] = t[29842] ^ n[29843];
assign t[29844] = t[29843] ^ n[29844];
assign t[29845] = t[29844] ^ n[29845];
assign t[29846] = t[29845] ^ n[29846];
assign t[29847] = t[29846] ^ n[29847];
assign t[29848] = t[29847] ^ n[29848];
assign t[29849] = t[29848] ^ n[29849];
assign t[29850] = t[29849] ^ n[29850];
assign t[29851] = t[29850] ^ n[29851];
assign t[29852] = t[29851] ^ n[29852];
assign t[29853] = t[29852] ^ n[29853];
assign t[29854] = t[29853] ^ n[29854];
assign t[29855] = t[29854] ^ n[29855];
assign t[29856] = t[29855] ^ n[29856];
assign t[29857] = t[29856] ^ n[29857];
assign t[29858] = t[29857] ^ n[29858];
assign t[29859] = t[29858] ^ n[29859];
assign t[29860] = t[29859] ^ n[29860];
assign t[29861] = t[29860] ^ n[29861];
assign t[29862] = t[29861] ^ n[29862];
assign t[29863] = t[29862] ^ n[29863];
assign t[29864] = t[29863] ^ n[29864];
assign t[29865] = t[29864] ^ n[29865];
assign t[29866] = t[29865] ^ n[29866];
assign t[29867] = t[29866] ^ n[29867];
assign t[29868] = t[29867] ^ n[29868];
assign t[29869] = t[29868] ^ n[29869];
assign t[29870] = t[29869] ^ n[29870];
assign t[29871] = t[29870] ^ n[29871];
assign t[29872] = t[29871] ^ n[29872];
assign t[29873] = t[29872] ^ n[29873];
assign t[29874] = t[29873] ^ n[29874];
assign t[29875] = t[29874] ^ n[29875];
assign t[29876] = t[29875] ^ n[29876];
assign t[29877] = t[29876] ^ n[29877];
assign t[29878] = t[29877] ^ n[29878];
assign t[29879] = t[29878] ^ n[29879];
assign t[29880] = t[29879] ^ n[29880];
assign t[29881] = t[29880] ^ n[29881];
assign t[29882] = t[29881] ^ n[29882];
assign t[29883] = t[29882] ^ n[29883];
assign t[29884] = t[29883] ^ n[29884];
assign t[29885] = t[29884] ^ n[29885];
assign t[29886] = t[29885] ^ n[29886];
assign t[29887] = t[29886] ^ n[29887];
assign t[29888] = t[29887] ^ n[29888];
assign t[29889] = t[29888] ^ n[29889];
assign t[29890] = t[29889] ^ n[29890];
assign t[29891] = t[29890] ^ n[29891];
assign t[29892] = t[29891] ^ n[29892];
assign t[29893] = t[29892] ^ n[29893];
assign t[29894] = t[29893] ^ n[29894];
assign t[29895] = t[29894] ^ n[29895];
assign t[29896] = t[29895] ^ n[29896];
assign t[29897] = t[29896] ^ n[29897];
assign t[29898] = t[29897] ^ n[29898];
assign t[29899] = t[29898] ^ n[29899];
assign t[29900] = t[29899] ^ n[29900];
assign t[29901] = t[29900] ^ n[29901];
assign t[29902] = t[29901] ^ n[29902];
assign t[29903] = t[29902] ^ n[29903];
assign t[29904] = t[29903] ^ n[29904];
assign t[29905] = t[29904] ^ n[29905];
assign t[29906] = t[29905] ^ n[29906];
assign t[29907] = t[29906] ^ n[29907];
assign t[29908] = t[29907] ^ n[29908];
assign t[29909] = t[29908] ^ n[29909];
assign t[29910] = t[29909] ^ n[29910];
assign t[29911] = t[29910] ^ n[29911];
assign t[29912] = t[29911] ^ n[29912];
assign t[29913] = t[29912] ^ n[29913];
assign t[29914] = t[29913] ^ n[29914];
assign t[29915] = t[29914] ^ n[29915];
assign t[29916] = t[29915] ^ n[29916];
assign t[29917] = t[29916] ^ n[29917];
assign t[29918] = t[29917] ^ n[29918];
assign t[29919] = t[29918] ^ n[29919];
assign t[29920] = t[29919] ^ n[29920];
assign t[29921] = t[29920] ^ n[29921];
assign t[29922] = t[29921] ^ n[29922];
assign t[29923] = t[29922] ^ n[29923];
assign t[29924] = t[29923] ^ n[29924];
assign t[29925] = t[29924] ^ n[29925];
assign t[29926] = t[29925] ^ n[29926];
assign t[29927] = t[29926] ^ n[29927];
assign t[29928] = t[29927] ^ n[29928];
assign t[29929] = t[29928] ^ n[29929];
assign t[29930] = t[29929] ^ n[29930];
assign t[29931] = t[29930] ^ n[29931];
assign t[29932] = t[29931] ^ n[29932];
assign t[29933] = t[29932] ^ n[29933];
assign t[29934] = t[29933] ^ n[29934];
assign t[29935] = t[29934] ^ n[29935];
assign t[29936] = t[29935] ^ n[29936];
assign t[29937] = t[29936] ^ n[29937];
assign t[29938] = t[29937] ^ n[29938];
assign t[29939] = t[29938] ^ n[29939];
assign t[29940] = t[29939] ^ n[29940];
assign t[29941] = t[29940] ^ n[29941];
assign t[29942] = t[29941] ^ n[29942];
assign t[29943] = t[29942] ^ n[29943];
assign t[29944] = t[29943] ^ n[29944];
assign t[29945] = t[29944] ^ n[29945];
assign t[29946] = t[29945] ^ n[29946];
assign t[29947] = t[29946] ^ n[29947];
assign t[29948] = t[29947] ^ n[29948];
assign t[29949] = t[29948] ^ n[29949];
assign t[29950] = t[29949] ^ n[29950];
assign t[29951] = t[29950] ^ n[29951];
assign t[29952] = t[29951] ^ n[29952];
assign t[29953] = t[29952] ^ n[29953];
assign t[29954] = t[29953] ^ n[29954];
assign t[29955] = t[29954] ^ n[29955];
assign t[29956] = t[29955] ^ n[29956];
assign t[29957] = t[29956] ^ n[29957];
assign t[29958] = t[29957] ^ n[29958];
assign t[29959] = t[29958] ^ n[29959];
assign t[29960] = t[29959] ^ n[29960];
assign t[29961] = t[29960] ^ n[29961];
assign t[29962] = t[29961] ^ n[29962];
assign t[29963] = t[29962] ^ n[29963];
assign t[29964] = t[29963] ^ n[29964];
assign t[29965] = t[29964] ^ n[29965];
assign t[29966] = t[29965] ^ n[29966];
assign t[29967] = t[29966] ^ n[29967];
assign t[29968] = t[29967] ^ n[29968];
assign t[29969] = t[29968] ^ n[29969];
assign t[29970] = t[29969] ^ n[29970];
assign t[29971] = t[29970] ^ n[29971];
assign t[29972] = t[29971] ^ n[29972];
assign t[29973] = t[29972] ^ n[29973];
assign t[29974] = t[29973] ^ n[29974];
assign t[29975] = t[29974] ^ n[29975];
assign t[29976] = t[29975] ^ n[29976];
assign t[29977] = t[29976] ^ n[29977];
assign t[29978] = t[29977] ^ n[29978];
assign t[29979] = t[29978] ^ n[29979];
assign t[29980] = t[29979] ^ n[29980];
assign t[29981] = t[29980] ^ n[29981];
assign t[29982] = t[29981] ^ n[29982];
assign t[29983] = t[29982] ^ n[29983];
assign t[29984] = t[29983] ^ n[29984];
assign t[29985] = t[29984] ^ n[29985];
assign t[29986] = t[29985] ^ n[29986];
assign t[29987] = t[29986] ^ n[29987];
assign t[29988] = t[29987] ^ n[29988];
assign t[29989] = t[29988] ^ n[29989];
assign t[29990] = t[29989] ^ n[29990];
assign t[29991] = t[29990] ^ n[29991];
assign t[29992] = t[29991] ^ n[29992];
assign t[29993] = t[29992] ^ n[29993];
assign t[29994] = t[29993] ^ n[29994];
assign t[29995] = t[29994] ^ n[29995];
assign t[29996] = t[29995] ^ n[29996];
assign t[29997] = t[29996] ^ n[29997];
assign t[29998] = t[29997] ^ n[29998];
assign t[29999] = t[29998] ^ n[29999];
assign t[30000] = t[29999] ^ n[30000];
assign t[30001] = t[30000] ^ n[30001];
assign t[30002] = t[30001] ^ n[30002];
assign t[30003] = t[30002] ^ n[30003];
assign t[30004] = t[30003] ^ n[30004];
assign t[30005] = t[30004] ^ n[30005];
assign t[30006] = t[30005] ^ n[30006];
assign t[30007] = t[30006] ^ n[30007];
assign t[30008] = t[30007] ^ n[30008];
assign t[30009] = t[30008] ^ n[30009];
assign t[30010] = t[30009] ^ n[30010];
assign t[30011] = t[30010] ^ n[30011];
assign t[30012] = t[30011] ^ n[30012];
assign t[30013] = t[30012] ^ n[30013];
assign t[30014] = t[30013] ^ n[30014];
assign t[30015] = t[30014] ^ n[30015];
assign t[30016] = t[30015] ^ n[30016];
assign t[30017] = t[30016] ^ n[30017];
assign t[30018] = t[30017] ^ n[30018];
assign t[30019] = t[30018] ^ n[30019];
assign t[30020] = t[30019] ^ n[30020];
assign t[30021] = t[30020] ^ n[30021];
assign t[30022] = t[30021] ^ n[30022];
assign t[30023] = t[30022] ^ n[30023];
assign t[30024] = t[30023] ^ n[30024];
assign t[30025] = t[30024] ^ n[30025];
assign t[30026] = t[30025] ^ n[30026];
assign t[30027] = t[30026] ^ n[30027];
assign t[30028] = t[30027] ^ n[30028];
assign t[30029] = t[30028] ^ n[30029];
assign t[30030] = t[30029] ^ n[30030];
assign t[30031] = t[30030] ^ n[30031];
assign t[30032] = t[30031] ^ n[30032];
assign t[30033] = t[30032] ^ n[30033];
assign t[30034] = t[30033] ^ n[30034];
assign t[30035] = t[30034] ^ n[30035];
assign t[30036] = t[30035] ^ n[30036];
assign t[30037] = t[30036] ^ n[30037];
assign t[30038] = t[30037] ^ n[30038];
assign t[30039] = t[30038] ^ n[30039];
assign t[30040] = t[30039] ^ n[30040];
assign t[30041] = t[30040] ^ n[30041];
assign t[30042] = t[30041] ^ n[30042];
assign t[30043] = t[30042] ^ n[30043];
assign t[30044] = t[30043] ^ n[30044];
assign t[30045] = t[30044] ^ n[30045];
assign t[30046] = t[30045] ^ n[30046];
assign t[30047] = t[30046] ^ n[30047];
assign t[30048] = t[30047] ^ n[30048];
assign t[30049] = t[30048] ^ n[30049];
assign t[30050] = t[30049] ^ n[30050];
assign t[30051] = t[30050] ^ n[30051];
assign t[30052] = t[30051] ^ n[30052];
assign t[30053] = t[30052] ^ n[30053];
assign t[30054] = t[30053] ^ n[30054];
assign t[30055] = t[30054] ^ n[30055];
assign t[30056] = t[30055] ^ n[30056];
assign t[30057] = t[30056] ^ n[30057];
assign t[30058] = t[30057] ^ n[30058];
assign t[30059] = t[30058] ^ n[30059];
assign t[30060] = t[30059] ^ n[30060];
assign t[30061] = t[30060] ^ n[30061];
assign t[30062] = t[30061] ^ n[30062];
assign t[30063] = t[30062] ^ n[30063];
assign t[30064] = t[30063] ^ n[30064];
assign t[30065] = t[30064] ^ n[30065];
assign t[30066] = t[30065] ^ n[30066];
assign t[30067] = t[30066] ^ n[30067];
assign t[30068] = t[30067] ^ n[30068];
assign t[30069] = t[30068] ^ n[30069];
assign t[30070] = t[30069] ^ n[30070];
assign t[30071] = t[30070] ^ n[30071];
assign t[30072] = t[30071] ^ n[30072];
assign t[30073] = t[30072] ^ n[30073];
assign t[30074] = t[30073] ^ n[30074];
assign t[30075] = t[30074] ^ n[30075];
assign t[30076] = t[30075] ^ n[30076];
assign t[30077] = t[30076] ^ n[30077];
assign t[30078] = t[30077] ^ n[30078];
assign t[30079] = t[30078] ^ n[30079];
assign t[30080] = t[30079] ^ n[30080];
assign t[30081] = t[30080] ^ n[30081];
assign t[30082] = t[30081] ^ n[30082];
assign t[30083] = t[30082] ^ n[30083];
assign t[30084] = t[30083] ^ n[30084];
assign t[30085] = t[30084] ^ n[30085];
assign t[30086] = t[30085] ^ n[30086];
assign t[30087] = t[30086] ^ n[30087];
assign t[30088] = t[30087] ^ n[30088];
assign t[30089] = t[30088] ^ n[30089];
assign t[30090] = t[30089] ^ n[30090];
assign t[30091] = t[30090] ^ n[30091];
assign t[30092] = t[30091] ^ n[30092];
assign t[30093] = t[30092] ^ n[30093];
assign t[30094] = t[30093] ^ n[30094];
assign t[30095] = t[30094] ^ n[30095];
assign t[30096] = t[30095] ^ n[30096];
assign t[30097] = t[30096] ^ n[30097];
assign t[30098] = t[30097] ^ n[30098];
assign t[30099] = t[30098] ^ n[30099];
assign t[30100] = t[30099] ^ n[30100];
assign t[30101] = t[30100] ^ n[30101];
assign t[30102] = t[30101] ^ n[30102];
assign t[30103] = t[30102] ^ n[30103];
assign t[30104] = t[30103] ^ n[30104];
assign t[30105] = t[30104] ^ n[30105];
assign t[30106] = t[30105] ^ n[30106];
assign t[30107] = t[30106] ^ n[30107];
assign t[30108] = t[30107] ^ n[30108];
assign t[30109] = t[30108] ^ n[30109];
assign t[30110] = t[30109] ^ n[30110];
assign t[30111] = t[30110] ^ n[30111];
assign t[30112] = t[30111] ^ n[30112];
assign t[30113] = t[30112] ^ n[30113];
assign t[30114] = t[30113] ^ n[30114];
assign t[30115] = t[30114] ^ n[30115];
assign t[30116] = t[30115] ^ n[30116];
assign t[30117] = t[30116] ^ n[30117];
assign t[30118] = t[30117] ^ n[30118];
assign t[30119] = t[30118] ^ n[30119];
assign t[30120] = t[30119] ^ n[30120];
assign t[30121] = t[30120] ^ n[30121];
assign t[30122] = t[30121] ^ n[30122];
assign t[30123] = t[30122] ^ n[30123];
assign t[30124] = t[30123] ^ n[30124];
assign t[30125] = t[30124] ^ n[30125];
assign t[30126] = t[30125] ^ n[30126];
assign t[30127] = t[30126] ^ n[30127];
assign t[30128] = t[30127] ^ n[30128];
assign t[30129] = t[30128] ^ n[30129];
assign t[30130] = t[30129] ^ n[30130];
assign t[30131] = t[30130] ^ n[30131];
assign t[30132] = t[30131] ^ n[30132];
assign t[30133] = t[30132] ^ n[30133];
assign t[30134] = t[30133] ^ n[30134];
assign t[30135] = t[30134] ^ n[30135];
assign t[30136] = t[30135] ^ n[30136];
assign t[30137] = t[30136] ^ n[30137];
assign t[30138] = t[30137] ^ n[30138];
assign t[30139] = t[30138] ^ n[30139];
assign t[30140] = t[30139] ^ n[30140];
assign t[30141] = t[30140] ^ n[30141];
assign t[30142] = t[30141] ^ n[30142];
assign t[30143] = t[30142] ^ n[30143];
assign t[30144] = t[30143] ^ n[30144];
assign t[30145] = t[30144] ^ n[30145];
assign t[30146] = t[30145] ^ n[30146];
assign t[30147] = t[30146] ^ n[30147];
assign t[30148] = t[30147] ^ n[30148];
assign t[30149] = t[30148] ^ n[30149];
assign t[30150] = t[30149] ^ n[30150];
assign t[30151] = t[30150] ^ n[30151];
assign t[30152] = t[30151] ^ n[30152];
assign t[30153] = t[30152] ^ n[30153];
assign t[30154] = t[30153] ^ n[30154];
assign t[30155] = t[30154] ^ n[30155];
assign t[30156] = t[30155] ^ n[30156];
assign t[30157] = t[30156] ^ n[30157];
assign t[30158] = t[30157] ^ n[30158];
assign t[30159] = t[30158] ^ n[30159];
assign t[30160] = t[30159] ^ n[30160];
assign t[30161] = t[30160] ^ n[30161];
assign t[30162] = t[30161] ^ n[30162];
assign t[30163] = t[30162] ^ n[30163];
assign t[30164] = t[30163] ^ n[30164];
assign t[30165] = t[30164] ^ n[30165];
assign t[30166] = t[30165] ^ n[30166];
assign t[30167] = t[30166] ^ n[30167];
assign t[30168] = t[30167] ^ n[30168];
assign t[30169] = t[30168] ^ n[30169];
assign t[30170] = t[30169] ^ n[30170];
assign t[30171] = t[30170] ^ n[30171];
assign t[30172] = t[30171] ^ n[30172];
assign t[30173] = t[30172] ^ n[30173];
assign t[30174] = t[30173] ^ n[30174];
assign t[30175] = t[30174] ^ n[30175];
assign t[30176] = t[30175] ^ n[30176];
assign t[30177] = t[30176] ^ n[30177];
assign t[30178] = t[30177] ^ n[30178];
assign t[30179] = t[30178] ^ n[30179];
assign t[30180] = t[30179] ^ n[30180];
assign t[30181] = t[30180] ^ n[30181];
assign t[30182] = t[30181] ^ n[30182];
assign t[30183] = t[30182] ^ n[30183];
assign t[30184] = t[30183] ^ n[30184];
assign t[30185] = t[30184] ^ n[30185];
assign t[30186] = t[30185] ^ n[30186];
assign t[30187] = t[30186] ^ n[30187];
assign t[30188] = t[30187] ^ n[30188];
assign t[30189] = t[30188] ^ n[30189];
assign t[30190] = t[30189] ^ n[30190];
assign t[30191] = t[30190] ^ n[30191];
assign t[30192] = t[30191] ^ n[30192];
assign t[30193] = t[30192] ^ n[30193];
assign t[30194] = t[30193] ^ n[30194];
assign t[30195] = t[30194] ^ n[30195];
assign t[30196] = t[30195] ^ n[30196];
assign t[30197] = t[30196] ^ n[30197];
assign t[30198] = t[30197] ^ n[30198];
assign t[30199] = t[30198] ^ n[30199];
assign t[30200] = t[30199] ^ n[30200];
assign t[30201] = t[30200] ^ n[30201];
assign t[30202] = t[30201] ^ n[30202];
assign t[30203] = t[30202] ^ n[30203];
assign t[30204] = t[30203] ^ n[30204];
assign t[30205] = t[30204] ^ n[30205];
assign t[30206] = t[30205] ^ n[30206];
assign t[30207] = t[30206] ^ n[30207];
assign t[30208] = t[30207] ^ n[30208];
assign t[30209] = t[30208] ^ n[30209];
assign t[30210] = t[30209] ^ n[30210];
assign t[30211] = t[30210] ^ n[30211];
assign t[30212] = t[30211] ^ n[30212];
assign t[30213] = t[30212] ^ n[30213];
assign t[30214] = t[30213] ^ n[30214];
assign t[30215] = t[30214] ^ n[30215];
assign t[30216] = t[30215] ^ n[30216];
assign t[30217] = t[30216] ^ n[30217];
assign t[30218] = t[30217] ^ n[30218];
assign t[30219] = t[30218] ^ n[30219];
assign t[30220] = t[30219] ^ n[30220];
assign t[30221] = t[30220] ^ n[30221];
assign t[30222] = t[30221] ^ n[30222];
assign t[30223] = t[30222] ^ n[30223];
assign t[30224] = t[30223] ^ n[30224];
assign t[30225] = t[30224] ^ n[30225];
assign t[30226] = t[30225] ^ n[30226];
assign t[30227] = t[30226] ^ n[30227];
assign t[30228] = t[30227] ^ n[30228];
assign t[30229] = t[30228] ^ n[30229];
assign t[30230] = t[30229] ^ n[30230];
assign t[30231] = t[30230] ^ n[30231];
assign t[30232] = t[30231] ^ n[30232];
assign t[30233] = t[30232] ^ n[30233];
assign t[30234] = t[30233] ^ n[30234];
assign t[30235] = t[30234] ^ n[30235];
assign t[30236] = t[30235] ^ n[30236];
assign t[30237] = t[30236] ^ n[30237];
assign t[30238] = t[30237] ^ n[30238];
assign t[30239] = t[30238] ^ n[30239];
assign t[30240] = t[30239] ^ n[30240];
assign t[30241] = t[30240] ^ n[30241];
assign t[30242] = t[30241] ^ n[30242];
assign t[30243] = t[30242] ^ n[30243];
assign t[30244] = t[30243] ^ n[30244];
assign t[30245] = t[30244] ^ n[30245];
assign t[30246] = t[30245] ^ n[30246];
assign t[30247] = t[30246] ^ n[30247];
assign t[30248] = t[30247] ^ n[30248];
assign t[30249] = t[30248] ^ n[30249];
assign t[30250] = t[30249] ^ n[30250];
assign t[30251] = t[30250] ^ n[30251];
assign t[30252] = t[30251] ^ n[30252];
assign t[30253] = t[30252] ^ n[30253];
assign t[30254] = t[30253] ^ n[30254];
assign t[30255] = t[30254] ^ n[30255];
assign t[30256] = t[30255] ^ n[30256];
assign t[30257] = t[30256] ^ n[30257];
assign t[30258] = t[30257] ^ n[30258];
assign t[30259] = t[30258] ^ n[30259];
assign t[30260] = t[30259] ^ n[30260];
assign t[30261] = t[30260] ^ n[30261];
assign t[30262] = t[30261] ^ n[30262];
assign t[30263] = t[30262] ^ n[30263];
assign t[30264] = t[30263] ^ n[30264];
assign t[30265] = t[30264] ^ n[30265];
assign t[30266] = t[30265] ^ n[30266];
assign t[30267] = t[30266] ^ n[30267];
assign t[30268] = t[30267] ^ n[30268];
assign t[30269] = t[30268] ^ n[30269];
assign t[30270] = t[30269] ^ n[30270];
assign t[30271] = t[30270] ^ n[30271];
assign t[30272] = t[30271] ^ n[30272];
assign t[30273] = t[30272] ^ n[30273];
assign t[30274] = t[30273] ^ n[30274];
assign t[30275] = t[30274] ^ n[30275];
assign t[30276] = t[30275] ^ n[30276];
assign t[30277] = t[30276] ^ n[30277];
assign t[30278] = t[30277] ^ n[30278];
assign t[30279] = t[30278] ^ n[30279];
assign t[30280] = t[30279] ^ n[30280];
assign t[30281] = t[30280] ^ n[30281];
assign t[30282] = t[30281] ^ n[30282];
assign t[30283] = t[30282] ^ n[30283];
assign t[30284] = t[30283] ^ n[30284];
assign t[30285] = t[30284] ^ n[30285];
assign t[30286] = t[30285] ^ n[30286];
assign t[30287] = t[30286] ^ n[30287];
assign t[30288] = t[30287] ^ n[30288];
assign t[30289] = t[30288] ^ n[30289];
assign t[30290] = t[30289] ^ n[30290];
assign t[30291] = t[30290] ^ n[30291];
assign t[30292] = t[30291] ^ n[30292];
assign t[30293] = t[30292] ^ n[30293];
assign t[30294] = t[30293] ^ n[30294];
assign t[30295] = t[30294] ^ n[30295];
assign t[30296] = t[30295] ^ n[30296];
assign t[30297] = t[30296] ^ n[30297];
assign t[30298] = t[30297] ^ n[30298];
assign t[30299] = t[30298] ^ n[30299];
assign t[30300] = t[30299] ^ n[30300];
assign t[30301] = t[30300] ^ n[30301];
assign t[30302] = t[30301] ^ n[30302];
assign t[30303] = t[30302] ^ n[30303];
assign t[30304] = t[30303] ^ n[30304];
assign t[30305] = t[30304] ^ n[30305];
assign t[30306] = t[30305] ^ n[30306];
assign t[30307] = t[30306] ^ n[30307];
assign t[30308] = t[30307] ^ n[30308];
assign t[30309] = t[30308] ^ n[30309];
assign t[30310] = t[30309] ^ n[30310];
assign t[30311] = t[30310] ^ n[30311];
assign t[30312] = t[30311] ^ n[30312];
assign t[30313] = t[30312] ^ n[30313];
assign t[30314] = t[30313] ^ n[30314];
assign t[30315] = t[30314] ^ n[30315];
assign t[30316] = t[30315] ^ n[30316];
assign t[30317] = t[30316] ^ n[30317];
assign t[30318] = t[30317] ^ n[30318];
assign t[30319] = t[30318] ^ n[30319];
assign t[30320] = t[30319] ^ n[30320];
assign t[30321] = t[30320] ^ n[30321];
assign t[30322] = t[30321] ^ n[30322];
assign t[30323] = t[30322] ^ n[30323];
assign t[30324] = t[30323] ^ n[30324];
assign t[30325] = t[30324] ^ n[30325];
assign t[30326] = t[30325] ^ n[30326];
assign t[30327] = t[30326] ^ n[30327];
assign t[30328] = t[30327] ^ n[30328];
assign t[30329] = t[30328] ^ n[30329];
assign t[30330] = t[30329] ^ n[30330];
assign t[30331] = t[30330] ^ n[30331];
assign t[30332] = t[30331] ^ n[30332];
assign t[30333] = t[30332] ^ n[30333];
assign t[30334] = t[30333] ^ n[30334];
assign t[30335] = t[30334] ^ n[30335];
assign t[30336] = t[30335] ^ n[30336];
assign t[30337] = t[30336] ^ n[30337];
assign t[30338] = t[30337] ^ n[30338];
assign t[30339] = t[30338] ^ n[30339];
assign t[30340] = t[30339] ^ n[30340];
assign t[30341] = t[30340] ^ n[30341];
assign t[30342] = t[30341] ^ n[30342];
assign t[30343] = t[30342] ^ n[30343];
assign t[30344] = t[30343] ^ n[30344];
assign t[30345] = t[30344] ^ n[30345];
assign t[30346] = t[30345] ^ n[30346];
assign t[30347] = t[30346] ^ n[30347];
assign t[30348] = t[30347] ^ n[30348];
assign t[30349] = t[30348] ^ n[30349];
assign t[30350] = t[30349] ^ n[30350];
assign t[30351] = t[30350] ^ n[30351];
assign t[30352] = t[30351] ^ n[30352];
assign t[30353] = t[30352] ^ n[30353];
assign t[30354] = t[30353] ^ n[30354];
assign t[30355] = t[30354] ^ n[30355];
assign t[30356] = t[30355] ^ n[30356];
assign t[30357] = t[30356] ^ n[30357];
assign t[30358] = t[30357] ^ n[30358];
assign t[30359] = t[30358] ^ n[30359];
assign t[30360] = t[30359] ^ n[30360];
assign t[30361] = t[30360] ^ n[30361];
assign t[30362] = t[30361] ^ n[30362];
assign t[30363] = t[30362] ^ n[30363];
assign t[30364] = t[30363] ^ n[30364];
assign t[30365] = t[30364] ^ n[30365];
assign t[30366] = t[30365] ^ n[30366];
assign t[30367] = t[30366] ^ n[30367];
assign t[30368] = t[30367] ^ n[30368];
assign t[30369] = t[30368] ^ n[30369];
assign t[30370] = t[30369] ^ n[30370];
assign t[30371] = t[30370] ^ n[30371];
assign t[30372] = t[30371] ^ n[30372];
assign t[30373] = t[30372] ^ n[30373];
assign t[30374] = t[30373] ^ n[30374];
assign t[30375] = t[30374] ^ n[30375];
assign t[30376] = t[30375] ^ n[30376];
assign t[30377] = t[30376] ^ n[30377];
assign t[30378] = t[30377] ^ n[30378];
assign t[30379] = t[30378] ^ n[30379];
assign t[30380] = t[30379] ^ n[30380];
assign t[30381] = t[30380] ^ n[30381];
assign t[30382] = t[30381] ^ n[30382];
assign t[30383] = t[30382] ^ n[30383];
assign t[30384] = t[30383] ^ n[30384];
assign t[30385] = t[30384] ^ n[30385];
assign t[30386] = t[30385] ^ n[30386];
assign t[30387] = t[30386] ^ n[30387];
assign t[30388] = t[30387] ^ n[30388];
assign t[30389] = t[30388] ^ n[30389];
assign t[30390] = t[30389] ^ n[30390];
assign t[30391] = t[30390] ^ n[30391];
assign t[30392] = t[30391] ^ n[30392];
assign t[30393] = t[30392] ^ n[30393];
assign t[30394] = t[30393] ^ n[30394];
assign t[30395] = t[30394] ^ n[30395];
assign t[30396] = t[30395] ^ n[30396];
assign t[30397] = t[30396] ^ n[30397];
assign t[30398] = t[30397] ^ n[30398];
assign t[30399] = t[30398] ^ n[30399];
assign t[30400] = t[30399] ^ n[30400];
assign t[30401] = t[30400] ^ n[30401];
assign t[30402] = t[30401] ^ n[30402];
assign t[30403] = t[30402] ^ n[30403];
assign t[30404] = t[30403] ^ n[30404];
assign t[30405] = t[30404] ^ n[30405];
assign t[30406] = t[30405] ^ n[30406];
assign t[30407] = t[30406] ^ n[30407];
assign t[30408] = t[30407] ^ n[30408];
assign t[30409] = t[30408] ^ n[30409];
assign t[30410] = t[30409] ^ n[30410];
assign t[30411] = t[30410] ^ n[30411];
assign t[30412] = t[30411] ^ n[30412];
assign t[30413] = t[30412] ^ n[30413];
assign t[30414] = t[30413] ^ n[30414];
assign t[30415] = t[30414] ^ n[30415];
assign t[30416] = t[30415] ^ n[30416];
assign t[30417] = t[30416] ^ n[30417];
assign t[30418] = t[30417] ^ n[30418];
assign t[30419] = t[30418] ^ n[30419];
assign t[30420] = t[30419] ^ n[30420];
assign t[30421] = t[30420] ^ n[30421];
assign t[30422] = t[30421] ^ n[30422];
assign t[30423] = t[30422] ^ n[30423];
assign t[30424] = t[30423] ^ n[30424];
assign t[30425] = t[30424] ^ n[30425];
assign t[30426] = t[30425] ^ n[30426];
assign t[30427] = t[30426] ^ n[30427];
assign t[30428] = t[30427] ^ n[30428];
assign t[30429] = t[30428] ^ n[30429];
assign t[30430] = t[30429] ^ n[30430];
assign t[30431] = t[30430] ^ n[30431];
assign t[30432] = t[30431] ^ n[30432];
assign t[30433] = t[30432] ^ n[30433];
assign t[30434] = t[30433] ^ n[30434];
assign t[30435] = t[30434] ^ n[30435];
assign t[30436] = t[30435] ^ n[30436];
assign t[30437] = t[30436] ^ n[30437];
assign t[30438] = t[30437] ^ n[30438];
assign t[30439] = t[30438] ^ n[30439];
assign t[30440] = t[30439] ^ n[30440];
assign t[30441] = t[30440] ^ n[30441];
assign t[30442] = t[30441] ^ n[30442];
assign t[30443] = t[30442] ^ n[30443];
assign t[30444] = t[30443] ^ n[30444];
assign t[30445] = t[30444] ^ n[30445];
assign t[30446] = t[30445] ^ n[30446];
assign t[30447] = t[30446] ^ n[30447];
assign t[30448] = t[30447] ^ n[30448];
assign t[30449] = t[30448] ^ n[30449];
assign t[30450] = t[30449] ^ n[30450];
assign t[30451] = t[30450] ^ n[30451];
assign t[30452] = t[30451] ^ n[30452];
assign t[30453] = t[30452] ^ n[30453];
assign t[30454] = t[30453] ^ n[30454];
assign t[30455] = t[30454] ^ n[30455];
assign t[30456] = t[30455] ^ n[30456];
assign t[30457] = t[30456] ^ n[30457];
assign t[30458] = t[30457] ^ n[30458];
assign t[30459] = t[30458] ^ n[30459];
assign t[30460] = t[30459] ^ n[30460];
assign t[30461] = t[30460] ^ n[30461];
assign t[30462] = t[30461] ^ n[30462];
assign t[30463] = t[30462] ^ n[30463];
assign t[30464] = t[30463] ^ n[30464];
assign t[30465] = t[30464] ^ n[30465];
assign t[30466] = t[30465] ^ n[30466];
assign t[30467] = t[30466] ^ n[30467];
assign t[30468] = t[30467] ^ n[30468];
assign t[30469] = t[30468] ^ n[30469];
assign t[30470] = t[30469] ^ n[30470];
assign t[30471] = t[30470] ^ n[30471];
assign t[30472] = t[30471] ^ n[30472];
assign t[30473] = t[30472] ^ n[30473];
assign t[30474] = t[30473] ^ n[30474];
assign t[30475] = t[30474] ^ n[30475];
assign t[30476] = t[30475] ^ n[30476];
assign t[30477] = t[30476] ^ n[30477];
assign t[30478] = t[30477] ^ n[30478];
assign t[30479] = t[30478] ^ n[30479];
assign t[30480] = t[30479] ^ n[30480];
assign t[30481] = t[30480] ^ n[30481];
assign t[30482] = t[30481] ^ n[30482];
assign t[30483] = t[30482] ^ n[30483];
assign t[30484] = t[30483] ^ n[30484];
assign t[30485] = t[30484] ^ n[30485];
assign t[30486] = t[30485] ^ n[30486];
assign t[30487] = t[30486] ^ n[30487];
assign t[30488] = t[30487] ^ n[30488];
assign t[30489] = t[30488] ^ n[30489];
assign t[30490] = t[30489] ^ n[30490];
assign t[30491] = t[30490] ^ n[30491];
assign t[30492] = t[30491] ^ n[30492];
assign t[30493] = t[30492] ^ n[30493];
assign t[30494] = t[30493] ^ n[30494];
assign t[30495] = t[30494] ^ n[30495];
assign t[30496] = t[30495] ^ n[30496];
assign t[30497] = t[30496] ^ n[30497];
assign t[30498] = t[30497] ^ n[30498];
assign t[30499] = t[30498] ^ n[30499];
assign t[30500] = t[30499] ^ n[30500];
assign t[30501] = t[30500] ^ n[30501];
assign t[30502] = t[30501] ^ n[30502];
assign t[30503] = t[30502] ^ n[30503];
assign t[30504] = t[30503] ^ n[30504];
assign t[30505] = t[30504] ^ n[30505];
assign t[30506] = t[30505] ^ n[30506];
assign t[30507] = t[30506] ^ n[30507];
assign t[30508] = t[30507] ^ n[30508];
assign t[30509] = t[30508] ^ n[30509];
assign t[30510] = t[30509] ^ n[30510];
assign t[30511] = t[30510] ^ n[30511];
assign t[30512] = t[30511] ^ n[30512];
assign t[30513] = t[30512] ^ n[30513];
assign t[30514] = t[30513] ^ n[30514];
assign t[30515] = t[30514] ^ n[30515];
assign t[30516] = t[30515] ^ n[30516];
assign t[30517] = t[30516] ^ n[30517];
assign t[30518] = t[30517] ^ n[30518];
assign t[30519] = t[30518] ^ n[30519];
assign t[30520] = t[30519] ^ n[30520];
assign t[30521] = t[30520] ^ n[30521];
assign t[30522] = t[30521] ^ n[30522];
assign t[30523] = t[30522] ^ n[30523];
assign t[30524] = t[30523] ^ n[30524];
assign t[30525] = t[30524] ^ n[30525];
assign t[30526] = t[30525] ^ n[30526];
assign t[30527] = t[30526] ^ n[30527];
assign t[30528] = t[30527] ^ n[30528];
assign t[30529] = t[30528] ^ n[30529];
assign t[30530] = t[30529] ^ n[30530];
assign t[30531] = t[30530] ^ n[30531];
assign t[30532] = t[30531] ^ n[30532];
assign t[30533] = t[30532] ^ n[30533];
assign t[30534] = t[30533] ^ n[30534];
assign t[30535] = t[30534] ^ n[30535];
assign t[30536] = t[30535] ^ n[30536];
assign t[30537] = t[30536] ^ n[30537];
assign t[30538] = t[30537] ^ n[30538];
assign t[30539] = t[30538] ^ n[30539];
assign t[30540] = t[30539] ^ n[30540];
assign t[30541] = t[30540] ^ n[30541];
assign t[30542] = t[30541] ^ n[30542];
assign t[30543] = t[30542] ^ n[30543];
assign t[30544] = t[30543] ^ n[30544];
assign t[30545] = t[30544] ^ n[30545];
assign t[30546] = t[30545] ^ n[30546];
assign t[30547] = t[30546] ^ n[30547];
assign t[30548] = t[30547] ^ n[30548];
assign t[30549] = t[30548] ^ n[30549];
assign t[30550] = t[30549] ^ n[30550];
assign t[30551] = t[30550] ^ n[30551];
assign t[30552] = t[30551] ^ n[30552];
assign t[30553] = t[30552] ^ n[30553];
assign t[30554] = t[30553] ^ n[30554];
assign t[30555] = t[30554] ^ n[30555];
assign t[30556] = t[30555] ^ n[30556];
assign t[30557] = t[30556] ^ n[30557];
assign t[30558] = t[30557] ^ n[30558];
assign t[30559] = t[30558] ^ n[30559];
assign t[30560] = t[30559] ^ n[30560];
assign t[30561] = t[30560] ^ n[30561];
assign t[30562] = t[30561] ^ n[30562];
assign t[30563] = t[30562] ^ n[30563];
assign t[30564] = t[30563] ^ n[30564];
assign t[30565] = t[30564] ^ n[30565];
assign t[30566] = t[30565] ^ n[30566];
assign t[30567] = t[30566] ^ n[30567];
assign t[30568] = t[30567] ^ n[30568];
assign t[30569] = t[30568] ^ n[30569];
assign t[30570] = t[30569] ^ n[30570];
assign t[30571] = t[30570] ^ n[30571];
assign t[30572] = t[30571] ^ n[30572];
assign t[30573] = t[30572] ^ n[30573];
assign t[30574] = t[30573] ^ n[30574];
assign t[30575] = t[30574] ^ n[30575];
assign t[30576] = t[30575] ^ n[30576];
assign t[30577] = t[30576] ^ n[30577];
assign t[30578] = t[30577] ^ n[30578];
assign t[30579] = t[30578] ^ n[30579];
assign t[30580] = t[30579] ^ n[30580];
assign t[30581] = t[30580] ^ n[30581];
assign t[30582] = t[30581] ^ n[30582];
assign t[30583] = t[30582] ^ n[30583];
assign t[30584] = t[30583] ^ n[30584];
assign t[30585] = t[30584] ^ n[30585];
assign t[30586] = t[30585] ^ n[30586];
assign t[30587] = t[30586] ^ n[30587];
assign t[30588] = t[30587] ^ n[30588];
assign t[30589] = t[30588] ^ n[30589];
assign t[30590] = t[30589] ^ n[30590];
assign t[30591] = t[30590] ^ n[30591];
assign t[30592] = t[30591] ^ n[30592];
assign t[30593] = t[30592] ^ n[30593];
assign t[30594] = t[30593] ^ n[30594];
assign t[30595] = t[30594] ^ n[30595];
assign t[30596] = t[30595] ^ n[30596];
assign t[30597] = t[30596] ^ n[30597];
assign t[30598] = t[30597] ^ n[30598];
assign t[30599] = t[30598] ^ n[30599];
assign t[30600] = t[30599] ^ n[30600];
assign t[30601] = t[30600] ^ n[30601];
assign t[30602] = t[30601] ^ n[30602];
assign t[30603] = t[30602] ^ n[30603];
assign t[30604] = t[30603] ^ n[30604];
assign t[30605] = t[30604] ^ n[30605];
assign t[30606] = t[30605] ^ n[30606];
assign t[30607] = t[30606] ^ n[30607];
assign t[30608] = t[30607] ^ n[30608];
assign t[30609] = t[30608] ^ n[30609];
assign t[30610] = t[30609] ^ n[30610];
assign t[30611] = t[30610] ^ n[30611];
assign t[30612] = t[30611] ^ n[30612];
assign t[30613] = t[30612] ^ n[30613];
assign t[30614] = t[30613] ^ n[30614];
assign t[30615] = t[30614] ^ n[30615];
assign t[30616] = t[30615] ^ n[30616];
assign t[30617] = t[30616] ^ n[30617];
assign t[30618] = t[30617] ^ n[30618];
assign t[30619] = t[30618] ^ n[30619];
assign t[30620] = t[30619] ^ n[30620];
assign t[30621] = t[30620] ^ n[30621];
assign t[30622] = t[30621] ^ n[30622];
assign t[30623] = t[30622] ^ n[30623];
assign t[30624] = t[30623] ^ n[30624];
assign t[30625] = t[30624] ^ n[30625];
assign t[30626] = t[30625] ^ n[30626];
assign t[30627] = t[30626] ^ n[30627];
assign t[30628] = t[30627] ^ n[30628];
assign t[30629] = t[30628] ^ n[30629];
assign t[30630] = t[30629] ^ n[30630];
assign t[30631] = t[30630] ^ n[30631];
assign t[30632] = t[30631] ^ n[30632];
assign t[30633] = t[30632] ^ n[30633];
assign t[30634] = t[30633] ^ n[30634];
assign t[30635] = t[30634] ^ n[30635];
assign t[30636] = t[30635] ^ n[30636];
assign t[30637] = t[30636] ^ n[30637];
assign t[30638] = t[30637] ^ n[30638];
assign t[30639] = t[30638] ^ n[30639];
assign t[30640] = t[30639] ^ n[30640];
assign t[30641] = t[30640] ^ n[30641];
assign t[30642] = t[30641] ^ n[30642];
assign t[30643] = t[30642] ^ n[30643];
assign t[30644] = t[30643] ^ n[30644];
assign t[30645] = t[30644] ^ n[30645];
assign t[30646] = t[30645] ^ n[30646];
assign t[30647] = t[30646] ^ n[30647];
assign t[30648] = t[30647] ^ n[30648];
assign t[30649] = t[30648] ^ n[30649];
assign t[30650] = t[30649] ^ n[30650];
assign t[30651] = t[30650] ^ n[30651];
assign t[30652] = t[30651] ^ n[30652];
assign t[30653] = t[30652] ^ n[30653];
assign t[30654] = t[30653] ^ n[30654];
assign t[30655] = t[30654] ^ n[30655];
assign t[30656] = t[30655] ^ n[30656];
assign t[30657] = t[30656] ^ n[30657];
assign t[30658] = t[30657] ^ n[30658];
assign t[30659] = t[30658] ^ n[30659];
assign t[30660] = t[30659] ^ n[30660];
assign t[30661] = t[30660] ^ n[30661];
assign t[30662] = t[30661] ^ n[30662];
assign t[30663] = t[30662] ^ n[30663];
assign t[30664] = t[30663] ^ n[30664];
assign t[30665] = t[30664] ^ n[30665];
assign t[30666] = t[30665] ^ n[30666];
assign t[30667] = t[30666] ^ n[30667];
assign t[30668] = t[30667] ^ n[30668];
assign t[30669] = t[30668] ^ n[30669];
assign t[30670] = t[30669] ^ n[30670];
assign t[30671] = t[30670] ^ n[30671];
assign t[30672] = t[30671] ^ n[30672];
assign t[30673] = t[30672] ^ n[30673];
assign t[30674] = t[30673] ^ n[30674];
assign t[30675] = t[30674] ^ n[30675];
assign t[30676] = t[30675] ^ n[30676];
assign t[30677] = t[30676] ^ n[30677];
assign t[30678] = t[30677] ^ n[30678];
assign t[30679] = t[30678] ^ n[30679];
assign t[30680] = t[30679] ^ n[30680];
assign t[30681] = t[30680] ^ n[30681];
assign t[30682] = t[30681] ^ n[30682];
assign t[30683] = t[30682] ^ n[30683];
assign t[30684] = t[30683] ^ n[30684];
assign t[30685] = t[30684] ^ n[30685];
assign t[30686] = t[30685] ^ n[30686];
assign t[30687] = t[30686] ^ n[30687];
assign t[30688] = t[30687] ^ n[30688];
assign t[30689] = t[30688] ^ n[30689];
assign t[30690] = t[30689] ^ n[30690];
assign t[30691] = t[30690] ^ n[30691];
assign t[30692] = t[30691] ^ n[30692];
assign t[30693] = t[30692] ^ n[30693];
assign t[30694] = t[30693] ^ n[30694];
assign t[30695] = t[30694] ^ n[30695];
assign t[30696] = t[30695] ^ n[30696];
assign t[30697] = t[30696] ^ n[30697];
assign t[30698] = t[30697] ^ n[30698];
assign t[30699] = t[30698] ^ n[30699];
assign t[30700] = t[30699] ^ n[30700];
assign t[30701] = t[30700] ^ n[30701];
assign t[30702] = t[30701] ^ n[30702];
assign t[30703] = t[30702] ^ n[30703];
assign t[30704] = t[30703] ^ n[30704];
assign t[30705] = t[30704] ^ n[30705];
assign t[30706] = t[30705] ^ n[30706];
assign t[30707] = t[30706] ^ n[30707];
assign t[30708] = t[30707] ^ n[30708];
assign t[30709] = t[30708] ^ n[30709];
assign t[30710] = t[30709] ^ n[30710];
assign t[30711] = t[30710] ^ n[30711];
assign t[30712] = t[30711] ^ n[30712];
assign t[30713] = t[30712] ^ n[30713];
assign t[30714] = t[30713] ^ n[30714];
assign t[30715] = t[30714] ^ n[30715];
assign t[30716] = t[30715] ^ n[30716];
assign t[30717] = t[30716] ^ n[30717];
assign t[30718] = t[30717] ^ n[30718];
assign t[30719] = t[30718] ^ n[30719];
assign t[30720] = t[30719] ^ n[30720];
assign t[30721] = t[30720] ^ n[30721];
assign t[30722] = t[30721] ^ n[30722];
assign t[30723] = t[30722] ^ n[30723];
assign t[30724] = t[30723] ^ n[30724];
assign t[30725] = t[30724] ^ n[30725];
assign t[30726] = t[30725] ^ n[30726];
assign t[30727] = t[30726] ^ n[30727];
assign t[30728] = t[30727] ^ n[30728];
assign t[30729] = t[30728] ^ n[30729];
assign t[30730] = t[30729] ^ n[30730];
assign t[30731] = t[30730] ^ n[30731];
assign t[30732] = t[30731] ^ n[30732];
assign t[30733] = t[30732] ^ n[30733];
assign t[30734] = t[30733] ^ n[30734];
assign t[30735] = t[30734] ^ n[30735];
assign t[30736] = t[30735] ^ n[30736];
assign t[30737] = t[30736] ^ n[30737];
assign t[30738] = t[30737] ^ n[30738];
assign t[30739] = t[30738] ^ n[30739];
assign t[30740] = t[30739] ^ n[30740];
assign t[30741] = t[30740] ^ n[30741];
assign t[30742] = t[30741] ^ n[30742];
assign t[30743] = t[30742] ^ n[30743];
assign t[30744] = t[30743] ^ n[30744];
assign t[30745] = t[30744] ^ n[30745];
assign t[30746] = t[30745] ^ n[30746];
assign t[30747] = t[30746] ^ n[30747];
assign t[30748] = t[30747] ^ n[30748];
assign t[30749] = t[30748] ^ n[30749];
assign t[30750] = t[30749] ^ n[30750];
assign t[30751] = t[30750] ^ n[30751];
assign t[30752] = t[30751] ^ n[30752];
assign t[30753] = t[30752] ^ n[30753];
assign t[30754] = t[30753] ^ n[30754];
assign t[30755] = t[30754] ^ n[30755];
assign t[30756] = t[30755] ^ n[30756];
assign t[30757] = t[30756] ^ n[30757];
assign t[30758] = t[30757] ^ n[30758];
assign t[30759] = t[30758] ^ n[30759];
assign t[30760] = t[30759] ^ n[30760];
assign t[30761] = t[30760] ^ n[30761];
assign t[30762] = t[30761] ^ n[30762];
assign t[30763] = t[30762] ^ n[30763];
assign t[30764] = t[30763] ^ n[30764];
assign t[30765] = t[30764] ^ n[30765];
assign t[30766] = t[30765] ^ n[30766];
assign t[30767] = t[30766] ^ n[30767];
assign t[30768] = t[30767] ^ n[30768];
assign t[30769] = t[30768] ^ n[30769];
assign t[30770] = t[30769] ^ n[30770];
assign t[30771] = t[30770] ^ n[30771];
assign t[30772] = t[30771] ^ n[30772];
assign t[30773] = t[30772] ^ n[30773];
assign t[30774] = t[30773] ^ n[30774];
assign t[30775] = t[30774] ^ n[30775];
assign t[30776] = t[30775] ^ n[30776];
assign t[30777] = t[30776] ^ n[30777];
assign t[30778] = t[30777] ^ n[30778];
assign t[30779] = t[30778] ^ n[30779];
assign t[30780] = t[30779] ^ n[30780];
assign t[30781] = t[30780] ^ n[30781];
assign t[30782] = t[30781] ^ n[30782];
assign t[30783] = t[30782] ^ n[30783];
assign t[30784] = t[30783] ^ n[30784];
assign t[30785] = t[30784] ^ n[30785];
assign t[30786] = t[30785] ^ n[30786];
assign t[30787] = t[30786] ^ n[30787];
assign t[30788] = t[30787] ^ n[30788];
assign t[30789] = t[30788] ^ n[30789];
assign t[30790] = t[30789] ^ n[30790];
assign t[30791] = t[30790] ^ n[30791];
assign t[30792] = t[30791] ^ n[30792];
assign t[30793] = t[30792] ^ n[30793];
assign t[30794] = t[30793] ^ n[30794];
assign t[30795] = t[30794] ^ n[30795];
assign t[30796] = t[30795] ^ n[30796];
assign t[30797] = t[30796] ^ n[30797];
assign t[30798] = t[30797] ^ n[30798];
assign t[30799] = t[30798] ^ n[30799];
assign t[30800] = t[30799] ^ n[30800];
assign t[30801] = t[30800] ^ n[30801];
assign t[30802] = t[30801] ^ n[30802];
assign t[30803] = t[30802] ^ n[30803];
assign t[30804] = t[30803] ^ n[30804];
assign t[30805] = t[30804] ^ n[30805];
assign t[30806] = t[30805] ^ n[30806];
assign t[30807] = t[30806] ^ n[30807];
assign t[30808] = t[30807] ^ n[30808];
assign t[30809] = t[30808] ^ n[30809];
assign t[30810] = t[30809] ^ n[30810];
assign t[30811] = t[30810] ^ n[30811];
assign t[30812] = t[30811] ^ n[30812];
assign t[30813] = t[30812] ^ n[30813];
assign t[30814] = t[30813] ^ n[30814];
assign t[30815] = t[30814] ^ n[30815];
assign t[30816] = t[30815] ^ n[30816];
assign t[30817] = t[30816] ^ n[30817];
assign t[30818] = t[30817] ^ n[30818];
assign t[30819] = t[30818] ^ n[30819];
assign t[30820] = t[30819] ^ n[30820];
assign t[30821] = t[30820] ^ n[30821];
assign t[30822] = t[30821] ^ n[30822];
assign t[30823] = t[30822] ^ n[30823];
assign t[30824] = t[30823] ^ n[30824];
assign t[30825] = t[30824] ^ n[30825];
assign t[30826] = t[30825] ^ n[30826];
assign t[30827] = t[30826] ^ n[30827];
assign t[30828] = t[30827] ^ n[30828];
assign t[30829] = t[30828] ^ n[30829];
assign t[30830] = t[30829] ^ n[30830];
assign t[30831] = t[30830] ^ n[30831];
assign t[30832] = t[30831] ^ n[30832];
assign t[30833] = t[30832] ^ n[30833];
assign t[30834] = t[30833] ^ n[30834];
assign t[30835] = t[30834] ^ n[30835];
assign t[30836] = t[30835] ^ n[30836];
assign t[30837] = t[30836] ^ n[30837];
assign t[30838] = t[30837] ^ n[30838];
assign t[30839] = t[30838] ^ n[30839];
assign t[30840] = t[30839] ^ n[30840];
assign t[30841] = t[30840] ^ n[30841];
assign t[30842] = t[30841] ^ n[30842];
assign t[30843] = t[30842] ^ n[30843];
assign t[30844] = t[30843] ^ n[30844];
assign t[30845] = t[30844] ^ n[30845];
assign t[30846] = t[30845] ^ n[30846];
assign t[30847] = t[30846] ^ n[30847];
assign t[30848] = t[30847] ^ n[30848];
assign t[30849] = t[30848] ^ n[30849];
assign t[30850] = t[30849] ^ n[30850];
assign t[30851] = t[30850] ^ n[30851];
assign t[30852] = t[30851] ^ n[30852];
assign t[30853] = t[30852] ^ n[30853];
assign t[30854] = t[30853] ^ n[30854];
assign t[30855] = t[30854] ^ n[30855];
assign t[30856] = t[30855] ^ n[30856];
assign t[30857] = t[30856] ^ n[30857];
assign t[30858] = t[30857] ^ n[30858];
assign t[30859] = t[30858] ^ n[30859];
assign t[30860] = t[30859] ^ n[30860];
assign t[30861] = t[30860] ^ n[30861];
assign t[30862] = t[30861] ^ n[30862];
assign t[30863] = t[30862] ^ n[30863];
assign t[30864] = t[30863] ^ n[30864];
assign t[30865] = t[30864] ^ n[30865];
assign t[30866] = t[30865] ^ n[30866];
assign t[30867] = t[30866] ^ n[30867];
assign t[30868] = t[30867] ^ n[30868];
assign t[30869] = t[30868] ^ n[30869];
assign t[30870] = t[30869] ^ n[30870];
assign t[30871] = t[30870] ^ n[30871];
assign t[30872] = t[30871] ^ n[30872];
assign t[30873] = t[30872] ^ n[30873];
assign t[30874] = t[30873] ^ n[30874];
assign t[30875] = t[30874] ^ n[30875];
assign t[30876] = t[30875] ^ n[30876];
assign t[30877] = t[30876] ^ n[30877];
assign t[30878] = t[30877] ^ n[30878];
assign t[30879] = t[30878] ^ n[30879];
assign t[30880] = t[30879] ^ n[30880];
assign t[30881] = t[30880] ^ n[30881];
assign t[30882] = t[30881] ^ n[30882];
assign t[30883] = t[30882] ^ n[30883];
assign t[30884] = t[30883] ^ n[30884];
assign t[30885] = t[30884] ^ n[30885];
assign t[30886] = t[30885] ^ n[30886];
assign t[30887] = t[30886] ^ n[30887];
assign t[30888] = t[30887] ^ n[30888];
assign t[30889] = t[30888] ^ n[30889];
assign t[30890] = t[30889] ^ n[30890];
assign t[30891] = t[30890] ^ n[30891];
assign t[30892] = t[30891] ^ n[30892];
assign t[30893] = t[30892] ^ n[30893];
assign t[30894] = t[30893] ^ n[30894];
assign t[30895] = t[30894] ^ n[30895];
assign t[30896] = t[30895] ^ n[30896];
assign t[30897] = t[30896] ^ n[30897];
assign t[30898] = t[30897] ^ n[30898];
assign t[30899] = t[30898] ^ n[30899];
assign t[30900] = t[30899] ^ n[30900];
assign t[30901] = t[30900] ^ n[30901];
assign t[30902] = t[30901] ^ n[30902];
assign t[30903] = t[30902] ^ n[30903];
assign t[30904] = t[30903] ^ n[30904];
assign t[30905] = t[30904] ^ n[30905];
assign t[30906] = t[30905] ^ n[30906];
assign t[30907] = t[30906] ^ n[30907];
assign t[30908] = t[30907] ^ n[30908];
assign t[30909] = t[30908] ^ n[30909];
assign t[30910] = t[30909] ^ n[30910];
assign t[30911] = t[30910] ^ n[30911];
assign t[30912] = t[30911] ^ n[30912];
assign t[30913] = t[30912] ^ n[30913];
assign t[30914] = t[30913] ^ n[30914];
assign t[30915] = t[30914] ^ n[30915];
assign t[30916] = t[30915] ^ n[30916];
assign t[30917] = t[30916] ^ n[30917];
assign t[30918] = t[30917] ^ n[30918];
assign t[30919] = t[30918] ^ n[30919];
assign t[30920] = t[30919] ^ n[30920];
assign t[30921] = t[30920] ^ n[30921];
assign t[30922] = t[30921] ^ n[30922];
assign t[30923] = t[30922] ^ n[30923];
assign t[30924] = t[30923] ^ n[30924];
assign t[30925] = t[30924] ^ n[30925];
assign t[30926] = t[30925] ^ n[30926];
assign t[30927] = t[30926] ^ n[30927];
assign t[30928] = t[30927] ^ n[30928];
assign t[30929] = t[30928] ^ n[30929];
assign t[30930] = t[30929] ^ n[30930];
assign t[30931] = t[30930] ^ n[30931];
assign t[30932] = t[30931] ^ n[30932];
assign t[30933] = t[30932] ^ n[30933];
assign t[30934] = t[30933] ^ n[30934];
assign t[30935] = t[30934] ^ n[30935];
assign t[30936] = t[30935] ^ n[30936];
assign t[30937] = t[30936] ^ n[30937];
assign t[30938] = t[30937] ^ n[30938];
assign t[30939] = t[30938] ^ n[30939];
assign t[30940] = t[30939] ^ n[30940];
assign t[30941] = t[30940] ^ n[30941];
assign t[30942] = t[30941] ^ n[30942];
assign t[30943] = t[30942] ^ n[30943];
assign t[30944] = t[30943] ^ n[30944];
assign t[30945] = t[30944] ^ n[30945];
assign t[30946] = t[30945] ^ n[30946];
assign t[30947] = t[30946] ^ n[30947];
assign t[30948] = t[30947] ^ n[30948];
assign t[30949] = t[30948] ^ n[30949];
assign t[30950] = t[30949] ^ n[30950];
assign t[30951] = t[30950] ^ n[30951];
assign t[30952] = t[30951] ^ n[30952];
assign t[30953] = t[30952] ^ n[30953];
assign t[30954] = t[30953] ^ n[30954];
assign t[30955] = t[30954] ^ n[30955];
assign t[30956] = t[30955] ^ n[30956];
assign t[30957] = t[30956] ^ n[30957];
assign t[30958] = t[30957] ^ n[30958];
assign t[30959] = t[30958] ^ n[30959];
assign t[30960] = t[30959] ^ n[30960];
assign t[30961] = t[30960] ^ n[30961];
assign t[30962] = t[30961] ^ n[30962];
assign t[30963] = t[30962] ^ n[30963];
assign t[30964] = t[30963] ^ n[30964];
assign t[30965] = t[30964] ^ n[30965];
assign t[30966] = t[30965] ^ n[30966];
assign t[30967] = t[30966] ^ n[30967];
assign t[30968] = t[30967] ^ n[30968];
assign t[30969] = t[30968] ^ n[30969];
assign t[30970] = t[30969] ^ n[30970];
assign t[30971] = t[30970] ^ n[30971];
assign t[30972] = t[30971] ^ n[30972];
assign t[30973] = t[30972] ^ n[30973];
assign t[30974] = t[30973] ^ n[30974];
assign t[30975] = t[30974] ^ n[30975];
assign t[30976] = t[30975] ^ n[30976];
assign t[30977] = t[30976] ^ n[30977];
assign t[30978] = t[30977] ^ n[30978];
assign t[30979] = t[30978] ^ n[30979];
assign t[30980] = t[30979] ^ n[30980];
assign t[30981] = t[30980] ^ n[30981];
assign t[30982] = t[30981] ^ n[30982];
assign t[30983] = t[30982] ^ n[30983];
assign t[30984] = t[30983] ^ n[30984];
assign t[30985] = t[30984] ^ n[30985];
assign t[30986] = t[30985] ^ n[30986];
assign t[30987] = t[30986] ^ n[30987];
assign t[30988] = t[30987] ^ n[30988];
assign t[30989] = t[30988] ^ n[30989];
assign t[30990] = t[30989] ^ n[30990];
assign t[30991] = t[30990] ^ n[30991];
assign t[30992] = t[30991] ^ n[30992];
assign t[30993] = t[30992] ^ n[30993];
assign t[30994] = t[30993] ^ n[30994];
assign t[30995] = t[30994] ^ n[30995];
assign t[30996] = t[30995] ^ n[30996];
assign t[30997] = t[30996] ^ n[30997];
assign t[30998] = t[30997] ^ n[30998];
assign t[30999] = t[30998] ^ n[30999];
assign t[31000] = t[30999] ^ n[31000];
assign t[31001] = t[31000] ^ n[31001];
assign t[31002] = t[31001] ^ n[31002];
assign t[31003] = t[31002] ^ n[31003];
assign t[31004] = t[31003] ^ n[31004];
assign t[31005] = t[31004] ^ n[31005];
assign t[31006] = t[31005] ^ n[31006];
assign t[31007] = t[31006] ^ n[31007];
assign t[31008] = t[31007] ^ n[31008];
assign t[31009] = t[31008] ^ n[31009];
assign t[31010] = t[31009] ^ n[31010];
assign t[31011] = t[31010] ^ n[31011];
assign t[31012] = t[31011] ^ n[31012];
assign t[31013] = t[31012] ^ n[31013];
assign t[31014] = t[31013] ^ n[31014];
assign t[31015] = t[31014] ^ n[31015];
assign t[31016] = t[31015] ^ n[31016];
assign t[31017] = t[31016] ^ n[31017];
assign t[31018] = t[31017] ^ n[31018];
assign t[31019] = t[31018] ^ n[31019];
assign t[31020] = t[31019] ^ n[31020];
assign t[31021] = t[31020] ^ n[31021];
assign t[31022] = t[31021] ^ n[31022];
assign t[31023] = t[31022] ^ n[31023];
assign t[31024] = t[31023] ^ n[31024];
assign t[31025] = t[31024] ^ n[31025];
assign t[31026] = t[31025] ^ n[31026];
assign t[31027] = t[31026] ^ n[31027];
assign t[31028] = t[31027] ^ n[31028];
assign t[31029] = t[31028] ^ n[31029];
assign t[31030] = t[31029] ^ n[31030];
assign t[31031] = t[31030] ^ n[31031];
assign t[31032] = t[31031] ^ n[31032];
assign t[31033] = t[31032] ^ n[31033];
assign t[31034] = t[31033] ^ n[31034];
assign t[31035] = t[31034] ^ n[31035];
assign t[31036] = t[31035] ^ n[31036];
assign t[31037] = t[31036] ^ n[31037];
assign t[31038] = t[31037] ^ n[31038];
assign t[31039] = t[31038] ^ n[31039];
assign t[31040] = t[31039] ^ n[31040];
assign t[31041] = t[31040] ^ n[31041];
assign t[31042] = t[31041] ^ n[31042];
assign t[31043] = t[31042] ^ n[31043];
assign t[31044] = t[31043] ^ n[31044];
assign t[31045] = t[31044] ^ n[31045];
assign t[31046] = t[31045] ^ n[31046];
assign t[31047] = t[31046] ^ n[31047];
assign t[31048] = t[31047] ^ n[31048];
assign t[31049] = t[31048] ^ n[31049];
assign t[31050] = t[31049] ^ n[31050];
assign t[31051] = t[31050] ^ n[31051];
assign t[31052] = t[31051] ^ n[31052];
assign t[31053] = t[31052] ^ n[31053];
assign t[31054] = t[31053] ^ n[31054];
assign t[31055] = t[31054] ^ n[31055];
assign t[31056] = t[31055] ^ n[31056];
assign t[31057] = t[31056] ^ n[31057];
assign t[31058] = t[31057] ^ n[31058];
assign t[31059] = t[31058] ^ n[31059];
assign t[31060] = t[31059] ^ n[31060];
assign t[31061] = t[31060] ^ n[31061];
assign t[31062] = t[31061] ^ n[31062];
assign t[31063] = t[31062] ^ n[31063];
assign t[31064] = t[31063] ^ n[31064];
assign t[31065] = t[31064] ^ n[31065];
assign t[31066] = t[31065] ^ n[31066];
assign t[31067] = t[31066] ^ n[31067];
assign t[31068] = t[31067] ^ n[31068];
assign t[31069] = t[31068] ^ n[31069];
assign t[31070] = t[31069] ^ n[31070];
assign t[31071] = t[31070] ^ n[31071];
assign t[31072] = t[31071] ^ n[31072];
assign t[31073] = t[31072] ^ n[31073];
assign t[31074] = t[31073] ^ n[31074];
assign t[31075] = t[31074] ^ n[31075];
assign t[31076] = t[31075] ^ n[31076];
assign t[31077] = t[31076] ^ n[31077];
assign t[31078] = t[31077] ^ n[31078];
assign t[31079] = t[31078] ^ n[31079];
assign t[31080] = t[31079] ^ n[31080];
assign t[31081] = t[31080] ^ n[31081];
assign t[31082] = t[31081] ^ n[31082];
assign t[31083] = t[31082] ^ n[31083];
assign t[31084] = t[31083] ^ n[31084];
assign t[31085] = t[31084] ^ n[31085];
assign t[31086] = t[31085] ^ n[31086];
assign t[31087] = t[31086] ^ n[31087];
assign t[31088] = t[31087] ^ n[31088];
assign t[31089] = t[31088] ^ n[31089];
assign t[31090] = t[31089] ^ n[31090];
assign t[31091] = t[31090] ^ n[31091];
assign t[31092] = t[31091] ^ n[31092];
assign t[31093] = t[31092] ^ n[31093];
assign t[31094] = t[31093] ^ n[31094];
assign t[31095] = t[31094] ^ n[31095];
assign t[31096] = t[31095] ^ n[31096];
assign t[31097] = t[31096] ^ n[31097];
assign t[31098] = t[31097] ^ n[31098];
assign t[31099] = t[31098] ^ n[31099];
assign t[31100] = t[31099] ^ n[31100];
assign t[31101] = t[31100] ^ n[31101];
assign t[31102] = t[31101] ^ n[31102];
assign t[31103] = t[31102] ^ n[31103];
assign t[31104] = t[31103] ^ n[31104];
assign t[31105] = t[31104] ^ n[31105];
assign t[31106] = t[31105] ^ n[31106];
assign t[31107] = t[31106] ^ n[31107];
assign t[31108] = t[31107] ^ n[31108];
assign t[31109] = t[31108] ^ n[31109];
assign t[31110] = t[31109] ^ n[31110];
assign t[31111] = t[31110] ^ n[31111];
assign t[31112] = t[31111] ^ n[31112];
assign t[31113] = t[31112] ^ n[31113];
assign t[31114] = t[31113] ^ n[31114];
assign t[31115] = t[31114] ^ n[31115];
assign t[31116] = t[31115] ^ n[31116];
assign t[31117] = t[31116] ^ n[31117];
assign t[31118] = t[31117] ^ n[31118];
assign t[31119] = t[31118] ^ n[31119];
assign t[31120] = t[31119] ^ n[31120];
assign t[31121] = t[31120] ^ n[31121];
assign t[31122] = t[31121] ^ n[31122];
assign t[31123] = t[31122] ^ n[31123];
assign t[31124] = t[31123] ^ n[31124];
assign t[31125] = t[31124] ^ n[31125];
assign t[31126] = t[31125] ^ n[31126];
assign t[31127] = t[31126] ^ n[31127];
assign t[31128] = t[31127] ^ n[31128];
assign t[31129] = t[31128] ^ n[31129];
assign t[31130] = t[31129] ^ n[31130];
assign t[31131] = t[31130] ^ n[31131];
assign t[31132] = t[31131] ^ n[31132];
assign t[31133] = t[31132] ^ n[31133];
assign t[31134] = t[31133] ^ n[31134];
assign t[31135] = t[31134] ^ n[31135];
assign t[31136] = t[31135] ^ n[31136];
assign t[31137] = t[31136] ^ n[31137];
assign t[31138] = t[31137] ^ n[31138];
assign t[31139] = t[31138] ^ n[31139];
assign t[31140] = t[31139] ^ n[31140];
assign t[31141] = t[31140] ^ n[31141];
assign t[31142] = t[31141] ^ n[31142];
assign t[31143] = t[31142] ^ n[31143];
assign t[31144] = t[31143] ^ n[31144];
assign t[31145] = t[31144] ^ n[31145];
assign t[31146] = t[31145] ^ n[31146];
assign t[31147] = t[31146] ^ n[31147];
assign t[31148] = t[31147] ^ n[31148];
assign t[31149] = t[31148] ^ n[31149];
assign t[31150] = t[31149] ^ n[31150];
assign t[31151] = t[31150] ^ n[31151];
assign t[31152] = t[31151] ^ n[31152];
assign t[31153] = t[31152] ^ n[31153];
assign t[31154] = t[31153] ^ n[31154];
assign t[31155] = t[31154] ^ n[31155];
assign t[31156] = t[31155] ^ n[31156];
assign t[31157] = t[31156] ^ n[31157];
assign t[31158] = t[31157] ^ n[31158];
assign t[31159] = t[31158] ^ n[31159];
assign t[31160] = t[31159] ^ n[31160];
assign t[31161] = t[31160] ^ n[31161];
assign t[31162] = t[31161] ^ n[31162];
assign t[31163] = t[31162] ^ n[31163];
assign t[31164] = t[31163] ^ n[31164];
assign t[31165] = t[31164] ^ n[31165];
assign t[31166] = t[31165] ^ n[31166];
assign t[31167] = t[31166] ^ n[31167];
assign t[31168] = t[31167] ^ n[31168];
assign t[31169] = t[31168] ^ n[31169];
assign t[31170] = t[31169] ^ n[31170];
assign t[31171] = t[31170] ^ n[31171];
assign t[31172] = t[31171] ^ n[31172];
assign t[31173] = t[31172] ^ n[31173];
assign t[31174] = t[31173] ^ n[31174];
assign t[31175] = t[31174] ^ n[31175];
assign t[31176] = t[31175] ^ n[31176];
assign t[31177] = t[31176] ^ n[31177];
assign t[31178] = t[31177] ^ n[31178];
assign t[31179] = t[31178] ^ n[31179];
assign t[31180] = t[31179] ^ n[31180];
assign t[31181] = t[31180] ^ n[31181];
assign t[31182] = t[31181] ^ n[31182];
assign t[31183] = t[31182] ^ n[31183];
assign t[31184] = t[31183] ^ n[31184];
assign t[31185] = t[31184] ^ n[31185];
assign t[31186] = t[31185] ^ n[31186];
assign t[31187] = t[31186] ^ n[31187];
assign t[31188] = t[31187] ^ n[31188];
assign t[31189] = t[31188] ^ n[31189];
assign t[31190] = t[31189] ^ n[31190];
assign t[31191] = t[31190] ^ n[31191];
assign t[31192] = t[31191] ^ n[31192];
assign t[31193] = t[31192] ^ n[31193];
assign t[31194] = t[31193] ^ n[31194];
assign t[31195] = t[31194] ^ n[31195];
assign t[31196] = t[31195] ^ n[31196];
assign t[31197] = t[31196] ^ n[31197];
assign t[31198] = t[31197] ^ n[31198];
assign t[31199] = t[31198] ^ n[31199];
assign t[31200] = t[31199] ^ n[31200];
assign t[31201] = t[31200] ^ n[31201];
assign t[31202] = t[31201] ^ n[31202];
assign t[31203] = t[31202] ^ n[31203];
assign t[31204] = t[31203] ^ n[31204];
assign t[31205] = t[31204] ^ n[31205];
assign t[31206] = t[31205] ^ n[31206];
assign t[31207] = t[31206] ^ n[31207];
assign t[31208] = t[31207] ^ n[31208];
assign t[31209] = t[31208] ^ n[31209];
assign t[31210] = t[31209] ^ n[31210];
assign t[31211] = t[31210] ^ n[31211];
assign t[31212] = t[31211] ^ n[31212];
assign t[31213] = t[31212] ^ n[31213];
assign t[31214] = t[31213] ^ n[31214];
assign t[31215] = t[31214] ^ n[31215];
assign t[31216] = t[31215] ^ n[31216];
assign t[31217] = t[31216] ^ n[31217];
assign t[31218] = t[31217] ^ n[31218];
assign t[31219] = t[31218] ^ n[31219];
assign t[31220] = t[31219] ^ n[31220];
assign t[31221] = t[31220] ^ n[31221];
assign t[31222] = t[31221] ^ n[31222];
assign t[31223] = t[31222] ^ n[31223];
assign t[31224] = t[31223] ^ n[31224];
assign t[31225] = t[31224] ^ n[31225];
assign t[31226] = t[31225] ^ n[31226];
assign t[31227] = t[31226] ^ n[31227];
assign t[31228] = t[31227] ^ n[31228];
assign t[31229] = t[31228] ^ n[31229];
assign t[31230] = t[31229] ^ n[31230];
assign t[31231] = t[31230] ^ n[31231];
assign t[31232] = t[31231] ^ n[31232];
assign t[31233] = t[31232] ^ n[31233];
assign t[31234] = t[31233] ^ n[31234];
assign t[31235] = t[31234] ^ n[31235];
assign t[31236] = t[31235] ^ n[31236];
assign t[31237] = t[31236] ^ n[31237];
assign t[31238] = t[31237] ^ n[31238];
assign t[31239] = t[31238] ^ n[31239];
assign t[31240] = t[31239] ^ n[31240];
assign t[31241] = t[31240] ^ n[31241];
assign t[31242] = t[31241] ^ n[31242];
assign t[31243] = t[31242] ^ n[31243];
assign t[31244] = t[31243] ^ n[31244];
assign t[31245] = t[31244] ^ n[31245];
assign t[31246] = t[31245] ^ n[31246];
assign t[31247] = t[31246] ^ n[31247];
assign t[31248] = t[31247] ^ n[31248];
assign t[31249] = t[31248] ^ n[31249];
assign t[31250] = t[31249] ^ n[31250];
assign t[31251] = t[31250] ^ n[31251];
assign t[31252] = t[31251] ^ n[31252];
assign t[31253] = t[31252] ^ n[31253];
assign t[31254] = t[31253] ^ n[31254];
assign t[31255] = t[31254] ^ n[31255];
assign t[31256] = t[31255] ^ n[31256];
assign t[31257] = t[31256] ^ n[31257];
assign t[31258] = t[31257] ^ n[31258];
assign t[31259] = t[31258] ^ n[31259];
assign t[31260] = t[31259] ^ n[31260];
assign t[31261] = t[31260] ^ n[31261];
assign t[31262] = t[31261] ^ n[31262];
assign t[31263] = t[31262] ^ n[31263];
assign t[31264] = t[31263] ^ n[31264];
assign t[31265] = t[31264] ^ n[31265];
assign t[31266] = t[31265] ^ n[31266];
assign t[31267] = t[31266] ^ n[31267];
assign t[31268] = t[31267] ^ n[31268];
assign t[31269] = t[31268] ^ n[31269];
assign t[31270] = t[31269] ^ n[31270];
assign t[31271] = t[31270] ^ n[31271];
assign t[31272] = t[31271] ^ n[31272];
assign t[31273] = t[31272] ^ n[31273];
assign t[31274] = t[31273] ^ n[31274];
assign t[31275] = t[31274] ^ n[31275];
assign t[31276] = t[31275] ^ n[31276];
assign t[31277] = t[31276] ^ n[31277];
assign t[31278] = t[31277] ^ n[31278];
assign t[31279] = t[31278] ^ n[31279];
assign t[31280] = t[31279] ^ n[31280];
assign t[31281] = t[31280] ^ n[31281];
assign t[31282] = t[31281] ^ n[31282];
assign t[31283] = t[31282] ^ n[31283];
assign t[31284] = t[31283] ^ n[31284];
assign t[31285] = t[31284] ^ n[31285];
assign t[31286] = t[31285] ^ n[31286];
assign t[31287] = t[31286] ^ n[31287];
assign t[31288] = t[31287] ^ n[31288];
assign t[31289] = t[31288] ^ n[31289];
assign t[31290] = t[31289] ^ n[31290];
assign t[31291] = t[31290] ^ n[31291];
assign t[31292] = t[31291] ^ n[31292];
assign t[31293] = t[31292] ^ n[31293];
assign t[31294] = t[31293] ^ n[31294];
assign t[31295] = t[31294] ^ n[31295];
assign t[31296] = t[31295] ^ n[31296];
assign t[31297] = t[31296] ^ n[31297];
assign t[31298] = t[31297] ^ n[31298];
assign t[31299] = t[31298] ^ n[31299];
assign t[31300] = t[31299] ^ n[31300];
assign t[31301] = t[31300] ^ n[31301];
assign t[31302] = t[31301] ^ n[31302];
assign t[31303] = t[31302] ^ n[31303];
assign t[31304] = t[31303] ^ n[31304];
assign t[31305] = t[31304] ^ n[31305];
assign t[31306] = t[31305] ^ n[31306];
assign t[31307] = t[31306] ^ n[31307];
assign t[31308] = t[31307] ^ n[31308];
assign t[31309] = t[31308] ^ n[31309];
assign t[31310] = t[31309] ^ n[31310];
assign t[31311] = t[31310] ^ n[31311];
assign t[31312] = t[31311] ^ n[31312];
assign t[31313] = t[31312] ^ n[31313];
assign t[31314] = t[31313] ^ n[31314];
assign t[31315] = t[31314] ^ n[31315];
assign t[31316] = t[31315] ^ n[31316];
assign t[31317] = t[31316] ^ n[31317];
assign t[31318] = t[31317] ^ n[31318];
assign t[31319] = t[31318] ^ n[31319];
assign t[31320] = t[31319] ^ n[31320];
assign t[31321] = t[31320] ^ n[31321];
assign t[31322] = t[31321] ^ n[31322];
assign t[31323] = t[31322] ^ n[31323];
assign t[31324] = t[31323] ^ n[31324];
assign t[31325] = t[31324] ^ n[31325];
assign t[31326] = t[31325] ^ n[31326];
assign t[31327] = t[31326] ^ n[31327];
assign t[31328] = t[31327] ^ n[31328];
assign t[31329] = t[31328] ^ n[31329];
assign t[31330] = t[31329] ^ n[31330];
assign t[31331] = t[31330] ^ n[31331];
assign t[31332] = t[31331] ^ n[31332];
assign t[31333] = t[31332] ^ n[31333];
assign t[31334] = t[31333] ^ n[31334];
assign t[31335] = t[31334] ^ n[31335];
assign t[31336] = t[31335] ^ n[31336];
assign t[31337] = t[31336] ^ n[31337];
assign t[31338] = t[31337] ^ n[31338];
assign t[31339] = t[31338] ^ n[31339];
assign t[31340] = t[31339] ^ n[31340];
assign t[31341] = t[31340] ^ n[31341];
assign t[31342] = t[31341] ^ n[31342];
assign t[31343] = t[31342] ^ n[31343];
assign t[31344] = t[31343] ^ n[31344];
assign t[31345] = t[31344] ^ n[31345];
assign t[31346] = t[31345] ^ n[31346];
assign t[31347] = t[31346] ^ n[31347];
assign t[31348] = t[31347] ^ n[31348];
assign t[31349] = t[31348] ^ n[31349];
assign t[31350] = t[31349] ^ n[31350];
assign t[31351] = t[31350] ^ n[31351];
assign t[31352] = t[31351] ^ n[31352];
assign t[31353] = t[31352] ^ n[31353];
assign t[31354] = t[31353] ^ n[31354];
assign t[31355] = t[31354] ^ n[31355];
assign t[31356] = t[31355] ^ n[31356];
assign t[31357] = t[31356] ^ n[31357];
assign t[31358] = t[31357] ^ n[31358];
assign t[31359] = t[31358] ^ n[31359];
assign t[31360] = t[31359] ^ n[31360];
assign t[31361] = t[31360] ^ n[31361];
assign t[31362] = t[31361] ^ n[31362];
assign t[31363] = t[31362] ^ n[31363];
assign t[31364] = t[31363] ^ n[31364];
assign t[31365] = t[31364] ^ n[31365];
assign t[31366] = t[31365] ^ n[31366];
assign t[31367] = t[31366] ^ n[31367];
assign t[31368] = t[31367] ^ n[31368];
assign t[31369] = t[31368] ^ n[31369];
assign t[31370] = t[31369] ^ n[31370];
assign t[31371] = t[31370] ^ n[31371];
assign t[31372] = t[31371] ^ n[31372];
assign t[31373] = t[31372] ^ n[31373];
assign t[31374] = t[31373] ^ n[31374];
assign t[31375] = t[31374] ^ n[31375];
assign t[31376] = t[31375] ^ n[31376];
assign t[31377] = t[31376] ^ n[31377];
assign t[31378] = t[31377] ^ n[31378];
assign t[31379] = t[31378] ^ n[31379];
assign t[31380] = t[31379] ^ n[31380];
assign t[31381] = t[31380] ^ n[31381];
assign t[31382] = t[31381] ^ n[31382];
assign t[31383] = t[31382] ^ n[31383];
assign t[31384] = t[31383] ^ n[31384];
assign t[31385] = t[31384] ^ n[31385];
assign t[31386] = t[31385] ^ n[31386];
assign t[31387] = t[31386] ^ n[31387];
assign t[31388] = t[31387] ^ n[31388];
assign t[31389] = t[31388] ^ n[31389];
assign t[31390] = t[31389] ^ n[31390];
assign t[31391] = t[31390] ^ n[31391];
assign t[31392] = t[31391] ^ n[31392];
assign t[31393] = t[31392] ^ n[31393];
assign t[31394] = t[31393] ^ n[31394];
assign t[31395] = t[31394] ^ n[31395];
assign t[31396] = t[31395] ^ n[31396];
assign t[31397] = t[31396] ^ n[31397];
assign t[31398] = t[31397] ^ n[31398];
assign t[31399] = t[31398] ^ n[31399];
assign t[31400] = t[31399] ^ n[31400];
assign t[31401] = t[31400] ^ n[31401];
assign t[31402] = t[31401] ^ n[31402];
assign t[31403] = t[31402] ^ n[31403];
assign t[31404] = t[31403] ^ n[31404];
assign t[31405] = t[31404] ^ n[31405];
assign t[31406] = t[31405] ^ n[31406];
assign t[31407] = t[31406] ^ n[31407];
assign t[31408] = t[31407] ^ n[31408];
assign t[31409] = t[31408] ^ n[31409];
assign t[31410] = t[31409] ^ n[31410];
assign t[31411] = t[31410] ^ n[31411];
assign t[31412] = t[31411] ^ n[31412];
assign t[31413] = t[31412] ^ n[31413];
assign t[31414] = t[31413] ^ n[31414];
assign t[31415] = t[31414] ^ n[31415];
assign t[31416] = t[31415] ^ n[31416];
assign t[31417] = t[31416] ^ n[31417];
assign t[31418] = t[31417] ^ n[31418];
assign t[31419] = t[31418] ^ n[31419];
assign t[31420] = t[31419] ^ n[31420];
assign t[31421] = t[31420] ^ n[31421];
assign t[31422] = t[31421] ^ n[31422];
assign t[31423] = t[31422] ^ n[31423];
assign t[31424] = t[31423] ^ n[31424];
assign t[31425] = t[31424] ^ n[31425];
assign t[31426] = t[31425] ^ n[31426];
assign t[31427] = t[31426] ^ n[31427];
assign t[31428] = t[31427] ^ n[31428];
assign t[31429] = t[31428] ^ n[31429];
assign t[31430] = t[31429] ^ n[31430];
assign t[31431] = t[31430] ^ n[31431];
assign t[31432] = t[31431] ^ n[31432];
assign t[31433] = t[31432] ^ n[31433];
assign t[31434] = t[31433] ^ n[31434];
assign t[31435] = t[31434] ^ n[31435];
assign t[31436] = t[31435] ^ n[31436];
assign t[31437] = t[31436] ^ n[31437];
assign t[31438] = t[31437] ^ n[31438];
assign t[31439] = t[31438] ^ n[31439];
assign t[31440] = t[31439] ^ n[31440];
assign t[31441] = t[31440] ^ n[31441];
assign t[31442] = t[31441] ^ n[31442];
assign t[31443] = t[31442] ^ n[31443];
assign t[31444] = t[31443] ^ n[31444];
assign t[31445] = t[31444] ^ n[31445];
assign t[31446] = t[31445] ^ n[31446];
assign t[31447] = t[31446] ^ n[31447];
assign t[31448] = t[31447] ^ n[31448];
assign t[31449] = t[31448] ^ n[31449];
assign t[31450] = t[31449] ^ n[31450];
assign t[31451] = t[31450] ^ n[31451];
assign t[31452] = t[31451] ^ n[31452];
assign t[31453] = t[31452] ^ n[31453];
assign t[31454] = t[31453] ^ n[31454];
assign t[31455] = t[31454] ^ n[31455];
assign t[31456] = t[31455] ^ n[31456];
assign t[31457] = t[31456] ^ n[31457];
assign t[31458] = t[31457] ^ n[31458];
assign t[31459] = t[31458] ^ n[31459];
assign t[31460] = t[31459] ^ n[31460];
assign t[31461] = t[31460] ^ n[31461];
assign t[31462] = t[31461] ^ n[31462];
assign t[31463] = t[31462] ^ n[31463];
assign t[31464] = t[31463] ^ n[31464];
assign t[31465] = t[31464] ^ n[31465];
assign t[31466] = t[31465] ^ n[31466];
assign t[31467] = t[31466] ^ n[31467];
assign t[31468] = t[31467] ^ n[31468];
assign t[31469] = t[31468] ^ n[31469];
assign t[31470] = t[31469] ^ n[31470];
assign t[31471] = t[31470] ^ n[31471];
assign t[31472] = t[31471] ^ n[31472];
assign t[31473] = t[31472] ^ n[31473];
assign t[31474] = t[31473] ^ n[31474];
assign t[31475] = t[31474] ^ n[31475];
assign t[31476] = t[31475] ^ n[31476];
assign t[31477] = t[31476] ^ n[31477];
assign t[31478] = t[31477] ^ n[31478];
assign t[31479] = t[31478] ^ n[31479];
assign t[31480] = t[31479] ^ n[31480];
assign t[31481] = t[31480] ^ n[31481];
assign t[31482] = t[31481] ^ n[31482];
assign t[31483] = t[31482] ^ n[31483];
assign t[31484] = t[31483] ^ n[31484];
assign t[31485] = t[31484] ^ n[31485];
assign t[31486] = t[31485] ^ n[31486];
assign t[31487] = t[31486] ^ n[31487];
assign t[31488] = t[31487] ^ n[31488];
assign t[31489] = t[31488] ^ n[31489];
assign t[31490] = t[31489] ^ n[31490];
assign t[31491] = t[31490] ^ n[31491];
assign t[31492] = t[31491] ^ n[31492];
assign t[31493] = t[31492] ^ n[31493];
assign t[31494] = t[31493] ^ n[31494];
assign t[31495] = t[31494] ^ n[31495];
assign t[31496] = t[31495] ^ n[31496];
assign t[31497] = t[31496] ^ n[31497];
assign t[31498] = t[31497] ^ n[31498];
assign t[31499] = t[31498] ^ n[31499];
assign t[31500] = t[31499] ^ n[31500];
assign t[31501] = t[31500] ^ n[31501];
assign t[31502] = t[31501] ^ n[31502];
assign t[31503] = t[31502] ^ n[31503];
assign t[31504] = t[31503] ^ n[31504];
assign t[31505] = t[31504] ^ n[31505];
assign t[31506] = t[31505] ^ n[31506];
assign t[31507] = t[31506] ^ n[31507];
assign t[31508] = t[31507] ^ n[31508];
assign t[31509] = t[31508] ^ n[31509];
assign t[31510] = t[31509] ^ n[31510];
assign t[31511] = t[31510] ^ n[31511];
assign t[31512] = t[31511] ^ n[31512];
assign t[31513] = t[31512] ^ n[31513];
assign t[31514] = t[31513] ^ n[31514];
assign t[31515] = t[31514] ^ n[31515];
assign t[31516] = t[31515] ^ n[31516];
assign t[31517] = t[31516] ^ n[31517];
assign t[31518] = t[31517] ^ n[31518];
assign t[31519] = t[31518] ^ n[31519];
assign t[31520] = t[31519] ^ n[31520];
assign t[31521] = t[31520] ^ n[31521];
assign t[31522] = t[31521] ^ n[31522];
assign t[31523] = t[31522] ^ n[31523];
assign t[31524] = t[31523] ^ n[31524];
assign t[31525] = t[31524] ^ n[31525];
assign t[31526] = t[31525] ^ n[31526];
assign t[31527] = t[31526] ^ n[31527];
assign t[31528] = t[31527] ^ n[31528];
assign t[31529] = t[31528] ^ n[31529];
assign t[31530] = t[31529] ^ n[31530];
assign t[31531] = t[31530] ^ n[31531];
assign t[31532] = t[31531] ^ n[31532];
assign t[31533] = t[31532] ^ n[31533];
assign t[31534] = t[31533] ^ n[31534];
assign t[31535] = t[31534] ^ n[31535];
assign t[31536] = t[31535] ^ n[31536];
assign t[31537] = t[31536] ^ n[31537];
assign t[31538] = t[31537] ^ n[31538];
assign t[31539] = t[31538] ^ n[31539];
assign t[31540] = t[31539] ^ n[31540];
assign t[31541] = t[31540] ^ n[31541];
assign t[31542] = t[31541] ^ n[31542];
assign t[31543] = t[31542] ^ n[31543];
assign t[31544] = t[31543] ^ n[31544];
assign t[31545] = t[31544] ^ n[31545];
assign t[31546] = t[31545] ^ n[31546];
assign t[31547] = t[31546] ^ n[31547];
assign t[31548] = t[31547] ^ n[31548];
assign t[31549] = t[31548] ^ n[31549];
assign t[31550] = t[31549] ^ n[31550];
assign t[31551] = t[31550] ^ n[31551];
assign t[31552] = t[31551] ^ n[31552];
assign t[31553] = t[31552] ^ n[31553];
assign t[31554] = t[31553] ^ n[31554];
assign t[31555] = t[31554] ^ n[31555];
assign t[31556] = t[31555] ^ n[31556];
assign t[31557] = t[31556] ^ n[31557];
assign t[31558] = t[31557] ^ n[31558];
assign t[31559] = t[31558] ^ n[31559];
assign t[31560] = t[31559] ^ n[31560];
assign t[31561] = t[31560] ^ n[31561];
assign t[31562] = t[31561] ^ n[31562];
assign t[31563] = t[31562] ^ n[31563];
assign t[31564] = t[31563] ^ n[31564];
assign t[31565] = t[31564] ^ n[31565];
assign t[31566] = t[31565] ^ n[31566];
assign t[31567] = t[31566] ^ n[31567];
assign t[31568] = t[31567] ^ n[31568];
assign t[31569] = t[31568] ^ n[31569];
assign t[31570] = t[31569] ^ n[31570];
assign t[31571] = t[31570] ^ n[31571];
assign t[31572] = t[31571] ^ n[31572];
assign t[31573] = t[31572] ^ n[31573];
assign t[31574] = t[31573] ^ n[31574];
assign t[31575] = t[31574] ^ n[31575];
assign t[31576] = t[31575] ^ n[31576];
assign t[31577] = t[31576] ^ n[31577];
assign t[31578] = t[31577] ^ n[31578];
assign t[31579] = t[31578] ^ n[31579];
assign t[31580] = t[31579] ^ n[31580];
assign t[31581] = t[31580] ^ n[31581];
assign t[31582] = t[31581] ^ n[31582];
assign t[31583] = t[31582] ^ n[31583];
assign t[31584] = t[31583] ^ n[31584];
assign t[31585] = t[31584] ^ n[31585];
assign t[31586] = t[31585] ^ n[31586];
assign t[31587] = t[31586] ^ n[31587];
assign t[31588] = t[31587] ^ n[31588];
assign t[31589] = t[31588] ^ n[31589];
assign t[31590] = t[31589] ^ n[31590];
assign t[31591] = t[31590] ^ n[31591];
assign t[31592] = t[31591] ^ n[31592];
assign t[31593] = t[31592] ^ n[31593];
assign t[31594] = t[31593] ^ n[31594];
assign t[31595] = t[31594] ^ n[31595];
assign t[31596] = t[31595] ^ n[31596];
assign t[31597] = t[31596] ^ n[31597];
assign t[31598] = t[31597] ^ n[31598];
assign t[31599] = t[31598] ^ n[31599];
assign t[31600] = t[31599] ^ n[31600];
assign t[31601] = t[31600] ^ n[31601];
assign t[31602] = t[31601] ^ n[31602];
assign t[31603] = t[31602] ^ n[31603];
assign t[31604] = t[31603] ^ n[31604];
assign t[31605] = t[31604] ^ n[31605];
assign t[31606] = t[31605] ^ n[31606];
assign t[31607] = t[31606] ^ n[31607];
assign t[31608] = t[31607] ^ n[31608];
assign t[31609] = t[31608] ^ n[31609];
assign t[31610] = t[31609] ^ n[31610];
assign t[31611] = t[31610] ^ n[31611];
assign t[31612] = t[31611] ^ n[31612];
assign t[31613] = t[31612] ^ n[31613];
assign t[31614] = t[31613] ^ n[31614];
assign t[31615] = t[31614] ^ n[31615];
assign t[31616] = t[31615] ^ n[31616];
assign t[31617] = t[31616] ^ n[31617];
assign t[31618] = t[31617] ^ n[31618];
assign t[31619] = t[31618] ^ n[31619];
assign t[31620] = t[31619] ^ n[31620];
assign t[31621] = t[31620] ^ n[31621];
assign t[31622] = t[31621] ^ n[31622];
assign t[31623] = t[31622] ^ n[31623];
assign t[31624] = t[31623] ^ n[31624];
assign t[31625] = t[31624] ^ n[31625];
assign t[31626] = t[31625] ^ n[31626];
assign t[31627] = t[31626] ^ n[31627];
assign t[31628] = t[31627] ^ n[31628];
assign t[31629] = t[31628] ^ n[31629];
assign t[31630] = t[31629] ^ n[31630];
assign t[31631] = t[31630] ^ n[31631];
assign t[31632] = t[31631] ^ n[31632];
assign t[31633] = t[31632] ^ n[31633];
assign t[31634] = t[31633] ^ n[31634];
assign t[31635] = t[31634] ^ n[31635];
assign t[31636] = t[31635] ^ n[31636];
assign t[31637] = t[31636] ^ n[31637];
assign t[31638] = t[31637] ^ n[31638];
assign t[31639] = t[31638] ^ n[31639];
assign t[31640] = t[31639] ^ n[31640];
assign t[31641] = t[31640] ^ n[31641];
assign t[31642] = t[31641] ^ n[31642];
assign t[31643] = t[31642] ^ n[31643];
assign t[31644] = t[31643] ^ n[31644];
assign t[31645] = t[31644] ^ n[31645];
assign t[31646] = t[31645] ^ n[31646];
assign t[31647] = t[31646] ^ n[31647];
assign t[31648] = t[31647] ^ n[31648];
assign t[31649] = t[31648] ^ n[31649];
assign t[31650] = t[31649] ^ n[31650];
assign t[31651] = t[31650] ^ n[31651];
assign t[31652] = t[31651] ^ n[31652];
assign t[31653] = t[31652] ^ n[31653];
assign t[31654] = t[31653] ^ n[31654];
assign t[31655] = t[31654] ^ n[31655];
assign t[31656] = t[31655] ^ n[31656];
assign t[31657] = t[31656] ^ n[31657];
assign t[31658] = t[31657] ^ n[31658];
assign t[31659] = t[31658] ^ n[31659];
assign t[31660] = t[31659] ^ n[31660];
assign t[31661] = t[31660] ^ n[31661];
assign t[31662] = t[31661] ^ n[31662];
assign t[31663] = t[31662] ^ n[31663];
assign t[31664] = t[31663] ^ n[31664];
assign t[31665] = t[31664] ^ n[31665];
assign t[31666] = t[31665] ^ n[31666];
assign t[31667] = t[31666] ^ n[31667];
assign t[31668] = t[31667] ^ n[31668];
assign t[31669] = t[31668] ^ n[31669];
assign t[31670] = t[31669] ^ n[31670];
assign t[31671] = t[31670] ^ n[31671];
assign t[31672] = t[31671] ^ n[31672];
assign t[31673] = t[31672] ^ n[31673];
assign t[31674] = t[31673] ^ n[31674];
assign t[31675] = t[31674] ^ n[31675];
assign t[31676] = t[31675] ^ n[31676];
assign t[31677] = t[31676] ^ n[31677];
assign t[31678] = t[31677] ^ n[31678];
assign t[31679] = t[31678] ^ n[31679];
assign t[31680] = t[31679] ^ n[31680];
assign t[31681] = t[31680] ^ n[31681];
assign t[31682] = t[31681] ^ n[31682];
assign t[31683] = t[31682] ^ n[31683];
assign t[31684] = t[31683] ^ n[31684];
assign t[31685] = t[31684] ^ n[31685];
assign t[31686] = t[31685] ^ n[31686];
assign t[31687] = t[31686] ^ n[31687];
assign t[31688] = t[31687] ^ n[31688];
assign t[31689] = t[31688] ^ n[31689];
assign t[31690] = t[31689] ^ n[31690];
assign t[31691] = t[31690] ^ n[31691];
assign t[31692] = t[31691] ^ n[31692];
assign t[31693] = t[31692] ^ n[31693];
assign t[31694] = t[31693] ^ n[31694];
assign t[31695] = t[31694] ^ n[31695];
assign t[31696] = t[31695] ^ n[31696];
assign t[31697] = t[31696] ^ n[31697];
assign t[31698] = t[31697] ^ n[31698];
assign t[31699] = t[31698] ^ n[31699];
assign t[31700] = t[31699] ^ n[31700];
assign t[31701] = t[31700] ^ n[31701];
assign t[31702] = t[31701] ^ n[31702];
assign t[31703] = t[31702] ^ n[31703];
assign t[31704] = t[31703] ^ n[31704];
assign t[31705] = t[31704] ^ n[31705];
assign t[31706] = t[31705] ^ n[31706];
assign t[31707] = t[31706] ^ n[31707];
assign t[31708] = t[31707] ^ n[31708];
assign t[31709] = t[31708] ^ n[31709];
assign t[31710] = t[31709] ^ n[31710];
assign t[31711] = t[31710] ^ n[31711];
assign t[31712] = t[31711] ^ n[31712];
assign t[31713] = t[31712] ^ n[31713];
assign t[31714] = t[31713] ^ n[31714];
assign t[31715] = t[31714] ^ n[31715];
assign t[31716] = t[31715] ^ n[31716];
assign t[31717] = t[31716] ^ n[31717];
assign t[31718] = t[31717] ^ n[31718];
assign t[31719] = t[31718] ^ n[31719];
assign t[31720] = t[31719] ^ n[31720];
assign t[31721] = t[31720] ^ n[31721];
assign t[31722] = t[31721] ^ n[31722];
assign t[31723] = t[31722] ^ n[31723];
assign t[31724] = t[31723] ^ n[31724];
assign t[31725] = t[31724] ^ n[31725];
assign t[31726] = t[31725] ^ n[31726];
assign t[31727] = t[31726] ^ n[31727];
assign t[31728] = t[31727] ^ n[31728];
assign t[31729] = t[31728] ^ n[31729];
assign t[31730] = t[31729] ^ n[31730];
assign t[31731] = t[31730] ^ n[31731];
assign t[31732] = t[31731] ^ n[31732];
assign t[31733] = t[31732] ^ n[31733];
assign t[31734] = t[31733] ^ n[31734];
assign t[31735] = t[31734] ^ n[31735];
assign t[31736] = t[31735] ^ n[31736];
assign t[31737] = t[31736] ^ n[31737];
assign t[31738] = t[31737] ^ n[31738];
assign t[31739] = t[31738] ^ n[31739];
assign t[31740] = t[31739] ^ n[31740];
assign t[31741] = t[31740] ^ n[31741];
assign t[31742] = t[31741] ^ n[31742];
assign t[31743] = t[31742] ^ n[31743];
assign t[31744] = t[31743] ^ n[31744];
assign t[31745] = t[31744] ^ n[31745];
assign t[31746] = t[31745] ^ n[31746];
assign t[31747] = t[31746] ^ n[31747];
assign t[31748] = t[31747] ^ n[31748];
assign t[31749] = t[31748] ^ n[31749];
assign t[31750] = t[31749] ^ n[31750];
assign t[31751] = t[31750] ^ n[31751];
assign t[31752] = t[31751] ^ n[31752];
assign t[31753] = t[31752] ^ n[31753];
assign t[31754] = t[31753] ^ n[31754];
assign t[31755] = t[31754] ^ n[31755];
assign t[31756] = t[31755] ^ n[31756];
assign t[31757] = t[31756] ^ n[31757];
assign t[31758] = t[31757] ^ n[31758];
assign t[31759] = t[31758] ^ n[31759];
assign t[31760] = t[31759] ^ n[31760];
assign t[31761] = t[31760] ^ n[31761];
assign t[31762] = t[31761] ^ n[31762];
assign t[31763] = t[31762] ^ n[31763];
assign t[31764] = t[31763] ^ n[31764];
assign t[31765] = t[31764] ^ n[31765];
assign t[31766] = t[31765] ^ n[31766];
assign t[31767] = t[31766] ^ n[31767];
assign t[31768] = t[31767] ^ n[31768];
assign t[31769] = t[31768] ^ n[31769];
assign t[31770] = t[31769] ^ n[31770];
assign t[31771] = t[31770] ^ n[31771];
assign t[31772] = t[31771] ^ n[31772];
assign t[31773] = t[31772] ^ n[31773];
assign t[31774] = t[31773] ^ n[31774];
assign t[31775] = t[31774] ^ n[31775];
assign t[31776] = t[31775] ^ n[31776];
assign t[31777] = t[31776] ^ n[31777];
assign t[31778] = t[31777] ^ n[31778];
assign t[31779] = t[31778] ^ n[31779];
assign t[31780] = t[31779] ^ n[31780];
assign t[31781] = t[31780] ^ n[31781];
assign t[31782] = t[31781] ^ n[31782];
assign t[31783] = t[31782] ^ n[31783];
assign t[31784] = t[31783] ^ n[31784];
assign t[31785] = t[31784] ^ n[31785];
assign t[31786] = t[31785] ^ n[31786];
assign t[31787] = t[31786] ^ n[31787];
assign t[31788] = t[31787] ^ n[31788];
assign t[31789] = t[31788] ^ n[31789];
assign t[31790] = t[31789] ^ n[31790];
assign t[31791] = t[31790] ^ n[31791];
assign t[31792] = t[31791] ^ n[31792];
assign t[31793] = t[31792] ^ n[31793];
assign t[31794] = t[31793] ^ n[31794];
assign t[31795] = t[31794] ^ n[31795];
assign t[31796] = t[31795] ^ n[31796];
assign t[31797] = t[31796] ^ n[31797];
assign t[31798] = t[31797] ^ n[31798];
assign t[31799] = t[31798] ^ n[31799];
assign t[31800] = t[31799] ^ n[31800];
assign t[31801] = t[31800] ^ n[31801];
assign t[31802] = t[31801] ^ n[31802];
assign t[31803] = t[31802] ^ n[31803];
assign t[31804] = t[31803] ^ n[31804];
assign t[31805] = t[31804] ^ n[31805];
assign t[31806] = t[31805] ^ n[31806];
assign t[31807] = t[31806] ^ n[31807];
assign t[31808] = t[31807] ^ n[31808];
assign t[31809] = t[31808] ^ n[31809];
assign t[31810] = t[31809] ^ n[31810];
assign t[31811] = t[31810] ^ n[31811];
assign t[31812] = t[31811] ^ n[31812];
assign t[31813] = t[31812] ^ n[31813];
assign t[31814] = t[31813] ^ n[31814];
assign t[31815] = t[31814] ^ n[31815];
assign t[31816] = t[31815] ^ n[31816];
assign t[31817] = t[31816] ^ n[31817];
assign t[31818] = t[31817] ^ n[31818];
assign t[31819] = t[31818] ^ n[31819];
assign t[31820] = t[31819] ^ n[31820];
assign t[31821] = t[31820] ^ n[31821];
assign t[31822] = t[31821] ^ n[31822];
assign t[31823] = t[31822] ^ n[31823];
assign t[31824] = t[31823] ^ n[31824];
assign t[31825] = t[31824] ^ n[31825];
assign t[31826] = t[31825] ^ n[31826];
assign t[31827] = t[31826] ^ n[31827];
assign t[31828] = t[31827] ^ n[31828];
assign t[31829] = t[31828] ^ n[31829];
assign t[31830] = t[31829] ^ n[31830];
assign t[31831] = t[31830] ^ n[31831];
assign t[31832] = t[31831] ^ n[31832];
assign t[31833] = t[31832] ^ n[31833];
assign t[31834] = t[31833] ^ n[31834];
assign t[31835] = t[31834] ^ n[31835];
assign t[31836] = t[31835] ^ n[31836];
assign t[31837] = t[31836] ^ n[31837];
assign t[31838] = t[31837] ^ n[31838];
assign t[31839] = t[31838] ^ n[31839];
assign t[31840] = t[31839] ^ n[31840];
assign t[31841] = t[31840] ^ n[31841];
assign t[31842] = t[31841] ^ n[31842];
assign t[31843] = t[31842] ^ n[31843];
assign t[31844] = t[31843] ^ n[31844];
assign t[31845] = t[31844] ^ n[31845];
assign t[31846] = t[31845] ^ n[31846];
assign t[31847] = t[31846] ^ n[31847];
assign t[31848] = t[31847] ^ n[31848];
assign t[31849] = t[31848] ^ n[31849];
assign t[31850] = t[31849] ^ n[31850];
assign t[31851] = t[31850] ^ n[31851];
assign t[31852] = t[31851] ^ n[31852];
assign t[31853] = t[31852] ^ n[31853];
assign t[31854] = t[31853] ^ n[31854];
assign t[31855] = t[31854] ^ n[31855];
assign t[31856] = t[31855] ^ n[31856];
assign t[31857] = t[31856] ^ n[31857];
assign t[31858] = t[31857] ^ n[31858];
assign t[31859] = t[31858] ^ n[31859];
assign t[31860] = t[31859] ^ n[31860];
assign t[31861] = t[31860] ^ n[31861];
assign t[31862] = t[31861] ^ n[31862];
assign t[31863] = t[31862] ^ n[31863];
assign t[31864] = t[31863] ^ n[31864];
assign t[31865] = t[31864] ^ n[31865];
assign t[31866] = t[31865] ^ n[31866];
assign t[31867] = t[31866] ^ n[31867];
assign t[31868] = t[31867] ^ n[31868];
assign t[31869] = t[31868] ^ n[31869];
assign t[31870] = t[31869] ^ n[31870];
assign t[31871] = t[31870] ^ n[31871];
assign t[31872] = t[31871] ^ n[31872];
assign t[31873] = t[31872] ^ n[31873];
assign t[31874] = t[31873] ^ n[31874];
assign t[31875] = t[31874] ^ n[31875];
assign t[31876] = t[31875] ^ n[31876];
assign t[31877] = t[31876] ^ n[31877];
assign t[31878] = t[31877] ^ n[31878];
assign t[31879] = t[31878] ^ n[31879];
assign t[31880] = t[31879] ^ n[31880];
assign t[31881] = t[31880] ^ n[31881];
assign t[31882] = t[31881] ^ n[31882];
assign t[31883] = t[31882] ^ n[31883];
assign t[31884] = t[31883] ^ n[31884];
assign t[31885] = t[31884] ^ n[31885];
assign t[31886] = t[31885] ^ n[31886];
assign t[31887] = t[31886] ^ n[31887];
assign t[31888] = t[31887] ^ n[31888];
assign t[31889] = t[31888] ^ n[31889];
assign t[31890] = t[31889] ^ n[31890];
assign t[31891] = t[31890] ^ n[31891];
assign t[31892] = t[31891] ^ n[31892];
assign t[31893] = t[31892] ^ n[31893];
assign t[31894] = t[31893] ^ n[31894];
assign t[31895] = t[31894] ^ n[31895];
assign t[31896] = t[31895] ^ n[31896];
assign t[31897] = t[31896] ^ n[31897];
assign t[31898] = t[31897] ^ n[31898];
assign t[31899] = t[31898] ^ n[31899];
assign t[31900] = t[31899] ^ n[31900];
assign t[31901] = t[31900] ^ n[31901];
assign t[31902] = t[31901] ^ n[31902];
assign t[31903] = t[31902] ^ n[31903];
assign t[31904] = t[31903] ^ n[31904];
assign t[31905] = t[31904] ^ n[31905];
assign t[31906] = t[31905] ^ n[31906];
assign t[31907] = t[31906] ^ n[31907];
assign t[31908] = t[31907] ^ n[31908];
assign t[31909] = t[31908] ^ n[31909];
assign t[31910] = t[31909] ^ n[31910];
assign t[31911] = t[31910] ^ n[31911];
assign t[31912] = t[31911] ^ n[31912];
assign t[31913] = t[31912] ^ n[31913];
assign t[31914] = t[31913] ^ n[31914];
assign t[31915] = t[31914] ^ n[31915];
assign t[31916] = t[31915] ^ n[31916];
assign t[31917] = t[31916] ^ n[31917];
assign t[31918] = t[31917] ^ n[31918];
assign t[31919] = t[31918] ^ n[31919];
assign t[31920] = t[31919] ^ n[31920];
assign t[31921] = t[31920] ^ n[31921];
assign t[31922] = t[31921] ^ n[31922];
assign t[31923] = t[31922] ^ n[31923];
assign t[31924] = t[31923] ^ n[31924];
assign t[31925] = t[31924] ^ n[31925];
assign t[31926] = t[31925] ^ n[31926];
assign t[31927] = t[31926] ^ n[31927];
assign t[31928] = t[31927] ^ n[31928];
assign t[31929] = t[31928] ^ n[31929];
assign t[31930] = t[31929] ^ n[31930];
assign t[31931] = t[31930] ^ n[31931];
assign t[31932] = t[31931] ^ n[31932];
assign t[31933] = t[31932] ^ n[31933];
assign t[31934] = t[31933] ^ n[31934];
assign t[31935] = t[31934] ^ n[31935];
assign t[31936] = t[31935] ^ n[31936];
assign t[31937] = t[31936] ^ n[31937];
assign t[31938] = t[31937] ^ n[31938];
assign t[31939] = t[31938] ^ n[31939];
assign t[31940] = t[31939] ^ n[31940];
assign t[31941] = t[31940] ^ n[31941];
assign t[31942] = t[31941] ^ n[31942];
assign t[31943] = t[31942] ^ n[31943];
assign t[31944] = t[31943] ^ n[31944];
assign t[31945] = t[31944] ^ n[31945];
assign t[31946] = t[31945] ^ n[31946];
assign t[31947] = t[31946] ^ n[31947];
assign t[31948] = t[31947] ^ n[31948];
assign t[31949] = t[31948] ^ n[31949];
assign t[31950] = t[31949] ^ n[31950];
assign t[31951] = t[31950] ^ n[31951];
assign t[31952] = t[31951] ^ n[31952];
assign t[31953] = t[31952] ^ n[31953];
assign t[31954] = t[31953] ^ n[31954];
assign t[31955] = t[31954] ^ n[31955];
assign t[31956] = t[31955] ^ n[31956];
assign t[31957] = t[31956] ^ n[31957];
assign t[31958] = t[31957] ^ n[31958];
assign t[31959] = t[31958] ^ n[31959];
assign t[31960] = t[31959] ^ n[31960];
assign t[31961] = t[31960] ^ n[31961];
assign t[31962] = t[31961] ^ n[31962];
assign t[31963] = t[31962] ^ n[31963];
assign t[31964] = t[31963] ^ n[31964];
assign t[31965] = t[31964] ^ n[31965];
assign t[31966] = t[31965] ^ n[31966];
assign t[31967] = t[31966] ^ n[31967];
assign t[31968] = t[31967] ^ n[31968];
assign t[31969] = t[31968] ^ n[31969];
assign t[31970] = t[31969] ^ n[31970];
assign t[31971] = t[31970] ^ n[31971];
assign t[31972] = t[31971] ^ n[31972];
assign t[31973] = t[31972] ^ n[31973];
assign t[31974] = t[31973] ^ n[31974];
assign t[31975] = t[31974] ^ n[31975];
assign t[31976] = t[31975] ^ n[31976];
assign t[31977] = t[31976] ^ n[31977];
assign t[31978] = t[31977] ^ n[31978];
assign t[31979] = t[31978] ^ n[31979];
assign t[31980] = t[31979] ^ n[31980];
assign t[31981] = t[31980] ^ n[31981];
assign t[31982] = t[31981] ^ n[31982];
assign t[31983] = t[31982] ^ n[31983];
assign t[31984] = t[31983] ^ n[31984];
assign t[31985] = t[31984] ^ n[31985];
assign t[31986] = t[31985] ^ n[31986];
assign t[31987] = t[31986] ^ n[31987];
assign t[31988] = t[31987] ^ n[31988];
assign t[31989] = t[31988] ^ n[31989];
assign t[31990] = t[31989] ^ n[31990];
assign t[31991] = t[31990] ^ n[31991];
assign t[31992] = t[31991] ^ n[31992];
assign t[31993] = t[31992] ^ n[31993];
assign t[31994] = t[31993] ^ n[31994];
assign t[31995] = t[31994] ^ n[31995];
assign t[31996] = t[31995] ^ n[31996];
assign t[31997] = t[31996] ^ n[31997];
assign t[31998] = t[31997] ^ n[31998];
assign t[31999] = t[31998] ^ n[31999];
assign t[32000] = t[31999] ^ n[32000];
assign t[32001] = t[32000] ^ n[32001];
assign t[32002] = t[32001] ^ n[32002];
assign t[32003] = t[32002] ^ n[32003];
assign t[32004] = t[32003] ^ n[32004];
assign t[32005] = t[32004] ^ n[32005];
assign t[32006] = t[32005] ^ n[32006];
assign t[32007] = t[32006] ^ n[32007];
assign t[32008] = t[32007] ^ n[32008];
assign t[32009] = t[32008] ^ n[32009];
assign t[32010] = t[32009] ^ n[32010];
assign t[32011] = t[32010] ^ n[32011];
assign t[32012] = t[32011] ^ n[32012];
assign t[32013] = t[32012] ^ n[32013];
assign t[32014] = t[32013] ^ n[32014];
assign t[32015] = t[32014] ^ n[32015];
assign t[32016] = t[32015] ^ n[32016];
assign t[32017] = t[32016] ^ n[32017];
assign t[32018] = t[32017] ^ n[32018];
assign t[32019] = t[32018] ^ n[32019];
assign t[32020] = t[32019] ^ n[32020];
assign t[32021] = t[32020] ^ n[32021];
assign t[32022] = t[32021] ^ n[32022];
assign t[32023] = t[32022] ^ n[32023];
assign t[32024] = t[32023] ^ n[32024];
assign t[32025] = t[32024] ^ n[32025];
assign t[32026] = t[32025] ^ n[32026];
assign t[32027] = t[32026] ^ n[32027];
assign t[32028] = t[32027] ^ n[32028];
assign t[32029] = t[32028] ^ n[32029];
assign t[32030] = t[32029] ^ n[32030];
assign t[32031] = t[32030] ^ n[32031];
assign t[32032] = t[32031] ^ n[32032];
assign t[32033] = t[32032] ^ n[32033];
assign t[32034] = t[32033] ^ n[32034];
assign t[32035] = t[32034] ^ n[32035];
assign t[32036] = t[32035] ^ n[32036];
assign t[32037] = t[32036] ^ n[32037];
assign t[32038] = t[32037] ^ n[32038];
assign t[32039] = t[32038] ^ n[32039];
assign t[32040] = t[32039] ^ n[32040];
assign t[32041] = t[32040] ^ n[32041];
assign t[32042] = t[32041] ^ n[32042];
assign t[32043] = t[32042] ^ n[32043];
assign t[32044] = t[32043] ^ n[32044];
assign t[32045] = t[32044] ^ n[32045];
assign t[32046] = t[32045] ^ n[32046];
assign t[32047] = t[32046] ^ n[32047];
assign t[32048] = t[32047] ^ n[32048];
assign t[32049] = t[32048] ^ n[32049];
assign t[32050] = t[32049] ^ n[32050];
assign t[32051] = t[32050] ^ n[32051];
assign t[32052] = t[32051] ^ n[32052];
assign t[32053] = t[32052] ^ n[32053];
assign t[32054] = t[32053] ^ n[32054];
assign t[32055] = t[32054] ^ n[32055];
assign t[32056] = t[32055] ^ n[32056];
assign t[32057] = t[32056] ^ n[32057];
assign t[32058] = t[32057] ^ n[32058];
assign t[32059] = t[32058] ^ n[32059];
assign t[32060] = t[32059] ^ n[32060];
assign t[32061] = t[32060] ^ n[32061];
assign t[32062] = t[32061] ^ n[32062];
assign t[32063] = t[32062] ^ n[32063];
assign t[32064] = t[32063] ^ n[32064];
assign t[32065] = t[32064] ^ n[32065];
assign t[32066] = t[32065] ^ n[32066];
assign t[32067] = t[32066] ^ n[32067];
assign t[32068] = t[32067] ^ n[32068];
assign t[32069] = t[32068] ^ n[32069];
assign t[32070] = t[32069] ^ n[32070];
assign t[32071] = t[32070] ^ n[32071];
assign t[32072] = t[32071] ^ n[32072];
assign t[32073] = t[32072] ^ n[32073];
assign t[32074] = t[32073] ^ n[32074];
assign t[32075] = t[32074] ^ n[32075];
assign t[32076] = t[32075] ^ n[32076];
assign t[32077] = t[32076] ^ n[32077];
assign t[32078] = t[32077] ^ n[32078];
assign t[32079] = t[32078] ^ n[32079];
assign t[32080] = t[32079] ^ n[32080];
assign t[32081] = t[32080] ^ n[32081];
assign t[32082] = t[32081] ^ n[32082];
assign t[32083] = t[32082] ^ n[32083];
assign t[32084] = t[32083] ^ n[32084];
assign t[32085] = t[32084] ^ n[32085];
assign t[32086] = t[32085] ^ n[32086];
assign t[32087] = t[32086] ^ n[32087];
assign t[32088] = t[32087] ^ n[32088];
assign t[32089] = t[32088] ^ n[32089];
assign t[32090] = t[32089] ^ n[32090];
assign t[32091] = t[32090] ^ n[32091];
assign t[32092] = t[32091] ^ n[32092];
assign t[32093] = t[32092] ^ n[32093];
assign t[32094] = t[32093] ^ n[32094];
assign t[32095] = t[32094] ^ n[32095];
assign t[32096] = t[32095] ^ n[32096];
assign t[32097] = t[32096] ^ n[32097];
assign t[32098] = t[32097] ^ n[32098];
assign t[32099] = t[32098] ^ n[32099];
assign t[32100] = t[32099] ^ n[32100];
assign t[32101] = t[32100] ^ n[32101];
assign t[32102] = t[32101] ^ n[32102];
assign t[32103] = t[32102] ^ n[32103];
assign t[32104] = t[32103] ^ n[32104];
assign t[32105] = t[32104] ^ n[32105];
assign t[32106] = t[32105] ^ n[32106];
assign t[32107] = t[32106] ^ n[32107];
assign t[32108] = t[32107] ^ n[32108];
assign t[32109] = t[32108] ^ n[32109];
assign t[32110] = t[32109] ^ n[32110];
assign t[32111] = t[32110] ^ n[32111];
assign t[32112] = t[32111] ^ n[32112];
assign t[32113] = t[32112] ^ n[32113];
assign t[32114] = t[32113] ^ n[32114];
assign t[32115] = t[32114] ^ n[32115];
assign t[32116] = t[32115] ^ n[32116];
assign t[32117] = t[32116] ^ n[32117];
assign t[32118] = t[32117] ^ n[32118];
assign t[32119] = t[32118] ^ n[32119];
assign t[32120] = t[32119] ^ n[32120];
assign t[32121] = t[32120] ^ n[32121];
assign t[32122] = t[32121] ^ n[32122];
assign t[32123] = t[32122] ^ n[32123];
assign t[32124] = t[32123] ^ n[32124];
assign t[32125] = t[32124] ^ n[32125];
assign t[32126] = t[32125] ^ n[32126];
assign t[32127] = t[32126] ^ n[32127];
assign t[32128] = t[32127] ^ n[32128];
assign t[32129] = t[32128] ^ n[32129];
assign t[32130] = t[32129] ^ n[32130];
assign t[32131] = t[32130] ^ n[32131];
assign t[32132] = t[32131] ^ n[32132];
assign t[32133] = t[32132] ^ n[32133];
assign t[32134] = t[32133] ^ n[32134];
assign t[32135] = t[32134] ^ n[32135];
assign t[32136] = t[32135] ^ n[32136];
assign t[32137] = t[32136] ^ n[32137];
assign t[32138] = t[32137] ^ n[32138];
assign t[32139] = t[32138] ^ n[32139];
assign t[32140] = t[32139] ^ n[32140];
assign t[32141] = t[32140] ^ n[32141];
assign t[32142] = t[32141] ^ n[32142];
assign t[32143] = t[32142] ^ n[32143];
assign t[32144] = t[32143] ^ n[32144];
assign t[32145] = t[32144] ^ n[32145];
assign t[32146] = t[32145] ^ n[32146];
assign t[32147] = t[32146] ^ n[32147];
assign t[32148] = t[32147] ^ n[32148];
assign t[32149] = t[32148] ^ n[32149];
assign t[32150] = t[32149] ^ n[32150];
assign t[32151] = t[32150] ^ n[32151];
assign t[32152] = t[32151] ^ n[32152];
assign t[32153] = t[32152] ^ n[32153];
assign t[32154] = t[32153] ^ n[32154];
assign t[32155] = t[32154] ^ n[32155];
assign t[32156] = t[32155] ^ n[32156];
assign t[32157] = t[32156] ^ n[32157];
assign t[32158] = t[32157] ^ n[32158];
assign t[32159] = t[32158] ^ n[32159];
assign t[32160] = t[32159] ^ n[32160];
assign t[32161] = t[32160] ^ n[32161];
assign t[32162] = t[32161] ^ n[32162];
assign t[32163] = t[32162] ^ n[32163];
assign t[32164] = t[32163] ^ n[32164];
assign t[32165] = t[32164] ^ n[32165];
assign t[32166] = t[32165] ^ n[32166];
assign t[32167] = t[32166] ^ n[32167];
assign t[32168] = t[32167] ^ n[32168];
assign t[32169] = t[32168] ^ n[32169];
assign t[32170] = t[32169] ^ n[32170];
assign t[32171] = t[32170] ^ n[32171];
assign t[32172] = t[32171] ^ n[32172];
assign t[32173] = t[32172] ^ n[32173];
assign t[32174] = t[32173] ^ n[32174];
assign t[32175] = t[32174] ^ n[32175];
assign t[32176] = t[32175] ^ n[32176];
assign t[32177] = t[32176] ^ n[32177];
assign t[32178] = t[32177] ^ n[32178];
assign t[32179] = t[32178] ^ n[32179];
assign t[32180] = t[32179] ^ n[32180];
assign t[32181] = t[32180] ^ n[32181];
assign t[32182] = t[32181] ^ n[32182];
assign t[32183] = t[32182] ^ n[32183];
assign t[32184] = t[32183] ^ n[32184];
assign t[32185] = t[32184] ^ n[32185];
assign t[32186] = t[32185] ^ n[32186];
assign t[32187] = t[32186] ^ n[32187];
assign t[32188] = t[32187] ^ n[32188];
assign t[32189] = t[32188] ^ n[32189];
assign t[32190] = t[32189] ^ n[32190];
assign t[32191] = t[32190] ^ n[32191];
assign t[32192] = t[32191] ^ n[32192];
assign t[32193] = t[32192] ^ n[32193];
assign t[32194] = t[32193] ^ n[32194];
assign t[32195] = t[32194] ^ n[32195];
assign t[32196] = t[32195] ^ n[32196];
assign t[32197] = t[32196] ^ n[32197];
assign t[32198] = t[32197] ^ n[32198];
assign t[32199] = t[32198] ^ n[32199];
assign t[32200] = t[32199] ^ n[32200];
assign t[32201] = t[32200] ^ n[32201];
assign t[32202] = t[32201] ^ n[32202];
assign t[32203] = t[32202] ^ n[32203];
assign t[32204] = t[32203] ^ n[32204];
assign t[32205] = t[32204] ^ n[32205];
assign t[32206] = t[32205] ^ n[32206];
assign t[32207] = t[32206] ^ n[32207];
assign t[32208] = t[32207] ^ n[32208];
assign t[32209] = t[32208] ^ n[32209];
assign t[32210] = t[32209] ^ n[32210];
assign t[32211] = t[32210] ^ n[32211];
assign t[32212] = t[32211] ^ n[32212];
assign t[32213] = t[32212] ^ n[32213];
assign t[32214] = t[32213] ^ n[32214];
assign t[32215] = t[32214] ^ n[32215];
assign t[32216] = t[32215] ^ n[32216];
assign t[32217] = t[32216] ^ n[32217];
assign t[32218] = t[32217] ^ n[32218];
assign t[32219] = t[32218] ^ n[32219];
assign t[32220] = t[32219] ^ n[32220];
assign t[32221] = t[32220] ^ n[32221];
assign t[32222] = t[32221] ^ n[32222];
assign t[32223] = t[32222] ^ n[32223];
assign t[32224] = t[32223] ^ n[32224];
assign t[32225] = t[32224] ^ n[32225];
assign t[32226] = t[32225] ^ n[32226];
assign t[32227] = t[32226] ^ n[32227];
assign t[32228] = t[32227] ^ n[32228];
assign t[32229] = t[32228] ^ n[32229];
assign t[32230] = t[32229] ^ n[32230];
assign t[32231] = t[32230] ^ n[32231];
assign t[32232] = t[32231] ^ n[32232];
assign t[32233] = t[32232] ^ n[32233];
assign t[32234] = t[32233] ^ n[32234];
assign t[32235] = t[32234] ^ n[32235];
assign t[32236] = t[32235] ^ n[32236];
assign t[32237] = t[32236] ^ n[32237];
assign t[32238] = t[32237] ^ n[32238];
assign t[32239] = t[32238] ^ n[32239];
assign t[32240] = t[32239] ^ n[32240];
assign t[32241] = t[32240] ^ n[32241];
assign t[32242] = t[32241] ^ n[32242];
assign t[32243] = t[32242] ^ n[32243];
assign t[32244] = t[32243] ^ n[32244];
assign t[32245] = t[32244] ^ n[32245];
assign t[32246] = t[32245] ^ n[32246];
assign t[32247] = t[32246] ^ n[32247];
assign t[32248] = t[32247] ^ n[32248];
assign t[32249] = t[32248] ^ n[32249];
assign t[32250] = t[32249] ^ n[32250];
assign t[32251] = t[32250] ^ n[32251];
assign t[32252] = t[32251] ^ n[32252];
assign t[32253] = t[32252] ^ n[32253];
assign t[32254] = t[32253] ^ n[32254];
assign t[32255] = t[32254] ^ n[32255];
assign t[32256] = t[32255] ^ n[32256];
assign t[32257] = t[32256] ^ n[32257];
assign t[32258] = t[32257] ^ n[32258];
assign t[32259] = t[32258] ^ n[32259];
assign t[32260] = t[32259] ^ n[32260];
assign t[32261] = t[32260] ^ n[32261];
assign t[32262] = t[32261] ^ n[32262];
assign t[32263] = t[32262] ^ n[32263];
assign t[32264] = t[32263] ^ n[32264];
assign t[32265] = t[32264] ^ n[32265];
assign t[32266] = t[32265] ^ n[32266];
assign t[32267] = t[32266] ^ n[32267];
assign t[32268] = t[32267] ^ n[32268];
assign t[32269] = t[32268] ^ n[32269];
assign t[32270] = t[32269] ^ n[32270];
assign t[32271] = t[32270] ^ n[32271];
assign t[32272] = t[32271] ^ n[32272];
assign t[32273] = t[32272] ^ n[32273];
assign t[32274] = t[32273] ^ n[32274];
assign t[32275] = t[32274] ^ n[32275];
assign t[32276] = t[32275] ^ n[32276];
assign t[32277] = t[32276] ^ n[32277];
assign t[32278] = t[32277] ^ n[32278];
assign t[32279] = t[32278] ^ n[32279];
assign t[32280] = t[32279] ^ n[32280];
assign t[32281] = t[32280] ^ n[32281];
assign t[32282] = t[32281] ^ n[32282];
assign t[32283] = t[32282] ^ n[32283];
assign t[32284] = t[32283] ^ n[32284];
assign t[32285] = t[32284] ^ n[32285];
assign t[32286] = t[32285] ^ n[32286];
assign t[32287] = t[32286] ^ n[32287];
assign t[32288] = t[32287] ^ n[32288];
assign t[32289] = t[32288] ^ n[32289];
assign t[32290] = t[32289] ^ n[32290];
assign t[32291] = t[32290] ^ n[32291];
assign t[32292] = t[32291] ^ n[32292];
assign t[32293] = t[32292] ^ n[32293];
assign t[32294] = t[32293] ^ n[32294];
assign t[32295] = t[32294] ^ n[32295];
assign t[32296] = t[32295] ^ n[32296];
assign t[32297] = t[32296] ^ n[32297];
assign t[32298] = t[32297] ^ n[32298];
assign t[32299] = t[32298] ^ n[32299];
assign t[32300] = t[32299] ^ n[32300];
assign t[32301] = t[32300] ^ n[32301];
assign t[32302] = t[32301] ^ n[32302];
assign t[32303] = t[32302] ^ n[32303];
assign t[32304] = t[32303] ^ n[32304];
assign t[32305] = t[32304] ^ n[32305];
assign t[32306] = t[32305] ^ n[32306];
assign t[32307] = t[32306] ^ n[32307];
assign t[32308] = t[32307] ^ n[32308];
assign t[32309] = t[32308] ^ n[32309];
assign t[32310] = t[32309] ^ n[32310];
assign t[32311] = t[32310] ^ n[32311];
assign t[32312] = t[32311] ^ n[32312];
assign t[32313] = t[32312] ^ n[32313];
assign t[32314] = t[32313] ^ n[32314];
assign t[32315] = t[32314] ^ n[32315];
assign t[32316] = t[32315] ^ n[32316];
assign t[32317] = t[32316] ^ n[32317];
assign t[32318] = t[32317] ^ n[32318];
assign t[32319] = t[32318] ^ n[32319];
assign t[32320] = t[32319] ^ n[32320];
assign t[32321] = t[32320] ^ n[32321];
assign t[32322] = t[32321] ^ n[32322];
assign t[32323] = t[32322] ^ n[32323];
assign t[32324] = t[32323] ^ n[32324];
assign t[32325] = t[32324] ^ n[32325];
assign t[32326] = t[32325] ^ n[32326];
assign t[32327] = t[32326] ^ n[32327];
assign t[32328] = t[32327] ^ n[32328];
assign t[32329] = t[32328] ^ n[32329];
assign t[32330] = t[32329] ^ n[32330];
assign t[32331] = t[32330] ^ n[32331];
assign t[32332] = t[32331] ^ n[32332];
assign t[32333] = t[32332] ^ n[32333];
assign t[32334] = t[32333] ^ n[32334];
assign t[32335] = t[32334] ^ n[32335];
assign t[32336] = t[32335] ^ n[32336];
assign t[32337] = t[32336] ^ n[32337];
assign t[32338] = t[32337] ^ n[32338];
assign t[32339] = t[32338] ^ n[32339];
assign t[32340] = t[32339] ^ n[32340];
assign t[32341] = t[32340] ^ n[32341];
assign t[32342] = t[32341] ^ n[32342];
assign t[32343] = t[32342] ^ n[32343];
assign t[32344] = t[32343] ^ n[32344];
assign t[32345] = t[32344] ^ n[32345];
assign t[32346] = t[32345] ^ n[32346];
assign t[32347] = t[32346] ^ n[32347];
assign t[32348] = t[32347] ^ n[32348];
assign t[32349] = t[32348] ^ n[32349];
assign t[32350] = t[32349] ^ n[32350];
assign t[32351] = t[32350] ^ n[32351];
assign t[32352] = t[32351] ^ n[32352];
assign t[32353] = t[32352] ^ n[32353];
assign t[32354] = t[32353] ^ n[32354];
assign t[32355] = t[32354] ^ n[32355];
assign t[32356] = t[32355] ^ n[32356];
assign t[32357] = t[32356] ^ n[32357];
assign t[32358] = t[32357] ^ n[32358];
assign t[32359] = t[32358] ^ n[32359];
assign t[32360] = t[32359] ^ n[32360];
assign t[32361] = t[32360] ^ n[32361];
assign t[32362] = t[32361] ^ n[32362];
assign t[32363] = t[32362] ^ n[32363];
assign t[32364] = t[32363] ^ n[32364];
assign t[32365] = t[32364] ^ n[32365];
assign t[32366] = t[32365] ^ n[32366];
assign t[32367] = t[32366] ^ n[32367];
assign t[32368] = t[32367] ^ n[32368];
assign t[32369] = t[32368] ^ n[32369];
assign t[32370] = t[32369] ^ n[32370];
assign t[32371] = t[32370] ^ n[32371];
assign t[32372] = t[32371] ^ n[32372];
assign t[32373] = t[32372] ^ n[32373];
assign t[32374] = t[32373] ^ n[32374];
assign t[32375] = t[32374] ^ n[32375];
assign t[32376] = t[32375] ^ n[32376];
assign t[32377] = t[32376] ^ n[32377];
assign t[32378] = t[32377] ^ n[32378];
assign t[32379] = t[32378] ^ n[32379];
assign t[32380] = t[32379] ^ n[32380];
assign t[32381] = t[32380] ^ n[32381];
assign t[32382] = t[32381] ^ n[32382];
assign t[32383] = t[32382] ^ n[32383];
assign t[32384] = t[32383] ^ n[32384];
assign t[32385] = t[32384] ^ n[32385];
assign t[32386] = t[32385] ^ n[32386];
assign t[32387] = t[32386] ^ n[32387];
assign t[32388] = t[32387] ^ n[32388];
assign t[32389] = t[32388] ^ n[32389];
assign t[32390] = t[32389] ^ n[32390];
assign t[32391] = t[32390] ^ n[32391];
assign t[32392] = t[32391] ^ n[32392];
assign t[32393] = t[32392] ^ n[32393];
assign t[32394] = t[32393] ^ n[32394];
assign t[32395] = t[32394] ^ n[32395];
assign t[32396] = t[32395] ^ n[32396];
assign t[32397] = t[32396] ^ n[32397];
assign t[32398] = t[32397] ^ n[32398];
assign t[32399] = t[32398] ^ n[32399];
assign t[32400] = t[32399] ^ n[32400];
assign t[32401] = t[32400] ^ n[32401];
assign t[32402] = t[32401] ^ n[32402];
assign t[32403] = t[32402] ^ n[32403];
assign t[32404] = t[32403] ^ n[32404];
assign t[32405] = t[32404] ^ n[32405];
assign t[32406] = t[32405] ^ n[32406];
assign t[32407] = t[32406] ^ n[32407];
assign t[32408] = t[32407] ^ n[32408];
assign t[32409] = t[32408] ^ n[32409];
assign t[32410] = t[32409] ^ n[32410];
assign t[32411] = t[32410] ^ n[32411];
assign t[32412] = t[32411] ^ n[32412];
assign t[32413] = t[32412] ^ n[32413];
assign t[32414] = t[32413] ^ n[32414];
assign t[32415] = t[32414] ^ n[32415];
assign t[32416] = t[32415] ^ n[32416];
assign t[32417] = t[32416] ^ n[32417];
assign t[32418] = t[32417] ^ n[32418];
assign t[32419] = t[32418] ^ n[32419];
assign t[32420] = t[32419] ^ n[32420];
assign t[32421] = t[32420] ^ n[32421];
assign t[32422] = t[32421] ^ n[32422];
assign t[32423] = t[32422] ^ n[32423];
assign t[32424] = t[32423] ^ n[32424];
assign t[32425] = t[32424] ^ n[32425];
assign t[32426] = t[32425] ^ n[32426];
assign t[32427] = t[32426] ^ n[32427];
assign t[32428] = t[32427] ^ n[32428];
assign t[32429] = t[32428] ^ n[32429];
assign t[32430] = t[32429] ^ n[32430];
assign t[32431] = t[32430] ^ n[32431];
assign t[32432] = t[32431] ^ n[32432];
assign t[32433] = t[32432] ^ n[32433];
assign t[32434] = t[32433] ^ n[32434];
assign t[32435] = t[32434] ^ n[32435];
assign t[32436] = t[32435] ^ n[32436];
assign t[32437] = t[32436] ^ n[32437];
assign t[32438] = t[32437] ^ n[32438];
assign t[32439] = t[32438] ^ n[32439];
assign t[32440] = t[32439] ^ n[32440];
assign t[32441] = t[32440] ^ n[32441];
assign t[32442] = t[32441] ^ n[32442];
assign t[32443] = t[32442] ^ n[32443];
assign t[32444] = t[32443] ^ n[32444];
assign t[32445] = t[32444] ^ n[32445];
assign t[32446] = t[32445] ^ n[32446];
assign t[32447] = t[32446] ^ n[32447];
assign t[32448] = t[32447] ^ n[32448];
assign t[32449] = t[32448] ^ n[32449];
assign t[32450] = t[32449] ^ n[32450];
assign t[32451] = t[32450] ^ n[32451];
assign t[32452] = t[32451] ^ n[32452];
assign t[32453] = t[32452] ^ n[32453];
assign t[32454] = t[32453] ^ n[32454];
assign t[32455] = t[32454] ^ n[32455];
assign t[32456] = t[32455] ^ n[32456];
assign t[32457] = t[32456] ^ n[32457];
assign t[32458] = t[32457] ^ n[32458];
assign t[32459] = t[32458] ^ n[32459];
assign t[32460] = t[32459] ^ n[32460];
assign t[32461] = t[32460] ^ n[32461];
assign t[32462] = t[32461] ^ n[32462];
assign t[32463] = t[32462] ^ n[32463];
assign t[32464] = t[32463] ^ n[32464];
assign t[32465] = t[32464] ^ n[32465];
assign t[32466] = t[32465] ^ n[32466];
assign t[32467] = t[32466] ^ n[32467];
assign t[32468] = t[32467] ^ n[32468];
assign t[32469] = t[32468] ^ n[32469];
assign t[32470] = t[32469] ^ n[32470];
assign t[32471] = t[32470] ^ n[32471];
assign t[32472] = t[32471] ^ n[32472];
assign t[32473] = t[32472] ^ n[32473];
assign t[32474] = t[32473] ^ n[32474];
assign t[32475] = t[32474] ^ n[32475];
assign t[32476] = t[32475] ^ n[32476];
assign t[32477] = t[32476] ^ n[32477];
assign t[32478] = t[32477] ^ n[32478];
assign t[32479] = t[32478] ^ n[32479];
assign t[32480] = t[32479] ^ n[32480];
assign t[32481] = t[32480] ^ n[32481];
assign t[32482] = t[32481] ^ n[32482];
assign t[32483] = t[32482] ^ n[32483];
assign t[32484] = t[32483] ^ n[32484];
assign t[32485] = t[32484] ^ n[32485];
assign t[32486] = t[32485] ^ n[32486];
assign t[32487] = t[32486] ^ n[32487];
assign t[32488] = t[32487] ^ n[32488];
assign t[32489] = t[32488] ^ n[32489];
assign t[32490] = t[32489] ^ n[32490];
assign t[32491] = t[32490] ^ n[32491];
assign t[32492] = t[32491] ^ n[32492];
assign t[32493] = t[32492] ^ n[32493];
assign t[32494] = t[32493] ^ n[32494];
assign t[32495] = t[32494] ^ n[32495];
assign t[32496] = t[32495] ^ n[32496];
assign t[32497] = t[32496] ^ n[32497];
assign t[32498] = t[32497] ^ n[32498];
assign t[32499] = t[32498] ^ n[32499];
assign t[32500] = t[32499] ^ n[32500];
assign t[32501] = t[32500] ^ n[32501];
assign t[32502] = t[32501] ^ n[32502];
assign t[32503] = t[32502] ^ n[32503];
assign t[32504] = t[32503] ^ n[32504];
assign t[32505] = t[32504] ^ n[32505];
assign t[32506] = t[32505] ^ n[32506];
assign t[32507] = t[32506] ^ n[32507];
assign t[32508] = t[32507] ^ n[32508];
assign t[32509] = t[32508] ^ n[32509];
assign t[32510] = t[32509] ^ n[32510];
assign t[32511] = t[32510] ^ n[32511];
assign t[32512] = t[32511] ^ n[32512];
assign t[32513] = t[32512] ^ n[32513];
assign t[32514] = t[32513] ^ n[32514];
assign t[32515] = t[32514] ^ n[32515];
assign t[32516] = t[32515] ^ n[32516];
assign t[32517] = t[32516] ^ n[32517];
assign t[32518] = t[32517] ^ n[32518];
assign t[32519] = t[32518] ^ n[32519];
assign t[32520] = t[32519] ^ n[32520];
assign t[32521] = t[32520] ^ n[32521];
assign t[32522] = t[32521] ^ n[32522];
assign t[32523] = t[32522] ^ n[32523];
assign t[32524] = t[32523] ^ n[32524];
assign t[32525] = t[32524] ^ n[32525];
assign t[32526] = t[32525] ^ n[32526];
assign t[32527] = t[32526] ^ n[32527];
assign t[32528] = t[32527] ^ n[32528];
assign t[32529] = t[32528] ^ n[32529];
assign t[32530] = t[32529] ^ n[32530];
assign t[32531] = t[32530] ^ n[32531];
assign t[32532] = t[32531] ^ n[32532];
assign t[32533] = t[32532] ^ n[32533];
assign t[32534] = t[32533] ^ n[32534];
assign t[32535] = t[32534] ^ n[32535];
assign t[32536] = t[32535] ^ n[32536];
assign t[32537] = t[32536] ^ n[32537];
assign t[32538] = t[32537] ^ n[32538];
assign t[32539] = t[32538] ^ n[32539];
assign t[32540] = t[32539] ^ n[32540];
assign t[32541] = t[32540] ^ n[32541];
assign t[32542] = t[32541] ^ n[32542];
assign t[32543] = t[32542] ^ n[32543];
assign t[32544] = t[32543] ^ n[32544];
assign t[32545] = t[32544] ^ n[32545];
assign t[32546] = t[32545] ^ n[32546];
assign t[32547] = t[32546] ^ n[32547];
assign t[32548] = t[32547] ^ n[32548];
assign t[32549] = t[32548] ^ n[32549];
assign t[32550] = t[32549] ^ n[32550];
assign t[32551] = t[32550] ^ n[32551];
assign t[32552] = t[32551] ^ n[32552];
assign t[32553] = t[32552] ^ n[32553];
assign t[32554] = t[32553] ^ n[32554];
assign t[32555] = t[32554] ^ n[32555];
assign t[32556] = t[32555] ^ n[32556];
assign t[32557] = t[32556] ^ n[32557];
assign t[32558] = t[32557] ^ n[32558];
assign t[32559] = t[32558] ^ n[32559];
assign t[32560] = t[32559] ^ n[32560];
assign t[32561] = t[32560] ^ n[32561];
assign t[32562] = t[32561] ^ n[32562];
assign t[32563] = t[32562] ^ n[32563];
assign t[32564] = t[32563] ^ n[32564];
assign t[32565] = t[32564] ^ n[32565];
assign t[32566] = t[32565] ^ n[32566];
assign t[32567] = t[32566] ^ n[32567];
assign t[32568] = t[32567] ^ n[32568];
assign t[32569] = t[32568] ^ n[32569];
assign t[32570] = t[32569] ^ n[32570];
assign t[32571] = t[32570] ^ n[32571];
assign t[32572] = t[32571] ^ n[32572];
assign t[32573] = t[32572] ^ n[32573];
assign t[32574] = t[32573] ^ n[32574];
assign t[32575] = t[32574] ^ n[32575];
assign t[32576] = t[32575] ^ n[32576];
assign t[32577] = t[32576] ^ n[32577];
assign t[32578] = t[32577] ^ n[32578];
assign t[32579] = t[32578] ^ n[32579];
assign t[32580] = t[32579] ^ n[32580];
assign t[32581] = t[32580] ^ n[32581];
assign t[32582] = t[32581] ^ n[32582];
assign t[32583] = t[32582] ^ n[32583];
assign t[32584] = t[32583] ^ n[32584];
assign t[32585] = t[32584] ^ n[32585];
assign t[32586] = t[32585] ^ n[32586];
assign t[32587] = t[32586] ^ n[32587];
assign t[32588] = t[32587] ^ n[32588];
assign t[32589] = t[32588] ^ n[32589];
assign t[32590] = t[32589] ^ n[32590];
assign t[32591] = t[32590] ^ n[32591];
assign t[32592] = t[32591] ^ n[32592];
assign t[32593] = t[32592] ^ n[32593];
assign t[32594] = t[32593] ^ n[32594];
assign t[32595] = t[32594] ^ n[32595];
assign t[32596] = t[32595] ^ n[32596];
assign t[32597] = t[32596] ^ n[32597];
assign t[32598] = t[32597] ^ n[32598];
assign t[32599] = t[32598] ^ n[32599];
assign t[32600] = t[32599] ^ n[32600];
assign t[32601] = t[32600] ^ n[32601];
assign t[32602] = t[32601] ^ n[32602];
assign t[32603] = t[32602] ^ n[32603];
assign t[32604] = t[32603] ^ n[32604];
assign t[32605] = t[32604] ^ n[32605];
assign t[32606] = t[32605] ^ n[32606];
assign t[32607] = t[32606] ^ n[32607];
assign t[32608] = t[32607] ^ n[32608];
assign t[32609] = t[32608] ^ n[32609];
assign t[32610] = t[32609] ^ n[32610];
assign t[32611] = t[32610] ^ n[32611];
assign t[32612] = t[32611] ^ n[32612];
assign t[32613] = t[32612] ^ n[32613];
assign t[32614] = t[32613] ^ n[32614];
assign t[32615] = t[32614] ^ n[32615];
assign t[32616] = t[32615] ^ n[32616];
assign t[32617] = t[32616] ^ n[32617];
assign t[32618] = t[32617] ^ n[32618];
assign t[32619] = t[32618] ^ n[32619];
assign t[32620] = t[32619] ^ n[32620];
assign t[32621] = t[32620] ^ n[32621];
assign t[32622] = t[32621] ^ n[32622];
assign t[32623] = t[32622] ^ n[32623];
assign t[32624] = t[32623] ^ n[32624];
assign t[32625] = t[32624] ^ n[32625];
assign t[32626] = t[32625] ^ n[32626];
assign t[32627] = t[32626] ^ n[32627];
assign t[32628] = t[32627] ^ n[32628];
assign t[32629] = t[32628] ^ n[32629];
assign t[32630] = t[32629] ^ n[32630];
assign t[32631] = t[32630] ^ n[32631];
assign t[32632] = t[32631] ^ n[32632];
assign t[32633] = t[32632] ^ n[32633];
assign t[32634] = t[32633] ^ n[32634];
assign t[32635] = t[32634] ^ n[32635];
assign t[32636] = t[32635] ^ n[32636];
assign t[32637] = t[32636] ^ n[32637];
assign t[32638] = t[32637] ^ n[32638];
assign t[32639] = t[32638] ^ n[32639];
assign t[32640] = t[32639] ^ n[32640];
assign t[32641] = t[32640] ^ n[32641];
assign t[32642] = t[32641] ^ n[32642];
assign t[32643] = t[32642] ^ n[32643];
assign t[32644] = t[32643] ^ n[32644];
assign t[32645] = t[32644] ^ n[32645];
assign t[32646] = t[32645] ^ n[32646];
assign t[32647] = t[32646] ^ n[32647];
assign t[32648] = t[32647] ^ n[32648];
assign t[32649] = t[32648] ^ n[32649];
assign t[32650] = t[32649] ^ n[32650];
assign t[32651] = t[32650] ^ n[32651];
assign t[32652] = t[32651] ^ n[32652];
assign t[32653] = t[32652] ^ n[32653];
assign t[32654] = t[32653] ^ n[32654];
assign t[32655] = t[32654] ^ n[32655];
assign t[32656] = t[32655] ^ n[32656];
assign t[32657] = t[32656] ^ n[32657];
assign t[32658] = t[32657] ^ n[32658];
assign t[32659] = t[32658] ^ n[32659];
assign t[32660] = t[32659] ^ n[32660];
assign t[32661] = t[32660] ^ n[32661];
assign t[32662] = t[32661] ^ n[32662];
assign t[32663] = t[32662] ^ n[32663];
assign t[32664] = t[32663] ^ n[32664];
assign t[32665] = t[32664] ^ n[32665];
assign t[32666] = t[32665] ^ n[32666];
assign t[32667] = t[32666] ^ n[32667];
assign t[32668] = t[32667] ^ n[32668];
assign t[32669] = t[32668] ^ n[32669];
assign t[32670] = t[32669] ^ n[32670];
assign t[32671] = t[32670] ^ n[32671];
assign t[32672] = t[32671] ^ n[32672];
assign t[32673] = t[32672] ^ n[32673];
assign t[32674] = t[32673] ^ n[32674];
assign t[32675] = t[32674] ^ n[32675];
assign t[32676] = t[32675] ^ n[32676];
assign t[32677] = t[32676] ^ n[32677];
assign t[32678] = t[32677] ^ n[32678];
assign t[32679] = t[32678] ^ n[32679];
assign t[32680] = t[32679] ^ n[32680];
assign t[32681] = t[32680] ^ n[32681];
assign t[32682] = t[32681] ^ n[32682];
assign t[32683] = t[32682] ^ n[32683];
assign t[32684] = t[32683] ^ n[32684];
assign t[32685] = t[32684] ^ n[32685];
assign t[32686] = t[32685] ^ n[32686];
assign t[32687] = t[32686] ^ n[32687];
assign t[32688] = t[32687] ^ n[32688];
assign t[32689] = t[32688] ^ n[32689];
assign t[32690] = t[32689] ^ n[32690];
assign t[32691] = t[32690] ^ n[32691];
assign t[32692] = t[32691] ^ n[32692];
assign t[32693] = t[32692] ^ n[32693];
assign t[32694] = t[32693] ^ n[32694];
assign t[32695] = t[32694] ^ n[32695];
assign t[32696] = t[32695] ^ n[32696];
assign t[32697] = t[32696] ^ n[32697];
assign t[32698] = t[32697] ^ n[32698];
assign t[32699] = t[32698] ^ n[32699];
assign t[32700] = t[32699] ^ n[32700];
assign t[32701] = t[32700] ^ n[32701];
assign t[32702] = t[32701] ^ n[32702];
assign t[32703] = t[32702] ^ n[32703];
assign t[32704] = t[32703] ^ n[32704];
assign t[32705] = t[32704] ^ n[32705];
assign t[32706] = t[32705] ^ n[32706];
assign t[32707] = t[32706] ^ n[32707];
assign t[32708] = t[32707] ^ n[32708];
assign t[32709] = t[32708] ^ n[32709];
assign t[32710] = t[32709] ^ n[32710];
assign t[32711] = t[32710] ^ n[32711];
assign t[32712] = t[32711] ^ n[32712];
assign t[32713] = t[32712] ^ n[32713];
assign t[32714] = t[32713] ^ n[32714];
assign t[32715] = t[32714] ^ n[32715];
assign t[32716] = t[32715] ^ n[32716];
assign t[32717] = t[32716] ^ n[32717];
assign t[32718] = t[32717] ^ n[32718];
assign t[32719] = t[32718] ^ n[32719];
assign t[32720] = t[32719] ^ n[32720];
assign t[32721] = t[32720] ^ n[32721];
assign t[32722] = t[32721] ^ n[32722];
assign t[32723] = t[32722] ^ n[32723];
assign t[32724] = t[32723] ^ n[32724];
assign t[32725] = t[32724] ^ n[32725];
assign t[32726] = t[32725] ^ n[32726];
assign t[32727] = t[32726] ^ n[32727];
assign t[32728] = t[32727] ^ n[32728];
assign t[32729] = t[32728] ^ n[32729];
assign t[32730] = t[32729] ^ n[32730];
assign t[32731] = t[32730] ^ n[32731];
assign t[32732] = t[32731] ^ n[32732];
assign t[32733] = t[32732] ^ n[32733];
assign t[32734] = t[32733] ^ n[32734];
assign t[32735] = t[32734] ^ n[32735];
assign t[32736] = t[32735] ^ n[32736];
assign t[32737] = t[32736] ^ n[32737];
assign t[32738] = t[32737] ^ n[32738];
assign t[32739] = t[32738] ^ n[32739];
assign t[32740] = t[32739] ^ n[32740];
assign t[32741] = t[32740] ^ n[32741];
assign t[32742] = t[32741] ^ n[32742];
assign t[32743] = t[32742] ^ n[32743];
assign t[32744] = t[32743] ^ n[32744];
assign t[32745] = t[32744] ^ n[32745];
assign t[32746] = t[32745] ^ n[32746];
assign t[32747] = t[32746] ^ n[32747];
assign t[32748] = t[32747] ^ n[32748];
assign t[32749] = t[32748] ^ n[32749];
assign t[32750] = t[32749] ^ n[32750];
assign t[32751] = t[32750] ^ n[32751];

//asigning bit 14
assign s[14] = ( a[14] ^ b [14] ) ^ t[32751];

assign t[32752] = n[32752];
assign t[32753] = t[32752] ^ n[32753];
assign t[32754] = t[32753] ^ n[32754];
assign t[32755] = t[32754] ^ n[32755];
assign t[32756] = t[32755] ^ n[32756];
assign t[32757] = t[32756] ^ n[32757];
assign t[32758] = t[32757] ^ n[32758];
assign t[32759] = t[32758] ^ n[32759];
assign t[32760] = t[32759] ^ n[32760];
assign t[32761] = t[32760] ^ n[32761];
assign t[32762] = t[32761] ^ n[32762];
assign t[32763] = t[32762] ^ n[32763];
assign t[32764] = t[32763] ^ n[32764];
assign t[32765] = t[32764] ^ n[32765];
assign t[32766] = t[32765] ^ n[32766];
assign t[32767] = t[32766] ^ n[32767];
assign t[32768] = t[32767] ^ n[32768];
assign t[32769] = t[32768] ^ n[32769];
assign t[32770] = t[32769] ^ n[32770];
assign t[32771] = t[32770] ^ n[32771];
assign t[32772] = t[32771] ^ n[32772];
assign t[32773] = t[32772] ^ n[32773];
assign t[32774] = t[32773] ^ n[32774];
assign t[32775] = t[32774] ^ n[32775];
assign t[32776] = t[32775] ^ n[32776];
assign t[32777] = t[32776] ^ n[32777];
assign t[32778] = t[32777] ^ n[32778];
assign t[32779] = t[32778] ^ n[32779];
assign t[32780] = t[32779] ^ n[32780];
assign t[32781] = t[32780] ^ n[32781];
assign t[32782] = t[32781] ^ n[32782];
assign t[32783] = t[32782] ^ n[32783];
assign t[32784] = t[32783] ^ n[32784];
assign t[32785] = t[32784] ^ n[32785];
assign t[32786] = t[32785] ^ n[32786];
assign t[32787] = t[32786] ^ n[32787];
assign t[32788] = t[32787] ^ n[32788];
assign t[32789] = t[32788] ^ n[32789];
assign t[32790] = t[32789] ^ n[32790];
assign t[32791] = t[32790] ^ n[32791];
assign t[32792] = t[32791] ^ n[32792];
assign t[32793] = t[32792] ^ n[32793];
assign t[32794] = t[32793] ^ n[32794];
assign t[32795] = t[32794] ^ n[32795];
assign t[32796] = t[32795] ^ n[32796];
assign t[32797] = t[32796] ^ n[32797];
assign t[32798] = t[32797] ^ n[32798];
assign t[32799] = t[32798] ^ n[32799];
assign t[32800] = t[32799] ^ n[32800];
assign t[32801] = t[32800] ^ n[32801];
assign t[32802] = t[32801] ^ n[32802];
assign t[32803] = t[32802] ^ n[32803];
assign t[32804] = t[32803] ^ n[32804];
assign t[32805] = t[32804] ^ n[32805];
assign t[32806] = t[32805] ^ n[32806];
assign t[32807] = t[32806] ^ n[32807];
assign t[32808] = t[32807] ^ n[32808];
assign t[32809] = t[32808] ^ n[32809];
assign t[32810] = t[32809] ^ n[32810];
assign t[32811] = t[32810] ^ n[32811];
assign t[32812] = t[32811] ^ n[32812];
assign t[32813] = t[32812] ^ n[32813];
assign t[32814] = t[32813] ^ n[32814];
assign t[32815] = t[32814] ^ n[32815];
assign t[32816] = t[32815] ^ n[32816];
assign t[32817] = t[32816] ^ n[32817];
assign t[32818] = t[32817] ^ n[32818];
assign t[32819] = t[32818] ^ n[32819];
assign t[32820] = t[32819] ^ n[32820];
assign t[32821] = t[32820] ^ n[32821];
assign t[32822] = t[32821] ^ n[32822];
assign t[32823] = t[32822] ^ n[32823];
assign t[32824] = t[32823] ^ n[32824];
assign t[32825] = t[32824] ^ n[32825];
assign t[32826] = t[32825] ^ n[32826];
assign t[32827] = t[32826] ^ n[32827];
assign t[32828] = t[32827] ^ n[32828];
assign t[32829] = t[32828] ^ n[32829];
assign t[32830] = t[32829] ^ n[32830];
assign t[32831] = t[32830] ^ n[32831];
assign t[32832] = t[32831] ^ n[32832];
assign t[32833] = t[32832] ^ n[32833];
assign t[32834] = t[32833] ^ n[32834];
assign t[32835] = t[32834] ^ n[32835];
assign t[32836] = t[32835] ^ n[32836];
assign t[32837] = t[32836] ^ n[32837];
assign t[32838] = t[32837] ^ n[32838];
assign t[32839] = t[32838] ^ n[32839];
assign t[32840] = t[32839] ^ n[32840];
assign t[32841] = t[32840] ^ n[32841];
assign t[32842] = t[32841] ^ n[32842];
assign t[32843] = t[32842] ^ n[32843];
assign t[32844] = t[32843] ^ n[32844];
assign t[32845] = t[32844] ^ n[32845];
assign t[32846] = t[32845] ^ n[32846];
assign t[32847] = t[32846] ^ n[32847];
assign t[32848] = t[32847] ^ n[32848];
assign t[32849] = t[32848] ^ n[32849];
assign t[32850] = t[32849] ^ n[32850];
assign t[32851] = t[32850] ^ n[32851];
assign t[32852] = t[32851] ^ n[32852];
assign t[32853] = t[32852] ^ n[32853];
assign t[32854] = t[32853] ^ n[32854];
assign t[32855] = t[32854] ^ n[32855];
assign t[32856] = t[32855] ^ n[32856];
assign t[32857] = t[32856] ^ n[32857];
assign t[32858] = t[32857] ^ n[32858];
assign t[32859] = t[32858] ^ n[32859];
assign t[32860] = t[32859] ^ n[32860];
assign t[32861] = t[32860] ^ n[32861];
assign t[32862] = t[32861] ^ n[32862];
assign t[32863] = t[32862] ^ n[32863];
assign t[32864] = t[32863] ^ n[32864];
assign t[32865] = t[32864] ^ n[32865];
assign t[32866] = t[32865] ^ n[32866];
assign t[32867] = t[32866] ^ n[32867];
assign t[32868] = t[32867] ^ n[32868];
assign t[32869] = t[32868] ^ n[32869];
assign t[32870] = t[32869] ^ n[32870];
assign t[32871] = t[32870] ^ n[32871];
assign t[32872] = t[32871] ^ n[32872];
assign t[32873] = t[32872] ^ n[32873];
assign t[32874] = t[32873] ^ n[32874];
assign t[32875] = t[32874] ^ n[32875];
assign t[32876] = t[32875] ^ n[32876];
assign t[32877] = t[32876] ^ n[32877];
assign t[32878] = t[32877] ^ n[32878];
assign t[32879] = t[32878] ^ n[32879];
assign t[32880] = t[32879] ^ n[32880];
assign t[32881] = t[32880] ^ n[32881];
assign t[32882] = t[32881] ^ n[32882];
assign t[32883] = t[32882] ^ n[32883];
assign t[32884] = t[32883] ^ n[32884];
assign t[32885] = t[32884] ^ n[32885];
assign t[32886] = t[32885] ^ n[32886];
assign t[32887] = t[32886] ^ n[32887];
assign t[32888] = t[32887] ^ n[32888];
assign t[32889] = t[32888] ^ n[32889];
assign t[32890] = t[32889] ^ n[32890];
assign t[32891] = t[32890] ^ n[32891];
assign t[32892] = t[32891] ^ n[32892];
assign t[32893] = t[32892] ^ n[32893];
assign t[32894] = t[32893] ^ n[32894];
assign t[32895] = t[32894] ^ n[32895];
assign t[32896] = t[32895] ^ n[32896];
assign t[32897] = t[32896] ^ n[32897];
assign t[32898] = t[32897] ^ n[32898];
assign t[32899] = t[32898] ^ n[32899];
assign t[32900] = t[32899] ^ n[32900];
assign t[32901] = t[32900] ^ n[32901];
assign t[32902] = t[32901] ^ n[32902];
assign t[32903] = t[32902] ^ n[32903];
assign t[32904] = t[32903] ^ n[32904];
assign t[32905] = t[32904] ^ n[32905];
assign t[32906] = t[32905] ^ n[32906];
assign t[32907] = t[32906] ^ n[32907];
assign t[32908] = t[32907] ^ n[32908];
assign t[32909] = t[32908] ^ n[32909];
assign t[32910] = t[32909] ^ n[32910];
assign t[32911] = t[32910] ^ n[32911];
assign t[32912] = t[32911] ^ n[32912];
assign t[32913] = t[32912] ^ n[32913];
assign t[32914] = t[32913] ^ n[32914];
assign t[32915] = t[32914] ^ n[32915];
assign t[32916] = t[32915] ^ n[32916];
assign t[32917] = t[32916] ^ n[32917];
assign t[32918] = t[32917] ^ n[32918];
assign t[32919] = t[32918] ^ n[32919];
assign t[32920] = t[32919] ^ n[32920];
assign t[32921] = t[32920] ^ n[32921];
assign t[32922] = t[32921] ^ n[32922];
assign t[32923] = t[32922] ^ n[32923];
assign t[32924] = t[32923] ^ n[32924];
assign t[32925] = t[32924] ^ n[32925];
assign t[32926] = t[32925] ^ n[32926];
assign t[32927] = t[32926] ^ n[32927];
assign t[32928] = t[32927] ^ n[32928];
assign t[32929] = t[32928] ^ n[32929];
assign t[32930] = t[32929] ^ n[32930];
assign t[32931] = t[32930] ^ n[32931];
assign t[32932] = t[32931] ^ n[32932];
assign t[32933] = t[32932] ^ n[32933];
assign t[32934] = t[32933] ^ n[32934];
assign t[32935] = t[32934] ^ n[32935];
assign t[32936] = t[32935] ^ n[32936];
assign t[32937] = t[32936] ^ n[32937];
assign t[32938] = t[32937] ^ n[32938];
assign t[32939] = t[32938] ^ n[32939];
assign t[32940] = t[32939] ^ n[32940];
assign t[32941] = t[32940] ^ n[32941];
assign t[32942] = t[32941] ^ n[32942];
assign t[32943] = t[32942] ^ n[32943];
assign t[32944] = t[32943] ^ n[32944];
assign t[32945] = t[32944] ^ n[32945];
assign t[32946] = t[32945] ^ n[32946];
assign t[32947] = t[32946] ^ n[32947];
assign t[32948] = t[32947] ^ n[32948];
assign t[32949] = t[32948] ^ n[32949];
assign t[32950] = t[32949] ^ n[32950];
assign t[32951] = t[32950] ^ n[32951];
assign t[32952] = t[32951] ^ n[32952];
assign t[32953] = t[32952] ^ n[32953];
assign t[32954] = t[32953] ^ n[32954];
assign t[32955] = t[32954] ^ n[32955];
assign t[32956] = t[32955] ^ n[32956];
assign t[32957] = t[32956] ^ n[32957];
assign t[32958] = t[32957] ^ n[32958];
assign t[32959] = t[32958] ^ n[32959];
assign t[32960] = t[32959] ^ n[32960];
assign t[32961] = t[32960] ^ n[32961];
assign t[32962] = t[32961] ^ n[32962];
assign t[32963] = t[32962] ^ n[32963];
assign t[32964] = t[32963] ^ n[32964];
assign t[32965] = t[32964] ^ n[32965];
assign t[32966] = t[32965] ^ n[32966];
assign t[32967] = t[32966] ^ n[32967];
assign t[32968] = t[32967] ^ n[32968];
assign t[32969] = t[32968] ^ n[32969];
assign t[32970] = t[32969] ^ n[32970];
assign t[32971] = t[32970] ^ n[32971];
assign t[32972] = t[32971] ^ n[32972];
assign t[32973] = t[32972] ^ n[32973];
assign t[32974] = t[32973] ^ n[32974];
assign t[32975] = t[32974] ^ n[32975];
assign t[32976] = t[32975] ^ n[32976];
assign t[32977] = t[32976] ^ n[32977];
assign t[32978] = t[32977] ^ n[32978];
assign t[32979] = t[32978] ^ n[32979];
assign t[32980] = t[32979] ^ n[32980];
assign t[32981] = t[32980] ^ n[32981];
assign t[32982] = t[32981] ^ n[32982];
assign t[32983] = t[32982] ^ n[32983];
assign t[32984] = t[32983] ^ n[32984];
assign t[32985] = t[32984] ^ n[32985];
assign t[32986] = t[32985] ^ n[32986];
assign t[32987] = t[32986] ^ n[32987];
assign t[32988] = t[32987] ^ n[32988];
assign t[32989] = t[32988] ^ n[32989];
assign t[32990] = t[32989] ^ n[32990];
assign t[32991] = t[32990] ^ n[32991];
assign t[32992] = t[32991] ^ n[32992];
assign t[32993] = t[32992] ^ n[32993];
assign t[32994] = t[32993] ^ n[32994];
assign t[32995] = t[32994] ^ n[32995];
assign t[32996] = t[32995] ^ n[32996];
assign t[32997] = t[32996] ^ n[32997];
assign t[32998] = t[32997] ^ n[32998];
assign t[32999] = t[32998] ^ n[32999];
assign t[33000] = t[32999] ^ n[33000];
assign t[33001] = t[33000] ^ n[33001];
assign t[33002] = t[33001] ^ n[33002];
assign t[33003] = t[33002] ^ n[33003];
assign t[33004] = t[33003] ^ n[33004];
assign t[33005] = t[33004] ^ n[33005];
assign t[33006] = t[33005] ^ n[33006];
assign t[33007] = t[33006] ^ n[33007];
assign t[33008] = t[33007] ^ n[33008];
assign t[33009] = t[33008] ^ n[33009];
assign t[33010] = t[33009] ^ n[33010];
assign t[33011] = t[33010] ^ n[33011];
assign t[33012] = t[33011] ^ n[33012];
assign t[33013] = t[33012] ^ n[33013];
assign t[33014] = t[33013] ^ n[33014];
assign t[33015] = t[33014] ^ n[33015];
assign t[33016] = t[33015] ^ n[33016];
assign t[33017] = t[33016] ^ n[33017];
assign t[33018] = t[33017] ^ n[33018];
assign t[33019] = t[33018] ^ n[33019];
assign t[33020] = t[33019] ^ n[33020];
assign t[33021] = t[33020] ^ n[33021];
assign t[33022] = t[33021] ^ n[33022];
assign t[33023] = t[33022] ^ n[33023];
assign t[33024] = t[33023] ^ n[33024];
assign t[33025] = t[33024] ^ n[33025];
assign t[33026] = t[33025] ^ n[33026];
assign t[33027] = t[33026] ^ n[33027];
assign t[33028] = t[33027] ^ n[33028];
assign t[33029] = t[33028] ^ n[33029];
assign t[33030] = t[33029] ^ n[33030];
assign t[33031] = t[33030] ^ n[33031];
assign t[33032] = t[33031] ^ n[33032];
assign t[33033] = t[33032] ^ n[33033];
assign t[33034] = t[33033] ^ n[33034];
assign t[33035] = t[33034] ^ n[33035];
assign t[33036] = t[33035] ^ n[33036];
assign t[33037] = t[33036] ^ n[33037];
assign t[33038] = t[33037] ^ n[33038];
assign t[33039] = t[33038] ^ n[33039];
assign t[33040] = t[33039] ^ n[33040];
assign t[33041] = t[33040] ^ n[33041];
assign t[33042] = t[33041] ^ n[33042];
assign t[33043] = t[33042] ^ n[33043];
assign t[33044] = t[33043] ^ n[33044];
assign t[33045] = t[33044] ^ n[33045];
assign t[33046] = t[33045] ^ n[33046];
assign t[33047] = t[33046] ^ n[33047];
assign t[33048] = t[33047] ^ n[33048];
assign t[33049] = t[33048] ^ n[33049];
assign t[33050] = t[33049] ^ n[33050];
assign t[33051] = t[33050] ^ n[33051];
assign t[33052] = t[33051] ^ n[33052];
assign t[33053] = t[33052] ^ n[33053];
assign t[33054] = t[33053] ^ n[33054];
assign t[33055] = t[33054] ^ n[33055];
assign t[33056] = t[33055] ^ n[33056];
assign t[33057] = t[33056] ^ n[33057];
assign t[33058] = t[33057] ^ n[33058];
assign t[33059] = t[33058] ^ n[33059];
assign t[33060] = t[33059] ^ n[33060];
assign t[33061] = t[33060] ^ n[33061];
assign t[33062] = t[33061] ^ n[33062];
assign t[33063] = t[33062] ^ n[33063];
assign t[33064] = t[33063] ^ n[33064];
assign t[33065] = t[33064] ^ n[33065];
assign t[33066] = t[33065] ^ n[33066];
assign t[33067] = t[33066] ^ n[33067];
assign t[33068] = t[33067] ^ n[33068];
assign t[33069] = t[33068] ^ n[33069];
assign t[33070] = t[33069] ^ n[33070];
assign t[33071] = t[33070] ^ n[33071];
assign t[33072] = t[33071] ^ n[33072];
assign t[33073] = t[33072] ^ n[33073];
assign t[33074] = t[33073] ^ n[33074];
assign t[33075] = t[33074] ^ n[33075];
assign t[33076] = t[33075] ^ n[33076];
assign t[33077] = t[33076] ^ n[33077];
assign t[33078] = t[33077] ^ n[33078];
assign t[33079] = t[33078] ^ n[33079];
assign t[33080] = t[33079] ^ n[33080];
assign t[33081] = t[33080] ^ n[33081];
assign t[33082] = t[33081] ^ n[33082];
assign t[33083] = t[33082] ^ n[33083];
assign t[33084] = t[33083] ^ n[33084];
assign t[33085] = t[33084] ^ n[33085];
assign t[33086] = t[33085] ^ n[33086];
assign t[33087] = t[33086] ^ n[33087];
assign t[33088] = t[33087] ^ n[33088];
assign t[33089] = t[33088] ^ n[33089];
assign t[33090] = t[33089] ^ n[33090];
assign t[33091] = t[33090] ^ n[33091];
assign t[33092] = t[33091] ^ n[33092];
assign t[33093] = t[33092] ^ n[33093];
assign t[33094] = t[33093] ^ n[33094];
assign t[33095] = t[33094] ^ n[33095];
assign t[33096] = t[33095] ^ n[33096];
assign t[33097] = t[33096] ^ n[33097];
assign t[33098] = t[33097] ^ n[33098];
assign t[33099] = t[33098] ^ n[33099];
assign t[33100] = t[33099] ^ n[33100];
assign t[33101] = t[33100] ^ n[33101];
assign t[33102] = t[33101] ^ n[33102];
assign t[33103] = t[33102] ^ n[33103];
assign t[33104] = t[33103] ^ n[33104];
assign t[33105] = t[33104] ^ n[33105];
assign t[33106] = t[33105] ^ n[33106];
assign t[33107] = t[33106] ^ n[33107];
assign t[33108] = t[33107] ^ n[33108];
assign t[33109] = t[33108] ^ n[33109];
assign t[33110] = t[33109] ^ n[33110];
assign t[33111] = t[33110] ^ n[33111];
assign t[33112] = t[33111] ^ n[33112];
assign t[33113] = t[33112] ^ n[33113];
assign t[33114] = t[33113] ^ n[33114];
assign t[33115] = t[33114] ^ n[33115];
assign t[33116] = t[33115] ^ n[33116];
assign t[33117] = t[33116] ^ n[33117];
assign t[33118] = t[33117] ^ n[33118];
assign t[33119] = t[33118] ^ n[33119];
assign t[33120] = t[33119] ^ n[33120];
assign t[33121] = t[33120] ^ n[33121];
assign t[33122] = t[33121] ^ n[33122];
assign t[33123] = t[33122] ^ n[33123];
assign t[33124] = t[33123] ^ n[33124];
assign t[33125] = t[33124] ^ n[33125];
assign t[33126] = t[33125] ^ n[33126];
assign t[33127] = t[33126] ^ n[33127];
assign t[33128] = t[33127] ^ n[33128];
assign t[33129] = t[33128] ^ n[33129];
assign t[33130] = t[33129] ^ n[33130];
assign t[33131] = t[33130] ^ n[33131];
assign t[33132] = t[33131] ^ n[33132];
assign t[33133] = t[33132] ^ n[33133];
assign t[33134] = t[33133] ^ n[33134];
assign t[33135] = t[33134] ^ n[33135];
assign t[33136] = t[33135] ^ n[33136];
assign t[33137] = t[33136] ^ n[33137];
assign t[33138] = t[33137] ^ n[33138];
assign t[33139] = t[33138] ^ n[33139];
assign t[33140] = t[33139] ^ n[33140];
assign t[33141] = t[33140] ^ n[33141];
assign t[33142] = t[33141] ^ n[33142];
assign t[33143] = t[33142] ^ n[33143];
assign t[33144] = t[33143] ^ n[33144];
assign t[33145] = t[33144] ^ n[33145];
assign t[33146] = t[33145] ^ n[33146];
assign t[33147] = t[33146] ^ n[33147];
assign t[33148] = t[33147] ^ n[33148];
assign t[33149] = t[33148] ^ n[33149];
assign t[33150] = t[33149] ^ n[33150];
assign t[33151] = t[33150] ^ n[33151];
assign t[33152] = t[33151] ^ n[33152];
assign t[33153] = t[33152] ^ n[33153];
assign t[33154] = t[33153] ^ n[33154];
assign t[33155] = t[33154] ^ n[33155];
assign t[33156] = t[33155] ^ n[33156];
assign t[33157] = t[33156] ^ n[33157];
assign t[33158] = t[33157] ^ n[33158];
assign t[33159] = t[33158] ^ n[33159];
assign t[33160] = t[33159] ^ n[33160];
assign t[33161] = t[33160] ^ n[33161];
assign t[33162] = t[33161] ^ n[33162];
assign t[33163] = t[33162] ^ n[33163];
assign t[33164] = t[33163] ^ n[33164];
assign t[33165] = t[33164] ^ n[33165];
assign t[33166] = t[33165] ^ n[33166];
assign t[33167] = t[33166] ^ n[33167];
assign t[33168] = t[33167] ^ n[33168];
assign t[33169] = t[33168] ^ n[33169];
assign t[33170] = t[33169] ^ n[33170];
assign t[33171] = t[33170] ^ n[33171];
assign t[33172] = t[33171] ^ n[33172];
assign t[33173] = t[33172] ^ n[33173];
assign t[33174] = t[33173] ^ n[33174];
assign t[33175] = t[33174] ^ n[33175];
assign t[33176] = t[33175] ^ n[33176];
assign t[33177] = t[33176] ^ n[33177];
assign t[33178] = t[33177] ^ n[33178];
assign t[33179] = t[33178] ^ n[33179];
assign t[33180] = t[33179] ^ n[33180];
assign t[33181] = t[33180] ^ n[33181];
assign t[33182] = t[33181] ^ n[33182];
assign t[33183] = t[33182] ^ n[33183];
assign t[33184] = t[33183] ^ n[33184];
assign t[33185] = t[33184] ^ n[33185];
assign t[33186] = t[33185] ^ n[33186];
assign t[33187] = t[33186] ^ n[33187];
assign t[33188] = t[33187] ^ n[33188];
assign t[33189] = t[33188] ^ n[33189];
assign t[33190] = t[33189] ^ n[33190];
assign t[33191] = t[33190] ^ n[33191];
assign t[33192] = t[33191] ^ n[33192];
assign t[33193] = t[33192] ^ n[33193];
assign t[33194] = t[33193] ^ n[33194];
assign t[33195] = t[33194] ^ n[33195];
assign t[33196] = t[33195] ^ n[33196];
assign t[33197] = t[33196] ^ n[33197];
assign t[33198] = t[33197] ^ n[33198];
assign t[33199] = t[33198] ^ n[33199];
assign t[33200] = t[33199] ^ n[33200];
assign t[33201] = t[33200] ^ n[33201];
assign t[33202] = t[33201] ^ n[33202];
assign t[33203] = t[33202] ^ n[33203];
assign t[33204] = t[33203] ^ n[33204];
assign t[33205] = t[33204] ^ n[33205];
assign t[33206] = t[33205] ^ n[33206];
assign t[33207] = t[33206] ^ n[33207];
assign t[33208] = t[33207] ^ n[33208];
assign t[33209] = t[33208] ^ n[33209];
assign t[33210] = t[33209] ^ n[33210];
assign t[33211] = t[33210] ^ n[33211];
assign t[33212] = t[33211] ^ n[33212];
assign t[33213] = t[33212] ^ n[33213];
assign t[33214] = t[33213] ^ n[33214];
assign t[33215] = t[33214] ^ n[33215];
assign t[33216] = t[33215] ^ n[33216];
assign t[33217] = t[33216] ^ n[33217];
assign t[33218] = t[33217] ^ n[33218];
assign t[33219] = t[33218] ^ n[33219];
assign t[33220] = t[33219] ^ n[33220];
assign t[33221] = t[33220] ^ n[33221];
assign t[33222] = t[33221] ^ n[33222];
assign t[33223] = t[33222] ^ n[33223];
assign t[33224] = t[33223] ^ n[33224];
assign t[33225] = t[33224] ^ n[33225];
assign t[33226] = t[33225] ^ n[33226];
assign t[33227] = t[33226] ^ n[33227];
assign t[33228] = t[33227] ^ n[33228];
assign t[33229] = t[33228] ^ n[33229];
assign t[33230] = t[33229] ^ n[33230];
assign t[33231] = t[33230] ^ n[33231];
assign t[33232] = t[33231] ^ n[33232];
assign t[33233] = t[33232] ^ n[33233];
assign t[33234] = t[33233] ^ n[33234];
assign t[33235] = t[33234] ^ n[33235];
assign t[33236] = t[33235] ^ n[33236];
assign t[33237] = t[33236] ^ n[33237];
assign t[33238] = t[33237] ^ n[33238];
assign t[33239] = t[33238] ^ n[33239];
assign t[33240] = t[33239] ^ n[33240];
assign t[33241] = t[33240] ^ n[33241];
assign t[33242] = t[33241] ^ n[33242];
assign t[33243] = t[33242] ^ n[33243];
assign t[33244] = t[33243] ^ n[33244];
assign t[33245] = t[33244] ^ n[33245];
assign t[33246] = t[33245] ^ n[33246];
assign t[33247] = t[33246] ^ n[33247];
assign t[33248] = t[33247] ^ n[33248];
assign t[33249] = t[33248] ^ n[33249];
assign t[33250] = t[33249] ^ n[33250];
assign t[33251] = t[33250] ^ n[33251];
assign t[33252] = t[33251] ^ n[33252];
assign t[33253] = t[33252] ^ n[33253];
assign t[33254] = t[33253] ^ n[33254];
assign t[33255] = t[33254] ^ n[33255];
assign t[33256] = t[33255] ^ n[33256];
assign t[33257] = t[33256] ^ n[33257];
assign t[33258] = t[33257] ^ n[33258];
assign t[33259] = t[33258] ^ n[33259];
assign t[33260] = t[33259] ^ n[33260];
assign t[33261] = t[33260] ^ n[33261];
assign t[33262] = t[33261] ^ n[33262];
assign t[33263] = t[33262] ^ n[33263];
assign t[33264] = t[33263] ^ n[33264];
assign t[33265] = t[33264] ^ n[33265];
assign t[33266] = t[33265] ^ n[33266];
assign t[33267] = t[33266] ^ n[33267];
assign t[33268] = t[33267] ^ n[33268];
assign t[33269] = t[33268] ^ n[33269];
assign t[33270] = t[33269] ^ n[33270];
assign t[33271] = t[33270] ^ n[33271];
assign t[33272] = t[33271] ^ n[33272];
assign t[33273] = t[33272] ^ n[33273];
assign t[33274] = t[33273] ^ n[33274];
assign t[33275] = t[33274] ^ n[33275];
assign t[33276] = t[33275] ^ n[33276];
assign t[33277] = t[33276] ^ n[33277];
assign t[33278] = t[33277] ^ n[33278];
assign t[33279] = t[33278] ^ n[33279];
assign t[33280] = t[33279] ^ n[33280];
assign t[33281] = t[33280] ^ n[33281];
assign t[33282] = t[33281] ^ n[33282];
assign t[33283] = t[33282] ^ n[33283];
assign t[33284] = t[33283] ^ n[33284];
assign t[33285] = t[33284] ^ n[33285];
assign t[33286] = t[33285] ^ n[33286];
assign t[33287] = t[33286] ^ n[33287];
assign t[33288] = t[33287] ^ n[33288];
assign t[33289] = t[33288] ^ n[33289];
assign t[33290] = t[33289] ^ n[33290];
assign t[33291] = t[33290] ^ n[33291];
assign t[33292] = t[33291] ^ n[33292];
assign t[33293] = t[33292] ^ n[33293];
assign t[33294] = t[33293] ^ n[33294];
assign t[33295] = t[33294] ^ n[33295];
assign t[33296] = t[33295] ^ n[33296];
assign t[33297] = t[33296] ^ n[33297];
assign t[33298] = t[33297] ^ n[33298];
assign t[33299] = t[33298] ^ n[33299];
assign t[33300] = t[33299] ^ n[33300];
assign t[33301] = t[33300] ^ n[33301];
assign t[33302] = t[33301] ^ n[33302];
assign t[33303] = t[33302] ^ n[33303];
assign t[33304] = t[33303] ^ n[33304];
assign t[33305] = t[33304] ^ n[33305];
assign t[33306] = t[33305] ^ n[33306];
assign t[33307] = t[33306] ^ n[33307];
assign t[33308] = t[33307] ^ n[33308];
assign t[33309] = t[33308] ^ n[33309];
assign t[33310] = t[33309] ^ n[33310];
assign t[33311] = t[33310] ^ n[33311];
assign t[33312] = t[33311] ^ n[33312];
assign t[33313] = t[33312] ^ n[33313];
assign t[33314] = t[33313] ^ n[33314];
assign t[33315] = t[33314] ^ n[33315];
assign t[33316] = t[33315] ^ n[33316];
assign t[33317] = t[33316] ^ n[33317];
assign t[33318] = t[33317] ^ n[33318];
assign t[33319] = t[33318] ^ n[33319];
assign t[33320] = t[33319] ^ n[33320];
assign t[33321] = t[33320] ^ n[33321];
assign t[33322] = t[33321] ^ n[33322];
assign t[33323] = t[33322] ^ n[33323];
assign t[33324] = t[33323] ^ n[33324];
assign t[33325] = t[33324] ^ n[33325];
assign t[33326] = t[33325] ^ n[33326];
assign t[33327] = t[33326] ^ n[33327];
assign t[33328] = t[33327] ^ n[33328];
assign t[33329] = t[33328] ^ n[33329];
assign t[33330] = t[33329] ^ n[33330];
assign t[33331] = t[33330] ^ n[33331];
assign t[33332] = t[33331] ^ n[33332];
assign t[33333] = t[33332] ^ n[33333];
assign t[33334] = t[33333] ^ n[33334];
assign t[33335] = t[33334] ^ n[33335];
assign t[33336] = t[33335] ^ n[33336];
assign t[33337] = t[33336] ^ n[33337];
assign t[33338] = t[33337] ^ n[33338];
assign t[33339] = t[33338] ^ n[33339];
assign t[33340] = t[33339] ^ n[33340];
assign t[33341] = t[33340] ^ n[33341];
assign t[33342] = t[33341] ^ n[33342];
assign t[33343] = t[33342] ^ n[33343];
assign t[33344] = t[33343] ^ n[33344];
assign t[33345] = t[33344] ^ n[33345];
assign t[33346] = t[33345] ^ n[33346];
assign t[33347] = t[33346] ^ n[33347];
assign t[33348] = t[33347] ^ n[33348];
assign t[33349] = t[33348] ^ n[33349];
assign t[33350] = t[33349] ^ n[33350];
assign t[33351] = t[33350] ^ n[33351];
assign t[33352] = t[33351] ^ n[33352];
assign t[33353] = t[33352] ^ n[33353];
assign t[33354] = t[33353] ^ n[33354];
assign t[33355] = t[33354] ^ n[33355];
assign t[33356] = t[33355] ^ n[33356];
assign t[33357] = t[33356] ^ n[33357];
assign t[33358] = t[33357] ^ n[33358];
assign t[33359] = t[33358] ^ n[33359];
assign t[33360] = t[33359] ^ n[33360];
assign t[33361] = t[33360] ^ n[33361];
assign t[33362] = t[33361] ^ n[33362];
assign t[33363] = t[33362] ^ n[33363];
assign t[33364] = t[33363] ^ n[33364];
assign t[33365] = t[33364] ^ n[33365];
assign t[33366] = t[33365] ^ n[33366];
assign t[33367] = t[33366] ^ n[33367];
assign t[33368] = t[33367] ^ n[33368];
assign t[33369] = t[33368] ^ n[33369];
assign t[33370] = t[33369] ^ n[33370];
assign t[33371] = t[33370] ^ n[33371];
assign t[33372] = t[33371] ^ n[33372];
assign t[33373] = t[33372] ^ n[33373];
assign t[33374] = t[33373] ^ n[33374];
assign t[33375] = t[33374] ^ n[33375];
assign t[33376] = t[33375] ^ n[33376];
assign t[33377] = t[33376] ^ n[33377];
assign t[33378] = t[33377] ^ n[33378];
assign t[33379] = t[33378] ^ n[33379];
assign t[33380] = t[33379] ^ n[33380];
assign t[33381] = t[33380] ^ n[33381];
assign t[33382] = t[33381] ^ n[33382];
assign t[33383] = t[33382] ^ n[33383];
assign t[33384] = t[33383] ^ n[33384];
assign t[33385] = t[33384] ^ n[33385];
assign t[33386] = t[33385] ^ n[33386];
assign t[33387] = t[33386] ^ n[33387];
assign t[33388] = t[33387] ^ n[33388];
assign t[33389] = t[33388] ^ n[33389];
assign t[33390] = t[33389] ^ n[33390];
assign t[33391] = t[33390] ^ n[33391];
assign t[33392] = t[33391] ^ n[33392];
assign t[33393] = t[33392] ^ n[33393];
assign t[33394] = t[33393] ^ n[33394];
assign t[33395] = t[33394] ^ n[33395];
assign t[33396] = t[33395] ^ n[33396];
assign t[33397] = t[33396] ^ n[33397];
assign t[33398] = t[33397] ^ n[33398];
assign t[33399] = t[33398] ^ n[33399];
assign t[33400] = t[33399] ^ n[33400];
assign t[33401] = t[33400] ^ n[33401];
assign t[33402] = t[33401] ^ n[33402];
assign t[33403] = t[33402] ^ n[33403];
assign t[33404] = t[33403] ^ n[33404];
assign t[33405] = t[33404] ^ n[33405];
assign t[33406] = t[33405] ^ n[33406];
assign t[33407] = t[33406] ^ n[33407];
assign t[33408] = t[33407] ^ n[33408];
assign t[33409] = t[33408] ^ n[33409];
assign t[33410] = t[33409] ^ n[33410];
assign t[33411] = t[33410] ^ n[33411];
assign t[33412] = t[33411] ^ n[33412];
assign t[33413] = t[33412] ^ n[33413];
assign t[33414] = t[33413] ^ n[33414];
assign t[33415] = t[33414] ^ n[33415];
assign t[33416] = t[33415] ^ n[33416];
assign t[33417] = t[33416] ^ n[33417];
assign t[33418] = t[33417] ^ n[33418];
assign t[33419] = t[33418] ^ n[33419];
assign t[33420] = t[33419] ^ n[33420];
assign t[33421] = t[33420] ^ n[33421];
assign t[33422] = t[33421] ^ n[33422];
assign t[33423] = t[33422] ^ n[33423];
assign t[33424] = t[33423] ^ n[33424];
assign t[33425] = t[33424] ^ n[33425];
assign t[33426] = t[33425] ^ n[33426];
assign t[33427] = t[33426] ^ n[33427];
assign t[33428] = t[33427] ^ n[33428];
assign t[33429] = t[33428] ^ n[33429];
assign t[33430] = t[33429] ^ n[33430];
assign t[33431] = t[33430] ^ n[33431];
assign t[33432] = t[33431] ^ n[33432];
assign t[33433] = t[33432] ^ n[33433];
assign t[33434] = t[33433] ^ n[33434];
assign t[33435] = t[33434] ^ n[33435];
assign t[33436] = t[33435] ^ n[33436];
assign t[33437] = t[33436] ^ n[33437];
assign t[33438] = t[33437] ^ n[33438];
assign t[33439] = t[33438] ^ n[33439];
assign t[33440] = t[33439] ^ n[33440];
assign t[33441] = t[33440] ^ n[33441];
assign t[33442] = t[33441] ^ n[33442];
assign t[33443] = t[33442] ^ n[33443];
assign t[33444] = t[33443] ^ n[33444];
assign t[33445] = t[33444] ^ n[33445];
assign t[33446] = t[33445] ^ n[33446];
assign t[33447] = t[33446] ^ n[33447];
assign t[33448] = t[33447] ^ n[33448];
assign t[33449] = t[33448] ^ n[33449];
assign t[33450] = t[33449] ^ n[33450];
assign t[33451] = t[33450] ^ n[33451];
assign t[33452] = t[33451] ^ n[33452];
assign t[33453] = t[33452] ^ n[33453];
assign t[33454] = t[33453] ^ n[33454];
assign t[33455] = t[33454] ^ n[33455];
assign t[33456] = t[33455] ^ n[33456];
assign t[33457] = t[33456] ^ n[33457];
assign t[33458] = t[33457] ^ n[33458];
assign t[33459] = t[33458] ^ n[33459];
assign t[33460] = t[33459] ^ n[33460];
assign t[33461] = t[33460] ^ n[33461];
assign t[33462] = t[33461] ^ n[33462];
assign t[33463] = t[33462] ^ n[33463];
assign t[33464] = t[33463] ^ n[33464];
assign t[33465] = t[33464] ^ n[33465];
assign t[33466] = t[33465] ^ n[33466];
assign t[33467] = t[33466] ^ n[33467];
assign t[33468] = t[33467] ^ n[33468];
assign t[33469] = t[33468] ^ n[33469];
assign t[33470] = t[33469] ^ n[33470];
assign t[33471] = t[33470] ^ n[33471];
assign t[33472] = t[33471] ^ n[33472];
assign t[33473] = t[33472] ^ n[33473];
assign t[33474] = t[33473] ^ n[33474];
assign t[33475] = t[33474] ^ n[33475];
assign t[33476] = t[33475] ^ n[33476];
assign t[33477] = t[33476] ^ n[33477];
assign t[33478] = t[33477] ^ n[33478];
assign t[33479] = t[33478] ^ n[33479];
assign t[33480] = t[33479] ^ n[33480];
assign t[33481] = t[33480] ^ n[33481];
assign t[33482] = t[33481] ^ n[33482];
assign t[33483] = t[33482] ^ n[33483];
assign t[33484] = t[33483] ^ n[33484];
assign t[33485] = t[33484] ^ n[33485];
assign t[33486] = t[33485] ^ n[33486];
assign t[33487] = t[33486] ^ n[33487];
assign t[33488] = t[33487] ^ n[33488];
assign t[33489] = t[33488] ^ n[33489];
assign t[33490] = t[33489] ^ n[33490];
assign t[33491] = t[33490] ^ n[33491];
assign t[33492] = t[33491] ^ n[33492];
assign t[33493] = t[33492] ^ n[33493];
assign t[33494] = t[33493] ^ n[33494];
assign t[33495] = t[33494] ^ n[33495];
assign t[33496] = t[33495] ^ n[33496];
assign t[33497] = t[33496] ^ n[33497];
assign t[33498] = t[33497] ^ n[33498];
assign t[33499] = t[33498] ^ n[33499];
assign t[33500] = t[33499] ^ n[33500];
assign t[33501] = t[33500] ^ n[33501];
assign t[33502] = t[33501] ^ n[33502];
assign t[33503] = t[33502] ^ n[33503];
assign t[33504] = t[33503] ^ n[33504];
assign t[33505] = t[33504] ^ n[33505];
assign t[33506] = t[33505] ^ n[33506];
assign t[33507] = t[33506] ^ n[33507];
assign t[33508] = t[33507] ^ n[33508];
assign t[33509] = t[33508] ^ n[33509];
assign t[33510] = t[33509] ^ n[33510];
assign t[33511] = t[33510] ^ n[33511];
assign t[33512] = t[33511] ^ n[33512];
assign t[33513] = t[33512] ^ n[33513];
assign t[33514] = t[33513] ^ n[33514];
assign t[33515] = t[33514] ^ n[33515];
assign t[33516] = t[33515] ^ n[33516];
assign t[33517] = t[33516] ^ n[33517];
assign t[33518] = t[33517] ^ n[33518];
assign t[33519] = t[33518] ^ n[33519];
assign t[33520] = t[33519] ^ n[33520];
assign t[33521] = t[33520] ^ n[33521];
assign t[33522] = t[33521] ^ n[33522];
assign t[33523] = t[33522] ^ n[33523];
assign t[33524] = t[33523] ^ n[33524];
assign t[33525] = t[33524] ^ n[33525];
assign t[33526] = t[33525] ^ n[33526];
assign t[33527] = t[33526] ^ n[33527];
assign t[33528] = t[33527] ^ n[33528];
assign t[33529] = t[33528] ^ n[33529];
assign t[33530] = t[33529] ^ n[33530];
assign t[33531] = t[33530] ^ n[33531];
assign t[33532] = t[33531] ^ n[33532];
assign t[33533] = t[33532] ^ n[33533];
assign t[33534] = t[33533] ^ n[33534];
assign t[33535] = t[33534] ^ n[33535];
assign t[33536] = t[33535] ^ n[33536];
assign t[33537] = t[33536] ^ n[33537];
assign t[33538] = t[33537] ^ n[33538];
assign t[33539] = t[33538] ^ n[33539];
assign t[33540] = t[33539] ^ n[33540];
assign t[33541] = t[33540] ^ n[33541];
assign t[33542] = t[33541] ^ n[33542];
assign t[33543] = t[33542] ^ n[33543];
assign t[33544] = t[33543] ^ n[33544];
assign t[33545] = t[33544] ^ n[33545];
assign t[33546] = t[33545] ^ n[33546];
assign t[33547] = t[33546] ^ n[33547];
assign t[33548] = t[33547] ^ n[33548];
assign t[33549] = t[33548] ^ n[33549];
assign t[33550] = t[33549] ^ n[33550];
assign t[33551] = t[33550] ^ n[33551];
assign t[33552] = t[33551] ^ n[33552];
assign t[33553] = t[33552] ^ n[33553];
assign t[33554] = t[33553] ^ n[33554];
assign t[33555] = t[33554] ^ n[33555];
assign t[33556] = t[33555] ^ n[33556];
assign t[33557] = t[33556] ^ n[33557];
assign t[33558] = t[33557] ^ n[33558];
assign t[33559] = t[33558] ^ n[33559];
assign t[33560] = t[33559] ^ n[33560];
assign t[33561] = t[33560] ^ n[33561];
assign t[33562] = t[33561] ^ n[33562];
assign t[33563] = t[33562] ^ n[33563];
assign t[33564] = t[33563] ^ n[33564];
assign t[33565] = t[33564] ^ n[33565];
assign t[33566] = t[33565] ^ n[33566];
assign t[33567] = t[33566] ^ n[33567];
assign t[33568] = t[33567] ^ n[33568];
assign t[33569] = t[33568] ^ n[33569];
assign t[33570] = t[33569] ^ n[33570];
assign t[33571] = t[33570] ^ n[33571];
assign t[33572] = t[33571] ^ n[33572];
assign t[33573] = t[33572] ^ n[33573];
assign t[33574] = t[33573] ^ n[33574];
assign t[33575] = t[33574] ^ n[33575];
assign t[33576] = t[33575] ^ n[33576];
assign t[33577] = t[33576] ^ n[33577];
assign t[33578] = t[33577] ^ n[33578];
assign t[33579] = t[33578] ^ n[33579];
assign t[33580] = t[33579] ^ n[33580];
assign t[33581] = t[33580] ^ n[33581];
assign t[33582] = t[33581] ^ n[33582];
assign t[33583] = t[33582] ^ n[33583];
assign t[33584] = t[33583] ^ n[33584];
assign t[33585] = t[33584] ^ n[33585];
assign t[33586] = t[33585] ^ n[33586];
assign t[33587] = t[33586] ^ n[33587];
assign t[33588] = t[33587] ^ n[33588];
assign t[33589] = t[33588] ^ n[33589];
assign t[33590] = t[33589] ^ n[33590];
assign t[33591] = t[33590] ^ n[33591];
assign t[33592] = t[33591] ^ n[33592];
assign t[33593] = t[33592] ^ n[33593];
assign t[33594] = t[33593] ^ n[33594];
assign t[33595] = t[33594] ^ n[33595];
assign t[33596] = t[33595] ^ n[33596];
assign t[33597] = t[33596] ^ n[33597];
assign t[33598] = t[33597] ^ n[33598];
assign t[33599] = t[33598] ^ n[33599];
assign t[33600] = t[33599] ^ n[33600];
assign t[33601] = t[33600] ^ n[33601];
assign t[33602] = t[33601] ^ n[33602];
assign t[33603] = t[33602] ^ n[33603];
assign t[33604] = t[33603] ^ n[33604];
assign t[33605] = t[33604] ^ n[33605];
assign t[33606] = t[33605] ^ n[33606];
assign t[33607] = t[33606] ^ n[33607];
assign t[33608] = t[33607] ^ n[33608];
assign t[33609] = t[33608] ^ n[33609];
assign t[33610] = t[33609] ^ n[33610];
assign t[33611] = t[33610] ^ n[33611];
assign t[33612] = t[33611] ^ n[33612];
assign t[33613] = t[33612] ^ n[33613];
assign t[33614] = t[33613] ^ n[33614];
assign t[33615] = t[33614] ^ n[33615];
assign t[33616] = t[33615] ^ n[33616];
assign t[33617] = t[33616] ^ n[33617];
assign t[33618] = t[33617] ^ n[33618];
assign t[33619] = t[33618] ^ n[33619];
assign t[33620] = t[33619] ^ n[33620];
assign t[33621] = t[33620] ^ n[33621];
assign t[33622] = t[33621] ^ n[33622];
assign t[33623] = t[33622] ^ n[33623];
assign t[33624] = t[33623] ^ n[33624];
assign t[33625] = t[33624] ^ n[33625];
assign t[33626] = t[33625] ^ n[33626];
assign t[33627] = t[33626] ^ n[33627];
assign t[33628] = t[33627] ^ n[33628];
assign t[33629] = t[33628] ^ n[33629];
assign t[33630] = t[33629] ^ n[33630];
assign t[33631] = t[33630] ^ n[33631];
assign t[33632] = t[33631] ^ n[33632];
assign t[33633] = t[33632] ^ n[33633];
assign t[33634] = t[33633] ^ n[33634];
assign t[33635] = t[33634] ^ n[33635];
assign t[33636] = t[33635] ^ n[33636];
assign t[33637] = t[33636] ^ n[33637];
assign t[33638] = t[33637] ^ n[33638];
assign t[33639] = t[33638] ^ n[33639];
assign t[33640] = t[33639] ^ n[33640];
assign t[33641] = t[33640] ^ n[33641];
assign t[33642] = t[33641] ^ n[33642];
assign t[33643] = t[33642] ^ n[33643];
assign t[33644] = t[33643] ^ n[33644];
assign t[33645] = t[33644] ^ n[33645];
assign t[33646] = t[33645] ^ n[33646];
assign t[33647] = t[33646] ^ n[33647];
assign t[33648] = t[33647] ^ n[33648];
assign t[33649] = t[33648] ^ n[33649];
assign t[33650] = t[33649] ^ n[33650];
assign t[33651] = t[33650] ^ n[33651];
assign t[33652] = t[33651] ^ n[33652];
assign t[33653] = t[33652] ^ n[33653];
assign t[33654] = t[33653] ^ n[33654];
assign t[33655] = t[33654] ^ n[33655];
assign t[33656] = t[33655] ^ n[33656];
assign t[33657] = t[33656] ^ n[33657];
assign t[33658] = t[33657] ^ n[33658];
assign t[33659] = t[33658] ^ n[33659];
assign t[33660] = t[33659] ^ n[33660];
assign t[33661] = t[33660] ^ n[33661];
assign t[33662] = t[33661] ^ n[33662];
assign t[33663] = t[33662] ^ n[33663];
assign t[33664] = t[33663] ^ n[33664];
assign t[33665] = t[33664] ^ n[33665];
assign t[33666] = t[33665] ^ n[33666];
assign t[33667] = t[33666] ^ n[33667];
assign t[33668] = t[33667] ^ n[33668];
assign t[33669] = t[33668] ^ n[33669];
assign t[33670] = t[33669] ^ n[33670];
assign t[33671] = t[33670] ^ n[33671];
assign t[33672] = t[33671] ^ n[33672];
assign t[33673] = t[33672] ^ n[33673];
assign t[33674] = t[33673] ^ n[33674];
assign t[33675] = t[33674] ^ n[33675];
assign t[33676] = t[33675] ^ n[33676];
assign t[33677] = t[33676] ^ n[33677];
assign t[33678] = t[33677] ^ n[33678];
assign t[33679] = t[33678] ^ n[33679];
assign t[33680] = t[33679] ^ n[33680];
assign t[33681] = t[33680] ^ n[33681];
assign t[33682] = t[33681] ^ n[33682];
assign t[33683] = t[33682] ^ n[33683];
assign t[33684] = t[33683] ^ n[33684];
assign t[33685] = t[33684] ^ n[33685];
assign t[33686] = t[33685] ^ n[33686];
assign t[33687] = t[33686] ^ n[33687];
assign t[33688] = t[33687] ^ n[33688];
assign t[33689] = t[33688] ^ n[33689];
assign t[33690] = t[33689] ^ n[33690];
assign t[33691] = t[33690] ^ n[33691];
assign t[33692] = t[33691] ^ n[33692];
assign t[33693] = t[33692] ^ n[33693];
assign t[33694] = t[33693] ^ n[33694];
assign t[33695] = t[33694] ^ n[33695];
assign t[33696] = t[33695] ^ n[33696];
assign t[33697] = t[33696] ^ n[33697];
assign t[33698] = t[33697] ^ n[33698];
assign t[33699] = t[33698] ^ n[33699];
assign t[33700] = t[33699] ^ n[33700];
assign t[33701] = t[33700] ^ n[33701];
assign t[33702] = t[33701] ^ n[33702];
assign t[33703] = t[33702] ^ n[33703];
assign t[33704] = t[33703] ^ n[33704];
assign t[33705] = t[33704] ^ n[33705];
assign t[33706] = t[33705] ^ n[33706];
assign t[33707] = t[33706] ^ n[33707];
assign t[33708] = t[33707] ^ n[33708];
assign t[33709] = t[33708] ^ n[33709];
assign t[33710] = t[33709] ^ n[33710];
assign t[33711] = t[33710] ^ n[33711];
assign t[33712] = t[33711] ^ n[33712];
assign t[33713] = t[33712] ^ n[33713];
assign t[33714] = t[33713] ^ n[33714];
assign t[33715] = t[33714] ^ n[33715];
assign t[33716] = t[33715] ^ n[33716];
assign t[33717] = t[33716] ^ n[33717];
assign t[33718] = t[33717] ^ n[33718];
assign t[33719] = t[33718] ^ n[33719];
assign t[33720] = t[33719] ^ n[33720];
assign t[33721] = t[33720] ^ n[33721];
assign t[33722] = t[33721] ^ n[33722];
assign t[33723] = t[33722] ^ n[33723];
assign t[33724] = t[33723] ^ n[33724];
assign t[33725] = t[33724] ^ n[33725];
assign t[33726] = t[33725] ^ n[33726];
assign t[33727] = t[33726] ^ n[33727];
assign t[33728] = t[33727] ^ n[33728];
assign t[33729] = t[33728] ^ n[33729];
assign t[33730] = t[33729] ^ n[33730];
assign t[33731] = t[33730] ^ n[33731];
assign t[33732] = t[33731] ^ n[33732];
assign t[33733] = t[33732] ^ n[33733];
assign t[33734] = t[33733] ^ n[33734];
assign t[33735] = t[33734] ^ n[33735];
assign t[33736] = t[33735] ^ n[33736];
assign t[33737] = t[33736] ^ n[33737];
assign t[33738] = t[33737] ^ n[33738];
assign t[33739] = t[33738] ^ n[33739];
assign t[33740] = t[33739] ^ n[33740];
assign t[33741] = t[33740] ^ n[33741];
assign t[33742] = t[33741] ^ n[33742];
assign t[33743] = t[33742] ^ n[33743];
assign t[33744] = t[33743] ^ n[33744];
assign t[33745] = t[33744] ^ n[33745];
assign t[33746] = t[33745] ^ n[33746];
assign t[33747] = t[33746] ^ n[33747];
assign t[33748] = t[33747] ^ n[33748];
assign t[33749] = t[33748] ^ n[33749];
assign t[33750] = t[33749] ^ n[33750];
assign t[33751] = t[33750] ^ n[33751];
assign t[33752] = t[33751] ^ n[33752];
assign t[33753] = t[33752] ^ n[33753];
assign t[33754] = t[33753] ^ n[33754];
assign t[33755] = t[33754] ^ n[33755];
assign t[33756] = t[33755] ^ n[33756];
assign t[33757] = t[33756] ^ n[33757];
assign t[33758] = t[33757] ^ n[33758];
assign t[33759] = t[33758] ^ n[33759];
assign t[33760] = t[33759] ^ n[33760];
assign t[33761] = t[33760] ^ n[33761];
assign t[33762] = t[33761] ^ n[33762];
assign t[33763] = t[33762] ^ n[33763];
assign t[33764] = t[33763] ^ n[33764];
assign t[33765] = t[33764] ^ n[33765];
assign t[33766] = t[33765] ^ n[33766];
assign t[33767] = t[33766] ^ n[33767];
assign t[33768] = t[33767] ^ n[33768];
assign t[33769] = t[33768] ^ n[33769];
assign t[33770] = t[33769] ^ n[33770];
assign t[33771] = t[33770] ^ n[33771];
assign t[33772] = t[33771] ^ n[33772];
assign t[33773] = t[33772] ^ n[33773];
assign t[33774] = t[33773] ^ n[33774];
assign t[33775] = t[33774] ^ n[33775];
assign t[33776] = t[33775] ^ n[33776];
assign t[33777] = t[33776] ^ n[33777];
assign t[33778] = t[33777] ^ n[33778];
assign t[33779] = t[33778] ^ n[33779];
assign t[33780] = t[33779] ^ n[33780];
assign t[33781] = t[33780] ^ n[33781];
assign t[33782] = t[33781] ^ n[33782];
assign t[33783] = t[33782] ^ n[33783];
assign t[33784] = t[33783] ^ n[33784];
assign t[33785] = t[33784] ^ n[33785];
assign t[33786] = t[33785] ^ n[33786];
assign t[33787] = t[33786] ^ n[33787];
assign t[33788] = t[33787] ^ n[33788];
assign t[33789] = t[33788] ^ n[33789];
assign t[33790] = t[33789] ^ n[33790];
assign t[33791] = t[33790] ^ n[33791];
assign t[33792] = t[33791] ^ n[33792];
assign t[33793] = t[33792] ^ n[33793];
assign t[33794] = t[33793] ^ n[33794];
assign t[33795] = t[33794] ^ n[33795];
assign t[33796] = t[33795] ^ n[33796];
assign t[33797] = t[33796] ^ n[33797];
assign t[33798] = t[33797] ^ n[33798];
assign t[33799] = t[33798] ^ n[33799];
assign t[33800] = t[33799] ^ n[33800];
assign t[33801] = t[33800] ^ n[33801];
assign t[33802] = t[33801] ^ n[33802];
assign t[33803] = t[33802] ^ n[33803];
assign t[33804] = t[33803] ^ n[33804];
assign t[33805] = t[33804] ^ n[33805];
assign t[33806] = t[33805] ^ n[33806];
assign t[33807] = t[33806] ^ n[33807];
assign t[33808] = t[33807] ^ n[33808];
assign t[33809] = t[33808] ^ n[33809];
assign t[33810] = t[33809] ^ n[33810];
assign t[33811] = t[33810] ^ n[33811];
assign t[33812] = t[33811] ^ n[33812];
assign t[33813] = t[33812] ^ n[33813];
assign t[33814] = t[33813] ^ n[33814];
assign t[33815] = t[33814] ^ n[33815];
assign t[33816] = t[33815] ^ n[33816];
assign t[33817] = t[33816] ^ n[33817];
assign t[33818] = t[33817] ^ n[33818];
assign t[33819] = t[33818] ^ n[33819];
assign t[33820] = t[33819] ^ n[33820];
assign t[33821] = t[33820] ^ n[33821];
assign t[33822] = t[33821] ^ n[33822];
assign t[33823] = t[33822] ^ n[33823];
assign t[33824] = t[33823] ^ n[33824];
assign t[33825] = t[33824] ^ n[33825];
assign t[33826] = t[33825] ^ n[33826];
assign t[33827] = t[33826] ^ n[33827];
assign t[33828] = t[33827] ^ n[33828];
assign t[33829] = t[33828] ^ n[33829];
assign t[33830] = t[33829] ^ n[33830];
assign t[33831] = t[33830] ^ n[33831];
assign t[33832] = t[33831] ^ n[33832];
assign t[33833] = t[33832] ^ n[33833];
assign t[33834] = t[33833] ^ n[33834];
assign t[33835] = t[33834] ^ n[33835];
assign t[33836] = t[33835] ^ n[33836];
assign t[33837] = t[33836] ^ n[33837];
assign t[33838] = t[33837] ^ n[33838];
assign t[33839] = t[33838] ^ n[33839];
assign t[33840] = t[33839] ^ n[33840];
assign t[33841] = t[33840] ^ n[33841];
assign t[33842] = t[33841] ^ n[33842];
assign t[33843] = t[33842] ^ n[33843];
assign t[33844] = t[33843] ^ n[33844];
assign t[33845] = t[33844] ^ n[33845];
assign t[33846] = t[33845] ^ n[33846];
assign t[33847] = t[33846] ^ n[33847];
assign t[33848] = t[33847] ^ n[33848];
assign t[33849] = t[33848] ^ n[33849];
assign t[33850] = t[33849] ^ n[33850];
assign t[33851] = t[33850] ^ n[33851];
assign t[33852] = t[33851] ^ n[33852];
assign t[33853] = t[33852] ^ n[33853];
assign t[33854] = t[33853] ^ n[33854];
assign t[33855] = t[33854] ^ n[33855];
assign t[33856] = t[33855] ^ n[33856];
assign t[33857] = t[33856] ^ n[33857];
assign t[33858] = t[33857] ^ n[33858];
assign t[33859] = t[33858] ^ n[33859];
assign t[33860] = t[33859] ^ n[33860];
assign t[33861] = t[33860] ^ n[33861];
assign t[33862] = t[33861] ^ n[33862];
assign t[33863] = t[33862] ^ n[33863];
assign t[33864] = t[33863] ^ n[33864];
assign t[33865] = t[33864] ^ n[33865];
assign t[33866] = t[33865] ^ n[33866];
assign t[33867] = t[33866] ^ n[33867];
assign t[33868] = t[33867] ^ n[33868];
assign t[33869] = t[33868] ^ n[33869];
assign t[33870] = t[33869] ^ n[33870];
assign t[33871] = t[33870] ^ n[33871];
assign t[33872] = t[33871] ^ n[33872];
assign t[33873] = t[33872] ^ n[33873];
assign t[33874] = t[33873] ^ n[33874];
assign t[33875] = t[33874] ^ n[33875];
assign t[33876] = t[33875] ^ n[33876];
assign t[33877] = t[33876] ^ n[33877];
assign t[33878] = t[33877] ^ n[33878];
assign t[33879] = t[33878] ^ n[33879];
assign t[33880] = t[33879] ^ n[33880];
assign t[33881] = t[33880] ^ n[33881];
assign t[33882] = t[33881] ^ n[33882];
assign t[33883] = t[33882] ^ n[33883];
assign t[33884] = t[33883] ^ n[33884];
assign t[33885] = t[33884] ^ n[33885];
assign t[33886] = t[33885] ^ n[33886];
assign t[33887] = t[33886] ^ n[33887];
assign t[33888] = t[33887] ^ n[33888];
assign t[33889] = t[33888] ^ n[33889];
assign t[33890] = t[33889] ^ n[33890];
assign t[33891] = t[33890] ^ n[33891];
assign t[33892] = t[33891] ^ n[33892];
assign t[33893] = t[33892] ^ n[33893];
assign t[33894] = t[33893] ^ n[33894];
assign t[33895] = t[33894] ^ n[33895];
assign t[33896] = t[33895] ^ n[33896];
assign t[33897] = t[33896] ^ n[33897];
assign t[33898] = t[33897] ^ n[33898];
assign t[33899] = t[33898] ^ n[33899];
assign t[33900] = t[33899] ^ n[33900];
assign t[33901] = t[33900] ^ n[33901];
assign t[33902] = t[33901] ^ n[33902];
assign t[33903] = t[33902] ^ n[33903];
assign t[33904] = t[33903] ^ n[33904];
assign t[33905] = t[33904] ^ n[33905];
assign t[33906] = t[33905] ^ n[33906];
assign t[33907] = t[33906] ^ n[33907];
assign t[33908] = t[33907] ^ n[33908];
assign t[33909] = t[33908] ^ n[33909];
assign t[33910] = t[33909] ^ n[33910];
assign t[33911] = t[33910] ^ n[33911];
assign t[33912] = t[33911] ^ n[33912];
assign t[33913] = t[33912] ^ n[33913];
assign t[33914] = t[33913] ^ n[33914];
assign t[33915] = t[33914] ^ n[33915];
assign t[33916] = t[33915] ^ n[33916];
assign t[33917] = t[33916] ^ n[33917];
assign t[33918] = t[33917] ^ n[33918];
assign t[33919] = t[33918] ^ n[33919];
assign t[33920] = t[33919] ^ n[33920];
assign t[33921] = t[33920] ^ n[33921];
assign t[33922] = t[33921] ^ n[33922];
assign t[33923] = t[33922] ^ n[33923];
assign t[33924] = t[33923] ^ n[33924];
assign t[33925] = t[33924] ^ n[33925];
assign t[33926] = t[33925] ^ n[33926];
assign t[33927] = t[33926] ^ n[33927];
assign t[33928] = t[33927] ^ n[33928];
assign t[33929] = t[33928] ^ n[33929];
assign t[33930] = t[33929] ^ n[33930];
assign t[33931] = t[33930] ^ n[33931];
assign t[33932] = t[33931] ^ n[33932];
assign t[33933] = t[33932] ^ n[33933];
assign t[33934] = t[33933] ^ n[33934];
assign t[33935] = t[33934] ^ n[33935];
assign t[33936] = t[33935] ^ n[33936];
assign t[33937] = t[33936] ^ n[33937];
assign t[33938] = t[33937] ^ n[33938];
assign t[33939] = t[33938] ^ n[33939];
assign t[33940] = t[33939] ^ n[33940];
assign t[33941] = t[33940] ^ n[33941];
assign t[33942] = t[33941] ^ n[33942];
assign t[33943] = t[33942] ^ n[33943];
assign t[33944] = t[33943] ^ n[33944];
assign t[33945] = t[33944] ^ n[33945];
assign t[33946] = t[33945] ^ n[33946];
assign t[33947] = t[33946] ^ n[33947];
assign t[33948] = t[33947] ^ n[33948];
assign t[33949] = t[33948] ^ n[33949];
assign t[33950] = t[33949] ^ n[33950];
assign t[33951] = t[33950] ^ n[33951];
assign t[33952] = t[33951] ^ n[33952];
assign t[33953] = t[33952] ^ n[33953];
assign t[33954] = t[33953] ^ n[33954];
assign t[33955] = t[33954] ^ n[33955];
assign t[33956] = t[33955] ^ n[33956];
assign t[33957] = t[33956] ^ n[33957];
assign t[33958] = t[33957] ^ n[33958];
assign t[33959] = t[33958] ^ n[33959];
assign t[33960] = t[33959] ^ n[33960];
assign t[33961] = t[33960] ^ n[33961];
assign t[33962] = t[33961] ^ n[33962];
assign t[33963] = t[33962] ^ n[33963];
assign t[33964] = t[33963] ^ n[33964];
assign t[33965] = t[33964] ^ n[33965];
assign t[33966] = t[33965] ^ n[33966];
assign t[33967] = t[33966] ^ n[33967];
assign t[33968] = t[33967] ^ n[33968];
assign t[33969] = t[33968] ^ n[33969];
assign t[33970] = t[33969] ^ n[33970];
assign t[33971] = t[33970] ^ n[33971];
assign t[33972] = t[33971] ^ n[33972];
assign t[33973] = t[33972] ^ n[33973];
assign t[33974] = t[33973] ^ n[33974];
assign t[33975] = t[33974] ^ n[33975];
assign t[33976] = t[33975] ^ n[33976];
assign t[33977] = t[33976] ^ n[33977];
assign t[33978] = t[33977] ^ n[33978];
assign t[33979] = t[33978] ^ n[33979];
assign t[33980] = t[33979] ^ n[33980];
assign t[33981] = t[33980] ^ n[33981];
assign t[33982] = t[33981] ^ n[33982];
assign t[33983] = t[33982] ^ n[33983];
assign t[33984] = t[33983] ^ n[33984];
assign t[33985] = t[33984] ^ n[33985];
assign t[33986] = t[33985] ^ n[33986];
assign t[33987] = t[33986] ^ n[33987];
assign t[33988] = t[33987] ^ n[33988];
assign t[33989] = t[33988] ^ n[33989];
assign t[33990] = t[33989] ^ n[33990];
assign t[33991] = t[33990] ^ n[33991];
assign t[33992] = t[33991] ^ n[33992];
assign t[33993] = t[33992] ^ n[33993];
assign t[33994] = t[33993] ^ n[33994];
assign t[33995] = t[33994] ^ n[33995];
assign t[33996] = t[33995] ^ n[33996];
assign t[33997] = t[33996] ^ n[33997];
assign t[33998] = t[33997] ^ n[33998];
assign t[33999] = t[33998] ^ n[33999];
assign t[34000] = t[33999] ^ n[34000];
assign t[34001] = t[34000] ^ n[34001];
assign t[34002] = t[34001] ^ n[34002];
assign t[34003] = t[34002] ^ n[34003];
assign t[34004] = t[34003] ^ n[34004];
assign t[34005] = t[34004] ^ n[34005];
assign t[34006] = t[34005] ^ n[34006];
assign t[34007] = t[34006] ^ n[34007];
assign t[34008] = t[34007] ^ n[34008];
assign t[34009] = t[34008] ^ n[34009];
assign t[34010] = t[34009] ^ n[34010];
assign t[34011] = t[34010] ^ n[34011];
assign t[34012] = t[34011] ^ n[34012];
assign t[34013] = t[34012] ^ n[34013];
assign t[34014] = t[34013] ^ n[34014];
assign t[34015] = t[34014] ^ n[34015];
assign t[34016] = t[34015] ^ n[34016];
assign t[34017] = t[34016] ^ n[34017];
assign t[34018] = t[34017] ^ n[34018];
assign t[34019] = t[34018] ^ n[34019];
assign t[34020] = t[34019] ^ n[34020];
assign t[34021] = t[34020] ^ n[34021];
assign t[34022] = t[34021] ^ n[34022];
assign t[34023] = t[34022] ^ n[34023];
assign t[34024] = t[34023] ^ n[34024];
assign t[34025] = t[34024] ^ n[34025];
assign t[34026] = t[34025] ^ n[34026];
assign t[34027] = t[34026] ^ n[34027];
assign t[34028] = t[34027] ^ n[34028];
assign t[34029] = t[34028] ^ n[34029];
assign t[34030] = t[34029] ^ n[34030];
assign t[34031] = t[34030] ^ n[34031];
assign t[34032] = t[34031] ^ n[34032];
assign t[34033] = t[34032] ^ n[34033];
assign t[34034] = t[34033] ^ n[34034];
assign t[34035] = t[34034] ^ n[34035];
assign t[34036] = t[34035] ^ n[34036];
assign t[34037] = t[34036] ^ n[34037];
assign t[34038] = t[34037] ^ n[34038];
assign t[34039] = t[34038] ^ n[34039];
assign t[34040] = t[34039] ^ n[34040];
assign t[34041] = t[34040] ^ n[34041];
assign t[34042] = t[34041] ^ n[34042];
assign t[34043] = t[34042] ^ n[34043];
assign t[34044] = t[34043] ^ n[34044];
assign t[34045] = t[34044] ^ n[34045];
assign t[34046] = t[34045] ^ n[34046];
assign t[34047] = t[34046] ^ n[34047];
assign t[34048] = t[34047] ^ n[34048];
assign t[34049] = t[34048] ^ n[34049];
assign t[34050] = t[34049] ^ n[34050];
assign t[34051] = t[34050] ^ n[34051];
assign t[34052] = t[34051] ^ n[34052];
assign t[34053] = t[34052] ^ n[34053];
assign t[34054] = t[34053] ^ n[34054];
assign t[34055] = t[34054] ^ n[34055];
assign t[34056] = t[34055] ^ n[34056];
assign t[34057] = t[34056] ^ n[34057];
assign t[34058] = t[34057] ^ n[34058];
assign t[34059] = t[34058] ^ n[34059];
assign t[34060] = t[34059] ^ n[34060];
assign t[34061] = t[34060] ^ n[34061];
assign t[34062] = t[34061] ^ n[34062];
assign t[34063] = t[34062] ^ n[34063];
assign t[34064] = t[34063] ^ n[34064];
assign t[34065] = t[34064] ^ n[34065];
assign t[34066] = t[34065] ^ n[34066];
assign t[34067] = t[34066] ^ n[34067];
assign t[34068] = t[34067] ^ n[34068];
assign t[34069] = t[34068] ^ n[34069];
assign t[34070] = t[34069] ^ n[34070];
assign t[34071] = t[34070] ^ n[34071];
assign t[34072] = t[34071] ^ n[34072];
assign t[34073] = t[34072] ^ n[34073];
assign t[34074] = t[34073] ^ n[34074];
assign t[34075] = t[34074] ^ n[34075];
assign t[34076] = t[34075] ^ n[34076];
assign t[34077] = t[34076] ^ n[34077];
assign t[34078] = t[34077] ^ n[34078];
assign t[34079] = t[34078] ^ n[34079];
assign t[34080] = t[34079] ^ n[34080];
assign t[34081] = t[34080] ^ n[34081];
assign t[34082] = t[34081] ^ n[34082];
assign t[34083] = t[34082] ^ n[34083];
assign t[34084] = t[34083] ^ n[34084];
assign t[34085] = t[34084] ^ n[34085];
assign t[34086] = t[34085] ^ n[34086];
assign t[34087] = t[34086] ^ n[34087];
assign t[34088] = t[34087] ^ n[34088];
assign t[34089] = t[34088] ^ n[34089];
assign t[34090] = t[34089] ^ n[34090];
assign t[34091] = t[34090] ^ n[34091];
assign t[34092] = t[34091] ^ n[34092];
assign t[34093] = t[34092] ^ n[34093];
assign t[34094] = t[34093] ^ n[34094];
assign t[34095] = t[34094] ^ n[34095];
assign t[34096] = t[34095] ^ n[34096];
assign t[34097] = t[34096] ^ n[34097];
assign t[34098] = t[34097] ^ n[34098];
assign t[34099] = t[34098] ^ n[34099];
assign t[34100] = t[34099] ^ n[34100];
assign t[34101] = t[34100] ^ n[34101];
assign t[34102] = t[34101] ^ n[34102];
assign t[34103] = t[34102] ^ n[34103];
assign t[34104] = t[34103] ^ n[34104];
assign t[34105] = t[34104] ^ n[34105];
assign t[34106] = t[34105] ^ n[34106];
assign t[34107] = t[34106] ^ n[34107];
assign t[34108] = t[34107] ^ n[34108];
assign t[34109] = t[34108] ^ n[34109];
assign t[34110] = t[34109] ^ n[34110];
assign t[34111] = t[34110] ^ n[34111];
assign t[34112] = t[34111] ^ n[34112];
assign t[34113] = t[34112] ^ n[34113];
assign t[34114] = t[34113] ^ n[34114];
assign t[34115] = t[34114] ^ n[34115];
assign t[34116] = t[34115] ^ n[34116];
assign t[34117] = t[34116] ^ n[34117];
assign t[34118] = t[34117] ^ n[34118];
assign t[34119] = t[34118] ^ n[34119];
assign t[34120] = t[34119] ^ n[34120];
assign t[34121] = t[34120] ^ n[34121];
assign t[34122] = t[34121] ^ n[34122];
assign t[34123] = t[34122] ^ n[34123];
assign t[34124] = t[34123] ^ n[34124];
assign t[34125] = t[34124] ^ n[34125];
assign t[34126] = t[34125] ^ n[34126];
assign t[34127] = t[34126] ^ n[34127];
assign t[34128] = t[34127] ^ n[34128];
assign t[34129] = t[34128] ^ n[34129];
assign t[34130] = t[34129] ^ n[34130];
assign t[34131] = t[34130] ^ n[34131];
assign t[34132] = t[34131] ^ n[34132];
assign t[34133] = t[34132] ^ n[34133];
assign t[34134] = t[34133] ^ n[34134];
assign t[34135] = t[34134] ^ n[34135];
assign t[34136] = t[34135] ^ n[34136];
assign t[34137] = t[34136] ^ n[34137];
assign t[34138] = t[34137] ^ n[34138];
assign t[34139] = t[34138] ^ n[34139];
assign t[34140] = t[34139] ^ n[34140];
assign t[34141] = t[34140] ^ n[34141];
assign t[34142] = t[34141] ^ n[34142];
assign t[34143] = t[34142] ^ n[34143];
assign t[34144] = t[34143] ^ n[34144];
assign t[34145] = t[34144] ^ n[34145];
assign t[34146] = t[34145] ^ n[34146];
assign t[34147] = t[34146] ^ n[34147];
assign t[34148] = t[34147] ^ n[34148];
assign t[34149] = t[34148] ^ n[34149];
assign t[34150] = t[34149] ^ n[34150];
assign t[34151] = t[34150] ^ n[34151];
assign t[34152] = t[34151] ^ n[34152];
assign t[34153] = t[34152] ^ n[34153];
assign t[34154] = t[34153] ^ n[34154];
assign t[34155] = t[34154] ^ n[34155];
assign t[34156] = t[34155] ^ n[34156];
assign t[34157] = t[34156] ^ n[34157];
assign t[34158] = t[34157] ^ n[34158];
assign t[34159] = t[34158] ^ n[34159];
assign t[34160] = t[34159] ^ n[34160];
assign t[34161] = t[34160] ^ n[34161];
assign t[34162] = t[34161] ^ n[34162];
assign t[34163] = t[34162] ^ n[34163];
assign t[34164] = t[34163] ^ n[34164];
assign t[34165] = t[34164] ^ n[34165];
assign t[34166] = t[34165] ^ n[34166];
assign t[34167] = t[34166] ^ n[34167];
assign t[34168] = t[34167] ^ n[34168];
assign t[34169] = t[34168] ^ n[34169];
assign t[34170] = t[34169] ^ n[34170];
assign t[34171] = t[34170] ^ n[34171];
assign t[34172] = t[34171] ^ n[34172];
assign t[34173] = t[34172] ^ n[34173];
assign t[34174] = t[34173] ^ n[34174];
assign t[34175] = t[34174] ^ n[34175];
assign t[34176] = t[34175] ^ n[34176];
assign t[34177] = t[34176] ^ n[34177];
assign t[34178] = t[34177] ^ n[34178];
assign t[34179] = t[34178] ^ n[34179];
assign t[34180] = t[34179] ^ n[34180];
assign t[34181] = t[34180] ^ n[34181];
assign t[34182] = t[34181] ^ n[34182];
assign t[34183] = t[34182] ^ n[34183];
assign t[34184] = t[34183] ^ n[34184];
assign t[34185] = t[34184] ^ n[34185];
assign t[34186] = t[34185] ^ n[34186];
assign t[34187] = t[34186] ^ n[34187];
assign t[34188] = t[34187] ^ n[34188];
assign t[34189] = t[34188] ^ n[34189];
assign t[34190] = t[34189] ^ n[34190];
assign t[34191] = t[34190] ^ n[34191];
assign t[34192] = t[34191] ^ n[34192];
assign t[34193] = t[34192] ^ n[34193];
assign t[34194] = t[34193] ^ n[34194];
assign t[34195] = t[34194] ^ n[34195];
assign t[34196] = t[34195] ^ n[34196];
assign t[34197] = t[34196] ^ n[34197];
assign t[34198] = t[34197] ^ n[34198];
assign t[34199] = t[34198] ^ n[34199];
assign t[34200] = t[34199] ^ n[34200];
assign t[34201] = t[34200] ^ n[34201];
assign t[34202] = t[34201] ^ n[34202];
assign t[34203] = t[34202] ^ n[34203];
assign t[34204] = t[34203] ^ n[34204];
assign t[34205] = t[34204] ^ n[34205];
assign t[34206] = t[34205] ^ n[34206];
assign t[34207] = t[34206] ^ n[34207];
assign t[34208] = t[34207] ^ n[34208];
assign t[34209] = t[34208] ^ n[34209];
assign t[34210] = t[34209] ^ n[34210];
assign t[34211] = t[34210] ^ n[34211];
assign t[34212] = t[34211] ^ n[34212];
assign t[34213] = t[34212] ^ n[34213];
assign t[34214] = t[34213] ^ n[34214];
assign t[34215] = t[34214] ^ n[34215];
assign t[34216] = t[34215] ^ n[34216];
assign t[34217] = t[34216] ^ n[34217];
assign t[34218] = t[34217] ^ n[34218];
assign t[34219] = t[34218] ^ n[34219];
assign t[34220] = t[34219] ^ n[34220];
assign t[34221] = t[34220] ^ n[34221];
assign t[34222] = t[34221] ^ n[34222];
assign t[34223] = t[34222] ^ n[34223];
assign t[34224] = t[34223] ^ n[34224];
assign t[34225] = t[34224] ^ n[34225];
assign t[34226] = t[34225] ^ n[34226];
assign t[34227] = t[34226] ^ n[34227];
assign t[34228] = t[34227] ^ n[34228];
assign t[34229] = t[34228] ^ n[34229];
assign t[34230] = t[34229] ^ n[34230];
assign t[34231] = t[34230] ^ n[34231];
assign t[34232] = t[34231] ^ n[34232];
assign t[34233] = t[34232] ^ n[34233];
assign t[34234] = t[34233] ^ n[34234];
assign t[34235] = t[34234] ^ n[34235];
assign t[34236] = t[34235] ^ n[34236];
assign t[34237] = t[34236] ^ n[34237];
assign t[34238] = t[34237] ^ n[34238];
assign t[34239] = t[34238] ^ n[34239];
assign t[34240] = t[34239] ^ n[34240];
assign t[34241] = t[34240] ^ n[34241];
assign t[34242] = t[34241] ^ n[34242];
assign t[34243] = t[34242] ^ n[34243];
assign t[34244] = t[34243] ^ n[34244];
assign t[34245] = t[34244] ^ n[34245];
assign t[34246] = t[34245] ^ n[34246];
assign t[34247] = t[34246] ^ n[34247];
assign t[34248] = t[34247] ^ n[34248];
assign t[34249] = t[34248] ^ n[34249];
assign t[34250] = t[34249] ^ n[34250];
assign t[34251] = t[34250] ^ n[34251];
assign t[34252] = t[34251] ^ n[34252];
assign t[34253] = t[34252] ^ n[34253];
assign t[34254] = t[34253] ^ n[34254];
assign t[34255] = t[34254] ^ n[34255];
assign t[34256] = t[34255] ^ n[34256];
assign t[34257] = t[34256] ^ n[34257];
assign t[34258] = t[34257] ^ n[34258];
assign t[34259] = t[34258] ^ n[34259];
assign t[34260] = t[34259] ^ n[34260];
assign t[34261] = t[34260] ^ n[34261];
assign t[34262] = t[34261] ^ n[34262];
assign t[34263] = t[34262] ^ n[34263];
assign t[34264] = t[34263] ^ n[34264];
assign t[34265] = t[34264] ^ n[34265];
assign t[34266] = t[34265] ^ n[34266];
assign t[34267] = t[34266] ^ n[34267];
assign t[34268] = t[34267] ^ n[34268];
assign t[34269] = t[34268] ^ n[34269];
assign t[34270] = t[34269] ^ n[34270];
assign t[34271] = t[34270] ^ n[34271];
assign t[34272] = t[34271] ^ n[34272];
assign t[34273] = t[34272] ^ n[34273];
assign t[34274] = t[34273] ^ n[34274];
assign t[34275] = t[34274] ^ n[34275];
assign t[34276] = t[34275] ^ n[34276];
assign t[34277] = t[34276] ^ n[34277];
assign t[34278] = t[34277] ^ n[34278];
assign t[34279] = t[34278] ^ n[34279];
assign t[34280] = t[34279] ^ n[34280];
assign t[34281] = t[34280] ^ n[34281];
assign t[34282] = t[34281] ^ n[34282];
assign t[34283] = t[34282] ^ n[34283];
assign t[34284] = t[34283] ^ n[34284];
assign t[34285] = t[34284] ^ n[34285];
assign t[34286] = t[34285] ^ n[34286];
assign t[34287] = t[34286] ^ n[34287];
assign t[34288] = t[34287] ^ n[34288];
assign t[34289] = t[34288] ^ n[34289];
assign t[34290] = t[34289] ^ n[34290];
assign t[34291] = t[34290] ^ n[34291];
assign t[34292] = t[34291] ^ n[34292];
assign t[34293] = t[34292] ^ n[34293];
assign t[34294] = t[34293] ^ n[34294];
assign t[34295] = t[34294] ^ n[34295];
assign t[34296] = t[34295] ^ n[34296];
assign t[34297] = t[34296] ^ n[34297];
assign t[34298] = t[34297] ^ n[34298];
assign t[34299] = t[34298] ^ n[34299];
assign t[34300] = t[34299] ^ n[34300];
assign t[34301] = t[34300] ^ n[34301];
assign t[34302] = t[34301] ^ n[34302];
assign t[34303] = t[34302] ^ n[34303];
assign t[34304] = t[34303] ^ n[34304];
assign t[34305] = t[34304] ^ n[34305];
assign t[34306] = t[34305] ^ n[34306];
assign t[34307] = t[34306] ^ n[34307];
assign t[34308] = t[34307] ^ n[34308];
assign t[34309] = t[34308] ^ n[34309];
assign t[34310] = t[34309] ^ n[34310];
assign t[34311] = t[34310] ^ n[34311];
assign t[34312] = t[34311] ^ n[34312];
assign t[34313] = t[34312] ^ n[34313];
assign t[34314] = t[34313] ^ n[34314];
assign t[34315] = t[34314] ^ n[34315];
assign t[34316] = t[34315] ^ n[34316];
assign t[34317] = t[34316] ^ n[34317];
assign t[34318] = t[34317] ^ n[34318];
assign t[34319] = t[34318] ^ n[34319];
assign t[34320] = t[34319] ^ n[34320];
assign t[34321] = t[34320] ^ n[34321];
assign t[34322] = t[34321] ^ n[34322];
assign t[34323] = t[34322] ^ n[34323];
assign t[34324] = t[34323] ^ n[34324];
assign t[34325] = t[34324] ^ n[34325];
assign t[34326] = t[34325] ^ n[34326];
assign t[34327] = t[34326] ^ n[34327];
assign t[34328] = t[34327] ^ n[34328];
assign t[34329] = t[34328] ^ n[34329];
assign t[34330] = t[34329] ^ n[34330];
assign t[34331] = t[34330] ^ n[34331];
assign t[34332] = t[34331] ^ n[34332];
assign t[34333] = t[34332] ^ n[34333];
assign t[34334] = t[34333] ^ n[34334];
assign t[34335] = t[34334] ^ n[34335];
assign t[34336] = t[34335] ^ n[34336];
assign t[34337] = t[34336] ^ n[34337];
assign t[34338] = t[34337] ^ n[34338];
assign t[34339] = t[34338] ^ n[34339];
assign t[34340] = t[34339] ^ n[34340];
assign t[34341] = t[34340] ^ n[34341];
assign t[34342] = t[34341] ^ n[34342];
assign t[34343] = t[34342] ^ n[34343];
assign t[34344] = t[34343] ^ n[34344];
assign t[34345] = t[34344] ^ n[34345];
assign t[34346] = t[34345] ^ n[34346];
assign t[34347] = t[34346] ^ n[34347];
assign t[34348] = t[34347] ^ n[34348];
assign t[34349] = t[34348] ^ n[34349];
assign t[34350] = t[34349] ^ n[34350];
assign t[34351] = t[34350] ^ n[34351];
assign t[34352] = t[34351] ^ n[34352];
assign t[34353] = t[34352] ^ n[34353];
assign t[34354] = t[34353] ^ n[34354];
assign t[34355] = t[34354] ^ n[34355];
assign t[34356] = t[34355] ^ n[34356];
assign t[34357] = t[34356] ^ n[34357];
assign t[34358] = t[34357] ^ n[34358];
assign t[34359] = t[34358] ^ n[34359];
assign t[34360] = t[34359] ^ n[34360];
assign t[34361] = t[34360] ^ n[34361];
assign t[34362] = t[34361] ^ n[34362];
assign t[34363] = t[34362] ^ n[34363];
assign t[34364] = t[34363] ^ n[34364];
assign t[34365] = t[34364] ^ n[34365];
assign t[34366] = t[34365] ^ n[34366];
assign t[34367] = t[34366] ^ n[34367];
assign t[34368] = t[34367] ^ n[34368];
assign t[34369] = t[34368] ^ n[34369];
assign t[34370] = t[34369] ^ n[34370];
assign t[34371] = t[34370] ^ n[34371];
assign t[34372] = t[34371] ^ n[34372];
assign t[34373] = t[34372] ^ n[34373];
assign t[34374] = t[34373] ^ n[34374];
assign t[34375] = t[34374] ^ n[34375];
assign t[34376] = t[34375] ^ n[34376];
assign t[34377] = t[34376] ^ n[34377];
assign t[34378] = t[34377] ^ n[34378];
assign t[34379] = t[34378] ^ n[34379];
assign t[34380] = t[34379] ^ n[34380];
assign t[34381] = t[34380] ^ n[34381];
assign t[34382] = t[34381] ^ n[34382];
assign t[34383] = t[34382] ^ n[34383];
assign t[34384] = t[34383] ^ n[34384];
assign t[34385] = t[34384] ^ n[34385];
assign t[34386] = t[34385] ^ n[34386];
assign t[34387] = t[34386] ^ n[34387];
assign t[34388] = t[34387] ^ n[34388];
assign t[34389] = t[34388] ^ n[34389];
assign t[34390] = t[34389] ^ n[34390];
assign t[34391] = t[34390] ^ n[34391];
assign t[34392] = t[34391] ^ n[34392];
assign t[34393] = t[34392] ^ n[34393];
assign t[34394] = t[34393] ^ n[34394];
assign t[34395] = t[34394] ^ n[34395];
assign t[34396] = t[34395] ^ n[34396];
assign t[34397] = t[34396] ^ n[34397];
assign t[34398] = t[34397] ^ n[34398];
assign t[34399] = t[34398] ^ n[34399];
assign t[34400] = t[34399] ^ n[34400];
assign t[34401] = t[34400] ^ n[34401];
assign t[34402] = t[34401] ^ n[34402];
assign t[34403] = t[34402] ^ n[34403];
assign t[34404] = t[34403] ^ n[34404];
assign t[34405] = t[34404] ^ n[34405];
assign t[34406] = t[34405] ^ n[34406];
assign t[34407] = t[34406] ^ n[34407];
assign t[34408] = t[34407] ^ n[34408];
assign t[34409] = t[34408] ^ n[34409];
assign t[34410] = t[34409] ^ n[34410];
assign t[34411] = t[34410] ^ n[34411];
assign t[34412] = t[34411] ^ n[34412];
assign t[34413] = t[34412] ^ n[34413];
assign t[34414] = t[34413] ^ n[34414];
assign t[34415] = t[34414] ^ n[34415];
assign t[34416] = t[34415] ^ n[34416];
assign t[34417] = t[34416] ^ n[34417];
assign t[34418] = t[34417] ^ n[34418];
assign t[34419] = t[34418] ^ n[34419];
assign t[34420] = t[34419] ^ n[34420];
assign t[34421] = t[34420] ^ n[34421];
assign t[34422] = t[34421] ^ n[34422];
assign t[34423] = t[34422] ^ n[34423];
assign t[34424] = t[34423] ^ n[34424];
assign t[34425] = t[34424] ^ n[34425];
assign t[34426] = t[34425] ^ n[34426];
assign t[34427] = t[34426] ^ n[34427];
assign t[34428] = t[34427] ^ n[34428];
assign t[34429] = t[34428] ^ n[34429];
assign t[34430] = t[34429] ^ n[34430];
assign t[34431] = t[34430] ^ n[34431];
assign t[34432] = t[34431] ^ n[34432];
assign t[34433] = t[34432] ^ n[34433];
assign t[34434] = t[34433] ^ n[34434];
assign t[34435] = t[34434] ^ n[34435];
assign t[34436] = t[34435] ^ n[34436];
assign t[34437] = t[34436] ^ n[34437];
assign t[34438] = t[34437] ^ n[34438];
assign t[34439] = t[34438] ^ n[34439];
assign t[34440] = t[34439] ^ n[34440];
assign t[34441] = t[34440] ^ n[34441];
assign t[34442] = t[34441] ^ n[34442];
assign t[34443] = t[34442] ^ n[34443];
assign t[34444] = t[34443] ^ n[34444];
assign t[34445] = t[34444] ^ n[34445];
assign t[34446] = t[34445] ^ n[34446];
assign t[34447] = t[34446] ^ n[34447];
assign t[34448] = t[34447] ^ n[34448];
assign t[34449] = t[34448] ^ n[34449];
assign t[34450] = t[34449] ^ n[34450];
assign t[34451] = t[34450] ^ n[34451];
assign t[34452] = t[34451] ^ n[34452];
assign t[34453] = t[34452] ^ n[34453];
assign t[34454] = t[34453] ^ n[34454];
assign t[34455] = t[34454] ^ n[34455];
assign t[34456] = t[34455] ^ n[34456];
assign t[34457] = t[34456] ^ n[34457];
assign t[34458] = t[34457] ^ n[34458];
assign t[34459] = t[34458] ^ n[34459];
assign t[34460] = t[34459] ^ n[34460];
assign t[34461] = t[34460] ^ n[34461];
assign t[34462] = t[34461] ^ n[34462];
assign t[34463] = t[34462] ^ n[34463];
assign t[34464] = t[34463] ^ n[34464];
assign t[34465] = t[34464] ^ n[34465];
assign t[34466] = t[34465] ^ n[34466];
assign t[34467] = t[34466] ^ n[34467];
assign t[34468] = t[34467] ^ n[34468];
assign t[34469] = t[34468] ^ n[34469];
assign t[34470] = t[34469] ^ n[34470];
assign t[34471] = t[34470] ^ n[34471];
assign t[34472] = t[34471] ^ n[34472];
assign t[34473] = t[34472] ^ n[34473];
assign t[34474] = t[34473] ^ n[34474];
assign t[34475] = t[34474] ^ n[34475];
assign t[34476] = t[34475] ^ n[34476];
assign t[34477] = t[34476] ^ n[34477];
assign t[34478] = t[34477] ^ n[34478];
assign t[34479] = t[34478] ^ n[34479];
assign t[34480] = t[34479] ^ n[34480];
assign t[34481] = t[34480] ^ n[34481];
assign t[34482] = t[34481] ^ n[34482];
assign t[34483] = t[34482] ^ n[34483];
assign t[34484] = t[34483] ^ n[34484];
assign t[34485] = t[34484] ^ n[34485];
assign t[34486] = t[34485] ^ n[34486];
assign t[34487] = t[34486] ^ n[34487];
assign t[34488] = t[34487] ^ n[34488];
assign t[34489] = t[34488] ^ n[34489];
assign t[34490] = t[34489] ^ n[34490];
assign t[34491] = t[34490] ^ n[34491];
assign t[34492] = t[34491] ^ n[34492];
assign t[34493] = t[34492] ^ n[34493];
assign t[34494] = t[34493] ^ n[34494];
assign t[34495] = t[34494] ^ n[34495];
assign t[34496] = t[34495] ^ n[34496];
assign t[34497] = t[34496] ^ n[34497];
assign t[34498] = t[34497] ^ n[34498];
assign t[34499] = t[34498] ^ n[34499];
assign t[34500] = t[34499] ^ n[34500];
assign t[34501] = t[34500] ^ n[34501];
assign t[34502] = t[34501] ^ n[34502];
assign t[34503] = t[34502] ^ n[34503];
assign t[34504] = t[34503] ^ n[34504];
assign t[34505] = t[34504] ^ n[34505];
assign t[34506] = t[34505] ^ n[34506];
assign t[34507] = t[34506] ^ n[34507];
assign t[34508] = t[34507] ^ n[34508];
assign t[34509] = t[34508] ^ n[34509];
assign t[34510] = t[34509] ^ n[34510];
assign t[34511] = t[34510] ^ n[34511];
assign t[34512] = t[34511] ^ n[34512];
assign t[34513] = t[34512] ^ n[34513];
assign t[34514] = t[34513] ^ n[34514];
assign t[34515] = t[34514] ^ n[34515];
assign t[34516] = t[34515] ^ n[34516];
assign t[34517] = t[34516] ^ n[34517];
assign t[34518] = t[34517] ^ n[34518];
assign t[34519] = t[34518] ^ n[34519];
assign t[34520] = t[34519] ^ n[34520];
assign t[34521] = t[34520] ^ n[34521];
assign t[34522] = t[34521] ^ n[34522];
assign t[34523] = t[34522] ^ n[34523];
assign t[34524] = t[34523] ^ n[34524];
assign t[34525] = t[34524] ^ n[34525];
assign t[34526] = t[34525] ^ n[34526];
assign t[34527] = t[34526] ^ n[34527];
assign t[34528] = t[34527] ^ n[34528];
assign t[34529] = t[34528] ^ n[34529];
assign t[34530] = t[34529] ^ n[34530];
assign t[34531] = t[34530] ^ n[34531];
assign t[34532] = t[34531] ^ n[34532];
assign t[34533] = t[34532] ^ n[34533];
assign t[34534] = t[34533] ^ n[34534];
assign t[34535] = t[34534] ^ n[34535];
assign t[34536] = t[34535] ^ n[34536];
assign t[34537] = t[34536] ^ n[34537];
assign t[34538] = t[34537] ^ n[34538];
assign t[34539] = t[34538] ^ n[34539];
assign t[34540] = t[34539] ^ n[34540];
assign t[34541] = t[34540] ^ n[34541];
assign t[34542] = t[34541] ^ n[34542];
assign t[34543] = t[34542] ^ n[34543];
assign t[34544] = t[34543] ^ n[34544];
assign t[34545] = t[34544] ^ n[34545];
assign t[34546] = t[34545] ^ n[34546];
assign t[34547] = t[34546] ^ n[34547];
assign t[34548] = t[34547] ^ n[34548];
assign t[34549] = t[34548] ^ n[34549];
assign t[34550] = t[34549] ^ n[34550];
assign t[34551] = t[34550] ^ n[34551];
assign t[34552] = t[34551] ^ n[34552];
assign t[34553] = t[34552] ^ n[34553];
assign t[34554] = t[34553] ^ n[34554];
assign t[34555] = t[34554] ^ n[34555];
assign t[34556] = t[34555] ^ n[34556];
assign t[34557] = t[34556] ^ n[34557];
assign t[34558] = t[34557] ^ n[34558];
assign t[34559] = t[34558] ^ n[34559];
assign t[34560] = t[34559] ^ n[34560];
assign t[34561] = t[34560] ^ n[34561];
assign t[34562] = t[34561] ^ n[34562];
assign t[34563] = t[34562] ^ n[34563];
assign t[34564] = t[34563] ^ n[34564];
assign t[34565] = t[34564] ^ n[34565];
assign t[34566] = t[34565] ^ n[34566];
assign t[34567] = t[34566] ^ n[34567];
assign t[34568] = t[34567] ^ n[34568];
assign t[34569] = t[34568] ^ n[34569];
assign t[34570] = t[34569] ^ n[34570];
assign t[34571] = t[34570] ^ n[34571];
assign t[34572] = t[34571] ^ n[34572];
assign t[34573] = t[34572] ^ n[34573];
assign t[34574] = t[34573] ^ n[34574];
assign t[34575] = t[34574] ^ n[34575];
assign t[34576] = t[34575] ^ n[34576];
assign t[34577] = t[34576] ^ n[34577];
assign t[34578] = t[34577] ^ n[34578];
assign t[34579] = t[34578] ^ n[34579];
assign t[34580] = t[34579] ^ n[34580];
assign t[34581] = t[34580] ^ n[34581];
assign t[34582] = t[34581] ^ n[34582];
assign t[34583] = t[34582] ^ n[34583];
assign t[34584] = t[34583] ^ n[34584];
assign t[34585] = t[34584] ^ n[34585];
assign t[34586] = t[34585] ^ n[34586];
assign t[34587] = t[34586] ^ n[34587];
assign t[34588] = t[34587] ^ n[34588];
assign t[34589] = t[34588] ^ n[34589];
assign t[34590] = t[34589] ^ n[34590];
assign t[34591] = t[34590] ^ n[34591];
assign t[34592] = t[34591] ^ n[34592];
assign t[34593] = t[34592] ^ n[34593];
assign t[34594] = t[34593] ^ n[34594];
assign t[34595] = t[34594] ^ n[34595];
assign t[34596] = t[34595] ^ n[34596];
assign t[34597] = t[34596] ^ n[34597];
assign t[34598] = t[34597] ^ n[34598];
assign t[34599] = t[34598] ^ n[34599];
assign t[34600] = t[34599] ^ n[34600];
assign t[34601] = t[34600] ^ n[34601];
assign t[34602] = t[34601] ^ n[34602];
assign t[34603] = t[34602] ^ n[34603];
assign t[34604] = t[34603] ^ n[34604];
assign t[34605] = t[34604] ^ n[34605];
assign t[34606] = t[34605] ^ n[34606];
assign t[34607] = t[34606] ^ n[34607];
assign t[34608] = t[34607] ^ n[34608];
assign t[34609] = t[34608] ^ n[34609];
assign t[34610] = t[34609] ^ n[34610];
assign t[34611] = t[34610] ^ n[34611];
assign t[34612] = t[34611] ^ n[34612];
assign t[34613] = t[34612] ^ n[34613];
assign t[34614] = t[34613] ^ n[34614];
assign t[34615] = t[34614] ^ n[34615];
assign t[34616] = t[34615] ^ n[34616];
assign t[34617] = t[34616] ^ n[34617];
assign t[34618] = t[34617] ^ n[34618];
assign t[34619] = t[34618] ^ n[34619];
assign t[34620] = t[34619] ^ n[34620];
assign t[34621] = t[34620] ^ n[34621];
assign t[34622] = t[34621] ^ n[34622];
assign t[34623] = t[34622] ^ n[34623];
assign t[34624] = t[34623] ^ n[34624];
assign t[34625] = t[34624] ^ n[34625];
assign t[34626] = t[34625] ^ n[34626];
assign t[34627] = t[34626] ^ n[34627];
assign t[34628] = t[34627] ^ n[34628];
assign t[34629] = t[34628] ^ n[34629];
assign t[34630] = t[34629] ^ n[34630];
assign t[34631] = t[34630] ^ n[34631];
assign t[34632] = t[34631] ^ n[34632];
assign t[34633] = t[34632] ^ n[34633];
assign t[34634] = t[34633] ^ n[34634];
assign t[34635] = t[34634] ^ n[34635];
assign t[34636] = t[34635] ^ n[34636];
assign t[34637] = t[34636] ^ n[34637];
assign t[34638] = t[34637] ^ n[34638];
assign t[34639] = t[34638] ^ n[34639];
assign t[34640] = t[34639] ^ n[34640];
assign t[34641] = t[34640] ^ n[34641];
assign t[34642] = t[34641] ^ n[34642];
assign t[34643] = t[34642] ^ n[34643];
assign t[34644] = t[34643] ^ n[34644];
assign t[34645] = t[34644] ^ n[34645];
assign t[34646] = t[34645] ^ n[34646];
assign t[34647] = t[34646] ^ n[34647];
assign t[34648] = t[34647] ^ n[34648];
assign t[34649] = t[34648] ^ n[34649];
assign t[34650] = t[34649] ^ n[34650];
assign t[34651] = t[34650] ^ n[34651];
assign t[34652] = t[34651] ^ n[34652];
assign t[34653] = t[34652] ^ n[34653];
assign t[34654] = t[34653] ^ n[34654];
assign t[34655] = t[34654] ^ n[34655];
assign t[34656] = t[34655] ^ n[34656];
assign t[34657] = t[34656] ^ n[34657];
assign t[34658] = t[34657] ^ n[34658];
assign t[34659] = t[34658] ^ n[34659];
assign t[34660] = t[34659] ^ n[34660];
assign t[34661] = t[34660] ^ n[34661];
assign t[34662] = t[34661] ^ n[34662];
assign t[34663] = t[34662] ^ n[34663];
assign t[34664] = t[34663] ^ n[34664];
assign t[34665] = t[34664] ^ n[34665];
assign t[34666] = t[34665] ^ n[34666];
assign t[34667] = t[34666] ^ n[34667];
assign t[34668] = t[34667] ^ n[34668];
assign t[34669] = t[34668] ^ n[34669];
assign t[34670] = t[34669] ^ n[34670];
assign t[34671] = t[34670] ^ n[34671];
assign t[34672] = t[34671] ^ n[34672];
assign t[34673] = t[34672] ^ n[34673];
assign t[34674] = t[34673] ^ n[34674];
assign t[34675] = t[34674] ^ n[34675];
assign t[34676] = t[34675] ^ n[34676];
assign t[34677] = t[34676] ^ n[34677];
assign t[34678] = t[34677] ^ n[34678];
assign t[34679] = t[34678] ^ n[34679];
assign t[34680] = t[34679] ^ n[34680];
assign t[34681] = t[34680] ^ n[34681];
assign t[34682] = t[34681] ^ n[34682];
assign t[34683] = t[34682] ^ n[34683];
assign t[34684] = t[34683] ^ n[34684];
assign t[34685] = t[34684] ^ n[34685];
assign t[34686] = t[34685] ^ n[34686];
assign t[34687] = t[34686] ^ n[34687];
assign t[34688] = t[34687] ^ n[34688];
assign t[34689] = t[34688] ^ n[34689];
assign t[34690] = t[34689] ^ n[34690];
assign t[34691] = t[34690] ^ n[34691];
assign t[34692] = t[34691] ^ n[34692];
assign t[34693] = t[34692] ^ n[34693];
assign t[34694] = t[34693] ^ n[34694];
assign t[34695] = t[34694] ^ n[34695];
assign t[34696] = t[34695] ^ n[34696];
assign t[34697] = t[34696] ^ n[34697];
assign t[34698] = t[34697] ^ n[34698];
assign t[34699] = t[34698] ^ n[34699];
assign t[34700] = t[34699] ^ n[34700];
assign t[34701] = t[34700] ^ n[34701];
assign t[34702] = t[34701] ^ n[34702];
assign t[34703] = t[34702] ^ n[34703];
assign t[34704] = t[34703] ^ n[34704];
assign t[34705] = t[34704] ^ n[34705];
assign t[34706] = t[34705] ^ n[34706];
assign t[34707] = t[34706] ^ n[34707];
assign t[34708] = t[34707] ^ n[34708];
assign t[34709] = t[34708] ^ n[34709];
assign t[34710] = t[34709] ^ n[34710];
assign t[34711] = t[34710] ^ n[34711];
assign t[34712] = t[34711] ^ n[34712];
assign t[34713] = t[34712] ^ n[34713];
assign t[34714] = t[34713] ^ n[34714];
assign t[34715] = t[34714] ^ n[34715];
assign t[34716] = t[34715] ^ n[34716];
assign t[34717] = t[34716] ^ n[34717];
assign t[34718] = t[34717] ^ n[34718];
assign t[34719] = t[34718] ^ n[34719];
assign t[34720] = t[34719] ^ n[34720];
assign t[34721] = t[34720] ^ n[34721];
assign t[34722] = t[34721] ^ n[34722];
assign t[34723] = t[34722] ^ n[34723];
assign t[34724] = t[34723] ^ n[34724];
assign t[34725] = t[34724] ^ n[34725];
assign t[34726] = t[34725] ^ n[34726];
assign t[34727] = t[34726] ^ n[34727];
assign t[34728] = t[34727] ^ n[34728];
assign t[34729] = t[34728] ^ n[34729];
assign t[34730] = t[34729] ^ n[34730];
assign t[34731] = t[34730] ^ n[34731];
assign t[34732] = t[34731] ^ n[34732];
assign t[34733] = t[34732] ^ n[34733];
assign t[34734] = t[34733] ^ n[34734];
assign t[34735] = t[34734] ^ n[34735];
assign t[34736] = t[34735] ^ n[34736];
assign t[34737] = t[34736] ^ n[34737];
assign t[34738] = t[34737] ^ n[34738];
assign t[34739] = t[34738] ^ n[34739];
assign t[34740] = t[34739] ^ n[34740];
assign t[34741] = t[34740] ^ n[34741];
assign t[34742] = t[34741] ^ n[34742];
assign t[34743] = t[34742] ^ n[34743];
assign t[34744] = t[34743] ^ n[34744];
assign t[34745] = t[34744] ^ n[34745];
assign t[34746] = t[34745] ^ n[34746];
assign t[34747] = t[34746] ^ n[34747];
assign t[34748] = t[34747] ^ n[34748];
assign t[34749] = t[34748] ^ n[34749];
assign t[34750] = t[34749] ^ n[34750];
assign t[34751] = t[34750] ^ n[34751];
assign t[34752] = t[34751] ^ n[34752];
assign t[34753] = t[34752] ^ n[34753];
assign t[34754] = t[34753] ^ n[34754];
assign t[34755] = t[34754] ^ n[34755];
assign t[34756] = t[34755] ^ n[34756];
assign t[34757] = t[34756] ^ n[34757];
assign t[34758] = t[34757] ^ n[34758];
assign t[34759] = t[34758] ^ n[34759];
assign t[34760] = t[34759] ^ n[34760];
assign t[34761] = t[34760] ^ n[34761];
assign t[34762] = t[34761] ^ n[34762];
assign t[34763] = t[34762] ^ n[34763];
assign t[34764] = t[34763] ^ n[34764];
assign t[34765] = t[34764] ^ n[34765];
assign t[34766] = t[34765] ^ n[34766];
assign t[34767] = t[34766] ^ n[34767];
assign t[34768] = t[34767] ^ n[34768];
assign t[34769] = t[34768] ^ n[34769];
assign t[34770] = t[34769] ^ n[34770];
assign t[34771] = t[34770] ^ n[34771];
assign t[34772] = t[34771] ^ n[34772];
assign t[34773] = t[34772] ^ n[34773];
assign t[34774] = t[34773] ^ n[34774];
assign t[34775] = t[34774] ^ n[34775];
assign t[34776] = t[34775] ^ n[34776];
assign t[34777] = t[34776] ^ n[34777];
assign t[34778] = t[34777] ^ n[34778];
assign t[34779] = t[34778] ^ n[34779];
assign t[34780] = t[34779] ^ n[34780];
assign t[34781] = t[34780] ^ n[34781];
assign t[34782] = t[34781] ^ n[34782];
assign t[34783] = t[34782] ^ n[34783];
assign t[34784] = t[34783] ^ n[34784];
assign t[34785] = t[34784] ^ n[34785];
assign t[34786] = t[34785] ^ n[34786];
assign t[34787] = t[34786] ^ n[34787];
assign t[34788] = t[34787] ^ n[34788];
assign t[34789] = t[34788] ^ n[34789];
assign t[34790] = t[34789] ^ n[34790];
assign t[34791] = t[34790] ^ n[34791];
assign t[34792] = t[34791] ^ n[34792];
assign t[34793] = t[34792] ^ n[34793];
assign t[34794] = t[34793] ^ n[34794];
assign t[34795] = t[34794] ^ n[34795];
assign t[34796] = t[34795] ^ n[34796];
assign t[34797] = t[34796] ^ n[34797];
assign t[34798] = t[34797] ^ n[34798];
assign t[34799] = t[34798] ^ n[34799];
assign t[34800] = t[34799] ^ n[34800];
assign t[34801] = t[34800] ^ n[34801];
assign t[34802] = t[34801] ^ n[34802];
assign t[34803] = t[34802] ^ n[34803];
assign t[34804] = t[34803] ^ n[34804];
assign t[34805] = t[34804] ^ n[34805];
assign t[34806] = t[34805] ^ n[34806];
assign t[34807] = t[34806] ^ n[34807];
assign t[34808] = t[34807] ^ n[34808];
assign t[34809] = t[34808] ^ n[34809];
assign t[34810] = t[34809] ^ n[34810];
assign t[34811] = t[34810] ^ n[34811];
assign t[34812] = t[34811] ^ n[34812];
assign t[34813] = t[34812] ^ n[34813];
assign t[34814] = t[34813] ^ n[34814];
assign t[34815] = t[34814] ^ n[34815];
assign t[34816] = t[34815] ^ n[34816];
assign t[34817] = t[34816] ^ n[34817];
assign t[34818] = t[34817] ^ n[34818];
assign t[34819] = t[34818] ^ n[34819];
assign t[34820] = t[34819] ^ n[34820];
assign t[34821] = t[34820] ^ n[34821];
assign t[34822] = t[34821] ^ n[34822];
assign t[34823] = t[34822] ^ n[34823];
assign t[34824] = t[34823] ^ n[34824];
assign t[34825] = t[34824] ^ n[34825];
assign t[34826] = t[34825] ^ n[34826];
assign t[34827] = t[34826] ^ n[34827];
assign t[34828] = t[34827] ^ n[34828];
assign t[34829] = t[34828] ^ n[34829];
assign t[34830] = t[34829] ^ n[34830];
assign t[34831] = t[34830] ^ n[34831];
assign t[34832] = t[34831] ^ n[34832];
assign t[34833] = t[34832] ^ n[34833];
assign t[34834] = t[34833] ^ n[34834];
assign t[34835] = t[34834] ^ n[34835];
assign t[34836] = t[34835] ^ n[34836];
assign t[34837] = t[34836] ^ n[34837];
assign t[34838] = t[34837] ^ n[34838];
assign t[34839] = t[34838] ^ n[34839];
assign t[34840] = t[34839] ^ n[34840];
assign t[34841] = t[34840] ^ n[34841];
assign t[34842] = t[34841] ^ n[34842];
assign t[34843] = t[34842] ^ n[34843];
assign t[34844] = t[34843] ^ n[34844];
assign t[34845] = t[34844] ^ n[34845];
assign t[34846] = t[34845] ^ n[34846];
assign t[34847] = t[34846] ^ n[34847];
assign t[34848] = t[34847] ^ n[34848];
assign t[34849] = t[34848] ^ n[34849];
assign t[34850] = t[34849] ^ n[34850];
assign t[34851] = t[34850] ^ n[34851];
assign t[34852] = t[34851] ^ n[34852];
assign t[34853] = t[34852] ^ n[34853];
assign t[34854] = t[34853] ^ n[34854];
assign t[34855] = t[34854] ^ n[34855];
assign t[34856] = t[34855] ^ n[34856];
assign t[34857] = t[34856] ^ n[34857];
assign t[34858] = t[34857] ^ n[34858];
assign t[34859] = t[34858] ^ n[34859];
assign t[34860] = t[34859] ^ n[34860];
assign t[34861] = t[34860] ^ n[34861];
assign t[34862] = t[34861] ^ n[34862];
assign t[34863] = t[34862] ^ n[34863];
assign t[34864] = t[34863] ^ n[34864];
assign t[34865] = t[34864] ^ n[34865];
assign t[34866] = t[34865] ^ n[34866];
assign t[34867] = t[34866] ^ n[34867];
assign t[34868] = t[34867] ^ n[34868];
assign t[34869] = t[34868] ^ n[34869];
assign t[34870] = t[34869] ^ n[34870];
assign t[34871] = t[34870] ^ n[34871];
assign t[34872] = t[34871] ^ n[34872];
assign t[34873] = t[34872] ^ n[34873];
assign t[34874] = t[34873] ^ n[34874];
assign t[34875] = t[34874] ^ n[34875];
assign t[34876] = t[34875] ^ n[34876];
assign t[34877] = t[34876] ^ n[34877];
assign t[34878] = t[34877] ^ n[34878];
assign t[34879] = t[34878] ^ n[34879];
assign t[34880] = t[34879] ^ n[34880];
assign t[34881] = t[34880] ^ n[34881];
assign t[34882] = t[34881] ^ n[34882];
assign t[34883] = t[34882] ^ n[34883];
assign t[34884] = t[34883] ^ n[34884];
assign t[34885] = t[34884] ^ n[34885];
assign t[34886] = t[34885] ^ n[34886];
assign t[34887] = t[34886] ^ n[34887];
assign t[34888] = t[34887] ^ n[34888];
assign t[34889] = t[34888] ^ n[34889];
assign t[34890] = t[34889] ^ n[34890];
assign t[34891] = t[34890] ^ n[34891];
assign t[34892] = t[34891] ^ n[34892];
assign t[34893] = t[34892] ^ n[34893];
assign t[34894] = t[34893] ^ n[34894];
assign t[34895] = t[34894] ^ n[34895];
assign t[34896] = t[34895] ^ n[34896];
assign t[34897] = t[34896] ^ n[34897];
assign t[34898] = t[34897] ^ n[34898];
assign t[34899] = t[34898] ^ n[34899];
assign t[34900] = t[34899] ^ n[34900];
assign t[34901] = t[34900] ^ n[34901];
assign t[34902] = t[34901] ^ n[34902];
assign t[34903] = t[34902] ^ n[34903];
assign t[34904] = t[34903] ^ n[34904];
assign t[34905] = t[34904] ^ n[34905];
assign t[34906] = t[34905] ^ n[34906];
assign t[34907] = t[34906] ^ n[34907];
assign t[34908] = t[34907] ^ n[34908];
assign t[34909] = t[34908] ^ n[34909];
assign t[34910] = t[34909] ^ n[34910];
assign t[34911] = t[34910] ^ n[34911];
assign t[34912] = t[34911] ^ n[34912];
assign t[34913] = t[34912] ^ n[34913];
assign t[34914] = t[34913] ^ n[34914];
assign t[34915] = t[34914] ^ n[34915];
assign t[34916] = t[34915] ^ n[34916];
assign t[34917] = t[34916] ^ n[34917];
assign t[34918] = t[34917] ^ n[34918];
assign t[34919] = t[34918] ^ n[34919];
assign t[34920] = t[34919] ^ n[34920];
assign t[34921] = t[34920] ^ n[34921];
assign t[34922] = t[34921] ^ n[34922];
assign t[34923] = t[34922] ^ n[34923];
assign t[34924] = t[34923] ^ n[34924];
assign t[34925] = t[34924] ^ n[34925];
assign t[34926] = t[34925] ^ n[34926];
assign t[34927] = t[34926] ^ n[34927];
assign t[34928] = t[34927] ^ n[34928];
assign t[34929] = t[34928] ^ n[34929];
assign t[34930] = t[34929] ^ n[34930];
assign t[34931] = t[34930] ^ n[34931];
assign t[34932] = t[34931] ^ n[34932];
assign t[34933] = t[34932] ^ n[34933];
assign t[34934] = t[34933] ^ n[34934];
assign t[34935] = t[34934] ^ n[34935];
assign t[34936] = t[34935] ^ n[34936];
assign t[34937] = t[34936] ^ n[34937];
assign t[34938] = t[34937] ^ n[34938];
assign t[34939] = t[34938] ^ n[34939];
assign t[34940] = t[34939] ^ n[34940];
assign t[34941] = t[34940] ^ n[34941];
assign t[34942] = t[34941] ^ n[34942];
assign t[34943] = t[34942] ^ n[34943];
assign t[34944] = t[34943] ^ n[34944];
assign t[34945] = t[34944] ^ n[34945];
assign t[34946] = t[34945] ^ n[34946];
assign t[34947] = t[34946] ^ n[34947];
assign t[34948] = t[34947] ^ n[34948];
assign t[34949] = t[34948] ^ n[34949];
assign t[34950] = t[34949] ^ n[34950];
assign t[34951] = t[34950] ^ n[34951];
assign t[34952] = t[34951] ^ n[34952];
assign t[34953] = t[34952] ^ n[34953];
assign t[34954] = t[34953] ^ n[34954];
assign t[34955] = t[34954] ^ n[34955];
assign t[34956] = t[34955] ^ n[34956];
assign t[34957] = t[34956] ^ n[34957];
assign t[34958] = t[34957] ^ n[34958];
assign t[34959] = t[34958] ^ n[34959];
assign t[34960] = t[34959] ^ n[34960];
assign t[34961] = t[34960] ^ n[34961];
assign t[34962] = t[34961] ^ n[34962];
assign t[34963] = t[34962] ^ n[34963];
assign t[34964] = t[34963] ^ n[34964];
assign t[34965] = t[34964] ^ n[34965];
assign t[34966] = t[34965] ^ n[34966];
assign t[34967] = t[34966] ^ n[34967];
assign t[34968] = t[34967] ^ n[34968];
assign t[34969] = t[34968] ^ n[34969];
assign t[34970] = t[34969] ^ n[34970];
assign t[34971] = t[34970] ^ n[34971];
assign t[34972] = t[34971] ^ n[34972];
assign t[34973] = t[34972] ^ n[34973];
assign t[34974] = t[34973] ^ n[34974];
assign t[34975] = t[34974] ^ n[34975];
assign t[34976] = t[34975] ^ n[34976];
assign t[34977] = t[34976] ^ n[34977];
assign t[34978] = t[34977] ^ n[34978];
assign t[34979] = t[34978] ^ n[34979];
assign t[34980] = t[34979] ^ n[34980];
assign t[34981] = t[34980] ^ n[34981];
assign t[34982] = t[34981] ^ n[34982];
assign t[34983] = t[34982] ^ n[34983];
assign t[34984] = t[34983] ^ n[34984];
assign t[34985] = t[34984] ^ n[34985];
assign t[34986] = t[34985] ^ n[34986];
assign t[34987] = t[34986] ^ n[34987];
assign t[34988] = t[34987] ^ n[34988];
assign t[34989] = t[34988] ^ n[34989];
assign t[34990] = t[34989] ^ n[34990];
assign t[34991] = t[34990] ^ n[34991];
assign t[34992] = t[34991] ^ n[34992];
assign t[34993] = t[34992] ^ n[34993];
assign t[34994] = t[34993] ^ n[34994];
assign t[34995] = t[34994] ^ n[34995];
assign t[34996] = t[34995] ^ n[34996];
assign t[34997] = t[34996] ^ n[34997];
assign t[34998] = t[34997] ^ n[34998];
assign t[34999] = t[34998] ^ n[34999];
assign t[35000] = t[34999] ^ n[35000];
assign t[35001] = t[35000] ^ n[35001];
assign t[35002] = t[35001] ^ n[35002];
assign t[35003] = t[35002] ^ n[35003];
assign t[35004] = t[35003] ^ n[35004];
assign t[35005] = t[35004] ^ n[35005];
assign t[35006] = t[35005] ^ n[35006];
assign t[35007] = t[35006] ^ n[35007];
assign t[35008] = t[35007] ^ n[35008];
assign t[35009] = t[35008] ^ n[35009];
assign t[35010] = t[35009] ^ n[35010];
assign t[35011] = t[35010] ^ n[35011];
assign t[35012] = t[35011] ^ n[35012];
assign t[35013] = t[35012] ^ n[35013];
assign t[35014] = t[35013] ^ n[35014];
assign t[35015] = t[35014] ^ n[35015];
assign t[35016] = t[35015] ^ n[35016];
assign t[35017] = t[35016] ^ n[35017];
assign t[35018] = t[35017] ^ n[35018];
assign t[35019] = t[35018] ^ n[35019];
assign t[35020] = t[35019] ^ n[35020];
assign t[35021] = t[35020] ^ n[35021];
assign t[35022] = t[35021] ^ n[35022];
assign t[35023] = t[35022] ^ n[35023];
assign t[35024] = t[35023] ^ n[35024];
assign t[35025] = t[35024] ^ n[35025];
assign t[35026] = t[35025] ^ n[35026];
assign t[35027] = t[35026] ^ n[35027];
assign t[35028] = t[35027] ^ n[35028];
assign t[35029] = t[35028] ^ n[35029];
assign t[35030] = t[35029] ^ n[35030];
assign t[35031] = t[35030] ^ n[35031];
assign t[35032] = t[35031] ^ n[35032];
assign t[35033] = t[35032] ^ n[35033];
assign t[35034] = t[35033] ^ n[35034];
assign t[35035] = t[35034] ^ n[35035];
assign t[35036] = t[35035] ^ n[35036];
assign t[35037] = t[35036] ^ n[35037];
assign t[35038] = t[35037] ^ n[35038];
assign t[35039] = t[35038] ^ n[35039];
assign t[35040] = t[35039] ^ n[35040];
assign t[35041] = t[35040] ^ n[35041];
assign t[35042] = t[35041] ^ n[35042];
assign t[35043] = t[35042] ^ n[35043];
assign t[35044] = t[35043] ^ n[35044];
assign t[35045] = t[35044] ^ n[35045];
assign t[35046] = t[35045] ^ n[35046];
assign t[35047] = t[35046] ^ n[35047];
assign t[35048] = t[35047] ^ n[35048];
assign t[35049] = t[35048] ^ n[35049];
assign t[35050] = t[35049] ^ n[35050];
assign t[35051] = t[35050] ^ n[35051];
assign t[35052] = t[35051] ^ n[35052];
assign t[35053] = t[35052] ^ n[35053];
assign t[35054] = t[35053] ^ n[35054];
assign t[35055] = t[35054] ^ n[35055];
assign t[35056] = t[35055] ^ n[35056];
assign t[35057] = t[35056] ^ n[35057];
assign t[35058] = t[35057] ^ n[35058];
assign t[35059] = t[35058] ^ n[35059];
assign t[35060] = t[35059] ^ n[35060];
assign t[35061] = t[35060] ^ n[35061];
assign t[35062] = t[35061] ^ n[35062];
assign t[35063] = t[35062] ^ n[35063];
assign t[35064] = t[35063] ^ n[35064];
assign t[35065] = t[35064] ^ n[35065];
assign t[35066] = t[35065] ^ n[35066];
assign t[35067] = t[35066] ^ n[35067];
assign t[35068] = t[35067] ^ n[35068];
assign t[35069] = t[35068] ^ n[35069];
assign t[35070] = t[35069] ^ n[35070];
assign t[35071] = t[35070] ^ n[35071];
assign t[35072] = t[35071] ^ n[35072];
assign t[35073] = t[35072] ^ n[35073];
assign t[35074] = t[35073] ^ n[35074];
assign t[35075] = t[35074] ^ n[35075];
assign t[35076] = t[35075] ^ n[35076];
assign t[35077] = t[35076] ^ n[35077];
assign t[35078] = t[35077] ^ n[35078];
assign t[35079] = t[35078] ^ n[35079];
assign t[35080] = t[35079] ^ n[35080];
assign t[35081] = t[35080] ^ n[35081];
assign t[35082] = t[35081] ^ n[35082];
assign t[35083] = t[35082] ^ n[35083];
assign t[35084] = t[35083] ^ n[35084];
assign t[35085] = t[35084] ^ n[35085];
assign t[35086] = t[35085] ^ n[35086];
assign t[35087] = t[35086] ^ n[35087];
assign t[35088] = t[35087] ^ n[35088];
assign t[35089] = t[35088] ^ n[35089];
assign t[35090] = t[35089] ^ n[35090];
assign t[35091] = t[35090] ^ n[35091];
assign t[35092] = t[35091] ^ n[35092];
assign t[35093] = t[35092] ^ n[35093];
assign t[35094] = t[35093] ^ n[35094];
assign t[35095] = t[35094] ^ n[35095];
assign t[35096] = t[35095] ^ n[35096];
assign t[35097] = t[35096] ^ n[35097];
assign t[35098] = t[35097] ^ n[35098];
assign t[35099] = t[35098] ^ n[35099];
assign t[35100] = t[35099] ^ n[35100];
assign t[35101] = t[35100] ^ n[35101];
assign t[35102] = t[35101] ^ n[35102];
assign t[35103] = t[35102] ^ n[35103];
assign t[35104] = t[35103] ^ n[35104];
assign t[35105] = t[35104] ^ n[35105];
assign t[35106] = t[35105] ^ n[35106];
assign t[35107] = t[35106] ^ n[35107];
assign t[35108] = t[35107] ^ n[35108];
assign t[35109] = t[35108] ^ n[35109];
assign t[35110] = t[35109] ^ n[35110];
assign t[35111] = t[35110] ^ n[35111];
assign t[35112] = t[35111] ^ n[35112];
assign t[35113] = t[35112] ^ n[35113];
assign t[35114] = t[35113] ^ n[35114];
assign t[35115] = t[35114] ^ n[35115];
assign t[35116] = t[35115] ^ n[35116];
assign t[35117] = t[35116] ^ n[35117];
assign t[35118] = t[35117] ^ n[35118];
assign t[35119] = t[35118] ^ n[35119];
assign t[35120] = t[35119] ^ n[35120];
assign t[35121] = t[35120] ^ n[35121];
assign t[35122] = t[35121] ^ n[35122];
assign t[35123] = t[35122] ^ n[35123];
assign t[35124] = t[35123] ^ n[35124];
assign t[35125] = t[35124] ^ n[35125];
assign t[35126] = t[35125] ^ n[35126];
assign t[35127] = t[35126] ^ n[35127];
assign t[35128] = t[35127] ^ n[35128];
assign t[35129] = t[35128] ^ n[35129];
assign t[35130] = t[35129] ^ n[35130];
assign t[35131] = t[35130] ^ n[35131];
assign t[35132] = t[35131] ^ n[35132];
assign t[35133] = t[35132] ^ n[35133];
assign t[35134] = t[35133] ^ n[35134];
assign t[35135] = t[35134] ^ n[35135];
assign t[35136] = t[35135] ^ n[35136];
assign t[35137] = t[35136] ^ n[35137];
assign t[35138] = t[35137] ^ n[35138];
assign t[35139] = t[35138] ^ n[35139];
assign t[35140] = t[35139] ^ n[35140];
assign t[35141] = t[35140] ^ n[35141];
assign t[35142] = t[35141] ^ n[35142];
assign t[35143] = t[35142] ^ n[35143];
assign t[35144] = t[35143] ^ n[35144];
assign t[35145] = t[35144] ^ n[35145];
assign t[35146] = t[35145] ^ n[35146];
assign t[35147] = t[35146] ^ n[35147];
assign t[35148] = t[35147] ^ n[35148];
assign t[35149] = t[35148] ^ n[35149];
assign t[35150] = t[35149] ^ n[35150];
assign t[35151] = t[35150] ^ n[35151];
assign t[35152] = t[35151] ^ n[35152];
assign t[35153] = t[35152] ^ n[35153];
assign t[35154] = t[35153] ^ n[35154];
assign t[35155] = t[35154] ^ n[35155];
assign t[35156] = t[35155] ^ n[35156];
assign t[35157] = t[35156] ^ n[35157];
assign t[35158] = t[35157] ^ n[35158];
assign t[35159] = t[35158] ^ n[35159];
assign t[35160] = t[35159] ^ n[35160];
assign t[35161] = t[35160] ^ n[35161];
assign t[35162] = t[35161] ^ n[35162];
assign t[35163] = t[35162] ^ n[35163];
assign t[35164] = t[35163] ^ n[35164];
assign t[35165] = t[35164] ^ n[35165];
assign t[35166] = t[35165] ^ n[35166];
assign t[35167] = t[35166] ^ n[35167];
assign t[35168] = t[35167] ^ n[35168];
assign t[35169] = t[35168] ^ n[35169];
assign t[35170] = t[35169] ^ n[35170];
assign t[35171] = t[35170] ^ n[35171];
assign t[35172] = t[35171] ^ n[35172];
assign t[35173] = t[35172] ^ n[35173];
assign t[35174] = t[35173] ^ n[35174];
assign t[35175] = t[35174] ^ n[35175];
assign t[35176] = t[35175] ^ n[35176];
assign t[35177] = t[35176] ^ n[35177];
assign t[35178] = t[35177] ^ n[35178];
assign t[35179] = t[35178] ^ n[35179];
assign t[35180] = t[35179] ^ n[35180];
assign t[35181] = t[35180] ^ n[35181];
assign t[35182] = t[35181] ^ n[35182];
assign t[35183] = t[35182] ^ n[35183];
assign t[35184] = t[35183] ^ n[35184];
assign t[35185] = t[35184] ^ n[35185];
assign t[35186] = t[35185] ^ n[35186];
assign t[35187] = t[35186] ^ n[35187];
assign t[35188] = t[35187] ^ n[35188];
assign t[35189] = t[35188] ^ n[35189];
assign t[35190] = t[35189] ^ n[35190];
assign t[35191] = t[35190] ^ n[35191];
assign t[35192] = t[35191] ^ n[35192];
assign t[35193] = t[35192] ^ n[35193];
assign t[35194] = t[35193] ^ n[35194];
assign t[35195] = t[35194] ^ n[35195];
assign t[35196] = t[35195] ^ n[35196];
assign t[35197] = t[35196] ^ n[35197];
assign t[35198] = t[35197] ^ n[35198];
assign t[35199] = t[35198] ^ n[35199];
assign t[35200] = t[35199] ^ n[35200];
assign t[35201] = t[35200] ^ n[35201];
assign t[35202] = t[35201] ^ n[35202];
assign t[35203] = t[35202] ^ n[35203];
assign t[35204] = t[35203] ^ n[35204];
assign t[35205] = t[35204] ^ n[35205];
assign t[35206] = t[35205] ^ n[35206];
assign t[35207] = t[35206] ^ n[35207];
assign t[35208] = t[35207] ^ n[35208];
assign t[35209] = t[35208] ^ n[35209];
assign t[35210] = t[35209] ^ n[35210];
assign t[35211] = t[35210] ^ n[35211];
assign t[35212] = t[35211] ^ n[35212];
assign t[35213] = t[35212] ^ n[35213];
assign t[35214] = t[35213] ^ n[35214];
assign t[35215] = t[35214] ^ n[35215];
assign t[35216] = t[35215] ^ n[35216];
assign t[35217] = t[35216] ^ n[35217];
assign t[35218] = t[35217] ^ n[35218];
assign t[35219] = t[35218] ^ n[35219];
assign t[35220] = t[35219] ^ n[35220];
assign t[35221] = t[35220] ^ n[35221];
assign t[35222] = t[35221] ^ n[35222];
assign t[35223] = t[35222] ^ n[35223];
assign t[35224] = t[35223] ^ n[35224];
assign t[35225] = t[35224] ^ n[35225];
assign t[35226] = t[35225] ^ n[35226];
assign t[35227] = t[35226] ^ n[35227];
assign t[35228] = t[35227] ^ n[35228];
assign t[35229] = t[35228] ^ n[35229];
assign t[35230] = t[35229] ^ n[35230];
assign t[35231] = t[35230] ^ n[35231];
assign t[35232] = t[35231] ^ n[35232];
assign t[35233] = t[35232] ^ n[35233];
assign t[35234] = t[35233] ^ n[35234];
assign t[35235] = t[35234] ^ n[35235];
assign t[35236] = t[35235] ^ n[35236];
assign t[35237] = t[35236] ^ n[35237];
assign t[35238] = t[35237] ^ n[35238];
assign t[35239] = t[35238] ^ n[35239];
assign t[35240] = t[35239] ^ n[35240];
assign t[35241] = t[35240] ^ n[35241];
assign t[35242] = t[35241] ^ n[35242];
assign t[35243] = t[35242] ^ n[35243];
assign t[35244] = t[35243] ^ n[35244];
assign t[35245] = t[35244] ^ n[35245];
assign t[35246] = t[35245] ^ n[35246];
assign t[35247] = t[35246] ^ n[35247];
assign t[35248] = t[35247] ^ n[35248];
assign t[35249] = t[35248] ^ n[35249];
assign t[35250] = t[35249] ^ n[35250];
assign t[35251] = t[35250] ^ n[35251];
assign t[35252] = t[35251] ^ n[35252];
assign t[35253] = t[35252] ^ n[35253];
assign t[35254] = t[35253] ^ n[35254];
assign t[35255] = t[35254] ^ n[35255];
assign t[35256] = t[35255] ^ n[35256];
assign t[35257] = t[35256] ^ n[35257];
assign t[35258] = t[35257] ^ n[35258];
assign t[35259] = t[35258] ^ n[35259];
assign t[35260] = t[35259] ^ n[35260];
assign t[35261] = t[35260] ^ n[35261];
assign t[35262] = t[35261] ^ n[35262];
assign t[35263] = t[35262] ^ n[35263];
assign t[35264] = t[35263] ^ n[35264];
assign t[35265] = t[35264] ^ n[35265];
assign t[35266] = t[35265] ^ n[35266];
assign t[35267] = t[35266] ^ n[35267];
assign t[35268] = t[35267] ^ n[35268];
assign t[35269] = t[35268] ^ n[35269];
assign t[35270] = t[35269] ^ n[35270];
assign t[35271] = t[35270] ^ n[35271];
assign t[35272] = t[35271] ^ n[35272];
assign t[35273] = t[35272] ^ n[35273];
assign t[35274] = t[35273] ^ n[35274];
assign t[35275] = t[35274] ^ n[35275];
assign t[35276] = t[35275] ^ n[35276];
assign t[35277] = t[35276] ^ n[35277];
assign t[35278] = t[35277] ^ n[35278];
assign t[35279] = t[35278] ^ n[35279];
assign t[35280] = t[35279] ^ n[35280];
assign t[35281] = t[35280] ^ n[35281];
assign t[35282] = t[35281] ^ n[35282];
assign t[35283] = t[35282] ^ n[35283];
assign t[35284] = t[35283] ^ n[35284];
assign t[35285] = t[35284] ^ n[35285];
assign t[35286] = t[35285] ^ n[35286];
assign t[35287] = t[35286] ^ n[35287];
assign t[35288] = t[35287] ^ n[35288];
assign t[35289] = t[35288] ^ n[35289];
assign t[35290] = t[35289] ^ n[35290];
assign t[35291] = t[35290] ^ n[35291];
assign t[35292] = t[35291] ^ n[35292];
assign t[35293] = t[35292] ^ n[35293];
assign t[35294] = t[35293] ^ n[35294];
assign t[35295] = t[35294] ^ n[35295];
assign t[35296] = t[35295] ^ n[35296];
assign t[35297] = t[35296] ^ n[35297];
assign t[35298] = t[35297] ^ n[35298];
assign t[35299] = t[35298] ^ n[35299];
assign t[35300] = t[35299] ^ n[35300];
assign t[35301] = t[35300] ^ n[35301];
assign t[35302] = t[35301] ^ n[35302];
assign t[35303] = t[35302] ^ n[35303];
assign t[35304] = t[35303] ^ n[35304];
assign t[35305] = t[35304] ^ n[35305];
assign t[35306] = t[35305] ^ n[35306];
assign t[35307] = t[35306] ^ n[35307];
assign t[35308] = t[35307] ^ n[35308];
assign t[35309] = t[35308] ^ n[35309];
assign t[35310] = t[35309] ^ n[35310];
assign t[35311] = t[35310] ^ n[35311];
assign t[35312] = t[35311] ^ n[35312];
assign t[35313] = t[35312] ^ n[35313];
assign t[35314] = t[35313] ^ n[35314];
assign t[35315] = t[35314] ^ n[35315];
assign t[35316] = t[35315] ^ n[35316];
assign t[35317] = t[35316] ^ n[35317];
assign t[35318] = t[35317] ^ n[35318];
assign t[35319] = t[35318] ^ n[35319];
assign t[35320] = t[35319] ^ n[35320];
assign t[35321] = t[35320] ^ n[35321];
assign t[35322] = t[35321] ^ n[35322];
assign t[35323] = t[35322] ^ n[35323];
assign t[35324] = t[35323] ^ n[35324];
assign t[35325] = t[35324] ^ n[35325];
assign t[35326] = t[35325] ^ n[35326];
assign t[35327] = t[35326] ^ n[35327];
assign t[35328] = t[35327] ^ n[35328];
assign t[35329] = t[35328] ^ n[35329];
assign t[35330] = t[35329] ^ n[35330];
assign t[35331] = t[35330] ^ n[35331];
assign t[35332] = t[35331] ^ n[35332];
assign t[35333] = t[35332] ^ n[35333];
assign t[35334] = t[35333] ^ n[35334];
assign t[35335] = t[35334] ^ n[35335];
assign t[35336] = t[35335] ^ n[35336];
assign t[35337] = t[35336] ^ n[35337];
assign t[35338] = t[35337] ^ n[35338];
assign t[35339] = t[35338] ^ n[35339];
assign t[35340] = t[35339] ^ n[35340];
assign t[35341] = t[35340] ^ n[35341];
assign t[35342] = t[35341] ^ n[35342];
assign t[35343] = t[35342] ^ n[35343];
assign t[35344] = t[35343] ^ n[35344];
assign t[35345] = t[35344] ^ n[35345];
assign t[35346] = t[35345] ^ n[35346];
assign t[35347] = t[35346] ^ n[35347];
assign t[35348] = t[35347] ^ n[35348];
assign t[35349] = t[35348] ^ n[35349];
assign t[35350] = t[35349] ^ n[35350];
assign t[35351] = t[35350] ^ n[35351];
assign t[35352] = t[35351] ^ n[35352];
assign t[35353] = t[35352] ^ n[35353];
assign t[35354] = t[35353] ^ n[35354];
assign t[35355] = t[35354] ^ n[35355];
assign t[35356] = t[35355] ^ n[35356];
assign t[35357] = t[35356] ^ n[35357];
assign t[35358] = t[35357] ^ n[35358];
assign t[35359] = t[35358] ^ n[35359];
assign t[35360] = t[35359] ^ n[35360];
assign t[35361] = t[35360] ^ n[35361];
assign t[35362] = t[35361] ^ n[35362];
assign t[35363] = t[35362] ^ n[35363];
assign t[35364] = t[35363] ^ n[35364];
assign t[35365] = t[35364] ^ n[35365];
assign t[35366] = t[35365] ^ n[35366];
assign t[35367] = t[35366] ^ n[35367];
assign t[35368] = t[35367] ^ n[35368];
assign t[35369] = t[35368] ^ n[35369];
assign t[35370] = t[35369] ^ n[35370];
assign t[35371] = t[35370] ^ n[35371];
assign t[35372] = t[35371] ^ n[35372];
assign t[35373] = t[35372] ^ n[35373];
assign t[35374] = t[35373] ^ n[35374];
assign t[35375] = t[35374] ^ n[35375];
assign t[35376] = t[35375] ^ n[35376];
assign t[35377] = t[35376] ^ n[35377];
assign t[35378] = t[35377] ^ n[35378];
assign t[35379] = t[35378] ^ n[35379];
assign t[35380] = t[35379] ^ n[35380];
assign t[35381] = t[35380] ^ n[35381];
assign t[35382] = t[35381] ^ n[35382];
assign t[35383] = t[35382] ^ n[35383];
assign t[35384] = t[35383] ^ n[35384];
assign t[35385] = t[35384] ^ n[35385];
assign t[35386] = t[35385] ^ n[35386];
assign t[35387] = t[35386] ^ n[35387];
assign t[35388] = t[35387] ^ n[35388];
assign t[35389] = t[35388] ^ n[35389];
assign t[35390] = t[35389] ^ n[35390];
assign t[35391] = t[35390] ^ n[35391];
assign t[35392] = t[35391] ^ n[35392];
assign t[35393] = t[35392] ^ n[35393];
assign t[35394] = t[35393] ^ n[35394];
assign t[35395] = t[35394] ^ n[35395];
assign t[35396] = t[35395] ^ n[35396];
assign t[35397] = t[35396] ^ n[35397];
assign t[35398] = t[35397] ^ n[35398];
assign t[35399] = t[35398] ^ n[35399];
assign t[35400] = t[35399] ^ n[35400];
assign t[35401] = t[35400] ^ n[35401];
assign t[35402] = t[35401] ^ n[35402];
assign t[35403] = t[35402] ^ n[35403];
assign t[35404] = t[35403] ^ n[35404];
assign t[35405] = t[35404] ^ n[35405];
assign t[35406] = t[35405] ^ n[35406];
assign t[35407] = t[35406] ^ n[35407];
assign t[35408] = t[35407] ^ n[35408];
assign t[35409] = t[35408] ^ n[35409];
assign t[35410] = t[35409] ^ n[35410];
assign t[35411] = t[35410] ^ n[35411];
assign t[35412] = t[35411] ^ n[35412];
assign t[35413] = t[35412] ^ n[35413];
assign t[35414] = t[35413] ^ n[35414];
assign t[35415] = t[35414] ^ n[35415];
assign t[35416] = t[35415] ^ n[35416];
assign t[35417] = t[35416] ^ n[35417];
assign t[35418] = t[35417] ^ n[35418];
assign t[35419] = t[35418] ^ n[35419];
assign t[35420] = t[35419] ^ n[35420];
assign t[35421] = t[35420] ^ n[35421];
assign t[35422] = t[35421] ^ n[35422];
assign t[35423] = t[35422] ^ n[35423];
assign t[35424] = t[35423] ^ n[35424];
assign t[35425] = t[35424] ^ n[35425];
assign t[35426] = t[35425] ^ n[35426];
assign t[35427] = t[35426] ^ n[35427];
assign t[35428] = t[35427] ^ n[35428];
assign t[35429] = t[35428] ^ n[35429];
assign t[35430] = t[35429] ^ n[35430];
assign t[35431] = t[35430] ^ n[35431];
assign t[35432] = t[35431] ^ n[35432];
assign t[35433] = t[35432] ^ n[35433];
assign t[35434] = t[35433] ^ n[35434];
assign t[35435] = t[35434] ^ n[35435];
assign t[35436] = t[35435] ^ n[35436];
assign t[35437] = t[35436] ^ n[35437];
assign t[35438] = t[35437] ^ n[35438];
assign t[35439] = t[35438] ^ n[35439];
assign t[35440] = t[35439] ^ n[35440];
assign t[35441] = t[35440] ^ n[35441];
assign t[35442] = t[35441] ^ n[35442];
assign t[35443] = t[35442] ^ n[35443];
assign t[35444] = t[35443] ^ n[35444];
assign t[35445] = t[35444] ^ n[35445];
assign t[35446] = t[35445] ^ n[35446];
assign t[35447] = t[35446] ^ n[35447];
assign t[35448] = t[35447] ^ n[35448];
assign t[35449] = t[35448] ^ n[35449];
assign t[35450] = t[35449] ^ n[35450];
assign t[35451] = t[35450] ^ n[35451];
assign t[35452] = t[35451] ^ n[35452];
assign t[35453] = t[35452] ^ n[35453];
assign t[35454] = t[35453] ^ n[35454];
assign t[35455] = t[35454] ^ n[35455];
assign t[35456] = t[35455] ^ n[35456];
assign t[35457] = t[35456] ^ n[35457];
assign t[35458] = t[35457] ^ n[35458];
assign t[35459] = t[35458] ^ n[35459];
assign t[35460] = t[35459] ^ n[35460];
assign t[35461] = t[35460] ^ n[35461];
assign t[35462] = t[35461] ^ n[35462];
assign t[35463] = t[35462] ^ n[35463];
assign t[35464] = t[35463] ^ n[35464];
assign t[35465] = t[35464] ^ n[35465];
assign t[35466] = t[35465] ^ n[35466];
assign t[35467] = t[35466] ^ n[35467];
assign t[35468] = t[35467] ^ n[35468];
assign t[35469] = t[35468] ^ n[35469];
assign t[35470] = t[35469] ^ n[35470];
assign t[35471] = t[35470] ^ n[35471];
assign t[35472] = t[35471] ^ n[35472];
assign t[35473] = t[35472] ^ n[35473];
assign t[35474] = t[35473] ^ n[35474];
assign t[35475] = t[35474] ^ n[35475];
assign t[35476] = t[35475] ^ n[35476];
assign t[35477] = t[35476] ^ n[35477];
assign t[35478] = t[35477] ^ n[35478];
assign t[35479] = t[35478] ^ n[35479];
assign t[35480] = t[35479] ^ n[35480];
assign t[35481] = t[35480] ^ n[35481];
assign t[35482] = t[35481] ^ n[35482];
assign t[35483] = t[35482] ^ n[35483];
assign t[35484] = t[35483] ^ n[35484];
assign t[35485] = t[35484] ^ n[35485];
assign t[35486] = t[35485] ^ n[35486];
assign t[35487] = t[35486] ^ n[35487];
assign t[35488] = t[35487] ^ n[35488];
assign t[35489] = t[35488] ^ n[35489];
assign t[35490] = t[35489] ^ n[35490];
assign t[35491] = t[35490] ^ n[35491];
assign t[35492] = t[35491] ^ n[35492];
assign t[35493] = t[35492] ^ n[35493];
assign t[35494] = t[35493] ^ n[35494];
assign t[35495] = t[35494] ^ n[35495];
assign t[35496] = t[35495] ^ n[35496];
assign t[35497] = t[35496] ^ n[35497];
assign t[35498] = t[35497] ^ n[35498];
assign t[35499] = t[35498] ^ n[35499];
assign t[35500] = t[35499] ^ n[35500];
assign t[35501] = t[35500] ^ n[35501];
assign t[35502] = t[35501] ^ n[35502];
assign t[35503] = t[35502] ^ n[35503];
assign t[35504] = t[35503] ^ n[35504];
assign t[35505] = t[35504] ^ n[35505];
assign t[35506] = t[35505] ^ n[35506];
assign t[35507] = t[35506] ^ n[35507];
assign t[35508] = t[35507] ^ n[35508];
assign t[35509] = t[35508] ^ n[35509];
assign t[35510] = t[35509] ^ n[35510];
assign t[35511] = t[35510] ^ n[35511];
assign t[35512] = t[35511] ^ n[35512];
assign t[35513] = t[35512] ^ n[35513];
assign t[35514] = t[35513] ^ n[35514];
assign t[35515] = t[35514] ^ n[35515];
assign t[35516] = t[35515] ^ n[35516];
assign t[35517] = t[35516] ^ n[35517];
assign t[35518] = t[35517] ^ n[35518];
assign t[35519] = t[35518] ^ n[35519];
assign t[35520] = t[35519] ^ n[35520];
assign t[35521] = t[35520] ^ n[35521];
assign t[35522] = t[35521] ^ n[35522];
assign t[35523] = t[35522] ^ n[35523];
assign t[35524] = t[35523] ^ n[35524];
assign t[35525] = t[35524] ^ n[35525];
assign t[35526] = t[35525] ^ n[35526];
assign t[35527] = t[35526] ^ n[35527];
assign t[35528] = t[35527] ^ n[35528];
assign t[35529] = t[35528] ^ n[35529];
assign t[35530] = t[35529] ^ n[35530];
assign t[35531] = t[35530] ^ n[35531];
assign t[35532] = t[35531] ^ n[35532];
assign t[35533] = t[35532] ^ n[35533];
assign t[35534] = t[35533] ^ n[35534];
assign t[35535] = t[35534] ^ n[35535];
assign t[35536] = t[35535] ^ n[35536];
assign t[35537] = t[35536] ^ n[35537];
assign t[35538] = t[35537] ^ n[35538];
assign t[35539] = t[35538] ^ n[35539];
assign t[35540] = t[35539] ^ n[35540];
assign t[35541] = t[35540] ^ n[35541];
assign t[35542] = t[35541] ^ n[35542];
assign t[35543] = t[35542] ^ n[35543];
assign t[35544] = t[35543] ^ n[35544];
assign t[35545] = t[35544] ^ n[35545];
assign t[35546] = t[35545] ^ n[35546];
assign t[35547] = t[35546] ^ n[35547];
assign t[35548] = t[35547] ^ n[35548];
assign t[35549] = t[35548] ^ n[35549];
assign t[35550] = t[35549] ^ n[35550];
assign t[35551] = t[35550] ^ n[35551];
assign t[35552] = t[35551] ^ n[35552];
assign t[35553] = t[35552] ^ n[35553];
assign t[35554] = t[35553] ^ n[35554];
assign t[35555] = t[35554] ^ n[35555];
assign t[35556] = t[35555] ^ n[35556];
assign t[35557] = t[35556] ^ n[35557];
assign t[35558] = t[35557] ^ n[35558];
assign t[35559] = t[35558] ^ n[35559];
assign t[35560] = t[35559] ^ n[35560];
assign t[35561] = t[35560] ^ n[35561];
assign t[35562] = t[35561] ^ n[35562];
assign t[35563] = t[35562] ^ n[35563];
assign t[35564] = t[35563] ^ n[35564];
assign t[35565] = t[35564] ^ n[35565];
assign t[35566] = t[35565] ^ n[35566];
assign t[35567] = t[35566] ^ n[35567];
assign t[35568] = t[35567] ^ n[35568];
assign t[35569] = t[35568] ^ n[35569];
assign t[35570] = t[35569] ^ n[35570];
assign t[35571] = t[35570] ^ n[35571];
assign t[35572] = t[35571] ^ n[35572];
assign t[35573] = t[35572] ^ n[35573];
assign t[35574] = t[35573] ^ n[35574];
assign t[35575] = t[35574] ^ n[35575];
assign t[35576] = t[35575] ^ n[35576];
assign t[35577] = t[35576] ^ n[35577];
assign t[35578] = t[35577] ^ n[35578];
assign t[35579] = t[35578] ^ n[35579];
assign t[35580] = t[35579] ^ n[35580];
assign t[35581] = t[35580] ^ n[35581];
assign t[35582] = t[35581] ^ n[35582];
assign t[35583] = t[35582] ^ n[35583];
assign t[35584] = t[35583] ^ n[35584];
assign t[35585] = t[35584] ^ n[35585];
assign t[35586] = t[35585] ^ n[35586];
assign t[35587] = t[35586] ^ n[35587];
assign t[35588] = t[35587] ^ n[35588];
assign t[35589] = t[35588] ^ n[35589];
assign t[35590] = t[35589] ^ n[35590];
assign t[35591] = t[35590] ^ n[35591];
assign t[35592] = t[35591] ^ n[35592];
assign t[35593] = t[35592] ^ n[35593];
assign t[35594] = t[35593] ^ n[35594];
assign t[35595] = t[35594] ^ n[35595];
assign t[35596] = t[35595] ^ n[35596];
assign t[35597] = t[35596] ^ n[35597];
assign t[35598] = t[35597] ^ n[35598];
assign t[35599] = t[35598] ^ n[35599];
assign t[35600] = t[35599] ^ n[35600];
assign t[35601] = t[35600] ^ n[35601];
assign t[35602] = t[35601] ^ n[35602];
assign t[35603] = t[35602] ^ n[35603];
assign t[35604] = t[35603] ^ n[35604];
assign t[35605] = t[35604] ^ n[35605];
assign t[35606] = t[35605] ^ n[35606];
assign t[35607] = t[35606] ^ n[35607];
assign t[35608] = t[35607] ^ n[35608];
assign t[35609] = t[35608] ^ n[35609];
assign t[35610] = t[35609] ^ n[35610];
assign t[35611] = t[35610] ^ n[35611];
assign t[35612] = t[35611] ^ n[35612];
assign t[35613] = t[35612] ^ n[35613];
assign t[35614] = t[35613] ^ n[35614];
assign t[35615] = t[35614] ^ n[35615];
assign t[35616] = t[35615] ^ n[35616];
assign t[35617] = t[35616] ^ n[35617];
assign t[35618] = t[35617] ^ n[35618];
assign t[35619] = t[35618] ^ n[35619];
assign t[35620] = t[35619] ^ n[35620];
assign t[35621] = t[35620] ^ n[35621];
assign t[35622] = t[35621] ^ n[35622];
assign t[35623] = t[35622] ^ n[35623];
assign t[35624] = t[35623] ^ n[35624];
assign t[35625] = t[35624] ^ n[35625];
assign t[35626] = t[35625] ^ n[35626];
assign t[35627] = t[35626] ^ n[35627];
assign t[35628] = t[35627] ^ n[35628];
assign t[35629] = t[35628] ^ n[35629];
assign t[35630] = t[35629] ^ n[35630];
assign t[35631] = t[35630] ^ n[35631];
assign t[35632] = t[35631] ^ n[35632];
assign t[35633] = t[35632] ^ n[35633];
assign t[35634] = t[35633] ^ n[35634];
assign t[35635] = t[35634] ^ n[35635];
assign t[35636] = t[35635] ^ n[35636];
assign t[35637] = t[35636] ^ n[35637];
assign t[35638] = t[35637] ^ n[35638];
assign t[35639] = t[35638] ^ n[35639];
assign t[35640] = t[35639] ^ n[35640];
assign t[35641] = t[35640] ^ n[35641];
assign t[35642] = t[35641] ^ n[35642];
assign t[35643] = t[35642] ^ n[35643];
assign t[35644] = t[35643] ^ n[35644];
assign t[35645] = t[35644] ^ n[35645];
assign t[35646] = t[35645] ^ n[35646];
assign t[35647] = t[35646] ^ n[35647];
assign t[35648] = t[35647] ^ n[35648];
assign t[35649] = t[35648] ^ n[35649];
assign t[35650] = t[35649] ^ n[35650];
assign t[35651] = t[35650] ^ n[35651];
assign t[35652] = t[35651] ^ n[35652];
assign t[35653] = t[35652] ^ n[35653];
assign t[35654] = t[35653] ^ n[35654];
assign t[35655] = t[35654] ^ n[35655];
assign t[35656] = t[35655] ^ n[35656];
assign t[35657] = t[35656] ^ n[35657];
assign t[35658] = t[35657] ^ n[35658];
assign t[35659] = t[35658] ^ n[35659];
assign t[35660] = t[35659] ^ n[35660];
assign t[35661] = t[35660] ^ n[35661];
assign t[35662] = t[35661] ^ n[35662];
assign t[35663] = t[35662] ^ n[35663];
assign t[35664] = t[35663] ^ n[35664];
assign t[35665] = t[35664] ^ n[35665];
assign t[35666] = t[35665] ^ n[35666];
assign t[35667] = t[35666] ^ n[35667];
assign t[35668] = t[35667] ^ n[35668];
assign t[35669] = t[35668] ^ n[35669];
assign t[35670] = t[35669] ^ n[35670];
assign t[35671] = t[35670] ^ n[35671];
assign t[35672] = t[35671] ^ n[35672];
assign t[35673] = t[35672] ^ n[35673];
assign t[35674] = t[35673] ^ n[35674];
assign t[35675] = t[35674] ^ n[35675];
assign t[35676] = t[35675] ^ n[35676];
assign t[35677] = t[35676] ^ n[35677];
assign t[35678] = t[35677] ^ n[35678];
assign t[35679] = t[35678] ^ n[35679];
assign t[35680] = t[35679] ^ n[35680];
assign t[35681] = t[35680] ^ n[35681];
assign t[35682] = t[35681] ^ n[35682];
assign t[35683] = t[35682] ^ n[35683];
assign t[35684] = t[35683] ^ n[35684];
assign t[35685] = t[35684] ^ n[35685];
assign t[35686] = t[35685] ^ n[35686];
assign t[35687] = t[35686] ^ n[35687];
assign t[35688] = t[35687] ^ n[35688];
assign t[35689] = t[35688] ^ n[35689];
assign t[35690] = t[35689] ^ n[35690];
assign t[35691] = t[35690] ^ n[35691];
assign t[35692] = t[35691] ^ n[35692];
assign t[35693] = t[35692] ^ n[35693];
assign t[35694] = t[35693] ^ n[35694];
assign t[35695] = t[35694] ^ n[35695];
assign t[35696] = t[35695] ^ n[35696];
assign t[35697] = t[35696] ^ n[35697];
assign t[35698] = t[35697] ^ n[35698];
assign t[35699] = t[35698] ^ n[35699];
assign t[35700] = t[35699] ^ n[35700];
assign t[35701] = t[35700] ^ n[35701];
assign t[35702] = t[35701] ^ n[35702];
assign t[35703] = t[35702] ^ n[35703];
assign t[35704] = t[35703] ^ n[35704];
assign t[35705] = t[35704] ^ n[35705];
assign t[35706] = t[35705] ^ n[35706];
assign t[35707] = t[35706] ^ n[35707];
assign t[35708] = t[35707] ^ n[35708];
assign t[35709] = t[35708] ^ n[35709];
assign t[35710] = t[35709] ^ n[35710];
assign t[35711] = t[35710] ^ n[35711];
assign t[35712] = t[35711] ^ n[35712];
assign t[35713] = t[35712] ^ n[35713];
assign t[35714] = t[35713] ^ n[35714];
assign t[35715] = t[35714] ^ n[35715];
assign t[35716] = t[35715] ^ n[35716];
assign t[35717] = t[35716] ^ n[35717];
assign t[35718] = t[35717] ^ n[35718];
assign t[35719] = t[35718] ^ n[35719];
assign t[35720] = t[35719] ^ n[35720];
assign t[35721] = t[35720] ^ n[35721];
assign t[35722] = t[35721] ^ n[35722];
assign t[35723] = t[35722] ^ n[35723];
assign t[35724] = t[35723] ^ n[35724];
assign t[35725] = t[35724] ^ n[35725];
assign t[35726] = t[35725] ^ n[35726];
assign t[35727] = t[35726] ^ n[35727];
assign t[35728] = t[35727] ^ n[35728];
assign t[35729] = t[35728] ^ n[35729];
assign t[35730] = t[35729] ^ n[35730];
assign t[35731] = t[35730] ^ n[35731];
assign t[35732] = t[35731] ^ n[35732];
assign t[35733] = t[35732] ^ n[35733];
assign t[35734] = t[35733] ^ n[35734];
assign t[35735] = t[35734] ^ n[35735];
assign t[35736] = t[35735] ^ n[35736];
assign t[35737] = t[35736] ^ n[35737];
assign t[35738] = t[35737] ^ n[35738];
assign t[35739] = t[35738] ^ n[35739];
assign t[35740] = t[35739] ^ n[35740];
assign t[35741] = t[35740] ^ n[35741];
assign t[35742] = t[35741] ^ n[35742];
assign t[35743] = t[35742] ^ n[35743];
assign t[35744] = t[35743] ^ n[35744];
assign t[35745] = t[35744] ^ n[35745];
assign t[35746] = t[35745] ^ n[35746];
assign t[35747] = t[35746] ^ n[35747];
assign t[35748] = t[35747] ^ n[35748];
assign t[35749] = t[35748] ^ n[35749];
assign t[35750] = t[35749] ^ n[35750];
assign t[35751] = t[35750] ^ n[35751];
assign t[35752] = t[35751] ^ n[35752];
assign t[35753] = t[35752] ^ n[35753];
assign t[35754] = t[35753] ^ n[35754];
assign t[35755] = t[35754] ^ n[35755];
assign t[35756] = t[35755] ^ n[35756];
assign t[35757] = t[35756] ^ n[35757];
assign t[35758] = t[35757] ^ n[35758];
assign t[35759] = t[35758] ^ n[35759];
assign t[35760] = t[35759] ^ n[35760];
assign t[35761] = t[35760] ^ n[35761];
assign t[35762] = t[35761] ^ n[35762];
assign t[35763] = t[35762] ^ n[35763];
assign t[35764] = t[35763] ^ n[35764];
assign t[35765] = t[35764] ^ n[35765];
assign t[35766] = t[35765] ^ n[35766];
assign t[35767] = t[35766] ^ n[35767];
assign t[35768] = t[35767] ^ n[35768];
assign t[35769] = t[35768] ^ n[35769];
assign t[35770] = t[35769] ^ n[35770];
assign t[35771] = t[35770] ^ n[35771];
assign t[35772] = t[35771] ^ n[35772];
assign t[35773] = t[35772] ^ n[35773];
assign t[35774] = t[35773] ^ n[35774];
assign t[35775] = t[35774] ^ n[35775];
assign t[35776] = t[35775] ^ n[35776];
assign t[35777] = t[35776] ^ n[35777];
assign t[35778] = t[35777] ^ n[35778];
assign t[35779] = t[35778] ^ n[35779];
assign t[35780] = t[35779] ^ n[35780];
assign t[35781] = t[35780] ^ n[35781];
assign t[35782] = t[35781] ^ n[35782];
assign t[35783] = t[35782] ^ n[35783];
assign t[35784] = t[35783] ^ n[35784];
assign t[35785] = t[35784] ^ n[35785];
assign t[35786] = t[35785] ^ n[35786];
assign t[35787] = t[35786] ^ n[35787];
assign t[35788] = t[35787] ^ n[35788];
assign t[35789] = t[35788] ^ n[35789];
assign t[35790] = t[35789] ^ n[35790];
assign t[35791] = t[35790] ^ n[35791];
assign t[35792] = t[35791] ^ n[35792];
assign t[35793] = t[35792] ^ n[35793];
assign t[35794] = t[35793] ^ n[35794];
assign t[35795] = t[35794] ^ n[35795];
assign t[35796] = t[35795] ^ n[35796];
assign t[35797] = t[35796] ^ n[35797];
assign t[35798] = t[35797] ^ n[35798];
assign t[35799] = t[35798] ^ n[35799];
assign t[35800] = t[35799] ^ n[35800];
assign t[35801] = t[35800] ^ n[35801];
assign t[35802] = t[35801] ^ n[35802];
assign t[35803] = t[35802] ^ n[35803];
assign t[35804] = t[35803] ^ n[35804];
assign t[35805] = t[35804] ^ n[35805];
assign t[35806] = t[35805] ^ n[35806];
assign t[35807] = t[35806] ^ n[35807];
assign t[35808] = t[35807] ^ n[35808];
assign t[35809] = t[35808] ^ n[35809];
assign t[35810] = t[35809] ^ n[35810];
assign t[35811] = t[35810] ^ n[35811];
assign t[35812] = t[35811] ^ n[35812];
assign t[35813] = t[35812] ^ n[35813];
assign t[35814] = t[35813] ^ n[35814];
assign t[35815] = t[35814] ^ n[35815];
assign t[35816] = t[35815] ^ n[35816];
assign t[35817] = t[35816] ^ n[35817];
assign t[35818] = t[35817] ^ n[35818];
assign t[35819] = t[35818] ^ n[35819];
assign t[35820] = t[35819] ^ n[35820];
assign t[35821] = t[35820] ^ n[35821];
assign t[35822] = t[35821] ^ n[35822];
assign t[35823] = t[35822] ^ n[35823];
assign t[35824] = t[35823] ^ n[35824];
assign t[35825] = t[35824] ^ n[35825];
assign t[35826] = t[35825] ^ n[35826];
assign t[35827] = t[35826] ^ n[35827];
assign t[35828] = t[35827] ^ n[35828];
assign t[35829] = t[35828] ^ n[35829];
assign t[35830] = t[35829] ^ n[35830];
assign t[35831] = t[35830] ^ n[35831];
assign t[35832] = t[35831] ^ n[35832];
assign t[35833] = t[35832] ^ n[35833];
assign t[35834] = t[35833] ^ n[35834];
assign t[35835] = t[35834] ^ n[35835];
assign t[35836] = t[35835] ^ n[35836];
assign t[35837] = t[35836] ^ n[35837];
assign t[35838] = t[35837] ^ n[35838];
assign t[35839] = t[35838] ^ n[35839];
assign t[35840] = t[35839] ^ n[35840];
assign t[35841] = t[35840] ^ n[35841];
assign t[35842] = t[35841] ^ n[35842];
assign t[35843] = t[35842] ^ n[35843];
assign t[35844] = t[35843] ^ n[35844];
assign t[35845] = t[35844] ^ n[35845];
assign t[35846] = t[35845] ^ n[35846];
assign t[35847] = t[35846] ^ n[35847];
assign t[35848] = t[35847] ^ n[35848];
assign t[35849] = t[35848] ^ n[35849];
assign t[35850] = t[35849] ^ n[35850];
assign t[35851] = t[35850] ^ n[35851];
assign t[35852] = t[35851] ^ n[35852];
assign t[35853] = t[35852] ^ n[35853];
assign t[35854] = t[35853] ^ n[35854];
assign t[35855] = t[35854] ^ n[35855];
assign t[35856] = t[35855] ^ n[35856];
assign t[35857] = t[35856] ^ n[35857];
assign t[35858] = t[35857] ^ n[35858];
assign t[35859] = t[35858] ^ n[35859];
assign t[35860] = t[35859] ^ n[35860];
assign t[35861] = t[35860] ^ n[35861];
assign t[35862] = t[35861] ^ n[35862];
assign t[35863] = t[35862] ^ n[35863];
assign t[35864] = t[35863] ^ n[35864];
assign t[35865] = t[35864] ^ n[35865];
assign t[35866] = t[35865] ^ n[35866];
assign t[35867] = t[35866] ^ n[35867];
assign t[35868] = t[35867] ^ n[35868];
assign t[35869] = t[35868] ^ n[35869];
assign t[35870] = t[35869] ^ n[35870];
assign t[35871] = t[35870] ^ n[35871];
assign t[35872] = t[35871] ^ n[35872];
assign t[35873] = t[35872] ^ n[35873];
assign t[35874] = t[35873] ^ n[35874];
assign t[35875] = t[35874] ^ n[35875];
assign t[35876] = t[35875] ^ n[35876];
assign t[35877] = t[35876] ^ n[35877];
assign t[35878] = t[35877] ^ n[35878];
assign t[35879] = t[35878] ^ n[35879];
assign t[35880] = t[35879] ^ n[35880];
assign t[35881] = t[35880] ^ n[35881];
assign t[35882] = t[35881] ^ n[35882];
assign t[35883] = t[35882] ^ n[35883];
assign t[35884] = t[35883] ^ n[35884];
assign t[35885] = t[35884] ^ n[35885];
assign t[35886] = t[35885] ^ n[35886];
assign t[35887] = t[35886] ^ n[35887];
assign t[35888] = t[35887] ^ n[35888];
assign t[35889] = t[35888] ^ n[35889];
assign t[35890] = t[35889] ^ n[35890];
assign t[35891] = t[35890] ^ n[35891];
assign t[35892] = t[35891] ^ n[35892];
assign t[35893] = t[35892] ^ n[35893];
assign t[35894] = t[35893] ^ n[35894];
assign t[35895] = t[35894] ^ n[35895];
assign t[35896] = t[35895] ^ n[35896];
assign t[35897] = t[35896] ^ n[35897];
assign t[35898] = t[35897] ^ n[35898];
assign t[35899] = t[35898] ^ n[35899];
assign t[35900] = t[35899] ^ n[35900];
assign t[35901] = t[35900] ^ n[35901];
assign t[35902] = t[35901] ^ n[35902];
assign t[35903] = t[35902] ^ n[35903];
assign t[35904] = t[35903] ^ n[35904];
assign t[35905] = t[35904] ^ n[35905];
assign t[35906] = t[35905] ^ n[35906];
assign t[35907] = t[35906] ^ n[35907];
assign t[35908] = t[35907] ^ n[35908];
assign t[35909] = t[35908] ^ n[35909];
assign t[35910] = t[35909] ^ n[35910];
assign t[35911] = t[35910] ^ n[35911];
assign t[35912] = t[35911] ^ n[35912];
assign t[35913] = t[35912] ^ n[35913];
assign t[35914] = t[35913] ^ n[35914];
assign t[35915] = t[35914] ^ n[35915];
assign t[35916] = t[35915] ^ n[35916];
assign t[35917] = t[35916] ^ n[35917];
assign t[35918] = t[35917] ^ n[35918];
assign t[35919] = t[35918] ^ n[35919];
assign t[35920] = t[35919] ^ n[35920];
assign t[35921] = t[35920] ^ n[35921];
assign t[35922] = t[35921] ^ n[35922];
assign t[35923] = t[35922] ^ n[35923];
assign t[35924] = t[35923] ^ n[35924];
assign t[35925] = t[35924] ^ n[35925];
assign t[35926] = t[35925] ^ n[35926];
assign t[35927] = t[35926] ^ n[35927];
assign t[35928] = t[35927] ^ n[35928];
assign t[35929] = t[35928] ^ n[35929];
assign t[35930] = t[35929] ^ n[35930];
assign t[35931] = t[35930] ^ n[35931];
assign t[35932] = t[35931] ^ n[35932];
assign t[35933] = t[35932] ^ n[35933];
assign t[35934] = t[35933] ^ n[35934];
assign t[35935] = t[35934] ^ n[35935];
assign t[35936] = t[35935] ^ n[35936];
assign t[35937] = t[35936] ^ n[35937];
assign t[35938] = t[35937] ^ n[35938];
assign t[35939] = t[35938] ^ n[35939];
assign t[35940] = t[35939] ^ n[35940];
assign t[35941] = t[35940] ^ n[35941];
assign t[35942] = t[35941] ^ n[35942];
assign t[35943] = t[35942] ^ n[35943];
assign t[35944] = t[35943] ^ n[35944];
assign t[35945] = t[35944] ^ n[35945];
assign t[35946] = t[35945] ^ n[35946];
assign t[35947] = t[35946] ^ n[35947];
assign t[35948] = t[35947] ^ n[35948];
assign t[35949] = t[35948] ^ n[35949];
assign t[35950] = t[35949] ^ n[35950];
assign t[35951] = t[35950] ^ n[35951];
assign t[35952] = t[35951] ^ n[35952];
assign t[35953] = t[35952] ^ n[35953];
assign t[35954] = t[35953] ^ n[35954];
assign t[35955] = t[35954] ^ n[35955];
assign t[35956] = t[35955] ^ n[35956];
assign t[35957] = t[35956] ^ n[35957];
assign t[35958] = t[35957] ^ n[35958];
assign t[35959] = t[35958] ^ n[35959];
assign t[35960] = t[35959] ^ n[35960];
assign t[35961] = t[35960] ^ n[35961];
assign t[35962] = t[35961] ^ n[35962];
assign t[35963] = t[35962] ^ n[35963];
assign t[35964] = t[35963] ^ n[35964];
assign t[35965] = t[35964] ^ n[35965];
assign t[35966] = t[35965] ^ n[35966];
assign t[35967] = t[35966] ^ n[35967];
assign t[35968] = t[35967] ^ n[35968];
assign t[35969] = t[35968] ^ n[35969];
assign t[35970] = t[35969] ^ n[35970];
assign t[35971] = t[35970] ^ n[35971];
assign t[35972] = t[35971] ^ n[35972];
assign t[35973] = t[35972] ^ n[35973];
assign t[35974] = t[35973] ^ n[35974];
assign t[35975] = t[35974] ^ n[35975];
assign t[35976] = t[35975] ^ n[35976];
assign t[35977] = t[35976] ^ n[35977];
assign t[35978] = t[35977] ^ n[35978];
assign t[35979] = t[35978] ^ n[35979];
assign t[35980] = t[35979] ^ n[35980];
assign t[35981] = t[35980] ^ n[35981];
assign t[35982] = t[35981] ^ n[35982];
assign t[35983] = t[35982] ^ n[35983];
assign t[35984] = t[35983] ^ n[35984];
assign t[35985] = t[35984] ^ n[35985];
assign t[35986] = t[35985] ^ n[35986];
assign t[35987] = t[35986] ^ n[35987];
assign t[35988] = t[35987] ^ n[35988];
assign t[35989] = t[35988] ^ n[35989];
assign t[35990] = t[35989] ^ n[35990];
assign t[35991] = t[35990] ^ n[35991];
assign t[35992] = t[35991] ^ n[35992];
assign t[35993] = t[35992] ^ n[35993];
assign t[35994] = t[35993] ^ n[35994];
assign t[35995] = t[35994] ^ n[35995];
assign t[35996] = t[35995] ^ n[35996];
assign t[35997] = t[35996] ^ n[35997];
assign t[35998] = t[35997] ^ n[35998];
assign t[35999] = t[35998] ^ n[35999];
assign t[36000] = t[35999] ^ n[36000];
assign t[36001] = t[36000] ^ n[36001];
assign t[36002] = t[36001] ^ n[36002];
assign t[36003] = t[36002] ^ n[36003];
assign t[36004] = t[36003] ^ n[36004];
assign t[36005] = t[36004] ^ n[36005];
assign t[36006] = t[36005] ^ n[36006];
assign t[36007] = t[36006] ^ n[36007];
assign t[36008] = t[36007] ^ n[36008];
assign t[36009] = t[36008] ^ n[36009];
assign t[36010] = t[36009] ^ n[36010];
assign t[36011] = t[36010] ^ n[36011];
assign t[36012] = t[36011] ^ n[36012];
assign t[36013] = t[36012] ^ n[36013];
assign t[36014] = t[36013] ^ n[36014];
assign t[36015] = t[36014] ^ n[36015];
assign t[36016] = t[36015] ^ n[36016];
assign t[36017] = t[36016] ^ n[36017];
assign t[36018] = t[36017] ^ n[36018];
assign t[36019] = t[36018] ^ n[36019];
assign t[36020] = t[36019] ^ n[36020];
assign t[36021] = t[36020] ^ n[36021];
assign t[36022] = t[36021] ^ n[36022];
assign t[36023] = t[36022] ^ n[36023];
assign t[36024] = t[36023] ^ n[36024];
assign t[36025] = t[36024] ^ n[36025];
assign t[36026] = t[36025] ^ n[36026];
assign t[36027] = t[36026] ^ n[36027];
assign t[36028] = t[36027] ^ n[36028];
assign t[36029] = t[36028] ^ n[36029];
assign t[36030] = t[36029] ^ n[36030];
assign t[36031] = t[36030] ^ n[36031];
assign t[36032] = t[36031] ^ n[36032];
assign t[36033] = t[36032] ^ n[36033];
assign t[36034] = t[36033] ^ n[36034];
assign t[36035] = t[36034] ^ n[36035];
assign t[36036] = t[36035] ^ n[36036];
assign t[36037] = t[36036] ^ n[36037];
assign t[36038] = t[36037] ^ n[36038];
assign t[36039] = t[36038] ^ n[36039];
assign t[36040] = t[36039] ^ n[36040];
assign t[36041] = t[36040] ^ n[36041];
assign t[36042] = t[36041] ^ n[36042];
assign t[36043] = t[36042] ^ n[36043];
assign t[36044] = t[36043] ^ n[36044];
assign t[36045] = t[36044] ^ n[36045];
assign t[36046] = t[36045] ^ n[36046];
assign t[36047] = t[36046] ^ n[36047];
assign t[36048] = t[36047] ^ n[36048];
assign t[36049] = t[36048] ^ n[36049];
assign t[36050] = t[36049] ^ n[36050];
assign t[36051] = t[36050] ^ n[36051];
assign t[36052] = t[36051] ^ n[36052];
assign t[36053] = t[36052] ^ n[36053];
assign t[36054] = t[36053] ^ n[36054];
assign t[36055] = t[36054] ^ n[36055];
assign t[36056] = t[36055] ^ n[36056];
assign t[36057] = t[36056] ^ n[36057];
assign t[36058] = t[36057] ^ n[36058];
assign t[36059] = t[36058] ^ n[36059];
assign t[36060] = t[36059] ^ n[36060];
assign t[36061] = t[36060] ^ n[36061];
assign t[36062] = t[36061] ^ n[36062];
assign t[36063] = t[36062] ^ n[36063];
assign t[36064] = t[36063] ^ n[36064];
assign t[36065] = t[36064] ^ n[36065];
assign t[36066] = t[36065] ^ n[36066];
assign t[36067] = t[36066] ^ n[36067];
assign t[36068] = t[36067] ^ n[36068];
assign t[36069] = t[36068] ^ n[36069];
assign t[36070] = t[36069] ^ n[36070];
assign t[36071] = t[36070] ^ n[36071];
assign t[36072] = t[36071] ^ n[36072];
assign t[36073] = t[36072] ^ n[36073];
assign t[36074] = t[36073] ^ n[36074];
assign t[36075] = t[36074] ^ n[36075];
assign t[36076] = t[36075] ^ n[36076];
assign t[36077] = t[36076] ^ n[36077];
assign t[36078] = t[36077] ^ n[36078];
assign t[36079] = t[36078] ^ n[36079];
assign t[36080] = t[36079] ^ n[36080];
assign t[36081] = t[36080] ^ n[36081];
assign t[36082] = t[36081] ^ n[36082];
assign t[36083] = t[36082] ^ n[36083];
assign t[36084] = t[36083] ^ n[36084];
assign t[36085] = t[36084] ^ n[36085];
assign t[36086] = t[36085] ^ n[36086];
assign t[36087] = t[36086] ^ n[36087];
assign t[36088] = t[36087] ^ n[36088];
assign t[36089] = t[36088] ^ n[36089];
assign t[36090] = t[36089] ^ n[36090];
assign t[36091] = t[36090] ^ n[36091];
assign t[36092] = t[36091] ^ n[36092];
assign t[36093] = t[36092] ^ n[36093];
assign t[36094] = t[36093] ^ n[36094];
assign t[36095] = t[36094] ^ n[36095];
assign t[36096] = t[36095] ^ n[36096];
assign t[36097] = t[36096] ^ n[36097];
assign t[36098] = t[36097] ^ n[36098];
assign t[36099] = t[36098] ^ n[36099];
assign t[36100] = t[36099] ^ n[36100];
assign t[36101] = t[36100] ^ n[36101];
assign t[36102] = t[36101] ^ n[36102];
assign t[36103] = t[36102] ^ n[36103];
assign t[36104] = t[36103] ^ n[36104];
assign t[36105] = t[36104] ^ n[36105];
assign t[36106] = t[36105] ^ n[36106];
assign t[36107] = t[36106] ^ n[36107];
assign t[36108] = t[36107] ^ n[36108];
assign t[36109] = t[36108] ^ n[36109];
assign t[36110] = t[36109] ^ n[36110];
assign t[36111] = t[36110] ^ n[36111];
assign t[36112] = t[36111] ^ n[36112];
assign t[36113] = t[36112] ^ n[36113];
assign t[36114] = t[36113] ^ n[36114];
assign t[36115] = t[36114] ^ n[36115];
assign t[36116] = t[36115] ^ n[36116];
assign t[36117] = t[36116] ^ n[36117];
assign t[36118] = t[36117] ^ n[36118];
assign t[36119] = t[36118] ^ n[36119];
assign t[36120] = t[36119] ^ n[36120];
assign t[36121] = t[36120] ^ n[36121];
assign t[36122] = t[36121] ^ n[36122];
assign t[36123] = t[36122] ^ n[36123];
assign t[36124] = t[36123] ^ n[36124];
assign t[36125] = t[36124] ^ n[36125];
assign t[36126] = t[36125] ^ n[36126];
assign t[36127] = t[36126] ^ n[36127];
assign t[36128] = t[36127] ^ n[36128];
assign t[36129] = t[36128] ^ n[36129];
assign t[36130] = t[36129] ^ n[36130];
assign t[36131] = t[36130] ^ n[36131];
assign t[36132] = t[36131] ^ n[36132];
assign t[36133] = t[36132] ^ n[36133];
assign t[36134] = t[36133] ^ n[36134];
assign t[36135] = t[36134] ^ n[36135];
assign t[36136] = t[36135] ^ n[36136];
assign t[36137] = t[36136] ^ n[36137];
assign t[36138] = t[36137] ^ n[36138];
assign t[36139] = t[36138] ^ n[36139];
assign t[36140] = t[36139] ^ n[36140];
assign t[36141] = t[36140] ^ n[36141];
assign t[36142] = t[36141] ^ n[36142];
assign t[36143] = t[36142] ^ n[36143];
assign t[36144] = t[36143] ^ n[36144];
assign t[36145] = t[36144] ^ n[36145];
assign t[36146] = t[36145] ^ n[36146];
assign t[36147] = t[36146] ^ n[36147];
assign t[36148] = t[36147] ^ n[36148];
assign t[36149] = t[36148] ^ n[36149];
assign t[36150] = t[36149] ^ n[36150];
assign t[36151] = t[36150] ^ n[36151];
assign t[36152] = t[36151] ^ n[36152];
assign t[36153] = t[36152] ^ n[36153];
assign t[36154] = t[36153] ^ n[36154];
assign t[36155] = t[36154] ^ n[36155];
assign t[36156] = t[36155] ^ n[36156];
assign t[36157] = t[36156] ^ n[36157];
assign t[36158] = t[36157] ^ n[36158];
assign t[36159] = t[36158] ^ n[36159];
assign t[36160] = t[36159] ^ n[36160];
assign t[36161] = t[36160] ^ n[36161];
assign t[36162] = t[36161] ^ n[36162];
assign t[36163] = t[36162] ^ n[36163];
assign t[36164] = t[36163] ^ n[36164];
assign t[36165] = t[36164] ^ n[36165];
assign t[36166] = t[36165] ^ n[36166];
assign t[36167] = t[36166] ^ n[36167];
assign t[36168] = t[36167] ^ n[36168];
assign t[36169] = t[36168] ^ n[36169];
assign t[36170] = t[36169] ^ n[36170];
assign t[36171] = t[36170] ^ n[36171];
assign t[36172] = t[36171] ^ n[36172];
assign t[36173] = t[36172] ^ n[36173];
assign t[36174] = t[36173] ^ n[36174];
assign t[36175] = t[36174] ^ n[36175];
assign t[36176] = t[36175] ^ n[36176];
assign t[36177] = t[36176] ^ n[36177];
assign t[36178] = t[36177] ^ n[36178];
assign t[36179] = t[36178] ^ n[36179];
assign t[36180] = t[36179] ^ n[36180];
assign t[36181] = t[36180] ^ n[36181];
assign t[36182] = t[36181] ^ n[36182];
assign t[36183] = t[36182] ^ n[36183];
assign t[36184] = t[36183] ^ n[36184];
assign t[36185] = t[36184] ^ n[36185];
assign t[36186] = t[36185] ^ n[36186];
assign t[36187] = t[36186] ^ n[36187];
assign t[36188] = t[36187] ^ n[36188];
assign t[36189] = t[36188] ^ n[36189];
assign t[36190] = t[36189] ^ n[36190];
assign t[36191] = t[36190] ^ n[36191];
assign t[36192] = t[36191] ^ n[36192];
assign t[36193] = t[36192] ^ n[36193];
assign t[36194] = t[36193] ^ n[36194];
assign t[36195] = t[36194] ^ n[36195];
assign t[36196] = t[36195] ^ n[36196];
assign t[36197] = t[36196] ^ n[36197];
assign t[36198] = t[36197] ^ n[36198];
assign t[36199] = t[36198] ^ n[36199];
assign t[36200] = t[36199] ^ n[36200];
assign t[36201] = t[36200] ^ n[36201];
assign t[36202] = t[36201] ^ n[36202];
assign t[36203] = t[36202] ^ n[36203];
assign t[36204] = t[36203] ^ n[36204];
assign t[36205] = t[36204] ^ n[36205];
assign t[36206] = t[36205] ^ n[36206];
assign t[36207] = t[36206] ^ n[36207];
assign t[36208] = t[36207] ^ n[36208];
assign t[36209] = t[36208] ^ n[36209];
assign t[36210] = t[36209] ^ n[36210];
assign t[36211] = t[36210] ^ n[36211];
assign t[36212] = t[36211] ^ n[36212];
assign t[36213] = t[36212] ^ n[36213];
assign t[36214] = t[36213] ^ n[36214];
assign t[36215] = t[36214] ^ n[36215];
assign t[36216] = t[36215] ^ n[36216];
assign t[36217] = t[36216] ^ n[36217];
assign t[36218] = t[36217] ^ n[36218];
assign t[36219] = t[36218] ^ n[36219];
assign t[36220] = t[36219] ^ n[36220];
assign t[36221] = t[36220] ^ n[36221];
assign t[36222] = t[36221] ^ n[36222];
assign t[36223] = t[36222] ^ n[36223];
assign t[36224] = t[36223] ^ n[36224];
assign t[36225] = t[36224] ^ n[36225];
assign t[36226] = t[36225] ^ n[36226];
assign t[36227] = t[36226] ^ n[36227];
assign t[36228] = t[36227] ^ n[36228];
assign t[36229] = t[36228] ^ n[36229];
assign t[36230] = t[36229] ^ n[36230];
assign t[36231] = t[36230] ^ n[36231];
assign t[36232] = t[36231] ^ n[36232];
assign t[36233] = t[36232] ^ n[36233];
assign t[36234] = t[36233] ^ n[36234];
assign t[36235] = t[36234] ^ n[36235];
assign t[36236] = t[36235] ^ n[36236];
assign t[36237] = t[36236] ^ n[36237];
assign t[36238] = t[36237] ^ n[36238];
assign t[36239] = t[36238] ^ n[36239];
assign t[36240] = t[36239] ^ n[36240];
assign t[36241] = t[36240] ^ n[36241];
assign t[36242] = t[36241] ^ n[36242];
assign t[36243] = t[36242] ^ n[36243];
assign t[36244] = t[36243] ^ n[36244];
assign t[36245] = t[36244] ^ n[36245];
assign t[36246] = t[36245] ^ n[36246];
assign t[36247] = t[36246] ^ n[36247];
assign t[36248] = t[36247] ^ n[36248];
assign t[36249] = t[36248] ^ n[36249];
assign t[36250] = t[36249] ^ n[36250];
assign t[36251] = t[36250] ^ n[36251];
assign t[36252] = t[36251] ^ n[36252];
assign t[36253] = t[36252] ^ n[36253];
assign t[36254] = t[36253] ^ n[36254];
assign t[36255] = t[36254] ^ n[36255];
assign t[36256] = t[36255] ^ n[36256];
assign t[36257] = t[36256] ^ n[36257];
assign t[36258] = t[36257] ^ n[36258];
assign t[36259] = t[36258] ^ n[36259];
assign t[36260] = t[36259] ^ n[36260];
assign t[36261] = t[36260] ^ n[36261];
assign t[36262] = t[36261] ^ n[36262];
assign t[36263] = t[36262] ^ n[36263];
assign t[36264] = t[36263] ^ n[36264];
assign t[36265] = t[36264] ^ n[36265];
assign t[36266] = t[36265] ^ n[36266];
assign t[36267] = t[36266] ^ n[36267];
assign t[36268] = t[36267] ^ n[36268];
assign t[36269] = t[36268] ^ n[36269];
assign t[36270] = t[36269] ^ n[36270];
assign t[36271] = t[36270] ^ n[36271];
assign t[36272] = t[36271] ^ n[36272];
assign t[36273] = t[36272] ^ n[36273];
assign t[36274] = t[36273] ^ n[36274];
assign t[36275] = t[36274] ^ n[36275];
assign t[36276] = t[36275] ^ n[36276];
assign t[36277] = t[36276] ^ n[36277];
assign t[36278] = t[36277] ^ n[36278];
assign t[36279] = t[36278] ^ n[36279];
assign t[36280] = t[36279] ^ n[36280];
assign t[36281] = t[36280] ^ n[36281];
assign t[36282] = t[36281] ^ n[36282];
assign t[36283] = t[36282] ^ n[36283];
assign t[36284] = t[36283] ^ n[36284];
assign t[36285] = t[36284] ^ n[36285];
assign t[36286] = t[36285] ^ n[36286];
assign t[36287] = t[36286] ^ n[36287];
assign t[36288] = t[36287] ^ n[36288];
assign t[36289] = t[36288] ^ n[36289];
assign t[36290] = t[36289] ^ n[36290];
assign t[36291] = t[36290] ^ n[36291];
assign t[36292] = t[36291] ^ n[36292];
assign t[36293] = t[36292] ^ n[36293];
assign t[36294] = t[36293] ^ n[36294];
assign t[36295] = t[36294] ^ n[36295];
assign t[36296] = t[36295] ^ n[36296];
assign t[36297] = t[36296] ^ n[36297];
assign t[36298] = t[36297] ^ n[36298];
assign t[36299] = t[36298] ^ n[36299];
assign t[36300] = t[36299] ^ n[36300];
assign t[36301] = t[36300] ^ n[36301];
assign t[36302] = t[36301] ^ n[36302];
assign t[36303] = t[36302] ^ n[36303];
assign t[36304] = t[36303] ^ n[36304];
assign t[36305] = t[36304] ^ n[36305];
assign t[36306] = t[36305] ^ n[36306];
assign t[36307] = t[36306] ^ n[36307];
assign t[36308] = t[36307] ^ n[36308];
assign t[36309] = t[36308] ^ n[36309];
assign t[36310] = t[36309] ^ n[36310];
assign t[36311] = t[36310] ^ n[36311];
assign t[36312] = t[36311] ^ n[36312];
assign t[36313] = t[36312] ^ n[36313];
assign t[36314] = t[36313] ^ n[36314];
assign t[36315] = t[36314] ^ n[36315];
assign t[36316] = t[36315] ^ n[36316];
assign t[36317] = t[36316] ^ n[36317];
assign t[36318] = t[36317] ^ n[36318];
assign t[36319] = t[36318] ^ n[36319];
assign t[36320] = t[36319] ^ n[36320];
assign t[36321] = t[36320] ^ n[36321];
assign t[36322] = t[36321] ^ n[36322];
assign t[36323] = t[36322] ^ n[36323];
assign t[36324] = t[36323] ^ n[36324];
assign t[36325] = t[36324] ^ n[36325];
assign t[36326] = t[36325] ^ n[36326];
assign t[36327] = t[36326] ^ n[36327];
assign t[36328] = t[36327] ^ n[36328];
assign t[36329] = t[36328] ^ n[36329];
assign t[36330] = t[36329] ^ n[36330];
assign t[36331] = t[36330] ^ n[36331];
assign t[36332] = t[36331] ^ n[36332];
assign t[36333] = t[36332] ^ n[36333];
assign t[36334] = t[36333] ^ n[36334];
assign t[36335] = t[36334] ^ n[36335];
assign t[36336] = t[36335] ^ n[36336];
assign t[36337] = t[36336] ^ n[36337];
assign t[36338] = t[36337] ^ n[36338];
assign t[36339] = t[36338] ^ n[36339];
assign t[36340] = t[36339] ^ n[36340];
assign t[36341] = t[36340] ^ n[36341];
assign t[36342] = t[36341] ^ n[36342];
assign t[36343] = t[36342] ^ n[36343];
assign t[36344] = t[36343] ^ n[36344];
assign t[36345] = t[36344] ^ n[36345];
assign t[36346] = t[36345] ^ n[36346];
assign t[36347] = t[36346] ^ n[36347];
assign t[36348] = t[36347] ^ n[36348];
assign t[36349] = t[36348] ^ n[36349];
assign t[36350] = t[36349] ^ n[36350];
assign t[36351] = t[36350] ^ n[36351];
assign t[36352] = t[36351] ^ n[36352];
assign t[36353] = t[36352] ^ n[36353];
assign t[36354] = t[36353] ^ n[36354];
assign t[36355] = t[36354] ^ n[36355];
assign t[36356] = t[36355] ^ n[36356];
assign t[36357] = t[36356] ^ n[36357];
assign t[36358] = t[36357] ^ n[36358];
assign t[36359] = t[36358] ^ n[36359];
assign t[36360] = t[36359] ^ n[36360];
assign t[36361] = t[36360] ^ n[36361];
assign t[36362] = t[36361] ^ n[36362];
assign t[36363] = t[36362] ^ n[36363];
assign t[36364] = t[36363] ^ n[36364];
assign t[36365] = t[36364] ^ n[36365];
assign t[36366] = t[36365] ^ n[36366];
assign t[36367] = t[36366] ^ n[36367];
assign t[36368] = t[36367] ^ n[36368];
assign t[36369] = t[36368] ^ n[36369];
assign t[36370] = t[36369] ^ n[36370];
assign t[36371] = t[36370] ^ n[36371];
assign t[36372] = t[36371] ^ n[36372];
assign t[36373] = t[36372] ^ n[36373];
assign t[36374] = t[36373] ^ n[36374];
assign t[36375] = t[36374] ^ n[36375];
assign t[36376] = t[36375] ^ n[36376];
assign t[36377] = t[36376] ^ n[36377];
assign t[36378] = t[36377] ^ n[36378];
assign t[36379] = t[36378] ^ n[36379];
assign t[36380] = t[36379] ^ n[36380];
assign t[36381] = t[36380] ^ n[36381];
assign t[36382] = t[36381] ^ n[36382];
assign t[36383] = t[36382] ^ n[36383];
assign t[36384] = t[36383] ^ n[36384];
assign t[36385] = t[36384] ^ n[36385];
assign t[36386] = t[36385] ^ n[36386];
assign t[36387] = t[36386] ^ n[36387];
assign t[36388] = t[36387] ^ n[36388];
assign t[36389] = t[36388] ^ n[36389];
assign t[36390] = t[36389] ^ n[36390];
assign t[36391] = t[36390] ^ n[36391];
assign t[36392] = t[36391] ^ n[36392];
assign t[36393] = t[36392] ^ n[36393];
assign t[36394] = t[36393] ^ n[36394];
assign t[36395] = t[36394] ^ n[36395];
assign t[36396] = t[36395] ^ n[36396];
assign t[36397] = t[36396] ^ n[36397];
assign t[36398] = t[36397] ^ n[36398];
assign t[36399] = t[36398] ^ n[36399];
assign t[36400] = t[36399] ^ n[36400];
assign t[36401] = t[36400] ^ n[36401];
assign t[36402] = t[36401] ^ n[36402];
assign t[36403] = t[36402] ^ n[36403];
assign t[36404] = t[36403] ^ n[36404];
assign t[36405] = t[36404] ^ n[36405];
assign t[36406] = t[36405] ^ n[36406];
assign t[36407] = t[36406] ^ n[36407];
assign t[36408] = t[36407] ^ n[36408];
assign t[36409] = t[36408] ^ n[36409];
assign t[36410] = t[36409] ^ n[36410];
assign t[36411] = t[36410] ^ n[36411];
assign t[36412] = t[36411] ^ n[36412];
assign t[36413] = t[36412] ^ n[36413];
assign t[36414] = t[36413] ^ n[36414];
assign t[36415] = t[36414] ^ n[36415];
assign t[36416] = t[36415] ^ n[36416];
assign t[36417] = t[36416] ^ n[36417];
assign t[36418] = t[36417] ^ n[36418];
assign t[36419] = t[36418] ^ n[36419];
assign t[36420] = t[36419] ^ n[36420];
assign t[36421] = t[36420] ^ n[36421];
assign t[36422] = t[36421] ^ n[36422];
assign t[36423] = t[36422] ^ n[36423];
assign t[36424] = t[36423] ^ n[36424];
assign t[36425] = t[36424] ^ n[36425];
assign t[36426] = t[36425] ^ n[36426];
assign t[36427] = t[36426] ^ n[36427];
assign t[36428] = t[36427] ^ n[36428];
assign t[36429] = t[36428] ^ n[36429];
assign t[36430] = t[36429] ^ n[36430];
assign t[36431] = t[36430] ^ n[36431];
assign t[36432] = t[36431] ^ n[36432];
assign t[36433] = t[36432] ^ n[36433];
assign t[36434] = t[36433] ^ n[36434];
assign t[36435] = t[36434] ^ n[36435];
assign t[36436] = t[36435] ^ n[36436];
assign t[36437] = t[36436] ^ n[36437];
assign t[36438] = t[36437] ^ n[36438];
assign t[36439] = t[36438] ^ n[36439];
assign t[36440] = t[36439] ^ n[36440];
assign t[36441] = t[36440] ^ n[36441];
assign t[36442] = t[36441] ^ n[36442];
assign t[36443] = t[36442] ^ n[36443];
assign t[36444] = t[36443] ^ n[36444];
assign t[36445] = t[36444] ^ n[36445];
assign t[36446] = t[36445] ^ n[36446];
assign t[36447] = t[36446] ^ n[36447];
assign t[36448] = t[36447] ^ n[36448];
assign t[36449] = t[36448] ^ n[36449];
assign t[36450] = t[36449] ^ n[36450];
assign t[36451] = t[36450] ^ n[36451];
assign t[36452] = t[36451] ^ n[36452];
assign t[36453] = t[36452] ^ n[36453];
assign t[36454] = t[36453] ^ n[36454];
assign t[36455] = t[36454] ^ n[36455];
assign t[36456] = t[36455] ^ n[36456];
assign t[36457] = t[36456] ^ n[36457];
assign t[36458] = t[36457] ^ n[36458];
assign t[36459] = t[36458] ^ n[36459];
assign t[36460] = t[36459] ^ n[36460];
assign t[36461] = t[36460] ^ n[36461];
assign t[36462] = t[36461] ^ n[36462];
assign t[36463] = t[36462] ^ n[36463];
assign t[36464] = t[36463] ^ n[36464];
assign t[36465] = t[36464] ^ n[36465];
assign t[36466] = t[36465] ^ n[36466];
assign t[36467] = t[36466] ^ n[36467];
assign t[36468] = t[36467] ^ n[36468];
assign t[36469] = t[36468] ^ n[36469];
assign t[36470] = t[36469] ^ n[36470];
assign t[36471] = t[36470] ^ n[36471];
assign t[36472] = t[36471] ^ n[36472];
assign t[36473] = t[36472] ^ n[36473];
assign t[36474] = t[36473] ^ n[36474];
assign t[36475] = t[36474] ^ n[36475];
assign t[36476] = t[36475] ^ n[36476];
assign t[36477] = t[36476] ^ n[36477];
assign t[36478] = t[36477] ^ n[36478];
assign t[36479] = t[36478] ^ n[36479];
assign t[36480] = t[36479] ^ n[36480];
assign t[36481] = t[36480] ^ n[36481];
assign t[36482] = t[36481] ^ n[36482];
assign t[36483] = t[36482] ^ n[36483];
assign t[36484] = t[36483] ^ n[36484];
assign t[36485] = t[36484] ^ n[36485];
assign t[36486] = t[36485] ^ n[36486];
assign t[36487] = t[36486] ^ n[36487];
assign t[36488] = t[36487] ^ n[36488];
assign t[36489] = t[36488] ^ n[36489];
assign t[36490] = t[36489] ^ n[36490];
assign t[36491] = t[36490] ^ n[36491];
assign t[36492] = t[36491] ^ n[36492];
assign t[36493] = t[36492] ^ n[36493];
assign t[36494] = t[36493] ^ n[36494];
assign t[36495] = t[36494] ^ n[36495];
assign t[36496] = t[36495] ^ n[36496];
assign t[36497] = t[36496] ^ n[36497];
assign t[36498] = t[36497] ^ n[36498];
assign t[36499] = t[36498] ^ n[36499];
assign t[36500] = t[36499] ^ n[36500];
assign t[36501] = t[36500] ^ n[36501];
assign t[36502] = t[36501] ^ n[36502];
assign t[36503] = t[36502] ^ n[36503];
assign t[36504] = t[36503] ^ n[36504];
assign t[36505] = t[36504] ^ n[36505];
assign t[36506] = t[36505] ^ n[36506];
assign t[36507] = t[36506] ^ n[36507];
assign t[36508] = t[36507] ^ n[36508];
assign t[36509] = t[36508] ^ n[36509];
assign t[36510] = t[36509] ^ n[36510];
assign t[36511] = t[36510] ^ n[36511];
assign t[36512] = t[36511] ^ n[36512];
assign t[36513] = t[36512] ^ n[36513];
assign t[36514] = t[36513] ^ n[36514];
assign t[36515] = t[36514] ^ n[36515];
assign t[36516] = t[36515] ^ n[36516];
assign t[36517] = t[36516] ^ n[36517];
assign t[36518] = t[36517] ^ n[36518];
assign t[36519] = t[36518] ^ n[36519];
assign t[36520] = t[36519] ^ n[36520];
assign t[36521] = t[36520] ^ n[36521];
assign t[36522] = t[36521] ^ n[36522];
assign t[36523] = t[36522] ^ n[36523];
assign t[36524] = t[36523] ^ n[36524];
assign t[36525] = t[36524] ^ n[36525];
assign t[36526] = t[36525] ^ n[36526];
assign t[36527] = t[36526] ^ n[36527];
assign t[36528] = t[36527] ^ n[36528];
assign t[36529] = t[36528] ^ n[36529];
assign t[36530] = t[36529] ^ n[36530];
assign t[36531] = t[36530] ^ n[36531];
assign t[36532] = t[36531] ^ n[36532];
assign t[36533] = t[36532] ^ n[36533];
assign t[36534] = t[36533] ^ n[36534];
assign t[36535] = t[36534] ^ n[36535];
assign t[36536] = t[36535] ^ n[36536];
assign t[36537] = t[36536] ^ n[36537];
assign t[36538] = t[36537] ^ n[36538];
assign t[36539] = t[36538] ^ n[36539];
assign t[36540] = t[36539] ^ n[36540];
assign t[36541] = t[36540] ^ n[36541];
assign t[36542] = t[36541] ^ n[36542];
assign t[36543] = t[36542] ^ n[36543];
assign t[36544] = t[36543] ^ n[36544];
assign t[36545] = t[36544] ^ n[36545];
assign t[36546] = t[36545] ^ n[36546];
assign t[36547] = t[36546] ^ n[36547];
assign t[36548] = t[36547] ^ n[36548];
assign t[36549] = t[36548] ^ n[36549];
assign t[36550] = t[36549] ^ n[36550];
assign t[36551] = t[36550] ^ n[36551];
assign t[36552] = t[36551] ^ n[36552];
assign t[36553] = t[36552] ^ n[36553];
assign t[36554] = t[36553] ^ n[36554];
assign t[36555] = t[36554] ^ n[36555];
assign t[36556] = t[36555] ^ n[36556];
assign t[36557] = t[36556] ^ n[36557];
assign t[36558] = t[36557] ^ n[36558];
assign t[36559] = t[36558] ^ n[36559];
assign t[36560] = t[36559] ^ n[36560];
assign t[36561] = t[36560] ^ n[36561];
assign t[36562] = t[36561] ^ n[36562];
assign t[36563] = t[36562] ^ n[36563];
assign t[36564] = t[36563] ^ n[36564];
assign t[36565] = t[36564] ^ n[36565];
assign t[36566] = t[36565] ^ n[36566];
assign t[36567] = t[36566] ^ n[36567];
assign t[36568] = t[36567] ^ n[36568];
assign t[36569] = t[36568] ^ n[36569];
assign t[36570] = t[36569] ^ n[36570];
assign t[36571] = t[36570] ^ n[36571];
assign t[36572] = t[36571] ^ n[36572];
assign t[36573] = t[36572] ^ n[36573];
assign t[36574] = t[36573] ^ n[36574];
assign t[36575] = t[36574] ^ n[36575];
assign t[36576] = t[36575] ^ n[36576];
assign t[36577] = t[36576] ^ n[36577];
assign t[36578] = t[36577] ^ n[36578];
assign t[36579] = t[36578] ^ n[36579];
assign t[36580] = t[36579] ^ n[36580];
assign t[36581] = t[36580] ^ n[36581];
assign t[36582] = t[36581] ^ n[36582];
assign t[36583] = t[36582] ^ n[36583];
assign t[36584] = t[36583] ^ n[36584];
assign t[36585] = t[36584] ^ n[36585];
assign t[36586] = t[36585] ^ n[36586];
assign t[36587] = t[36586] ^ n[36587];
assign t[36588] = t[36587] ^ n[36588];
assign t[36589] = t[36588] ^ n[36589];
assign t[36590] = t[36589] ^ n[36590];
assign t[36591] = t[36590] ^ n[36591];
assign t[36592] = t[36591] ^ n[36592];
assign t[36593] = t[36592] ^ n[36593];
assign t[36594] = t[36593] ^ n[36594];
assign t[36595] = t[36594] ^ n[36595];
assign t[36596] = t[36595] ^ n[36596];
assign t[36597] = t[36596] ^ n[36597];
assign t[36598] = t[36597] ^ n[36598];
assign t[36599] = t[36598] ^ n[36599];
assign t[36600] = t[36599] ^ n[36600];
assign t[36601] = t[36600] ^ n[36601];
assign t[36602] = t[36601] ^ n[36602];
assign t[36603] = t[36602] ^ n[36603];
assign t[36604] = t[36603] ^ n[36604];
assign t[36605] = t[36604] ^ n[36605];
assign t[36606] = t[36605] ^ n[36606];
assign t[36607] = t[36606] ^ n[36607];
assign t[36608] = t[36607] ^ n[36608];
assign t[36609] = t[36608] ^ n[36609];
assign t[36610] = t[36609] ^ n[36610];
assign t[36611] = t[36610] ^ n[36611];
assign t[36612] = t[36611] ^ n[36612];
assign t[36613] = t[36612] ^ n[36613];
assign t[36614] = t[36613] ^ n[36614];
assign t[36615] = t[36614] ^ n[36615];
assign t[36616] = t[36615] ^ n[36616];
assign t[36617] = t[36616] ^ n[36617];
assign t[36618] = t[36617] ^ n[36618];
assign t[36619] = t[36618] ^ n[36619];
assign t[36620] = t[36619] ^ n[36620];
assign t[36621] = t[36620] ^ n[36621];
assign t[36622] = t[36621] ^ n[36622];
assign t[36623] = t[36622] ^ n[36623];
assign t[36624] = t[36623] ^ n[36624];
assign t[36625] = t[36624] ^ n[36625];
assign t[36626] = t[36625] ^ n[36626];
assign t[36627] = t[36626] ^ n[36627];
assign t[36628] = t[36627] ^ n[36628];
assign t[36629] = t[36628] ^ n[36629];
assign t[36630] = t[36629] ^ n[36630];
assign t[36631] = t[36630] ^ n[36631];
assign t[36632] = t[36631] ^ n[36632];
assign t[36633] = t[36632] ^ n[36633];
assign t[36634] = t[36633] ^ n[36634];
assign t[36635] = t[36634] ^ n[36635];
assign t[36636] = t[36635] ^ n[36636];
assign t[36637] = t[36636] ^ n[36637];
assign t[36638] = t[36637] ^ n[36638];
assign t[36639] = t[36638] ^ n[36639];
assign t[36640] = t[36639] ^ n[36640];
assign t[36641] = t[36640] ^ n[36641];
assign t[36642] = t[36641] ^ n[36642];
assign t[36643] = t[36642] ^ n[36643];
assign t[36644] = t[36643] ^ n[36644];
assign t[36645] = t[36644] ^ n[36645];
assign t[36646] = t[36645] ^ n[36646];
assign t[36647] = t[36646] ^ n[36647];
assign t[36648] = t[36647] ^ n[36648];
assign t[36649] = t[36648] ^ n[36649];
assign t[36650] = t[36649] ^ n[36650];
assign t[36651] = t[36650] ^ n[36651];
assign t[36652] = t[36651] ^ n[36652];
assign t[36653] = t[36652] ^ n[36653];
assign t[36654] = t[36653] ^ n[36654];
assign t[36655] = t[36654] ^ n[36655];
assign t[36656] = t[36655] ^ n[36656];
assign t[36657] = t[36656] ^ n[36657];
assign t[36658] = t[36657] ^ n[36658];
assign t[36659] = t[36658] ^ n[36659];
assign t[36660] = t[36659] ^ n[36660];
assign t[36661] = t[36660] ^ n[36661];
assign t[36662] = t[36661] ^ n[36662];
assign t[36663] = t[36662] ^ n[36663];
assign t[36664] = t[36663] ^ n[36664];
assign t[36665] = t[36664] ^ n[36665];
assign t[36666] = t[36665] ^ n[36666];
assign t[36667] = t[36666] ^ n[36667];
assign t[36668] = t[36667] ^ n[36668];
assign t[36669] = t[36668] ^ n[36669];
assign t[36670] = t[36669] ^ n[36670];
assign t[36671] = t[36670] ^ n[36671];
assign t[36672] = t[36671] ^ n[36672];
assign t[36673] = t[36672] ^ n[36673];
assign t[36674] = t[36673] ^ n[36674];
assign t[36675] = t[36674] ^ n[36675];
assign t[36676] = t[36675] ^ n[36676];
assign t[36677] = t[36676] ^ n[36677];
assign t[36678] = t[36677] ^ n[36678];
assign t[36679] = t[36678] ^ n[36679];
assign t[36680] = t[36679] ^ n[36680];
assign t[36681] = t[36680] ^ n[36681];
assign t[36682] = t[36681] ^ n[36682];
assign t[36683] = t[36682] ^ n[36683];
assign t[36684] = t[36683] ^ n[36684];
assign t[36685] = t[36684] ^ n[36685];
assign t[36686] = t[36685] ^ n[36686];
assign t[36687] = t[36686] ^ n[36687];
assign t[36688] = t[36687] ^ n[36688];
assign t[36689] = t[36688] ^ n[36689];
assign t[36690] = t[36689] ^ n[36690];
assign t[36691] = t[36690] ^ n[36691];
assign t[36692] = t[36691] ^ n[36692];
assign t[36693] = t[36692] ^ n[36693];
assign t[36694] = t[36693] ^ n[36694];
assign t[36695] = t[36694] ^ n[36695];
assign t[36696] = t[36695] ^ n[36696];
assign t[36697] = t[36696] ^ n[36697];
assign t[36698] = t[36697] ^ n[36698];
assign t[36699] = t[36698] ^ n[36699];
assign t[36700] = t[36699] ^ n[36700];
assign t[36701] = t[36700] ^ n[36701];
assign t[36702] = t[36701] ^ n[36702];
assign t[36703] = t[36702] ^ n[36703];
assign t[36704] = t[36703] ^ n[36704];
assign t[36705] = t[36704] ^ n[36705];
assign t[36706] = t[36705] ^ n[36706];
assign t[36707] = t[36706] ^ n[36707];
assign t[36708] = t[36707] ^ n[36708];
assign t[36709] = t[36708] ^ n[36709];
assign t[36710] = t[36709] ^ n[36710];
assign t[36711] = t[36710] ^ n[36711];
assign t[36712] = t[36711] ^ n[36712];
assign t[36713] = t[36712] ^ n[36713];
assign t[36714] = t[36713] ^ n[36714];
assign t[36715] = t[36714] ^ n[36715];
assign t[36716] = t[36715] ^ n[36716];
assign t[36717] = t[36716] ^ n[36717];
assign t[36718] = t[36717] ^ n[36718];
assign t[36719] = t[36718] ^ n[36719];
assign t[36720] = t[36719] ^ n[36720];
assign t[36721] = t[36720] ^ n[36721];
assign t[36722] = t[36721] ^ n[36722];
assign t[36723] = t[36722] ^ n[36723];
assign t[36724] = t[36723] ^ n[36724];
assign t[36725] = t[36724] ^ n[36725];
assign t[36726] = t[36725] ^ n[36726];
assign t[36727] = t[36726] ^ n[36727];
assign t[36728] = t[36727] ^ n[36728];
assign t[36729] = t[36728] ^ n[36729];
assign t[36730] = t[36729] ^ n[36730];
assign t[36731] = t[36730] ^ n[36731];
assign t[36732] = t[36731] ^ n[36732];
assign t[36733] = t[36732] ^ n[36733];
assign t[36734] = t[36733] ^ n[36734];
assign t[36735] = t[36734] ^ n[36735];
assign t[36736] = t[36735] ^ n[36736];
assign t[36737] = t[36736] ^ n[36737];
assign t[36738] = t[36737] ^ n[36738];
assign t[36739] = t[36738] ^ n[36739];
assign t[36740] = t[36739] ^ n[36740];
assign t[36741] = t[36740] ^ n[36741];
assign t[36742] = t[36741] ^ n[36742];
assign t[36743] = t[36742] ^ n[36743];
assign t[36744] = t[36743] ^ n[36744];
assign t[36745] = t[36744] ^ n[36745];
assign t[36746] = t[36745] ^ n[36746];
assign t[36747] = t[36746] ^ n[36747];
assign t[36748] = t[36747] ^ n[36748];
assign t[36749] = t[36748] ^ n[36749];
assign t[36750] = t[36749] ^ n[36750];
assign t[36751] = t[36750] ^ n[36751];
assign t[36752] = t[36751] ^ n[36752];
assign t[36753] = t[36752] ^ n[36753];
assign t[36754] = t[36753] ^ n[36754];
assign t[36755] = t[36754] ^ n[36755];
assign t[36756] = t[36755] ^ n[36756];
assign t[36757] = t[36756] ^ n[36757];
assign t[36758] = t[36757] ^ n[36758];
assign t[36759] = t[36758] ^ n[36759];
assign t[36760] = t[36759] ^ n[36760];
assign t[36761] = t[36760] ^ n[36761];
assign t[36762] = t[36761] ^ n[36762];
assign t[36763] = t[36762] ^ n[36763];
assign t[36764] = t[36763] ^ n[36764];
assign t[36765] = t[36764] ^ n[36765];
assign t[36766] = t[36765] ^ n[36766];
assign t[36767] = t[36766] ^ n[36767];
assign t[36768] = t[36767] ^ n[36768];
assign t[36769] = t[36768] ^ n[36769];
assign t[36770] = t[36769] ^ n[36770];
assign t[36771] = t[36770] ^ n[36771];
assign t[36772] = t[36771] ^ n[36772];
assign t[36773] = t[36772] ^ n[36773];
assign t[36774] = t[36773] ^ n[36774];
assign t[36775] = t[36774] ^ n[36775];
assign t[36776] = t[36775] ^ n[36776];
assign t[36777] = t[36776] ^ n[36777];
assign t[36778] = t[36777] ^ n[36778];
assign t[36779] = t[36778] ^ n[36779];
assign t[36780] = t[36779] ^ n[36780];
assign t[36781] = t[36780] ^ n[36781];
assign t[36782] = t[36781] ^ n[36782];
assign t[36783] = t[36782] ^ n[36783];
assign t[36784] = t[36783] ^ n[36784];
assign t[36785] = t[36784] ^ n[36785];
assign t[36786] = t[36785] ^ n[36786];
assign t[36787] = t[36786] ^ n[36787];
assign t[36788] = t[36787] ^ n[36788];
assign t[36789] = t[36788] ^ n[36789];
assign t[36790] = t[36789] ^ n[36790];
assign t[36791] = t[36790] ^ n[36791];
assign t[36792] = t[36791] ^ n[36792];
assign t[36793] = t[36792] ^ n[36793];
assign t[36794] = t[36793] ^ n[36794];
assign t[36795] = t[36794] ^ n[36795];
assign t[36796] = t[36795] ^ n[36796];
assign t[36797] = t[36796] ^ n[36797];
assign t[36798] = t[36797] ^ n[36798];
assign t[36799] = t[36798] ^ n[36799];
assign t[36800] = t[36799] ^ n[36800];
assign t[36801] = t[36800] ^ n[36801];
assign t[36802] = t[36801] ^ n[36802];
assign t[36803] = t[36802] ^ n[36803];
assign t[36804] = t[36803] ^ n[36804];
assign t[36805] = t[36804] ^ n[36805];
assign t[36806] = t[36805] ^ n[36806];
assign t[36807] = t[36806] ^ n[36807];
assign t[36808] = t[36807] ^ n[36808];
assign t[36809] = t[36808] ^ n[36809];
assign t[36810] = t[36809] ^ n[36810];
assign t[36811] = t[36810] ^ n[36811];
assign t[36812] = t[36811] ^ n[36812];
assign t[36813] = t[36812] ^ n[36813];
assign t[36814] = t[36813] ^ n[36814];
assign t[36815] = t[36814] ^ n[36815];
assign t[36816] = t[36815] ^ n[36816];
assign t[36817] = t[36816] ^ n[36817];
assign t[36818] = t[36817] ^ n[36818];
assign t[36819] = t[36818] ^ n[36819];
assign t[36820] = t[36819] ^ n[36820];
assign t[36821] = t[36820] ^ n[36821];
assign t[36822] = t[36821] ^ n[36822];
assign t[36823] = t[36822] ^ n[36823];
assign t[36824] = t[36823] ^ n[36824];
assign t[36825] = t[36824] ^ n[36825];
assign t[36826] = t[36825] ^ n[36826];
assign t[36827] = t[36826] ^ n[36827];
assign t[36828] = t[36827] ^ n[36828];
assign t[36829] = t[36828] ^ n[36829];
assign t[36830] = t[36829] ^ n[36830];
assign t[36831] = t[36830] ^ n[36831];
assign t[36832] = t[36831] ^ n[36832];
assign t[36833] = t[36832] ^ n[36833];
assign t[36834] = t[36833] ^ n[36834];
assign t[36835] = t[36834] ^ n[36835];
assign t[36836] = t[36835] ^ n[36836];
assign t[36837] = t[36836] ^ n[36837];
assign t[36838] = t[36837] ^ n[36838];
assign t[36839] = t[36838] ^ n[36839];
assign t[36840] = t[36839] ^ n[36840];
assign t[36841] = t[36840] ^ n[36841];
assign t[36842] = t[36841] ^ n[36842];
assign t[36843] = t[36842] ^ n[36843];
assign t[36844] = t[36843] ^ n[36844];
assign t[36845] = t[36844] ^ n[36845];
assign t[36846] = t[36845] ^ n[36846];
assign t[36847] = t[36846] ^ n[36847];
assign t[36848] = t[36847] ^ n[36848];
assign t[36849] = t[36848] ^ n[36849];
assign t[36850] = t[36849] ^ n[36850];
assign t[36851] = t[36850] ^ n[36851];
assign t[36852] = t[36851] ^ n[36852];
assign t[36853] = t[36852] ^ n[36853];
assign t[36854] = t[36853] ^ n[36854];
assign t[36855] = t[36854] ^ n[36855];
assign t[36856] = t[36855] ^ n[36856];
assign t[36857] = t[36856] ^ n[36857];
assign t[36858] = t[36857] ^ n[36858];
assign t[36859] = t[36858] ^ n[36859];
assign t[36860] = t[36859] ^ n[36860];
assign t[36861] = t[36860] ^ n[36861];
assign t[36862] = t[36861] ^ n[36862];
assign t[36863] = t[36862] ^ n[36863];
assign t[36864] = t[36863] ^ n[36864];
assign t[36865] = t[36864] ^ n[36865];
assign t[36866] = t[36865] ^ n[36866];
assign t[36867] = t[36866] ^ n[36867];
assign t[36868] = t[36867] ^ n[36868];
assign t[36869] = t[36868] ^ n[36869];
assign t[36870] = t[36869] ^ n[36870];
assign t[36871] = t[36870] ^ n[36871];
assign t[36872] = t[36871] ^ n[36872];
assign t[36873] = t[36872] ^ n[36873];
assign t[36874] = t[36873] ^ n[36874];
assign t[36875] = t[36874] ^ n[36875];
assign t[36876] = t[36875] ^ n[36876];
assign t[36877] = t[36876] ^ n[36877];
assign t[36878] = t[36877] ^ n[36878];
assign t[36879] = t[36878] ^ n[36879];
assign t[36880] = t[36879] ^ n[36880];
assign t[36881] = t[36880] ^ n[36881];
assign t[36882] = t[36881] ^ n[36882];
assign t[36883] = t[36882] ^ n[36883];
assign t[36884] = t[36883] ^ n[36884];
assign t[36885] = t[36884] ^ n[36885];
assign t[36886] = t[36885] ^ n[36886];
assign t[36887] = t[36886] ^ n[36887];
assign t[36888] = t[36887] ^ n[36888];
assign t[36889] = t[36888] ^ n[36889];
assign t[36890] = t[36889] ^ n[36890];
assign t[36891] = t[36890] ^ n[36891];
assign t[36892] = t[36891] ^ n[36892];
assign t[36893] = t[36892] ^ n[36893];
assign t[36894] = t[36893] ^ n[36894];
assign t[36895] = t[36894] ^ n[36895];
assign t[36896] = t[36895] ^ n[36896];
assign t[36897] = t[36896] ^ n[36897];
assign t[36898] = t[36897] ^ n[36898];
assign t[36899] = t[36898] ^ n[36899];
assign t[36900] = t[36899] ^ n[36900];
assign t[36901] = t[36900] ^ n[36901];
assign t[36902] = t[36901] ^ n[36902];
assign t[36903] = t[36902] ^ n[36903];
assign t[36904] = t[36903] ^ n[36904];
assign t[36905] = t[36904] ^ n[36905];
assign t[36906] = t[36905] ^ n[36906];
assign t[36907] = t[36906] ^ n[36907];
assign t[36908] = t[36907] ^ n[36908];
assign t[36909] = t[36908] ^ n[36909];
assign t[36910] = t[36909] ^ n[36910];
assign t[36911] = t[36910] ^ n[36911];
assign t[36912] = t[36911] ^ n[36912];
assign t[36913] = t[36912] ^ n[36913];
assign t[36914] = t[36913] ^ n[36914];
assign t[36915] = t[36914] ^ n[36915];
assign t[36916] = t[36915] ^ n[36916];
assign t[36917] = t[36916] ^ n[36917];
assign t[36918] = t[36917] ^ n[36918];
assign t[36919] = t[36918] ^ n[36919];
assign t[36920] = t[36919] ^ n[36920];
assign t[36921] = t[36920] ^ n[36921];
assign t[36922] = t[36921] ^ n[36922];
assign t[36923] = t[36922] ^ n[36923];
assign t[36924] = t[36923] ^ n[36924];
assign t[36925] = t[36924] ^ n[36925];
assign t[36926] = t[36925] ^ n[36926];
assign t[36927] = t[36926] ^ n[36927];
assign t[36928] = t[36927] ^ n[36928];
assign t[36929] = t[36928] ^ n[36929];
assign t[36930] = t[36929] ^ n[36930];
assign t[36931] = t[36930] ^ n[36931];
assign t[36932] = t[36931] ^ n[36932];
assign t[36933] = t[36932] ^ n[36933];
assign t[36934] = t[36933] ^ n[36934];
assign t[36935] = t[36934] ^ n[36935];
assign t[36936] = t[36935] ^ n[36936];
assign t[36937] = t[36936] ^ n[36937];
assign t[36938] = t[36937] ^ n[36938];
assign t[36939] = t[36938] ^ n[36939];
assign t[36940] = t[36939] ^ n[36940];
assign t[36941] = t[36940] ^ n[36941];
assign t[36942] = t[36941] ^ n[36942];
assign t[36943] = t[36942] ^ n[36943];
assign t[36944] = t[36943] ^ n[36944];
assign t[36945] = t[36944] ^ n[36945];
assign t[36946] = t[36945] ^ n[36946];
assign t[36947] = t[36946] ^ n[36947];
assign t[36948] = t[36947] ^ n[36948];
assign t[36949] = t[36948] ^ n[36949];
assign t[36950] = t[36949] ^ n[36950];
assign t[36951] = t[36950] ^ n[36951];
assign t[36952] = t[36951] ^ n[36952];
assign t[36953] = t[36952] ^ n[36953];
assign t[36954] = t[36953] ^ n[36954];
assign t[36955] = t[36954] ^ n[36955];
assign t[36956] = t[36955] ^ n[36956];
assign t[36957] = t[36956] ^ n[36957];
assign t[36958] = t[36957] ^ n[36958];
assign t[36959] = t[36958] ^ n[36959];
assign t[36960] = t[36959] ^ n[36960];
assign t[36961] = t[36960] ^ n[36961];
assign t[36962] = t[36961] ^ n[36962];
assign t[36963] = t[36962] ^ n[36963];
assign t[36964] = t[36963] ^ n[36964];
assign t[36965] = t[36964] ^ n[36965];
assign t[36966] = t[36965] ^ n[36966];
assign t[36967] = t[36966] ^ n[36967];
assign t[36968] = t[36967] ^ n[36968];
assign t[36969] = t[36968] ^ n[36969];
assign t[36970] = t[36969] ^ n[36970];
assign t[36971] = t[36970] ^ n[36971];
assign t[36972] = t[36971] ^ n[36972];
assign t[36973] = t[36972] ^ n[36973];
assign t[36974] = t[36973] ^ n[36974];
assign t[36975] = t[36974] ^ n[36975];
assign t[36976] = t[36975] ^ n[36976];
assign t[36977] = t[36976] ^ n[36977];
assign t[36978] = t[36977] ^ n[36978];
assign t[36979] = t[36978] ^ n[36979];
assign t[36980] = t[36979] ^ n[36980];
assign t[36981] = t[36980] ^ n[36981];
assign t[36982] = t[36981] ^ n[36982];
assign t[36983] = t[36982] ^ n[36983];
assign t[36984] = t[36983] ^ n[36984];
assign t[36985] = t[36984] ^ n[36985];
assign t[36986] = t[36985] ^ n[36986];
assign t[36987] = t[36986] ^ n[36987];
assign t[36988] = t[36987] ^ n[36988];
assign t[36989] = t[36988] ^ n[36989];
assign t[36990] = t[36989] ^ n[36990];
assign t[36991] = t[36990] ^ n[36991];
assign t[36992] = t[36991] ^ n[36992];
assign t[36993] = t[36992] ^ n[36993];
assign t[36994] = t[36993] ^ n[36994];
assign t[36995] = t[36994] ^ n[36995];
assign t[36996] = t[36995] ^ n[36996];
assign t[36997] = t[36996] ^ n[36997];
assign t[36998] = t[36997] ^ n[36998];
assign t[36999] = t[36998] ^ n[36999];
assign t[37000] = t[36999] ^ n[37000];
assign t[37001] = t[37000] ^ n[37001];
assign t[37002] = t[37001] ^ n[37002];
assign t[37003] = t[37002] ^ n[37003];
assign t[37004] = t[37003] ^ n[37004];
assign t[37005] = t[37004] ^ n[37005];
assign t[37006] = t[37005] ^ n[37006];
assign t[37007] = t[37006] ^ n[37007];
assign t[37008] = t[37007] ^ n[37008];
assign t[37009] = t[37008] ^ n[37009];
assign t[37010] = t[37009] ^ n[37010];
assign t[37011] = t[37010] ^ n[37011];
assign t[37012] = t[37011] ^ n[37012];
assign t[37013] = t[37012] ^ n[37013];
assign t[37014] = t[37013] ^ n[37014];
assign t[37015] = t[37014] ^ n[37015];
assign t[37016] = t[37015] ^ n[37016];
assign t[37017] = t[37016] ^ n[37017];
assign t[37018] = t[37017] ^ n[37018];
assign t[37019] = t[37018] ^ n[37019];
assign t[37020] = t[37019] ^ n[37020];
assign t[37021] = t[37020] ^ n[37021];
assign t[37022] = t[37021] ^ n[37022];
assign t[37023] = t[37022] ^ n[37023];
assign t[37024] = t[37023] ^ n[37024];
assign t[37025] = t[37024] ^ n[37025];
assign t[37026] = t[37025] ^ n[37026];
assign t[37027] = t[37026] ^ n[37027];
assign t[37028] = t[37027] ^ n[37028];
assign t[37029] = t[37028] ^ n[37029];
assign t[37030] = t[37029] ^ n[37030];
assign t[37031] = t[37030] ^ n[37031];
assign t[37032] = t[37031] ^ n[37032];
assign t[37033] = t[37032] ^ n[37033];
assign t[37034] = t[37033] ^ n[37034];
assign t[37035] = t[37034] ^ n[37035];
assign t[37036] = t[37035] ^ n[37036];
assign t[37037] = t[37036] ^ n[37037];
assign t[37038] = t[37037] ^ n[37038];
assign t[37039] = t[37038] ^ n[37039];
assign t[37040] = t[37039] ^ n[37040];
assign t[37041] = t[37040] ^ n[37041];
assign t[37042] = t[37041] ^ n[37042];
assign t[37043] = t[37042] ^ n[37043];
assign t[37044] = t[37043] ^ n[37044];
assign t[37045] = t[37044] ^ n[37045];
assign t[37046] = t[37045] ^ n[37046];
assign t[37047] = t[37046] ^ n[37047];
assign t[37048] = t[37047] ^ n[37048];
assign t[37049] = t[37048] ^ n[37049];
assign t[37050] = t[37049] ^ n[37050];
assign t[37051] = t[37050] ^ n[37051];
assign t[37052] = t[37051] ^ n[37052];
assign t[37053] = t[37052] ^ n[37053];
assign t[37054] = t[37053] ^ n[37054];
assign t[37055] = t[37054] ^ n[37055];
assign t[37056] = t[37055] ^ n[37056];
assign t[37057] = t[37056] ^ n[37057];
assign t[37058] = t[37057] ^ n[37058];
assign t[37059] = t[37058] ^ n[37059];
assign t[37060] = t[37059] ^ n[37060];
assign t[37061] = t[37060] ^ n[37061];
assign t[37062] = t[37061] ^ n[37062];
assign t[37063] = t[37062] ^ n[37063];
assign t[37064] = t[37063] ^ n[37064];
assign t[37065] = t[37064] ^ n[37065];
assign t[37066] = t[37065] ^ n[37066];
assign t[37067] = t[37066] ^ n[37067];
assign t[37068] = t[37067] ^ n[37068];
assign t[37069] = t[37068] ^ n[37069];
assign t[37070] = t[37069] ^ n[37070];
assign t[37071] = t[37070] ^ n[37071];
assign t[37072] = t[37071] ^ n[37072];
assign t[37073] = t[37072] ^ n[37073];
assign t[37074] = t[37073] ^ n[37074];
assign t[37075] = t[37074] ^ n[37075];
assign t[37076] = t[37075] ^ n[37076];
assign t[37077] = t[37076] ^ n[37077];
assign t[37078] = t[37077] ^ n[37078];
assign t[37079] = t[37078] ^ n[37079];
assign t[37080] = t[37079] ^ n[37080];
assign t[37081] = t[37080] ^ n[37081];
assign t[37082] = t[37081] ^ n[37082];
assign t[37083] = t[37082] ^ n[37083];
assign t[37084] = t[37083] ^ n[37084];
assign t[37085] = t[37084] ^ n[37085];
assign t[37086] = t[37085] ^ n[37086];
assign t[37087] = t[37086] ^ n[37087];
assign t[37088] = t[37087] ^ n[37088];
assign t[37089] = t[37088] ^ n[37089];
assign t[37090] = t[37089] ^ n[37090];
assign t[37091] = t[37090] ^ n[37091];
assign t[37092] = t[37091] ^ n[37092];
assign t[37093] = t[37092] ^ n[37093];
assign t[37094] = t[37093] ^ n[37094];
assign t[37095] = t[37094] ^ n[37095];
assign t[37096] = t[37095] ^ n[37096];
assign t[37097] = t[37096] ^ n[37097];
assign t[37098] = t[37097] ^ n[37098];
assign t[37099] = t[37098] ^ n[37099];
assign t[37100] = t[37099] ^ n[37100];
assign t[37101] = t[37100] ^ n[37101];
assign t[37102] = t[37101] ^ n[37102];
assign t[37103] = t[37102] ^ n[37103];
assign t[37104] = t[37103] ^ n[37104];
assign t[37105] = t[37104] ^ n[37105];
assign t[37106] = t[37105] ^ n[37106];
assign t[37107] = t[37106] ^ n[37107];
assign t[37108] = t[37107] ^ n[37108];
assign t[37109] = t[37108] ^ n[37109];
assign t[37110] = t[37109] ^ n[37110];
assign t[37111] = t[37110] ^ n[37111];
assign t[37112] = t[37111] ^ n[37112];
assign t[37113] = t[37112] ^ n[37113];
assign t[37114] = t[37113] ^ n[37114];
assign t[37115] = t[37114] ^ n[37115];
assign t[37116] = t[37115] ^ n[37116];
assign t[37117] = t[37116] ^ n[37117];
assign t[37118] = t[37117] ^ n[37118];
assign t[37119] = t[37118] ^ n[37119];
assign t[37120] = t[37119] ^ n[37120];
assign t[37121] = t[37120] ^ n[37121];
assign t[37122] = t[37121] ^ n[37122];
assign t[37123] = t[37122] ^ n[37123];
assign t[37124] = t[37123] ^ n[37124];
assign t[37125] = t[37124] ^ n[37125];
assign t[37126] = t[37125] ^ n[37126];
assign t[37127] = t[37126] ^ n[37127];
assign t[37128] = t[37127] ^ n[37128];
assign t[37129] = t[37128] ^ n[37129];
assign t[37130] = t[37129] ^ n[37130];
assign t[37131] = t[37130] ^ n[37131];
assign t[37132] = t[37131] ^ n[37132];
assign t[37133] = t[37132] ^ n[37133];
assign t[37134] = t[37133] ^ n[37134];
assign t[37135] = t[37134] ^ n[37135];
assign t[37136] = t[37135] ^ n[37136];
assign t[37137] = t[37136] ^ n[37137];
assign t[37138] = t[37137] ^ n[37138];
assign t[37139] = t[37138] ^ n[37139];
assign t[37140] = t[37139] ^ n[37140];
assign t[37141] = t[37140] ^ n[37141];
assign t[37142] = t[37141] ^ n[37142];
assign t[37143] = t[37142] ^ n[37143];
assign t[37144] = t[37143] ^ n[37144];
assign t[37145] = t[37144] ^ n[37145];
assign t[37146] = t[37145] ^ n[37146];
assign t[37147] = t[37146] ^ n[37147];
assign t[37148] = t[37147] ^ n[37148];
assign t[37149] = t[37148] ^ n[37149];
assign t[37150] = t[37149] ^ n[37150];
assign t[37151] = t[37150] ^ n[37151];
assign t[37152] = t[37151] ^ n[37152];
assign t[37153] = t[37152] ^ n[37153];
assign t[37154] = t[37153] ^ n[37154];
assign t[37155] = t[37154] ^ n[37155];
assign t[37156] = t[37155] ^ n[37156];
assign t[37157] = t[37156] ^ n[37157];
assign t[37158] = t[37157] ^ n[37158];
assign t[37159] = t[37158] ^ n[37159];
assign t[37160] = t[37159] ^ n[37160];
assign t[37161] = t[37160] ^ n[37161];
assign t[37162] = t[37161] ^ n[37162];
assign t[37163] = t[37162] ^ n[37163];
assign t[37164] = t[37163] ^ n[37164];
assign t[37165] = t[37164] ^ n[37165];
assign t[37166] = t[37165] ^ n[37166];
assign t[37167] = t[37166] ^ n[37167];
assign t[37168] = t[37167] ^ n[37168];
assign t[37169] = t[37168] ^ n[37169];
assign t[37170] = t[37169] ^ n[37170];
assign t[37171] = t[37170] ^ n[37171];
assign t[37172] = t[37171] ^ n[37172];
assign t[37173] = t[37172] ^ n[37173];
assign t[37174] = t[37173] ^ n[37174];
assign t[37175] = t[37174] ^ n[37175];
assign t[37176] = t[37175] ^ n[37176];
assign t[37177] = t[37176] ^ n[37177];
assign t[37178] = t[37177] ^ n[37178];
assign t[37179] = t[37178] ^ n[37179];
assign t[37180] = t[37179] ^ n[37180];
assign t[37181] = t[37180] ^ n[37181];
assign t[37182] = t[37181] ^ n[37182];
assign t[37183] = t[37182] ^ n[37183];
assign t[37184] = t[37183] ^ n[37184];
assign t[37185] = t[37184] ^ n[37185];
assign t[37186] = t[37185] ^ n[37186];
assign t[37187] = t[37186] ^ n[37187];
assign t[37188] = t[37187] ^ n[37188];
assign t[37189] = t[37188] ^ n[37189];
assign t[37190] = t[37189] ^ n[37190];
assign t[37191] = t[37190] ^ n[37191];
assign t[37192] = t[37191] ^ n[37192];
assign t[37193] = t[37192] ^ n[37193];
assign t[37194] = t[37193] ^ n[37194];
assign t[37195] = t[37194] ^ n[37195];
assign t[37196] = t[37195] ^ n[37196];
assign t[37197] = t[37196] ^ n[37197];
assign t[37198] = t[37197] ^ n[37198];
assign t[37199] = t[37198] ^ n[37199];
assign t[37200] = t[37199] ^ n[37200];
assign t[37201] = t[37200] ^ n[37201];
assign t[37202] = t[37201] ^ n[37202];
assign t[37203] = t[37202] ^ n[37203];
assign t[37204] = t[37203] ^ n[37204];
assign t[37205] = t[37204] ^ n[37205];
assign t[37206] = t[37205] ^ n[37206];
assign t[37207] = t[37206] ^ n[37207];
assign t[37208] = t[37207] ^ n[37208];
assign t[37209] = t[37208] ^ n[37209];
assign t[37210] = t[37209] ^ n[37210];
assign t[37211] = t[37210] ^ n[37211];
assign t[37212] = t[37211] ^ n[37212];
assign t[37213] = t[37212] ^ n[37213];
assign t[37214] = t[37213] ^ n[37214];
assign t[37215] = t[37214] ^ n[37215];
assign t[37216] = t[37215] ^ n[37216];
assign t[37217] = t[37216] ^ n[37217];
assign t[37218] = t[37217] ^ n[37218];
assign t[37219] = t[37218] ^ n[37219];
assign t[37220] = t[37219] ^ n[37220];
assign t[37221] = t[37220] ^ n[37221];
assign t[37222] = t[37221] ^ n[37222];
assign t[37223] = t[37222] ^ n[37223];
assign t[37224] = t[37223] ^ n[37224];
assign t[37225] = t[37224] ^ n[37225];
assign t[37226] = t[37225] ^ n[37226];
assign t[37227] = t[37226] ^ n[37227];
assign t[37228] = t[37227] ^ n[37228];
assign t[37229] = t[37228] ^ n[37229];
assign t[37230] = t[37229] ^ n[37230];
assign t[37231] = t[37230] ^ n[37231];
assign t[37232] = t[37231] ^ n[37232];
assign t[37233] = t[37232] ^ n[37233];
assign t[37234] = t[37233] ^ n[37234];
assign t[37235] = t[37234] ^ n[37235];
assign t[37236] = t[37235] ^ n[37236];
assign t[37237] = t[37236] ^ n[37237];
assign t[37238] = t[37237] ^ n[37238];
assign t[37239] = t[37238] ^ n[37239];
assign t[37240] = t[37239] ^ n[37240];
assign t[37241] = t[37240] ^ n[37241];
assign t[37242] = t[37241] ^ n[37242];
assign t[37243] = t[37242] ^ n[37243];
assign t[37244] = t[37243] ^ n[37244];
assign t[37245] = t[37244] ^ n[37245];
assign t[37246] = t[37245] ^ n[37246];
assign t[37247] = t[37246] ^ n[37247];
assign t[37248] = t[37247] ^ n[37248];
assign t[37249] = t[37248] ^ n[37249];
assign t[37250] = t[37249] ^ n[37250];
assign t[37251] = t[37250] ^ n[37251];
assign t[37252] = t[37251] ^ n[37252];
assign t[37253] = t[37252] ^ n[37253];
assign t[37254] = t[37253] ^ n[37254];
assign t[37255] = t[37254] ^ n[37255];
assign t[37256] = t[37255] ^ n[37256];
assign t[37257] = t[37256] ^ n[37257];
assign t[37258] = t[37257] ^ n[37258];
assign t[37259] = t[37258] ^ n[37259];
assign t[37260] = t[37259] ^ n[37260];
assign t[37261] = t[37260] ^ n[37261];
assign t[37262] = t[37261] ^ n[37262];
assign t[37263] = t[37262] ^ n[37263];
assign t[37264] = t[37263] ^ n[37264];
assign t[37265] = t[37264] ^ n[37265];
assign t[37266] = t[37265] ^ n[37266];
assign t[37267] = t[37266] ^ n[37267];
assign t[37268] = t[37267] ^ n[37268];
assign t[37269] = t[37268] ^ n[37269];
assign t[37270] = t[37269] ^ n[37270];
assign t[37271] = t[37270] ^ n[37271];
assign t[37272] = t[37271] ^ n[37272];
assign t[37273] = t[37272] ^ n[37273];
assign t[37274] = t[37273] ^ n[37274];
assign t[37275] = t[37274] ^ n[37275];
assign t[37276] = t[37275] ^ n[37276];
assign t[37277] = t[37276] ^ n[37277];
assign t[37278] = t[37277] ^ n[37278];
assign t[37279] = t[37278] ^ n[37279];
assign t[37280] = t[37279] ^ n[37280];
assign t[37281] = t[37280] ^ n[37281];
assign t[37282] = t[37281] ^ n[37282];
assign t[37283] = t[37282] ^ n[37283];
assign t[37284] = t[37283] ^ n[37284];
assign t[37285] = t[37284] ^ n[37285];
assign t[37286] = t[37285] ^ n[37286];
assign t[37287] = t[37286] ^ n[37287];
assign t[37288] = t[37287] ^ n[37288];
assign t[37289] = t[37288] ^ n[37289];
assign t[37290] = t[37289] ^ n[37290];
assign t[37291] = t[37290] ^ n[37291];
assign t[37292] = t[37291] ^ n[37292];
assign t[37293] = t[37292] ^ n[37293];
assign t[37294] = t[37293] ^ n[37294];
assign t[37295] = t[37294] ^ n[37295];
assign t[37296] = t[37295] ^ n[37296];
assign t[37297] = t[37296] ^ n[37297];
assign t[37298] = t[37297] ^ n[37298];
assign t[37299] = t[37298] ^ n[37299];
assign t[37300] = t[37299] ^ n[37300];
assign t[37301] = t[37300] ^ n[37301];
assign t[37302] = t[37301] ^ n[37302];
assign t[37303] = t[37302] ^ n[37303];
assign t[37304] = t[37303] ^ n[37304];
assign t[37305] = t[37304] ^ n[37305];
assign t[37306] = t[37305] ^ n[37306];
assign t[37307] = t[37306] ^ n[37307];
assign t[37308] = t[37307] ^ n[37308];
assign t[37309] = t[37308] ^ n[37309];
assign t[37310] = t[37309] ^ n[37310];
assign t[37311] = t[37310] ^ n[37311];
assign t[37312] = t[37311] ^ n[37312];
assign t[37313] = t[37312] ^ n[37313];
assign t[37314] = t[37313] ^ n[37314];
assign t[37315] = t[37314] ^ n[37315];
assign t[37316] = t[37315] ^ n[37316];
assign t[37317] = t[37316] ^ n[37317];
assign t[37318] = t[37317] ^ n[37318];
assign t[37319] = t[37318] ^ n[37319];
assign t[37320] = t[37319] ^ n[37320];
assign t[37321] = t[37320] ^ n[37321];
assign t[37322] = t[37321] ^ n[37322];
assign t[37323] = t[37322] ^ n[37323];
assign t[37324] = t[37323] ^ n[37324];
assign t[37325] = t[37324] ^ n[37325];
assign t[37326] = t[37325] ^ n[37326];
assign t[37327] = t[37326] ^ n[37327];
assign t[37328] = t[37327] ^ n[37328];
assign t[37329] = t[37328] ^ n[37329];
assign t[37330] = t[37329] ^ n[37330];
assign t[37331] = t[37330] ^ n[37331];
assign t[37332] = t[37331] ^ n[37332];
assign t[37333] = t[37332] ^ n[37333];
assign t[37334] = t[37333] ^ n[37334];
assign t[37335] = t[37334] ^ n[37335];
assign t[37336] = t[37335] ^ n[37336];
assign t[37337] = t[37336] ^ n[37337];
assign t[37338] = t[37337] ^ n[37338];
assign t[37339] = t[37338] ^ n[37339];
assign t[37340] = t[37339] ^ n[37340];
assign t[37341] = t[37340] ^ n[37341];
assign t[37342] = t[37341] ^ n[37342];
assign t[37343] = t[37342] ^ n[37343];
assign t[37344] = t[37343] ^ n[37344];
assign t[37345] = t[37344] ^ n[37345];
assign t[37346] = t[37345] ^ n[37346];
assign t[37347] = t[37346] ^ n[37347];
assign t[37348] = t[37347] ^ n[37348];
assign t[37349] = t[37348] ^ n[37349];
assign t[37350] = t[37349] ^ n[37350];
assign t[37351] = t[37350] ^ n[37351];
assign t[37352] = t[37351] ^ n[37352];
assign t[37353] = t[37352] ^ n[37353];
assign t[37354] = t[37353] ^ n[37354];
assign t[37355] = t[37354] ^ n[37355];
assign t[37356] = t[37355] ^ n[37356];
assign t[37357] = t[37356] ^ n[37357];
assign t[37358] = t[37357] ^ n[37358];
assign t[37359] = t[37358] ^ n[37359];
assign t[37360] = t[37359] ^ n[37360];
assign t[37361] = t[37360] ^ n[37361];
assign t[37362] = t[37361] ^ n[37362];
assign t[37363] = t[37362] ^ n[37363];
assign t[37364] = t[37363] ^ n[37364];
assign t[37365] = t[37364] ^ n[37365];
assign t[37366] = t[37365] ^ n[37366];
assign t[37367] = t[37366] ^ n[37367];
assign t[37368] = t[37367] ^ n[37368];
assign t[37369] = t[37368] ^ n[37369];
assign t[37370] = t[37369] ^ n[37370];
assign t[37371] = t[37370] ^ n[37371];
assign t[37372] = t[37371] ^ n[37372];
assign t[37373] = t[37372] ^ n[37373];
assign t[37374] = t[37373] ^ n[37374];
assign t[37375] = t[37374] ^ n[37375];
assign t[37376] = t[37375] ^ n[37376];
assign t[37377] = t[37376] ^ n[37377];
assign t[37378] = t[37377] ^ n[37378];
assign t[37379] = t[37378] ^ n[37379];
assign t[37380] = t[37379] ^ n[37380];
assign t[37381] = t[37380] ^ n[37381];
assign t[37382] = t[37381] ^ n[37382];
assign t[37383] = t[37382] ^ n[37383];
assign t[37384] = t[37383] ^ n[37384];
assign t[37385] = t[37384] ^ n[37385];
assign t[37386] = t[37385] ^ n[37386];
assign t[37387] = t[37386] ^ n[37387];
assign t[37388] = t[37387] ^ n[37388];
assign t[37389] = t[37388] ^ n[37389];
assign t[37390] = t[37389] ^ n[37390];
assign t[37391] = t[37390] ^ n[37391];
assign t[37392] = t[37391] ^ n[37392];
assign t[37393] = t[37392] ^ n[37393];
assign t[37394] = t[37393] ^ n[37394];
assign t[37395] = t[37394] ^ n[37395];
assign t[37396] = t[37395] ^ n[37396];
assign t[37397] = t[37396] ^ n[37397];
assign t[37398] = t[37397] ^ n[37398];
assign t[37399] = t[37398] ^ n[37399];
assign t[37400] = t[37399] ^ n[37400];
assign t[37401] = t[37400] ^ n[37401];
assign t[37402] = t[37401] ^ n[37402];
assign t[37403] = t[37402] ^ n[37403];
assign t[37404] = t[37403] ^ n[37404];
assign t[37405] = t[37404] ^ n[37405];
assign t[37406] = t[37405] ^ n[37406];
assign t[37407] = t[37406] ^ n[37407];
assign t[37408] = t[37407] ^ n[37408];
assign t[37409] = t[37408] ^ n[37409];
assign t[37410] = t[37409] ^ n[37410];
assign t[37411] = t[37410] ^ n[37411];
assign t[37412] = t[37411] ^ n[37412];
assign t[37413] = t[37412] ^ n[37413];
assign t[37414] = t[37413] ^ n[37414];
assign t[37415] = t[37414] ^ n[37415];
assign t[37416] = t[37415] ^ n[37416];
assign t[37417] = t[37416] ^ n[37417];
assign t[37418] = t[37417] ^ n[37418];
assign t[37419] = t[37418] ^ n[37419];
assign t[37420] = t[37419] ^ n[37420];
assign t[37421] = t[37420] ^ n[37421];
assign t[37422] = t[37421] ^ n[37422];
assign t[37423] = t[37422] ^ n[37423];
assign t[37424] = t[37423] ^ n[37424];
assign t[37425] = t[37424] ^ n[37425];
assign t[37426] = t[37425] ^ n[37426];
assign t[37427] = t[37426] ^ n[37427];
assign t[37428] = t[37427] ^ n[37428];
assign t[37429] = t[37428] ^ n[37429];
assign t[37430] = t[37429] ^ n[37430];
assign t[37431] = t[37430] ^ n[37431];
assign t[37432] = t[37431] ^ n[37432];
assign t[37433] = t[37432] ^ n[37433];
assign t[37434] = t[37433] ^ n[37434];
assign t[37435] = t[37434] ^ n[37435];
assign t[37436] = t[37435] ^ n[37436];
assign t[37437] = t[37436] ^ n[37437];
assign t[37438] = t[37437] ^ n[37438];
assign t[37439] = t[37438] ^ n[37439];
assign t[37440] = t[37439] ^ n[37440];
assign t[37441] = t[37440] ^ n[37441];
assign t[37442] = t[37441] ^ n[37442];
assign t[37443] = t[37442] ^ n[37443];
assign t[37444] = t[37443] ^ n[37444];
assign t[37445] = t[37444] ^ n[37445];
assign t[37446] = t[37445] ^ n[37446];
assign t[37447] = t[37446] ^ n[37447];
assign t[37448] = t[37447] ^ n[37448];
assign t[37449] = t[37448] ^ n[37449];
assign t[37450] = t[37449] ^ n[37450];
assign t[37451] = t[37450] ^ n[37451];
assign t[37452] = t[37451] ^ n[37452];
assign t[37453] = t[37452] ^ n[37453];
assign t[37454] = t[37453] ^ n[37454];
assign t[37455] = t[37454] ^ n[37455];
assign t[37456] = t[37455] ^ n[37456];
assign t[37457] = t[37456] ^ n[37457];
assign t[37458] = t[37457] ^ n[37458];
assign t[37459] = t[37458] ^ n[37459];
assign t[37460] = t[37459] ^ n[37460];
assign t[37461] = t[37460] ^ n[37461];
assign t[37462] = t[37461] ^ n[37462];
assign t[37463] = t[37462] ^ n[37463];
assign t[37464] = t[37463] ^ n[37464];
assign t[37465] = t[37464] ^ n[37465];
assign t[37466] = t[37465] ^ n[37466];
assign t[37467] = t[37466] ^ n[37467];
assign t[37468] = t[37467] ^ n[37468];
assign t[37469] = t[37468] ^ n[37469];
assign t[37470] = t[37469] ^ n[37470];
assign t[37471] = t[37470] ^ n[37471];
assign t[37472] = t[37471] ^ n[37472];
assign t[37473] = t[37472] ^ n[37473];
assign t[37474] = t[37473] ^ n[37474];
assign t[37475] = t[37474] ^ n[37475];
assign t[37476] = t[37475] ^ n[37476];
assign t[37477] = t[37476] ^ n[37477];
assign t[37478] = t[37477] ^ n[37478];
assign t[37479] = t[37478] ^ n[37479];
assign t[37480] = t[37479] ^ n[37480];
assign t[37481] = t[37480] ^ n[37481];
assign t[37482] = t[37481] ^ n[37482];
assign t[37483] = t[37482] ^ n[37483];
assign t[37484] = t[37483] ^ n[37484];
assign t[37485] = t[37484] ^ n[37485];
assign t[37486] = t[37485] ^ n[37486];
assign t[37487] = t[37486] ^ n[37487];
assign t[37488] = t[37487] ^ n[37488];
assign t[37489] = t[37488] ^ n[37489];
assign t[37490] = t[37489] ^ n[37490];
assign t[37491] = t[37490] ^ n[37491];
assign t[37492] = t[37491] ^ n[37492];
assign t[37493] = t[37492] ^ n[37493];
assign t[37494] = t[37493] ^ n[37494];
assign t[37495] = t[37494] ^ n[37495];
assign t[37496] = t[37495] ^ n[37496];
assign t[37497] = t[37496] ^ n[37497];
assign t[37498] = t[37497] ^ n[37498];
assign t[37499] = t[37498] ^ n[37499];
assign t[37500] = t[37499] ^ n[37500];
assign t[37501] = t[37500] ^ n[37501];
assign t[37502] = t[37501] ^ n[37502];
assign t[37503] = t[37502] ^ n[37503];
assign t[37504] = t[37503] ^ n[37504];
assign t[37505] = t[37504] ^ n[37505];
assign t[37506] = t[37505] ^ n[37506];
assign t[37507] = t[37506] ^ n[37507];
assign t[37508] = t[37507] ^ n[37508];
assign t[37509] = t[37508] ^ n[37509];
assign t[37510] = t[37509] ^ n[37510];
assign t[37511] = t[37510] ^ n[37511];
assign t[37512] = t[37511] ^ n[37512];
assign t[37513] = t[37512] ^ n[37513];
assign t[37514] = t[37513] ^ n[37514];
assign t[37515] = t[37514] ^ n[37515];
assign t[37516] = t[37515] ^ n[37516];
assign t[37517] = t[37516] ^ n[37517];
assign t[37518] = t[37517] ^ n[37518];
assign t[37519] = t[37518] ^ n[37519];
assign t[37520] = t[37519] ^ n[37520];
assign t[37521] = t[37520] ^ n[37521];
assign t[37522] = t[37521] ^ n[37522];
assign t[37523] = t[37522] ^ n[37523];
assign t[37524] = t[37523] ^ n[37524];
assign t[37525] = t[37524] ^ n[37525];
assign t[37526] = t[37525] ^ n[37526];
assign t[37527] = t[37526] ^ n[37527];
assign t[37528] = t[37527] ^ n[37528];
assign t[37529] = t[37528] ^ n[37529];
assign t[37530] = t[37529] ^ n[37530];
assign t[37531] = t[37530] ^ n[37531];
assign t[37532] = t[37531] ^ n[37532];
assign t[37533] = t[37532] ^ n[37533];
assign t[37534] = t[37533] ^ n[37534];
assign t[37535] = t[37534] ^ n[37535];
assign t[37536] = t[37535] ^ n[37536];
assign t[37537] = t[37536] ^ n[37537];
assign t[37538] = t[37537] ^ n[37538];
assign t[37539] = t[37538] ^ n[37539];
assign t[37540] = t[37539] ^ n[37540];
assign t[37541] = t[37540] ^ n[37541];
assign t[37542] = t[37541] ^ n[37542];
assign t[37543] = t[37542] ^ n[37543];
assign t[37544] = t[37543] ^ n[37544];
assign t[37545] = t[37544] ^ n[37545];
assign t[37546] = t[37545] ^ n[37546];
assign t[37547] = t[37546] ^ n[37547];
assign t[37548] = t[37547] ^ n[37548];
assign t[37549] = t[37548] ^ n[37549];
assign t[37550] = t[37549] ^ n[37550];
assign t[37551] = t[37550] ^ n[37551];
assign t[37552] = t[37551] ^ n[37552];
assign t[37553] = t[37552] ^ n[37553];
assign t[37554] = t[37553] ^ n[37554];
assign t[37555] = t[37554] ^ n[37555];
assign t[37556] = t[37555] ^ n[37556];
assign t[37557] = t[37556] ^ n[37557];
assign t[37558] = t[37557] ^ n[37558];
assign t[37559] = t[37558] ^ n[37559];
assign t[37560] = t[37559] ^ n[37560];
assign t[37561] = t[37560] ^ n[37561];
assign t[37562] = t[37561] ^ n[37562];
assign t[37563] = t[37562] ^ n[37563];
assign t[37564] = t[37563] ^ n[37564];
assign t[37565] = t[37564] ^ n[37565];
assign t[37566] = t[37565] ^ n[37566];
assign t[37567] = t[37566] ^ n[37567];
assign t[37568] = t[37567] ^ n[37568];
assign t[37569] = t[37568] ^ n[37569];
assign t[37570] = t[37569] ^ n[37570];
assign t[37571] = t[37570] ^ n[37571];
assign t[37572] = t[37571] ^ n[37572];
assign t[37573] = t[37572] ^ n[37573];
assign t[37574] = t[37573] ^ n[37574];
assign t[37575] = t[37574] ^ n[37575];
assign t[37576] = t[37575] ^ n[37576];
assign t[37577] = t[37576] ^ n[37577];
assign t[37578] = t[37577] ^ n[37578];
assign t[37579] = t[37578] ^ n[37579];
assign t[37580] = t[37579] ^ n[37580];
assign t[37581] = t[37580] ^ n[37581];
assign t[37582] = t[37581] ^ n[37582];
assign t[37583] = t[37582] ^ n[37583];
assign t[37584] = t[37583] ^ n[37584];
assign t[37585] = t[37584] ^ n[37585];
assign t[37586] = t[37585] ^ n[37586];
assign t[37587] = t[37586] ^ n[37587];
assign t[37588] = t[37587] ^ n[37588];
assign t[37589] = t[37588] ^ n[37589];
assign t[37590] = t[37589] ^ n[37590];
assign t[37591] = t[37590] ^ n[37591];
assign t[37592] = t[37591] ^ n[37592];
assign t[37593] = t[37592] ^ n[37593];
assign t[37594] = t[37593] ^ n[37594];
assign t[37595] = t[37594] ^ n[37595];
assign t[37596] = t[37595] ^ n[37596];
assign t[37597] = t[37596] ^ n[37597];
assign t[37598] = t[37597] ^ n[37598];
assign t[37599] = t[37598] ^ n[37599];
assign t[37600] = t[37599] ^ n[37600];
assign t[37601] = t[37600] ^ n[37601];
assign t[37602] = t[37601] ^ n[37602];
assign t[37603] = t[37602] ^ n[37603];
assign t[37604] = t[37603] ^ n[37604];
assign t[37605] = t[37604] ^ n[37605];
assign t[37606] = t[37605] ^ n[37606];
assign t[37607] = t[37606] ^ n[37607];
assign t[37608] = t[37607] ^ n[37608];
assign t[37609] = t[37608] ^ n[37609];
assign t[37610] = t[37609] ^ n[37610];
assign t[37611] = t[37610] ^ n[37611];
assign t[37612] = t[37611] ^ n[37612];
assign t[37613] = t[37612] ^ n[37613];
assign t[37614] = t[37613] ^ n[37614];
assign t[37615] = t[37614] ^ n[37615];
assign t[37616] = t[37615] ^ n[37616];
assign t[37617] = t[37616] ^ n[37617];
assign t[37618] = t[37617] ^ n[37618];
assign t[37619] = t[37618] ^ n[37619];
assign t[37620] = t[37619] ^ n[37620];
assign t[37621] = t[37620] ^ n[37621];
assign t[37622] = t[37621] ^ n[37622];
assign t[37623] = t[37622] ^ n[37623];
assign t[37624] = t[37623] ^ n[37624];
assign t[37625] = t[37624] ^ n[37625];
assign t[37626] = t[37625] ^ n[37626];
assign t[37627] = t[37626] ^ n[37627];
assign t[37628] = t[37627] ^ n[37628];
assign t[37629] = t[37628] ^ n[37629];
assign t[37630] = t[37629] ^ n[37630];
assign t[37631] = t[37630] ^ n[37631];
assign t[37632] = t[37631] ^ n[37632];
assign t[37633] = t[37632] ^ n[37633];
assign t[37634] = t[37633] ^ n[37634];
assign t[37635] = t[37634] ^ n[37635];
assign t[37636] = t[37635] ^ n[37636];
assign t[37637] = t[37636] ^ n[37637];
assign t[37638] = t[37637] ^ n[37638];
assign t[37639] = t[37638] ^ n[37639];
assign t[37640] = t[37639] ^ n[37640];
assign t[37641] = t[37640] ^ n[37641];
assign t[37642] = t[37641] ^ n[37642];
assign t[37643] = t[37642] ^ n[37643];
assign t[37644] = t[37643] ^ n[37644];
assign t[37645] = t[37644] ^ n[37645];
assign t[37646] = t[37645] ^ n[37646];
assign t[37647] = t[37646] ^ n[37647];
assign t[37648] = t[37647] ^ n[37648];
assign t[37649] = t[37648] ^ n[37649];
assign t[37650] = t[37649] ^ n[37650];
assign t[37651] = t[37650] ^ n[37651];
assign t[37652] = t[37651] ^ n[37652];
assign t[37653] = t[37652] ^ n[37653];
assign t[37654] = t[37653] ^ n[37654];
assign t[37655] = t[37654] ^ n[37655];
assign t[37656] = t[37655] ^ n[37656];
assign t[37657] = t[37656] ^ n[37657];
assign t[37658] = t[37657] ^ n[37658];
assign t[37659] = t[37658] ^ n[37659];
assign t[37660] = t[37659] ^ n[37660];
assign t[37661] = t[37660] ^ n[37661];
assign t[37662] = t[37661] ^ n[37662];
assign t[37663] = t[37662] ^ n[37663];
assign t[37664] = t[37663] ^ n[37664];
assign t[37665] = t[37664] ^ n[37665];
assign t[37666] = t[37665] ^ n[37666];
assign t[37667] = t[37666] ^ n[37667];
assign t[37668] = t[37667] ^ n[37668];
assign t[37669] = t[37668] ^ n[37669];
assign t[37670] = t[37669] ^ n[37670];
assign t[37671] = t[37670] ^ n[37671];
assign t[37672] = t[37671] ^ n[37672];
assign t[37673] = t[37672] ^ n[37673];
assign t[37674] = t[37673] ^ n[37674];
assign t[37675] = t[37674] ^ n[37675];
assign t[37676] = t[37675] ^ n[37676];
assign t[37677] = t[37676] ^ n[37677];
assign t[37678] = t[37677] ^ n[37678];
assign t[37679] = t[37678] ^ n[37679];
assign t[37680] = t[37679] ^ n[37680];
assign t[37681] = t[37680] ^ n[37681];
assign t[37682] = t[37681] ^ n[37682];
assign t[37683] = t[37682] ^ n[37683];
assign t[37684] = t[37683] ^ n[37684];
assign t[37685] = t[37684] ^ n[37685];
assign t[37686] = t[37685] ^ n[37686];
assign t[37687] = t[37686] ^ n[37687];
assign t[37688] = t[37687] ^ n[37688];
assign t[37689] = t[37688] ^ n[37689];
assign t[37690] = t[37689] ^ n[37690];
assign t[37691] = t[37690] ^ n[37691];
assign t[37692] = t[37691] ^ n[37692];
assign t[37693] = t[37692] ^ n[37693];
assign t[37694] = t[37693] ^ n[37694];
assign t[37695] = t[37694] ^ n[37695];
assign t[37696] = t[37695] ^ n[37696];
assign t[37697] = t[37696] ^ n[37697];
assign t[37698] = t[37697] ^ n[37698];
assign t[37699] = t[37698] ^ n[37699];
assign t[37700] = t[37699] ^ n[37700];
assign t[37701] = t[37700] ^ n[37701];
assign t[37702] = t[37701] ^ n[37702];
assign t[37703] = t[37702] ^ n[37703];
assign t[37704] = t[37703] ^ n[37704];
assign t[37705] = t[37704] ^ n[37705];
assign t[37706] = t[37705] ^ n[37706];
assign t[37707] = t[37706] ^ n[37707];
assign t[37708] = t[37707] ^ n[37708];
assign t[37709] = t[37708] ^ n[37709];
assign t[37710] = t[37709] ^ n[37710];
assign t[37711] = t[37710] ^ n[37711];
assign t[37712] = t[37711] ^ n[37712];
assign t[37713] = t[37712] ^ n[37713];
assign t[37714] = t[37713] ^ n[37714];
assign t[37715] = t[37714] ^ n[37715];
assign t[37716] = t[37715] ^ n[37716];
assign t[37717] = t[37716] ^ n[37717];
assign t[37718] = t[37717] ^ n[37718];
assign t[37719] = t[37718] ^ n[37719];
assign t[37720] = t[37719] ^ n[37720];
assign t[37721] = t[37720] ^ n[37721];
assign t[37722] = t[37721] ^ n[37722];
assign t[37723] = t[37722] ^ n[37723];
assign t[37724] = t[37723] ^ n[37724];
assign t[37725] = t[37724] ^ n[37725];
assign t[37726] = t[37725] ^ n[37726];
assign t[37727] = t[37726] ^ n[37727];
assign t[37728] = t[37727] ^ n[37728];
assign t[37729] = t[37728] ^ n[37729];
assign t[37730] = t[37729] ^ n[37730];
assign t[37731] = t[37730] ^ n[37731];
assign t[37732] = t[37731] ^ n[37732];
assign t[37733] = t[37732] ^ n[37733];
assign t[37734] = t[37733] ^ n[37734];
assign t[37735] = t[37734] ^ n[37735];
assign t[37736] = t[37735] ^ n[37736];
assign t[37737] = t[37736] ^ n[37737];
assign t[37738] = t[37737] ^ n[37738];
assign t[37739] = t[37738] ^ n[37739];
assign t[37740] = t[37739] ^ n[37740];
assign t[37741] = t[37740] ^ n[37741];
assign t[37742] = t[37741] ^ n[37742];
assign t[37743] = t[37742] ^ n[37743];
assign t[37744] = t[37743] ^ n[37744];
assign t[37745] = t[37744] ^ n[37745];
assign t[37746] = t[37745] ^ n[37746];
assign t[37747] = t[37746] ^ n[37747];
assign t[37748] = t[37747] ^ n[37748];
assign t[37749] = t[37748] ^ n[37749];
assign t[37750] = t[37749] ^ n[37750];
assign t[37751] = t[37750] ^ n[37751];
assign t[37752] = t[37751] ^ n[37752];
assign t[37753] = t[37752] ^ n[37753];
assign t[37754] = t[37753] ^ n[37754];
assign t[37755] = t[37754] ^ n[37755];
assign t[37756] = t[37755] ^ n[37756];
assign t[37757] = t[37756] ^ n[37757];
assign t[37758] = t[37757] ^ n[37758];
assign t[37759] = t[37758] ^ n[37759];
assign t[37760] = t[37759] ^ n[37760];
assign t[37761] = t[37760] ^ n[37761];
assign t[37762] = t[37761] ^ n[37762];
assign t[37763] = t[37762] ^ n[37763];
assign t[37764] = t[37763] ^ n[37764];
assign t[37765] = t[37764] ^ n[37765];
assign t[37766] = t[37765] ^ n[37766];
assign t[37767] = t[37766] ^ n[37767];
assign t[37768] = t[37767] ^ n[37768];
assign t[37769] = t[37768] ^ n[37769];
assign t[37770] = t[37769] ^ n[37770];
assign t[37771] = t[37770] ^ n[37771];
assign t[37772] = t[37771] ^ n[37772];
assign t[37773] = t[37772] ^ n[37773];
assign t[37774] = t[37773] ^ n[37774];
assign t[37775] = t[37774] ^ n[37775];
assign t[37776] = t[37775] ^ n[37776];
assign t[37777] = t[37776] ^ n[37777];
assign t[37778] = t[37777] ^ n[37778];
assign t[37779] = t[37778] ^ n[37779];
assign t[37780] = t[37779] ^ n[37780];
assign t[37781] = t[37780] ^ n[37781];
assign t[37782] = t[37781] ^ n[37782];
assign t[37783] = t[37782] ^ n[37783];
assign t[37784] = t[37783] ^ n[37784];
assign t[37785] = t[37784] ^ n[37785];
assign t[37786] = t[37785] ^ n[37786];
assign t[37787] = t[37786] ^ n[37787];
assign t[37788] = t[37787] ^ n[37788];
assign t[37789] = t[37788] ^ n[37789];
assign t[37790] = t[37789] ^ n[37790];
assign t[37791] = t[37790] ^ n[37791];
assign t[37792] = t[37791] ^ n[37792];
assign t[37793] = t[37792] ^ n[37793];
assign t[37794] = t[37793] ^ n[37794];
assign t[37795] = t[37794] ^ n[37795];
assign t[37796] = t[37795] ^ n[37796];
assign t[37797] = t[37796] ^ n[37797];
assign t[37798] = t[37797] ^ n[37798];
assign t[37799] = t[37798] ^ n[37799];
assign t[37800] = t[37799] ^ n[37800];
assign t[37801] = t[37800] ^ n[37801];
assign t[37802] = t[37801] ^ n[37802];
assign t[37803] = t[37802] ^ n[37803];
assign t[37804] = t[37803] ^ n[37804];
assign t[37805] = t[37804] ^ n[37805];
assign t[37806] = t[37805] ^ n[37806];
assign t[37807] = t[37806] ^ n[37807];
assign t[37808] = t[37807] ^ n[37808];
assign t[37809] = t[37808] ^ n[37809];
assign t[37810] = t[37809] ^ n[37810];
assign t[37811] = t[37810] ^ n[37811];
assign t[37812] = t[37811] ^ n[37812];
assign t[37813] = t[37812] ^ n[37813];
assign t[37814] = t[37813] ^ n[37814];
assign t[37815] = t[37814] ^ n[37815];
assign t[37816] = t[37815] ^ n[37816];
assign t[37817] = t[37816] ^ n[37817];
assign t[37818] = t[37817] ^ n[37818];
assign t[37819] = t[37818] ^ n[37819];
assign t[37820] = t[37819] ^ n[37820];
assign t[37821] = t[37820] ^ n[37821];
assign t[37822] = t[37821] ^ n[37822];
assign t[37823] = t[37822] ^ n[37823];
assign t[37824] = t[37823] ^ n[37824];
assign t[37825] = t[37824] ^ n[37825];
assign t[37826] = t[37825] ^ n[37826];
assign t[37827] = t[37826] ^ n[37827];
assign t[37828] = t[37827] ^ n[37828];
assign t[37829] = t[37828] ^ n[37829];
assign t[37830] = t[37829] ^ n[37830];
assign t[37831] = t[37830] ^ n[37831];
assign t[37832] = t[37831] ^ n[37832];
assign t[37833] = t[37832] ^ n[37833];
assign t[37834] = t[37833] ^ n[37834];
assign t[37835] = t[37834] ^ n[37835];
assign t[37836] = t[37835] ^ n[37836];
assign t[37837] = t[37836] ^ n[37837];
assign t[37838] = t[37837] ^ n[37838];
assign t[37839] = t[37838] ^ n[37839];
assign t[37840] = t[37839] ^ n[37840];
assign t[37841] = t[37840] ^ n[37841];
assign t[37842] = t[37841] ^ n[37842];
assign t[37843] = t[37842] ^ n[37843];
assign t[37844] = t[37843] ^ n[37844];
assign t[37845] = t[37844] ^ n[37845];
assign t[37846] = t[37845] ^ n[37846];
assign t[37847] = t[37846] ^ n[37847];
assign t[37848] = t[37847] ^ n[37848];
assign t[37849] = t[37848] ^ n[37849];
assign t[37850] = t[37849] ^ n[37850];
assign t[37851] = t[37850] ^ n[37851];
assign t[37852] = t[37851] ^ n[37852];
assign t[37853] = t[37852] ^ n[37853];
assign t[37854] = t[37853] ^ n[37854];
assign t[37855] = t[37854] ^ n[37855];
assign t[37856] = t[37855] ^ n[37856];
assign t[37857] = t[37856] ^ n[37857];
assign t[37858] = t[37857] ^ n[37858];
assign t[37859] = t[37858] ^ n[37859];
assign t[37860] = t[37859] ^ n[37860];
assign t[37861] = t[37860] ^ n[37861];
assign t[37862] = t[37861] ^ n[37862];
assign t[37863] = t[37862] ^ n[37863];
assign t[37864] = t[37863] ^ n[37864];
assign t[37865] = t[37864] ^ n[37865];
assign t[37866] = t[37865] ^ n[37866];
assign t[37867] = t[37866] ^ n[37867];
assign t[37868] = t[37867] ^ n[37868];
assign t[37869] = t[37868] ^ n[37869];
assign t[37870] = t[37869] ^ n[37870];
assign t[37871] = t[37870] ^ n[37871];
assign t[37872] = t[37871] ^ n[37872];
assign t[37873] = t[37872] ^ n[37873];
assign t[37874] = t[37873] ^ n[37874];
assign t[37875] = t[37874] ^ n[37875];
assign t[37876] = t[37875] ^ n[37876];
assign t[37877] = t[37876] ^ n[37877];
assign t[37878] = t[37877] ^ n[37878];
assign t[37879] = t[37878] ^ n[37879];
assign t[37880] = t[37879] ^ n[37880];
assign t[37881] = t[37880] ^ n[37881];
assign t[37882] = t[37881] ^ n[37882];
assign t[37883] = t[37882] ^ n[37883];
assign t[37884] = t[37883] ^ n[37884];
assign t[37885] = t[37884] ^ n[37885];
assign t[37886] = t[37885] ^ n[37886];
assign t[37887] = t[37886] ^ n[37887];
assign t[37888] = t[37887] ^ n[37888];
assign t[37889] = t[37888] ^ n[37889];
assign t[37890] = t[37889] ^ n[37890];
assign t[37891] = t[37890] ^ n[37891];
assign t[37892] = t[37891] ^ n[37892];
assign t[37893] = t[37892] ^ n[37893];
assign t[37894] = t[37893] ^ n[37894];
assign t[37895] = t[37894] ^ n[37895];
assign t[37896] = t[37895] ^ n[37896];
assign t[37897] = t[37896] ^ n[37897];
assign t[37898] = t[37897] ^ n[37898];
assign t[37899] = t[37898] ^ n[37899];
assign t[37900] = t[37899] ^ n[37900];
assign t[37901] = t[37900] ^ n[37901];
assign t[37902] = t[37901] ^ n[37902];
assign t[37903] = t[37902] ^ n[37903];
assign t[37904] = t[37903] ^ n[37904];
assign t[37905] = t[37904] ^ n[37905];
assign t[37906] = t[37905] ^ n[37906];
assign t[37907] = t[37906] ^ n[37907];
assign t[37908] = t[37907] ^ n[37908];
assign t[37909] = t[37908] ^ n[37909];
assign t[37910] = t[37909] ^ n[37910];
assign t[37911] = t[37910] ^ n[37911];
assign t[37912] = t[37911] ^ n[37912];
assign t[37913] = t[37912] ^ n[37913];
assign t[37914] = t[37913] ^ n[37914];
assign t[37915] = t[37914] ^ n[37915];
assign t[37916] = t[37915] ^ n[37916];
assign t[37917] = t[37916] ^ n[37917];
assign t[37918] = t[37917] ^ n[37918];
assign t[37919] = t[37918] ^ n[37919];
assign t[37920] = t[37919] ^ n[37920];
assign t[37921] = t[37920] ^ n[37921];
assign t[37922] = t[37921] ^ n[37922];
assign t[37923] = t[37922] ^ n[37923];
assign t[37924] = t[37923] ^ n[37924];
assign t[37925] = t[37924] ^ n[37925];
assign t[37926] = t[37925] ^ n[37926];
assign t[37927] = t[37926] ^ n[37927];
assign t[37928] = t[37927] ^ n[37928];
assign t[37929] = t[37928] ^ n[37929];
assign t[37930] = t[37929] ^ n[37930];
assign t[37931] = t[37930] ^ n[37931];
assign t[37932] = t[37931] ^ n[37932];
assign t[37933] = t[37932] ^ n[37933];
assign t[37934] = t[37933] ^ n[37934];
assign t[37935] = t[37934] ^ n[37935];
assign t[37936] = t[37935] ^ n[37936];
assign t[37937] = t[37936] ^ n[37937];
assign t[37938] = t[37937] ^ n[37938];
assign t[37939] = t[37938] ^ n[37939];
assign t[37940] = t[37939] ^ n[37940];
assign t[37941] = t[37940] ^ n[37941];
assign t[37942] = t[37941] ^ n[37942];
assign t[37943] = t[37942] ^ n[37943];
assign t[37944] = t[37943] ^ n[37944];
assign t[37945] = t[37944] ^ n[37945];
assign t[37946] = t[37945] ^ n[37946];
assign t[37947] = t[37946] ^ n[37947];
assign t[37948] = t[37947] ^ n[37948];
assign t[37949] = t[37948] ^ n[37949];
assign t[37950] = t[37949] ^ n[37950];
assign t[37951] = t[37950] ^ n[37951];
assign t[37952] = t[37951] ^ n[37952];
assign t[37953] = t[37952] ^ n[37953];
assign t[37954] = t[37953] ^ n[37954];
assign t[37955] = t[37954] ^ n[37955];
assign t[37956] = t[37955] ^ n[37956];
assign t[37957] = t[37956] ^ n[37957];
assign t[37958] = t[37957] ^ n[37958];
assign t[37959] = t[37958] ^ n[37959];
assign t[37960] = t[37959] ^ n[37960];
assign t[37961] = t[37960] ^ n[37961];
assign t[37962] = t[37961] ^ n[37962];
assign t[37963] = t[37962] ^ n[37963];
assign t[37964] = t[37963] ^ n[37964];
assign t[37965] = t[37964] ^ n[37965];
assign t[37966] = t[37965] ^ n[37966];
assign t[37967] = t[37966] ^ n[37967];
assign t[37968] = t[37967] ^ n[37968];
assign t[37969] = t[37968] ^ n[37969];
assign t[37970] = t[37969] ^ n[37970];
assign t[37971] = t[37970] ^ n[37971];
assign t[37972] = t[37971] ^ n[37972];
assign t[37973] = t[37972] ^ n[37973];
assign t[37974] = t[37973] ^ n[37974];
assign t[37975] = t[37974] ^ n[37975];
assign t[37976] = t[37975] ^ n[37976];
assign t[37977] = t[37976] ^ n[37977];
assign t[37978] = t[37977] ^ n[37978];
assign t[37979] = t[37978] ^ n[37979];
assign t[37980] = t[37979] ^ n[37980];
assign t[37981] = t[37980] ^ n[37981];
assign t[37982] = t[37981] ^ n[37982];
assign t[37983] = t[37982] ^ n[37983];
assign t[37984] = t[37983] ^ n[37984];
assign t[37985] = t[37984] ^ n[37985];
assign t[37986] = t[37985] ^ n[37986];
assign t[37987] = t[37986] ^ n[37987];
assign t[37988] = t[37987] ^ n[37988];
assign t[37989] = t[37988] ^ n[37989];
assign t[37990] = t[37989] ^ n[37990];
assign t[37991] = t[37990] ^ n[37991];
assign t[37992] = t[37991] ^ n[37992];
assign t[37993] = t[37992] ^ n[37993];
assign t[37994] = t[37993] ^ n[37994];
assign t[37995] = t[37994] ^ n[37995];
assign t[37996] = t[37995] ^ n[37996];
assign t[37997] = t[37996] ^ n[37997];
assign t[37998] = t[37997] ^ n[37998];
assign t[37999] = t[37998] ^ n[37999];
assign t[38000] = t[37999] ^ n[38000];
assign t[38001] = t[38000] ^ n[38001];
assign t[38002] = t[38001] ^ n[38002];
assign t[38003] = t[38002] ^ n[38003];
assign t[38004] = t[38003] ^ n[38004];
assign t[38005] = t[38004] ^ n[38005];
assign t[38006] = t[38005] ^ n[38006];
assign t[38007] = t[38006] ^ n[38007];
assign t[38008] = t[38007] ^ n[38008];
assign t[38009] = t[38008] ^ n[38009];
assign t[38010] = t[38009] ^ n[38010];
assign t[38011] = t[38010] ^ n[38011];
assign t[38012] = t[38011] ^ n[38012];
assign t[38013] = t[38012] ^ n[38013];
assign t[38014] = t[38013] ^ n[38014];
assign t[38015] = t[38014] ^ n[38015];
assign t[38016] = t[38015] ^ n[38016];
assign t[38017] = t[38016] ^ n[38017];
assign t[38018] = t[38017] ^ n[38018];
assign t[38019] = t[38018] ^ n[38019];
assign t[38020] = t[38019] ^ n[38020];
assign t[38021] = t[38020] ^ n[38021];
assign t[38022] = t[38021] ^ n[38022];
assign t[38023] = t[38022] ^ n[38023];
assign t[38024] = t[38023] ^ n[38024];
assign t[38025] = t[38024] ^ n[38025];
assign t[38026] = t[38025] ^ n[38026];
assign t[38027] = t[38026] ^ n[38027];
assign t[38028] = t[38027] ^ n[38028];
assign t[38029] = t[38028] ^ n[38029];
assign t[38030] = t[38029] ^ n[38030];
assign t[38031] = t[38030] ^ n[38031];
assign t[38032] = t[38031] ^ n[38032];
assign t[38033] = t[38032] ^ n[38033];
assign t[38034] = t[38033] ^ n[38034];
assign t[38035] = t[38034] ^ n[38035];
assign t[38036] = t[38035] ^ n[38036];
assign t[38037] = t[38036] ^ n[38037];
assign t[38038] = t[38037] ^ n[38038];
assign t[38039] = t[38038] ^ n[38039];
assign t[38040] = t[38039] ^ n[38040];
assign t[38041] = t[38040] ^ n[38041];
assign t[38042] = t[38041] ^ n[38042];
assign t[38043] = t[38042] ^ n[38043];
assign t[38044] = t[38043] ^ n[38044];
assign t[38045] = t[38044] ^ n[38045];
assign t[38046] = t[38045] ^ n[38046];
assign t[38047] = t[38046] ^ n[38047];
assign t[38048] = t[38047] ^ n[38048];
assign t[38049] = t[38048] ^ n[38049];
assign t[38050] = t[38049] ^ n[38050];
assign t[38051] = t[38050] ^ n[38051];
assign t[38052] = t[38051] ^ n[38052];
assign t[38053] = t[38052] ^ n[38053];
assign t[38054] = t[38053] ^ n[38054];
assign t[38055] = t[38054] ^ n[38055];
assign t[38056] = t[38055] ^ n[38056];
assign t[38057] = t[38056] ^ n[38057];
assign t[38058] = t[38057] ^ n[38058];
assign t[38059] = t[38058] ^ n[38059];
assign t[38060] = t[38059] ^ n[38060];
assign t[38061] = t[38060] ^ n[38061];
assign t[38062] = t[38061] ^ n[38062];
assign t[38063] = t[38062] ^ n[38063];
assign t[38064] = t[38063] ^ n[38064];
assign t[38065] = t[38064] ^ n[38065];
assign t[38066] = t[38065] ^ n[38066];
assign t[38067] = t[38066] ^ n[38067];
assign t[38068] = t[38067] ^ n[38068];
assign t[38069] = t[38068] ^ n[38069];
assign t[38070] = t[38069] ^ n[38070];
assign t[38071] = t[38070] ^ n[38071];
assign t[38072] = t[38071] ^ n[38072];
assign t[38073] = t[38072] ^ n[38073];
assign t[38074] = t[38073] ^ n[38074];
assign t[38075] = t[38074] ^ n[38075];
assign t[38076] = t[38075] ^ n[38076];
assign t[38077] = t[38076] ^ n[38077];
assign t[38078] = t[38077] ^ n[38078];
assign t[38079] = t[38078] ^ n[38079];
assign t[38080] = t[38079] ^ n[38080];
assign t[38081] = t[38080] ^ n[38081];
assign t[38082] = t[38081] ^ n[38082];
assign t[38083] = t[38082] ^ n[38083];
assign t[38084] = t[38083] ^ n[38084];
assign t[38085] = t[38084] ^ n[38085];
assign t[38086] = t[38085] ^ n[38086];
assign t[38087] = t[38086] ^ n[38087];
assign t[38088] = t[38087] ^ n[38088];
assign t[38089] = t[38088] ^ n[38089];
assign t[38090] = t[38089] ^ n[38090];
assign t[38091] = t[38090] ^ n[38091];
assign t[38092] = t[38091] ^ n[38092];
assign t[38093] = t[38092] ^ n[38093];
assign t[38094] = t[38093] ^ n[38094];
assign t[38095] = t[38094] ^ n[38095];
assign t[38096] = t[38095] ^ n[38096];
assign t[38097] = t[38096] ^ n[38097];
assign t[38098] = t[38097] ^ n[38098];
assign t[38099] = t[38098] ^ n[38099];
assign t[38100] = t[38099] ^ n[38100];
assign t[38101] = t[38100] ^ n[38101];
assign t[38102] = t[38101] ^ n[38102];
assign t[38103] = t[38102] ^ n[38103];
assign t[38104] = t[38103] ^ n[38104];
assign t[38105] = t[38104] ^ n[38105];
assign t[38106] = t[38105] ^ n[38106];
assign t[38107] = t[38106] ^ n[38107];
assign t[38108] = t[38107] ^ n[38108];
assign t[38109] = t[38108] ^ n[38109];
assign t[38110] = t[38109] ^ n[38110];
assign t[38111] = t[38110] ^ n[38111];
assign t[38112] = t[38111] ^ n[38112];
assign t[38113] = t[38112] ^ n[38113];
assign t[38114] = t[38113] ^ n[38114];
assign t[38115] = t[38114] ^ n[38115];
assign t[38116] = t[38115] ^ n[38116];
assign t[38117] = t[38116] ^ n[38117];
assign t[38118] = t[38117] ^ n[38118];
assign t[38119] = t[38118] ^ n[38119];
assign t[38120] = t[38119] ^ n[38120];
assign t[38121] = t[38120] ^ n[38121];
assign t[38122] = t[38121] ^ n[38122];
assign t[38123] = t[38122] ^ n[38123];
assign t[38124] = t[38123] ^ n[38124];
assign t[38125] = t[38124] ^ n[38125];
assign t[38126] = t[38125] ^ n[38126];
assign t[38127] = t[38126] ^ n[38127];
assign t[38128] = t[38127] ^ n[38128];
assign t[38129] = t[38128] ^ n[38129];
assign t[38130] = t[38129] ^ n[38130];
assign t[38131] = t[38130] ^ n[38131];
assign t[38132] = t[38131] ^ n[38132];
assign t[38133] = t[38132] ^ n[38133];
assign t[38134] = t[38133] ^ n[38134];
assign t[38135] = t[38134] ^ n[38135];
assign t[38136] = t[38135] ^ n[38136];
assign t[38137] = t[38136] ^ n[38137];
assign t[38138] = t[38137] ^ n[38138];
assign t[38139] = t[38138] ^ n[38139];
assign t[38140] = t[38139] ^ n[38140];
assign t[38141] = t[38140] ^ n[38141];
assign t[38142] = t[38141] ^ n[38142];
assign t[38143] = t[38142] ^ n[38143];
assign t[38144] = t[38143] ^ n[38144];
assign t[38145] = t[38144] ^ n[38145];
assign t[38146] = t[38145] ^ n[38146];
assign t[38147] = t[38146] ^ n[38147];
assign t[38148] = t[38147] ^ n[38148];
assign t[38149] = t[38148] ^ n[38149];
assign t[38150] = t[38149] ^ n[38150];
assign t[38151] = t[38150] ^ n[38151];
assign t[38152] = t[38151] ^ n[38152];
assign t[38153] = t[38152] ^ n[38153];
assign t[38154] = t[38153] ^ n[38154];
assign t[38155] = t[38154] ^ n[38155];
assign t[38156] = t[38155] ^ n[38156];
assign t[38157] = t[38156] ^ n[38157];
assign t[38158] = t[38157] ^ n[38158];
assign t[38159] = t[38158] ^ n[38159];
assign t[38160] = t[38159] ^ n[38160];
assign t[38161] = t[38160] ^ n[38161];
assign t[38162] = t[38161] ^ n[38162];
assign t[38163] = t[38162] ^ n[38163];
assign t[38164] = t[38163] ^ n[38164];
assign t[38165] = t[38164] ^ n[38165];
assign t[38166] = t[38165] ^ n[38166];
assign t[38167] = t[38166] ^ n[38167];
assign t[38168] = t[38167] ^ n[38168];
assign t[38169] = t[38168] ^ n[38169];
assign t[38170] = t[38169] ^ n[38170];
assign t[38171] = t[38170] ^ n[38171];
assign t[38172] = t[38171] ^ n[38172];
assign t[38173] = t[38172] ^ n[38173];
assign t[38174] = t[38173] ^ n[38174];
assign t[38175] = t[38174] ^ n[38175];
assign t[38176] = t[38175] ^ n[38176];
assign t[38177] = t[38176] ^ n[38177];
assign t[38178] = t[38177] ^ n[38178];
assign t[38179] = t[38178] ^ n[38179];
assign t[38180] = t[38179] ^ n[38180];
assign t[38181] = t[38180] ^ n[38181];
assign t[38182] = t[38181] ^ n[38182];
assign t[38183] = t[38182] ^ n[38183];
assign t[38184] = t[38183] ^ n[38184];
assign t[38185] = t[38184] ^ n[38185];
assign t[38186] = t[38185] ^ n[38186];
assign t[38187] = t[38186] ^ n[38187];
assign t[38188] = t[38187] ^ n[38188];
assign t[38189] = t[38188] ^ n[38189];
assign t[38190] = t[38189] ^ n[38190];
assign t[38191] = t[38190] ^ n[38191];
assign t[38192] = t[38191] ^ n[38192];
assign t[38193] = t[38192] ^ n[38193];
assign t[38194] = t[38193] ^ n[38194];
assign t[38195] = t[38194] ^ n[38195];
assign t[38196] = t[38195] ^ n[38196];
assign t[38197] = t[38196] ^ n[38197];
assign t[38198] = t[38197] ^ n[38198];
assign t[38199] = t[38198] ^ n[38199];
assign t[38200] = t[38199] ^ n[38200];
assign t[38201] = t[38200] ^ n[38201];
assign t[38202] = t[38201] ^ n[38202];
assign t[38203] = t[38202] ^ n[38203];
assign t[38204] = t[38203] ^ n[38204];
assign t[38205] = t[38204] ^ n[38205];
assign t[38206] = t[38205] ^ n[38206];
assign t[38207] = t[38206] ^ n[38207];
assign t[38208] = t[38207] ^ n[38208];
assign t[38209] = t[38208] ^ n[38209];
assign t[38210] = t[38209] ^ n[38210];
assign t[38211] = t[38210] ^ n[38211];
assign t[38212] = t[38211] ^ n[38212];
assign t[38213] = t[38212] ^ n[38213];
assign t[38214] = t[38213] ^ n[38214];
assign t[38215] = t[38214] ^ n[38215];
assign t[38216] = t[38215] ^ n[38216];
assign t[38217] = t[38216] ^ n[38217];
assign t[38218] = t[38217] ^ n[38218];
assign t[38219] = t[38218] ^ n[38219];
assign t[38220] = t[38219] ^ n[38220];
assign t[38221] = t[38220] ^ n[38221];
assign t[38222] = t[38221] ^ n[38222];
assign t[38223] = t[38222] ^ n[38223];
assign t[38224] = t[38223] ^ n[38224];
assign t[38225] = t[38224] ^ n[38225];
assign t[38226] = t[38225] ^ n[38226];
assign t[38227] = t[38226] ^ n[38227];
assign t[38228] = t[38227] ^ n[38228];
assign t[38229] = t[38228] ^ n[38229];
assign t[38230] = t[38229] ^ n[38230];
assign t[38231] = t[38230] ^ n[38231];
assign t[38232] = t[38231] ^ n[38232];
assign t[38233] = t[38232] ^ n[38233];
assign t[38234] = t[38233] ^ n[38234];
assign t[38235] = t[38234] ^ n[38235];
assign t[38236] = t[38235] ^ n[38236];
assign t[38237] = t[38236] ^ n[38237];
assign t[38238] = t[38237] ^ n[38238];
assign t[38239] = t[38238] ^ n[38239];
assign t[38240] = t[38239] ^ n[38240];
assign t[38241] = t[38240] ^ n[38241];
assign t[38242] = t[38241] ^ n[38242];
assign t[38243] = t[38242] ^ n[38243];
assign t[38244] = t[38243] ^ n[38244];
assign t[38245] = t[38244] ^ n[38245];
assign t[38246] = t[38245] ^ n[38246];
assign t[38247] = t[38246] ^ n[38247];
assign t[38248] = t[38247] ^ n[38248];
assign t[38249] = t[38248] ^ n[38249];
assign t[38250] = t[38249] ^ n[38250];
assign t[38251] = t[38250] ^ n[38251];
assign t[38252] = t[38251] ^ n[38252];
assign t[38253] = t[38252] ^ n[38253];
assign t[38254] = t[38253] ^ n[38254];
assign t[38255] = t[38254] ^ n[38255];
assign t[38256] = t[38255] ^ n[38256];
assign t[38257] = t[38256] ^ n[38257];
assign t[38258] = t[38257] ^ n[38258];
assign t[38259] = t[38258] ^ n[38259];
assign t[38260] = t[38259] ^ n[38260];
assign t[38261] = t[38260] ^ n[38261];
assign t[38262] = t[38261] ^ n[38262];
assign t[38263] = t[38262] ^ n[38263];
assign t[38264] = t[38263] ^ n[38264];
assign t[38265] = t[38264] ^ n[38265];
assign t[38266] = t[38265] ^ n[38266];
assign t[38267] = t[38266] ^ n[38267];
assign t[38268] = t[38267] ^ n[38268];
assign t[38269] = t[38268] ^ n[38269];
assign t[38270] = t[38269] ^ n[38270];
assign t[38271] = t[38270] ^ n[38271];
assign t[38272] = t[38271] ^ n[38272];
assign t[38273] = t[38272] ^ n[38273];
assign t[38274] = t[38273] ^ n[38274];
assign t[38275] = t[38274] ^ n[38275];
assign t[38276] = t[38275] ^ n[38276];
assign t[38277] = t[38276] ^ n[38277];
assign t[38278] = t[38277] ^ n[38278];
assign t[38279] = t[38278] ^ n[38279];
assign t[38280] = t[38279] ^ n[38280];
assign t[38281] = t[38280] ^ n[38281];
assign t[38282] = t[38281] ^ n[38282];
assign t[38283] = t[38282] ^ n[38283];
assign t[38284] = t[38283] ^ n[38284];
assign t[38285] = t[38284] ^ n[38285];
assign t[38286] = t[38285] ^ n[38286];
assign t[38287] = t[38286] ^ n[38287];
assign t[38288] = t[38287] ^ n[38288];
assign t[38289] = t[38288] ^ n[38289];
assign t[38290] = t[38289] ^ n[38290];
assign t[38291] = t[38290] ^ n[38291];
assign t[38292] = t[38291] ^ n[38292];
assign t[38293] = t[38292] ^ n[38293];
assign t[38294] = t[38293] ^ n[38294];
assign t[38295] = t[38294] ^ n[38295];
assign t[38296] = t[38295] ^ n[38296];
assign t[38297] = t[38296] ^ n[38297];
assign t[38298] = t[38297] ^ n[38298];
assign t[38299] = t[38298] ^ n[38299];
assign t[38300] = t[38299] ^ n[38300];
assign t[38301] = t[38300] ^ n[38301];
assign t[38302] = t[38301] ^ n[38302];
assign t[38303] = t[38302] ^ n[38303];
assign t[38304] = t[38303] ^ n[38304];
assign t[38305] = t[38304] ^ n[38305];
assign t[38306] = t[38305] ^ n[38306];
assign t[38307] = t[38306] ^ n[38307];
assign t[38308] = t[38307] ^ n[38308];
assign t[38309] = t[38308] ^ n[38309];
assign t[38310] = t[38309] ^ n[38310];
assign t[38311] = t[38310] ^ n[38311];
assign t[38312] = t[38311] ^ n[38312];
assign t[38313] = t[38312] ^ n[38313];
assign t[38314] = t[38313] ^ n[38314];
assign t[38315] = t[38314] ^ n[38315];
assign t[38316] = t[38315] ^ n[38316];
assign t[38317] = t[38316] ^ n[38317];
assign t[38318] = t[38317] ^ n[38318];
assign t[38319] = t[38318] ^ n[38319];
assign t[38320] = t[38319] ^ n[38320];
assign t[38321] = t[38320] ^ n[38321];
assign t[38322] = t[38321] ^ n[38322];
assign t[38323] = t[38322] ^ n[38323];
assign t[38324] = t[38323] ^ n[38324];
assign t[38325] = t[38324] ^ n[38325];
assign t[38326] = t[38325] ^ n[38326];
assign t[38327] = t[38326] ^ n[38327];
assign t[38328] = t[38327] ^ n[38328];
assign t[38329] = t[38328] ^ n[38329];
assign t[38330] = t[38329] ^ n[38330];
assign t[38331] = t[38330] ^ n[38331];
assign t[38332] = t[38331] ^ n[38332];
assign t[38333] = t[38332] ^ n[38333];
assign t[38334] = t[38333] ^ n[38334];
assign t[38335] = t[38334] ^ n[38335];
assign t[38336] = t[38335] ^ n[38336];
assign t[38337] = t[38336] ^ n[38337];
assign t[38338] = t[38337] ^ n[38338];
assign t[38339] = t[38338] ^ n[38339];
assign t[38340] = t[38339] ^ n[38340];
assign t[38341] = t[38340] ^ n[38341];
assign t[38342] = t[38341] ^ n[38342];
assign t[38343] = t[38342] ^ n[38343];
assign t[38344] = t[38343] ^ n[38344];
assign t[38345] = t[38344] ^ n[38345];
assign t[38346] = t[38345] ^ n[38346];
assign t[38347] = t[38346] ^ n[38347];
assign t[38348] = t[38347] ^ n[38348];
assign t[38349] = t[38348] ^ n[38349];
assign t[38350] = t[38349] ^ n[38350];
assign t[38351] = t[38350] ^ n[38351];
assign t[38352] = t[38351] ^ n[38352];
assign t[38353] = t[38352] ^ n[38353];
assign t[38354] = t[38353] ^ n[38354];
assign t[38355] = t[38354] ^ n[38355];
assign t[38356] = t[38355] ^ n[38356];
assign t[38357] = t[38356] ^ n[38357];
assign t[38358] = t[38357] ^ n[38358];
assign t[38359] = t[38358] ^ n[38359];
assign t[38360] = t[38359] ^ n[38360];
assign t[38361] = t[38360] ^ n[38361];
assign t[38362] = t[38361] ^ n[38362];
assign t[38363] = t[38362] ^ n[38363];
assign t[38364] = t[38363] ^ n[38364];
assign t[38365] = t[38364] ^ n[38365];
assign t[38366] = t[38365] ^ n[38366];
assign t[38367] = t[38366] ^ n[38367];
assign t[38368] = t[38367] ^ n[38368];
assign t[38369] = t[38368] ^ n[38369];
assign t[38370] = t[38369] ^ n[38370];
assign t[38371] = t[38370] ^ n[38371];
assign t[38372] = t[38371] ^ n[38372];
assign t[38373] = t[38372] ^ n[38373];
assign t[38374] = t[38373] ^ n[38374];
assign t[38375] = t[38374] ^ n[38375];
assign t[38376] = t[38375] ^ n[38376];
assign t[38377] = t[38376] ^ n[38377];
assign t[38378] = t[38377] ^ n[38378];
assign t[38379] = t[38378] ^ n[38379];
assign t[38380] = t[38379] ^ n[38380];
assign t[38381] = t[38380] ^ n[38381];
assign t[38382] = t[38381] ^ n[38382];
assign t[38383] = t[38382] ^ n[38383];
assign t[38384] = t[38383] ^ n[38384];
assign t[38385] = t[38384] ^ n[38385];
assign t[38386] = t[38385] ^ n[38386];
assign t[38387] = t[38386] ^ n[38387];
assign t[38388] = t[38387] ^ n[38388];
assign t[38389] = t[38388] ^ n[38389];
assign t[38390] = t[38389] ^ n[38390];
assign t[38391] = t[38390] ^ n[38391];
assign t[38392] = t[38391] ^ n[38392];
assign t[38393] = t[38392] ^ n[38393];
assign t[38394] = t[38393] ^ n[38394];
assign t[38395] = t[38394] ^ n[38395];
assign t[38396] = t[38395] ^ n[38396];
assign t[38397] = t[38396] ^ n[38397];
assign t[38398] = t[38397] ^ n[38398];
assign t[38399] = t[38398] ^ n[38399];
assign t[38400] = t[38399] ^ n[38400];
assign t[38401] = t[38400] ^ n[38401];
assign t[38402] = t[38401] ^ n[38402];
assign t[38403] = t[38402] ^ n[38403];
assign t[38404] = t[38403] ^ n[38404];
assign t[38405] = t[38404] ^ n[38405];
assign t[38406] = t[38405] ^ n[38406];
assign t[38407] = t[38406] ^ n[38407];
assign t[38408] = t[38407] ^ n[38408];
assign t[38409] = t[38408] ^ n[38409];
assign t[38410] = t[38409] ^ n[38410];
assign t[38411] = t[38410] ^ n[38411];
assign t[38412] = t[38411] ^ n[38412];
assign t[38413] = t[38412] ^ n[38413];
assign t[38414] = t[38413] ^ n[38414];
assign t[38415] = t[38414] ^ n[38415];
assign t[38416] = t[38415] ^ n[38416];
assign t[38417] = t[38416] ^ n[38417];
assign t[38418] = t[38417] ^ n[38418];
assign t[38419] = t[38418] ^ n[38419];
assign t[38420] = t[38419] ^ n[38420];
assign t[38421] = t[38420] ^ n[38421];
assign t[38422] = t[38421] ^ n[38422];
assign t[38423] = t[38422] ^ n[38423];
assign t[38424] = t[38423] ^ n[38424];
assign t[38425] = t[38424] ^ n[38425];
assign t[38426] = t[38425] ^ n[38426];
assign t[38427] = t[38426] ^ n[38427];
assign t[38428] = t[38427] ^ n[38428];
assign t[38429] = t[38428] ^ n[38429];
assign t[38430] = t[38429] ^ n[38430];
assign t[38431] = t[38430] ^ n[38431];
assign t[38432] = t[38431] ^ n[38432];
assign t[38433] = t[38432] ^ n[38433];
assign t[38434] = t[38433] ^ n[38434];
assign t[38435] = t[38434] ^ n[38435];
assign t[38436] = t[38435] ^ n[38436];
assign t[38437] = t[38436] ^ n[38437];
assign t[38438] = t[38437] ^ n[38438];
assign t[38439] = t[38438] ^ n[38439];
assign t[38440] = t[38439] ^ n[38440];
assign t[38441] = t[38440] ^ n[38441];
assign t[38442] = t[38441] ^ n[38442];
assign t[38443] = t[38442] ^ n[38443];
assign t[38444] = t[38443] ^ n[38444];
assign t[38445] = t[38444] ^ n[38445];
assign t[38446] = t[38445] ^ n[38446];
assign t[38447] = t[38446] ^ n[38447];
assign t[38448] = t[38447] ^ n[38448];
assign t[38449] = t[38448] ^ n[38449];
assign t[38450] = t[38449] ^ n[38450];
assign t[38451] = t[38450] ^ n[38451];
assign t[38452] = t[38451] ^ n[38452];
assign t[38453] = t[38452] ^ n[38453];
assign t[38454] = t[38453] ^ n[38454];
assign t[38455] = t[38454] ^ n[38455];
assign t[38456] = t[38455] ^ n[38456];
assign t[38457] = t[38456] ^ n[38457];
assign t[38458] = t[38457] ^ n[38458];
assign t[38459] = t[38458] ^ n[38459];
assign t[38460] = t[38459] ^ n[38460];
assign t[38461] = t[38460] ^ n[38461];
assign t[38462] = t[38461] ^ n[38462];
assign t[38463] = t[38462] ^ n[38463];
assign t[38464] = t[38463] ^ n[38464];
assign t[38465] = t[38464] ^ n[38465];
assign t[38466] = t[38465] ^ n[38466];
assign t[38467] = t[38466] ^ n[38467];
assign t[38468] = t[38467] ^ n[38468];
assign t[38469] = t[38468] ^ n[38469];
assign t[38470] = t[38469] ^ n[38470];
assign t[38471] = t[38470] ^ n[38471];
assign t[38472] = t[38471] ^ n[38472];
assign t[38473] = t[38472] ^ n[38473];
assign t[38474] = t[38473] ^ n[38474];
assign t[38475] = t[38474] ^ n[38475];
assign t[38476] = t[38475] ^ n[38476];
assign t[38477] = t[38476] ^ n[38477];
assign t[38478] = t[38477] ^ n[38478];
assign t[38479] = t[38478] ^ n[38479];
assign t[38480] = t[38479] ^ n[38480];
assign t[38481] = t[38480] ^ n[38481];
assign t[38482] = t[38481] ^ n[38482];
assign t[38483] = t[38482] ^ n[38483];
assign t[38484] = t[38483] ^ n[38484];
assign t[38485] = t[38484] ^ n[38485];
assign t[38486] = t[38485] ^ n[38486];
assign t[38487] = t[38486] ^ n[38487];
assign t[38488] = t[38487] ^ n[38488];
assign t[38489] = t[38488] ^ n[38489];
assign t[38490] = t[38489] ^ n[38490];
assign t[38491] = t[38490] ^ n[38491];
assign t[38492] = t[38491] ^ n[38492];
assign t[38493] = t[38492] ^ n[38493];
assign t[38494] = t[38493] ^ n[38494];
assign t[38495] = t[38494] ^ n[38495];
assign t[38496] = t[38495] ^ n[38496];
assign t[38497] = t[38496] ^ n[38497];
assign t[38498] = t[38497] ^ n[38498];
assign t[38499] = t[38498] ^ n[38499];
assign t[38500] = t[38499] ^ n[38500];
assign t[38501] = t[38500] ^ n[38501];
assign t[38502] = t[38501] ^ n[38502];
assign t[38503] = t[38502] ^ n[38503];
assign t[38504] = t[38503] ^ n[38504];
assign t[38505] = t[38504] ^ n[38505];
assign t[38506] = t[38505] ^ n[38506];
assign t[38507] = t[38506] ^ n[38507];
assign t[38508] = t[38507] ^ n[38508];
assign t[38509] = t[38508] ^ n[38509];
assign t[38510] = t[38509] ^ n[38510];
assign t[38511] = t[38510] ^ n[38511];
assign t[38512] = t[38511] ^ n[38512];
assign t[38513] = t[38512] ^ n[38513];
assign t[38514] = t[38513] ^ n[38514];
assign t[38515] = t[38514] ^ n[38515];
assign t[38516] = t[38515] ^ n[38516];
assign t[38517] = t[38516] ^ n[38517];
assign t[38518] = t[38517] ^ n[38518];
assign t[38519] = t[38518] ^ n[38519];
assign t[38520] = t[38519] ^ n[38520];
assign t[38521] = t[38520] ^ n[38521];
assign t[38522] = t[38521] ^ n[38522];
assign t[38523] = t[38522] ^ n[38523];
assign t[38524] = t[38523] ^ n[38524];
assign t[38525] = t[38524] ^ n[38525];
assign t[38526] = t[38525] ^ n[38526];
assign t[38527] = t[38526] ^ n[38527];
assign t[38528] = t[38527] ^ n[38528];
assign t[38529] = t[38528] ^ n[38529];
assign t[38530] = t[38529] ^ n[38530];
assign t[38531] = t[38530] ^ n[38531];
assign t[38532] = t[38531] ^ n[38532];
assign t[38533] = t[38532] ^ n[38533];
assign t[38534] = t[38533] ^ n[38534];
assign t[38535] = t[38534] ^ n[38535];
assign t[38536] = t[38535] ^ n[38536];
assign t[38537] = t[38536] ^ n[38537];
assign t[38538] = t[38537] ^ n[38538];
assign t[38539] = t[38538] ^ n[38539];
assign t[38540] = t[38539] ^ n[38540];
assign t[38541] = t[38540] ^ n[38541];
assign t[38542] = t[38541] ^ n[38542];
assign t[38543] = t[38542] ^ n[38543];
assign t[38544] = t[38543] ^ n[38544];
assign t[38545] = t[38544] ^ n[38545];
assign t[38546] = t[38545] ^ n[38546];
assign t[38547] = t[38546] ^ n[38547];
assign t[38548] = t[38547] ^ n[38548];
assign t[38549] = t[38548] ^ n[38549];
assign t[38550] = t[38549] ^ n[38550];
assign t[38551] = t[38550] ^ n[38551];
assign t[38552] = t[38551] ^ n[38552];
assign t[38553] = t[38552] ^ n[38553];
assign t[38554] = t[38553] ^ n[38554];
assign t[38555] = t[38554] ^ n[38555];
assign t[38556] = t[38555] ^ n[38556];
assign t[38557] = t[38556] ^ n[38557];
assign t[38558] = t[38557] ^ n[38558];
assign t[38559] = t[38558] ^ n[38559];
assign t[38560] = t[38559] ^ n[38560];
assign t[38561] = t[38560] ^ n[38561];
assign t[38562] = t[38561] ^ n[38562];
assign t[38563] = t[38562] ^ n[38563];
assign t[38564] = t[38563] ^ n[38564];
assign t[38565] = t[38564] ^ n[38565];
assign t[38566] = t[38565] ^ n[38566];
assign t[38567] = t[38566] ^ n[38567];
assign t[38568] = t[38567] ^ n[38568];
assign t[38569] = t[38568] ^ n[38569];
assign t[38570] = t[38569] ^ n[38570];
assign t[38571] = t[38570] ^ n[38571];
assign t[38572] = t[38571] ^ n[38572];
assign t[38573] = t[38572] ^ n[38573];
assign t[38574] = t[38573] ^ n[38574];
assign t[38575] = t[38574] ^ n[38575];
assign t[38576] = t[38575] ^ n[38576];
assign t[38577] = t[38576] ^ n[38577];
assign t[38578] = t[38577] ^ n[38578];
assign t[38579] = t[38578] ^ n[38579];
assign t[38580] = t[38579] ^ n[38580];
assign t[38581] = t[38580] ^ n[38581];
assign t[38582] = t[38581] ^ n[38582];
assign t[38583] = t[38582] ^ n[38583];
assign t[38584] = t[38583] ^ n[38584];
assign t[38585] = t[38584] ^ n[38585];
assign t[38586] = t[38585] ^ n[38586];
assign t[38587] = t[38586] ^ n[38587];
assign t[38588] = t[38587] ^ n[38588];
assign t[38589] = t[38588] ^ n[38589];
assign t[38590] = t[38589] ^ n[38590];
assign t[38591] = t[38590] ^ n[38591];
assign t[38592] = t[38591] ^ n[38592];
assign t[38593] = t[38592] ^ n[38593];
assign t[38594] = t[38593] ^ n[38594];
assign t[38595] = t[38594] ^ n[38595];
assign t[38596] = t[38595] ^ n[38596];
assign t[38597] = t[38596] ^ n[38597];
assign t[38598] = t[38597] ^ n[38598];
assign t[38599] = t[38598] ^ n[38599];
assign t[38600] = t[38599] ^ n[38600];
assign t[38601] = t[38600] ^ n[38601];
assign t[38602] = t[38601] ^ n[38602];
assign t[38603] = t[38602] ^ n[38603];
assign t[38604] = t[38603] ^ n[38604];
assign t[38605] = t[38604] ^ n[38605];
assign t[38606] = t[38605] ^ n[38606];
assign t[38607] = t[38606] ^ n[38607];
assign t[38608] = t[38607] ^ n[38608];
assign t[38609] = t[38608] ^ n[38609];
assign t[38610] = t[38609] ^ n[38610];
assign t[38611] = t[38610] ^ n[38611];
assign t[38612] = t[38611] ^ n[38612];
assign t[38613] = t[38612] ^ n[38613];
assign t[38614] = t[38613] ^ n[38614];
assign t[38615] = t[38614] ^ n[38615];
assign t[38616] = t[38615] ^ n[38616];
assign t[38617] = t[38616] ^ n[38617];
assign t[38618] = t[38617] ^ n[38618];
assign t[38619] = t[38618] ^ n[38619];
assign t[38620] = t[38619] ^ n[38620];
assign t[38621] = t[38620] ^ n[38621];
assign t[38622] = t[38621] ^ n[38622];
assign t[38623] = t[38622] ^ n[38623];
assign t[38624] = t[38623] ^ n[38624];
assign t[38625] = t[38624] ^ n[38625];
assign t[38626] = t[38625] ^ n[38626];
assign t[38627] = t[38626] ^ n[38627];
assign t[38628] = t[38627] ^ n[38628];
assign t[38629] = t[38628] ^ n[38629];
assign t[38630] = t[38629] ^ n[38630];
assign t[38631] = t[38630] ^ n[38631];
assign t[38632] = t[38631] ^ n[38632];
assign t[38633] = t[38632] ^ n[38633];
assign t[38634] = t[38633] ^ n[38634];
assign t[38635] = t[38634] ^ n[38635];
assign t[38636] = t[38635] ^ n[38636];
assign t[38637] = t[38636] ^ n[38637];
assign t[38638] = t[38637] ^ n[38638];
assign t[38639] = t[38638] ^ n[38639];
assign t[38640] = t[38639] ^ n[38640];
assign t[38641] = t[38640] ^ n[38641];
assign t[38642] = t[38641] ^ n[38642];
assign t[38643] = t[38642] ^ n[38643];
assign t[38644] = t[38643] ^ n[38644];
assign t[38645] = t[38644] ^ n[38645];
assign t[38646] = t[38645] ^ n[38646];
assign t[38647] = t[38646] ^ n[38647];
assign t[38648] = t[38647] ^ n[38648];
assign t[38649] = t[38648] ^ n[38649];
assign t[38650] = t[38649] ^ n[38650];
assign t[38651] = t[38650] ^ n[38651];
assign t[38652] = t[38651] ^ n[38652];
assign t[38653] = t[38652] ^ n[38653];
assign t[38654] = t[38653] ^ n[38654];
assign t[38655] = t[38654] ^ n[38655];
assign t[38656] = t[38655] ^ n[38656];
assign t[38657] = t[38656] ^ n[38657];
assign t[38658] = t[38657] ^ n[38658];
assign t[38659] = t[38658] ^ n[38659];
assign t[38660] = t[38659] ^ n[38660];
assign t[38661] = t[38660] ^ n[38661];
assign t[38662] = t[38661] ^ n[38662];
assign t[38663] = t[38662] ^ n[38663];
assign t[38664] = t[38663] ^ n[38664];
assign t[38665] = t[38664] ^ n[38665];
assign t[38666] = t[38665] ^ n[38666];
assign t[38667] = t[38666] ^ n[38667];
assign t[38668] = t[38667] ^ n[38668];
assign t[38669] = t[38668] ^ n[38669];
assign t[38670] = t[38669] ^ n[38670];
assign t[38671] = t[38670] ^ n[38671];
assign t[38672] = t[38671] ^ n[38672];
assign t[38673] = t[38672] ^ n[38673];
assign t[38674] = t[38673] ^ n[38674];
assign t[38675] = t[38674] ^ n[38675];
assign t[38676] = t[38675] ^ n[38676];
assign t[38677] = t[38676] ^ n[38677];
assign t[38678] = t[38677] ^ n[38678];
assign t[38679] = t[38678] ^ n[38679];
assign t[38680] = t[38679] ^ n[38680];
assign t[38681] = t[38680] ^ n[38681];
assign t[38682] = t[38681] ^ n[38682];
assign t[38683] = t[38682] ^ n[38683];
assign t[38684] = t[38683] ^ n[38684];
assign t[38685] = t[38684] ^ n[38685];
assign t[38686] = t[38685] ^ n[38686];
assign t[38687] = t[38686] ^ n[38687];
assign t[38688] = t[38687] ^ n[38688];
assign t[38689] = t[38688] ^ n[38689];
assign t[38690] = t[38689] ^ n[38690];
assign t[38691] = t[38690] ^ n[38691];
assign t[38692] = t[38691] ^ n[38692];
assign t[38693] = t[38692] ^ n[38693];
assign t[38694] = t[38693] ^ n[38694];
assign t[38695] = t[38694] ^ n[38695];
assign t[38696] = t[38695] ^ n[38696];
assign t[38697] = t[38696] ^ n[38697];
assign t[38698] = t[38697] ^ n[38698];
assign t[38699] = t[38698] ^ n[38699];
assign t[38700] = t[38699] ^ n[38700];
assign t[38701] = t[38700] ^ n[38701];
assign t[38702] = t[38701] ^ n[38702];
assign t[38703] = t[38702] ^ n[38703];
assign t[38704] = t[38703] ^ n[38704];
assign t[38705] = t[38704] ^ n[38705];
assign t[38706] = t[38705] ^ n[38706];
assign t[38707] = t[38706] ^ n[38707];
assign t[38708] = t[38707] ^ n[38708];
assign t[38709] = t[38708] ^ n[38709];
assign t[38710] = t[38709] ^ n[38710];
assign t[38711] = t[38710] ^ n[38711];
assign t[38712] = t[38711] ^ n[38712];
assign t[38713] = t[38712] ^ n[38713];
assign t[38714] = t[38713] ^ n[38714];
assign t[38715] = t[38714] ^ n[38715];
assign t[38716] = t[38715] ^ n[38716];
assign t[38717] = t[38716] ^ n[38717];
assign t[38718] = t[38717] ^ n[38718];
assign t[38719] = t[38718] ^ n[38719];
assign t[38720] = t[38719] ^ n[38720];
assign t[38721] = t[38720] ^ n[38721];
assign t[38722] = t[38721] ^ n[38722];
assign t[38723] = t[38722] ^ n[38723];
assign t[38724] = t[38723] ^ n[38724];
assign t[38725] = t[38724] ^ n[38725];
assign t[38726] = t[38725] ^ n[38726];
assign t[38727] = t[38726] ^ n[38727];
assign t[38728] = t[38727] ^ n[38728];
assign t[38729] = t[38728] ^ n[38729];
assign t[38730] = t[38729] ^ n[38730];
assign t[38731] = t[38730] ^ n[38731];
assign t[38732] = t[38731] ^ n[38732];
assign t[38733] = t[38732] ^ n[38733];
assign t[38734] = t[38733] ^ n[38734];
assign t[38735] = t[38734] ^ n[38735];
assign t[38736] = t[38735] ^ n[38736];
assign t[38737] = t[38736] ^ n[38737];
assign t[38738] = t[38737] ^ n[38738];
assign t[38739] = t[38738] ^ n[38739];
assign t[38740] = t[38739] ^ n[38740];
assign t[38741] = t[38740] ^ n[38741];
assign t[38742] = t[38741] ^ n[38742];
assign t[38743] = t[38742] ^ n[38743];
assign t[38744] = t[38743] ^ n[38744];
assign t[38745] = t[38744] ^ n[38745];
assign t[38746] = t[38745] ^ n[38746];
assign t[38747] = t[38746] ^ n[38747];
assign t[38748] = t[38747] ^ n[38748];
assign t[38749] = t[38748] ^ n[38749];
assign t[38750] = t[38749] ^ n[38750];
assign t[38751] = t[38750] ^ n[38751];
assign t[38752] = t[38751] ^ n[38752];
assign t[38753] = t[38752] ^ n[38753];
assign t[38754] = t[38753] ^ n[38754];
assign t[38755] = t[38754] ^ n[38755];
assign t[38756] = t[38755] ^ n[38756];
assign t[38757] = t[38756] ^ n[38757];
assign t[38758] = t[38757] ^ n[38758];
assign t[38759] = t[38758] ^ n[38759];
assign t[38760] = t[38759] ^ n[38760];
assign t[38761] = t[38760] ^ n[38761];
assign t[38762] = t[38761] ^ n[38762];
assign t[38763] = t[38762] ^ n[38763];
assign t[38764] = t[38763] ^ n[38764];
assign t[38765] = t[38764] ^ n[38765];
assign t[38766] = t[38765] ^ n[38766];
assign t[38767] = t[38766] ^ n[38767];
assign t[38768] = t[38767] ^ n[38768];
assign t[38769] = t[38768] ^ n[38769];
assign t[38770] = t[38769] ^ n[38770];
assign t[38771] = t[38770] ^ n[38771];
assign t[38772] = t[38771] ^ n[38772];
assign t[38773] = t[38772] ^ n[38773];
assign t[38774] = t[38773] ^ n[38774];
assign t[38775] = t[38774] ^ n[38775];
assign t[38776] = t[38775] ^ n[38776];
assign t[38777] = t[38776] ^ n[38777];
assign t[38778] = t[38777] ^ n[38778];
assign t[38779] = t[38778] ^ n[38779];
assign t[38780] = t[38779] ^ n[38780];
assign t[38781] = t[38780] ^ n[38781];
assign t[38782] = t[38781] ^ n[38782];
assign t[38783] = t[38782] ^ n[38783];
assign t[38784] = t[38783] ^ n[38784];
assign t[38785] = t[38784] ^ n[38785];
assign t[38786] = t[38785] ^ n[38786];
assign t[38787] = t[38786] ^ n[38787];
assign t[38788] = t[38787] ^ n[38788];
assign t[38789] = t[38788] ^ n[38789];
assign t[38790] = t[38789] ^ n[38790];
assign t[38791] = t[38790] ^ n[38791];
assign t[38792] = t[38791] ^ n[38792];
assign t[38793] = t[38792] ^ n[38793];
assign t[38794] = t[38793] ^ n[38794];
assign t[38795] = t[38794] ^ n[38795];
assign t[38796] = t[38795] ^ n[38796];
assign t[38797] = t[38796] ^ n[38797];
assign t[38798] = t[38797] ^ n[38798];
assign t[38799] = t[38798] ^ n[38799];
assign t[38800] = t[38799] ^ n[38800];
assign t[38801] = t[38800] ^ n[38801];
assign t[38802] = t[38801] ^ n[38802];
assign t[38803] = t[38802] ^ n[38803];
assign t[38804] = t[38803] ^ n[38804];
assign t[38805] = t[38804] ^ n[38805];
assign t[38806] = t[38805] ^ n[38806];
assign t[38807] = t[38806] ^ n[38807];
assign t[38808] = t[38807] ^ n[38808];
assign t[38809] = t[38808] ^ n[38809];
assign t[38810] = t[38809] ^ n[38810];
assign t[38811] = t[38810] ^ n[38811];
assign t[38812] = t[38811] ^ n[38812];
assign t[38813] = t[38812] ^ n[38813];
assign t[38814] = t[38813] ^ n[38814];
assign t[38815] = t[38814] ^ n[38815];
assign t[38816] = t[38815] ^ n[38816];
assign t[38817] = t[38816] ^ n[38817];
assign t[38818] = t[38817] ^ n[38818];
assign t[38819] = t[38818] ^ n[38819];
assign t[38820] = t[38819] ^ n[38820];
assign t[38821] = t[38820] ^ n[38821];
assign t[38822] = t[38821] ^ n[38822];
assign t[38823] = t[38822] ^ n[38823];
assign t[38824] = t[38823] ^ n[38824];
assign t[38825] = t[38824] ^ n[38825];
assign t[38826] = t[38825] ^ n[38826];
assign t[38827] = t[38826] ^ n[38827];
assign t[38828] = t[38827] ^ n[38828];
assign t[38829] = t[38828] ^ n[38829];
assign t[38830] = t[38829] ^ n[38830];
assign t[38831] = t[38830] ^ n[38831];
assign t[38832] = t[38831] ^ n[38832];
assign t[38833] = t[38832] ^ n[38833];
assign t[38834] = t[38833] ^ n[38834];
assign t[38835] = t[38834] ^ n[38835];
assign t[38836] = t[38835] ^ n[38836];
assign t[38837] = t[38836] ^ n[38837];
assign t[38838] = t[38837] ^ n[38838];
assign t[38839] = t[38838] ^ n[38839];
assign t[38840] = t[38839] ^ n[38840];
assign t[38841] = t[38840] ^ n[38841];
assign t[38842] = t[38841] ^ n[38842];
assign t[38843] = t[38842] ^ n[38843];
assign t[38844] = t[38843] ^ n[38844];
assign t[38845] = t[38844] ^ n[38845];
assign t[38846] = t[38845] ^ n[38846];
assign t[38847] = t[38846] ^ n[38847];
assign t[38848] = t[38847] ^ n[38848];
assign t[38849] = t[38848] ^ n[38849];
assign t[38850] = t[38849] ^ n[38850];
assign t[38851] = t[38850] ^ n[38851];
assign t[38852] = t[38851] ^ n[38852];
assign t[38853] = t[38852] ^ n[38853];
assign t[38854] = t[38853] ^ n[38854];
assign t[38855] = t[38854] ^ n[38855];
assign t[38856] = t[38855] ^ n[38856];
assign t[38857] = t[38856] ^ n[38857];
assign t[38858] = t[38857] ^ n[38858];
assign t[38859] = t[38858] ^ n[38859];
assign t[38860] = t[38859] ^ n[38860];
assign t[38861] = t[38860] ^ n[38861];
assign t[38862] = t[38861] ^ n[38862];
assign t[38863] = t[38862] ^ n[38863];
assign t[38864] = t[38863] ^ n[38864];
assign t[38865] = t[38864] ^ n[38865];
assign t[38866] = t[38865] ^ n[38866];
assign t[38867] = t[38866] ^ n[38867];
assign t[38868] = t[38867] ^ n[38868];
assign t[38869] = t[38868] ^ n[38869];
assign t[38870] = t[38869] ^ n[38870];
assign t[38871] = t[38870] ^ n[38871];
assign t[38872] = t[38871] ^ n[38872];
assign t[38873] = t[38872] ^ n[38873];
assign t[38874] = t[38873] ^ n[38874];
assign t[38875] = t[38874] ^ n[38875];
assign t[38876] = t[38875] ^ n[38876];
assign t[38877] = t[38876] ^ n[38877];
assign t[38878] = t[38877] ^ n[38878];
assign t[38879] = t[38878] ^ n[38879];
assign t[38880] = t[38879] ^ n[38880];
assign t[38881] = t[38880] ^ n[38881];
assign t[38882] = t[38881] ^ n[38882];
assign t[38883] = t[38882] ^ n[38883];
assign t[38884] = t[38883] ^ n[38884];
assign t[38885] = t[38884] ^ n[38885];
assign t[38886] = t[38885] ^ n[38886];
assign t[38887] = t[38886] ^ n[38887];
assign t[38888] = t[38887] ^ n[38888];
assign t[38889] = t[38888] ^ n[38889];
assign t[38890] = t[38889] ^ n[38890];
assign t[38891] = t[38890] ^ n[38891];
assign t[38892] = t[38891] ^ n[38892];
assign t[38893] = t[38892] ^ n[38893];
assign t[38894] = t[38893] ^ n[38894];
assign t[38895] = t[38894] ^ n[38895];
assign t[38896] = t[38895] ^ n[38896];
assign t[38897] = t[38896] ^ n[38897];
assign t[38898] = t[38897] ^ n[38898];
assign t[38899] = t[38898] ^ n[38899];
assign t[38900] = t[38899] ^ n[38900];
assign t[38901] = t[38900] ^ n[38901];
assign t[38902] = t[38901] ^ n[38902];
assign t[38903] = t[38902] ^ n[38903];
assign t[38904] = t[38903] ^ n[38904];
assign t[38905] = t[38904] ^ n[38905];
assign t[38906] = t[38905] ^ n[38906];
assign t[38907] = t[38906] ^ n[38907];
assign t[38908] = t[38907] ^ n[38908];
assign t[38909] = t[38908] ^ n[38909];
assign t[38910] = t[38909] ^ n[38910];
assign t[38911] = t[38910] ^ n[38911];
assign t[38912] = t[38911] ^ n[38912];
assign t[38913] = t[38912] ^ n[38913];
assign t[38914] = t[38913] ^ n[38914];
assign t[38915] = t[38914] ^ n[38915];
assign t[38916] = t[38915] ^ n[38916];
assign t[38917] = t[38916] ^ n[38917];
assign t[38918] = t[38917] ^ n[38918];
assign t[38919] = t[38918] ^ n[38919];
assign t[38920] = t[38919] ^ n[38920];
assign t[38921] = t[38920] ^ n[38921];
assign t[38922] = t[38921] ^ n[38922];
assign t[38923] = t[38922] ^ n[38923];
assign t[38924] = t[38923] ^ n[38924];
assign t[38925] = t[38924] ^ n[38925];
assign t[38926] = t[38925] ^ n[38926];
assign t[38927] = t[38926] ^ n[38927];
assign t[38928] = t[38927] ^ n[38928];
assign t[38929] = t[38928] ^ n[38929];
assign t[38930] = t[38929] ^ n[38930];
assign t[38931] = t[38930] ^ n[38931];
assign t[38932] = t[38931] ^ n[38932];
assign t[38933] = t[38932] ^ n[38933];
assign t[38934] = t[38933] ^ n[38934];
assign t[38935] = t[38934] ^ n[38935];
assign t[38936] = t[38935] ^ n[38936];
assign t[38937] = t[38936] ^ n[38937];
assign t[38938] = t[38937] ^ n[38938];
assign t[38939] = t[38938] ^ n[38939];
assign t[38940] = t[38939] ^ n[38940];
assign t[38941] = t[38940] ^ n[38941];
assign t[38942] = t[38941] ^ n[38942];
assign t[38943] = t[38942] ^ n[38943];
assign t[38944] = t[38943] ^ n[38944];
assign t[38945] = t[38944] ^ n[38945];
assign t[38946] = t[38945] ^ n[38946];
assign t[38947] = t[38946] ^ n[38947];
assign t[38948] = t[38947] ^ n[38948];
assign t[38949] = t[38948] ^ n[38949];
assign t[38950] = t[38949] ^ n[38950];
assign t[38951] = t[38950] ^ n[38951];
assign t[38952] = t[38951] ^ n[38952];
assign t[38953] = t[38952] ^ n[38953];
assign t[38954] = t[38953] ^ n[38954];
assign t[38955] = t[38954] ^ n[38955];
assign t[38956] = t[38955] ^ n[38956];
assign t[38957] = t[38956] ^ n[38957];
assign t[38958] = t[38957] ^ n[38958];
assign t[38959] = t[38958] ^ n[38959];
assign t[38960] = t[38959] ^ n[38960];
assign t[38961] = t[38960] ^ n[38961];
assign t[38962] = t[38961] ^ n[38962];
assign t[38963] = t[38962] ^ n[38963];
assign t[38964] = t[38963] ^ n[38964];
assign t[38965] = t[38964] ^ n[38965];
assign t[38966] = t[38965] ^ n[38966];
assign t[38967] = t[38966] ^ n[38967];
assign t[38968] = t[38967] ^ n[38968];
assign t[38969] = t[38968] ^ n[38969];
assign t[38970] = t[38969] ^ n[38970];
assign t[38971] = t[38970] ^ n[38971];
assign t[38972] = t[38971] ^ n[38972];
assign t[38973] = t[38972] ^ n[38973];
assign t[38974] = t[38973] ^ n[38974];
assign t[38975] = t[38974] ^ n[38975];
assign t[38976] = t[38975] ^ n[38976];
assign t[38977] = t[38976] ^ n[38977];
assign t[38978] = t[38977] ^ n[38978];
assign t[38979] = t[38978] ^ n[38979];
assign t[38980] = t[38979] ^ n[38980];
assign t[38981] = t[38980] ^ n[38981];
assign t[38982] = t[38981] ^ n[38982];
assign t[38983] = t[38982] ^ n[38983];
assign t[38984] = t[38983] ^ n[38984];
assign t[38985] = t[38984] ^ n[38985];
assign t[38986] = t[38985] ^ n[38986];
assign t[38987] = t[38986] ^ n[38987];
assign t[38988] = t[38987] ^ n[38988];
assign t[38989] = t[38988] ^ n[38989];
assign t[38990] = t[38989] ^ n[38990];
assign t[38991] = t[38990] ^ n[38991];
assign t[38992] = t[38991] ^ n[38992];
assign t[38993] = t[38992] ^ n[38993];
assign t[38994] = t[38993] ^ n[38994];
assign t[38995] = t[38994] ^ n[38995];
assign t[38996] = t[38995] ^ n[38996];
assign t[38997] = t[38996] ^ n[38997];
assign t[38998] = t[38997] ^ n[38998];
assign t[38999] = t[38998] ^ n[38999];
assign t[39000] = t[38999] ^ n[39000];
assign t[39001] = t[39000] ^ n[39001];
assign t[39002] = t[39001] ^ n[39002];
assign t[39003] = t[39002] ^ n[39003];
assign t[39004] = t[39003] ^ n[39004];
assign t[39005] = t[39004] ^ n[39005];
assign t[39006] = t[39005] ^ n[39006];
assign t[39007] = t[39006] ^ n[39007];
assign t[39008] = t[39007] ^ n[39008];
assign t[39009] = t[39008] ^ n[39009];
assign t[39010] = t[39009] ^ n[39010];
assign t[39011] = t[39010] ^ n[39011];
assign t[39012] = t[39011] ^ n[39012];
assign t[39013] = t[39012] ^ n[39013];
assign t[39014] = t[39013] ^ n[39014];
assign t[39015] = t[39014] ^ n[39015];
assign t[39016] = t[39015] ^ n[39016];
assign t[39017] = t[39016] ^ n[39017];
assign t[39018] = t[39017] ^ n[39018];
assign t[39019] = t[39018] ^ n[39019];
assign t[39020] = t[39019] ^ n[39020];
assign t[39021] = t[39020] ^ n[39021];
assign t[39022] = t[39021] ^ n[39022];
assign t[39023] = t[39022] ^ n[39023];
assign t[39024] = t[39023] ^ n[39024];
assign t[39025] = t[39024] ^ n[39025];
assign t[39026] = t[39025] ^ n[39026];
assign t[39027] = t[39026] ^ n[39027];
assign t[39028] = t[39027] ^ n[39028];
assign t[39029] = t[39028] ^ n[39029];
assign t[39030] = t[39029] ^ n[39030];
assign t[39031] = t[39030] ^ n[39031];
assign t[39032] = t[39031] ^ n[39032];
assign t[39033] = t[39032] ^ n[39033];
assign t[39034] = t[39033] ^ n[39034];
assign t[39035] = t[39034] ^ n[39035];
assign t[39036] = t[39035] ^ n[39036];
assign t[39037] = t[39036] ^ n[39037];
assign t[39038] = t[39037] ^ n[39038];
assign t[39039] = t[39038] ^ n[39039];
assign t[39040] = t[39039] ^ n[39040];
assign t[39041] = t[39040] ^ n[39041];
assign t[39042] = t[39041] ^ n[39042];
assign t[39043] = t[39042] ^ n[39043];
assign t[39044] = t[39043] ^ n[39044];
assign t[39045] = t[39044] ^ n[39045];
assign t[39046] = t[39045] ^ n[39046];
assign t[39047] = t[39046] ^ n[39047];
assign t[39048] = t[39047] ^ n[39048];
assign t[39049] = t[39048] ^ n[39049];
assign t[39050] = t[39049] ^ n[39050];
assign t[39051] = t[39050] ^ n[39051];
assign t[39052] = t[39051] ^ n[39052];
assign t[39053] = t[39052] ^ n[39053];
assign t[39054] = t[39053] ^ n[39054];
assign t[39055] = t[39054] ^ n[39055];
assign t[39056] = t[39055] ^ n[39056];
assign t[39057] = t[39056] ^ n[39057];
assign t[39058] = t[39057] ^ n[39058];
assign t[39059] = t[39058] ^ n[39059];
assign t[39060] = t[39059] ^ n[39060];
assign t[39061] = t[39060] ^ n[39061];
assign t[39062] = t[39061] ^ n[39062];
assign t[39063] = t[39062] ^ n[39063];
assign t[39064] = t[39063] ^ n[39064];
assign t[39065] = t[39064] ^ n[39065];
assign t[39066] = t[39065] ^ n[39066];
assign t[39067] = t[39066] ^ n[39067];
assign t[39068] = t[39067] ^ n[39068];
assign t[39069] = t[39068] ^ n[39069];
assign t[39070] = t[39069] ^ n[39070];
assign t[39071] = t[39070] ^ n[39071];
assign t[39072] = t[39071] ^ n[39072];
assign t[39073] = t[39072] ^ n[39073];
assign t[39074] = t[39073] ^ n[39074];
assign t[39075] = t[39074] ^ n[39075];
assign t[39076] = t[39075] ^ n[39076];
assign t[39077] = t[39076] ^ n[39077];
assign t[39078] = t[39077] ^ n[39078];
assign t[39079] = t[39078] ^ n[39079];
assign t[39080] = t[39079] ^ n[39080];
assign t[39081] = t[39080] ^ n[39081];
assign t[39082] = t[39081] ^ n[39082];
assign t[39083] = t[39082] ^ n[39083];
assign t[39084] = t[39083] ^ n[39084];
assign t[39085] = t[39084] ^ n[39085];
assign t[39086] = t[39085] ^ n[39086];
assign t[39087] = t[39086] ^ n[39087];
assign t[39088] = t[39087] ^ n[39088];
assign t[39089] = t[39088] ^ n[39089];
assign t[39090] = t[39089] ^ n[39090];
assign t[39091] = t[39090] ^ n[39091];
assign t[39092] = t[39091] ^ n[39092];
assign t[39093] = t[39092] ^ n[39093];
assign t[39094] = t[39093] ^ n[39094];
assign t[39095] = t[39094] ^ n[39095];
assign t[39096] = t[39095] ^ n[39096];
assign t[39097] = t[39096] ^ n[39097];
assign t[39098] = t[39097] ^ n[39098];
assign t[39099] = t[39098] ^ n[39099];
assign t[39100] = t[39099] ^ n[39100];
assign t[39101] = t[39100] ^ n[39101];
assign t[39102] = t[39101] ^ n[39102];
assign t[39103] = t[39102] ^ n[39103];
assign t[39104] = t[39103] ^ n[39104];
assign t[39105] = t[39104] ^ n[39105];
assign t[39106] = t[39105] ^ n[39106];
assign t[39107] = t[39106] ^ n[39107];
assign t[39108] = t[39107] ^ n[39108];
assign t[39109] = t[39108] ^ n[39109];
assign t[39110] = t[39109] ^ n[39110];
assign t[39111] = t[39110] ^ n[39111];
assign t[39112] = t[39111] ^ n[39112];
assign t[39113] = t[39112] ^ n[39113];
assign t[39114] = t[39113] ^ n[39114];
assign t[39115] = t[39114] ^ n[39115];
assign t[39116] = t[39115] ^ n[39116];
assign t[39117] = t[39116] ^ n[39117];
assign t[39118] = t[39117] ^ n[39118];
assign t[39119] = t[39118] ^ n[39119];
assign t[39120] = t[39119] ^ n[39120];
assign t[39121] = t[39120] ^ n[39121];
assign t[39122] = t[39121] ^ n[39122];
assign t[39123] = t[39122] ^ n[39123];
assign t[39124] = t[39123] ^ n[39124];
assign t[39125] = t[39124] ^ n[39125];
assign t[39126] = t[39125] ^ n[39126];
assign t[39127] = t[39126] ^ n[39127];
assign t[39128] = t[39127] ^ n[39128];
assign t[39129] = t[39128] ^ n[39129];
assign t[39130] = t[39129] ^ n[39130];
assign t[39131] = t[39130] ^ n[39131];
assign t[39132] = t[39131] ^ n[39132];
assign t[39133] = t[39132] ^ n[39133];
assign t[39134] = t[39133] ^ n[39134];
assign t[39135] = t[39134] ^ n[39135];
assign t[39136] = t[39135] ^ n[39136];
assign t[39137] = t[39136] ^ n[39137];
assign t[39138] = t[39137] ^ n[39138];
assign t[39139] = t[39138] ^ n[39139];
assign t[39140] = t[39139] ^ n[39140];
assign t[39141] = t[39140] ^ n[39141];
assign t[39142] = t[39141] ^ n[39142];
assign t[39143] = t[39142] ^ n[39143];
assign t[39144] = t[39143] ^ n[39144];
assign t[39145] = t[39144] ^ n[39145];
assign t[39146] = t[39145] ^ n[39146];
assign t[39147] = t[39146] ^ n[39147];
assign t[39148] = t[39147] ^ n[39148];
assign t[39149] = t[39148] ^ n[39149];
assign t[39150] = t[39149] ^ n[39150];
assign t[39151] = t[39150] ^ n[39151];
assign t[39152] = t[39151] ^ n[39152];
assign t[39153] = t[39152] ^ n[39153];
assign t[39154] = t[39153] ^ n[39154];
assign t[39155] = t[39154] ^ n[39155];
assign t[39156] = t[39155] ^ n[39156];
assign t[39157] = t[39156] ^ n[39157];
assign t[39158] = t[39157] ^ n[39158];
assign t[39159] = t[39158] ^ n[39159];
assign t[39160] = t[39159] ^ n[39160];
assign t[39161] = t[39160] ^ n[39161];
assign t[39162] = t[39161] ^ n[39162];
assign t[39163] = t[39162] ^ n[39163];
assign t[39164] = t[39163] ^ n[39164];
assign t[39165] = t[39164] ^ n[39165];
assign t[39166] = t[39165] ^ n[39166];
assign t[39167] = t[39166] ^ n[39167];
assign t[39168] = t[39167] ^ n[39168];
assign t[39169] = t[39168] ^ n[39169];
assign t[39170] = t[39169] ^ n[39170];
assign t[39171] = t[39170] ^ n[39171];
assign t[39172] = t[39171] ^ n[39172];
assign t[39173] = t[39172] ^ n[39173];
assign t[39174] = t[39173] ^ n[39174];
assign t[39175] = t[39174] ^ n[39175];
assign t[39176] = t[39175] ^ n[39176];
assign t[39177] = t[39176] ^ n[39177];
assign t[39178] = t[39177] ^ n[39178];
assign t[39179] = t[39178] ^ n[39179];
assign t[39180] = t[39179] ^ n[39180];
assign t[39181] = t[39180] ^ n[39181];
assign t[39182] = t[39181] ^ n[39182];
assign t[39183] = t[39182] ^ n[39183];
assign t[39184] = t[39183] ^ n[39184];
assign t[39185] = t[39184] ^ n[39185];
assign t[39186] = t[39185] ^ n[39186];
assign t[39187] = t[39186] ^ n[39187];
assign t[39188] = t[39187] ^ n[39188];
assign t[39189] = t[39188] ^ n[39189];
assign t[39190] = t[39189] ^ n[39190];
assign t[39191] = t[39190] ^ n[39191];
assign t[39192] = t[39191] ^ n[39192];
assign t[39193] = t[39192] ^ n[39193];
assign t[39194] = t[39193] ^ n[39194];
assign t[39195] = t[39194] ^ n[39195];
assign t[39196] = t[39195] ^ n[39196];
assign t[39197] = t[39196] ^ n[39197];
assign t[39198] = t[39197] ^ n[39198];
assign t[39199] = t[39198] ^ n[39199];
assign t[39200] = t[39199] ^ n[39200];
assign t[39201] = t[39200] ^ n[39201];
assign t[39202] = t[39201] ^ n[39202];
assign t[39203] = t[39202] ^ n[39203];
assign t[39204] = t[39203] ^ n[39204];
assign t[39205] = t[39204] ^ n[39205];
assign t[39206] = t[39205] ^ n[39206];
assign t[39207] = t[39206] ^ n[39207];
assign t[39208] = t[39207] ^ n[39208];
assign t[39209] = t[39208] ^ n[39209];
assign t[39210] = t[39209] ^ n[39210];
assign t[39211] = t[39210] ^ n[39211];
assign t[39212] = t[39211] ^ n[39212];
assign t[39213] = t[39212] ^ n[39213];
assign t[39214] = t[39213] ^ n[39214];
assign t[39215] = t[39214] ^ n[39215];
assign t[39216] = t[39215] ^ n[39216];
assign t[39217] = t[39216] ^ n[39217];
assign t[39218] = t[39217] ^ n[39218];
assign t[39219] = t[39218] ^ n[39219];
assign t[39220] = t[39219] ^ n[39220];
assign t[39221] = t[39220] ^ n[39221];
assign t[39222] = t[39221] ^ n[39222];
assign t[39223] = t[39222] ^ n[39223];
assign t[39224] = t[39223] ^ n[39224];
assign t[39225] = t[39224] ^ n[39225];
assign t[39226] = t[39225] ^ n[39226];
assign t[39227] = t[39226] ^ n[39227];
assign t[39228] = t[39227] ^ n[39228];
assign t[39229] = t[39228] ^ n[39229];
assign t[39230] = t[39229] ^ n[39230];
assign t[39231] = t[39230] ^ n[39231];
assign t[39232] = t[39231] ^ n[39232];
assign t[39233] = t[39232] ^ n[39233];
assign t[39234] = t[39233] ^ n[39234];
assign t[39235] = t[39234] ^ n[39235];
assign t[39236] = t[39235] ^ n[39236];
assign t[39237] = t[39236] ^ n[39237];
assign t[39238] = t[39237] ^ n[39238];
assign t[39239] = t[39238] ^ n[39239];
assign t[39240] = t[39239] ^ n[39240];
assign t[39241] = t[39240] ^ n[39241];
assign t[39242] = t[39241] ^ n[39242];
assign t[39243] = t[39242] ^ n[39243];
assign t[39244] = t[39243] ^ n[39244];
assign t[39245] = t[39244] ^ n[39245];
assign t[39246] = t[39245] ^ n[39246];
assign t[39247] = t[39246] ^ n[39247];
assign t[39248] = t[39247] ^ n[39248];
assign t[39249] = t[39248] ^ n[39249];
assign t[39250] = t[39249] ^ n[39250];
assign t[39251] = t[39250] ^ n[39251];
assign t[39252] = t[39251] ^ n[39252];
assign t[39253] = t[39252] ^ n[39253];
assign t[39254] = t[39253] ^ n[39254];
assign t[39255] = t[39254] ^ n[39255];
assign t[39256] = t[39255] ^ n[39256];
assign t[39257] = t[39256] ^ n[39257];
assign t[39258] = t[39257] ^ n[39258];
assign t[39259] = t[39258] ^ n[39259];
assign t[39260] = t[39259] ^ n[39260];
assign t[39261] = t[39260] ^ n[39261];
assign t[39262] = t[39261] ^ n[39262];
assign t[39263] = t[39262] ^ n[39263];
assign t[39264] = t[39263] ^ n[39264];
assign t[39265] = t[39264] ^ n[39265];
assign t[39266] = t[39265] ^ n[39266];
assign t[39267] = t[39266] ^ n[39267];
assign t[39268] = t[39267] ^ n[39268];
assign t[39269] = t[39268] ^ n[39269];
assign t[39270] = t[39269] ^ n[39270];
assign t[39271] = t[39270] ^ n[39271];
assign t[39272] = t[39271] ^ n[39272];
assign t[39273] = t[39272] ^ n[39273];
assign t[39274] = t[39273] ^ n[39274];
assign t[39275] = t[39274] ^ n[39275];
assign t[39276] = t[39275] ^ n[39276];
assign t[39277] = t[39276] ^ n[39277];
assign t[39278] = t[39277] ^ n[39278];
assign t[39279] = t[39278] ^ n[39279];
assign t[39280] = t[39279] ^ n[39280];
assign t[39281] = t[39280] ^ n[39281];
assign t[39282] = t[39281] ^ n[39282];
assign t[39283] = t[39282] ^ n[39283];
assign t[39284] = t[39283] ^ n[39284];
assign t[39285] = t[39284] ^ n[39285];
assign t[39286] = t[39285] ^ n[39286];
assign t[39287] = t[39286] ^ n[39287];
assign t[39288] = t[39287] ^ n[39288];
assign t[39289] = t[39288] ^ n[39289];
assign t[39290] = t[39289] ^ n[39290];
assign t[39291] = t[39290] ^ n[39291];
assign t[39292] = t[39291] ^ n[39292];
assign t[39293] = t[39292] ^ n[39293];
assign t[39294] = t[39293] ^ n[39294];
assign t[39295] = t[39294] ^ n[39295];
assign t[39296] = t[39295] ^ n[39296];
assign t[39297] = t[39296] ^ n[39297];
assign t[39298] = t[39297] ^ n[39298];
assign t[39299] = t[39298] ^ n[39299];
assign t[39300] = t[39299] ^ n[39300];
assign t[39301] = t[39300] ^ n[39301];
assign t[39302] = t[39301] ^ n[39302];
assign t[39303] = t[39302] ^ n[39303];
assign t[39304] = t[39303] ^ n[39304];
assign t[39305] = t[39304] ^ n[39305];
assign t[39306] = t[39305] ^ n[39306];
assign t[39307] = t[39306] ^ n[39307];
assign t[39308] = t[39307] ^ n[39308];
assign t[39309] = t[39308] ^ n[39309];
assign t[39310] = t[39309] ^ n[39310];
assign t[39311] = t[39310] ^ n[39311];
assign t[39312] = t[39311] ^ n[39312];
assign t[39313] = t[39312] ^ n[39313];
assign t[39314] = t[39313] ^ n[39314];
assign t[39315] = t[39314] ^ n[39315];
assign t[39316] = t[39315] ^ n[39316];
assign t[39317] = t[39316] ^ n[39317];
assign t[39318] = t[39317] ^ n[39318];
assign t[39319] = t[39318] ^ n[39319];
assign t[39320] = t[39319] ^ n[39320];
assign t[39321] = t[39320] ^ n[39321];
assign t[39322] = t[39321] ^ n[39322];
assign t[39323] = t[39322] ^ n[39323];
assign t[39324] = t[39323] ^ n[39324];
assign t[39325] = t[39324] ^ n[39325];
assign t[39326] = t[39325] ^ n[39326];
assign t[39327] = t[39326] ^ n[39327];
assign t[39328] = t[39327] ^ n[39328];
assign t[39329] = t[39328] ^ n[39329];
assign t[39330] = t[39329] ^ n[39330];
assign t[39331] = t[39330] ^ n[39331];
assign t[39332] = t[39331] ^ n[39332];
assign t[39333] = t[39332] ^ n[39333];
assign t[39334] = t[39333] ^ n[39334];
assign t[39335] = t[39334] ^ n[39335];
assign t[39336] = t[39335] ^ n[39336];
assign t[39337] = t[39336] ^ n[39337];
assign t[39338] = t[39337] ^ n[39338];
assign t[39339] = t[39338] ^ n[39339];
assign t[39340] = t[39339] ^ n[39340];
assign t[39341] = t[39340] ^ n[39341];
assign t[39342] = t[39341] ^ n[39342];
assign t[39343] = t[39342] ^ n[39343];
assign t[39344] = t[39343] ^ n[39344];
assign t[39345] = t[39344] ^ n[39345];
assign t[39346] = t[39345] ^ n[39346];
assign t[39347] = t[39346] ^ n[39347];
assign t[39348] = t[39347] ^ n[39348];
assign t[39349] = t[39348] ^ n[39349];
assign t[39350] = t[39349] ^ n[39350];
assign t[39351] = t[39350] ^ n[39351];
assign t[39352] = t[39351] ^ n[39352];
assign t[39353] = t[39352] ^ n[39353];
assign t[39354] = t[39353] ^ n[39354];
assign t[39355] = t[39354] ^ n[39355];
assign t[39356] = t[39355] ^ n[39356];
assign t[39357] = t[39356] ^ n[39357];
assign t[39358] = t[39357] ^ n[39358];
assign t[39359] = t[39358] ^ n[39359];
assign t[39360] = t[39359] ^ n[39360];
assign t[39361] = t[39360] ^ n[39361];
assign t[39362] = t[39361] ^ n[39362];
assign t[39363] = t[39362] ^ n[39363];
assign t[39364] = t[39363] ^ n[39364];
assign t[39365] = t[39364] ^ n[39365];
assign t[39366] = t[39365] ^ n[39366];
assign t[39367] = t[39366] ^ n[39367];
assign t[39368] = t[39367] ^ n[39368];
assign t[39369] = t[39368] ^ n[39369];
assign t[39370] = t[39369] ^ n[39370];
assign t[39371] = t[39370] ^ n[39371];
assign t[39372] = t[39371] ^ n[39372];
assign t[39373] = t[39372] ^ n[39373];
assign t[39374] = t[39373] ^ n[39374];
assign t[39375] = t[39374] ^ n[39375];
assign t[39376] = t[39375] ^ n[39376];
assign t[39377] = t[39376] ^ n[39377];
assign t[39378] = t[39377] ^ n[39378];
assign t[39379] = t[39378] ^ n[39379];
assign t[39380] = t[39379] ^ n[39380];
assign t[39381] = t[39380] ^ n[39381];
assign t[39382] = t[39381] ^ n[39382];
assign t[39383] = t[39382] ^ n[39383];
assign t[39384] = t[39383] ^ n[39384];
assign t[39385] = t[39384] ^ n[39385];
assign t[39386] = t[39385] ^ n[39386];
assign t[39387] = t[39386] ^ n[39387];
assign t[39388] = t[39387] ^ n[39388];
assign t[39389] = t[39388] ^ n[39389];
assign t[39390] = t[39389] ^ n[39390];
assign t[39391] = t[39390] ^ n[39391];
assign t[39392] = t[39391] ^ n[39392];
assign t[39393] = t[39392] ^ n[39393];
assign t[39394] = t[39393] ^ n[39394];
assign t[39395] = t[39394] ^ n[39395];
assign t[39396] = t[39395] ^ n[39396];
assign t[39397] = t[39396] ^ n[39397];
assign t[39398] = t[39397] ^ n[39398];
assign t[39399] = t[39398] ^ n[39399];
assign t[39400] = t[39399] ^ n[39400];
assign t[39401] = t[39400] ^ n[39401];
assign t[39402] = t[39401] ^ n[39402];
assign t[39403] = t[39402] ^ n[39403];
assign t[39404] = t[39403] ^ n[39404];
assign t[39405] = t[39404] ^ n[39405];
assign t[39406] = t[39405] ^ n[39406];
assign t[39407] = t[39406] ^ n[39407];
assign t[39408] = t[39407] ^ n[39408];
assign t[39409] = t[39408] ^ n[39409];
assign t[39410] = t[39409] ^ n[39410];
assign t[39411] = t[39410] ^ n[39411];
assign t[39412] = t[39411] ^ n[39412];
assign t[39413] = t[39412] ^ n[39413];
assign t[39414] = t[39413] ^ n[39414];
assign t[39415] = t[39414] ^ n[39415];
assign t[39416] = t[39415] ^ n[39416];
assign t[39417] = t[39416] ^ n[39417];
assign t[39418] = t[39417] ^ n[39418];
assign t[39419] = t[39418] ^ n[39419];
assign t[39420] = t[39419] ^ n[39420];
assign t[39421] = t[39420] ^ n[39421];
assign t[39422] = t[39421] ^ n[39422];
assign t[39423] = t[39422] ^ n[39423];
assign t[39424] = t[39423] ^ n[39424];
assign t[39425] = t[39424] ^ n[39425];
assign t[39426] = t[39425] ^ n[39426];
assign t[39427] = t[39426] ^ n[39427];
assign t[39428] = t[39427] ^ n[39428];
assign t[39429] = t[39428] ^ n[39429];
assign t[39430] = t[39429] ^ n[39430];
assign t[39431] = t[39430] ^ n[39431];
assign t[39432] = t[39431] ^ n[39432];
assign t[39433] = t[39432] ^ n[39433];
assign t[39434] = t[39433] ^ n[39434];
assign t[39435] = t[39434] ^ n[39435];
assign t[39436] = t[39435] ^ n[39436];
assign t[39437] = t[39436] ^ n[39437];
assign t[39438] = t[39437] ^ n[39438];
assign t[39439] = t[39438] ^ n[39439];
assign t[39440] = t[39439] ^ n[39440];
assign t[39441] = t[39440] ^ n[39441];
assign t[39442] = t[39441] ^ n[39442];
assign t[39443] = t[39442] ^ n[39443];
assign t[39444] = t[39443] ^ n[39444];
assign t[39445] = t[39444] ^ n[39445];
assign t[39446] = t[39445] ^ n[39446];
assign t[39447] = t[39446] ^ n[39447];
assign t[39448] = t[39447] ^ n[39448];
assign t[39449] = t[39448] ^ n[39449];
assign t[39450] = t[39449] ^ n[39450];
assign t[39451] = t[39450] ^ n[39451];
assign t[39452] = t[39451] ^ n[39452];
assign t[39453] = t[39452] ^ n[39453];
assign t[39454] = t[39453] ^ n[39454];
assign t[39455] = t[39454] ^ n[39455];
assign t[39456] = t[39455] ^ n[39456];
assign t[39457] = t[39456] ^ n[39457];
assign t[39458] = t[39457] ^ n[39458];
assign t[39459] = t[39458] ^ n[39459];
assign t[39460] = t[39459] ^ n[39460];
assign t[39461] = t[39460] ^ n[39461];
assign t[39462] = t[39461] ^ n[39462];
assign t[39463] = t[39462] ^ n[39463];
assign t[39464] = t[39463] ^ n[39464];
assign t[39465] = t[39464] ^ n[39465];
assign t[39466] = t[39465] ^ n[39466];
assign t[39467] = t[39466] ^ n[39467];
assign t[39468] = t[39467] ^ n[39468];
assign t[39469] = t[39468] ^ n[39469];
assign t[39470] = t[39469] ^ n[39470];
assign t[39471] = t[39470] ^ n[39471];
assign t[39472] = t[39471] ^ n[39472];
assign t[39473] = t[39472] ^ n[39473];
assign t[39474] = t[39473] ^ n[39474];
assign t[39475] = t[39474] ^ n[39475];
assign t[39476] = t[39475] ^ n[39476];
assign t[39477] = t[39476] ^ n[39477];
assign t[39478] = t[39477] ^ n[39478];
assign t[39479] = t[39478] ^ n[39479];
assign t[39480] = t[39479] ^ n[39480];
assign t[39481] = t[39480] ^ n[39481];
assign t[39482] = t[39481] ^ n[39482];
assign t[39483] = t[39482] ^ n[39483];
assign t[39484] = t[39483] ^ n[39484];
assign t[39485] = t[39484] ^ n[39485];
assign t[39486] = t[39485] ^ n[39486];
assign t[39487] = t[39486] ^ n[39487];
assign t[39488] = t[39487] ^ n[39488];
assign t[39489] = t[39488] ^ n[39489];
assign t[39490] = t[39489] ^ n[39490];
assign t[39491] = t[39490] ^ n[39491];
assign t[39492] = t[39491] ^ n[39492];
assign t[39493] = t[39492] ^ n[39493];
assign t[39494] = t[39493] ^ n[39494];
assign t[39495] = t[39494] ^ n[39495];
assign t[39496] = t[39495] ^ n[39496];
assign t[39497] = t[39496] ^ n[39497];
assign t[39498] = t[39497] ^ n[39498];
assign t[39499] = t[39498] ^ n[39499];
assign t[39500] = t[39499] ^ n[39500];
assign t[39501] = t[39500] ^ n[39501];
assign t[39502] = t[39501] ^ n[39502];
assign t[39503] = t[39502] ^ n[39503];
assign t[39504] = t[39503] ^ n[39504];
assign t[39505] = t[39504] ^ n[39505];
assign t[39506] = t[39505] ^ n[39506];
assign t[39507] = t[39506] ^ n[39507];
assign t[39508] = t[39507] ^ n[39508];
assign t[39509] = t[39508] ^ n[39509];
assign t[39510] = t[39509] ^ n[39510];
assign t[39511] = t[39510] ^ n[39511];
assign t[39512] = t[39511] ^ n[39512];
assign t[39513] = t[39512] ^ n[39513];
assign t[39514] = t[39513] ^ n[39514];
assign t[39515] = t[39514] ^ n[39515];
assign t[39516] = t[39515] ^ n[39516];
assign t[39517] = t[39516] ^ n[39517];
assign t[39518] = t[39517] ^ n[39518];
assign t[39519] = t[39518] ^ n[39519];
assign t[39520] = t[39519] ^ n[39520];
assign t[39521] = t[39520] ^ n[39521];
assign t[39522] = t[39521] ^ n[39522];
assign t[39523] = t[39522] ^ n[39523];
assign t[39524] = t[39523] ^ n[39524];
assign t[39525] = t[39524] ^ n[39525];
assign t[39526] = t[39525] ^ n[39526];
assign t[39527] = t[39526] ^ n[39527];
assign t[39528] = t[39527] ^ n[39528];
assign t[39529] = t[39528] ^ n[39529];
assign t[39530] = t[39529] ^ n[39530];
assign t[39531] = t[39530] ^ n[39531];
assign t[39532] = t[39531] ^ n[39532];
assign t[39533] = t[39532] ^ n[39533];
assign t[39534] = t[39533] ^ n[39534];
assign t[39535] = t[39534] ^ n[39535];
assign t[39536] = t[39535] ^ n[39536];
assign t[39537] = t[39536] ^ n[39537];
assign t[39538] = t[39537] ^ n[39538];
assign t[39539] = t[39538] ^ n[39539];
assign t[39540] = t[39539] ^ n[39540];
assign t[39541] = t[39540] ^ n[39541];
assign t[39542] = t[39541] ^ n[39542];
assign t[39543] = t[39542] ^ n[39543];
assign t[39544] = t[39543] ^ n[39544];
assign t[39545] = t[39544] ^ n[39545];
assign t[39546] = t[39545] ^ n[39546];
assign t[39547] = t[39546] ^ n[39547];
assign t[39548] = t[39547] ^ n[39548];
assign t[39549] = t[39548] ^ n[39549];
assign t[39550] = t[39549] ^ n[39550];
assign t[39551] = t[39550] ^ n[39551];
assign t[39552] = t[39551] ^ n[39552];
assign t[39553] = t[39552] ^ n[39553];
assign t[39554] = t[39553] ^ n[39554];
assign t[39555] = t[39554] ^ n[39555];
assign t[39556] = t[39555] ^ n[39556];
assign t[39557] = t[39556] ^ n[39557];
assign t[39558] = t[39557] ^ n[39558];
assign t[39559] = t[39558] ^ n[39559];
assign t[39560] = t[39559] ^ n[39560];
assign t[39561] = t[39560] ^ n[39561];
assign t[39562] = t[39561] ^ n[39562];
assign t[39563] = t[39562] ^ n[39563];
assign t[39564] = t[39563] ^ n[39564];
assign t[39565] = t[39564] ^ n[39565];
assign t[39566] = t[39565] ^ n[39566];
assign t[39567] = t[39566] ^ n[39567];
assign t[39568] = t[39567] ^ n[39568];
assign t[39569] = t[39568] ^ n[39569];
assign t[39570] = t[39569] ^ n[39570];
assign t[39571] = t[39570] ^ n[39571];
assign t[39572] = t[39571] ^ n[39572];
assign t[39573] = t[39572] ^ n[39573];
assign t[39574] = t[39573] ^ n[39574];
assign t[39575] = t[39574] ^ n[39575];
assign t[39576] = t[39575] ^ n[39576];
assign t[39577] = t[39576] ^ n[39577];
assign t[39578] = t[39577] ^ n[39578];
assign t[39579] = t[39578] ^ n[39579];
assign t[39580] = t[39579] ^ n[39580];
assign t[39581] = t[39580] ^ n[39581];
assign t[39582] = t[39581] ^ n[39582];
assign t[39583] = t[39582] ^ n[39583];
assign t[39584] = t[39583] ^ n[39584];
assign t[39585] = t[39584] ^ n[39585];
assign t[39586] = t[39585] ^ n[39586];
assign t[39587] = t[39586] ^ n[39587];
assign t[39588] = t[39587] ^ n[39588];
assign t[39589] = t[39588] ^ n[39589];
assign t[39590] = t[39589] ^ n[39590];
assign t[39591] = t[39590] ^ n[39591];
assign t[39592] = t[39591] ^ n[39592];
assign t[39593] = t[39592] ^ n[39593];
assign t[39594] = t[39593] ^ n[39594];
assign t[39595] = t[39594] ^ n[39595];
assign t[39596] = t[39595] ^ n[39596];
assign t[39597] = t[39596] ^ n[39597];
assign t[39598] = t[39597] ^ n[39598];
assign t[39599] = t[39598] ^ n[39599];
assign t[39600] = t[39599] ^ n[39600];
assign t[39601] = t[39600] ^ n[39601];
assign t[39602] = t[39601] ^ n[39602];
assign t[39603] = t[39602] ^ n[39603];
assign t[39604] = t[39603] ^ n[39604];
assign t[39605] = t[39604] ^ n[39605];
assign t[39606] = t[39605] ^ n[39606];
assign t[39607] = t[39606] ^ n[39607];
assign t[39608] = t[39607] ^ n[39608];
assign t[39609] = t[39608] ^ n[39609];
assign t[39610] = t[39609] ^ n[39610];
assign t[39611] = t[39610] ^ n[39611];
assign t[39612] = t[39611] ^ n[39612];
assign t[39613] = t[39612] ^ n[39613];
assign t[39614] = t[39613] ^ n[39614];
assign t[39615] = t[39614] ^ n[39615];
assign t[39616] = t[39615] ^ n[39616];
assign t[39617] = t[39616] ^ n[39617];
assign t[39618] = t[39617] ^ n[39618];
assign t[39619] = t[39618] ^ n[39619];
assign t[39620] = t[39619] ^ n[39620];
assign t[39621] = t[39620] ^ n[39621];
assign t[39622] = t[39621] ^ n[39622];
assign t[39623] = t[39622] ^ n[39623];
assign t[39624] = t[39623] ^ n[39624];
assign t[39625] = t[39624] ^ n[39625];
assign t[39626] = t[39625] ^ n[39626];
assign t[39627] = t[39626] ^ n[39627];
assign t[39628] = t[39627] ^ n[39628];
assign t[39629] = t[39628] ^ n[39629];
assign t[39630] = t[39629] ^ n[39630];
assign t[39631] = t[39630] ^ n[39631];
assign t[39632] = t[39631] ^ n[39632];
assign t[39633] = t[39632] ^ n[39633];
assign t[39634] = t[39633] ^ n[39634];
assign t[39635] = t[39634] ^ n[39635];
assign t[39636] = t[39635] ^ n[39636];
assign t[39637] = t[39636] ^ n[39637];
assign t[39638] = t[39637] ^ n[39638];
assign t[39639] = t[39638] ^ n[39639];
assign t[39640] = t[39639] ^ n[39640];
assign t[39641] = t[39640] ^ n[39641];
assign t[39642] = t[39641] ^ n[39642];
assign t[39643] = t[39642] ^ n[39643];
assign t[39644] = t[39643] ^ n[39644];
assign t[39645] = t[39644] ^ n[39645];
assign t[39646] = t[39645] ^ n[39646];
assign t[39647] = t[39646] ^ n[39647];
assign t[39648] = t[39647] ^ n[39648];
assign t[39649] = t[39648] ^ n[39649];
assign t[39650] = t[39649] ^ n[39650];
assign t[39651] = t[39650] ^ n[39651];
assign t[39652] = t[39651] ^ n[39652];
assign t[39653] = t[39652] ^ n[39653];
assign t[39654] = t[39653] ^ n[39654];
assign t[39655] = t[39654] ^ n[39655];
assign t[39656] = t[39655] ^ n[39656];
assign t[39657] = t[39656] ^ n[39657];
assign t[39658] = t[39657] ^ n[39658];
assign t[39659] = t[39658] ^ n[39659];
assign t[39660] = t[39659] ^ n[39660];
assign t[39661] = t[39660] ^ n[39661];
assign t[39662] = t[39661] ^ n[39662];
assign t[39663] = t[39662] ^ n[39663];
assign t[39664] = t[39663] ^ n[39664];
assign t[39665] = t[39664] ^ n[39665];
assign t[39666] = t[39665] ^ n[39666];
assign t[39667] = t[39666] ^ n[39667];
assign t[39668] = t[39667] ^ n[39668];
assign t[39669] = t[39668] ^ n[39669];
assign t[39670] = t[39669] ^ n[39670];
assign t[39671] = t[39670] ^ n[39671];
assign t[39672] = t[39671] ^ n[39672];
assign t[39673] = t[39672] ^ n[39673];
assign t[39674] = t[39673] ^ n[39674];
assign t[39675] = t[39674] ^ n[39675];
assign t[39676] = t[39675] ^ n[39676];
assign t[39677] = t[39676] ^ n[39677];
assign t[39678] = t[39677] ^ n[39678];
assign t[39679] = t[39678] ^ n[39679];
assign t[39680] = t[39679] ^ n[39680];
assign t[39681] = t[39680] ^ n[39681];
assign t[39682] = t[39681] ^ n[39682];
assign t[39683] = t[39682] ^ n[39683];
assign t[39684] = t[39683] ^ n[39684];
assign t[39685] = t[39684] ^ n[39685];
assign t[39686] = t[39685] ^ n[39686];
assign t[39687] = t[39686] ^ n[39687];
assign t[39688] = t[39687] ^ n[39688];
assign t[39689] = t[39688] ^ n[39689];
assign t[39690] = t[39689] ^ n[39690];
assign t[39691] = t[39690] ^ n[39691];
assign t[39692] = t[39691] ^ n[39692];
assign t[39693] = t[39692] ^ n[39693];
assign t[39694] = t[39693] ^ n[39694];
assign t[39695] = t[39694] ^ n[39695];
assign t[39696] = t[39695] ^ n[39696];
assign t[39697] = t[39696] ^ n[39697];
assign t[39698] = t[39697] ^ n[39698];
assign t[39699] = t[39698] ^ n[39699];
assign t[39700] = t[39699] ^ n[39700];
assign t[39701] = t[39700] ^ n[39701];
assign t[39702] = t[39701] ^ n[39702];
assign t[39703] = t[39702] ^ n[39703];
assign t[39704] = t[39703] ^ n[39704];
assign t[39705] = t[39704] ^ n[39705];
assign t[39706] = t[39705] ^ n[39706];
assign t[39707] = t[39706] ^ n[39707];
assign t[39708] = t[39707] ^ n[39708];
assign t[39709] = t[39708] ^ n[39709];
assign t[39710] = t[39709] ^ n[39710];
assign t[39711] = t[39710] ^ n[39711];
assign t[39712] = t[39711] ^ n[39712];
assign t[39713] = t[39712] ^ n[39713];
assign t[39714] = t[39713] ^ n[39714];
assign t[39715] = t[39714] ^ n[39715];
assign t[39716] = t[39715] ^ n[39716];
assign t[39717] = t[39716] ^ n[39717];
assign t[39718] = t[39717] ^ n[39718];
assign t[39719] = t[39718] ^ n[39719];
assign t[39720] = t[39719] ^ n[39720];
assign t[39721] = t[39720] ^ n[39721];
assign t[39722] = t[39721] ^ n[39722];
assign t[39723] = t[39722] ^ n[39723];
assign t[39724] = t[39723] ^ n[39724];
assign t[39725] = t[39724] ^ n[39725];
assign t[39726] = t[39725] ^ n[39726];
assign t[39727] = t[39726] ^ n[39727];
assign t[39728] = t[39727] ^ n[39728];
assign t[39729] = t[39728] ^ n[39729];
assign t[39730] = t[39729] ^ n[39730];
assign t[39731] = t[39730] ^ n[39731];
assign t[39732] = t[39731] ^ n[39732];
assign t[39733] = t[39732] ^ n[39733];
assign t[39734] = t[39733] ^ n[39734];
assign t[39735] = t[39734] ^ n[39735];
assign t[39736] = t[39735] ^ n[39736];
assign t[39737] = t[39736] ^ n[39737];
assign t[39738] = t[39737] ^ n[39738];
assign t[39739] = t[39738] ^ n[39739];
assign t[39740] = t[39739] ^ n[39740];
assign t[39741] = t[39740] ^ n[39741];
assign t[39742] = t[39741] ^ n[39742];
assign t[39743] = t[39742] ^ n[39743];
assign t[39744] = t[39743] ^ n[39744];
assign t[39745] = t[39744] ^ n[39745];
assign t[39746] = t[39745] ^ n[39746];
assign t[39747] = t[39746] ^ n[39747];
assign t[39748] = t[39747] ^ n[39748];
assign t[39749] = t[39748] ^ n[39749];
assign t[39750] = t[39749] ^ n[39750];
assign t[39751] = t[39750] ^ n[39751];
assign t[39752] = t[39751] ^ n[39752];
assign t[39753] = t[39752] ^ n[39753];
assign t[39754] = t[39753] ^ n[39754];
assign t[39755] = t[39754] ^ n[39755];
assign t[39756] = t[39755] ^ n[39756];
assign t[39757] = t[39756] ^ n[39757];
assign t[39758] = t[39757] ^ n[39758];
assign t[39759] = t[39758] ^ n[39759];
assign t[39760] = t[39759] ^ n[39760];
assign t[39761] = t[39760] ^ n[39761];
assign t[39762] = t[39761] ^ n[39762];
assign t[39763] = t[39762] ^ n[39763];
assign t[39764] = t[39763] ^ n[39764];
assign t[39765] = t[39764] ^ n[39765];
assign t[39766] = t[39765] ^ n[39766];
assign t[39767] = t[39766] ^ n[39767];
assign t[39768] = t[39767] ^ n[39768];
assign t[39769] = t[39768] ^ n[39769];
assign t[39770] = t[39769] ^ n[39770];
assign t[39771] = t[39770] ^ n[39771];
assign t[39772] = t[39771] ^ n[39772];
assign t[39773] = t[39772] ^ n[39773];
assign t[39774] = t[39773] ^ n[39774];
assign t[39775] = t[39774] ^ n[39775];
assign t[39776] = t[39775] ^ n[39776];
assign t[39777] = t[39776] ^ n[39777];
assign t[39778] = t[39777] ^ n[39778];
assign t[39779] = t[39778] ^ n[39779];
assign t[39780] = t[39779] ^ n[39780];
assign t[39781] = t[39780] ^ n[39781];
assign t[39782] = t[39781] ^ n[39782];
assign t[39783] = t[39782] ^ n[39783];
assign t[39784] = t[39783] ^ n[39784];
assign t[39785] = t[39784] ^ n[39785];
assign t[39786] = t[39785] ^ n[39786];
assign t[39787] = t[39786] ^ n[39787];
assign t[39788] = t[39787] ^ n[39788];
assign t[39789] = t[39788] ^ n[39789];
assign t[39790] = t[39789] ^ n[39790];
assign t[39791] = t[39790] ^ n[39791];
assign t[39792] = t[39791] ^ n[39792];
assign t[39793] = t[39792] ^ n[39793];
assign t[39794] = t[39793] ^ n[39794];
assign t[39795] = t[39794] ^ n[39795];
assign t[39796] = t[39795] ^ n[39796];
assign t[39797] = t[39796] ^ n[39797];
assign t[39798] = t[39797] ^ n[39798];
assign t[39799] = t[39798] ^ n[39799];
assign t[39800] = t[39799] ^ n[39800];
assign t[39801] = t[39800] ^ n[39801];
assign t[39802] = t[39801] ^ n[39802];
assign t[39803] = t[39802] ^ n[39803];
assign t[39804] = t[39803] ^ n[39804];
assign t[39805] = t[39804] ^ n[39805];
assign t[39806] = t[39805] ^ n[39806];
assign t[39807] = t[39806] ^ n[39807];
assign t[39808] = t[39807] ^ n[39808];
assign t[39809] = t[39808] ^ n[39809];
assign t[39810] = t[39809] ^ n[39810];
assign t[39811] = t[39810] ^ n[39811];
assign t[39812] = t[39811] ^ n[39812];
assign t[39813] = t[39812] ^ n[39813];
assign t[39814] = t[39813] ^ n[39814];
assign t[39815] = t[39814] ^ n[39815];
assign t[39816] = t[39815] ^ n[39816];
assign t[39817] = t[39816] ^ n[39817];
assign t[39818] = t[39817] ^ n[39818];
assign t[39819] = t[39818] ^ n[39819];
assign t[39820] = t[39819] ^ n[39820];
assign t[39821] = t[39820] ^ n[39821];
assign t[39822] = t[39821] ^ n[39822];
assign t[39823] = t[39822] ^ n[39823];
assign t[39824] = t[39823] ^ n[39824];
assign t[39825] = t[39824] ^ n[39825];
assign t[39826] = t[39825] ^ n[39826];
assign t[39827] = t[39826] ^ n[39827];
assign t[39828] = t[39827] ^ n[39828];
assign t[39829] = t[39828] ^ n[39829];
assign t[39830] = t[39829] ^ n[39830];
assign t[39831] = t[39830] ^ n[39831];
assign t[39832] = t[39831] ^ n[39832];
assign t[39833] = t[39832] ^ n[39833];
assign t[39834] = t[39833] ^ n[39834];
assign t[39835] = t[39834] ^ n[39835];
assign t[39836] = t[39835] ^ n[39836];
assign t[39837] = t[39836] ^ n[39837];
assign t[39838] = t[39837] ^ n[39838];
assign t[39839] = t[39838] ^ n[39839];
assign t[39840] = t[39839] ^ n[39840];
assign t[39841] = t[39840] ^ n[39841];
assign t[39842] = t[39841] ^ n[39842];
assign t[39843] = t[39842] ^ n[39843];
assign t[39844] = t[39843] ^ n[39844];
assign t[39845] = t[39844] ^ n[39845];
assign t[39846] = t[39845] ^ n[39846];
assign t[39847] = t[39846] ^ n[39847];
assign t[39848] = t[39847] ^ n[39848];
assign t[39849] = t[39848] ^ n[39849];
assign t[39850] = t[39849] ^ n[39850];
assign t[39851] = t[39850] ^ n[39851];
assign t[39852] = t[39851] ^ n[39852];
assign t[39853] = t[39852] ^ n[39853];
assign t[39854] = t[39853] ^ n[39854];
assign t[39855] = t[39854] ^ n[39855];
assign t[39856] = t[39855] ^ n[39856];
assign t[39857] = t[39856] ^ n[39857];
assign t[39858] = t[39857] ^ n[39858];
assign t[39859] = t[39858] ^ n[39859];
assign t[39860] = t[39859] ^ n[39860];
assign t[39861] = t[39860] ^ n[39861];
assign t[39862] = t[39861] ^ n[39862];
assign t[39863] = t[39862] ^ n[39863];
assign t[39864] = t[39863] ^ n[39864];
assign t[39865] = t[39864] ^ n[39865];
assign t[39866] = t[39865] ^ n[39866];
assign t[39867] = t[39866] ^ n[39867];
assign t[39868] = t[39867] ^ n[39868];
assign t[39869] = t[39868] ^ n[39869];
assign t[39870] = t[39869] ^ n[39870];
assign t[39871] = t[39870] ^ n[39871];
assign t[39872] = t[39871] ^ n[39872];
assign t[39873] = t[39872] ^ n[39873];
assign t[39874] = t[39873] ^ n[39874];
assign t[39875] = t[39874] ^ n[39875];
assign t[39876] = t[39875] ^ n[39876];
assign t[39877] = t[39876] ^ n[39877];
assign t[39878] = t[39877] ^ n[39878];
assign t[39879] = t[39878] ^ n[39879];
assign t[39880] = t[39879] ^ n[39880];
assign t[39881] = t[39880] ^ n[39881];
assign t[39882] = t[39881] ^ n[39882];
assign t[39883] = t[39882] ^ n[39883];
assign t[39884] = t[39883] ^ n[39884];
assign t[39885] = t[39884] ^ n[39885];
assign t[39886] = t[39885] ^ n[39886];
assign t[39887] = t[39886] ^ n[39887];
assign t[39888] = t[39887] ^ n[39888];
assign t[39889] = t[39888] ^ n[39889];
assign t[39890] = t[39889] ^ n[39890];
assign t[39891] = t[39890] ^ n[39891];
assign t[39892] = t[39891] ^ n[39892];
assign t[39893] = t[39892] ^ n[39893];
assign t[39894] = t[39893] ^ n[39894];
assign t[39895] = t[39894] ^ n[39895];
assign t[39896] = t[39895] ^ n[39896];
assign t[39897] = t[39896] ^ n[39897];
assign t[39898] = t[39897] ^ n[39898];
assign t[39899] = t[39898] ^ n[39899];
assign t[39900] = t[39899] ^ n[39900];
assign t[39901] = t[39900] ^ n[39901];
assign t[39902] = t[39901] ^ n[39902];
assign t[39903] = t[39902] ^ n[39903];
assign t[39904] = t[39903] ^ n[39904];
assign t[39905] = t[39904] ^ n[39905];
assign t[39906] = t[39905] ^ n[39906];
assign t[39907] = t[39906] ^ n[39907];
assign t[39908] = t[39907] ^ n[39908];
assign t[39909] = t[39908] ^ n[39909];
assign t[39910] = t[39909] ^ n[39910];
assign t[39911] = t[39910] ^ n[39911];
assign t[39912] = t[39911] ^ n[39912];
assign t[39913] = t[39912] ^ n[39913];
assign t[39914] = t[39913] ^ n[39914];
assign t[39915] = t[39914] ^ n[39915];
assign t[39916] = t[39915] ^ n[39916];
assign t[39917] = t[39916] ^ n[39917];
assign t[39918] = t[39917] ^ n[39918];
assign t[39919] = t[39918] ^ n[39919];
assign t[39920] = t[39919] ^ n[39920];
assign t[39921] = t[39920] ^ n[39921];
assign t[39922] = t[39921] ^ n[39922];
assign t[39923] = t[39922] ^ n[39923];
assign t[39924] = t[39923] ^ n[39924];
assign t[39925] = t[39924] ^ n[39925];
assign t[39926] = t[39925] ^ n[39926];
assign t[39927] = t[39926] ^ n[39927];
assign t[39928] = t[39927] ^ n[39928];
assign t[39929] = t[39928] ^ n[39929];
assign t[39930] = t[39929] ^ n[39930];
assign t[39931] = t[39930] ^ n[39931];
assign t[39932] = t[39931] ^ n[39932];
assign t[39933] = t[39932] ^ n[39933];
assign t[39934] = t[39933] ^ n[39934];
assign t[39935] = t[39934] ^ n[39935];
assign t[39936] = t[39935] ^ n[39936];
assign t[39937] = t[39936] ^ n[39937];
assign t[39938] = t[39937] ^ n[39938];
assign t[39939] = t[39938] ^ n[39939];
assign t[39940] = t[39939] ^ n[39940];
assign t[39941] = t[39940] ^ n[39941];
assign t[39942] = t[39941] ^ n[39942];
assign t[39943] = t[39942] ^ n[39943];
assign t[39944] = t[39943] ^ n[39944];
assign t[39945] = t[39944] ^ n[39945];
assign t[39946] = t[39945] ^ n[39946];
assign t[39947] = t[39946] ^ n[39947];
assign t[39948] = t[39947] ^ n[39948];
assign t[39949] = t[39948] ^ n[39949];
assign t[39950] = t[39949] ^ n[39950];
assign t[39951] = t[39950] ^ n[39951];
assign t[39952] = t[39951] ^ n[39952];
assign t[39953] = t[39952] ^ n[39953];
assign t[39954] = t[39953] ^ n[39954];
assign t[39955] = t[39954] ^ n[39955];
assign t[39956] = t[39955] ^ n[39956];
assign t[39957] = t[39956] ^ n[39957];
assign t[39958] = t[39957] ^ n[39958];
assign t[39959] = t[39958] ^ n[39959];
assign t[39960] = t[39959] ^ n[39960];
assign t[39961] = t[39960] ^ n[39961];
assign t[39962] = t[39961] ^ n[39962];
assign t[39963] = t[39962] ^ n[39963];
assign t[39964] = t[39963] ^ n[39964];
assign t[39965] = t[39964] ^ n[39965];
assign t[39966] = t[39965] ^ n[39966];
assign t[39967] = t[39966] ^ n[39967];
assign t[39968] = t[39967] ^ n[39968];
assign t[39969] = t[39968] ^ n[39969];
assign t[39970] = t[39969] ^ n[39970];
assign t[39971] = t[39970] ^ n[39971];
assign t[39972] = t[39971] ^ n[39972];
assign t[39973] = t[39972] ^ n[39973];
assign t[39974] = t[39973] ^ n[39974];
assign t[39975] = t[39974] ^ n[39975];
assign t[39976] = t[39975] ^ n[39976];
assign t[39977] = t[39976] ^ n[39977];
assign t[39978] = t[39977] ^ n[39978];
assign t[39979] = t[39978] ^ n[39979];
assign t[39980] = t[39979] ^ n[39980];
assign t[39981] = t[39980] ^ n[39981];
assign t[39982] = t[39981] ^ n[39982];
assign t[39983] = t[39982] ^ n[39983];
assign t[39984] = t[39983] ^ n[39984];
assign t[39985] = t[39984] ^ n[39985];
assign t[39986] = t[39985] ^ n[39986];
assign t[39987] = t[39986] ^ n[39987];
assign t[39988] = t[39987] ^ n[39988];
assign t[39989] = t[39988] ^ n[39989];
assign t[39990] = t[39989] ^ n[39990];
assign t[39991] = t[39990] ^ n[39991];
assign t[39992] = t[39991] ^ n[39992];
assign t[39993] = t[39992] ^ n[39993];
assign t[39994] = t[39993] ^ n[39994];
assign t[39995] = t[39994] ^ n[39995];
assign t[39996] = t[39995] ^ n[39996];
assign t[39997] = t[39996] ^ n[39997];
assign t[39998] = t[39997] ^ n[39998];
assign t[39999] = t[39998] ^ n[39999];
assign t[40000] = t[39999] ^ n[40000];
assign t[40001] = t[40000] ^ n[40001];
assign t[40002] = t[40001] ^ n[40002];
assign t[40003] = t[40002] ^ n[40003];
assign t[40004] = t[40003] ^ n[40004];
assign t[40005] = t[40004] ^ n[40005];
assign t[40006] = t[40005] ^ n[40006];
assign t[40007] = t[40006] ^ n[40007];
assign t[40008] = t[40007] ^ n[40008];
assign t[40009] = t[40008] ^ n[40009];
assign t[40010] = t[40009] ^ n[40010];
assign t[40011] = t[40010] ^ n[40011];
assign t[40012] = t[40011] ^ n[40012];
assign t[40013] = t[40012] ^ n[40013];
assign t[40014] = t[40013] ^ n[40014];
assign t[40015] = t[40014] ^ n[40015];
assign t[40016] = t[40015] ^ n[40016];
assign t[40017] = t[40016] ^ n[40017];
assign t[40018] = t[40017] ^ n[40018];
assign t[40019] = t[40018] ^ n[40019];
assign t[40020] = t[40019] ^ n[40020];
assign t[40021] = t[40020] ^ n[40021];
assign t[40022] = t[40021] ^ n[40022];
assign t[40023] = t[40022] ^ n[40023];
assign t[40024] = t[40023] ^ n[40024];
assign t[40025] = t[40024] ^ n[40025];
assign t[40026] = t[40025] ^ n[40026];
assign t[40027] = t[40026] ^ n[40027];
assign t[40028] = t[40027] ^ n[40028];
assign t[40029] = t[40028] ^ n[40029];
assign t[40030] = t[40029] ^ n[40030];
assign t[40031] = t[40030] ^ n[40031];
assign t[40032] = t[40031] ^ n[40032];
assign t[40033] = t[40032] ^ n[40033];
assign t[40034] = t[40033] ^ n[40034];
assign t[40035] = t[40034] ^ n[40035];
assign t[40036] = t[40035] ^ n[40036];
assign t[40037] = t[40036] ^ n[40037];
assign t[40038] = t[40037] ^ n[40038];
assign t[40039] = t[40038] ^ n[40039];
assign t[40040] = t[40039] ^ n[40040];
assign t[40041] = t[40040] ^ n[40041];
assign t[40042] = t[40041] ^ n[40042];
assign t[40043] = t[40042] ^ n[40043];
assign t[40044] = t[40043] ^ n[40044];
assign t[40045] = t[40044] ^ n[40045];
assign t[40046] = t[40045] ^ n[40046];
assign t[40047] = t[40046] ^ n[40047];
assign t[40048] = t[40047] ^ n[40048];
assign t[40049] = t[40048] ^ n[40049];
assign t[40050] = t[40049] ^ n[40050];
assign t[40051] = t[40050] ^ n[40051];
assign t[40052] = t[40051] ^ n[40052];
assign t[40053] = t[40052] ^ n[40053];
assign t[40054] = t[40053] ^ n[40054];
assign t[40055] = t[40054] ^ n[40055];
assign t[40056] = t[40055] ^ n[40056];
assign t[40057] = t[40056] ^ n[40057];
assign t[40058] = t[40057] ^ n[40058];
assign t[40059] = t[40058] ^ n[40059];
assign t[40060] = t[40059] ^ n[40060];
assign t[40061] = t[40060] ^ n[40061];
assign t[40062] = t[40061] ^ n[40062];
assign t[40063] = t[40062] ^ n[40063];
assign t[40064] = t[40063] ^ n[40064];
assign t[40065] = t[40064] ^ n[40065];
assign t[40066] = t[40065] ^ n[40066];
assign t[40067] = t[40066] ^ n[40067];
assign t[40068] = t[40067] ^ n[40068];
assign t[40069] = t[40068] ^ n[40069];
assign t[40070] = t[40069] ^ n[40070];
assign t[40071] = t[40070] ^ n[40071];
assign t[40072] = t[40071] ^ n[40072];
assign t[40073] = t[40072] ^ n[40073];
assign t[40074] = t[40073] ^ n[40074];
assign t[40075] = t[40074] ^ n[40075];
assign t[40076] = t[40075] ^ n[40076];
assign t[40077] = t[40076] ^ n[40077];
assign t[40078] = t[40077] ^ n[40078];
assign t[40079] = t[40078] ^ n[40079];
assign t[40080] = t[40079] ^ n[40080];
assign t[40081] = t[40080] ^ n[40081];
assign t[40082] = t[40081] ^ n[40082];
assign t[40083] = t[40082] ^ n[40083];
assign t[40084] = t[40083] ^ n[40084];
assign t[40085] = t[40084] ^ n[40085];
assign t[40086] = t[40085] ^ n[40086];
assign t[40087] = t[40086] ^ n[40087];
assign t[40088] = t[40087] ^ n[40088];
assign t[40089] = t[40088] ^ n[40089];
assign t[40090] = t[40089] ^ n[40090];
assign t[40091] = t[40090] ^ n[40091];
assign t[40092] = t[40091] ^ n[40092];
assign t[40093] = t[40092] ^ n[40093];
assign t[40094] = t[40093] ^ n[40094];
assign t[40095] = t[40094] ^ n[40095];
assign t[40096] = t[40095] ^ n[40096];
assign t[40097] = t[40096] ^ n[40097];
assign t[40098] = t[40097] ^ n[40098];
assign t[40099] = t[40098] ^ n[40099];
assign t[40100] = t[40099] ^ n[40100];
assign t[40101] = t[40100] ^ n[40101];
assign t[40102] = t[40101] ^ n[40102];
assign t[40103] = t[40102] ^ n[40103];
assign t[40104] = t[40103] ^ n[40104];
assign t[40105] = t[40104] ^ n[40105];
assign t[40106] = t[40105] ^ n[40106];
assign t[40107] = t[40106] ^ n[40107];
assign t[40108] = t[40107] ^ n[40108];
assign t[40109] = t[40108] ^ n[40109];
assign t[40110] = t[40109] ^ n[40110];
assign t[40111] = t[40110] ^ n[40111];
assign t[40112] = t[40111] ^ n[40112];
assign t[40113] = t[40112] ^ n[40113];
assign t[40114] = t[40113] ^ n[40114];
assign t[40115] = t[40114] ^ n[40115];
assign t[40116] = t[40115] ^ n[40116];
assign t[40117] = t[40116] ^ n[40117];
assign t[40118] = t[40117] ^ n[40118];
assign t[40119] = t[40118] ^ n[40119];
assign t[40120] = t[40119] ^ n[40120];
assign t[40121] = t[40120] ^ n[40121];
assign t[40122] = t[40121] ^ n[40122];
assign t[40123] = t[40122] ^ n[40123];
assign t[40124] = t[40123] ^ n[40124];
assign t[40125] = t[40124] ^ n[40125];
assign t[40126] = t[40125] ^ n[40126];
assign t[40127] = t[40126] ^ n[40127];
assign t[40128] = t[40127] ^ n[40128];
assign t[40129] = t[40128] ^ n[40129];
assign t[40130] = t[40129] ^ n[40130];
assign t[40131] = t[40130] ^ n[40131];
assign t[40132] = t[40131] ^ n[40132];
assign t[40133] = t[40132] ^ n[40133];
assign t[40134] = t[40133] ^ n[40134];
assign t[40135] = t[40134] ^ n[40135];
assign t[40136] = t[40135] ^ n[40136];
assign t[40137] = t[40136] ^ n[40137];
assign t[40138] = t[40137] ^ n[40138];
assign t[40139] = t[40138] ^ n[40139];
assign t[40140] = t[40139] ^ n[40140];
assign t[40141] = t[40140] ^ n[40141];
assign t[40142] = t[40141] ^ n[40142];
assign t[40143] = t[40142] ^ n[40143];
assign t[40144] = t[40143] ^ n[40144];
assign t[40145] = t[40144] ^ n[40145];
assign t[40146] = t[40145] ^ n[40146];
assign t[40147] = t[40146] ^ n[40147];
assign t[40148] = t[40147] ^ n[40148];
assign t[40149] = t[40148] ^ n[40149];
assign t[40150] = t[40149] ^ n[40150];
assign t[40151] = t[40150] ^ n[40151];
assign t[40152] = t[40151] ^ n[40152];
assign t[40153] = t[40152] ^ n[40153];
assign t[40154] = t[40153] ^ n[40154];
assign t[40155] = t[40154] ^ n[40155];
assign t[40156] = t[40155] ^ n[40156];
assign t[40157] = t[40156] ^ n[40157];
assign t[40158] = t[40157] ^ n[40158];
assign t[40159] = t[40158] ^ n[40159];
assign t[40160] = t[40159] ^ n[40160];
assign t[40161] = t[40160] ^ n[40161];
assign t[40162] = t[40161] ^ n[40162];
assign t[40163] = t[40162] ^ n[40163];
assign t[40164] = t[40163] ^ n[40164];
assign t[40165] = t[40164] ^ n[40165];
assign t[40166] = t[40165] ^ n[40166];
assign t[40167] = t[40166] ^ n[40167];
assign t[40168] = t[40167] ^ n[40168];
assign t[40169] = t[40168] ^ n[40169];
assign t[40170] = t[40169] ^ n[40170];
assign t[40171] = t[40170] ^ n[40171];
assign t[40172] = t[40171] ^ n[40172];
assign t[40173] = t[40172] ^ n[40173];
assign t[40174] = t[40173] ^ n[40174];
assign t[40175] = t[40174] ^ n[40175];
assign t[40176] = t[40175] ^ n[40176];
assign t[40177] = t[40176] ^ n[40177];
assign t[40178] = t[40177] ^ n[40178];
assign t[40179] = t[40178] ^ n[40179];
assign t[40180] = t[40179] ^ n[40180];
assign t[40181] = t[40180] ^ n[40181];
assign t[40182] = t[40181] ^ n[40182];
assign t[40183] = t[40182] ^ n[40183];
assign t[40184] = t[40183] ^ n[40184];
assign t[40185] = t[40184] ^ n[40185];
assign t[40186] = t[40185] ^ n[40186];
assign t[40187] = t[40186] ^ n[40187];
assign t[40188] = t[40187] ^ n[40188];
assign t[40189] = t[40188] ^ n[40189];
assign t[40190] = t[40189] ^ n[40190];
assign t[40191] = t[40190] ^ n[40191];
assign t[40192] = t[40191] ^ n[40192];
assign t[40193] = t[40192] ^ n[40193];
assign t[40194] = t[40193] ^ n[40194];
assign t[40195] = t[40194] ^ n[40195];
assign t[40196] = t[40195] ^ n[40196];
assign t[40197] = t[40196] ^ n[40197];
assign t[40198] = t[40197] ^ n[40198];
assign t[40199] = t[40198] ^ n[40199];
assign t[40200] = t[40199] ^ n[40200];
assign t[40201] = t[40200] ^ n[40201];
assign t[40202] = t[40201] ^ n[40202];
assign t[40203] = t[40202] ^ n[40203];
assign t[40204] = t[40203] ^ n[40204];
assign t[40205] = t[40204] ^ n[40205];
assign t[40206] = t[40205] ^ n[40206];
assign t[40207] = t[40206] ^ n[40207];
assign t[40208] = t[40207] ^ n[40208];
assign t[40209] = t[40208] ^ n[40209];
assign t[40210] = t[40209] ^ n[40210];
assign t[40211] = t[40210] ^ n[40211];
assign t[40212] = t[40211] ^ n[40212];
assign t[40213] = t[40212] ^ n[40213];
assign t[40214] = t[40213] ^ n[40214];
assign t[40215] = t[40214] ^ n[40215];
assign t[40216] = t[40215] ^ n[40216];
assign t[40217] = t[40216] ^ n[40217];
assign t[40218] = t[40217] ^ n[40218];
assign t[40219] = t[40218] ^ n[40219];
assign t[40220] = t[40219] ^ n[40220];
assign t[40221] = t[40220] ^ n[40221];
assign t[40222] = t[40221] ^ n[40222];
assign t[40223] = t[40222] ^ n[40223];
assign t[40224] = t[40223] ^ n[40224];
assign t[40225] = t[40224] ^ n[40225];
assign t[40226] = t[40225] ^ n[40226];
assign t[40227] = t[40226] ^ n[40227];
assign t[40228] = t[40227] ^ n[40228];
assign t[40229] = t[40228] ^ n[40229];
assign t[40230] = t[40229] ^ n[40230];
assign t[40231] = t[40230] ^ n[40231];
assign t[40232] = t[40231] ^ n[40232];
assign t[40233] = t[40232] ^ n[40233];
assign t[40234] = t[40233] ^ n[40234];
assign t[40235] = t[40234] ^ n[40235];
assign t[40236] = t[40235] ^ n[40236];
assign t[40237] = t[40236] ^ n[40237];
assign t[40238] = t[40237] ^ n[40238];
assign t[40239] = t[40238] ^ n[40239];
assign t[40240] = t[40239] ^ n[40240];
assign t[40241] = t[40240] ^ n[40241];
assign t[40242] = t[40241] ^ n[40242];
assign t[40243] = t[40242] ^ n[40243];
assign t[40244] = t[40243] ^ n[40244];
assign t[40245] = t[40244] ^ n[40245];
assign t[40246] = t[40245] ^ n[40246];
assign t[40247] = t[40246] ^ n[40247];
assign t[40248] = t[40247] ^ n[40248];
assign t[40249] = t[40248] ^ n[40249];
assign t[40250] = t[40249] ^ n[40250];
assign t[40251] = t[40250] ^ n[40251];
assign t[40252] = t[40251] ^ n[40252];
assign t[40253] = t[40252] ^ n[40253];
assign t[40254] = t[40253] ^ n[40254];
assign t[40255] = t[40254] ^ n[40255];
assign t[40256] = t[40255] ^ n[40256];
assign t[40257] = t[40256] ^ n[40257];
assign t[40258] = t[40257] ^ n[40258];
assign t[40259] = t[40258] ^ n[40259];
assign t[40260] = t[40259] ^ n[40260];
assign t[40261] = t[40260] ^ n[40261];
assign t[40262] = t[40261] ^ n[40262];
assign t[40263] = t[40262] ^ n[40263];
assign t[40264] = t[40263] ^ n[40264];
assign t[40265] = t[40264] ^ n[40265];
assign t[40266] = t[40265] ^ n[40266];
assign t[40267] = t[40266] ^ n[40267];
assign t[40268] = t[40267] ^ n[40268];
assign t[40269] = t[40268] ^ n[40269];
assign t[40270] = t[40269] ^ n[40270];
assign t[40271] = t[40270] ^ n[40271];
assign t[40272] = t[40271] ^ n[40272];
assign t[40273] = t[40272] ^ n[40273];
assign t[40274] = t[40273] ^ n[40274];
assign t[40275] = t[40274] ^ n[40275];
assign t[40276] = t[40275] ^ n[40276];
assign t[40277] = t[40276] ^ n[40277];
assign t[40278] = t[40277] ^ n[40278];
assign t[40279] = t[40278] ^ n[40279];
assign t[40280] = t[40279] ^ n[40280];
assign t[40281] = t[40280] ^ n[40281];
assign t[40282] = t[40281] ^ n[40282];
assign t[40283] = t[40282] ^ n[40283];
assign t[40284] = t[40283] ^ n[40284];
assign t[40285] = t[40284] ^ n[40285];
assign t[40286] = t[40285] ^ n[40286];
assign t[40287] = t[40286] ^ n[40287];
assign t[40288] = t[40287] ^ n[40288];
assign t[40289] = t[40288] ^ n[40289];
assign t[40290] = t[40289] ^ n[40290];
assign t[40291] = t[40290] ^ n[40291];
assign t[40292] = t[40291] ^ n[40292];
assign t[40293] = t[40292] ^ n[40293];
assign t[40294] = t[40293] ^ n[40294];
assign t[40295] = t[40294] ^ n[40295];
assign t[40296] = t[40295] ^ n[40296];
assign t[40297] = t[40296] ^ n[40297];
assign t[40298] = t[40297] ^ n[40298];
assign t[40299] = t[40298] ^ n[40299];
assign t[40300] = t[40299] ^ n[40300];
assign t[40301] = t[40300] ^ n[40301];
assign t[40302] = t[40301] ^ n[40302];
assign t[40303] = t[40302] ^ n[40303];
assign t[40304] = t[40303] ^ n[40304];
assign t[40305] = t[40304] ^ n[40305];
assign t[40306] = t[40305] ^ n[40306];
assign t[40307] = t[40306] ^ n[40307];
assign t[40308] = t[40307] ^ n[40308];
assign t[40309] = t[40308] ^ n[40309];
assign t[40310] = t[40309] ^ n[40310];
assign t[40311] = t[40310] ^ n[40311];
assign t[40312] = t[40311] ^ n[40312];
assign t[40313] = t[40312] ^ n[40313];
assign t[40314] = t[40313] ^ n[40314];
assign t[40315] = t[40314] ^ n[40315];
assign t[40316] = t[40315] ^ n[40316];
assign t[40317] = t[40316] ^ n[40317];
assign t[40318] = t[40317] ^ n[40318];
assign t[40319] = t[40318] ^ n[40319];
assign t[40320] = t[40319] ^ n[40320];
assign t[40321] = t[40320] ^ n[40321];
assign t[40322] = t[40321] ^ n[40322];
assign t[40323] = t[40322] ^ n[40323];
assign t[40324] = t[40323] ^ n[40324];
assign t[40325] = t[40324] ^ n[40325];
assign t[40326] = t[40325] ^ n[40326];
assign t[40327] = t[40326] ^ n[40327];
assign t[40328] = t[40327] ^ n[40328];
assign t[40329] = t[40328] ^ n[40329];
assign t[40330] = t[40329] ^ n[40330];
assign t[40331] = t[40330] ^ n[40331];
assign t[40332] = t[40331] ^ n[40332];
assign t[40333] = t[40332] ^ n[40333];
assign t[40334] = t[40333] ^ n[40334];
assign t[40335] = t[40334] ^ n[40335];
assign t[40336] = t[40335] ^ n[40336];
assign t[40337] = t[40336] ^ n[40337];
assign t[40338] = t[40337] ^ n[40338];
assign t[40339] = t[40338] ^ n[40339];
assign t[40340] = t[40339] ^ n[40340];
assign t[40341] = t[40340] ^ n[40341];
assign t[40342] = t[40341] ^ n[40342];
assign t[40343] = t[40342] ^ n[40343];
assign t[40344] = t[40343] ^ n[40344];
assign t[40345] = t[40344] ^ n[40345];
assign t[40346] = t[40345] ^ n[40346];
assign t[40347] = t[40346] ^ n[40347];
assign t[40348] = t[40347] ^ n[40348];
assign t[40349] = t[40348] ^ n[40349];
assign t[40350] = t[40349] ^ n[40350];
assign t[40351] = t[40350] ^ n[40351];
assign t[40352] = t[40351] ^ n[40352];
assign t[40353] = t[40352] ^ n[40353];
assign t[40354] = t[40353] ^ n[40354];
assign t[40355] = t[40354] ^ n[40355];
assign t[40356] = t[40355] ^ n[40356];
assign t[40357] = t[40356] ^ n[40357];
assign t[40358] = t[40357] ^ n[40358];
assign t[40359] = t[40358] ^ n[40359];
assign t[40360] = t[40359] ^ n[40360];
assign t[40361] = t[40360] ^ n[40361];
assign t[40362] = t[40361] ^ n[40362];
assign t[40363] = t[40362] ^ n[40363];
assign t[40364] = t[40363] ^ n[40364];
assign t[40365] = t[40364] ^ n[40365];
assign t[40366] = t[40365] ^ n[40366];
assign t[40367] = t[40366] ^ n[40367];
assign t[40368] = t[40367] ^ n[40368];
assign t[40369] = t[40368] ^ n[40369];
assign t[40370] = t[40369] ^ n[40370];
assign t[40371] = t[40370] ^ n[40371];
assign t[40372] = t[40371] ^ n[40372];
assign t[40373] = t[40372] ^ n[40373];
assign t[40374] = t[40373] ^ n[40374];
assign t[40375] = t[40374] ^ n[40375];
assign t[40376] = t[40375] ^ n[40376];
assign t[40377] = t[40376] ^ n[40377];
assign t[40378] = t[40377] ^ n[40378];
assign t[40379] = t[40378] ^ n[40379];
assign t[40380] = t[40379] ^ n[40380];
assign t[40381] = t[40380] ^ n[40381];
assign t[40382] = t[40381] ^ n[40382];
assign t[40383] = t[40382] ^ n[40383];
assign t[40384] = t[40383] ^ n[40384];
assign t[40385] = t[40384] ^ n[40385];
assign t[40386] = t[40385] ^ n[40386];
assign t[40387] = t[40386] ^ n[40387];
assign t[40388] = t[40387] ^ n[40388];
assign t[40389] = t[40388] ^ n[40389];
assign t[40390] = t[40389] ^ n[40390];
assign t[40391] = t[40390] ^ n[40391];
assign t[40392] = t[40391] ^ n[40392];
assign t[40393] = t[40392] ^ n[40393];
assign t[40394] = t[40393] ^ n[40394];
assign t[40395] = t[40394] ^ n[40395];
assign t[40396] = t[40395] ^ n[40396];
assign t[40397] = t[40396] ^ n[40397];
assign t[40398] = t[40397] ^ n[40398];
assign t[40399] = t[40398] ^ n[40399];
assign t[40400] = t[40399] ^ n[40400];
assign t[40401] = t[40400] ^ n[40401];
assign t[40402] = t[40401] ^ n[40402];
assign t[40403] = t[40402] ^ n[40403];
assign t[40404] = t[40403] ^ n[40404];
assign t[40405] = t[40404] ^ n[40405];
assign t[40406] = t[40405] ^ n[40406];
assign t[40407] = t[40406] ^ n[40407];
assign t[40408] = t[40407] ^ n[40408];
assign t[40409] = t[40408] ^ n[40409];
assign t[40410] = t[40409] ^ n[40410];
assign t[40411] = t[40410] ^ n[40411];
assign t[40412] = t[40411] ^ n[40412];
assign t[40413] = t[40412] ^ n[40413];
assign t[40414] = t[40413] ^ n[40414];
assign t[40415] = t[40414] ^ n[40415];
assign t[40416] = t[40415] ^ n[40416];
assign t[40417] = t[40416] ^ n[40417];
assign t[40418] = t[40417] ^ n[40418];
assign t[40419] = t[40418] ^ n[40419];
assign t[40420] = t[40419] ^ n[40420];
assign t[40421] = t[40420] ^ n[40421];
assign t[40422] = t[40421] ^ n[40422];
assign t[40423] = t[40422] ^ n[40423];
assign t[40424] = t[40423] ^ n[40424];
assign t[40425] = t[40424] ^ n[40425];
assign t[40426] = t[40425] ^ n[40426];
assign t[40427] = t[40426] ^ n[40427];
assign t[40428] = t[40427] ^ n[40428];
assign t[40429] = t[40428] ^ n[40429];
assign t[40430] = t[40429] ^ n[40430];
assign t[40431] = t[40430] ^ n[40431];
assign t[40432] = t[40431] ^ n[40432];
assign t[40433] = t[40432] ^ n[40433];
assign t[40434] = t[40433] ^ n[40434];
assign t[40435] = t[40434] ^ n[40435];
assign t[40436] = t[40435] ^ n[40436];
assign t[40437] = t[40436] ^ n[40437];
assign t[40438] = t[40437] ^ n[40438];
assign t[40439] = t[40438] ^ n[40439];
assign t[40440] = t[40439] ^ n[40440];
assign t[40441] = t[40440] ^ n[40441];
assign t[40442] = t[40441] ^ n[40442];
assign t[40443] = t[40442] ^ n[40443];
assign t[40444] = t[40443] ^ n[40444];
assign t[40445] = t[40444] ^ n[40445];
assign t[40446] = t[40445] ^ n[40446];
assign t[40447] = t[40446] ^ n[40447];
assign t[40448] = t[40447] ^ n[40448];
assign t[40449] = t[40448] ^ n[40449];
assign t[40450] = t[40449] ^ n[40450];
assign t[40451] = t[40450] ^ n[40451];
assign t[40452] = t[40451] ^ n[40452];
assign t[40453] = t[40452] ^ n[40453];
assign t[40454] = t[40453] ^ n[40454];
assign t[40455] = t[40454] ^ n[40455];
assign t[40456] = t[40455] ^ n[40456];
assign t[40457] = t[40456] ^ n[40457];
assign t[40458] = t[40457] ^ n[40458];
assign t[40459] = t[40458] ^ n[40459];
assign t[40460] = t[40459] ^ n[40460];
assign t[40461] = t[40460] ^ n[40461];
assign t[40462] = t[40461] ^ n[40462];
assign t[40463] = t[40462] ^ n[40463];
assign t[40464] = t[40463] ^ n[40464];
assign t[40465] = t[40464] ^ n[40465];
assign t[40466] = t[40465] ^ n[40466];
assign t[40467] = t[40466] ^ n[40467];
assign t[40468] = t[40467] ^ n[40468];
assign t[40469] = t[40468] ^ n[40469];
assign t[40470] = t[40469] ^ n[40470];
assign t[40471] = t[40470] ^ n[40471];
assign t[40472] = t[40471] ^ n[40472];
assign t[40473] = t[40472] ^ n[40473];
assign t[40474] = t[40473] ^ n[40474];
assign t[40475] = t[40474] ^ n[40475];
assign t[40476] = t[40475] ^ n[40476];
assign t[40477] = t[40476] ^ n[40477];
assign t[40478] = t[40477] ^ n[40478];
assign t[40479] = t[40478] ^ n[40479];
assign t[40480] = t[40479] ^ n[40480];
assign t[40481] = t[40480] ^ n[40481];
assign t[40482] = t[40481] ^ n[40482];
assign t[40483] = t[40482] ^ n[40483];
assign t[40484] = t[40483] ^ n[40484];
assign t[40485] = t[40484] ^ n[40485];
assign t[40486] = t[40485] ^ n[40486];
assign t[40487] = t[40486] ^ n[40487];
assign t[40488] = t[40487] ^ n[40488];
assign t[40489] = t[40488] ^ n[40489];
assign t[40490] = t[40489] ^ n[40490];
assign t[40491] = t[40490] ^ n[40491];
assign t[40492] = t[40491] ^ n[40492];
assign t[40493] = t[40492] ^ n[40493];
assign t[40494] = t[40493] ^ n[40494];
assign t[40495] = t[40494] ^ n[40495];
assign t[40496] = t[40495] ^ n[40496];
assign t[40497] = t[40496] ^ n[40497];
assign t[40498] = t[40497] ^ n[40498];
assign t[40499] = t[40498] ^ n[40499];
assign t[40500] = t[40499] ^ n[40500];
assign t[40501] = t[40500] ^ n[40501];
assign t[40502] = t[40501] ^ n[40502];
assign t[40503] = t[40502] ^ n[40503];
assign t[40504] = t[40503] ^ n[40504];
assign t[40505] = t[40504] ^ n[40505];
assign t[40506] = t[40505] ^ n[40506];
assign t[40507] = t[40506] ^ n[40507];
assign t[40508] = t[40507] ^ n[40508];
assign t[40509] = t[40508] ^ n[40509];
assign t[40510] = t[40509] ^ n[40510];
assign t[40511] = t[40510] ^ n[40511];
assign t[40512] = t[40511] ^ n[40512];
assign t[40513] = t[40512] ^ n[40513];
assign t[40514] = t[40513] ^ n[40514];
assign t[40515] = t[40514] ^ n[40515];
assign t[40516] = t[40515] ^ n[40516];
assign t[40517] = t[40516] ^ n[40517];
assign t[40518] = t[40517] ^ n[40518];
assign t[40519] = t[40518] ^ n[40519];
assign t[40520] = t[40519] ^ n[40520];
assign t[40521] = t[40520] ^ n[40521];
assign t[40522] = t[40521] ^ n[40522];
assign t[40523] = t[40522] ^ n[40523];
assign t[40524] = t[40523] ^ n[40524];
assign t[40525] = t[40524] ^ n[40525];
assign t[40526] = t[40525] ^ n[40526];
assign t[40527] = t[40526] ^ n[40527];
assign t[40528] = t[40527] ^ n[40528];
assign t[40529] = t[40528] ^ n[40529];
assign t[40530] = t[40529] ^ n[40530];
assign t[40531] = t[40530] ^ n[40531];
assign t[40532] = t[40531] ^ n[40532];
assign t[40533] = t[40532] ^ n[40533];
assign t[40534] = t[40533] ^ n[40534];
assign t[40535] = t[40534] ^ n[40535];
assign t[40536] = t[40535] ^ n[40536];
assign t[40537] = t[40536] ^ n[40537];
assign t[40538] = t[40537] ^ n[40538];
assign t[40539] = t[40538] ^ n[40539];
assign t[40540] = t[40539] ^ n[40540];
assign t[40541] = t[40540] ^ n[40541];
assign t[40542] = t[40541] ^ n[40542];
assign t[40543] = t[40542] ^ n[40543];
assign t[40544] = t[40543] ^ n[40544];
assign t[40545] = t[40544] ^ n[40545];
assign t[40546] = t[40545] ^ n[40546];
assign t[40547] = t[40546] ^ n[40547];
assign t[40548] = t[40547] ^ n[40548];
assign t[40549] = t[40548] ^ n[40549];
assign t[40550] = t[40549] ^ n[40550];
assign t[40551] = t[40550] ^ n[40551];
assign t[40552] = t[40551] ^ n[40552];
assign t[40553] = t[40552] ^ n[40553];
assign t[40554] = t[40553] ^ n[40554];
assign t[40555] = t[40554] ^ n[40555];
assign t[40556] = t[40555] ^ n[40556];
assign t[40557] = t[40556] ^ n[40557];
assign t[40558] = t[40557] ^ n[40558];
assign t[40559] = t[40558] ^ n[40559];
assign t[40560] = t[40559] ^ n[40560];
assign t[40561] = t[40560] ^ n[40561];
assign t[40562] = t[40561] ^ n[40562];
assign t[40563] = t[40562] ^ n[40563];
assign t[40564] = t[40563] ^ n[40564];
assign t[40565] = t[40564] ^ n[40565];
assign t[40566] = t[40565] ^ n[40566];
assign t[40567] = t[40566] ^ n[40567];
assign t[40568] = t[40567] ^ n[40568];
assign t[40569] = t[40568] ^ n[40569];
assign t[40570] = t[40569] ^ n[40570];
assign t[40571] = t[40570] ^ n[40571];
assign t[40572] = t[40571] ^ n[40572];
assign t[40573] = t[40572] ^ n[40573];
assign t[40574] = t[40573] ^ n[40574];
assign t[40575] = t[40574] ^ n[40575];
assign t[40576] = t[40575] ^ n[40576];
assign t[40577] = t[40576] ^ n[40577];
assign t[40578] = t[40577] ^ n[40578];
assign t[40579] = t[40578] ^ n[40579];
assign t[40580] = t[40579] ^ n[40580];
assign t[40581] = t[40580] ^ n[40581];
assign t[40582] = t[40581] ^ n[40582];
assign t[40583] = t[40582] ^ n[40583];
assign t[40584] = t[40583] ^ n[40584];
assign t[40585] = t[40584] ^ n[40585];
assign t[40586] = t[40585] ^ n[40586];
assign t[40587] = t[40586] ^ n[40587];
assign t[40588] = t[40587] ^ n[40588];
assign t[40589] = t[40588] ^ n[40589];
assign t[40590] = t[40589] ^ n[40590];
assign t[40591] = t[40590] ^ n[40591];
assign t[40592] = t[40591] ^ n[40592];
assign t[40593] = t[40592] ^ n[40593];
assign t[40594] = t[40593] ^ n[40594];
assign t[40595] = t[40594] ^ n[40595];
assign t[40596] = t[40595] ^ n[40596];
assign t[40597] = t[40596] ^ n[40597];
assign t[40598] = t[40597] ^ n[40598];
assign t[40599] = t[40598] ^ n[40599];
assign t[40600] = t[40599] ^ n[40600];
assign t[40601] = t[40600] ^ n[40601];
assign t[40602] = t[40601] ^ n[40602];
assign t[40603] = t[40602] ^ n[40603];
assign t[40604] = t[40603] ^ n[40604];
assign t[40605] = t[40604] ^ n[40605];
assign t[40606] = t[40605] ^ n[40606];
assign t[40607] = t[40606] ^ n[40607];
assign t[40608] = t[40607] ^ n[40608];
assign t[40609] = t[40608] ^ n[40609];
assign t[40610] = t[40609] ^ n[40610];
assign t[40611] = t[40610] ^ n[40611];
assign t[40612] = t[40611] ^ n[40612];
assign t[40613] = t[40612] ^ n[40613];
assign t[40614] = t[40613] ^ n[40614];
assign t[40615] = t[40614] ^ n[40615];
assign t[40616] = t[40615] ^ n[40616];
assign t[40617] = t[40616] ^ n[40617];
assign t[40618] = t[40617] ^ n[40618];
assign t[40619] = t[40618] ^ n[40619];
assign t[40620] = t[40619] ^ n[40620];
assign t[40621] = t[40620] ^ n[40621];
assign t[40622] = t[40621] ^ n[40622];
assign t[40623] = t[40622] ^ n[40623];
assign t[40624] = t[40623] ^ n[40624];
assign t[40625] = t[40624] ^ n[40625];
assign t[40626] = t[40625] ^ n[40626];
assign t[40627] = t[40626] ^ n[40627];
assign t[40628] = t[40627] ^ n[40628];
assign t[40629] = t[40628] ^ n[40629];
assign t[40630] = t[40629] ^ n[40630];
assign t[40631] = t[40630] ^ n[40631];
assign t[40632] = t[40631] ^ n[40632];
assign t[40633] = t[40632] ^ n[40633];
assign t[40634] = t[40633] ^ n[40634];
assign t[40635] = t[40634] ^ n[40635];
assign t[40636] = t[40635] ^ n[40636];
assign t[40637] = t[40636] ^ n[40637];
assign t[40638] = t[40637] ^ n[40638];
assign t[40639] = t[40638] ^ n[40639];
assign t[40640] = t[40639] ^ n[40640];
assign t[40641] = t[40640] ^ n[40641];
assign t[40642] = t[40641] ^ n[40642];
assign t[40643] = t[40642] ^ n[40643];
assign t[40644] = t[40643] ^ n[40644];
assign t[40645] = t[40644] ^ n[40645];
assign t[40646] = t[40645] ^ n[40646];
assign t[40647] = t[40646] ^ n[40647];
assign t[40648] = t[40647] ^ n[40648];
assign t[40649] = t[40648] ^ n[40649];
assign t[40650] = t[40649] ^ n[40650];
assign t[40651] = t[40650] ^ n[40651];
assign t[40652] = t[40651] ^ n[40652];
assign t[40653] = t[40652] ^ n[40653];
assign t[40654] = t[40653] ^ n[40654];
assign t[40655] = t[40654] ^ n[40655];
assign t[40656] = t[40655] ^ n[40656];
assign t[40657] = t[40656] ^ n[40657];
assign t[40658] = t[40657] ^ n[40658];
assign t[40659] = t[40658] ^ n[40659];
assign t[40660] = t[40659] ^ n[40660];
assign t[40661] = t[40660] ^ n[40661];
assign t[40662] = t[40661] ^ n[40662];
assign t[40663] = t[40662] ^ n[40663];
assign t[40664] = t[40663] ^ n[40664];
assign t[40665] = t[40664] ^ n[40665];
assign t[40666] = t[40665] ^ n[40666];
assign t[40667] = t[40666] ^ n[40667];
assign t[40668] = t[40667] ^ n[40668];
assign t[40669] = t[40668] ^ n[40669];
assign t[40670] = t[40669] ^ n[40670];
assign t[40671] = t[40670] ^ n[40671];
assign t[40672] = t[40671] ^ n[40672];
assign t[40673] = t[40672] ^ n[40673];
assign t[40674] = t[40673] ^ n[40674];
assign t[40675] = t[40674] ^ n[40675];
assign t[40676] = t[40675] ^ n[40676];
assign t[40677] = t[40676] ^ n[40677];
assign t[40678] = t[40677] ^ n[40678];
assign t[40679] = t[40678] ^ n[40679];
assign t[40680] = t[40679] ^ n[40680];
assign t[40681] = t[40680] ^ n[40681];
assign t[40682] = t[40681] ^ n[40682];
assign t[40683] = t[40682] ^ n[40683];
assign t[40684] = t[40683] ^ n[40684];
assign t[40685] = t[40684] ^ n[40685];
assign t[40686] = t[40685] ^ n[40686];
assign t[40687] = t[40686] ^ n[40687];
assign t[40688] = t[40687] ^ n[40688];
assign t[40689] = t[40688] ^ n[40689];
assign t[40690] = t[40689] ^ n[40690];
assign t[40691] = t[40690] ^ n[40691];
assign t[40692] = t[40691] ^ n[40692];
assign t[40693] = t[40692] ^ n[40693];
assign t[40694] = t[40693] ^ n[40694];
assign t[40695] = t[40694] ^ n[40695];
assign t[40696] = t[40695] ^ n[40696];
assign t[40697] = t[40696] ^ n[40697];
assign t[40698] = t[40697] ^ n[40698];
assign t[40699] = t[40698] ^ n[40699];
assign t[40700] = t[40699] ^ n[40700];
assign t[40701] = t[40700] ^ n[40701];
assign t[40702] = t[40701] ^ n[40702];
assign t[40703] = t[40702] ^ n[40703];
assign t[40704] = t[40703] ^ n[40704];
assign t[40705] = t[40704] ^ n[40705];
assign t[40706] = t[40705] ^ n[40706];
assign t[40707] = t[40706] ^ n[40707];
assign t[40708] = t[40707] ^ n[40708];
assign t[40709] = t[40708] ^ n[40709];
assign t[40710] = t[40709] ^ n[40710];
assign t[40711] = t[40710] ^ n[40711];
assign t[40712] = t[40711] ^ n[40712];
assign t[40713] = t[40712] ^ n[40713];
assign t[40714] = t[40713] ^ n[40714];
assign t[40715] = t[40714] ^ n[40715];
assign t[40716] = t[40715] ^ n[40716];
assign t[40717] = t[40716] ^ n[40717];
assign t[40718] = t[40717] ^ n[40718];
assign t[40719] = t[40718] ^ n[40719];
assign t[40720] = t[40719] ^ n[40720];
assign t[40721] = t[40720] ^ n[40721];
assign t[40722] = t[40721] ^ n[40722];
assign t[40723] = t[40722] ^ n[40723];
assign t[40724] = t[40723] ^ n[40724];
assign t[40725] = t[40724] ^ n[40725];
assign t[40726] = t[40725] ^ n[40726];
assign t[40727] = t[40726] ^ n[40727];
assign t[40728] = t[40727] ^ n[40728];
assign t[40729] = t[40728] ^ n[40729];
assign t[40730] = t[40729] ^ n[40730];
assign t[40731] = t[40730] ^ n[40731];
assign t[40732] = t[40731] ^ n[40732];
assign t[40733] = t[40732] ^ n[40733];
assign t[40734] = t[40733] ^ n[40734];
assign t[40735] = t[40734] ^ n[40735];
assign t[40736] = t[40735] ^ n[40736];
assign t[40737] = t[40736] ^ n[40737];
assign t[40738] = t[40737] ^ n[40738];
assign t[40739] = t[40738] ^ n[40739];
assign t[40740] = t[40739] ^ n[40740];
assign t[40741] = t[40740] ^ n[40741];
assign t[40742] = t[40741] ^ n[40742];
assign t[40743] = t[40742] ^ n[40743];
assign t[40744] = t[40743] ^ n[40744];
assign t[40745] = t[40744] ^ n[40745];
assign t[40746] = t[40745] ^ n[40746];
assign t[40747] = t[40746] ^ n[40747];
assign t[40748] = t[40747] ^ n[40748];
assign t[40749] = t[40748] ^ n[40749];
assign t[40750] = t[40749] ^ n[40750];
assign t[40751] = t[40750] ^ n[40751];
assign t[40752] = t[40751] ^ n[40752];
assign t[40753] = t[40752] ^ n[40753];
assign t[40754] = t[40753] ^ n[40754];
assign t[40755] = t[40754] ^ n[40755];
assign t[40756] = t[40755] ^ n[40756];
assign t[40757] = t[40756] ^ n[40757];
assign t[40758] = t[40757] ^ n[40758];
assign t[40759] = t[40758] ^ n[40759];
assign t[40760] = t[40759] ^ n[40760];
assign t[40761] = t[40760] ^ n[40761];
assign t[40762] = t[40761] ^ n[40762];
assign t[40763] = t[40762] ^ n[40763];
assign t[40764] = t[40763] ^ n[40764];
assign t[40765] = t[40764] ^ n[40765];
assign t[40766] = t[40765] ^ n[40766];
assign t[40767] = t[40766] ^ n[40767];
assign t[40768] = t[40767] ^ n[40768];
assign t[40769] = t[40768] ^ n[40769];
assign t[40770] = t[40769] ^ n[40770];
assign t[40771] = t[40770] ^ n[40771];
assign t[40772] = t[40771] ^ n[40772];
assign t[40773] = t[40772] ^ n[40773];
assign t[40774] = t[40773] ^ n[40774];
assign t[40775] = t[40774] ^ n[40775];
assign t[40776] = t[40775] ^ n[40776];
assign t[40777] = t[40776] ^ n[40777];
assign t[40778] = t[40777] ^ n[40778];
assign t[40779] = t[40778] ^ n[40779];
assign t[40780] = t[40779] ^ n[40780];
assign t[40781] = t[40780] ^ n[40781];
assign t[40782] = t[40781] ^ n[40782];
assign t[40783] = t[40782] ^ n[40783];
assign t[40784] = t[40783] ^ n[40784];
assign t[40785] = t[40784] ^ n[40785];
assign t[40786] = t[40785] ^ n[40786];
assign t[40787] = t[40786] ^ n[40787];
assign t[40788] = t[40787] ^ n[40788];
assign t[40789] = t[40788] ^ n[40789];
assign t[40790] = t[40789] ^ n[40790];
assign t[40791] = t[40790] ^ n[40791];
assign t[40792] = t[40791] ^ n[40792];
assign t[40793] = t[40792] ^ n[40793];
assign t[40794] = t[40793] ^ n[40794];
assign t[40795] = t[40794] ^ n[40795];
assign t[40796] = t[40795] ^ n[40796];
assign t[40797] = t[40796] ^ n[40797];
assign t[40798] = t[40797] ^ n[40798];
assign t[40799] = t[40798] ^ n[40799];
assign t[40800] = t[40799] ^ n[40800];
assign t[40801] = t[40800] ^ n[40801];
assign t[40802] = t[40801] ^ n[40802];
assign t[40803] = t[40802] ^ n[40803];
assign t[40804] = t[40803] ^ n[40804];
assign t[40805] = t[40804] ^ n[40805];
assign t[40806] = t[40805] ^ n[40806];
assign t[40807] = t[40806] ^ n[40807];
assign t[40808] = t[40807] ^ n[40808];
assign t[40809] = t[40808] ^ n[40809];
assign t[40810] = t[40809] ^ n[40810];
assign t[40811] = t[40810] ^ n[40811];
assign t[40812] = t[40811] ^ n[40812];
assign t[40813] = t[40812] ^ n[40813];
assign t[40814] = t[40813] ^ n[40814];
assign t[40815] = t[40814] ^ n[40815];
assign t[40816] = t[40815] ^ n[40816];
assign t[40817] = t[40816] ^ n[40817];
assign t[40818] = t[40817] ^ n[40818];
assign t[40819] = t[40818] ^ n[40819];
assign t[40820] = t[40819] ^ n[40820];
assign t[40821] = t[40820] ^ n[40821];
assign t[40822] = t[40821] ^ n[40822];
assign t[40823] = t[40822] ^ n[40823];
assign t[40824] = t[40823] ^ n[40824];
assign t[40825] = t[40824] ^ n[40825];
assign t[40826] = t[40825] ^ n[40826];
assign t[40827] = t[40826] ^ n[40827];
assign t[40828] = t[40827] ^ n[40828];
assign t[40829] = t[40828] ^ n[40829];
assign t[40830] = t[40829] ^ n[40830];
assign t[40831] = t[40830] ^ n[40831];
assign t[40832] = t[40831] ^ n[40832];
assign t[40833] = t[40832] ^ n[40833];
assign t[40834] = t[40833] ^ n[40834];
assign t[40835] = t[40834] ^ n[40835];
assign t[40836] = t[40835] ^ n[40836];
assign t[40837] = t[40836] ^ n[40837];
assign t[40838] = t[40837] ^ n[40838];
assign t[40839] = t[40838] ^ n[40839];
assign t[40840] = t[40839] ^ n[40840];
assign t[40841] = t[40840] ^ n[40841];
assign t[40842] = t[40841] ^ n[40842];
assign t[40843] = t[40842] ^ n[40843];
assign t[40844] = t[40843] ^ n[40844];
assign t[40845] = t[40844] ^ n[40845];
assign t[40846] = t[40845] ^ n[40846];
assign t[40847] = t[40846] ^ n[40847];
assign t[40848] = t[40847] ^ n[40848];
assign t[40849] = t[40848] ^ n[40849];
assign t[40850] = t[40849] ^ n[40850];
assign t[40851] = t[40850] ^ n[40851];
assign t[40852] = t[40851] ^ n[40852];
assign t[40853] = t[40852] ^ n[40853];
assign t[40854] = t[40853] ^ n[40854];
assign t[40855] = t[40854] ^ n[40855];
assign t[40856] = t[40855] ^ n[40856];
assign t[40857] = t[40856] ^ n[40857];
assign t[40858] = t[40857] ^ n[40858];
assign t[40859] = t[40858] ^ n[40859];
assign t[40860] = t[40859] ^ n[40860];
assign t[40861] = t[40860] ^ n[40861];
assign t[40862] = t[40861] ^ n[40862];
assign t[40863] = t[40862] ^ n[40863];
assign t[40864] = t[40863] ^ n[40864];
assign t[40865] = t[40864] ^ n[40865];
assign t[40866] = t[40865] ^ n[40866];
assign t[40867] = t[40866] ^ n[40867];
assign t[40868] = t[40867] ^ n[40868];
assign t[40869] = t[40868] ^ n[40869];
assign t[40870] = t[40869] ^ n[40870];
assign t[40871] = t[40870] ^ n[40871];
assign t[40872] = t[40871] ^ n[40872];
assign t[40873] = t[40872] ^ n[40873];
assign t[40874] = t[40873] ^ n[40874];
assign t[40875] = t[40874] ^ n[40875];
assign t[40876] = t[40875] ^ n[40876];
assign t[40877] = t[40876] ^ n[40877];
assign t[40878] = t[40877] ^ n[40878];
assign t[40879] = t[40878] ^ n[40879];
assign t[40880] = t[40879] ^ n[40880];
assign t[40881] = t[40880] ^ n[40881];
assign t[40882] = t[40881] ^ n[40882];
assign t[40883] = t[40882] ^ n[40883];
assign t[40884] = t[40883] ^ n[40884];
assign t[40885] = t[40884] ^ n[40885];
assign t[40886] = t[40885] ^ n[40886];
assign t[40887] = t[40886] ^ n[40887];
assign t[40888] = t[40887] ^ n[40888];
assign t[40889] = t[40888] ^ n[40889];
assign t[40890] = t[40889] ^ n[40890];
assign t[40891] = t[40890] ^ n[40891];
assign t[40892] = t[40891] ^ n[40892];
assign t[40893] = t[40892] ^ n[40893];
assign t[40894] = t[40893] ^ n[40894];
assign t[40895] = t[40894] ^ n[40895];
assign t[40896] = t[40895] ^ n[40896];
assign t[40897] = t[40896] ^ n[40897];
assign t[40898] = t[40897] ^ n[40898];
assign t[40899] = t[40898] ^ n[40899];
assign t[40900] = t[40899] ^ n[40900];
assign t[40901] = t[40900] ^ n[40901];
assign t[40902] = t[40901] ^ n[40902];
assign t[40903] = t[40902] ^ n[40903];
assign t[40904] = t[40903] ^ n[40904];
assign t[40905] = t[40904] ^ n[40905];
assign t[40906] = t[40905] ^ n[40906];
assign t[40907] = t[40906] ^ n[40907];
assign t[40908] = t[40907] ^ n[40908];
assign t[40909] = t[40908] ^ n[40909];
assign t[40910] = t[40909] ^ n[40910];
assign t[40911] = t[40910] ^ n[40911];
assign t[40912] = t[40911] ^ n[40912];
assign t[40913] = t[40912] ^ n[40913];
assign t[40914] = t[40913] ^ n[40914];
assign t[40915] = t[40914] ^ n[40915];
assign t[40916] = t[40915] ^ n[40916];
assign t[40917] = t[40916] ^ n[40917];
assign t[40918] = t[40917] ^ n[40918];
assign t[40919] = t[40918] ^ n[40919];
assign t[40920] = t[40919] ^ n[40920];
assign t[40921] = t[40920] ^ n[40921];
assign t[40922] = t[40921] ^ n[40922];
assign t[40923] = t[40922] ^ n[40923];
assign t[40924] = t[40923] ^ n[40924];
assign t[40925] = t[40924] ^ n[40925];
assign t[40926] = t[40925] ^ n[40926];
assign t[40927] = t[40926] ^ n[40927];
assign t[40928] = t[40927] ^ n[40928];
assign t[40929] = t[40928] ^ n[40929];
assign t[40930] = t[40929] ^ n[40930];
assign t[40931] = t[40930] ^ n[40931];
assign t[40932] = t[40931] ^ n[40932];
assign t[40933] = t[40932] ^ n[40933];
assign t[40934] = t[40933] ^ n[40934];
assign t[40935] = t[40934] ^ n[40935];
assign t[40936] = t[40935] ^ n[40936];
assign t[40937] = t[40936] ^ n[40937];
assign t[40938] = t[40937] ^ n[40938];
assign t[40939] = t[40938] ^ n[40939];
assign t[40940] = t[40939] ^ n[40940];
assign t[40941] = t[40940] ^ n[40941];
assign t[40942] = t[40941] ^ n[40942];
assign t[40943] = t[40942] ^ n[40943];
assign t[40944] = t[40943] ^ n[40944];
assign t[40945] = t[40944] ^ n[40945];
assign t[40946] = t[40945] ^ n[40946];
assign t[40947] = t[40946] ^ n[40947];
assign t[40948] = t[40947] ^ n[40948];
assign t[40949] = t[40948] ^ n[40949];
assign t[40950] = t[40949] ^ n[40950];
assign t[40951] = t[40950] ^ n[40951];
assign t[40952] = t[40951] ^ n[40952];
assign t[40953] = t[40952] ^ n[40953];
assign t[40954] = t[40953] ^ n[40954];
assign t[40955] = t[40954] ^ n[40955];
assign t[40956] = t[40955] ^ n[40956];
assign t[40957] = t[40956] ^ n[40957];
assign t[40958] = t[40957] ^ n[40958];
assign t[40959] = t[40958] ^ n[40959];
assign t[40960] = t[40959] ^ n[40960];
assign t[40961] = t[40960] ^ n[40961];
assign t[40962] = t[40961] ^ n[40962];
assign t[40963] = t[40962] ^ n[40963];
assign t[40964] = t[40963] ^ n[40964];
assign t[40965] = t[40964] ^ n[40965];
assign t[40966] = t[40965] ^ n[40966];
assign t[40967] = t[40966] ^ n[40967];
assign t[40968] = t[40967] ^ n[40968];
assign t[40969] = t[40968] ^ n[40969];
assign t[40970] = t[40969] ^ n[40970];
assign t[40971] = t[40970] ^ n[40971];
assign t[40972] = t[40971] ^ n[40972];
assign t[40973] = t[40972] ^ n[40973];
assign t[40974] = t[40973] ^ n[40974];
assign t[40975] = t[40974] ^ n[40975];
assign t[40976] = t[40975] ^ n[40976];
assign t[40977] = t[40976] ^ n[40977];
assign t[40978] = t[40977] ^ n[40978];
assign t[40979] = t[40978] ^ n[40979];
assign t[40980] = t[40979] ^ n[40980];
assign t[40981] = t[40980] ^ n[40981];
assign t[40982] = t[40981] ^ n[40982];
assign t[40983] = t[40982] ^ n[40983];
assign t[40984] = t[40983] ^ n[40984];
assign t[40985] = t[40984] ^ n[40985];
assign t[40986] = t[40985] ^ n[40986];
assign t[40987] = t[40986] ^ n[40987];
assign t[40988] = t[40987] ^ n[40988];
assign t[40989] = t[40988] ^ n[40989];
assign t[40990] = t[40989] ^ n[40990];
assign t[40991] = t[40990] ^ n[40991];
assign t[40992] = t[40991] ^ n[40992];
assign t[40993] = t[40992] ^ n[40993];
assign t[40994] = t[40993] ^ n[40994];
assign t[40995] = t[40994] ^ n[40995];
assign t[40996] = t[40995] ^ n[40996];
assign t[40997] = t[40996] ^ n[40997];
assign t[40998] = t[40997] ^ n[40998];
assign t[40999] = t[40998] ^ n[40999];
assign t[41000] = t[40999] ^ n[41000];
assign t[41001] = t[41000] ^ n[41001];
assign t[41002] = t[41001] ^ n[41002];
assign t[41003] = t[41002] ^ n[41003];
assign t[41004] = t[41003] ^ n[41004];
assign t[41005] = t[41004] ^ n[41005];
assign t[41006] = t[41005] ^ n[41006];
assign t[41007] = t[41006] ^ n[41007];
assign t[41008] = t[41007] ^ n[41008];
assign t[41009] = t[41008] ^ n[41009];
assign t[41010] = t[41009] ^ n[41010];
assign t[41011] = t[41010] ^ n[41011];
assign t[41012] = t[41011] ^ n[41012];
assign t[41013] = t[41012] ^ n[41013];
assign t[41014] = t[41013] ^ n[41014];
assign t[41015] = t[41014] ^ n[41015];
assign t[41016] = t[41015] ^ n[41016];
assign t[41017] = t[41016] ^ n[41017];
assign t[41018] = t[41017] ^ n[41018];
assign t[41019] = t[41018] ^ n[41019];
assign t[41020] = t[41019] ^ n[41020];
assign t[41021] = t[41020] ^ n[41021];
assign t[41022] = t[41021] ^ n[41022];
assign t[41023] = t[41022] ^ n[41023];
assign t[41024] = t[41023] ^ n[41024];
assign t[41025] = t[41024] ^ n[41025];
assign t[41026] = t[41025] ^ n[41026];
assign t[41027] = t[41026] ^ n[41027];
assign t[41028] = t[41027] ^ n[41028];
assign t[41029] = t[41028] ^ n[41029];
assign t[41030] = t[41029] ^ n[41030];
assign t[41031] = t[41030] ^ n[41031];
assign t[41032] = t[41031] ^ n[41032];
assign t[41033] = t[41032] ^ n[41033];
assign t[41034] = t[41033] ^ n[41034];
assign t[41035] = t[41034] ^ n[41035];
assign t[41036] = t[41035] ^ n[41036];
assign t[41037] = t[41036] ^ n[41037];
assign t[41038] = t[41037] ^ n[41038];
assign t[41039] = t[41038] ^ n[41039];
assign t[41040] = t[41039] ^ n[41040];
assign t[41041] = t[41040] ^ n[41041];
assign t[41042] = t[41041] ^ n[41042];
assign t[41043] = t[41042] ^ n[41043];
assign t[41044] = t[41043] ^ n[41044];
assign t[41045] = t[41044] ^ n[41045];
assign t[41046] = t[41045] ^ n[41046];
assign t[41047] = t[41046] ^ n[41047];
assign t[41048] = t[41047] ^ n[41048];
assign t[41049] = t[41048] ^ n[41049];
assign t[41050] = t[41049] ^ n[41050];
assign t[41051] = t[41050] ^ n[41051];
assign t[41052] = t[41051] ^ n[41052];
assign t[41053] = t[41052] ^ n[41053];
assign t[41054] = t[41053] ^ n[41054];
assign t[41055] = t[41054] ^ n[41055];
assign t[41056] = t[41055] ^ n[41056];
assign t[41057] = t[41056] ^ n[41057];
assign t[41058] = t[41057] ^ n[41058];
assign t[41059] = t[41058] ^ n[41059];
assign t[41060] = t[41059] ^ n[41060];
assign t[41061] = t[41060] ^ n[41061];
assign t[41062] = t[41061] ^ n[41062];
assign t[41063] = t[41062] ^ n[41063];
assign t[41064] = t[41063] ^ n[41064];
assign t[41065] = t[41064] ^ n[41065];
assign t[41066] = t[41065] ^ n[41066];
assign t[41067] = t[41066] ^ n[41067];
assign t[41068] = t[41067] ^ n[41068];
assign t[41069] = t[41068] ^ n[41069];
assign t[41070] = t[41069] ^ n[41070];
assign t[41071] = t[41070] ^ n[41071];
assign t[41072] = t[41071] ^ n[41072];
assign t[41073] = t[41072] ^ n[41073];
assign t[41074] = t[41073] ^ n[41074];
assign t[41075] = t[41074] ^ n[41075];
assign t[41076] = t[41075] ^ n[41076];
assign t[41077] = t[41076] ^ n[41077];
assign t[41078] = t[41077] ^ n[41078];
assign t[41079] = t[41078] ^ n[41079];
assign t[41080] = t[41079] ^ n[41080];
assign t[41081] = t[41080] ^ n[41081];
assign t[41082] = t[41081] ^ n[41082];
assign t[41083] = t[41082] ^ n[41083];
assign t[41084] = t[41083] ^ n[41084];
assign t[41085] = t[41084] ^ n[41085];
assign t[41086] = t[41085] ^ n[41086];
assign t[41087] = t[41086] ^ n[41087];
assign t[41088] = t[41087] ^ n[41088];
assign t[41089] = t[41088] ^ n[41089];
assign t[41090] = t[41089] ^ n[41090];
assign t[41091] = t[41090] ^ n[41091];
assign t[41092] = t[41091] ^ n[41092];
assign t[41093] = t[41092] ^ n[41093];
assign t[41094] = t[41093] ^ n[41094];
assign t[41095] = t[41094] ^ n[41095];
assign t[41096] = t[41095] ^ n[41096];
assign t[41097] = t[41096] ^ n[41097];
assign t[41098] = t[41097] ^ n[41098];
assign t[41099] = t[41098] ^ n[41099];
assign t[41100] = t[41099] ^ n[41100];
assign t[41101] = t[41100] ^ n[41101];
assign t[41102] = t[41101] ^ n[41102];
assign t[41103] = t[41102] ^ n[41103];
assign t[41104] = t[41103] ^ n[41104];
assign t[41105] = t[41104] ^ n[41105];
assign t[41106] = t[41105] ^ n[41106];
assign t[41107] = t[41106] ^ n[41107];
assign t[41108] = t[41107] ^ n[41108];
assign t[41109] = t[41108] ^ n[41109];
assign t[41110] = t[41109] ^ n[41110];
assign t[41111] = t[41110] ^ n[41111];
assign t[41112] = t[41111] ^ n[41112];
assign t[41113] = t[41112] ^ n[41113];
assign t[41114] = t[41113] ^ n[41114];
assign t[41115] = t[41114] ^ n[41115];
assign t[41116] = t[41115] ^ n[41116];
assign t[41117] = t[41116] ^ n[41117];
assign t[41118] = t[41117] ^ n[41118];
assign t[41119] = t[41118] ^ n[41119];
assign t[41120] = t[41119] ^ n[41120];
assign t[41121] = t[41120] ^ n[41121];
assign t[41122] = t[41121] ^ n[41122];
assign t[41123] = t[41122] ^ n[41123];
assign t[41124] = t[41123] ^ n[41124];
assign t[41125] = t[41124] ^ n[41125];
assign t[41126] = t[41125] ^ n[41126];
assign t[41127] = t[41126] ^ n[41127];
assign t[41128] = t[41127] ^ n[41128];
assign t[41129] = t[41128] ^ n[41129];
assign t[41130] = t[41129] ^ n[41130];
assign t[41131] = t[41130] ^ n[41131];
assign t[41132] = t[41131] ^ n[41132];
assign t[41133] = t[41132] ^ n[41133];
assign t[41134] = t[41133] ^ n[41134];
assign t[41135] = t[41134] ^ n[41135];
assign t[41136] = t[41135] ^ n[41136];
assign t[41137] = t[41136] ^ n[41137];
assign t[41138] = t[41137] ^ n[41138];
assign t[41139] = t[41138] ^ n[41139];
assign t[41140] = t[41139] ^ n[41140];
assign t[41141] = t[41140] ^ n[41141];
assign t[41142] = t[41141] ^ n[41142];
assign t[41143] = t[41142] ^ n[41143];
assign t[41144] = t[41143] ^ n[41144];
assign t[41145] = t[41144] ^ n[41145];
assign t[41146] = t[41145] ^ n[41146];
assign t[41147] = t[41146] ^ n[41147];
assign t[41148] = t[41147] ^ n[41148];
assign t[41149] = t[41148] ^ n[41149];
assign t[41150] = t[41149] ^ n[41150];
assign t[41151] = t[41150] ^ n[41151];
assign t[41152] = t[41151] ^ n[41152];
assign t[41153] = t[41152] ^ n[41153];
assign t[41154] = t[41153] ^ n[41154];
assign t[41155] = t[41154] ^ n[41155];
assign t[41156] = t[41155] ^ n[41156];
assign t[41157] = t[41156] ^ n[41157];
assign t[41158] = t[41157] ^ n[41158];
assign t[41159] = t[41158] ^ n[41159];
assign t[41160] = t[41159] ^ n[41160];
assign t[41161] = t[41160] ^ n[41161];
assign t[41162] = t[41161] ^ n[41162];
assign t[41163] = t[41162] ^ n[41163];
assign t[41164] = t[41163] ^ n[41164];
assign t[41165] = t[41164] ^ n[41165];
assign t[41166] = t[41165] ^ n[41166];
assign t[41167] = t[41166] ^ n[41167];
assign t[41168] = t[41167] ^ n[41168];
assign t[41169] = t[41168] ^ n[41169];
assign t[41170] = t[41169] ^ n[41170];
assign t[41171] = t[41170] ^ n[41171];
assign t[41172] = t[41171] ^ n[41172];
assign t[41173] = t[41172] ^ n[41173];
assign t[41174] = t[41173] ^ n[41174];
assign t[41175] = t[41174] ^ n[41175];
assign t[41176] = t[41175] ^ n[41176];
assign t[41177] = t[41176] ^ n[41177];
assign t[41178] = t[41177] ^ n[41178];
assign t[41179] = t[41178] ^ n[41179];
assign t[41180] = t[41179] ^ n[41180];
assign t[41181] = t[41180] ^ n[41181];
assign t[41182] = t[41181] ^ n[41182];
assign t[41183] = t[41182] ^ n[41183];
assign t[41184] = t[41183] ^ n[41184];
assign t[41185] = t[41184] ^ n[41185];
assign t[41186] = t[41185] ^ n[41186];
assign t[41187] = t[41186] ^ n[41187];
assign t[41188] = t[41187] ^ n[41188];
assign t[41189] = t[41188] ^ n[41189];
assign t[41190] = t[41189] ^ n[41190];
assign t[41191] = t[41190] ^ n[41191];
assign t[41192] = t[41191] ^ n[41192];
assign t[41193] = t[41192] ^ n[41193];
assign t[41194] = t[41193] ^ n[41194];
assign t[41195] = t[41194] ^ n[41195];
assign t[41196] = t[41195] ^ n[41196];
assign t[41197] = t[41196] ^ n[41197];
assign t[41198] = t[41197] ^ n[41198];
assign t[41199] = t[41198] ^ n[41199];
assign t[41200] = t[41199] ^ n[41200];
assign t[41201] = t[41200] ^ n[41201];
assign t[41202] = t[41201] ^ n[41202];
assign t[41203] = t[41202] ^ n[41203];
assign t[41204] = t[41203] ^ n[41204];
assign t[41205] = t[41204] ^ n[41205];
assign t[41206] = t[41205] ^ n[41206];
assign t[41207] = t[41206] ^ n[41207];
assign t[41208] = t[41207] ^ n[41208];
assign t[41209] = t[41208] ^ n[41209];
assign t[41210] = t[41209] ^ n[41210];
assign t[41211] = t[41210] ^ n[41211];
assign t[41212] = t[41211] ^ n[41212];
assign t[41213] = t[41212] ^ n[41213];
assign t[41214] = t[41213] ^ n[41214];
assign t[41215] = t[41214] ^ n[41215];
assign t[41216] = t[41215] ^ n[41216];
assign t[41217] = t[41216] ^ n[41217];
assign t[41218] = t[41217] ^ n[41218];
assign t[41219] = t[41218] ^ n[41219];
assign t[41220] = t[41219] ^ n[41220];
assign t[41221] = t[41220] ^ n[41221];
assign t[41222] = t[41221] ^ n[41222];
assign t[41223] = t[41222] ^ n[41223];
assign t[41224] = t[41223] ^ n[41224];
assign t[41225] = t[41224] ^ n[41225];
assign t[41226] = t[41225] ^ n[41226];
assign t[41227] = t[41226] ^ n[41227];
assign t[41228] = t[41227] ^ n[41228];
assign t[41229] = t[41228] ^ n[41229];
assign t[41230] = t[41229] ^ n[41230];
assign t[41231] = t[41230] ^ n[41231];
assign t[41232] = t[41231] ^ n[41232];
assign t[41233] = t[41232] ^ n[41233];
assign t[41234] = t[41233] ^ n[41234];
assign t[41235] = t[41234] ^ n[41235];
assign t[41236] = t[41235] ^ n[41236];
assign t[41237] = t[41236] ^ n[41237];
assign t[41238] = t[41237] ^ n[41238];
assign t[41239] = t[41238] ^ n[41239];
assign t[41240] = t[41239] ^ n[41240];
assign t[41241] = t[41240] ^ n[41241];
assign t[41242] = t[41241] ^ n[41242];
assign t[41243] = t[41242] ^ n[41243];
assign t[41244] = t[41243] ^ n[41244];
assign t[41245] = t[41244] ^ n[41245];
assign t[41246] = t[41245] ^ n[41246];
assign t[41247] = t[41246] ^ n[41247];
assign t[41248] = t[41247] ^ n[41248];
assign t[41249] = t[41248] ^ n[41249];
assign t[41250] = t[41249] ^ n[41250];
assign t[41251] = t[41250] ^ n[41251];
assign t[41252] = t[41251] ^ n[41252];
assign t[41253] = t[41252] ^ n[41253];
assign t[41254] = t[41253] ^ n[41254];
assign t[41255] = t[41254] ^ n[41255];
assign t[41256] = t[41255] ^ n[41256];
assign t[41257] = t[41256] ^ n[41257];
assign t[41258] = t[41257] ^ n[41258];
assign t[41259] = t[41258] ^ n[41259];
assign t[41260] = t[41259] ^ n[41260];
assign t[41261] = t[41260] ^ n[41261];
assign t[41262] = t[41261] ^ n[41262];
assign t[41263] = t[41262] ^ n[41263];
assign t[41264] = t[41263] ^ n[41264];
assign t[41265] = t[41264] ^ n[41265];
assign t[41266] = t[41265] ^ n[41266];
assign t[41267] = t[41266] ^ n[41267];
assign t[41268] = t[41267] ^ n[41268];
assign t[41269] = t[41268] ^ n[41269];
assign t[41270] = t[41269] ^ n[41270];
assign t[41271] = t[41270] ^ n[41271];
assign t[41272] = t[41271] ^ n[41272];
assign t[41273] = t[41272] ^ n[41273];
assign t[41274] = t[41273] ^ n[41274];
assign t[41275] = t[41274] ^ n[41275];
assign t[41276] = t[41275] ^ n[41276];
assign t[41277] = t[41276] ^ n[41277];
assign t[41278] = t[41277] ^ n[41278];
assign t[41279] = t[41278] ^ n[41279];
assign t[41280] = t[41279] ^ n[41280];
assign t[41281] = t[41280] ^ n[41281];
assign t[41282] = t[41281] ^ n[41282];
assign t[41283] = t[41282] ^ n[41283];
assign t[41284] = t[41283] ^ n[41284];
assign t[41285] = t[41284] ^ n[41285];
assign t[41286] = t[41285] ^ n[41286];
assign t[41287] = t[41286] ^ n[41287];
assign t[41288] = t[41287] ^ n[41288];
assign t[41289] = t[41288] ^ n[41289];
assign t[41290] = t[41289] ^ n[41290];
assign t[41291] = t[41290] ^ n[41291];
assign t[41292] = t[41291] ^ n[41292];
assign t[41293] = t[41292] ^ n[41293];
assign t[41294] = t[41293] ^ n[41294];
assign t[41295] = t[41294] ^ n[41295];
assign t[41296] = t[41295] ^ n[41296];
assign t[41297] = t[41296] ^ n[41297];
assign t[41298] = t[41297] ^ n[41298];
assign t[41299] = t[41298] ^ n[41299];
assign t[41300] = t[41299] ^ n[41300];
assign t[41301] = t[41300] ^ n[41301];
assign t[41302] = t[41301] ^ n[41302];
assign t[41303] = t[41302] ^ n[41303];
assign t[41304] = t[41303] ^ n[41304];
assign t[41305] = t[41304] ^ n[41305];
assign t[41306] = t[41305] ^ n[41306];
assign t[41307] = t[41306] ^ n[41307];
assign t[41308] = t[41307] ^ n[41308];
assign t[41309] = t[41308] ^ n[41309];
assign t[41310] = t[41309] ^ n[41310];
assign t[41311] = t[41310] ^ n[41311];
assign t[41312] = t[41311] ^ n[41312];
assign t[41313] = t[41312] ^ n[41313];
assign t[41314] = t[41313] ^ n[41314];
assign t[41315] = t[41314] ^ n[41315];
assign t[41316] = t[41315] ^ n[41316];
assign t[41317] = t[41316] ^ n[41317];
assign t[41318] = t[41317] ^ n[41318];
assign t[41319] = t[41318] ^ n[41319];
assign t[41320] = t[41319] ^ n[41320];
assign t[41321] = t[41320] ^ n[41321];
assign t[41322] = t[41321] ^ n[41322];
assign t[41323] = t[41322] ^ n[41323];
assign t[41324] = t[41323] ^ n[41324];
assign t[41325] = t[41324] ^ n[41325];
assign t[41326] = t[41325] ^ n[41326];
assign t[41327] = t[41326] ^ n[41327];
assign t[41328] = t[41327] ^ n[41328];
assign t[41329] = t[41328] ^ n[41329];
assign t[41330] = t[41329] ^ n[41330];
assign t[41331] = t[41330] ^ n[41331];
assign t[41332] = t[41331] ^ n[41332];
assign t[41333] = t[41332] ^ n[41333];
assign t[41334] = t[41333] ^ n[41334];
assign t[41335] = t[41334] ^ n[41335];
assign t[41336] = t[41335] ^ n[41336];
assign t[41337] = t[41336] ^ n[41337];
assign t[41338] = t[41337] ^ n[41338];
assign t[41339] = t[41338] ^ n[41339];
assign t[41340] = t[41339] ^ n[41340];
assign t[41341] = t[41340] ^ n[41341];
assign t[41342] = t[41341] ^ n[41342];
assign t[41343] = t[41342] ^ n[41343];
assign t[41344] = t[41343] ^ n[41344];
assign t[41345] = t[41344] ^ n[41345];
assign t[41346] = t[41345] ^ n[41346];
assign t[41347] = t[41346] ^ n[41347];
assign t[41348] = t[41347] ^ n[41348];
assign t[41349] = t[41348] ^ n[41349];
assign t[41350] = t[41349] ^ n[41350];
assign t[41351] = t[41350] ^ n[41351];
assign t[41352] = t[41351] ^ n[41352];
assign t[41353] = t[41352] ^ n[41353];
assign t[41354] = t[41353] ^ n[41354];
assign t[41355] = t[41354] ^ n[41355];
assign t[41356] = t[41355] ^ n[41356];
assign t[41357] = t[41356] ^ n[41357];
assign t[41358] = t[41357] ^ n[41358];
assign t[41359] = t[41358] ^ n[41359];
assign t[41360] = t[41359] ^ n[41360];
assign t[41361] = t[41360] ^ n[41361];
assign t[41362] = t[41361] ^ n[41362];
assign t[41363] = t[41362] ^ n[41363];
assign t[41364] = t[41363] ^ n[41364];
assign t[41365] = t[41364] ^ n[41365];
assign t[41366] = t[41365] ^ n[41366];
assign t[41367] = t[41366] ^ n[41367];
assign t[41368] = t[41367] ^ n[41368];
assign t[41369] = t[41368] ^ n[41369];
assign t[41370] = t[41369] ^ n[41370];
assign t[41371] = t[41370] ^ n[41371];
assign t[41372] = t[41371] ^ n[41372];
assign t[41373] = t[41372] ^ n[41373];
assign t[41374] = t[41373] ^ n[41374];
assign t[41375] = t[41374] ^ n[41375];
assign t[41376] = t[41375] ^ n[41376];
assign t[41377] = t[41376] ^ n[41377];
assign t[41378] = t[41377] ^ n[41378];
assign t[41379] = t[41378] ^ n[41379];
assign t[41380] = t[41379] ^ n[41380];
assign t[41381] = t[41380] ^ n[41381];
assign t[41382] = t[41381] ^ n[41382];
assign t[41383] = t[41382] ^ n[41383];
assign t[41384] = t[41383] ^ n[41384];
assign t[41385] = t[41384] ^ n[41385];
assign t[41386] = t[41385] ^ n[41386];
assign t[41387] = t[41386] ^ n[41387];
assign t[41388] = t[41387] ^ n[41388];
assign t[41389] = t[41388] ^ n[41389];
assign t[41390] = t[41389] ^ n[41390];
assign t[41391] = t[41390] ^ n[41391];
assign t[41392] = t[41391] ^ n[41392];
assign t[41393] = t[41392] ^ n[41393];
assign t[41394] = t[41393] ^ n[41394];
assign t[41395] = t[41394] ^ n[41395];
assign t[41396] = t[41395] ^ n[41396];
assign t[41397] = t[41396] ^ n[41397];
assign t[41398] = t[41397] ^ n[41398];
assign t[41399] = t[41398] ^ n[41399];
assign t[41400] = t[41399] ^ n[41400];
assign t[41401] = t[41400] ^ n[41401];
assign t[41402] = t[41401] ^ n[41402];
assign t[41403] = t[41402] ^ n[41403];
assign t[41404] = t[41403] ^ n[41404];
assign t[41405] = t[41404] ^ n[41405];
assign t[41406] = t[41405] ^ n[41406];
assign t[41407] = t[41406] ^ n[41407];
assign t[41408] = t[41407] ^ n[41408];
assign t[41409] = t[41408] ^ n[41409];
assign t[41410] = t[41409] ^ n[41410];
assign t[41411] = t[41410] ^ n[41411];
assign t[41412] = t[41411] ^ n[41412];
assign t[41413] = t[41412] ^ n[41413];
assign t[41414] = t[41413] ^ n[41414];
assign t[41415] = t[41414] ^ n[41415];
assign t[41416] = t[41415] ^ n[41416];
assign t[41417] = t[41416] ^ n[41417];
assign t[41418] = t[41417] ^ n[41418];
assign t[41419] = t[41418] ^ n[41419];
assign t[41420] = t[41419] ^ n[41420];
assign t[41421] = t[41420] ^ n[41421];
assign t[41422] = t[41421] ^ n[41422];
assign t[41423] = t[41422] ^ n[41423];
assign t[41424] = t[41423] ^ n[41424];
assign t[41425] = t[41424] ^ n[41425];
assign t[41426] = t[41425] ^ n[41426];
assign t[41427] = t[41426] ^ n[41427];
assign t[41428] = t[41427] ^ n[41428];
assign t[41429] = t[41428] ^ n[41429];
assign t[41430] = t[41429] ^ n[41430];
assign t[41431] = t[41430] ^ n[41431];
assign t[41432] = t[41431] ^ n[41432];
assign t[41433] = t[41432] ^ n[41433];
assign t[41434] = t[41433] ^ n[41434];
assign t[41435] = t[41434] ^ n[41435];
assign t[41436] = t[41435] ^ n[41436];
assign t[41437] = t[41436] ^ n[41437];
assign t[41438] = t[41437] ^ n[41438];
assign t[41439] = t[41438] ^ n[41439];
assign t[41440] = t[41439] ^ n[41440];
assign t[41441] = t[41440] ^ n[41441];
assign t[41442] = t[41441] ^ n[41442];
assign t[41443] = t[41442] ^ n[41443];
assign t[41444] = t[41443] ^ n[41444];
assign t[41445] = t[41444] ^ n[41445];
assign t[41446] = t[41445] ^ n[41446];
assign t[41447] = t[41446] ^ n[41447];
assign t[41448] = t[41447] ^ n[41448];
assign t[41449] = t[41448] ^ n[41449];
assign t[41450] = t[41449] ^ n[41450];
assign t[41451] = t[41450] ^ n[41451];
assign t[41452] = t[41451] ^ n[41452];
assign t[41453] = t[41452] ^ n[41453];
assign t[41454] = t[41453] ^ n[41454];
assign t[41455] = t[41454] ^ n[41455];
assign t[41456] = t[41455] ^ n[41456];
assign t[41457] = t[41456] ^ n[41457];
assign t[41458] = t[41457] ^ n[41458];
assign t[41459] = t[41458] ^ n[41459];
assign t[41460] = t[41459] ^ n[41460];
assign t[41461] = t[41460] ^ n[41461];
assign t[41462] = t[41461] ^ n[41462];
assign t[41463] = t[41462] ^ n[41463];
assign t[41464] = t[41463] ^ n[41464];
assign t[41465] = t[41464] ^ n[41465];
assign t[41466] = t[41465] ^ n[41466];
assign t[41467] = t[41466] ^ n[41467];
assign t[41468] = t[41467] ^ n[41468];
assign t[41469] = t[41468] ^ n[41469];
assign t[41470] = t[41469] ^ n[41470];
assign t[41471] = t[41470] ^ n[41471];
assign t[41472] = t[41471] ^ n[41472];
assign t[41473] = t[41472] ^ n[41473];
assign t[41474] = t[41473] ^ n[41474];
assign t[41475] = t[41474] ^ n[41475];
assign t[41476] = t[41475] ^ n[41476];
assign t[41477] = t[41476] ^ n[41477];
assign t[41478] = t[41477] ^ n[41478];
assign t[41479] = t[41478] ^ n[41479];
assign t[41480] = t[41479] ^ n[41480];
assign t[41481] = t[41480] ^ n[41481];
assign t[41482] = t[41481] ^ n[41482];
assign t[41483] = t[41482] ^ n[41483];
assign t[41484] = t[41483] ^ n[41484];
assign t[41485] = t[41484] ^ n[41485];
assign t[41486] = t[41485] ^ n[41486];
assign t[41487] = t[41486] ^ n[41487];
assign t[41488] = t[41487] ^ n[41488];
assign t[41489] = t[41488] ^ n[41489];
assign t[41490] = t[41489] ^ n[41490];
assign t[41491] = t[41490] ^ n[41491];
assign t[41492] = t[41491] ^ n[41492];
assign t[41493] = t[41492] ^ n[41493];
assign t[41494] = t[41493] ^ n[41494];
assign t[41495] = t[41494] ^ n[41495];
assign t[41496] = t[41495] ^ n[41496];
assign t[41497] = t[41496] ^ n[41497];
assign t[41498] = t[41497] ^ n[41498];
assign t[41499] = t[41498] ^ n[41499];
assign t[41500] = t[41499] ^ n[41500];
assign t[41501] = t[41500] ^ n[41501];
assign t[41502] = t[41501] ^ n[41502];
assign t[41503] = t[41502] ^ n[41503];
assign t[41504] = t[41503] ^ n[41504];
assign t[41505] = t[41504] ^ n[41505];
assign t[41506] = t[41505] ^ n[41506];
assign t[41507] = t[41506] ^ n[41507];
assign t[41508] = t[41507] ^ n[41508];
assign t[41509] = t[41508] ^ n[41509];
assign t[41510] = t[41509] ^ n[41510];
assign t[41511] = t[41510] ^ n[41511];
assign t[41512] = t[41511] ^ n[41512];
assign t[41513] = t[41512] ^ n[41513];
assign t[41514] = t[41513] ^ n[41514];
assign t[41515] = t[41514] ^ n[41515];
assign t[41516] = t[41515] ^ n[41516];
assign t[41517] = t[41516] ^ n[41517];
assign t[41518] = t[41517] ^ n[41518];
assign t[41519] = t[41518] ^ n[41519];
assign t[41520] = t[41519] ^ n[41520];
assign t[41521] = t[41520] ^ n[41521];
assign t[41522] = t[41521] ^ n[41522];
assign t[41523] = t[41522] ^ n[41523];
assign t[41524] = t[41523] ^ n[41524];
assign t[41525] = t[41524] ^ n[41525];
assign t[41526] = t[41525] ^ n[41526];
assign t[41527] = t[41526] ^ n[41527];
assign t[41528] = t[41527] ^ n[41528];
assign t[41529] = t[41528] ^ n[41529];
assign t[41530] = t[41529] ^ n[41530];
assign t[41531] = t[41530] ^ n[41531];
assign t[41532] = t[41531] ^ n[41532];
assign t[41533] = t[41532] ^ n[41533];
assign t[41534] = t[41533] ^ n[41534];
assign t[41535] = t[41534] ^ n[41535];
assign t[41536] = t[41535] ^ n[41536];
assign t[41537] = t[41536] ^ n[41537];
assign t[41538] = t[41537] ^ n[41538];
assign t[41539] = t[41538] ^ n[41539];
assign t[41540] = t[41539] ^ n[41540];
assign t[41541] = t[41540] ^ n[41541];
assign t[41542] = t[41541] ^ n[41542];
assign t[41543] = t[41542] ^ n[41543];
assign t[41544] = t[41543] ^ n[41544];
assign t[41545] = t[41544] ^ n[41545];
assign t[41546] = t[41545] ^ n[41546];
assign t[41547] = t[41546] ^ n[41547];
assign t[41548] = t[41547] ^ n[41548];
assign t[41549] = t[41548] ^ n[41549];
assign t[41550] = t[41549] ^ n[41550];
assign t[41551] = t[41550] ^ n[41551];
assign t[41552] = t[41551] ^ n[41552];
assign t[41553] = t[41552] ^ n[41553];
assign t[41554] = t[41553] ^ n[41554];
assign t[41555] = t[41554] ^ n[41555];
assign t[41556] = t[41555] ^ n[41556];
assign t[41557] = t[41556] ^ n[41557];
assign t[41558] = t[41557] ^ n[41558];
assign t[41559] = t[41558] ^ n[41559];
assign t[41560] = t[41559] ^ n[41560];
assign t[41561] = t[41560] ^ n[41561];
assign t[41562] = t[41561] ^ n[41562];
assign t[41563] = t[41562] ^ n[41563];
assign t[41564] = t[41563] ^ n[41564];
assign t[41565] = t[41564] ^ n[41565];
assign t[41566] = t[41565] ^ n[41566];
assign t[41567] = t[41566] ^ n[41567];
assign t[41568] = t[41567] ^ n[41568];
assign t[41569] = t[41568] ^ n[41569];
assign t[41570] = t[41569] ^ n[41570];
assign t[41571] = t[41570] ^ n[41571];
assign t[41572] = t[41571] ^ n[41572];
assign t[41573] = t[41572] ^ n[41573];
assign t[41574] = t[41573] ^ n[41574];
assign t[41575] = t[41574] ^ n[41575];
assign t[41576] = t[41575] ^ n[41576];
assign t[41577] = t[41576] ^ n[41577];
assign t[41578] = t[41577] ^ n[41578];
assign t[41579] = t[41578] ^ n[41579];
assign t[41580] = t[41579] ^ n[41580];
assign t[41581] = t[41580] ^ n[41581];
assign t[41582] = t[41581] ^ n[41582];
assign t[41583] = t[41582] ^ n[41583];
assign t[41584] = t[41583] ^ n[41584];
assign t[41585] = t[41584] ^ n[41585];
assign t[41586] = t[41585] ^ n[41586];
assign t[41587] = t[41586] ^ n[41587];
assign t[41588] = t[41587] ^ n[41588];
assign t[41589] = t[41588] ^ n[41589];
assign t[41590] = t[41589] ^ n[41590];
assign t[41591] = t[41590] ^ n[41591];
assign t[41592] = t[41591] ^ n[41592];
assign t[41593] = t[41592] ^ n[41593];
assign t[41594] = t[41593] ^ n[41594];
assign t[41595] = t[41594] ^ n[41595];
assign t[41596] = t[41595] ^ n[41596];
assign t[41597] = t[41596] ^ n[41597];
assign t[41598] = t[41597] ^ n[41598];
assign t[41599] = t[41598] ^ n[41599];
assign t[41600] = t[41599] ^ n[41600];
assign t[41601] = t[41600] ^ n[41601];
assign t[41602] = t[41601] ^ n[41602];
assign t[41603] = t[41602] ^ n[41603];
assign t[41604] = t[41603] ^ n[41604];
assign t[41605] = t[41604] ^ n[41605];
assign t[41606] = t[41605] ^ n[41606];
assign t[41607] = t[41606] ^ n[41607];
assign t[41608] = t[41607] ^ n[41608];
assign t[41609] = t[41608] ^ n[41609];
assign t[41610] = t[41609] ^ n[41610];
assign t[41611] = t[41610] ^ n[41611];
assign t[41612] = t[41611] ^ n[41612];
assign t[41613] = t[41612] ^ n[41613];
assign t[41614] = t[41613] ^ n[41614];
assign t[41615] = t[41614] ^ n[41615];
assign t[41616] = t[41615] ^ n[41616];
assign t[41617] = t[41616] ^ n[41617];
assign t[41618] = t[41617] ^ n[41618];
assign t[41619] = t[41618] ^ n[41619];
assign t[41620] = t[41619] ^ n[41620];
assign t[41621] = t[41620] ^ n[41621];
assign t[41622] = t[41621] ^ n[41622];
assign t[41623] = t[41622] ^ n[41623];
assign t[41624] = t[41623] ^ n[41624];
assign t[41625] = t[41624] ^ n[41625];
assign t[41626] = t[41625] ^ n[41626];
assign t[41627] = t[41626] ^ n[41627];
assign t[41628] = t[41627] ^ n[41628];
assign t[41629] = t[41628] ^ n[41629];
assign t[41630] = t[41629] ^ n[41630];
assign t[41631] = t[41630] ^ n[41631];
assign t[41632] = t[41631] ^ n[41632];
assign t[41633] = t[41632] ^ n[41633];
assign t[41634] = t[41633] ^ n[41634];
assign t[41635] = t[41634] ^ n[41635];
assign t[41636] = t[41635] ^ n[41636];
assign t[41637] = t[41636] ^ n[41637];
assign t[41638] = t[41637] ^ n[41638];
assign t[41639] = t[41638] ^ n[41639];
assign t[41640] = t[41639] ^ n[41640];
assign t[41641] = t[41640] ^ n[41641];
assign t[41642] = t[41641] ^ n[41642];
assign t[41643] = t[41642] ^ n[41643];
assign t[41644] = t[41643] ^ n[41644];
assign t[41645] = t[41644] ^ n[41645];
assign t[41646] = t[41645] ^ n[41646];
assign t[41647] = t[41646] ^ n[41647];
assign t[41648] = t[41647] ^ n[41648];
assign t[41649] = t[41648] ^ n[41649];
assign t[41650] = t[41649] ^ n[41650];
assign t[41651] = t[41650] ^ n[41651];
assign t[41652] = t[41651] ^ n[41652];
assign t[41653] = t[41652] ^ n[41653];
assign t[41654] = t[41653] ^ n[41654];
assign t[41655] = t[41654] ^ n[41655];
assign t[41656] = t[41655] ^ n[41656];
assign t[41657] = t[41656] ^ n[41657];
assign t[41658] = t[41657] ^ n[41658];
assign t[41659] = t[41658] ^ n[41659];
assign t[41660] = t[41659] ^ n[41660];
assign t[41661] = t[41660] ^ n[41661];
assign t[41662] = t[41661] ^ n[41662];
assign t[41663] = t[41662] ^ n[41663];
assign t[41664] = t[41663] ^ n[41664];
assign t[41665] = t[41664] ^ n[41665];
assign t[41666] = t[41665] ^ n[41666];
assign t[41667] = t[41666] ^ n[41667];
assign t[41668] = t[41667] ^ n[41668];
assign t[41669] = t[41668] ^ n[41669];
assign t[41670] = t[41669] ^ n[41670];
assign t[41671] = t[41670] ^ n[41671];
assign t[41672] = t[41671] ^ n[41672];
assign t[41673] = t[41672] ^ n[41673];
assign t[41674] = t[41673] ^ n[41674];
assign t[41675] = t[41674] ^ n[41675];
assign t[41676] = t[41675] ^ n[41676];
assign t[41677] = t[41676] ^ n[41677];
assign t[41678] = t[41677] ^ n[41678];
assign t[41679] = t[41678] ^ n[41679];
assign t[41680] = t[41679] ^ n[41680];
assign t[41681] = t[41680] ^ n[41681];
assign t[41682] = t[41681] ^ n[41682];
assign t[41683] = t[41682] ^ n[41683];
assign t[41684] = t[41683] ^ n[41684];
assign t[41685] = t[41684] ^ n[41685];
assign t[41686] = t[41685] ^ n[41686];
assign t[41687] = t[41686] ^ n[41687];
assign t[41688] = t[41687] ^ n[41688];
assign t[41689] = t[41688] ^ n[41689];
assign t[41690] = t[41689] ^ n[41690];
assign t[41691] = t[41690] ^ n[41691];
assign t[41692] = t[41691] ^ n[41692];
assign t[41693] = t[41692] ^ n[41693];
assign t[41694] = t[41693] ^ n[41694];
assign t[41695] = t[41694] ^ n[41695];
assign t[41696] = t[41695] ^ n[41696];
assign t[41697] = t[41696] ^ n[41697];
assign t[41698] = t[41697] ^ n[41698];
assign t[41699] = t[41698] ^ n[41699];
assign t[41700] = t[41699] ^ n[41700];
assign t[41701] = t[41700] ^ n[41701];
assign t[41702] = t[41701] ^ n[41702];
assign t[41703] = t[41702] ^ n[41703];
assign t[41704] = t[41703] ^ n[41704];
assign t[41705] = t[41704] ^ n[41705];
assign t[41706] = t[41705] ^ n[41706];
assign t[41707] = t[41706] ^ n[41707];
assign t[41708] = t[41707] ^ n[41708];
assign t[41709] = t[41708] ^ n[41709];
assign t[41710] = t[41709] ^ n[41710];
assign t[41711] = t[41710] ^ n[41711];
assign t[41712] = t[41711] ^ n[41712];
assign t[41713] = t[41712] ^ n[41713];
assign t[41714] = t[41713] ^ n[41714];
assign t[41715] = t[41714] ^ n[41715];
assign t[41716] = t[41715] ^ n[41716];
assign t[41717] = t[41716] ^ n[41717];
assign t[41718] = t[41717] ^ n[41718];
assign t[41719] = t[41718] ^ n[41719];
assign t[41720] = t[41719] ^ n[41720];
assign t[41721] = t[41720] ^ n[41721];
assign t[41722] = t[41721] ^ n[41722];
assign t[41723] = t[41722] ^ n[41723];
assign t[41724] = t[41723] ^ n[41724];
assign t[41725] = t[41724] ^ n[41725];
assign t[41726] = t[41725] ^ n[41726];
assign t[41727] = t[41726] ^ n[41727];
assign t[41728] = t[41727] ^ n[41728];
assign t[41729] = t[41728] ^ n[41729];
assign t[41730] = t[41729] ^ n[41730];
assign t[41731] = t[41730] ^ n[41731];
assign t[41732] = t[41731] ^ n[41732];
assign t[41733] = t[41732] ^ n[41733];
assign t[41734] = t[41733] ^ n[41734];
assign t[41735] = t[41734] ^ n[41735];
assign t[41736] = t[41735] ^ n[41736];
assign t[41737] = t[41736] ^ n[41737];
assign t[41738] = t[41737] ^ n[41738];
assign t[41739] = t[41738] ^ n[41739];
assign t[41740] = t[41739] ^ n[41740];
assign t[41741] = t[41740] ^ n[41741];
assign t[41742] = t[41741] ^ n[41742];
assign t[41743] = t[41742] ^ n[41743];
assign t[41744] = t[41743] ^ n[41744];
assign t[41745] = t[41744] ^ n[41745];
assign t[41746] = t[41745] ^ n[41746];
assign t[41747] = t[41746] ^ n[41747];
assign t[41748] = t[41747] ^ n[41748];
assign t[41749] = t[41748] ^ n[41749];
assign t[41750] = t[41749] ^ n[41750];
assign t[41751] = t[41750] ^ n[41751];
assign t[41752] = t[41751] ^ n[41752];
assign t[41753] = t[41752] ^ n[41753];
assign t[41754] = t[41753] ^ n[41754];
assign t[41755] = t[41754] ^ n[41755];
assign t[41756] = t[41755] ^ n[41756];
assign t[41757] = t[41756] ^ n[41757];
assign t[41758] = t[41757] ^ n[41758];
assign t[41759] = t[41758] ^ n[41759];
assign t[41760] = t[41759] ^ n[41760];
assign t[41761] = t[41760] ^ n[41761];
assign t[41762] = t[41761] ^ n[41762];
assign t[41763] = t[41762] ^ n[41763];
assign t[41764] = t[41763] ^ n[41764];
assign t[41765] = t[41764] ^ n[41765];
assign t[41766] = t[41765] ^ n[41766];
assign t[41767] = t[41766] ^ n[41767];
assign t[41768] = t[41767] ^ n[41768];
assign t[41769] = t[41768] ^ n[41769];
assign t[41770] = t[41769] ^ n[41770];
assign t[41771] = t[41770] ^ n[41771];
assign t[41772] = t[41771] ^ n[41772];
assign t[41773] = t[41772] ^ n[41773];
assign t[41774] = t[41773] ^ n[41774];
assign t[41775] = t[41774] ^ n[41775];
assign t[41776] = t[41775] ^ n[41776];
assign t[41777] = t[41776] ^ n[41777];
assign t[41778] = t[41777] ^ n[41778];
assign t[41779] = t[41778] ^ n[41779];
assign t[41780] = t[41779] ^ n[41780];
assign t[41781] = t[41780] ^ n[41781];
assign t[41782] = t[41781] ^ n[41782];
assign t[41783] = t[41782] ^ n[41783];
assign t[41784] = t[41783] ^ n[41784];
assign t[41785] = t[41784] ^ n[41785];
assign t[41786] = t[41785] ^ n[41786];
assign t[41787] = t[41786] ^ n[41787];
assign t[41788] = t[41787] ^ n[41788];
assign t[41789] = t[41788] ^ n[41789];
assign t[41790] = t[41789] ^ n[41790];
assign t[41791] = t[41790] ^ n[41791];
assign t[41792] = t[41791] ^ n[41792];
assign t[41793] = t[41792] ^ n[41793];
assign t[41794] = t[41793] ^ n[41794];
assign t[41795] = t[41794] ^ n[41795];
assign t[41796] = t[41795] ^ n[41796];
assign t[41797] = t[41796] ^ n[41797];
assign t[41798] = t[41797] ^ n[41798];
assign t[41799] = t[41798] ^ n[41799];
assign t[41800] = t[41799] ^ n[41800];
assign t[41801] = t[41800] ^ n[41801];
assign t[41802] = t[41801] ^ n[41802];
assign t[41803] = t[41802] ^ n[41803];
assign t[41804] = t[41803] ^ n[41804];
assign t[41805] = t[41804] ^ n[41805];
assign t[41806] = t[41805] ^ n[41806];
assign t[41807] = t[41806] ^ n[41807];
assign t[41808] = t[41807] ^ n[41808];
assign t[41809] = t[41808] ^ n[41809];
assign t[41810] = t[41809] ^ n[41810];
assign t[41811] = t[41810] ^ n[41811];
assign t[41812] = t[41811] ^ n[41812];
assign t[41813] = t[41812] ^ n[41813];
assign t[41814] = t[41813] ^ n[41814];
assign t[41815] = t[41814] ^ n[41815];
assign t[41816] = t[41815] ^ n[41816];
assign t[41817] = t[41816] ^ n[41817];
assign t[41818] = t[41817] ^ n[41818];
assign t[41819] = t[41818] ^ n[41819];
assign t[41820] = t[41819] ^ n[41820];
assign t[41821] = t[41820] ^ n[41821];
assign t[41822] = t[41821] ^ n[41822];
assign t[41823] = t[41822] ^ n[41823];
assign t[41824] = t[41823] ^ n[41824];
assign t[41825] = t[41824] ^ n[41825];
assign t[41826] = t[41825] ^ n[41826];
assign t[41827] = t[41826] ^ n[41827];
assign t[41828] = t[41827] ^ n[41828];
assign t[41829] = t[41828] ^ n[41829];
assign t[41830] = t[41829] ^ n[41830];
assign t[41831] = t[41830] ^ n[41831];
assign t[41832] = t[41831] ^ n[41832];
assign t[41833] = t[41832] ^ n[41833];
assign t[41834] = t[41833] ^ n[41834];
assign t[41835] = t[41834] ^ n[41835];
assign t[41836] = t[41835] ^ n[41836];
assign t[41837] = t[41836] ^ n[41837];
assign t[41838] = t[41837] ^ n[41838];
assign t[41839] = t[41838] ^ n[41839];
assign t[41840] = t[41839] ^ n[41840];
assign t[41841] = t[41840] ^ n[41841];
assign t[41842] = t[41841] ^ n[41842];
assign t[41843] = t[41842] ^ n[41843];
assign t[41844] = t[41843] ^ n[41844];
assign t[41845] = t[41844] ^ n[41845];
assign t[41846] = t[41845] ^ n[41846];
assign t[41847] = t[41846] ^ n[41847];
assign t[41848] = t[41847] ^ n[41848];
assign t[41849] = t[41848] ^ n[41849];
assign t[41850] = t[41849] ^ n[41850];
assign t[41851] = t[41850] ^ n[41851];
assign t[41852] = t[41851] ^ n[41852];
assign t[41853] = t[41852] ^ n[41853];
assign t[41854] = t[41853] ^ n[41854];
assign t[41855] = t[41854] ^ n[41855];
assign t[41856] = t[41855] ^ n[41856];
assign t[41857] = t[41856] ^ n[41857];
assign t[41858] = t[41857] ^ n[41858];
assign t[41859] = t[41858] ^ n[41859];
assign t[41860] = t[41859] ^ n[41860];
assign t[41861] = t[41860] ^ n[41861];
assign t[41862] = t[41861] ^ n[41862];
assign t[41863] = t[41862] ^ n[41863];
assign t[41864] = t[41863] ^ n[41864];
assign t[41865] = t[41864] ^ n[41865];
assign t[41866] = t[41865] ^ n[41866];
assign t[41867] = t[41866] ^ n[41867];
assign t[41868] = t[41867] ^ n[41868];
assign t[41869] = t[41868] ^ n[41869];
assign t[41870] = t[41869] ^ n[41870];
assign t[41871] = t[41870] ^ n[41871];
assign t[41872] = t[41871] ^ n[41872];
assign t[41873] = t[41872] ^ n[41873];
assign t[41874] = t[41873] ^ n[41874];
assign t[41875] = t[41874] ^ n[41875];
assign t[41876] = t[41875] ^ n[41876];
assign t[41877] = t[41876] ^ n[41877];
assign t[41878] = t[41877] ^ n[41878];
assign t[41879] = t[41878] ^ n[41879];
assign t[41880] = t[41879] ^ n[41880];
assign t[41881] = t[41880] ^ n[41881];
assign t[41882] = t[41881] ^ n[41882];
assign t[41883] = t[41882] ^ n[41883];
assign t[41884] = t[41883] ^ n[41884];
assign t[41885] = t[41884] ^ n[41885];
assign t[41886] = t[41885] ^ n[41886];
assign t[41887] = t[41886] ^ n[41887];
assign t[41888] = t[41887] ^ n[41888];
assign t[41889] = t[41888] ^ n[41889];
assign t[41890] = t[41889] ^ n[41890];
assign t[41891] = t[41890] ^ n[41891];
assign t[41892] = t[41891] ^ n[41892];
assign t[41893] = t[41892] ^ n[41893];
assign t[41894] = t[41893] ^ n[41894];
assign t[41895] = t[41894] ^ n[41895];
assign t[41896] = t[41895] ^ n[41896];
assign t[41897] = t[41896] ^ n[41897];
assign t[41898] = t[41897] ^ n[41898];
assign t[41899] = t[41898] ^ n[41899];
assign t[41900] = t[41899] ^ n[41900];
assign t[41901] = t[41900] ^ n[41901];
assign t[41902] = t[41901] ^ n[41902];
assign t[41903] = t[41902] ^ n[41903];
assign t[41904] = t[41903] ^ n[41904];
assign t[41905] = t[41904] ^ n[41905];
assign t[41906] = t[41905] ^ n[41906];
assign t[41907] = t[41906] ^ n[41907];
assign t[41908] = t[41907] ^ n[41908];
assign t[41909] = t[41908] ^ n[41909];
assign t[41910] = t[41909] ^ n[41910];
assign t[41911] = t[41910] ^ n[41911];
assign t[41912] = t[41911] ^ n[41912];
assign t[41913] = t[41912] ^ n[41913];
assign t[41914] = t[41913] ^ n[41914];
assign t[41915] = t[41914] ^ n[41915];
assign t[41916] = t[41915] ^ n[41916];
assign t[41917] = t[41916] ^ n[41917];
assign t[41918] = t[41917] ^ n[41918];
assign t[41919] = t[41918] ^ n[41919];
assign t[41920] = t[41919] ^ n[41920];
assign t[41921] = t[41920] ^ n[41921];
assign t[41922] = t[41921] ^ n[41922];
assign t[41923] = t[41922] ^ n[41923];
assign t[41924] = t[41923] ^ n[41924];
assign t[41925] = t[41924] ^ n[41925];
assign t[41926] = t[41925] ^ n[41926];
assign t[41927] = t[41926] ^ n[41927];
assign t[41928] = t[41927] ^ n[41928];
assign t[41929] = t[41928] ^ n[41929];
assign t[41930] = t[41929] ^ n[41930];
assign t[41931] = t[41930] ^ n[41931];
assign t[41932] = t[41931] ^ n[41932];
assign t[41933] = t[41932] ^ n[41933];
assign t[41934] = t[41933] ^ n[41934];
assign t[41935] = t[41934] ^ n[41935];
assign t[41936] = t[41935] ^ n[41936];
assign t[41937] = t[41936] ^ n[41937];
assign t[41938] = t[41937] ^ n[41938];
assign t[41939] = t[41938] ^ n[41939];
assign t[41940] = t[41939] ^ n[41940];
assign t[41941] = t[41940] ^ n[41941];
assign t[41942] = t[41941] ^ n[41942];
assign t[41943] = t[41942] ^ n[41943];
assign t[41944] = t[41943] ^ n[41944];
assign t[41945] = t[41944] ^ n[41945];
assign t[41946] = t[41945] ^ n[41946];
assign t[41947] = t[41946] ^ n[41947];
assign t[41948] = t[41947] ^ n[41948];
assign t[41949] = t[41948] ^ n[41949];
assign t[41950] = t[41949] ^ n[41950];
assign t[41951] = t[41950] ^ n[41951];
assign t[41952] = t[41951] ^ n[41952];
assign t[41953] = t[41952] ^ n[41953];
assign t[41954] = t[41953] ^ n[41954];
assign t[41955] = t[41954] ^ n[41955];
assign t[41956] = t[41955] ^ n[41956];
assign t[41957] = t[41956] ^ n[41957];
assign t[41958] = t[41957] ^ n[41958];
assign t[41959] = t[41958] ^ n[41959];
assign t[41960] = t[41959] ^ n[41960];
assign t[41961] = t[41960] ^ n[41961];
assign t[41962] = t[41961] ^ n[41962];
assign t[41963] = t[41962] ^ n[41963];
assign t[41964] = t[41963] ^ n[41964];
assign t[41965] = t[41964] ^ n[41965];
assign t[41966] = t[41965] ^ n[41966];
assign t[41967] = t[41966] ^ n[41967];
assign t[41968] = t[41967] ^ n[41968];
assign t[41969] = t[41968] ^ n[41969];
assign t[41970] = t[41969] ^ n[41970];
assign t[41971] = t[41970] ^ n[41971];
assign t[41972] = t[41971] ^ n[41972];
assign t[41973] = t[41972] ^ n[41973];
assign t[41974] = t[41973] ^ n[41974];
assign t[41975] = t[41974] ^ n[41975];
assign t[41976] = t[41975] ^ n[41976];
assign t[41977] = t[41976] ^ n[41977];
assign t[41978] = t[41977] ^ n[41978];
assign t[41979] = t[41978] ^ n[41979];
assign t[41980] = t[41979] ^ n[41980];
assign t[41981] = t[41980] ^ n[41981];
assign t[41982] = t[41981] ^ n[41982];
assign t[41983] = t[41982] ^ n[41983];
assign t[41984] = t[41983] ^ n[41984];
assign t[41985] = t[41984] ^ n[41985];
assign t[41986] = t[41985] ^ n[41986];
assign t[41987] = t[41986] ^ n[41987];
assign t[41988] = t[41987] ^ n[41988];
assign t[41989] = t[41988] ^ n[41989];
assign t[41990] = t[41989] ^ n[41990];
assign t[41991] = t[41990] ^ n[41991];
assign t[41992] = t[41991] ^ n[41992];
assign t[41993] = t[41992] ^ n[41993];
assign t[41994] = t[41993] ^ n[41994];
assign t[41995] = t[41994] ^ n[41995];
assign t[41996] = t[41995] ^ n[41996];
assign t[41997] = t[41996] ^ n[41997];
assign t[41998] = t[41997] ^ n[41998];
assign t[41999] = t[41998] ^ n[41999];
assign t[42000] = t[41999] ^ n[42000];
assign t[42001] = t[42000] ^ n[42001];
assign t[42002] = t[42001] ^ n[42002];
assign t[42003] = t[42002] ^ n[42003];
assign t[42004] = t[42003] ^ n[42004];
assign t[42005] = t[42004] ^ n[42005];
assign t[42006] = t[42005] ^ n[42006];
assign t[42007] = t[42006] ^ n[42007];
assign t[42008] = t[42007] ^ n[42008];
assign t[42009] = t[42008] ^ n[42009];
assign t[42010] = t[42009] ^ n[42010];
assign t[42011] = t[42010] ^ n[42011];
assign t[42012] = t[42011] ^ n[42012];
assign t[42013] = t[42012] ^ n[42013];
assign t[42014] = t[42013] ^ n[42014];
assign t[42015] = t[42014] ^ n[42015];
assign t[42016] = t[42015] ^ n[42016];
assign t[42017] = t[42016] ^ n[42017];
assign t[42018] = t[42017] ^ n[42018];
assign t[42019] = t[42018] ^ n[42019];
assign t[42020] = t[42019] ^ n[42020];
assign t[42021] = t[42020] ^ n[42021];
assign t[42022] = t[42021] ^ n[42022];
assign t[42023] = t[42022] ^ n[42023];
assign t[42024] = t[42023] ^ n[42024];
assign t[42025] = t[42024] ^ n[42025];
assign t[42026] = t[42025] ^ n[42026];
assign t[42027] = t[42026] ^ n[42027];
assign t[42028] = t[42027] ^ n[42028];
assign t[42029] = t[42028] ^ n[42029];
assign t[42030] = t[42029] ^ n[42030];
assign t[42031] = t[42030] ^ n[42031];
assign t[42032] = t[42031] ^ n[42032];
assign t[42033] = t[42032] ^ n[42033];
assign t[42034] = t[42033] ^ n[42034];
assign t[42035] = t[42034] ^ n[42035];
assign t[42036] = t[42035] ^ n[42036];
assign t[42037] = t[42036] ^ n[42037];
assign t[42038] = t[42037] ^ n[42038];
assign t[42039] = t[42038] ^ n[42039];
assign t[42040] = t[42039] ^ n[42040];
assign t[42041] = t[42040] ^ n[42041];
assign t[42042] = t[42041] ^ n[42042];
assign t[42043] = t[42042] ^ n[42043];
assign t[42044] = t[42043] ^ n[42044];
assign t[42045] = t[42044] ^ n[42045];
assign t[42046] = t[42045] ^ n[42046];
assign t[42047] = t[42046] ^ n[42047];
assign t[42048] = t[42047] ^ n[42048];
assign t[42049] = t[42048] ^ n[42049];
assign t[42050] = t[42049] ^ n[42050];
assign t[42051] = t[42050] ^ n[42051];
assign t[42052] = t[42051] ^ n[42052];
assign t[42053] = t[42052] ^ n[42053];
assign t[42054] = t[42053] ^ n[42054];
assign t[42055] = t[42054] ^ n[42055];
assign t[42056] = t[42055] ^ n[42056];
assign t[42057] = t[42056] ^ n[42057];
assign t[42058] = t[42057] ^ n[42058];
assign t[42059] = t[42058] ^ n[42059];
assign t[42060] = t[42059] ^ n[42060];
assign t[42061] = t[42060] ^ n[42061];
assign t[42062] = t[42061] ^ n[42062];
assign t[42063] = t[42062] ^ n[42063];
assign t[42064] = t[42063] ^ n[42064];
assign t[42065] = t[42064] ^ n[42065];
assign t[42066] = t[42065] ^ n[42066];
assign t[42067] = t[42066] ^ n[42067];
assign t[42068] = t[42067] ^ n[42068];
assign t[42069] = t[42068] ^ n[42069];
assign t[42070] = t[42069] ^ n[42070];
assign t[42071] = t[42070] ^ n[42071];
assign t[42072] = t[42071] ^ n[42072];
assign t[42073] = t[42072] ^ n[42073];
assign t[42074] = t[42073] ^ n[42074];
assign t[42075] = t[42074] ^ n[42075];
assign t[42076] = t[42075] ^ n[42076];
assign t[42077] = t[42076] ^ n[42077];
assign t[42078] = t[42077] ^ n[42078];
assign t[42079] = t[42078] ^ n[42079];
assign t[42080] = t[42079] ^ n[42080];
assign t[42081] = t[42080] ^ n[42081];
assign t[42082] = t[42081] ^ n[42082];
assign t[42083] = t[42082] ^ n[42083];
assign t[42084] = t[42083] ^ n[42084];
assign t[42085] = t[42084] ^ n[42085];
assign t[42086] = t[42085] ^ n[42086];
assign t[42087] = t[42086] ^ n[42087];
assign t[42088] = t[42087] ^ n[42088];
assign t[42089] = t[42088] ^ n[42089];
assign t[42090] = t[42089] ^ n[42090];
assign t[42091] = t[42090] ^ n[42091];
assign t[42092] = t[42091] ^ n[42092];
assign t[42093] = t[42092] ^ n[42093];
assign t[42094] = t[42093] ^ n[42094];
assign t[42095] = t[42094] ^ n[42095];
assign t[42096] = t[42095] ^ n[42096];
assign t[42097] = t[42096] ^ n[42097];
assign t[42098] = t[42097] ^ n[42098];
assign t[42099] = t[42098] ^ n[42099];
assign t[42100] = t[42099] ^ n[42100];
assign t[42101] = t[42100] ^ n[42101];
assign t[42102] = t[42101] ^ n[42102];
assign t[42103] = t[42102] ^ n[42103];
assign t[42104] = t[42103] ^ n[42104];
assign t[42105] = t[42104] ^ n[42105];
assign t[42106] = t[42105] ^ n[42106];
assign t[42107] = t[42106] ^ n[42107];
assign t[42108] = t[42107] ^ n[42108];
assign t[42109] = t[42108] ^ n[42109];
assign t[42110] = t[42109] ^ n[42110];
assign t[42111] = t[42110] ^ n[42111];
assign t[42112] = t[42111] ^ n[42112];
assign t[42113] = t[42112] ^ n[42113];
assign t[42114] = t[42113] ^ n[42114];
assign t[42115] = t[42114] ^ n[42115];
assign t[42116] = t[42115] ^ n[42116];
assign t[42117] = t[42116] ^ n[42117];
assign t[42118] = t[42117] ^ n[42118];
assign t[42119] = t[42118] ^ n[42119];
assign t[42120] = t[42119] ^ n[42120];
assign t[42121] = t[42120] ^ n[42121];
assign t[42122] = t[42121] ^ n[42122];
assign t[42123] = t[42122] ^ n[42123];
assign t[42124] = t[42123] ^ n[42124];
assign t[42125] = t[42124] ^ n[42125];
assign t[42126] = t[42125] ^ n[42126];
assign t[42127] = t[42126] ^ n[42127];
assign t[42128] = t[42127] ^ n[42128];
assign t[42129] = t[42128] ^ n[42129];
assign t[42130] = t[42129] ^ n[42130];
assign t[42131] = t[42130] ^ n[42131];
assign t[42132] = t[42131] ^ n[42132];
assign t[42133] = t[42132] ^ n[42133];
assign t[42134] = t[42133] ^ n[42134];
assign t[42135] = t[42134] ^ n[42135];
assign t[42136] = t[42135] ^ n[42136];
assign t[42137] = t[42136] ^ n[42137];
assign t[42138] = t[42137] ^ n[42138];
assign t[42139] = t[42138] ^ n[42139];
assign t[42140] = t[42139] ^ n[42140];
assign t[42141] = t[42140] ^ n[42141];
assign t[42142] = t[42141] ^ n[42142];
assign t[42143] = t[42142] ^ n[42143];
assign t[42144] = t[42143] ^ n[42144];
assign t[42145] = t[42144] ^ n[42145];
assign t[42146] = t[42145] ^ n[42146];
assign t[42147] = t[42146] ^ n[42147];
assign t[42148] = t[42147] ^ n[42148];
assign t[42149] = t[42148] ^ n[42149];
assign t[42150] = t[42149] ^ n[42150];
assign t[42151] = t[42150] ^ n[42151];
assign t[42152] = t[42151] ^ n[42152];
assign t[42153] = t[42152] ^ n[42153];
assign t[42154] = t[42153] ^ n[42154];
assign t[42155] = t[42154] ^ n[42155];
assign t[42156] = t[42155] ^ n[42156];
assign t[42157] = t[42156] ^ n[42157];
assign t[42158] = t[42157] ^ n[42158];
assign t[42159] = t[42158] ^ n[42159];
assign t[42160] = t[42159] ^ n[42160];
assign t[42161] = t[42160] ^ n[42161];
assign t[42162] = t[42161] ^ n[42162];
assign t[42163] = t[42162] ^ n[42163];
assign t[42164] = t[42163] ^ n[42164];
assign t[42165] = t[42164] ^ n[42165];
assign t[42166] = t[42165] ^ n[42166];
assign t[42167] = t[42166] ^ n[42167];
assign t[42168] = t[42167] ^ n[42168];
assign t[42169] = t[42168] ^ n[42169];
assign t[42170] = t[42169] ^ n[42170];
assign t[42171] = t[42170] ^ n[42171];
assign t[42172] = t[42171] ^ n[42172];
assign t[42173] = t[42172] ^ n[42173];
assign t[42174] = t[42173] ^ n[42174];
assign t[42175] = t[42174] ^ n[42175];
assign t[42176] = t[42175] ^ n[42176];
assign t[42177] = t[42176] ^ n[42177];
assign t[42178] = t[42177] ^ n[42178];
assign t[42179] = t[42178] ^ n[42179];
assign t[42180] = t[42179] ^ n[42180];
assign t[42181] = t[42180] ^ n[42181];
assign t[42182] = t[42181] ^ n[42182];
assign t[42183] = t[42182] ^ n[42183];
assign t[42184] = t[42183] ^ n[42184];
assign t[42185] = t[42184] ^ n[42185];
assign t[42186] = t[42185] ^ n[42186];
assign t[42187] = t[42186] ^ n[42187];
assign t[42188] = t[42187] ^ n[42188];
assign t[42189] = t[42188] ^ n[42189];
assign t[42190] = t[42189] ^ n[42190];
assign t[42191] = t[42190] ^ n[42191];
assign t[42192] = t[42191] ^ n[42192];
assign t[42193] = t[42192] ^ n[42193];
assign t[42194] = t[42193] ^ n[42194];
assign t[42195] = t[42194] ^ n[42195];
assign t[42196] = t[42195] ^ n[42196];
assign t[42197] = t[42196] ^ n[42197];
assign t[42198] = t[42197] ^ n[42198];
assign t[42199] = t[42198] ^ n[42199];
assign t[42200] = t[42199] ^ n[42200];
assign t[42201] = t[42200] ^ n[42201];
assign t[42202] = t[42201] ^ n[42202];
assign t[42203] = t[42202] ^ n[42203];
assign t[42204] = t[42203] ^ n[42204];
assign t[42205] = t[42204] ^ n[42205];
assign t[42206] = t[42205] ^ n[42206];
assign t[42207] = t[42206] ^ n[42207];
assign t[42208] = t[42207] ^ n[42208];
assign t[42209] = t[42208] ^ n[42209];
assign t[42210] = t[42209] ^ n[42210];
assign t[42211] = t[42210] ^ n[42211];
assign t[42212] = t[42211] ^ n[42212];
assign t[42213] = t[42212] ^ n[42213];
assign t[42214] = t[42213] ^ n[42214];
assign t[42215] = t[42214] ^ n[42215];
assign t[42216] = t[42215] ^ n[42216];
assign t[42217] = t[42216] ^ n[42217];
assign t[42218] = t[42217] ^ n[42218];
assign t[42219] = t[42218] ^ n[42219];
assign t[42220] = t[42219] ^ n[42220];
assign t[42221] = t[42220] ^ n[42221];
assign t[42222] = t[42221] ^ n[42222];
assign t[42223] = t[42222] ^ n[42223];
assign t[42224] = t[42223] ^ n[42224];
assign t[42225] = t[42224] ^ n[42225];
assign t[42226] = t[42225] ^ n[42226];
assign t[42227] = t[42226] ^ n[42227];
assign t[42228] = t[42227] ^ n[42228];
assign t[42229] = t[42228] ^ n[42229];
assign t[42230] = t[42229] ^ n[42230];
assign t[42231] = t[42230] ^ n[42231];
assign t[42232] = t[42231] ^ n[42232];
assign t[42233] = t[42232] ^ n[42233];
assign t[42234] = t[42233] ^ n[42234];
assign t[42235] = t[42234] ^ n[42235];
assign t[42236] = t[42235] ^ n[42236];
assign t[42237] = t[42236] ^ n[42237];
assign t[42238] = t[42237] ^ n[42238];
assign t[42239] = t[42238] ^ n[42239];
assign t[42240] = t[42239] ^ n[42240];
assign t[42241] = t[42240] ^ n[42241];
assign t[42242] = t[42241] ^ n[42242];
assign t[42243] = t[42242] ^ n[42243];
assign t[42244] = t[42243] ^ n[42244];
assign t[42245] = t[42244] ^ n[42245];
assign t[42246] = t[42245] ^ n[42246];
assign t[42247] = t[42246] ^ n[42247];
assign t[42248] = t[42247] ^ n[42248];
assign t[42249] = t[42248] ^ n[42249];
assign t[42250] = t[42249] ^ n[42250];
assign t[42251] = t[42250] ^ n[42251];
assign t[42252] = t[42251] ^ n[42252];
assign t[42253] = t[42252] ^ n[42253];
assign t[42254] = t[42253] ^ n[42254];
assign t[42255] = t[42254] ^ n[42255];
assign t[42256] = t[42255] ^ n[42256];
assign t[42257] = t[42256] ^ n[42257];
assign t[42258] = t[42257] ^ n[42258];
assign t[42259] = t[42258] ^ n[42259];
assign t[42260] = t[42259] ^ n[42260];
assign t[42261] = t[42260] ^ n[42261];
assign t[42262] = t[42261] ^ n[42262];
assign t[42263] = t[42262] ^ n[42263];
assign t[42264] = t[42263] ^ n[42264];
assign t[42265] = t[42264] ^ n[42265];
assign t[42266] = t[42265] ^ n[42266];
assign t[42267] = t[42266] ^ n[42267];
assign t[42268] = t[42267] ^ n[42268];
assign t[42269] = t[42268] ^ n[42269];
assign t[42270] = t[42269] ^ n[42270];
assign t[42271] = t[42270] ^ n[42271];
assign t[42272] = t[42271] ^ n[42272];
assign t[42273] = t[42272] ^ n[42273];
assign t[42274] = t[42273] ^ n[42274];
assign t[42275] = t[42274] ^ n[42275];
assign t[42276] = t[42275] ^ n[42276];
assign t[42277] = t[42276] ^ n[42277];
assign t[42278] = t[42277] ^ n[42278];
assign t[42279] = t[42278] ^ n[42279];
assign t[42280] = t[42279] ^ n[42280];
assign t[42281] = t[42280] ^ n[42281];
assign t[42282] = t[42281] ^ n[42282];
assign t[42283] = t[42282] ^ n[42283];
assign t[42284] = t[42283] ^ n[42284];
assign t[42285] = t[42284] ^ n[42285];
assign t[42286] = t[42285] ^ n[42286];
assign t[42287] = t[42286] ^ n[42287];
assign t[42288] = t[42287] ^ n[42288];
assign t[42289] = t[42288] ^ n[42289];
assign t[42290] = t[42289] ^ n[42290];
assign t[42291] = t[42290] ^ n[42291];
assign t[42292] = t[42291] ^ n[42292];
assign t[42293] = t[42292] ^ n[42293];
assign t[42294] = t[42293] ^ n[42294];
assign t[42295] = t[42294] ^ n[42295];
assign t[42296] = t[42295] ^ n[42296];
assign t[42297] = t[42296] ^ n[42297];
assign t[42298] = t[42297] ^ n[42298];
assign t[42299] = t[42298] ^ n[42299];
assign t[42300] = t[42299] ^ n[42300];
assign t[42301] = t[42300] ^ n[42301];
assign t[42302] = t[42301] ^ n[42302];
assign t[42303] = t[42302] ^ n[42303];
assign t[42304] = t[42303] ^ n[42304];
assign t[42305] = t[42304] ^ n[42305];
assign t[42306] = t[42305] ^ n[42306];
assign t[42307] = t[42306] ^ n[42307];
assign t[42308] = t[42307] ^ n[42308];
assign t[42309] = t[42308] ^ n[42309];
assign t[42310] = t[42309] ^ n[42310];
assign t[42311] = t[42310] ^ n[42311];
assign t[42312] = t[42311] ^ n[42312];
assign t[42313] = t[42312] ^ n[42313];
assign t[42314] = t[42313] ^ n[42314];
assign t[42315] = t[42314] ^ n[42315];
assign t[42316] = t[42315] ^ n[42316];
assign t[42317] = t[42316] ^ n[42317];
assign t[42318] = t[42317] ^ n[42318];
assign t[42319] = t[42318] ^ n[42319];
assign t[42320] = t[42319] ^ n[42320];
assign t[42321] = t[42320] ^ n[42321];
assign t[42322] = t[42321] ^ n[42322];
assign t[42323] = t[42322] ^ n[42323];
assign t[42324] = t[42323] ^ n[42324];
assign t[42325] = t[42324] ^ n[42325];
assign t[42326] = t[42325] ^ n[42326];
assign t[42327] = t[42326] ^ n[42327];
assign t[42328] = t[42327] ^ n[42328];
assign t[42329] = t[42328] ^ n[42329];
assign t[42330] = t[42329] ^ n[42330];
assign t[42331] = t[42330] ^ n[42331];
assign t[42332] = t[42331] ^ n[42332];
assign t[42333] = t[42332] ^ n[42333];
assign t[42334] = t[42333] ^ n[42334];
assign t[42335] = t[42334] ^ n[42335];
assign t[42336] = t[42335] ^ n[42336];
assign t[42337] = t[42336] ^ n[42337];
assign t[42338] = t[42337] ^ n[42338];
assign t[42339] = t[42338] ^ n[42339];
assign t[42340] = t[42339] ^ n[42340];
assign t[42341] = t[42340] ^ n[42341];
assign t[42342] = t[42341] ^ n[42342];
assign t[42343] = t[42342] ^ n[42343];
assign t[42344] = t[42343] ^ n[42344];
assign t[42345] = t[42344] ^ n[42345];
assign t[42346] = t[42345] ^ n[42346];
assign t[42347] = t[42346] ^ n[42347];
assign t[42348] = t[42347] ^ n[42348];
assign t[42349] = t[42348] ^ n[42349];
assign t[42350] = t[42349] ^ n[42350];
assign t[42351] = t[42350] ^ n[42351];
assign t[42352] = t[42351] ^ n[42352];
assign t[42353] = t[42352] ^ n[42353];
assign t[42354] = t[42353] ^ n[42354];
assign t[42355] = t[42354] ^ n[42355];
assign t[42356] = t[42355] ^ n[42356];
assign t[42357] = t[42356] ^ n[42357];
assign t[42358] = t[42357] ^ n[42358];
assign t[42359] = t[42358] ^ n[42359];
assign t[42360] = t[42359] ^ n[42360];
assign t[42361] = t[42360] ^ n[42361];
assign t[42362] = t[42361] ^ n[42362];
assign t[42363] = t[42362] ^ n[42363];
assign t[42364] = t[42363] ^ n[42364];
assign t[42365] = t[42364] ^ n[42365];
assign t[42366] = t[42365] ^ n[42366];
assign t[42367] = t[42366] ^ n[42367];
assign t[42368] = t[42367] ^ n[42368];
assign t[42369] = t[42368] ^ n[42369];
assign t[42370] = t[42369] ^ n[42370];
assign t[42371] = t[42370] ^ n[42371];
assign t[42372] = t[42371] ^ n[42372];
assign t[42373] = t[42372] ^ n[42373];
assign t[42374] = t[42373] ^ n[42374];
assign t[42375] = t[42374] ^ n[42375];
assign t[42376] = t[42375] ^ n[42376];
assign t[42377] = t[42376] ^ n[42377];
assign t[42378] = t[42377] ^ n[42378];
assign t[42379] = t[42378] ^ n[42379];
assign t[42380] = t[42379] ^ n[42380];
assign t[42381] = t[42380] ^ n[42381];
assign t[42382] = t[42381] ^ n[42382];
assign t[42383] = t[42382] ^ n[42383];
assign t[42384] = t[42383] ^ n[42384];
assign t[42385] = t[42384] ^ n[42385];
assign t[42386] = t[42385] ^ n[42386];
assign t[42387] = t[42386] ^ n[42387];
assign t[42388] = t[42387] ^ n[42388];
assign t[42389] = t[42388] ^ n[42389];
assign t[42390] = t[42389] ^ n[42390];
assign t[42391] = t[42390] ^ n[42391];
assign t[42392] = t[42391] ^ n[42392];
assign t[42393] = t[42392] ^ n[42393];
assign t[42394] = t[42393] ^ n[42394];
assign t[42395] = t[42394] ^ n[42395];
assign t[42396] = t[42395] ^ n[42396];
assign t[42397] = t[42396] ^ n[42397];
assign t[42398] = t[42397] ^ n[42398];
assign t[42399] = t[42398] ^ n[42399];
assign t[42400] = t[42399] ^ n[42400];
assign t[42401] = t[42400] ^ n[42401];
assign t[42402] = t[42401] ^ n[42402];
assign t[42403] = t[42402] ^ n[42403];
assign t[42404] = t[42403] ^ n[42404];
assign t[42405] = t[42404] ^ n[42405];
assign t[42406] = t[42405] ^ n[42406];
assign t[42407] = t[42406] ^ n[42407];
assign t[42408] = t[42407] ^ n[42408];
assign t[42409] = t[42408] ^ n[42409];
assign t[42410] = t[42409] ^ n[42410];
assign t[42411] = t[42410] ^ n[42411];
assign t[42412] = t[42411] ^ n[42412];
assign t[42413] = t[42412] ^ n[42413];
assign t[42414] = t[42413] ^ n[42414];
assign t[42415] = t[42414] ^ n[42415];
assign t[42416] = t[42415] ^ n[42416];
assign t[42417] = t[42416] ^ n[42417];
assign t[42418] = t[42417] ^ n[42418];
assign t[42419] = t[42418] ^ n[42419];
assign t[42420] = t[42419] ^ n[42420];
assign t[42421] = t[42420] ^ n[42421];
assign t[42422] = t[42421] ^ n[42422];
assign t[42423] = t[42422] ^ n[42423];
assign t[42424] = t[42423] ^ n[42424];
assign t[42425] = t[42424] ^ n[42425];
assign t[42426] = t[42425] ^ n[42426];
assign t[42427] = t[42426] ^ n[42427];
assign t[42428] = t[42427] ^ n[42428];
assign t[42429] = t[42428] ^ n[42429];
assign t[42430] = t[42429] ^ n[42430];
assign t[42431] = t[42430] ^ n[42431];
assign t[42432] = t[42431] ^ n[42432];
assign t[42433] = t[42432] ^ n[42433];
assign t[42434] = t[42433] ^ n[42434];
assign t[42435] = t[42434] ^ n[42435];
assign t[42436] = t[42435] ^ n[42436];
assign t[42437] = t[42436] ^ n[42437];
assign t[42438] = t[42437] ^ n[42438];
assign t[42439] = t[42438] ^ n[42439];
assign t[42440] = t[42439] ^ n[42440];
assign t[42441] = t[42440] ^ n[42441];
assign t[42442] = t[42441] ^ n[42442];
assign t[42443] = t[42442] ^ n[42443];
assign t[42444] = t[42443] ^ n[42444];
assign t[42445] = t[42444] ^ n[42445];
assign t[42446] = t[42445] ^ n[42446];
assign t[42447] = t[42446] ^ n[42447];
assign t[42448] = t[42447] ^ n[42448];
assign t[42449] = t[42448] ^ n[42449];
assign t[42450] = t[42449] ^ n[42450];
assign t[42451] = t[42450] ^ n[42451];
assign t[42452] = t[42451] ^ n[42452];
assign t[42453] = t[42452] ^ n[42453];
assign t[42454] = t[42453] ^ n[42454];
assign t[42455] = t[42454] ^ n[42455];
assign t[42456] = t[42455] ^ n[42456];
assign t[42457] = t[42456] ^ n[42457];
assign t[42458] = t[42457] ^ n[42458];
assign t[42459] = t[42458] ^ n[42459];
assign t[42460] = t[42459] ^ n[42460];
assign t[42461] = t[42460] ^ n[42461];
assign t[42462] = t[42461] ^ n[42462];
assign t[42463] = t[42462] ^ n[42463];
assign t[42464] = t[42463] ^ n[42464];
assign t[42465] = t[42464] ^ n[42465];
assign t[42466] = t[42465] ^ n[42466];
assign t[42467] = t[42466] ^ n[42467];
assign t[42468] = t[42467] ^ n[42468];
assign t[42469] = t[42468] ^ n[42469];
assign t[42470] = t[42469] ^ n[42470];
assign t[42471] = t[42470] ^ n[42471];
assign t[42472] = t[42471] ^ n[42472];
assign t[42473] = t[42472] ^ n[42473];
assign t[42474] = t[42473] ^ n[42474];
assign t[42475] = t[42474] ^ n[42475];
assign t[42476] = t[42475] ^ n[42476];
assign t[42477] = t[42476] ^ n[42477];
assign t[42478] = t[42477] ^ n[42478];
assign t[42479] = t[42478] ^ n[42479];
assign t[42480] = t[42479] ^ n[42480];
assign t[42481] = t[42480] ^ n[42481];
assign t[42482] = t[42481] ^ n[42482];
assign t[42483] = t[42482] ^ n[42483];
assign t[42484] = t[42483] ^ n[42484];
assign t[42485] = t[42484] ^ n[42485];
assign t[42486] = t[42485] ^ n[42486];
assign t[42487] = t[42486] ^ n[42487];
assign t[42488] = t[42487] ^ n[42488];
assign t[42489] = t[42488] ^ n[42489];
assign t[42490] = t[42489] ^ n[42490];
assign t[42491] = t[42490] ^ n[42491];
assign t[42492] = t[42491] ^ n[42492];
assign t[42493] = t[42492] ^ n[42493];
assign t[42494] = t[42493] ^ n[42494];
assign t[42495] = t[42494] ^ n[42495];
assign t[42496] = t[42495] ^ n[42496];
assign t[42497] = t[42496] ^ n[42497];
assign t[42498] = t[42497] ^ n[42498];
assign t[42499] = t[42498] ^ n[42499];
assign t[42500] = t[42499] ^ n[42500];
assign t[42501] = t[42500] ^ n[42501];
assign t[42502] = t[42501] ^ n[42502];
assign t[42503] = t[42502] ^ n[42503];
assign t[42504] = t[42503] ^ n[42504];
assign t[42505] = t[42504] ^ n[42505];
assign t[42506] = t[42505] ^ n[42506];
assign t[42507] = t[42506] ^ n[42507];
assign t[42508] = t[42507] ^ n[42508];
assign t[42509] = t[42508] ^ n[42509];
assign t[42510] = t[42509] ^ n[42510];
assign t[42511] = t[42510] ^ n[42511];
assign t[42512] = t[42511] ^ n[42512];
assign t[42513] = t[42512] ^ n[42513];
assign t[42514] = t[42513] ^ n[42514];
assign t[42515] = t[42514] ^ n[42515];
assign t[42516] = t[42515] ^ n[42516];
assign t[42517] = t[42516] ^ n[42517];
assign t[42518] = t[42517] ^ n[42518];
assign t[42519] = t[42518] ^ n[42519];
assign t[42520] = t[42519] ^ n[42520];
assign t[42521] = t[42520] ^ n[42521];
assign t[42522] = t[42521] ^ n[42522];
assign t[42523] = t[42522] ^ n[42523];
assign t[42524] = t[42523] ^ n[42524];
assign t[42525] = t[42524] ^ n[42525];
assign t[42526] = t[42525] ^ n[42526];
assign t[42527] = t[42526] ^ n[42527];
assign t[42528] = t[42527] ^ n[42528];
assign t[42529] = t[42528] ^ n[42529];
assign t[42530] = t[42529] ^ n[42530];
assign t[42531] = t[42530] ^ n[42531];
assign t[42532] = t[42531] ^ n[42532];
assign t[42533] = t[42532] ^ n[42533];
assign t[42534] = t[42533] ^ n[42534];
assign t[42535] = t[42534] ^ n[42535];
assign t[42536] = t[42535] ^ n[42536];
assign t[42537] = t[42536] ^ n[42537];
assign t[42538] = t[42537] ^ n[42538];
assign t[42539] = t[42538] ^ n[42539];
assign t[42540] = t[42539] ^ n[42540];
assign t[42541] = t[42540] ^ n[42541];
assign t[42542] = t[42541] ^ n[42542];
assign t[42543] = t[42542] ^ n[42543];
assign t[42544] = t[42543] ^ n[42544];
assign t[42545] = t[42544] ^ n[42545];
assign t[42546] = t[42545] ^ n[42546];
assign t[42547] = t[42546] ^ n[42547];
assign t[42548] = t[42547] ^ n[42548];
assign t[42549] = t[42548] ^ n[42549];
assign t[42550] = t[42549] ^ n[42550];
assign t[42551] = t[42550] ^ n[42551];
assign t[42552] = t[42551] ^ n[42552];
assign t[42553] = t[42552] ^ n[42553];
assign t[42554] = t[42553] ^ n[42554];
assign t[42555] = t[42554] ^ n[42555];
assign t[42556] = t[42555] ^ n[42556];
assign t[42557] = t[42556] ^ n[42557];
assign t[42558] = t[42557] ^ n[42558];
assign t[42559] = t[42558] ^ n[42559];
assign t[42560] = t[42559] ^ n[42560];
assign t[42561] = t[42560] ^ n[42561];
assign t[42562] = t[42561] ^ n[42562];
assign t[42563] = t[42562] ^ n[42563];
assign t[42564] = t[42563] ^ n[42564];
assign t[42565] = t[42564] ^ n[42565];
assign t[42566] = t[42565] ^ n[42566];
assign t[42567] = t[42566] ^ n[42567];
assign t[42568] = t[42567] ^ n[42568];
assign t[42569] = t[42568] ^ n[42569];
assign t[42570] = t[42569] ^ n[42570];
assign t[42571] = t[42570] ^ n[42571];
assign t[42572] = t[42571] ^ n[42572];
assign t[42573] = t[42572] ^ n[42573];
assign t[42574] = t[42573] ^ n[42574];
assign t[42575] = t[42574] ^ n[42575];
assign t[42576] = t[42575] ^ n[42576];
assign t[42577] = t[42576] ^ n[42577];
assign t[42578] = t[42577] ^ n[42578];
assign t[42579] = t[42578] ^ n[42579];
assign t[42580] = t[42579] ^ n[42580];
assign t[42581] = t[42580] ^ n[42581];
assign t[42582] = t[42581] ^ n[42582];
assign t[42583] = t[42582] ^ n[42583];
assign t[42584] = t[42583] ^ n[42584];
assign t[42585] = t[42584] ^ n[42585];
assign t[42586] = t[42585] ^ n[42586];
assign t[42587] = t[42586] ^ n[42587];
assign t[42588] = t[42587] ^ n[42588];
assign t[42589] = t[42588] ^ n[42589];
assign t[42590] = t[42589] ^ n[42590];
assign t[42591] = t[42590] ^ n[42591];
assign t[42592] = t[42591] ^ n[42592];
assign t[42593] = t[42592] ^ n[42593];
assign t[42594] = t[42593] ^ n[42594];
assign t[42595] = t[42594] ^ n[42595];
assign t[42596] = t[42595] ^ n[42596];
assign t[42597] = t[42596] ^ n[42597];
assign t[42598] = t[42597] ^ n[42598];
assign t[42599] = t[42598] ^ n[42599];
assign t[42600] = t[42599] ^ n[42600];
assign t[42601] = t[42600] ^ n[42601];
assign t[42602] = t[42601] ^ n[42602];
assign t[42603] = t[42602] ^ n[42603];
assign t[42604] = t[42603] ^ n[42604];
assign t[42605] = t[42604] ^ n[42605];
assign t[42606] = t[42605] ^ n[42606];
assign t[42607] = t[42606] ^ n[42607];
assign t[42608] = t[42607] ^ n[42608];
assign t[42609] = t[42608] ^ n[42609];
assign t[42610] = t[42609] ^ n[42610];
assign t[42611] = t[42610] ^ n[42611];
assign t[42612] = t[42611] ^ n[42612];
assign t[42613] = t[42612] ^ n[42613];
assign t[42614] = t[42613] ^ n[42614];
assign t[42615] = t[42614] ^ n[42615];
assign t[42616] = t[42615] ^ n[42616];
assign t[42617] = t[42616] ^ n[42617];
assign t[42618] = t[42617] ^ n[42618];
assign t[42619] = t[42618] ^ n[42619];
assign t[42620] = t[42619] ^ n[42620];
assign t[42621] = t[42620] ^ n[42621];
assign t[42622] = t[42621] ^ n[42622];
assign t[42623] = t[42622] ^ n[42623];
assign t[42624] = t[42623] ^ n[42624];
assign t[42625] = t[42624] ^ n[42625];
assign t[42626] = t[42625] ^ n[42626];
assign t[42627] = t[42626] ^ n[42627];
assign t[42628] = t[42627] ^ n[42628];
assign t[42629] = t[42628] ^ n[42629];
assign t[42630] = t[42629] ^ n[42630];
assign t[42631] = t[42630] ^ n[42631];
assign t[42632] = t[42631] ^ n[42632];
assign t[42633] = t[42632] ^ n[42633];
assign t[42634] = t[42633] ^ n[42634];
assign t[42635] = t[42634] ^ n[42635];
assign t[42636] = t[42635] ^ n[42636];
assign t[42637] = t[42636] ^ n[42637];
assign t[42638] = t[42637] ^ n[42638];
assign t[42639] = t[42638] ^ n[42639];
assign t[42640] = t[42639] ^ n[42640];
assign t[42641] = t[42640] ^ n[42641];
assign t[42642] = t[42641] ^ n[42642];
assign t[42643] = t[42642] ^ n[42643];
assign t[42644] = t[42643] ^ n[42644];
assign t[42645] = t[42644] ^ n[42645];
assign t[42646] = t[42645] ^ n[42646];
assign t[42647] = t[42646] ^ n[42647];
assign t[42648] = t[42647] ^ n[42648];
assign t[42649] = t[42648] ^ n[42649];
assign t[42650] = t[42649] ^ n[42650];
assign t[42651] = t[42650] ^ n[42651];
assign t[42652] = t[42651] ^ n[42652];
assign t[42653] = t[42652] ^ n[42653];
assign t[42654] = t[42653] ^ n[42654];
assign t[42655] = t[42654] ^ n[42655];
assign t[42656] = t[42655] ^ n[42656];
assign t[42657] = t[42656] ^ n[42657];
assign t[42658] = t[42657] ^ n[42658];
assign t[42659] = t[42658] ^ n[42659];
assign t[42660] = t[42659] ^ n[42660];
assign t[42661] = t[42660] ^ n[42661];
assign t[42662] = t[42661] ^ n[42662];
assign t[42663] = t[42662] ^ n[42663];
assign t[42664] = t[42663] ^ n[42664];
assign t[42665] = t[42664] ^ n[42665];
assign t[42666] = t[42665] ^ n[42666];
assign t[42667] = t[42666] ^ n[42667];
assign t[42668] = t[42667] ^ n[42668];
assign t[42669] = t[42668] ^ n[42669];
assign t[42670] = t[42669] ^ n[42670];
assign t[42671] = t[42670] ^ n[42671];
assign t[42672] = t[42671] ^ n[42672];
assign t[42673] = t[42672] ^ n[42673];
assign t[42674] = t[42673] ^ n[42674];
assign t[42675] = t[42674] ^ n[42675];
assign t[42676] = t[42675] ^ n[42676];
assign t[42677] = t[42676] ^ n[42677];
assign t[42678] = t[42677] ^ n[42678];
assign t[42679] = t[42678] ^ n[42679];
assign t[42680] = t[42679] ^ n[42680];
assign t[42681] = t[42680] ^ n[42681];
assign t[42682] = t[42681] ^ n[42682];
assign t[42683] = t[42682] ^ n[42683];
assign t[42684] = t[42683] ^ n[42684];
assign t[42685] = t[42684] ^ n[42685];
assign t[42686] = t[42685] ^ n[42686];
assign t[42687] = t[42686] ^ n[42687];
assign t[42688] = t[42687] ^ n[42688];
assign t[42689] = t[42688] ^ n[42689];
assign t[42690] = t[42689] ^ n[42690];
assign t[42691] = t[42690] ^ n[42691];
assign t[42692] = t[42691] ^ n[42692];
assign t[42693] = t[42692] ^ n[42693];
assign t[42694] = t[42693] ^ n[42694];
assign t[42695] = t[42694] ^ n[42695];
assign t[42696] = t[42695] ^ n[42696];
assign t[42697] = t[42696] ^ n[42697];
assign t[42698] = t[42697] ^ n[42698];
assign t[42699] = t[42698] ^ n[42699];
assign t[42700] = t[42699] ^ n[42700];
assign t[42701] = t[42700] ^ n[42701];
assign t[42702] = t[42701] ^ n[42702];
assign t[42703] = t[42702] ^ n[42703];
assign t[42704] = t[42703] ^ n[42704];
assign t[42705] = t[42704] ^ n[42705];
assign t[42706] = t[42705] ^ n[42706];
assign t[42707] = t[42706] ^ n[42707];
assign t[42708] = t[42707] ^ n[42708];
assign t[42709] = t[42708] ^ n[42709];
assign t[42710] = t[42709] ^ n[42710];
assign t[42711] = t[42710] ^ n[42711];
assign t[42712] = t[42711] ^ n[42712];
assign t[42713] = t[42712] ^ n[42713];
assign t[42714] = t[42713] ^ n[42714];
assign t[42715] = t[42714] ^ n[42715];
assign t[42716] = t[42715] ^ n[42716];
assign t[42717] = t[42716] ^ n[42717];
assign t[42718] = t[42717] ^ n[42718];
assign t[42719] = t[42718] ^ n[42719];
assign t[42720] = t[42719] ^ n[42720];
assign t[42721] = t[42720] ^ n[42721];
assign t[42722] = t[42721] ^ n[42722];
assign t[42723] = t[42722] ^ n[42723];
assign t[42724] = t[42723] ^ n[42724];
assign t[42725] = t[42724] ^ n[42725];
assign t[42726] = t[42725] ^ n[42726];
assign t[42727] = t[42726] ^ n[42727];
assign t[42728] = t[42727] ^ n[42728];
assign t[42729] = t[42728] ^ n[42729];
assign t[42730] = t[42729] ^ n[42730];
assign t[42731] = t[42730] ^ n[42731];
assign t[42732] = t[42731] ^ n[42732];
assign t[42733] = t[42732] ^ n[42733];
assign t[42734] = t[42733] ^ n[42734];
assign t[42735] = t[42734] ^ n[42735];
assign t[42736] = t[42735] ^ n[42736];
assign t[42737] = t[42736] ^ n[42737];
assign t[42738] = t[42737] ^ n[42738];
assign t[42739] = t[42738] ^ n[42739];
assign t[42740] = t[42739] ^ n[42740];
assign t[42741] = t[42740] ^ n[42741];
assign t[42742] = t[42741] ^ n[42742];
assign t[42743] = t[42742] ^ n[42743];
assign t[42744] = t[42743] ^ n[42744];
assign t[42745] = t[42744] ^ n[42745];
assign t[42746] = t[42745] ^ n[42746];
assign t[42747] = t[42746] ^ n[42747];
assign t[42748] = t[42747] ^ n[42748];
assign t[42749] = t[42748] ^ n[42749];
assign t[42750] = t[42749] ^ n[42750];
assign t[42751] = t[42750] ^ n[42751];
assign t[42752] = t[42751] ^ n[42752];
assign t[42753] = t[42752] ^ n[42753];
assign t[42754] = t[42753] ^ n[42754];
assign t[42755] = t[42754] ^ n[42755];
assign t[42756] = t[42755] ^ n[42756];
assign t[42757] = t[42756] ^ n[42757];
assign t[42758] = t[42757] ^ n[42758];
assign t[42759] = t[42758] ^ n[42759];
assign t[42760] = t[42759] ^ n[42760];
assign t[42761] = t[42760] ^ n[42761];
assign t[42762] = t[42761] ^ n[42762];
assign t[42763] = t[42762] ^ n[42763];
assign t[42764] = t[42763] ^ n[42764];
assign t[42765] = t[42764] ^ n[42765];
assign t[42766] = t[42765] ^ n[42766];
assign t[42767] = t[42766] ^ n[42767];
assign t[42768] = t[42767] ^ n[42768];
assign t[42769] = t[42768] ^ n[42769];
assign t[42770] = t[42769] ^ n[42770];
assign t[42771] = t[42770] ^ n[42771];
assign t[42772] = t[42771] ^ n[42772];
assign t[42773] = t[42772] ^ n[42773];
assign t[42774] = t[42773] ^ n[42774];
assign t[42775] = t[42774] ^ n[42775];
assign t[42776] = t[42775] ^ n[42776];
assign t[42777] = t[42776] ^ n[42777];
assign t[42778] = t[42777] ^ n[42778];
assign t[42779] = t[42778] ^ n[42779];
assign t[42780] = t[42779] ^ n[42780];
assign t[42781] = t[42780] ^ n[42781];
assign t[42782] = t[42781] ^ n[42782];
assign t[42783] = t[42782] ^ n[42783];
assign t[42784] = t[42783] ^ n[42784];
assign t[42785] = t[42784] ^ n[42785];
assign t[42786] = t[42785] ^ n[42786];
assign t[42787] = t[42786] ^ n[42787];
assign t[42788] = t[42787] ^ n[42788];
assign t[42789] = t[42788] ^ n[42789];
assign t[42790] = t[42789] ^ n[42790];
assign t[42791] = t[42790] ^ n[42791];
assign t[42792] = t[42791] ^ n[42792];
assign t[42793] = t[42792] ^ n[42793];
assign t[42794] = t[42793] ^ n[42794];
assign t[42795] = t[42794] ^ n[42795];
assign t[42796] = t[42795] ^ n[42796];
assign t[42797] = t[42796] ^ n[42797];
assign t[42798] = t[42797] ^ n[42798];
assign t[42799] = t[42798] ^ n[42799];
assign t[42800] = t[42799] ^ n[42800];
assign t[42801] = t[42800] ^ n[42801];
assign t[42802] = t[42801] ^ n[42802];
assign t[42803] = t[42802] ^ n[42803];
assign t[42804] = t[42803] ^ n[42804];
assign t[42805] = t[42804] ^ n[42805];
assign t[42806] = t[42805] ^ n[42806];
assign t[42807] = t[42806] ^ n[42807];
assign t[42808] = t[42807] ^ n[42808];
assign t[42809] = t[42808] ^ n[42809];
assign t[42810] = t[42809] ^ n[42810];
assign t[42811] = t[42810] ^ n[42811];
assign t[42812] = t[42811] ^ n[42812];
assign t[42813] = t[42812] ^ n[42813];
assign t[42814] = t[42813] ^ n[42814];
assign t[42815] = t[42814] ^ n[42815];
assign t[42816] = t[42815] ^ n[42816];
assign t[42817] = t[42816] ^ n[42817];
assign t[42818] = t[42817] ^ n[42818];
assign t[42819] = t[42818] ^ n[42819];
assign t[42820] = t[42819] ^ n[42820];
assign t[42821] = t[42820] ^ n[42821];
assign t[42822] = t[42821] ^ n[42822];
assign t[42823] = t[42822] ^ n[42823];
assign t[42824] = t[42823] ^ n[42824];
assign t[42825] = t[42824] ^ n[42825];
assign t[42826] = t[42825] ^ n[42826];
assign t[42827] = t[42826] ^ n[42827];
assign t[42828] = t[42827] ^ n[42828];
assign t[42829] = t[42828] ^ n[42829];
assign t[42830] = t[42829] ^ n[42830];
assign t[42831] = t[42830] ^ n[42831];
assign t[42832] = t[42831] ^ n[42832];
assign t[42833] = t[42832] ^ n[42833];
assign t[42834] = t[42833] ^ n[42834];
assign t[42835] = t[42834] ^ n[42835];
assign t[42836] = t[42835] ^ n[42836];
assign t[42837] = t[42836] ^ n[42837];
assign t[42838] = t[42837] ^ n[42838];
assign t[42839] = t[42838] ^ n[42839];
assign t[42840] = t[42839] ^ n[42840];
assign t[42841] = t[42840] ^ n[42841];
assign t[42842] = t[42841] ^ n[42842];
assign t[42843] = t[42842] ^ n[42843];
assign t[42844] = t[42843] ^ n[42844];
assign t[42845] = t[42844] ^ n[42845];
assign t[42846] = t[42845] ^ n[42846];
assign t[42847] = t[42846] ^ n[42847];
assign t[42848] = t[42847] ^ n[42848];
assign t[42849] = t[42848] ^ n[42849];
assign t[42850] = t[42849] ^ n[42850];
assign t[42851] = t[42850] ^ n[42851];
assign t[42852] = t[42851] ^ n[42852];
assign t[42853] = t[42852] ^ n[42853];
assign t[42854] = t[42853] ^ n[42854];
assign t[42855] = t[42854] ^ n[42855];
assign t[42856] = t[42855] ^ n[42856];
assign t[42857] = t[42856] ^ n[42857];
assign t[42858] = t[42857] ^ n[42858];
assign t[42859] = t[42858] ^ n[42859];
assign t[42860] = t[42859] ^ n[42860];
assign t[42861] = t[42860] ^ n[42861];
assign t[42862] = t[42861] ^ n[42862];
assign t[42863] = t[42862] ^ n[42863];
assign t[42864] = t[42863] ^ n[42864];
assign t[42865] = t[42864] ^ n[42865];
assign t[42866] = t[42865] ^ n[42866];
assign t[42867] = t[42866] ^ n[42867];
assign t[42868] = t[42867] ^ n[42868];
assign t[42869] = t[42868] ^ n[42869];
assign t[42870] = t[42869] ^ n[42870];
assign t[42871] = t[42870] ^ n[42871];
assign t[42872] = t[42871] ^ n[42872];
assign t[42873] = t[42872] ^ n[42873];
assign t[42874] = t[42873] ^ n[42874];
assign t[42875] = t[42874] ^ n[42875];
assign t[42876] = t[42875] ^ n[42876];
assign t[42877] = t[42876] ^ n[42877];
assign t[42878] = t[42877] ^ n[42878];
assign t[42879] = t[42878] ^ n[42879];
assign t[42880] = t[42879] ^ n[42880];
assign t[42881] = t[42880] ^ n[42881];
assign t[42882] = t[42881] ^ n[42882];
assign t[42883] = t[42882] ^ n[42883];
assign t[42884] = t[42883] ^ n[42884];
assign t[42885] = t[42884] ^ n[42885];
assign t[42886] = t[42885] ^ n[42886];
assign t[42887] = t[42886] ^ n[42887];
assign t[42888] = t[42887] ^ n[42888];
assign t[42889] = t[42888] ^ n[42889];
assign t[42890] = t[42889] ^ n[42890];
assign t[42891] = t[42890] ^ n[42891];
assign t[42892] = t[42891] ^ n[42892];
assign t[42893] = t[42892] ^ n[42893];
assign t[42894] = t[42893] ^ n[42894];
assign t[42895] = t[42894] ^ n[42895];
assign t[42896] = t[42895] ^ n[42896];
assign t[42897] = t[42896] ^ n[42897];
assign t[42898] = t[42897] ^ n[42898];
assign t[42899] = t[42898] ^ n[42899];
assign t[42900] = t[42899] ^ n[42900];
assign t[42901] = t[42900] ^ n[42901];
assign t[42902] = t[42901] ^ n[42902];
assign t[42903] = t[42902] ^ n[42903];
assign t[42904] = t[42903] ^ n[42904];
assign t[42905] = t[42904] ^ n[42905];
assign t[42906] = t[42905] ^ n[42906];
assign t[42907] = t[42906] ^ n[42907];
assign t[42908] = t[42907] ^ n[42908];
assign t[42909] = t[42908] ^ n[42909];
assign t[42910] = t[42909] ^ n[42910];
assign t[42911] = t[42910] ^ n[42911];
assign t[42912] = t[42911] ^ n[42912];
assign t[42913] = t[42912] ^ n[42913];
assign t[42914] = t[42913] ^ n[42914];
assign t[42915] = t[42914] ^ n[42915];
assign t[42916] = t[42915] ^ n[42916];
assign t[42917] = t[42916] ^ n[42917];
assign t[42918] = t[42917] ^ n[42918];
assign t[42919] = t[42918] ^ n[42919];
assign t[42920] = t[42919] ^ n[42920];
assign t[42921] = t[42920] ^ n[42921];
assign t[42922] = t[42921] ^ n[42922];
assign t[42923] = t[42922] ^ n[42923];
assign t[42924] = t[42923] ^ n[42924];
assign t[42925] = t[42924] ^ n[42925];
assign t[42926] = t[42925] ^ n[42926];
assign t[42927] = t[42926] ^ n[42927];
assign t[42928] = t[42927] ^ n[42928];
assign t[42929] = t[42928] ^ n[42929];
assign t[42930] = t[42929] ^ n[42930];
assign t[42931] = t[42930] ^ n[42931];
assign t[42932] = t[42931] ^ n[42932];
assign t[42933] = t[42932] ^ n[42933];
assign t[42934] = t[42933] ^ n[42934];
assign t[42935] = t[42934] ^ n[42935];
assign t[42936] = t[42935] ^ n[42936];
assign t[42937] = t[42936] ^ n[42937];
assign t[42938] = t[42937] ^ n[42938];
assign t[42939] = t[42938] ^ n[42939];
assign t[42940] = t[42939] ^ n[42940];
assign t[42941] = t[42940] ^ n[42941];
assign t[42942] = t[42941] ^ n[42942];
assign t[42943] = t[42942] ^ n[42943];
assign t[42944] = t[42943] ^ n[42944];
assign t[42945] = t[42944] ^ n[42945];
assign t[42946] = t[42945] ^ n[42946];
assign t[42947] = t[42946] ^ n[42947];
assign t[42948] = t[42947] ^ n[42948];
assign t[42949] = t[42948] ^ n[42949];
assign t[42950] = t[42949] ^ n[42950];
assign t[42951] = t[42950] ^ n[42951];
assign t[42952] = t[42951] ^ n[42952];
assign t[42953] = t[42952] ^ n[42953];
assign t[42954] = t[42953] ^ n[42954];
assign t[42955] = t[42954] ^ n[42955];
assign t[42956] = t[42955] ^ n[42956];
assign t[42957] = t[42956] ^ n[42957];
assign t[42958] = t[42957] ^ n[42958];
assign t[42959] = t[42958] ^ n[42959];
assign t[42960] = t[42959] ^ n[42960];
assign t[42961] = t[42960] ^ n[42961];
assign t[42962] = t[42961] ^ n[42962];
assign t[42963] = t[42962] ^ n[42963];
assign t[42964] = t[42963] ^ n[42964];
assign t[42965] = t[42964] ^ n[42965];
assign t[42966] = t[42965] ^ n[42966];
assign t[42967] = t[42966] ^ n[42967];
assign t[42968] = t[42967] ^ n[42968];
assign t[42969] = t[42968] ^ n[42969];
assign t[42970] = t[42969] ^ n[42970];
assign t[42971] = t[42970] ^ n[42971];
assign t[42972] = t[42971] ^ n[42972];
assign t[42973] = t[42972] ^ n[42973];
assign t[42974] = t[42973] ^ n[42974];
assign t[42975] = t[42974] ^ n[42975];
assign t[42976] = t[42975] ^ n[42976];
assign t[42977] = t[42976] ^ n[42977];
assign t[42978] = t[42977] ^ n[42978];
assign t[42979] = t[42978] ^ n[42979];
assign t[42980] = t[42979] ^ n[42980];
assign t[42981] = t[42980] ^ n[42981];
assign t[42982] = t[42981] ^ n[42982];
assign t[42983] = t[42982] ^ n[42983];
assign t[42984] = t[42983] ^ n[42984];
assign t[42985] = t[42984] ^ n[42985];
assign t[42986] = t[42985] ^ n[42986];
assign t[42987] = t[42986] ^ n[42987];
assign t[42988] = t[42987] ^ n[42988];
assign t[42989] = t[42988] ^ n[42989];
assign t[42990] = t[42989] ^ n[42990];
assign t[42991] = t[42990] ^ n[42991];
assign t[42992] = t[42991] ^ n[42992];
assign t[42993] = t[42992] ^ n[42993];
assign t[42994] = t[42993] ^ n[42994];
assign t[42995] = t[42994] ^ n[42995];
assign t[42996] = t[42995] ^ n[42996];
assign t[42997] = t[42996] ^ n[42997];
assign t[42998] = t[42997] ^ n[42998];
assign t[42999] = t[42998] ^ n[42999];
assign t[43000] = t[42999] ^ n[43000];
assign t[43001] = t[43000] ^ n[43001];
assign t[43002] = t[43001] ^ n[43002];
assign t[43003] = t[43002] ^ n[43003];
assign t[43004] = t[43003] ^ n[43004];
assign t[43005] = t[43004] ^ n[43005];
assign t[43006] = t[43005] ^ n[43006];
assign t[43007] = t[43006] ^ n[43007];
assign t[43008] = t[43007] ^ n[43008];
assign t[43009] = t[43008] ^ n[43009];
assign t[43010] = t[43009] ^ n[43010];
assign t[43011] = t[43010] ^ n[43011];
assign t[43012] = t[43011] ^ n[43012];
assign t[43013] = t[43012] ^ n[43013];
assign t[43014] = t[43013] ^ n[43014];
assign t[43015] = t[43014] ^ n[43015];
assign t[43016] = t[43015] ^ n[43016];
assign t[43017] = t[43016] ^ n[43017];
assign t[43018] = t[43017] ^ n[43018];
assign t[43019] = t[43018] ^ n[43019];
assign t[43020] = t[43019] ^ n[43020];
assign t[43021] = t[43020] ^ n[43021];
assign t[43022] = t[43021] ^ n[43022];
assign t[43023] = t[43022] ^ n[43023];
assign t[43024] = t[43023] ^ n[43024];
assign t[43025] = t[43024] ^ n[43025];
assign t[43026] = t[43025] ^ n[43026];
assign t[43027] = t[43026] ^ n[43027];
assign t[43028] = t[43027] ^ n[43028];
assign t[43029] = t[43028] ^ n[43029];
assign t[43030] = t[43029] ^ n[43030];
assign t[43031] = t[43030] ^ n[43031];
assign t[43032] = t[43031] ^ n[43032];
assign t[43033] = t[43032] ^ n[43033];
assign t[43034] = t[43033] ^ n[43034];
assign t[43035] = t[43034] ^ n[43035];
assign t[43036] = t[43035] ^ n[43036];
assign t[43037] = t[43036] ^ n[43037];
assign t[43038] = t[43037] ^ n[43038];
assign t[43039] = t[43038] ^ n[43039];
assign t[43040] = t[43039] ^ n[43040];
assign t[43041] = t[43040] ^ n[43041];
assign t[43042] = t[43041] ^ n[43042];
assign t[43043] = t[43042] ^ n[43043];
assign t[43044] = t[43043] ^ n[43044];
assign t[43045] = t[43044] ^ n[43045];
assign t[43046] = t[43045] ^ n[43046];
assign t[43047] = t[43046] ^ n[43047];
assign t[43048] = t[43047] ^ n[43048];
assign t[43049] = t[43048] ^ n[43049];
assign t[43050] = t[43049] ^ n[43050];
assign t[43051] = t[43050] ^ n[43051];
assign t[43052] = t[43051] ^ n[43052];
assign t[43053] = t[43052] ^ n[43053];
assign t[43054] = t[43053] ^ n[43054];
assign t[43055] = t[43054] ^ n[43055];
assign t[43056] = t[43055] ^ n[43056];
assign t[43057] = t[43056] ^ n[43057];
assign t[43058] = t[43057] ^ n[43058];
assign t[43059] = t[43058] ^ n[43059];
assign t[43060] = t[43059] ^ n[43060];
assign t[43061] = t[43060] ^ n[43061];
assign t[43062] = t[43061] ^ n[43062];
assign t[43063] = t[43062] ^ n[43063];
assign t[43064] = t[43063] ^ n[43064];
assign t[43065] = t[43064] ^ n[43065];
assign t[43066] = t[43065] ^ n[43066];
assign t[43067] = t[43066] ^ n[43067];
assign t[43068] = t[43067] ^ n[43068];
assign t[43069] = t[43068] ^ n[43069];
assign t[43070] = t[43069] ^ n[43070];
assign t[43071] = t[43070] ^ n[43071];
assign t[43072] = t[43071] ^ n[43072];
assign t[43073] = t[43072] ^ n[43073];
assign t[43074] = t[43073] ^ n[43074];
assign t[43075] = t[43074] ^ n[43075];
assign t[43076] = t[43075] ^ n[43076];
assign t[43077] = t[43076] ^ n[43077];
assign t[43078] = t[43077] ^ n[43078];
assign t[43079] = t[43078] ^ n[43079];
assign t[43080] = t[43079] ^ n[43080];
assign t[43081] = t[43080] ^ n[43081];
assign t[43082] = t[43081] ^ n[43082];
assign t[43083] = t[43082] ^ n[43083];
assign t[43084] = t[43083] ^ n[43084];
assign t[43085] = t[43084] ^ n[43085];
assign t[43086] = t[43085] ^ n[43086];
assign t[43087] = t[43086] ^ n[43087];
assign t[43088] = t[43087] ^ n[43088];
assign t[43089] = t[43088] ^ n[43089];
assign t[43090] = t[43089] ^ n[43090];
assign t[43091] = t[43090] ^ n[43091];
assign t[43092] = t[43091] ^ n[43092];
assign t[43093] = t[43092] ^ n[43093];
assign t[43094] = t[43093] ^ n[43094];
assign t[43095] = t[43094] ^ n[43095];
assign t[43096] = t[43095] ^ n[43096];
assign t[43097] = t[43096] ^ n[43097];
assign t[43098] = t[43097] ^ n[43098];
assign t[43099] = t[43098] ^ n[43099];
assign t[43100] = t[43099] ^ n[43100];
assign t[43101] = t[43100] ^ n[43101];
assign t[43102] = t[43101] ^ n[43102];
assign t[43103] = t[43102] ^ n[43103];
assign t[43104] = t[43103] ^ n[43104];
assign t[43105] = t[43104] ^ n[43105];
assign t[43106] = t[43105] ^ n[43106];
assign t[43107] = t[43106] ^ n[43107];
assign t[43108] = t[43107] ^ n[43108];
assign t[43109] = t[43108] ^ n[43109];
assign t[43110] = t[43109] ^ n[43110];
assign t[43111] = t[43110] ^ n[43111];
assign t[43112] = t[43111] ^ n[43112];
assign t[43113] = t[43112] ^ n[43113];
assign t[43114] = t[43113] ^ n[43114];
assign t[43115] = t[43114] ^ n[43115];
assign t[43116] = t[43115] ^ n[43116];
assign t[43117] = t[43116] ^ n[43117];
assign t[43118] = t[43117] ^ n[43118];
assign t[43119] = t[43118] ^ n[43119];
assign t[43120] = t[43119] ^ n[43120];
assign t[43121] = t[43120] ^ n[43121];
assign t[43122] = t[43121] ^ n[43122];
assign t[43123] = t[43122] ^ n[43123];
assign t[43124] = t[43123] ^ n[43124];
assign t[43125] = t[43124] ^ n[43125];
assign t[43126] = t[43125] ^ n[43126];
assign t[43127] = t[43126] ^ n[43127];
assign t[43128] = t[43127] ^ n[43128];
assign t[43129] = t[43128] ^ n[43129];
assign t[43130] = t[43129] ^ n[43130];
assign t[43131] = t[43130] ^ n[43131];
assign t[43132] = t[43131] ^ n[43132];
assign t[43133] = t[43132] ^ n[43133];
assign t[43134] = t[43133] ^ n[43134];
assign t[43135] = t[43134] ^ n[43135];
assign t[43136] = t[43135] ^ n[43136];
assign t[43137] = t[43136] ^ n[43137];
assign t[43138] = t[43137] ^ n[43138];
assign t[43139] = t[43138] ^ n[43139];
assign t[43140] = t[43139] ^ n[43140];
assign t[43141] = t[43140] ^ n[43141];
assign t[43142] = t[43141] ^ n[43142];
assign t[43143] = t[43142] ^ n[43143];
assign t[43144] = t[43143] ^ n[43144];
assign t[43145] = t[43144] ^ n[43145];
assign t[43146] = t[43145] ^ n[43146];
assign t[43147] = t[43146] ^ n[43147];
assign t[43148] = t[43147] ^ n[43148];
assign t[43149] = t[43148] ^ n[43149];
assign t[43150] = t[43149] ^ n[43150];
assign t[43151] = t[43150] ^ n[43151];
assign t[43152] = t[43151] ^ n[43152];
assign t[43153] = t[43152] ^ n[43153];
assign t[43154] = t[43153] ^ n[43154];
assign t[43155] = t[43154] ^ n[43155];
assign t[43156] = t[43155] ^ n[43156];
assign t[43157] = t[43156] ^ n[43157];
assign t[43158] = t[43157] ^ n[43158];
assign t[43159] = t[43158] ^ n[43159];
assign t[43160] = t[43159] ^ n[43160];
assign t[43161] = t[43160] ^ n[43161];
assign t[43162] = t[43161] ^ n[43162];
assign t[43163] = t[43162] ^ n[43163];
assign t[43164] = t[43163] ^ n[43164];
assign t[43165] = t[43164] ^ n[43165];
assign t[43166] = t[43165] ^ n[43166];
assign t[43167] = t[43166] ^ n[43167];
assign t[43168] = t[43167] ^ n[43168];
assign t[43169] = t[43168] ^ n[43169];
assign t[43170] = t[43169] ^ n[43170];
assign t[43171] = t[43170] ^ n[43171];
assign t[43172] = t[43171] ^ n[43172];
assign t[43173] = t[43172] ^ n[43173];
assign t[43174] = t[43173] ^ n[43174];
assign t[43175] = t[43174] ^ n[43175];
assign t[43176] = t[43175] ^ n[43176];
assign t[43177] = t[43176] ^ n[43177];
assign t[43178] = t[43177] ^ n[43178];
assign t[43179] = t[43178] ^ n[43179];
assign t[43180] = t[43179] ^ n[43180];
assign t[43181] = t[43180] ^ n[43181];
assign t[43182] = t[43181] ^ n[43182];
assign t[43183] = t[43182] ^ n[43183];
assign t[43184] = t[43183] ^ n[43184];
assign t[43185] = t[43184] ^ n[43185];
assign t[43186] = t[43185] ^ n[43186];
assign t[43187] = t[43186] ^ n[43187];
assign t[43188] = t[43187] ^ n[43188];
assign t[43189] = t[43188] ^ n[43189];
assign t[43190] = t[43189] ^ n[43190];
assign t[43191] = t[43190] ^ n[43191];
assign t[43192] = t[43191] ^ n[43192];
assign t[43193] = t[43192] ^ n[43193];
assign t[43194] = t[43193] ^ n[43194];
assign t[43195] = t[43194] ^ n[43195];
assign t[43196] = t[43195] ^ n[43196];
assign t[43197] = t[43196] ^ n[43197];
assign t[43198] = t[43197] ^ n[43198];
assign t[43199] = t[43198] ^ n[43199];
assign t[43200] = t[43199] ^ n[43200];
assign t[43201] = t[43200] ^ n[43201];
assign t[43202] = t[43201] ^ n[43202];
assign t[43203] = t[43202] ^ n[43203];
assign t[43204] = t[43203] ^ n[43204];
assign t[43205] = t[43204] ^ n[43205];
assign t[43206] = t[43205] ^ n[43206];
assign t[43207] = t[43206] ^ n[43207];
assign t[43208] = t[43207] ^ n[43208];
assign t[43209] = t[43208] ^ n[43209];
assign t[43210] = t[43209] ^ n[43210];
assign t[43211] = t[43210] ^ n[43211];
assign t[43212] = t[43211] ^ n[43212];
assign t[43213] = t[43212] ^ n[43213];
assign t[43214] = t[43213] ^ n[43214];
assign t[43215] = t[43214] ^ n[43215];
assign t[43216] = t[43215] ^ n[43216];
assign t[43217] = t[43216] ^ n[43217];
assign t[43218] = t[43217] ^ n[43218];
assign t[43219] = t[43218] ^ n[43219];
assign t[43220] = t[43219] ^ n[43220];
assign t[43221] = t[43220] ^ n[43221];
assign t[43222] = t[43221] ^ n[43222];
assign t[43223] = t[43222] ^ n[43223];
assign t[43224] = t[43223] ^ n[43224];
assign t[43225] = t[43224] ^ n[43225];
assign t[43226] = t[43225] ^ n[43226];
assign t[43227] = t[43226] ^ n[43227];
assign t[43228] = t[43227] ^ n[43228];
assign t[43229] = t[43228] ^ n[43229];
assign t[43230] = t[43229] ^ n[43230];
assign t[43231] = t[43230] ^ n[43231];
assign t[43232] = t[43231] ^ n[43232];
assign t[43233] = t[43232] ^ n[43233];
assign t[43234] = t[43233] ^ n[43234];
assign t[43235] = t[43234] ^ n[43235];
assign t[43236] = t[43235] ^ n[43236];
assign t[43237] = t[43236] ^ n[43237];
assign t[43238] = t[43237] ^ n[43238];
assign t[43239] = t[43238] ^ n[43239];
assign t[43240] = t[43239] ^ n[43240];
assign t[43241] = t[43240] ^ n[43241];
assign t[43242] = t[43241] ^ n[43242];
assign t[43243] = t[43242] ^ n[43243];
assign t[43244] = t[43243] ^ n[43244];
assign t[43245] = t[43244] ^ n[43245];
assign t[43246] = t[43245] ^ n[43246];
assign t[43247] = t[43246] ^ n[43247];
assign t[43248] = t[43247] ^ n[43248];
assign t[43249] = t[43248] ^ n[43249];
assign t[43250] = t[43249] ^ n[43250];
assign t[43251] = t[43250] ^ n[43251];
assign t[43252] = t[43251] ^ n[43252];
assign t[43253] = t[43252] ^ n[43253];
assign t[43254] = t[43253] ^ n[43254];
assign t[43255] = t[43254] ^ n[43255];
assign t[43256] = t[43255] ^ n[43256];
assign t[43257] = t[43256] ^ n[43257];
assign t[43258] = t[43257] ^ n[43258];
assign t[43259] = t[43258] ^ n[43259];
assign t[43260] = t[43259] ^ n[43260];
assign t[43261] = t[43260] ^ n[43261];
assign t[43262] = t[43261] ^ n[43262];
assign t[43263] = t[43262] ^ n[43263];
assign t[43264] = t[43263] ^ n[43264];
assign t[43265] = t[43264] ^ n[43265];
assign t[43266] = t[43265] ^ n[43266];
assign t[43267] = t[43266] ^ n[43267];
assign t[43268] = t[43267] ^ n[43268];
assign t[43269] = t[43268] ^ n[43269];
assign t[43270] = t[43269] ^ n[43270];
assign t[43271] = t[43270] ^ n[43271];
assign t[43272] = t[43271] ^ n[43272];
assign t[43273] = t[43272] ^ n[43273];
assign t[43274] = t[43273] ^ n[43274];
assign t[43275] = t[43274] ^ n[43275];
assign t[43276] = t[43275] ^ n[43276];
assign t[43277] = t[43276] ^ n[43277];
assign t[43278] = t[43277] ^ n[43278];
assign t[43279] = t[43278] ^ n[43279];
assign t[43280] = t[43279] ^ n[43280];
assign t[43281] = t[43280] ^ n[43281];
assign t[43282] = t[43281] ^ n[43282];
assign t[43283] = t[43282] ^ n[43283];
assign t[43284] = t[43283] ^ n[43284];
assign t[43285] = t[43284] ^ n[43285];
assign t[43286] = t[43285] ^ n[43286];
assign t[43287] = t[43286] ^ n[43287];
assign t[43288] = t[43287] ^ n[43288];
assign t[43289] = t[43288] ^ n[43289];
assign t[43290] = t[43289] ^ n[43290];
assign t[43291] = t[43290] ^ n[43291];
assign t[43292] = t[43291] ^ n[43292];
assign t[43293] = t[43292] ^ n[43293];
assign t[43294] = t[43293] ^ n[43294];
assign t[43295] = t[43294] ^ n[43295];
assign t[43296] = t[43295] ^ n[43296];
assign t[43297] = t[43296] ^ n[43297];
assign t[43298] = t[43297] ^ n[43298];
assign t[43299] = t[43298] ^ n[43299];
assign t[43300] = t[43299] ^ n[43300];
assign t[43301] = t[43300] ^ n[43301];
assign t[43302] = t[43301] ^ n[43302];
assign t[43303] = t[43302] ^ n[43303];
assign t[43304] = t[43303] ^ n[43304];
assign t[43305] = t[43304] ^ n[43305];
assign t[43306] = t[43305] ^ n[43306];
assign t[43307] = t[43306] ^ n[43307];
assign t[43308] = t[43307] ^ n[43308];
assign t[43309] = t[43308] ^ n[43309];
assign t[43310] = t[43309] ^ n[43310];
assign t[43311] = t[43310] ^ n[43311];
assign t[43312] = t[43311] ^ n[43312];
assign t[43313] = t[43312] ^ n[43313];
assign t[43314] = t[43313] ^ n[43314];
assign t[43315] = t[43314] ^ n[43315];
assign t[43316] = t[43315] ^ n[43316];
assign t[43317] = t[43316] ^ n[43317];
assign t[43318] = t[43317] ^ n[43318];
assign t[43319] = t[43318] ^ n[43319];
assign t[43320] = t[43319] ^ n[43320];
assign t[43321] = t[43320] ^ n[43321];
assign t[43322] = t[43321] ^ n[43322];
assign t[43323] = t[43322] ^ n[43323];
assign t[43324] = t[43323] ^ n[43324];
assign t[43325] = t[43324] ^ n[43325];
assign t[43326] = t[43325] ^ n[43326];
assign t[43327] = t[43326] ^ n[43327];
assign t[43328] = t[43327] ^ n[43328];
assign t[43329] = t[43328] ^ n[43329];
assign t[43330] = t[43329] ^ n[43330];
assign t[43331] = t[43330] ^ n[43331];
assign t[43332] = t[43331] ^ n[43332];
assign t[43333] = t[43332] ^ n[43333];
assign t[43334] = t[43333] ^ n[43334];
assign t[43335] = t[43334] ^ n[43335];
assign t[43336] = t[43335] ^ n[43336];
assign t[43337] = t[43336] ^ n[43337];
assign t[43338] = t[43337] ^ n[43338];
assign t[43339] = t[43338] ^ n[43339];
assign t[43340] = t[43339] ^ n[43340];
assign t[43341] = t[43340] ^ n[43341];
assign t[43342] = t[43341] ^ n[43342];
assign t[43343] = t[43342] ^ n[43343];
assign t[43344] = t[43343] ^ n[43344];
assign t[43345] = t[43344] ^ n[43345];
assign t[43346] = t[43345] ^ n[43346];
assign t[43347] = t[43346] ^ n[43347];
assign t[43348] = t[43347] ^ n[43348];
assign t[43349] = t[43348] ^ n[43349];
assign t[43350] = t[43349] ^ n[43350];
assign t[43351] = t[43350] ^ n[43351];
assign t[43352] = t[43351] ^ n[43352];
assign t[43353] = t[43352] ^ n[43353];
assign t[43354] = t[43353] ^ n[43354];
assign t[43355] = t[43354] ^ n[43355];
assign t[43356] = t[43355] ^ n[43356];
assign t[43357] = t[43356] ^ n[43357];
assign t[43358] = t[43357] ^ n[43358];
assign t[43359] = t[43358] ^ n[43359];
assign t[43360] = t[43359] ^ n[43360];
assign t[43361] = t[43360] ^ n[43361];
assign t[43362] = t[43361] ^ n[43362];
assign t[43363] = t[43362] ^ n[43363];
assign t[43364] = t[43363] ^ n[43364];
assign t[43365] = t[43364] ^ n[43365];
assign t[43366] = t[43365] ^ n[43366];
assign t[43367] = t[43366] ^ n[43367];
assign t[43368] = t[43367] ^ n[43368];
assign t[43369] = t[43368] ^ n[43369];
assign t[43370] = t[43369] ^ n[43370];
assign t[43371] = t[43370] ^ n[43371];
assign t[43372] = t[43371] ^ n[43372];
assign t[43373] = t[43372] ^ n[43373];
assign t[43374] = t[43373] ^ n[43374];
assign t[43375] = t[43374] ^ n[43375];
assign t[43376] = t[43375] ^ n[43376];
assign t[43377] = t[43376] ^ n[43377];
assign t[43378] = t[43377] ^ n[43378];
assign t[43379] = t[43378] ^ n[43379];
assign t[43380] = t[43379] ^ n[43380];
assign t[43381] = t[43380] ^ n[43381];
assign t[43382] = t[43381] ^ n[43382];
assign t[43383] = t[43382] ^ n[43383];
assign t[43384] = t[43383] ^ n[43384];
assign t[43385] = t[43384] ^ n[43385];
assign t[43386] = t[43385] ^ n[43386];
assign t[43387] = t[43386] ^ n[43387];
assign t[43388] = t[43387] ^ n[43388];
assign t[43389] = t[43388] ^ n[43389];
assign t[43390] = t[43389] ^ n[43390];
assign t[43391] = t[43390] ^ n[43391];
assign t[43392] = t[43391] ^ n[43392];
assign t[43393] = t[43392] ^ n[43393];
assign t[43394] = t[43393] ^ n[43394];
assign t[43395] = t[43394] ^ n[43395];
assign t[43396] = t[43395] ^ n[43396];
assign t[43397] = t[43396] ^ n[43397];
assign t[43398] = t[43397] ^ n[43398];
assign t[43399] = t[43398] ^ n[43399];
assign t[43400] = t[43399] ^ n[43400];
assign t[43401] = t[43400] ^ n[43401];
assign t[43402] = t[43401] ^ n[43402];
assign t[43403] = t[43402] ^ n[43403];
assign t[43404] = t[43403] ^ n[43404];
assign t[43405] = t[43404] ^ n[43405];
assign t[43406] = t[43405] ^ n[43406];
assign t[43407] = t[43406] ^ n[43407];
assign t[43408] = t[43407] ^ n[43408];
assign t[43409] = t[43408] ^ n[43409];
assign t[43410] = t[43409] ^ n[43410];
assign t[43411] = t[43410] ^ n[43411];
assign t[43412] = t[43411] ^ n[43412];
assign t[43413] = t[43412] ^ n[43413];
assign t[43414] = t[43413] ^ n[43414];
assign t[43415] = t[43414] ^ n[43415];
assign t[43416] = t[43415] ^ n[43416];
assign t[43417] = t[43416] ^ n[43417];
assign t[43418] = t[43417] ^ n[43418];
assign t[43419] = t[43418] ^ n[43419];
assign t[43420] = t[43419] ^ n[43420];
assign t[43421] = t[43420] ^ n[43421];
assign t[43422] = t[43421] ^ n[43422];
assign t[43423] = t[43422] ^ n[43423];
assign t[43424] = t[43423] ^ n[43424];
assign t[43425] = t[43424] ^ n[43425];
assign t[43426] = t[43425] ^ n[43426];
assign t[43427] = t[43426] ^ n[43427];
assign t[43428] = t[43427] ^ n[43428];
assign t[43429] = t[43428] ^ n[43429];
assign t[43430] = t[43429] ^ n[43430];
assign t[43431] = t[43430] ^ n[43431];
assign t[43432] = t[43431] ^ n[43432];
assign t[43433] = t[43432] ^ n[43433];
assign t[43434] = t[43433] ^ n[43434];
assign t[43435] = t[43434] ^ n[43435];
assign t[43436] = t[43435] ^ n[43436];
assign t[43437] = t[43436] ^ n[43437];
assign t[43438] = t[43437] ^ n[43438];
assign t[43439] = t[43438] ^ n[43439];
assign t[43440] = t[43439] ^ n[43440];
assign t[43441] = t[43440] ^ n[43441];
assign t[43442] = t[43441] ^ n[43442];
assign t[43443] = t[43442] ^ n[43443];
assign t[43444] = t[43443] ^ n[43444];
assign t[43445] = t[43444] ^ n[43445];
assign t[43446] = t[43445] ^ n[43446];
assign t[43447] = t[43446] ^ n[43447];
assign t[43448] = t[43447] ^ n[43448];
assign t[43449] = t[43448] ^ n[43449];
assign t[43450] = t[43449] ^ n[43450];
assign t[43451] = t[43450] ^ n[43451];
assign t[43452] = t[43451] ^ n[43452];
assign t[43453] = t[43452] ^ n[43453];
assign t[43454] = t[43453] ^ n[43454];
assign t[43455] = t[43454] ^ n[43455];
assign t[43456] = t[43455] ^ n[43456];
assign t[43457] = t[43456] ^ n[43457];
assign t[43458] = t[43457] ^ n[43458];
assign t[43459] = t[43458] ^ n[43459];
assign t[43460] = t[43459] ^ n[43460];
assign t[43461] = t[43460] ^ n[43461];
assign t[43462] = t[43461] ^ n[43462];
assign t[43463] = t[43462] ^ n[43463];
assign t[43464] = t[43463] ^ n[43464];
assign t[43465] = t[43464] ^ n[43465];
assign t[43466] = t[43465] ^ n[43466];
assign t[43467] = t[43466] ^ n[43467];
assign t[43468] = t[43467] ^ n[43468];
assign t[43469] = t[43468] ^ n[43469];
assign t[43470] = t[43469] ^ n[43470];
assign t[43471] = t[43470] ^ n[43471];
assign t[43472] = t[43471] ^ n[43472];
assign t[43473] = t[43472] ^ n[43473];
assign t[43474] = t[43473] ^ n[43474];
assign t[43475] = t[43474] ^ n[43475];
assign t[43476] = t[43475] ^ n[43476];
assign t[43477] = t[43476] ^ n[43477];
assign t[43478] = t[43477] ^ n[43478];
assign t[43479] = t[43478] ^ n[43479];
assign t[43480] = t[43479] ^ n[43480];
assign t[43481] = t[43480] ^ n[43481];
assign t[43482] = t[43481] ^ n[43482];
assign t[43483] = t[43482] ^ n[43483];
assign t[43484] = t[43483] ^ n[43484];
assign t[43485] = t[43484] ^ n[43485];
assign t[43486] = t[43485] ^ n[43486];
assign t[43487] = t[43486] ^ n[43487];
assign t[43488] = t[43487] ^ n[43488];
assign t[43489] = t[43488] ^ n[43489];
assign t[43490] = t[43489] ^ n[43490];
assign t[43491] = t[43490] ^ n[43491];
assign t[43492] = t[43491] ^ n[43492];
assign t[43493] = t[43492] ^ n[43493];
assign t[43494] = t[43493] ^ n[43494];
assign t[43495] = t[43494] ^ n[43495];
assign t[43496] = t[43495] ^ n[43496];
assign t[43497] = t[43496] ^ n[43497];
assign t[43498] = t[43497] ^ n[43498];
assign t[43499] = t[43498] ^ n[43499];
assign t[43500] = t[43499] ^ n[43500];
assign t[43501] = t[43500] ^ n[43501];
assign t[43502] = t[43501] ^ n[43502];
assign t[43503] = t[43502] ^ n[43503];
assign t[43504] = t[43503] ^ n[43504];
assign t[43505] = t[43504] ^ n[43505];
assign t[43506] = t[43505] ^ n[43506];
assign t[43507] = t[43506] ^ n[43507];
assign t[43508] = t[43507] ^ n[43508];
assign t[43509] = t[43508] ^ n[43509];
assign t[43510] = t[43509] ^ n[43510];
assign t[43511] = t[43510] ^ n[43511];
assign t[43512] = t[43511] ^ n[43512];
assign t[43513] = t[43512] ^ n[43513];
assign t[43514] = t[43513] ^ n[43514];
assign t[43515] = t[43514] ^ n[43515];
assign t[43516] = t[43515] ^ n[43516];
assign t[43517] = t[43516] ^ n[43517];
assign t[43518] = t[43517] ^ n[43518];
assign t[43519] = t[43518] ^ n[43519];
assign t[43520] = t[43519] ^ n[43520];
assign t[43521] = t[43520] ^ n[43521];
assign t[43522] = t[43521] ^ n[43522];
assign t[43523] = t[43522] ^ n[43523];
assign t[43524] = t[43523] ^ n[43524];
assign t[43525] = t[43524] ^ n[43525];
assign t[43526] = t[43525] ^ n[43526];
assign t[43527] = t[43526] ^ n[43527];
assign t[43528] = t[43527] ^ n[43528];
assign t[43529] = t[43528] ^ n[43529];
assign t[43530] = t[43529] ^ n[43530];
assign t[43531] = t[43530] ^ n[43531];
assign t[43532] = t[43531] ^ n[43532];
assign t[43533] = t[43532] ^ n[43533];
assign t[43534] = t[43533] ^ n[43534];
assign t[43535] = t[43534] ^ n[43535];
assign t[43536] = t[43535] ^ n[43536];
assign t[43537] = t[43536] ^ n[43537];
assign t[43538] = t[43537] ^ n[43538];
assign t[43539] = t[43538] ^ n[43539];
assign t[43540] = t[43539] ^ n[43540];
assign t[43541] = t[43540] ^ n[43541];
assign t[43542] = t[43541] ^ n[43542];
assign t[43543] = t[43542] ^ n[43543];
assign t[43544] = t[43543] ^ n[43544];
assign t[43545] = t[43544] ^ n[43545];
assign t[43546] = t[43545] ^ n[43546];
assign t[43547] = t[43546] ^ n[43547];
assign t[43548] = t[43547] ^ n[43548];
assign t[43549] = t[43548] ^ n[43549];
assign t[43550] = t[43549] ^ n[43550];
assign t[43551] = t[43550] ^ n[43551];
assign t[43552] = t[43551] ^ n[43552];
assign t[43553] = t[43552] ^ n[43553];
assign t[43554] = t[43553] ^ n[43554];
assign t[43555] = t[43554] ^ n[43555];
assign t[43556] = t[43555] ^ n[43556];
assign t[43557] = t[43556] ^ n[43557];
assign t[43558] = t[43557] ^ n[43558];
assign t[43559] = t[43558] ^ n[43559];
assign t[43560] = t[43559] ^ n[43560];
assign t[43561] = t[43560] ^ n[43561];
assign t[43562] = t[43561] ^ n[43562];
assign t[43563] = t[43562] ^ n[43563];
assign t[43564] = t[43563] ^ n[43564];
assign t[43565] = t[43564] ^ n[43565];
assign t[43566] = t[43565] ^ n[43566];
assign t[43567] = t[43566] ^ n[43567];
assign t[43568] = t[43567] ^ n[43568];
assign t[43569] = t[43568] ^ n[43569];
assign t[43570] = t[43569] ^ n[43570];
assign t[43571] = t[43570] ^ n[43571];
assign t[43572] = t[43571] ^ n[43572];
assign t[43573] = t[43572] ^ n[43573];
assign t[43574] = t[43573] ^ n[43574];
assign t[43575] = t[43574] ^ n[43575];
assign t[43576] = t[43575] ^ n[43576];
assign t[43577] = t[43576] ^ n[43577];
assign t[43578] = t[43577] ^ n[43578];
assign t[43579] = t[43578] ^ n[43579];
assign t[43580] = t[43579] ^ n[43580];
assign t[43581] = t[43580] ^ n[43581];
assign t[43582] = t[43581] ^ n[43582];
assign t[43583] = t[43582] ^ n[43583];
assign t[43584] = t[43583] ^ n[43584];
assign t[43585] = t[43584] ^ n[43585];
assign t[43586] = t[43585] ^ n[43586];
assign t[43587] = t[43586] ^ n[43587];
assign t[43588] = t[43587] ^ n[43588];
assign t[43589] = t[43588] ^ n[43589];
assign t[43590] = t[43589] ^ n[43590];
assign t[43591] = t[43590] ^ n[43591];
assign t[43592] = t[43591] ^ n[43592];
assign t[43593] = t[43592] ^ n[43593];
assign t[43594] = t[43593] ^ n[43594];
assign t[43595] = t[43594] ^ n[43595];
assign t[43596] = t[43595] ^ n[43596];
assign t[43597] = t[43596] ^ n[43597];
assign t[43598] = t[43597] ^ n[43598];
assign t[43599] = t[43598] ^ n[43599];
assign t[43600] = t[43599] ^ n[43600];
assign t[43601] = t[43600] ^ n[43601];
assign t[43602] = t[43601] ^ n[43602];
assign t[43603] = t[43602] ^ n[43603];
assign t[43604] = t[43603] ^ n[43604];
assign t[43605] = t[43604] ^ n[43605];
assign t[43606] = t[43605] ^ n[43606];
assign t[43607] = t[43606] ^ n[43607];
assign t[43608] = t[43607] ^ n[43608];
assign t[43609] = t[43608] ^ n[43609];
assign t[43610] = t[43609] ^ n[43610];
assign t[43611] = t[43610] ^ n[43611];
assign t[43612] = t[43611] ^ n[43612];
assign t[43613] = t[43612] ^ n[43613];
assign t[43614] = t[43613] ^ n[43614];
assign t[43615] = t[43614] ^ n[43615];
assign t[43616] = t[43615] ^ n[43616];
assign t[43617] = t[43616] ^ n[43617];
assign t[43618] = t[43617] ^ n[43618];
assign t[43619] = t[43618] ^ n[43619];
assign t[43620] = t[43619] ^ n[43620];
assign t[43621] = t[43620] ^ n[43621];
assign t[43622] = t[43621] ^ n[43622];
assign t[43623] = t[43622] ^ n[43623];
assign t[43624] = t[43623] ^ n[43624];
assign t[43625] = t[43624] ^ n[43625];
assign t[43626] = t[43625] ^ n[43626];
assign t[43627] = t[43626] ^ n[43627];
assign t[43628] = t[43627] ^ n[43628];
assign t[43629] = t[43628] ^ n[43629];
assign t[43630] = t[43629] ^ n[43630];
assign t[43631] = t[43630] ^ n[43631];
assign t[43632] = t[43631] ^ n[43632];
assign t[43633] = t[43632] ^ n[43633];
assign t[43634] = t[43633] ^ n[43634];
assign t[43635] = t[43634] ^ n[43635];
assign t[43636] = t[43635] ^ n[43636];
assign t[43637] = t[43636] ^ n[43637];
assign t[43638] = t[43637] ^ n[43638];
assign t[43639] = t[43638] ^ n[43639];
assign t[43640] = t[43639] ^ n[43640];
assign t[43641] = t[43640] ^ n[43641];
assign t[43642] = t[43641] ^ n[43642];
assign t[43643] = t[43642] ^ n[43643];
assign t[43644] = t[43643] ^ n[43644];
assign t[43645] = t[43644] ^ n[43645];
assign t[43646] = t[43645] ^ n[43646];
assign t[43647] = t[43646] ^ n[43647];
assign t[43648] = t[43647] ^ n[43648];
assign t[43649] = t[43648] ^ n[43649];
assign t[43650] = t[43649] ^ n[43650];
assign t[43651] = t[43650] ^ n[43651];
assign t[43652] = t[43651] ^ n[43652];
assign t[43653] = t[43652] ^ n[43653];
assign t[43654] = t[43653] ^ n[43654];
assign t[43655] = t[43654] ^ n[43655];
assign t[43656] = t[43655] ^ n[43656];
assign t[43657] = t[43656] ^ n[43657];
assign t[43658] = t[43657] ^ n[43658];
assign t[43659] = t[43658] ^ n[43659];
assign t[43660] = t[43659] ^ n[43660];
assign t[43661] = t[43660] ^ n[43661];
assign t[43662] = t[43661] ^ n[43662];
assign t[43663] = t[43662] ^ n[43663];
assign t[43664] = t[43663] ^ n[43664];
assign t[43665] = t[43664] ^ n[43665];
assign t[43666] = t[43665] ^ n[43666];
assign t[43667] = t[43666] ^ n[43667];
assign t[43668] = t[43667] ^ n[43668];
assign t[43669] = t[43668] ^ n[43669];
assign t[43670] = t[43669] ^ n[43670];
assign t[43671] = t[43670] ^ n[43671];
assign t[43672] = t[43671] ^ n[43672];
assign t[43673] = t[43672] ^ n[43673];
assign t[43674] = t[43673] ^ n[43674];
assign t[43675] = t[43674] ^ n[43675];
assign t[43676] = t[43675] ^ n[43676];
assign t[43677] = t[43676] ^ n[43677];
assign t[43678] = t[43677] ^ n[43678];
assign t[43679] = t[43678] ^ n[43679];
assign t[43680] = t[43679] ^ n[43680];
assign t[43681] = t[43680] ^ n[43681];
assign t[43682] = t[43681] ^ n[43682];
assign t[43683] = t[43682] ^ n[43683];
assign t[43684] = t[43683] ^ n[43684];
assign t[43685] = t[43684] ^ n[43685];
assign t[43686] = t[43685] ^ n[43686];
assign t[43687] = t[43686] ^ n[43687];
assign t[43688] = t[43687] ^ n[43688];
assign t[43689] = t[43688] ^ n[43689];
assign t[43690] = t[43689] ^ n[43690];
assign t[43691] = t[43690] ^ n[43691];
assign t[43692] = t[43691] ^ n[43692];
assign t[43693] = t[43692] ^ n[43693];
assign t[43694] = t[43693] ^ n[43694];
assign t[43695] = t[43694] ^ n[43695];
assign t[43696] = t[43695] ^ n[43696];
assign t[43697] = t[43696] ^ n[43697];
assign t[43698] = t[43697] ^ n[43698];
assign t[43699] = t[43698] ^ n[43699];
assign t[43700] = t[43699] ^ n[43700];
assign t[43701] = t[43700] ^ n[43701];
assign t[43702] = t[43701] ^ n[43702];
assign t[43703] = t[43702] ^ n[43703];
assign t[43704] = t[43703] ^ n[43704];
assign t[43705] = t[43704] ^ n[43705];
assign t[43706] = t[43705] ^ n[43706];
assign t[43707] = t[43706] ^ n[43707];
assign t[43708] = t[43707] ^ n[43708];
assign t[43709] = t[43708] ^ n[43709];
assign t[43710] = t[43709] ^ n[43710];
assign t[43711] = t[43710] ^ n[43711];
assign t[43712] = t[43711] ^ n[43712];
assign t[43713] = t[43712] ^ n[43713];
assign t[43714] = t[43713] ^ n[43714];
assign t[43715] = t[43714] ^ n[43715];
assign t[43716] = t[43715] ^ n[43716];
assign t[43717] = t[43716] ^ n[43717];
assign t[43718] = t[43717] ^ n[43718];
assign t[43719] = t[43718] ^ n[43719];
assign t[43720] = t[43719] ^ n[43720];
assign t[43721] = t[43720] ^ n[43721];
assign t[43722] = t[43721] ^ n[43722];
assign t[43723] = t[43722] ^ n[43723];
assign t[43724] = t[43723] ^ n[43724];
assign t[43725] = t[43724] ^ n[43725];
assign t[43726] = t[43725] ^ n[43726];
assign t[43727] = t[43726] ^ n[43727];
assign t[43728] = t[43727] ^ n[43728];
assign t[43729] = t[43728] ^ n[43729];
assign t[43730] = t[43729] ^ n[43730];
assign t[43731] = t[43730] ^ n[43731];
assign t[43732] = t[43731] ^ n[43732];
assign t[43733] = t[43732] ^ n[43733];
assign t[43734] = t[43733] ^ n[43734];
assign t[43735] = t[43734] ^ n[43735];
assign t[43736] = t[43735] ^ n[43736];
assign t[43737] = t[43736] ^ n[43737];
assign t[43738] = t[43737] ^ n[43738];
assign t[43739] = t[43738] ^ n[43739];
assign t[43740] = t[43739] ^ n[43740];
assign t[43741] = t[43740] ^ n[43741];
assign t[43742] = t[43741] ^ n[43742];
assign t[43743] = t[43742] ^ n[43743];
assign t[43744] = t[43743] ^ n[43744];
assign t[43745] = t[43744] ^ n[43745];
assign t[43746] = t[43745] ^ n[43746];
assign t[43747] = t[43746] ^ n[43747];
assign t[43748] = t[43747] ^ n[43748];
assign t[43749] = t[43748] ^ n[43749];
assign t[43750] = t[43749] ^ n[43750];
assign t[43751] = t[43750] ^ n[43751];
assign t[43752] = t[43751] ^ n[43752];
assign t[43753] = t[43752] ^ n[43753];
assign t[43754] = t[43753] ^ n[43754];
assign t[43755] = t[43754] ^ n[43755];
assign t[43756] = t[43755] ^ n[43756];
assign t[43757] = t[43756] ^ n[43757];
assign t[43758] = t[43757] ^ n[43758];
assign t[43759] = t[43758] ^ n[43759];
assign t[43760] = t[43759] ^ n[43760];
assign t[43761] = t[43760] ^ n[43761];
assign t[43762] = t[43761] ^ n[43762];
assign t[43763] = t[43762] ^ n[43763];
assign t[43764] = t[43763] ^ n[43764];
assign t[43765] = t[43764] ^ n[43765];
assign t[43766] = t[43765] ^ n[43766];
assign t[43767] = t[43766] ^ n[43767];
assign t[43768] = t[43767] ^ n[43768];
assign t[43769] = t[43768] ^ n[43769];
assign t[43770] = t[43769] ^ n[43770];
assign t[43771] = t[43770] ^ n[43771];
assign t[43772] = t[43771] ^ n[43772];
assign t[43773] = t[43772] ^ n[43773];
assign t[43774] = t[43773] ^ n[43774];
assign t[43775] = t[43774] ^ n[43775];
assign t[43776] = t[43775] ^ n[43776];
assign t[43777] = t[43776] ^ n[43777];
assign t[43778] = t[43777] ^ n[43778];
assign t[43779] = t[43778] ^ n[43779];
assign t[43780] = t[43779] ^ n[43780];
assign t[43781] = t[43780] ^ n[43781];
assign t[43782] = t[43781] ^ n[43782];
assign t[43783] = t[43782] ^ n[43783];
assign t[43784] = t[43783] ^ n[43784];
assign t[43785] = t[43784] ^ n[43785];
assign t[43786] = t[43785] ^ n[43786];
assign t[43787] = t[43786] ^ n[43787];
assign t[43788] = t[43787] ^ n[43788];
assign t[43789] = t[43788] ^ n[43789];
assign t[43790] = t[43789] ^ n[43790];
assign t[43791] = t[43790] ^ n[43791];
assign t[43792] = t[43791] ^ n[43792];
assign t[43793] = t[43792] ^ n[43793];
assign t[43794] = t[43793] ^ n[43794];
assign t[43795] = t[43794] ^ n[43795];
assign t[43796] = t[43795] ^ n[43796];
assign t[43797] = t[43796] ^ n[43797];
assign t[43798] = t[43797] ^ n[43798];
assign t[43799] = t[43798] ^ n[43799];
assign t[43800] = t[43799] ^ n[43800];
assign t[43801] = t[43800] ^ n[43801];
assign t[43802] = t[43801] ^ n[43802];
assign t[43803] = t[43802] ^ n[43803];
assign t[43804] = t[43803] ^ n[43804];
assign t[43805] = t[43804] ^ n[43805];
assign t[43806] = t[43805] ^ n[43806];
assign t[43807] = t[43806] ^ n[43807];
assign t[43808] = t[43807] ^ n[43808];
assign t[43809] = t[43808] ^ n[43809];
assign t[43810] = t[43809] ^ n[43810];
assign t[43811] = t[43810] ^ n[43811];
assign t[43812] = t[43811] ^ n[43812];
assign t[43813] = t[43812] ^ n[43813];
assign t[43814] = t[43813] ^ n[43814];
assign t[43815] = t[43814] ^ n[43815];
assign t[43816] = t[43815] ^ n[43816];
assign t[43817] = t[43816] ^ n[43817];
assign t[43818] = t[43817] ^ n[43818];
assign t[43819] = t[43818] ^ n[43819];
assign t[43820] = t[43819] ^ n[43820];
assign t[43821] = t[43820] ^ n[43821];
assign t[43822] = t[43821] ^ n[43822];
assign t[43823] = t[43822] ^ n[43823];
assign t[43824] = t[43823] ^ n[43824];
assign t[43825] = t[43824] ^ n[43825];
assign t[43826] = t[43825] ^ n[43826];
assign t[43827] = t[43826] ^ n[43827];
assign t[43828] = t[43827] ^ n[43828];
assign t[43829] = t[43828] ^ n[43829];
assign t[43830] = t[43829] ^ n[43830];
assign t[43831] = t[43830] ^ n[43831];
assign t[43832] = t[43831] ^ n[43832];
assign t[43833] = t[43832] ^ n[43833];
assign t[43834] = t[43833] ^ n[43834];
assign t[43835] = t[43834] ^ n[43835];
assign t[43836] = t[43835] ^ n[43836];
assign t[43837] = t[43836] ^ n[43837];
assign t[43838] = t[43837] ^ n[43838];
assign t[43839] = t[43838] ^ n[43839];
assign t[43840] = t[43839] ^ n[43840];
assign t[43841] = t[43840] ^ n[43841];
assign t[43842] = t[43841] ^ n[43842];
assign t[43843] = t[43842] ^ n[43843];
assign t[43844] = t[43843] ^ n[43844];
assign t[43845] = t[43844] ^ n[43845];
assign t[43846] = t[43845] ^ n[43846];
assign t[43847] = t[43846] ^ n[43847];
assign t[43848] = t[43847] ^ n[43848];
assign t[43849] = t[43848] ^ n[43849];
assign t[43850] = t[43849] ^ n[43850];
assign t[43851] = t[43850] ^ n[43851];
assign t[43852] = t[43851] ^ n[43852];
assign t[43853] = t[43852] ^ n[43853];
assign t[43854] = t[43853] ^ n[43854];
assign t[43855] = t[43854] ^ n[43855];
assign t[43856] = t[43855] ^ n[43856];
assign t[43857] = t[43856] ^ n[43857];
assign t[43858] = t[43857] ^ n[43858];
assign t[43859] = t[43858] ^ n[43859];
assign t[43860] = t[43859] ^ n[43860];
assign t[43861] = t[43860] ^ n[43861];
assign t[43862] = t[43861] ^ n[43862];
assign t[43863] = t[43862] ^ n[43863];
assign t[43864] = t[43863] ^ n[43864];
assign t[43865] = t[43864] ^ n[43865];
assign t[43866] = t[43865] ^ n[43866];
assign t[43867] = t[43866] ^ n[43867];
assign t[43868] = t[43867] ^ n[43868];
assign t[43869] = t[43868] ^ n[43869];
assign t[43870] = t[43869] ^ n[43870];
assign t[43871] = t[43870] ^ n[43871];
assign t[43872] = t[43871] ^ n[43872];
assign t[43873] = t[43872] ^ n[43873];
assign t[43874] = t[43873] ^ n[43874];
assign t[43875] = t[43874] ^ n[43875];
assign t[43876] = t[43875] ^ n[43876];
assign t[43877] = t[43876] ^ n[43877];
assign t[43878] = t[43877] ^ n[43878];
assign t[43879] = t[43878] ^ n[43879];
assign t[43880] = t[43879] ^ n[43880];
assign t[43881] = t[43880] ^ n[43881];
assign t[43882] = t[43881] ^ n[43882];
assign t[43883] = t[43882] ^ n[43883];
assign t[43884] = t[43883] ^ n[43884];
assign t[43885] = t[43884] ^ n[43885];
assign t[43886] = t[43885] ^ n[43886];
assign t[43887] = t[43886] ^ n[43887];
assign t[43888] = t[43887] ^ n[43888];
assign t[43889] = t[43888] ^ n[43889];
assign t[43890] = t[43889] ^ n[43890];
assign t[43891] = t[43890] ^ n[43891];
assign t[43892] = t[43891] ^ n[43892];
assign t[43893] = t[43892] ^ n[43893];
assign t[43894] = t[43893] ^ n[43894];
assign t[43895] = t[43894] ^ n[43895];
assign t[43896] = t[43895] ^ n[43896];
assign t[43897] = t[43896] ^ n[43897];
assign t[43898] = t[43897] ^ n[43898];
assign t[43899] = t[43898] ^ n[43899];
assign t[43900] = t[43899] ^ n[43900];
assign t[43901] = t[43900] ^ n[43901];
assign t[43902] = t[43901] ^ n[43902];
assign t[43903] = t[43902] ^ n[43903];
assign t[43904] = t[43903] ^ n[43904];
assign t[43905] = t[43904] ^ n[43905];
assign t[43906] = t[43905] ^ n[43906];
assign t[43907] = t[43906] ^ n[43907];
assign t[43908] = t[43907] ^ n[43908];
assign t[43909] = t[43908] ^ n[43909];
assign t[43910] = t[43909] ^ n[43910];
assign t[43911] = t[43910] ^ n[43911];
assign t[43912] = t[43911] ^ n[43912];
assign t[43913] = t[43912] ^ n[43913];
assign t[43914] = t[43913] ^ n[43914];
assign t[43915] = t[43914] ^ n[43915];
assign t[43916] = t[43915] ^ n[43916];
assign t[43917] = t[43916] ^ n[43917];
assign t[43918] = t[43917] ^ n[43918];
assign t[43919] = t[43918] ^ n[43919];
assign t[43920] = t[43919] ^ n[43920];
assign t[43921] = t[43920] ^ n[43921];
assign t[43922] = t[43921] ^ n[43922];
assign t[43923] = t[43922] ^ n[43923];
assign t[43924] = t[43923] ^ n[43924];
assign t[43925] = t[43924] ^ n[43925];
assign t[43926] = t[43925] ^ n[43926];
assign t[43927] = t[43926] ^ n[43927];
assign t[43928] = t[43927] ^ n[43928];
assign t[43929] = t[43928] ^ n[43929];
assign t[43930] = t[43929] ^ n[43930];
assign t[43931] = t[43930] ^ n[43931];
assign t[43932] = t[43931] ^ n[43932];
assign t[43933] = t[43932] ^ n[43933];
assign t[43934] = t[43933] ^ n[43934];
assign t[43935] = t[43934] ^ n[43935];
assign t[43936] = t[43935] ^ n[43936];
assign t[43937] = t[43936] ^ n[43937];
assign t[43938] = t[43937] ^ n[43938];
assign t[43939] = t[43938] ^ n[43939];
assign t[43940] = t[43939] ^ n[43940];
assign t[43941] = t[43940] ^ n[43941];
assign t[43942] = t[43941] ^ n[43942];
assign t[43943] = t[43942] ^ n[43943];
assign t[43944] = t[43943] ^ n[43944];
assign t[43945] = t[43944] ^ n[43945];
assign t[43946] = t[43945] ^ n[43946];
assign t[43947] = t[43946] ^ n[43947];
assign t[43948] = t[43947] ^ n[43948];
assign t[43949] = t[43948] ^ n[43949];
assign t[43950] = t[43949] ^ n[43950];
assign t[43951] = t[43950] ^ n[43951];
assign t[43952] = t[43951] ^ n[43952];
assign t[43953] = t[43952] ^ n[43953];
assign t[43954] = t[43953] ^ n[43954];
assign t[43955] = t[43954] ^ n[43955];
assign t[43956] = t[43955] ^ n[43956];
assign t[43957] = t[43956] ^ n[43957];
assign t[43958] = t[43957] ^ n[43958];
assign t[43959] = t[43958] ^ n[43959];
assign t[43960] = t[43959] ^ n[43960];
assign t[43961] = t[43960] ^ n[43961];
assign t[43962] = t[43961] ^ n[43962];
assign t[43963] = t[43962] ^ n[43963];
assign t[43964] = t[43963] ^ n[43964];
assign t[43965] = t[43964] ^ n[43965];
assign t[43966] = t[43965] ^ n[43966];
assign t[43967] = t[43966] ^ n[43967];
assign t[43968] = t[43967] ^ n[43968];
assign t[43969] = t[43968] ^ n[43969];
assign t[43970] = t[43969] ^ n[43970];
assign t[43971] = t[43970] ^ n[43971];
assign t[43972] = t[43971] ^ n[43972];
assign t[43973] = t[43972] ^ n[43973];
assign t[43974] = t[43973] ^ n[43974];
assign t[43975] = t[43974] ^ n[43975];
assign t[43976] = t[43975] ^ n[43976];
assign t[43977] = t[43976] ^ n[43977];
assign t[43978] = t[43977] ^ n[43978];
assign t[43979] = t[43978] ^ n[43979];
assign t[43980] = t[43979] ^ n[43980];
assign t[43981] = t[43980] ^ n[43981];
assign t[43982] = t[43981] ^ n[43982];
assign t[43983] = t[43982] ^ n[43983];
assign t[43984] = t[43983] ^ n[43984];
assign t[43985] = t[43984] ^ n[43985];
assign t[43986] = t[43985] ^ n[43986];
assign t[43987] = t[43986] ^ n[43987];
assign t[43988] = t[43987] ^ n[43988];
assign t[43989] = t[43988] ^ n[43989];
assign t[43990] = t[43989] ^ n[43990];
assign t[43991] = t[43990] ^ n[43991];
assign t[43992] = t[43991] ^ n[43992];
assign t[43993] = t[43992] ^ n[43993];
assign t[43994] = t[43993] ^ n[43994];
assign t[43995] = t[43994] ^ n[43995];
assign t[43996] = t[43995] ^ n[43996];
assign t[43997] = t[43996] ^ n[43997];
assign t[43998] = t[43997] ^ n[43998];
assign t[43999] = t[43998] ^ n[43999];
assign t[44000] = t[43999] ^ n[44000];
assign t[44001] = t[44000] ^ n[44001];
assign t[44002] = t[44001] ^ n[44002];
assign t[44003] = t[44002] ^ n[44003];
assign t[44004] = t[44003] ^ n[44004];
assign t[44005] = t[44004] ^ n[44005];
assign t[44006] = t[44005] ^ n[44006];
assign t[44007] = t[44006] ^ n[44007];
assign t[44008] = t[44007] ^ n[44008];
assign t[44009] = t[44008] ^ n[44009];
assign t[44010] = t[44009] ^ n[44010];
assign t[44011] = t[44010] ^ n[44011];
assign t[44012] = t[44011] ^ n[44012];
assign t[44013] = t[44012] ^ n[44013];
assign t[44014] = t[44013] ^ n[44014];
assign t[44015] = t[44014] ^ n[44015];
assign t[44016] = t[44015] ^ n[44016];
assign t[44017] = t[44016] ^ n[44017];
assign t[44018] = t[44017] ^ n[44018];
assign t[44019] = t[44018] ^ n[44019];
assign t[44020] = t[44019] ^ n[44020];
assign t[44021] = t[44020] ^ n[44021];
assign t[44022] = t[44021] ^ n[44022];
assign t[44023] = t[44022] ^ n[44023];
assign t[44024] = t[44023] ^ n[44024];
assign t[44025] = t[44024] ^ n[44025];
assign t[44026] = t[44025] ^ n[44026];
assign t[44027] = t[44026] ^ n[44027];
assign t[44028] = t[44027] ^ n[44028];
assign t[44029] = t[44028] ^ n[44029];
assign t[44030] = t[44029] ^ n[44030];
assign t[44031] = t[44030] ^ n[44031];
assign t[44032] = t[44031] ^ n[44032];
assign t[44033] = t[44032] ^ n[44033];
assign t[44034] = t[44033] ^ n[44034];
assign t[44035] = t[44034] ^ n[44035];
assign t[44036] = t[44035] ^ n[44036];
assign t[44037] = t[44036] ^ n[44037];
assign t[44038] = t[44037] ^ n[44038];
assign t[44039] = t[44038] ^ n[44039];
assign t[44040] = t[44039] ^ n[44040];
assign t[44041] = t[44040] ^ n[44041];
assign t[44042] = t[44041] ^ n[44042];
assign t[44043] = t[44042] ^ n[44043];
assign t[44044] = t[44043] ^ n[44044];
assign t[44045] = t[44044] ^ n[44045];
assign t[44046] = t[44045] ^ n[44046];
assign t[44047] = t[44046] ^ n[44047];
assign t[44048] = t[44047] ^ n[44048];
assign t[44049] = t[44048] ^ n[44049];
assign t[44050] = t[44049] ^ n[44050];
assign t[44051] = t[44050] ^ n[44051];
assign t[44052] = t[44051] ^ n[44052];
assign t[44053] = t[44052] ^ n[44053];
assign t[44054] = t[44053] ^ n[44054];
assign t[44055] = t[44054] ^ n[44055];
assign t[44056] = t[44055] ^ n[44056];
assign t[44057] = t[44056] ^ n[44057];
assign t[44058] = t[44057] ^ n[44058];
assign t[44059] = t[44058] ^ n[44059];
assign t[44060] = t[44059] ^ n[44060];
assign t[44061] = t[44060] ^ n[44061];
assign t[44062] = t[44061] ^ n[44062];
assign t[44063] = t[44062] ^ n[44063];
assign t[44064] = t[44063] ^ n[44064];
assign t[44065] = t[44064] ^ n[44065];
assign t[44066] = t[44065] ^ n[44066];
assign t[44067] = t[44066] ^ n[44067];
assign t[44068] = t[44067] ^ n[44068];
assign t[44069] = t[44068] ^ n[44069];
assign t[44070] = t[44069] ^ n[44070];
assign t[44071] = t[44070] ^ n[44071];
assign t[44072] = t[44071] ^ n[44072];
assign t[44073] = t[44072] ^ n[44073];
assign t[44074] = t[44073] ^ n[44074];
assign t[44075] = t[44074] ^ n[44075];
assign t[44076] = t[44075] ^ n[44076];
assign t[44077] = t[44076] ^ n[44077];
assign t[44078] = t[44077] ^ n[44078];
assign t[44079] = t[44078] ^ n[44079];
assign t[44080] = t[44079] ^ n[44080];
assign t[44081] = t[44080] ^ n[44081];
assign t[44082] = t[44081] ^ n[44082];
assign t[44083] = t[44082] ^ n[44083];
assign t[44084] = t[44083] ^ n[44084];
assign t[44085] = t[44084] ^ n[44085];
assign t[44086] = t[44085] ^ n[44086];
assign t[44087] = t[44086] ^ n[44087];
assign t[44088] = t[44087] ^ n[44088];
assign t[44089] = t[44088] ^ n[44089];
assign t[44090] = t[44089] ^ n[44090];
assign t[44091] = t[44090] ^ n[44091];
assign t[44092] = t[44091] ^ n[44092];
assign t[44093] = t[44092] ^ n[44093];
assign t[44094] = t[44093] ^ n[44094];
assign t[44095] = t[44094] ^ n[44095];
assign t[44096] = t[44095] ^ n[44096];
assign t[44097] = t[44096] ^ n[44097];
assign t[44098] = t[44097] ^ n[44098];
assign t[44099] = t[44098] ^ n[44099];
assign t[44100] = t[44099] ^ n[44100];
assign t[44101] = t[44100] ^ n[44101];
assign t[44102] = t[44101] ^ n[44102];
assign t[44103] = t[44102] ^ n[44103];
assign t[44104] = t[44103] ^ n[44104];
assign t[44105] = t[44104] ^ n[44105];
assign t[44106] = t[44105] ^ n[44106];
assign t[44107] = t[44106] ^ n[44107];
assign t[44108] = t[44107] ^ n[44108];
assign t[44109] = t[44108] ^ n[44109];
assign t[44110] = t[44109] ^ n[44110];
assign t[44111] = t[44110] ^ n[44111];
assign t[44112] = t[44111] ^ n[44112];
assign t[44113] = t[44112] ^ n[44113];
assign t[44114] = t[44113] ^ n[44114];
assign t[44115] = t[44114] ^ n[44115];
assign t[44116] = t[44115] ^ n[44116];
assign t[44117] = t[44116] ^ n[44117];
assign t[44118] = t[44117] ^ n[44118];
assign t[44119] = t[44118] ^ n[44119];
assign t[44120] = t[44119] ^ n[44120];
assign t[44121] = t[44120] ^ n[44121];
assign t[44122] = t[44121] ^ n[44122];
assign t[44123] = t[44122] ^ n[44123];
assign t[44124] = t[44123] ^ n[44124];
assign t[44125] = t[44124] ^ n[44125];
assign t[44126] = t[44125] ^ n[44126];
assign t[44127] = t[44126] ^ n[44127];
assign t[44128] = t[44127] ^ n[44128];
assign t[44129] = t[44128] ^ n[44129];
assign t[44130] = t[44129] ^ n[44130];
assign t[44131] = t[44130] ^ n[44131];
assign t[44132] = t[44131] ^ n[44132];
assign t[44133] = t[44132] ^ n[44133];
assign t[44134] = t[44133] ^ n[44134];
assign t[44135] = t[44134] ^ n[44135];
assign t[44136] = t[44135] ^ n[44136];
assign t[44137] = t[44136] ^ n[44137];
assign t[44138] = t[44137] ^ n[44138];
assign t[44139] = t[44138] ^ n[44139];
assign t[44140] = t[44139] ^ n[44140];
assign t[44141] = t[44140] ^ n[44141];
assign t[44142] = t[44141] ^ n[44142];
assign t[44143] = t[44142] ^ n[44143];
assign t[44144] = t[44143] ^ n[44144];
assign t[44145] = t[44144] ^ n[44145];
assign t[44146] = t[44145] ^ n[44146];
assign t[44147] = t[44146] ^ n[44147];
assign t[44148] = t[44147] ^ n[44148];
assign t[44149] = t[44148] ^ n[44149];
assign t[44150] = t[44149] ^ n[44150];
assign t[44151] = t[44150] ^ n[44151];
assign t[44152] = t[44151] ^ n[44152];
assign t[44153] = t[44152] ^ n[44153];
assign t[44154] = t[44153] ^ n[44154];
assign t[44155] = t[44154] ^ n[44155];
assign t[44156] = t[44155] ^ n[44156];
assign t[44157] = t[44156] ^ n[44157];
assign t[44158] = t[44157] ^ n[44158];
assign t[44159] = t[44158] ^ n[44159];
assign t[44160] = t[44159] ^ n[44160];
assign t[44161] = t[44160] ^ n[44161];
assign t[44162] = t[44161] ^ n[44162];
assign t[44163] = t[44162] ^ n[44163];
assign t[44164] = t[44163] ^ n[44164];
assign t[44165] = t[44164] ^ n[44165];
assign t[44166] = t[44165] ^ n[44166];
assign t[44167] = t[44166] ^ n[44167];
assign t[44168] = t[44167] ^ n[44168];
assign t[44169] = t[44168] ^ n[44169];
assign t[44170] = t[44169] ^ n[44170];
assign t[44171] = t[44170] ^ n[44171];
assign t[44172] = t[44171] ^ n[44172];
assign t[44173] = t[44172] ^ n[44173];
assign t[44174] = t[44173] ^ n[44174];
assign t[44175] = t[44174] ^ n[44175];
assign t[44176] = t[44175] ^ n[44176];
assign t[44177] = t[44176] ^ n[44177];
assign t[44178] = t[44177] ^ n[44178];
assign t[44179] = t[44178] ^ n[44179];
assign t[44180] = t[44179] ^ n[44180];
assign t[44181] = t[44180] ^ n[44181];
assign t[44182] = t[44181] ^ n[44182];
assign t[44183] = t[44182] ^ n[44183];
assign t[44184] = t[44183] ^ n[44184];
assign t[44185] = t[44184] ^ n[44185];
assign t[44186] = t[44185] ^ n[44186];
assign t[44187] = t[44186] ^ n[44187];
assign t[44188] = t[44187] ^ n[44188];
assign t[44189] = t[44188] ^ n[44189];
assign t[44190] = t[44189] ^ n[44190];
assign t[44191] = t[44190] ^ n[44191];
assign t[44192] = t[44191] ^ n[44192];
assign t[44193] = t[44192] ^ n[44193];
assign t[44194] = t[44193] ^ n[44194];
assign t[44195] = t[44194] ^ n[44195];
assign t[44196] = t[44195] ^ n[44196];
assign t[44197] = t[44196] ^ n[44197];
assign t[44198] = t[44197] ^ n[44198];
assign t[44199] = t[44198] ^ n[44199];
assign t[44200] = t[44199] ^ n[44200];
assign t[44201] = t[44200] ^ n[44201];
assign t[44202] = t[44201] ^ n[44202];
assign t[44203] = t[44202] ^ n[44203];
assign t[44204] = t[44203] ^ n[44204];
assign t[44205] = t[44204] ^ n[44205];
assign t[44206] = t[44205] ^ n[44206];
assign t[44207] = t[44206] ^ n[44207];
assign t[44208] = t[44207] ^ n[44208];
assign t[44209] = t[44208] ^ n[44209];
assign t[44210] = t[44209] ^ n[44210];
assign t[44211] = t[44210] ^ n[44211];
assign t[44212] = t[44211] ^ n[44212];
assign t[44213] = t[44212] ^ n[44213];
assign t[44214] = t[44213] ^ n[44214];
assign t[44215] = t[44214] ^ n[44215];
assign t[44216] = t[44215] ^ n[44216];
assign t[44217] = t[44216] ^ n[44217];
assign t[44218] = t[44217] ^ n[44218];
assign t[44219] = t[44218] ^ n[44219];
assign t[44220] = t[44219] ^ n[44220];
assign t[44221] = t[44220] ^ n[44221];
assign t[44222] = t[44221] ^ n[44222];
assign t[44223] = t[44222] ^ n[44223];
assign t[44224] = t[44223] ^ n[44224];
assign t[44225] = t[44224] ^ n[44225];
assign t[44226] = t[44225] ^ n[44226];
assign t[44227] = t[44226] ^ n[44227];
assign t[44228] = t[44227] ^ n[44228];
assign t[44229] = t[44228] ^ n[44229];
assign t[44230] = t[44229] ^ n[44230];
assign t[44231] = t[44230] ^ n[44231];
assign t[44232] = t[44231] ^ n[44232];
assign t[44233] = t[44232] ^ n[44233];
assign t[44234] = t[44233] ^ n[44234];
assign t[44235] = t[44234] ^ n[44235];
assign t[44236] = t[44235] ^ n[44236];
assign t[44237] = t[44236] ^ n[44237];
assign t[44238] = t[44237] ^ n[44238];
assign t[44239] = t[44238] ^ n[44239];
assign t[44240] = t[44239] ^ n[44240];
assign t[44241] = t[44240] ^ n[44241];
assign t[44242] = t[44241] ^ n[44242];
assign t[44243] = t[44242] ^ n[44243];
assign t[44244] = t[44243] ^ n[44244];
assign t[44245] = t[44244] ^ n[44245];
assign t[44246] = t[44245] ^ n[44246];
assign t[44247] = t[44246] ^ n[44247];
assign t[44248] = t[44247] ^ n[44248];
assign t[44249] = t[44248] ^ n[44249];
assign t[44250] = t[44249] ^ n[44250];
assign t[44251] = t[44250] ^ n[44251];
assign t[44252] = t[44251] ^ n[44252];
assign t[44253] = t[44252] ^ n[44253];
assign t[44254] = t[44253] ^ n[44254];
assign t[44255] = t[44254] ^ n[44255];
assign t[44256] = t[44255] ^ n[44256];
assign t[44257] = t[44256] ^ n[44257];
assign t[44258] = t[44257] ^ n[44258];
assign t[44259] = t[44258] ^ n[44259];
assign t[44260] = t[44259] ^ n[44260];
assign t[44261] = t[44260] ^ n[44261];
assign t[44262] = t[44261] ^ n[44262];
assign t[44263] = t[44262] ^ n[44263];
assign t[44264] = t[44263] ^ n[44264];
assign t[44265] = t[44264] ^ n[44265];
assign t[44266] = t[44265] ^ n[44266];
assign t[44267] = t[44266] ^ n[44267];
assign t[44268] = t[44267] ^ n[44268];
assign t[44269] = t[44268] ^ n[44269];
assign t[44270] = t[44269] ^ n[44270];
assign t[44271] = t[44270] ^ n[44271];
assign t[44272] = t[44271] ^ n[44272];
assign t[44273] = t[44272] ^ n[44273];
assign t[44274] = t[44273] ^ n[44274];
assign t[44275] = t[44274] ^ n[44275];
assign t[44276] = t[44275] ^ n[44276];
assign t[44277] = t[44276] ^ n[44277];
assign t[44278] = t[44277] ^ n[44278];
assign t[44279] = t[44278] ^ n[44279];
assign t[44280] = t[44279] ^ n[44280];
assign t[44281] = t[44280] ^ n[44281];
assign t[44282] = t[44281] ^ n[44282];
assign t[44283] = t[44282] ^ n[44283];
assign t[44284] = t[44283] ^ n[44284];
assign t[44285] = t[44284] ^ n[44285];
assign t[44286] = t[44285] ^ n[44286];
assign t[44287] = t[44286] ^ n[44287];
assign t[44288] = t[44287] ^ n[44288];
assign t[44289] = t[44288] ^ n[44289];
assign t[44290] = t[44289] ^ n[44290];
assign t[44291] = t[44290] ^ n[44291];
assign t[44292] = t[44291] ^ n[44292];
assign t[44293] = t[44292] ^ n[44293];
assign t[44294] = t[44293] ^ n[44294];
assign t[44295] = t[44294] ^ n[44295];
assign t[44296] = t[44295] ^ n[44296];
assign t[44297] = t[44296] ^ n[44297];
assign t[44298] = t[44297] ^ n[44298];
assign t[44299] = t[44298] ^ n[44299];
assign t[44300] = t[44299] ^ n[44300];
assign t[44301] = t[44300] ^ n[44301];
assign t[44302] = t[44301] ^ n[44302];
assign t[44303] = t[44302] ^ n[44303];
assign t[44304] = t[44303] ^ n[44304];
assign t[44305] = t[44304] ^ n[44305];
assign t[44306] = t[44305] ^ n[44306];
assign t[44307] = t[44306] ^ n[44307];
assign t[44308] = t[44307] ^ n[44308];
assign t[44309] = t[44308] ^ n[44309];
assign t[44310] = t[44309] ^ n[44310];
assign t[44311] = t[44310] ^ n[44311];
assign t[44312] = t[44311] ^ n[44312];
assign t[44313] = t[44312] ^ n[44313];
assign t[44314] = t[44313] ^ n[44314];
assign t[44315] = t[44314] ^ n[44315];
assign t[44316] = t[44315] ^ n[44316];
assign t[44317] = t[44316] ^ n[44317];
assign t[44318] = t[44317] ^ n[44318];
assign t[44319] = t[44318] ^ n[44319];
assign t[44320] = t[44319] ^ n[44320];
assign t[44321] = t[44320] ^ n[44321];
assign t[44322] = t[44321] ^ n[44322];
assign t[44323] = t[44322] ^ n[44323];
assign t[44324] = t[44323] ^ n[44324];
assign t[44325] = t[44324] ^ n[44325];
assign t[44326] = t[44325] ^ n[44326];
assign t[44327] = t[44326] ^ n[44327];
assign t[44328] = t[44327] ^ n[44328];
assign t[44329] = t[44328] ^ n[44329];
assign t[44330] = t[44329] ^ n[44330];
assign t[44331] = t[44330] ^ n[44331];
assign t[44332] = t[44331] ^ n[44332];
assign t[44333] = t[44332] ^ n[44333];
assign t[44334] = t[44333] ^ n[44334];
assign t[44335] = t[44334] ^ n[44335];
assign t[44336] = t[44335] ^ n[44336];
assign t[44337] = t[44336] ^ n[44337];
assign t[44338] = t[44337] ^ n[44338];
assign t[44339] = t[44338] ^ n[44339];
assign t[44340] = t[44339] ^ n[44340];
assign t[44341] = t[44340] ^ n[44341];
assign t[44342] = t[44341] ^ n[44342];
assign t[44343] = t[44342] ^ n[44343];
assign t[44344] = t[44343] ^ n[44344];
assign t[44345] = t[44344] ^ n[44345];
assign t[44346] = t[44345] ^ n[44346];
assign t[44347] = t[44346] ^ n[44347];
assign t[44348] = t[44347] ^ n[44348];
assign t[44349] = t[44348] ^ n[44349];
assign t[44350] = t[44349] ^ n[44350];
assign t[44351] = t[44350] ^ n[44351];
assign t[44352] = t[44351] ^ n[44352];
assign t[44353] = t[44352] ^ n[44353];
assign t[44354] = t[44353] ^ n[44354];
assign t[44355] = t[44354] ^ n[44355];
assign t[44356] = t[44355] ^ n[44356];
assign t[44357] = t[44356] ^ n[44357];
assign t[44358] = t[44357] ^ n[44358];
assign t[44359] = t[44358] ^ n[44359];
assign t[44360] = t[44359] ^ n[44360];
assign t[44361] = t[44360] ^ n[44361];
assign t[44362] = t[44361] ^ n[44362];
assign t[44363] = t[44362] ^ n[44363];
assign t[44364] = t[44363] ^ n[44364];
assign t[44365] = t[44364] ^ n[44365];
assign t[44366] = t[44365] ^ n[44366];
assign t[44367] = t[44366] ^ n[44367];
assign t[44368] = t[44367] ^ n[44368];
assign t[44369] = t[44368] ^ n[44369];
assign t[44370] = t[44369] ^ n[44370];
assign t[44371] = t[44370] ^ n[44371];
assign t[44372] = t[44371] ^ n[44372];
assign t[44373] = t[44372] ^ n[44373];
assign t[44374] = t[44373] ^ n[44374];
assign t[44375] = t[44374] ^ n[44375];
assign t[44376] = t[44375] ^ n[44376];
assign t[44377] = t[44376] ^ n[44377];
assign t[44378] = t[44377] ^ n[44378];
assign t[44379] = t[44378] ^ n[44379];
assign t[44380] = t[44379] ^ n[44380];
assign t[44381] = t[44380] ^ n[44381];
assign t[44382] = t[44381] ^ n[44382];
assign t[44383] = t[44382] ^ n[44383];
assign t[44384] = t[44383] ^ n[44384];
assign t[44385] = t[44384] ^ n[44385];
assign t[44386] = t[44385] ^ n[44386];
assign t[44387] = t[44386] ^ n[44387];
assign t[44388] = t[44387] ^ n[44388];
assign t[44389] = t[44388] ^ n[44389];
assign t[44390] = t[44389] ^ n[44390];
assign t[44391] = t[44390] ^ n[44391];
assign t[44392] = t[44391] ^ n[44392];
assign t[44393] = t[44392] ^ n[44393];
assign t[44394] = t[44393] ^ n[44394];
assign t[44395] = t[44394] ^ n[44395];
assign t[44396] = t[44395] ^ n[44396];
assign t[44397] = t[44396] ^ n[44397];
assign t[44398] = t[44397] ^ n[44398];
assign t[44399] = t[44398] ^ n[44399];
assign t[44400] = t[44399] ^ n[44400];
assign t[44401] = t[44400] ^ n[44401];
assign t[44402] = t[44401] ^ n[44402];
assign t[44403] = t[44402] ^ n[44403];
assign t[44404] = t[44403] ^ n[44404];
assign t[44405] = t[44404] ^ n[44405];
assign t[44406] = t[44405] ^ n[44406];
assign t[44407] = t[44406] ^ n[44407];
assign t[44408] = t[44407] ^ n[44408];
assign t[44409] = t[44408] ^ n[44409];
assign t[44410] = t[44409] ^ n[44410];
assign t[44411] = t[44410] ^ n[44411];
assign t[44412] = t[44411] ^ n[44412];
assign t[44413] = t[44412] ^ n[44413];
assign t[44414] = t[44413] ^ n[44414];
assign t[44415] = t[44414] ^ n[44415];
assign t[44416] = t[44415] ^ n[44416];
assign t[44417] = t[44416] ^ n[44417];
assign t[44418] = t[44417] ^ n[44418];
assign t[44419] = t[44418] ^ n[44419];
assign t[44420] = t[44419] ^ n[44420];
assign t[44421] = t[44420] ^ n[44421];
assign t[44422] = t[44421] ^ n[44422];
assign t[44423] = t[44422] ^ n[44423];
assign t[44424] = t[44423] ^ n[44424];
assign t[44425] = t[44424] ^ n[44425];
assign t[44426] = t[44425] ^ n[44426];
assign t[44427] = t[44426] ^ n[44427];
assign t[44428] = t[44427] ^ n[44428];
assign t[44429] = t[44428] ^ n[44429];
assign t[44430] = t[44429] ^ n[44430];
assign t[44431] = t[44430] ^ n[44431];
assign t[44432] = t[44431] ^ n[44432];
assign t[44433] = t[44432] ^ n[44433];
assign t[44434] = t[44433] ^ n[44434];
assign t[44435] = t[44434] ^ n[44435];
assign t[44436] = t[44435] ^ n[44436];
assign t[44437] = t[44436] ^ n[44437];
assign t[44438] = t[44437] ^ n[44438];
assign t[44439] = t[44438] ^ n[44439];
assign t[44440] = t[44439] ^ n[44440];
assign t[44441] = t[44440] ^ n[44441];
assign t[44442] = t[44441] ^ n[44442];
assign t[44443] = t[44442] ^ n[44443];
assign t[44444] = t[44443] ^ n[44444];
assign t[44445] = t[44444] ^ n[44445];
assign t[44446] = t[44445] ^ n[44446];
assign t[44447] = t[44446] ^ n[44447];
assign t[44448] = t[44447] ^ n[44448];
assign t[44449] = t[44448] ^ n[44449];
assign t[44450] = t[44449] ^ n[44450];
assign t[44451] = t[44450] ^ n[44451];
assign t[44452] = t[44451] ^ n[44452];
assign t[44453] = t[44452] ^ n[44453];
assign t[44454] = t[44453] ^ n[44454];
assign t[44455] = t[44454] ^ n[44455];
assign t[44456] = t[44455] ^ n[44456];
assign t[44457] = t[44456] ^ n[44457];
assign t[44458] = t[44457] ^ n[44458];
assign t[44459] = t[44458] ^ n[44459];
assign t[44460] = t[44459] ^ n[44460];
assign t[44461] = t[44460] ^ n[44461];
assign t[44462] = t[44461] ^ n[44462];
assign t[44463] = t[44462] ^ n[44463];
assign t[44464] = t[44463] ^ n[44464];
assign t[44465] = t[44464] ^ n[44465];
assign t[44466] = t[44465] ^ n[44466];
assign t[44467] = t[44466] ^ n[44467];
assign t[44468] = t[44467] ^ n[44468];
assign t[44469] = t[44468] ^ n[44469];
assign t[44470] = t[44469] ^ n[44470];
assign t[44471] = t[44470] ^ n[44471];
assign t[44472] = t[44471] ^ n[44472];
assign t[44473] = t[44472] ^ n[44473];
assign t[44474] = t[44473] ^ n[44474];
assign t[44475] = t[44474] ^ n[44475];
assign t[44476] = t[44475] ^ n[44476];
assign t[44477] = t[44476] ^ n[44477];
assign t[44478] = t[44477] ^ n[44478];
assign t[44479] = t[44478] ^ n[44479];
assign t[44480] = t[44479] ^ n[44480];
assign t[44481] = t[44480] ^ n[44481];
assign t[44482] = t[44481] ^ n[44482];
assign t[44483] = t[44482] ^ n[44483];
assign t[44484] = t[44483] ^ n[44484];
assign t[44485] = t[44484] ^ n[44485];
assign t[44486] = t[44485] ^ n[44486];
assign t[44487] = t[44486] ^ n[44487];
assign t[44488] = t[44487] ^ n[44488];
assign t[44489] = t[44488] ^ n[44489];
assign t[44490] = t[44489] ^ n[44490];
assign t[44491] = t[44490] ^ n[44491];
assign t[44492] = t[44491] ^ n[44492];
assign t[44493] = t[44492] ^ n[44493];
assign t[44494] = t[44493] ^ n[44494];
assign t[44495] = t[44494] ^ n[44495];
assign t[44496] = t[44495] ^ n[44496];
assign t[44497] = t[44496] ^ n[44497];
assign t[44498] = t[44497] ^ n[44498];
assign t[44499] = t[44498] ^ n[44499];
assign t[44500] = t[44499] ^ n[44500];
assign t[44501] = t[44500] ^ n[44501];
assign t[44502] = t[44501] ^ n[44502];
assign t[44503] = t[44502] ^ n[44503];
assign t[44504] = t[44503] ^ n[44504];
assign t[44505] = t[44504] ^ n[44505];
assign t[44506] = t[44505] ^ n[44506];
assign t[44507] = t[44506] ^ n[44507];
assign t[44508] = t[44507] ^ n[44508];
assign t[44509] = t[44508] ^ n[44509];
assign t[44510] = t[44509] ^ n[44510];
assign t[44511] = t[44510] ^ n[44511];
assign t[44512] = t[44511] ^ n[44512];
assign t[44513] = t[44512] ^ n[44513];
assign t[44514] = t[44513] ^ n[44514];
assign t[44515] = t[44514] ^ n[44515];
assign t[44516] = t[44515] ^ n[44516];
assign t[44517] = t[44516] ^ n[44517];
assign t[44518] = t[44517] ^ n[44518];
assign t[44519] = t[44518] ^ n[44519];
assign t[44520] = t[44519] ^ n[44520];
assign t[44521] = t[44520] ^ n[44521];
assign t[44522] = t[44521] ^ n[44522];
assign t[44523] = t[44522] ^ n[44523];
assign t[44524] = t[44523] ^ n[44524];
assign t[44525] = t[44524] ^ n[44525];
assign t[44526] = t[44525] ^ n[44526];
assign t[44527] = t[44526] ^ n[44527];
assign t[44528] = t[44527] ^ n[44528];
assign t[44529] = t[44528] ^ n[44529];
assign t[44530] = t[44529] ^ n[44530];
assign t[44531] = t[44530] ^ n[44531];
assign t[44532] = t[44531] ^ n[44532];
assign t[44533] = t[44532] ^ n[44533];
assign t[44534] = t[44533] ^ n[44534];
assign t[44535] = t[44534] ^ n[44535];
assign t[44536] = t[44535] ^ n[44536];
assign t[44537] = t[44536] ^ n[44537];
assign t[44538] = t[44537] ^ n[44538];
assign t[44539] = t[44538] ^ n[44539];
assign t[44540] = t[44539] ^ n[44540];
assign t[44541] = t[44540] ^ n[44541];
assign t[44542] = t[44541] ^ n[44542];
assign t[44543] = t[44542] ^ n[44543];
assign t[44544] = t[44543] ^ n[44544];
assign t[44545] = t[44544] ^ n[44545];
assign t[44546] = t[44545] ^ n[44546];
assign t[44547] = t[44546] ^ n[44547];
assign t[44548] = t[44547] ^ n[44548];
assign t[44549] = t[44548] ^ n[44549];
assign t[44550] = t[44549] ^ n[44550];
assign t[44551] = t[44550] ^ n[44551];
assign t[44552] = t[44551] ^ n[44552];
assign t[44553] = t[44552] ^ n[44553];
assign t[44554] = t[44553] ^ n[44554];
assign t[44555] = t[44554] ^ n[44555];
assign t[44556] = t[44555] ^ n[44556];
assign t[44557] = t[44556] ^ n[44557];
assign t[44558] = t[44557] ^ n[44558];
assign t[44559] = t[44558] ^ n[44559];
assign t[44560] = t[44559] ^ n[44560];
assign t[44561] = t[44560] ^ n[44561];
assign t[44562] = t[44561] ^ n[44562];
assign t[44563] = t[44562] ^ n[44563];
assign t[44564] = t[44563] ^ n[44564];
assign t[44565] = t[44564] ^ n[44565];
assign t[44566] = t[44565] ^ n[44566];
assign t[44567] = t[44566] ^ n[44567];
assign t[44568] = t[44567] ^ n[44568];
assign t[44569] = t[44568] ^ n[44569];
assign t[44570] = t[44569] ^ n[44570];
assign t[44571] = t[44570] ^ n[44571];
assign t[44572] = t[44571] ^ n[44572];
assign t[44573] = t[44572] ^ n[44573];
assign t[44574] = t[44573] ^ n[44574];
assign t[44575] = t[44574] ^ n[44575];
assign t[44576] = t[44575] ^ n[44576];
assign t[44577] = t[44576] ^ n[44577];
assign t[44578] = t[44577] ^ n[44578];
assign t[44579] = t[44578] ^ n[44579];
assign t[44580] = t[44579] ^ n[44580];
assign t[44581] = t[44580] ^ n[44581];
assign t[44582] = t[44581] ^ n[44582];
assign t[44583] = t[44582] ^ n[44583];
assign t[44584] = t[44583] ^ n[44584];
assign t[44585] = t[44584] ^ n[44585];
assign t[44586] = t[44585] ^ n[44586];
assign t[44587] = t[44586] ^ n[44587];
assign t[44588] = t[44587] ^ n[44588];
assign t[44589] = t[44588] ^ n[44589];
assign t[44590] = t[44589] ^ n[44590];
assign t[44591] = t[44590] ^ n[44591];
assign t[44592] = t[44591] ^ n[44592];
assign t[44593] = t[44592] ^ n[44593];
assign t[44594] = t[44593] ^ n[44594];
assign t[44595] = t[44594] ^ n[44595];
assign t[44596] = t[44595] ^ n[44596];
assign t[44597] = t[44596] ^ n[44597];
assign t[44598] = t[44597] ^ n[44598];
assign t[44599] = t[44598] ^ n[44599];
assign t[44600] = t[44599] ^ n[44600];
assign t[44601] = t[44600] ^ n[44601];
assign t[44602] = t[44601] ^ n[44602];
assign t[44603] = t[44602] ^ n[44603];
assign t[44604] = t[44603] ^ n[44604];
assign t[44605] = t[44604] ^ n[44605];
assign t[44606] = t[44605] ^ n[44606];
assign t[44607] = t[44606] ^ n[44607];
assign t[44608] = t[44607] ^ n[44608];
assign t[44609] = t[44608] ^ n[44609];
assign t[44610] = t[44609] ^ n[44610];
assign t[44611] = t[44610] ^ n[44611];
assign t[44612] = t[44611] ^ n[44612];
assign t[44613] = t[44612] ^ n[44613];
assign t[44614] = t[44613] ^ n[44614];
assign t[44615] = t[44614] ^ n[44615];
assign t[44616] = t[44615] ^ n[44616];
assign t[44617] = t[44616] ^ n[44617];
assign t[44618] = t[44617] ^ n[44618];
assign t[44619] = t[44618] ^ n[44619];
assign t[44620] = t[44619] ^ n[44620];
assign t[44621] = t[44620] ^ n[44621];
assign t[44622] = t[44621] ^ n[44622];
assign t[44623] = t[44622] ^ n[44623];
assign t[44624] = t[44623] ^ n[44624];
assign t[44625] = t[44624] ^ n[44625];
assign t[44626] = t[44625] ^ n[44626];
assign t[44627] = t[44626] ^ n[44627];
assign t[44628] = t[44627] ^ n[44628];
assign t[44629] = t[44628] ^ n[44629];
assign t[44630] = t[44629] ^ n[44630];
assign t[44631] = t[44630] ^ n[44631];
assign t[44632] = t[44631] ^ n[44632];
assign t[44633] = t[44632] ^ n[44633];
assign t[44634] = t[44633] ^ n[44634];
assign t[44635] = t[44634] ^ n[44635];
assign t[44636] = t[44635] ^ n[44636];
assign t[44637] = t[44636] ^ n[44637];
assign t[44638] = t[44637] ^ n[44638];
assign t[44639] = t[44638] ^ n[44639];
assign t[44640] = t[44639] ^ n[44640];
assign t[44641] = t[44640] ^ n[44641];
assign t[44642] = t[44641] ^ n[44642];
assign t[44643] = t[44642] ^ n[44643];
assign t[44644] = t[44643] ^ n[44644];
assign t[44645] = t[44644] ^ n[44645];
assign t[44646] = t[44645] ^ n[44646];
assign t[44647] = t[44646] ^ n[44647];
assign t[44648] = t[44647] ^ n[44648];
assign t[44649] = t[44648] ^ n[44649];
assign t[44650] = t[44649] ^ n[44650];
assign t[44651] = t[44650] ^ n[44651];
assign t[44652] = t[44651] ^ n[44652];
assign t[44653] = t[44652] ^ n[44653];
assign t[44654] = t[44653] ^ n[44654];
assign t[44655] = t[44654] ^ n[44655];
assign t[44656] = t[44655] ^ n[44656];
assign t[44657] = t[44656] ^ n[44657];
assign t[44658] = t[44657] ^ n[44658];
assign t[44659] = t[44658] ^ n[44659];
assign t[44660] = t[44659] ^ n[44660];
assign t[44661] = t[44660] ^ n[44661];
assign t[44662] = t[44661] ^ n[44662];
assign t[44663] = t[44662] ^ n[44663];
assign t[44664] = t[44663] ^ n[44664];
assign t[44665] = t[44664] ^ n[44665];
assign t[44666] = t[44665] ^ n[44666];
assign t[44667] = t[44666] ^ n[44667];
assign t[44668] = t[44667] ^ n[44668];
assign t[44669] = t[44668] ^ n[44669];
assign t[44670] = t[44669] ^ n[44670];
assign t[44671] = t[44670] ^ n[44671];
assign t[44672] = t[44671] ^ n[44672];
assign t[44673] = t[44672] ^ n[44673];
assign t[44674] = t[44673] ^ n[44674];
assign t[44675] = t[44674] ^ n[44675];
assign t[44676] = t[44675] ^ n[44676];
assign t[44677] = t[44676] ^ n[44677];
assign t[44678] = t[44677] ^ n[44678];
assign t[44679] = t[44678] ^ n[44679];
assign t[44680] = t[44679] ^ n[44680];
assign t[44681] = t[44680] ^ n[44681];
assign t[44682] = t[44681] ^ n[44682];
assign t[44683] = t[44682] ^ n[44683];
assign t[44684] = t[44683] ^ n[44684];
assign t[44685] = t[44684] ^ n[44685];
assign t[44686] = t[44685] ^ n[44686];
assign t[44687] = t[44686] ^ n[44687];
assign t[44688] = t[44687] ^ n[44688];
assign t[44689] = t[44688] ^ n[44689];
assign t[44690] = t[44689] ^ n[44690];
assign t[44691] = t[44690] ^ n[44691];
assign t[44692] = t[44691] ^ n[44692];
assign t[44693] = t[44692] ^ n[44693];
assign t[44694] = t[44693] ^ n[44694];
assign t[44695] = t[44694] ^ n[44695];
assign t[44696] = t[44695] ^ n[44696];
assign t[44697] = t[44696] ^ n[44697];
assign t[44698] = t[44697] ^ n[44698];
assign t[44699] = t[44698] ^ n[44699];
assign t[44700] = t[44699] ^ n[44700];
assign t[44701] = t[44700] ^ n[44701];
assign t[44702] = t[44701] ^ n[44702];
assign t[44703] = t[44702] ^ n[44703];
assign t[44704] = t[44703] ^ n[44704];
assign t[44705] = t[44704] ^ n[44705];
assign t[44706] = t[44705] ^ n[44706];
assign t[44707] = t[44706] ^ n[44707];
assign t[44708] = t[44707] ^ n[44708];
assign t[44709] = t[44708] ^ n[44709];
assign t[44710] = t[44709] ^ n[44710];
assign t[44711] = t[44710] ^ n[44711];
assign t[44712] = t[44711] ^ n[44712];
assign t[44713] = t[44712] ^ n[44713];
assign t[44714] = t[44713] ^ n[44714];
assign t[44715] = t[44714] ^ n[44715];
assign t[44716] = t[44715] ^ n[44716];
assign t[44717] = t[44716] ^ n[44717];
assign t[44718] = t[44717] ^ n[44718];
assign t[44719] = t[44718] ^ n[44719];
assign t[44720] = t[44719] ^ n[44720];
assign t[44721] = t[44720] ^ n[44721];
assign t[44722] = t[44721] ^ n[44722];
assign t[44723] = t[44722] ^ n[44723];
assign t[44724] = t[44723] ^ n[44724];
assign t[44725] = t[44724] ^ n[44725];
assign t[44726] = t[44725] ^ n[44726];
assign t[44727] = t[44726] ^ n[44727];
assign t[44728] = t[44727] ^ n[44728];
assign t[44729] = t[44728] ^ n[44729];
assign t[44730] = t[44729] ^ n[44730];
assign t[44731] = t[44730] ^ n[44731];
assign t[44732] = t[44731] ^ n[44732];
assign t[44733] = t[44732] ^ n[44733];
assign t[44734] = t[44733] ^ n[44734];
assign t[44735] = t[44734] ^ n[44735];
assign t[44736] = t[44735] ^ n[44736];
assign t[44737] = t[44736] ^ n[44737];
assign t[44738] = t[44737] ^ n[44738];
assign t[44739] = t[44738] ^ n[44739];
assign t[44740] = t[44739] ^ n[44740];
assign t[44741] = t[44740] ^ n[44741];
assign t[44742] = t[44741] ^ n[44742];
assign t[44743] = t[44742] ^ n[44743];
assign t[44744] = t[44743] ^ n[44744];
assign t[44745] = t[44744] ^ n[44745];
assign t[44746] = t[44745] ^ n[44746];
assign t[44747] = t[44746] ^ n[44747];
assign t[44748] = t[44747] ^ n[44748];
assign t[44749] = t[44748] ^ n[44749];
assign t[44750] = t[44749] ^ n[44750];
assign t[44751] = t[44750] ^ n[44751];
assign t[44752] = t[44751] ^ n[44752];
assign t[44753] = t[44752] ^ n[44753];
assign t[44754] = t[44753] ^ n[44754];
assign t[44755] = t[44754] ^ n[44755];
assign t[44756] = t[44755] ^ n[44756];
assign t[44757] = t[44756] ^ n[44757];
assign t[44758] = t[44757] ^ n[44758];
assign t[44759] = t[44758] ^ n[44759];
assign t[44760] = t[44759] ^ n[44760];
assign t[44761] = t[44760] ^ n[44761];
assign t[44762] = t[44761] ^ n[44762];
assign t[44763] = t[44762] ^ n[44763];
assign t[44764] = t[44763] ^ n[44764];
assign t[44765] = t[44764] ^ n[44765];
assign t[44766] = t[44765] ^ n[44766];
assign t[44767] = t[44766] ^ n[44767];
assign t[44768] = t[44767] ^ n[44768];
assign t[44769] = t[44768] ^ n[44769];
assign t[44770] = t[44769] ^ n[44770];
assign t[44771] = t[44770] ^ n[44771];
assign t[44772] = t[44771] ^ n[44772];
assign t[44773] = t[44772] ^ n[44773];
assign t[44774] = t[44773] ^ n[44774];
assign t[44775] = t[44774] ^ n[44775];
assign t[44776] = t[44775] ^ n[44776];
assign t[44777] = t[44776] ^ n[44777];
assign t[44778] = t[44777] ^ n[44778];
assign t[44779] = t[44778] ^ n[44779];
assign t[44780] = t[44779] ^ n[44780];
assign t[44781] = t[44780] ^ n[44781];
assign t[44782] = t[44781] ^ n[44782];
assign t[44783] = t[44782] ^ n[44783];
assign t[44784] = t[44783] ^ n[44784];
assign t[44785] = t[44784] ^ n[44785];
assign t[44786] = t[44785] ^ n[44786];
assign t[44787] = t[44786] ^ n[44787];
assign t[44788] = t[44787] ^ n[44788];
assign t[44789] = t[44788] ^ n[44789];
assign t[44790] = t[44789] ^ n[44790];
assign t[44791] = t[44790] ^ n[44791];
assign t[44792] = t[44791] ^ n[44792];
assign t[44793] = t[44792] ^ n[44793];
assign t[44794] = t[44793] ^ n[44794];
assign t[44795] = t[44794] ^ n[44795];
assign t[44796] = t[44795] ^ n[44796];
assign t[44797] = t[44796] ^ n[44797];
assign t[44798] = t[44797] ^ n[44798];
assign t[44799] = t[44798] ^ n[44799];
assign t[44800] = t[44799] ^ n[44800];
assign t[44801] = t[44800] ^ n[44801];
assign t[44802] = t[44801] ^ n[44802];
assign t[44803] = t[44802] ^ n[44803];
assign t[44804] = t[44803] ^ n[44804];
assign t[44805] = t[44804] ^ n[44805];
assign t[44806] = t[44805] ^ n[44806];
assign t[44807] = t[44806] ^ n[44807];
assign t[44808] = t[44807] ^ n[44808];
assign t[44809] = t[44808] ^ n[44809];
assign t[44810] = t[44809] ^ n[44810];
assign t[44811] = t[44810] ^ n[44811];
assign t[44812] = t[44811] ^ n[44812];
assign t[44813] = t[44812] ^ n[44813];
assign t[44814] = t[44813] ^ n[44814];
assign t[44815] = t[44814] ^ n[44815];
assign t[44816] = t[44815] ^ n[44816];
assign t[44817] = t[44816] ^ n[44817];
assign t[44818] = t[44817] ^ n[44818];
assign t[44819] = t[44818] ^ n[44819];
assign t[44820] = t[44819] ^ n[44820];
assign t[44821] = t[44820] ^ n[44821];
assign t[44822] = t[44821] ^ n[44822];
assign t[44823] = t[44822] ^ n[44823];
assign t[44824] = t[44823] ^ n[44824];
assign t[44825] = t[44824] ^ n[44825];
assign t[44826] = t[44825] ^ n[44826];
assign t[44827] = t[44826] ^ n[44827];
assign t[44828] = t[44827] ^ n[44828];
assign t[44829] = t[44828] ^ n[44829];
assign t[44830] = t[44829] ^ n[44830];
assign t[44831] = t[44830] ^ n[44831];
assign t[44832] = t[44831] ^ n[44832];
assign t[44833] = t[44832] ^ n[44833];
assign t[44834] = t[44833] ^ n[44834];
assign t[44835] = t[44834] ^ n[44835];
assign t[44836] = t[44835] ^ n[44836];
assign t[44837] = t[44836] ^ n[44837];
assign t[44838] = t[44837] ^ n[44838];
assign t[44839] = t[44838] ^ n[44839];
assign t[44840] = t[44839] ^ n[44840];
assign t[44841] = t[44840] ^ n[44841];
assign t[44842] = t[44841] ^ n[44842];
assign t[44843] = t[44842] ^ n[44843];
assign t[44844] = t[44843] ^ n[44844];
assign t[44845] = t[44844] ^ n[44845];
assign t[44846] = t[44845] ^ n[44846];
assign t[44847] = t[44846] ^ n[44847];
assign t[44848] = t[44847] ^ n[44848];
assign t[44849] = t[44848] ^ n[44849];
assign t[44850] = t[44849] ^ n[44850];
assign t[44851] = t[44850] ^ n[44851];
assign t[44852] = t[44851] ^ n[44852];
assign t[44853] = t[44852] ^ n[44853];
assign t[44854] = t[44853] ^ n[44854];
assign t[44855] = t[44854] ^ n[44855];
assign t[44856] = t[44855] ^ n[44856];
assign t[44857] = t[44856] ^ n[44857];
assign t[44858] = t[44857] ^ n[44858];
assign t[44859] = t[44858] ^ n[44859];
assign t[44860] = t[44859] ^ n[44860];
assign t[44861] = t[44860] ^ n[44861];
assign t[44862] = t[44861] ^ n[44862];
assign t[44863] = t[44862] ^ n[44863];
assign t[44864] = t[44863] ^ n[44864];
assign t[44865] = t[44864] ^ n[44865];
assign t[44866] = t[44865] ^ n[44866];
assign t[44867] = t[44866] ^ n[44867];
assign t[44868] = t[44867] ^ n[44868];
assign t[44869] = t[44868] ^ n[44869];
assign t[44870] = t[44869] ^ n[44870];
assign t[44871] = t[44870] ^ n[44871];
assign t[44872] = t[44871] ^ n[44872];
assign t[44873] = t[44872] ^ n[44873];
assign t[44874] = t[44873] ^ n[44874];
assign t[44875] = t[44874] ^ n[44875];
assign t[44876] = t[44875] ^ n[44876];
assign t[44877] = t[44876] ^ n[44877];
assign t[44878] = t[44877] ^ n[44878];
assign t[44879] = t[44878] ^ n[44879];
assign t[44880] = t[44879] ^ n[44880];
assign t[44881] = t[44880] ^ n[44881];
assign t[44882] = t[44881] ^ n[44882];
assign t[44883] = t[44882] ^ n[44883];
assign t[44884] = t[44883] ^ n[44884];
assign t[44885] = t[44884] ^ n[44885];
assign t[44886] = t[44885] ^ n[44886];
assign t[44887] = t[44886] ^ n[44887];
assign t[44888] = t[44887] ^ n[44888];
assign t[44889] = t[44888] ^ n[44889];
assign t[44890] = t[44889] ^ n[44890];
assign t[44891] = t[44890] ^ n[44891];
assign t[44892] = t[44891] ^ n[44892];
assign t[44893] = t[44892] ^ n[44893];
assign t[44894] = t[44893] ^ n[44894];
assign t[44895] = t[44894] ^ n[44895];
assign t[44896] = t[44895] ^ n[44896];
assign t[44897] = t[44896] ^ n[44897];
assign t[44898] = t[44897] ^ n[44898];
assign t[44899] = t[44898] ^ n[44899];
assign t[44900] = t[44899] ^ n[44900];
assign t[44901] = t[44900] ^ n[44901];
assign t[44902] = t[44901] ^ n[44902];
assign t[44903] = t[44902] ^ n[44903];
assign t[44904] = t[44903] ^ n[44904];
assign t[44905] = t[44904] ^ n[44905];
assign t[44906] = t[44905] ^ n[44906];
assign t[44907] = t[44906] ^ n[44907];
assign t[44908] = t[44907] ^ n[44908];
assign t[44909] = t[44908] ^ n[44909];
assign t[44910] = t[44909] ^ n[44910];
assign t[44911] = t[44910] ^ n[44911];
assign t[44912] = t[44911] ^ n[44912];
assign t[44913] = t[44912] ^ n[44913];
assign t[44914] = t[44913] ^ n[44914];
assign t[44915] = t[44914] ^ n[44915];
assign t[44916] = t[44915] ^ n[44916];
assign t[44917] = t[44916] ^ n[44917];
assign t[44918] = t[44917] ^ n[44918];
assign t[44919] = t[44918] ^ n[44919];
assign t[44920] = t[44919] ^ n[44920];
assign t[44921] = t[44920] ^ n[44921];
assign t[44922] = t[44921] ^ n[44922];
assign t[44923] = t[44922] ^ n[44923];
assign t[44924] = t[44923] ^ n[44924];
assign t[44925] = t[44924] ^ n[44925];
assign t[44926] = t[44925] ^ n[44926];
assign t[44927] = t[44926] ^ n[44927];
assign t[44928] = t[44927] ^ n[44928];
assign t[44929] = t[44928] ^ n[44929];
assign t[44930] = t[44929] ^ n[44930];
assign t[44931] = t[44930] ^ n[44931];
assign t[44932] = t[44931] ^ n[44932];
assign t[44933] = t[44932] ^ n[44933];
assign t[44934] = t[44933] ^ n[44934];
assign t[44935] = t[44934] ^ n[44935];
assign t[44936] = t[44935] ^ n[44936];
assign t[44937] = t[44936] ^ n[44937];
assign t[44938] = t[44937] ^ n[44938];
assign t[44939] = t[44938] ^ n[44939];
assign t[44940] = t[44939] ^ n[44940];
assign t[44941] = t[44940] ^ n[44941];
assign t[44942] = t[44941] ^ n[44942];
assign t[44943] = t[44942] ^ n[44943];
assign t[44944] = t[44943] ^ n[44944];
assign t[44945] = t[44944] ^ n[44945];
assign t[44946] = t[44945] ^ n[44946];
assign t[44947] = t[44946] ^ n[44947];
assign t[44948] = t[44947] ^ n[44948];
assign t[44949] = t[44948] ^ n[44949];
assign t[44950] = t[44949] ^ n[44950];
assign t[44951] = t[44950] ^ n[44951];
assign t[44952] = t[44951] ^ n[44952];
assign t[44953] = t[44952] ^ n[44953];
assign t[44954] = t[44953] ^ n[44954];
assign t[44955] = t[44954] ^ n[44955];
assign t[44956] = t[44955] ^ n[44956];
assign t[44957] = t[44956] ^ n[44957];
assign t[44958] = t[44957] ^ n[44958];
assign t[44959] = t[44958] ^ n[44959];
assign t[44960] = t[44959] ^ n[44960];
assign t[44961] = t[44960] ^ n[44961];
assign t[44962] = t[44961] ^ n[44962];
assign t[44963] = t[44962] ^ n[44963];
assign t[44964] = t[44963] ^ n[44964];
assign t[44965] = t[44964] ^ n[44965];
assign t[44966] = t[44965] ^ n[44966];
assign t[44967] = t[44966] ^ n[44967];
assign t[44968] = t[44967] ^ n[44968];
assign t[44969] = t[44968] ^ n[44969];
assign t[44970] = t[44969] ^ n[44970];
assign t[44971] = t[44970] ^ n[44971];
assign t[44972] = t[44971] ^ n[44972];
assign t[44973] = t[44972] ^ n[44973];
assign t[44974] = t[44973] ^ n[44974];
assign t[44975] = t[44974] ^ n[44975];
assign t[44976] = t[44975] ^ n[44976];
assign t[44977] = t[44976] ^ n[44977];
assign t[44978] = t[44977] ^ n[44978];
assign t[44979] = t[44978] ^ n[44979];
assign t[44980] = t[44979] ^ n[44980];
assign t[44981] = t[44980] ^ n[44981];
assign t[44982] = t[44981] ^ n[44982];
assign t[44983] = t[44982] ^ n[44983];
assign t[44984] = t[44983] ^ n[44984];
assign t[44985] = t[44984] ^ n[44985];
assign t[44986] = t[44985] ^ n[44986];
assign t[44987] = t[44986] ^ n[44987];
assign t[44988] = t[44987] ^ n[44988];
assign t[44989] = t[44988] ^ n[44989];
assign t[44990] = t[44989] ^ n[44990];
assign t[44991] = t[44990] ^ n[44991];
assign t[44992] = t[44991] ^ n[44992];
assign t[44993] = t[44992] ^ n[44993];
assign t[44994] = t[44993] ^ n[44994];
assign t[44995] = t[44994] ^ n[44995];
assign t[44996] = t[44995] ^ n[44996];
assign t[44997] = t[44996] ^ n[44997];
assign t[44998] = t[44997] ^ n[44998];
assign t[44999] = t[44998] ^ n[44999];
assign t[45000] = t[44999] ^ n[45000];
assign t[45001] = t[45000] ^ n[45001];
assign t[45002] = t[45001] ^ n[45002];
assign t[45003] = t[45002] ^ n[45003];
assign t[45004] = t[45003] ^ n[45004];
assign t[45005] = t[45004] ^ n[45005];
assign t[45006] = t[45005] ^ n[45006];
assign t[45007] = t[45006] ^ n[45007];
assign t[45008] = t[45007] ^ n[45008];
assign t[45009] = t[45008] ^ n[45009];
assign t[45010] = t[45009] ^ n[45010];
assign t[45011] = t[45010] ^ n[45011];
assign t[45012] = t[45011] ^ n[45012];
assign t[45013] = t[45012] ^ n[45013];
assign t[45014] = t[45013] ^ n[45014];
assign t[45015] = t[45014] ^ n[45015];
assign t[45016] = t[45015] ^ n[45016];
assign t[45017] = t[45016] ^ n[45017];
assign t[45018] = t[45017] ^ n[45018];
assign t[45019] = t[45018] ^ n[45019];
assign t[45020] = t[45019] ^ n[45020];
assign t[45021] = t[45020] ^ n[45021];
assign t[45022] = t[45021] ^ n[45022];
assign t[45023] = t[45022] ^ n[45023];
assign t[45024] = t[45023] ^ n[45024];
assign t[45025] = t[45024] ^ n[45025];
assign t[45026] = t[45025] ^ n[45026];
assign t[45027] = t[45026] ^ n[45027];
assign t[45028] = t[45027] ^ n[45028];
assign t[45029] = t[45028] ^ n[45029];
assign t[45030] = t[45029] ^ n[45030];
assign t[45031] = t[45030] ^ n[45031];
assign t[45032] = t[45031] ^ n[45032];
assign t[45033] = t[45032] ^ n[45033];
assign t[45034] = t[45033] ^ n[45034];
assign t[45035] = t[45034] ^ n[45035];
assign t[45036] = t[45035] ^ n[45036];
assign t[45037] = t[45036] ^ n[45037];
assign t[45038] = t[45037] ^ n[45038];
assign t[45039] = t[45038] ^ n[45039];
assign t[45040] = t[45039] ^ n[45040];
assign t[45041] = t[45040] ^ n[45041];
assign t[45042] = t[45041] ^ n[45042];
assign t[45043] = t[45042] ^ n[45043];
assign t[45044] = t[45043] ^ n[45044];
assign t[45045] = t[45044] ^ n[45045];
assign t[45046] = t[45045] ^ n[45046];
assign t[45047] = t[45046] ^ n[45047];
assign t[45048] = t[45047] ^ n[45048];
assign t[45049] = t[45048] ^ n[45049];
assign t[45050] = t[45049] ^ n[45050];
assign t[45051] = t[45050] ^ n[45051];
assign t[45052] = t[45051] ^ n[45052];
assign t[45053] = t[45052] ^ n[45053];
assign t[45054] = t[45053] ^ n[45054];
assign t[45055] = t[45054] ^ n[45055];
assign t[45056] = t[45055] ^ n[45056];
assign t[45057] = t[45056] ^ n[45057];
assign t[45058] = t[45057] ^ n[45058];
assign t[45059] = t[45058] ^ n[45059];
assign t[45060] = t[45059] ^ n[45060];
assign t[45061] = t[45060] ^ n[45061];
assign t[45062] = t[45061] ^ n[45062];
assign t[45063] = t[45062] ^ n[45063];
assign t[45064] = t[45063] ^ n[45064];
assign t[45065] = t[45064] ^ n[45065];
assign t[45066] = t[45065] ^ n[45066];
assign t[45067] = t[45066] ^ n[45067];
assign t[45068] = t[45067] ^ n[45068];
assign t[45069] = t[45068] ^ n[45069];
assign t[45070] = t[45069] ^ n[45070];
assign t[45071] = t[45070] ^ n[45071];
assign t[45072] = t[45071] ^ n[45072];
assign t[45073] = t[45072] ^ n[45073];
assign t[45074] = t[45073] ^ n[45074];
assign t[45075] = t[45074] ^ n[45075];
assign t[45076] = t[45075] ^ n[45076];
assign t[45077] = t[45076] ^ n[45077];
assign t[45078] = t[45077] ^ n[45078];
assign t[45079] = t[45078] ^ n[45079];
assign t[45080] = t[45079] ^ n[45080];
assign t[45081] = t[45080] ^ n[45081];
assign t[45082] = t[45081] ^ n[45082];
assign t[45083] = t[45082] ^ n[45083];
assign t[45084] = t[45083] ^ n[45084];
assign t[45085] = t[45084] ^ n[45085];
assign t[45086] = t[45085] ^ n[45086];
assign t[45087] = t[45086] ^ n[45087];
assign t[45088] = t[45087] ^ n[45088];
assign t[45089] = t[45088] ^ n[45089];
assign t[45090] = t[45089] ^ n[45090];
assign t[45091] = t[45090] ^ n[45091];
assign t[45092] = t[45091] ^ n[45092];
assign t[45093] = t[45092] ^ n[45093];
assign t[45094] = t[45093] ^ n[45094];
assign t[45095] = t[45094] ^ n[45095];
assign t[45096] = t[45095] ^ n[45096];
assign t[45097] = t[45096] ^ n[45097];
assign t[45098] = t[45097] ^ n[45098];
assign t[45099] = t[45098] ^ n[45099];
assign t[45100] = t[45099] ^ n[45100];
assign t[45101] = t[45100] ^ n[45101];
assign t[45102] = t[45101] ^ n[45102];
assign t[45103] = t[45102] ^ n[45103];
assign t[45104] = t[45103] ^ n[45104];
assign t[45105] = t[45104] ^ n[45105];
assign t[45106] = t[45105] ^ n[45106];
assign t[45107] = t[45106] ^ n[45107];
assign t[45108] = t[45107] ^ n[45108];
assign t[45109] = t[45108] ^ n[45109];
assign t[45110] = t[45109] ^ n[45110];
assign t[45111] = t[45110] ^ n[45111];
assign t[45112] = t[45111] ^ n[45112];
assign t[45113] = t[45112] ^ n[45113];
assign t[45114] = t[45113] ^ n[45114];
assign t[45115] = t[45114] ^ n[45115];
assign t[45116] = t[45115] ^ n[45116];
assign t[45117] = t[45116] ^ n[45117];
assign t[45118] = t[45117] ^ n[45118];
assign t[45119] = t[45118] ^ n[45119];
assign t[45120] = t[45119] ^ n[45120];
assign t[45121] = t[45120] ^ n[45121];
assign t[45122] = t[45121] ^ n[45122];
assign t[45123] = t[45122] ^ n[45123];
assign t[45124] = t[45123] ^ n[45124];
assign t[45125] = t[45124] ^ n[45125];
assign t[45126] = t[45125] ^ n[45126];
assign t[45127] = t[45126] ^ n[45127];
assign t[45128] = t[45127] ^ n[45128];
assign t[45129] = t[45128] ^ n[45129];
assign t[45130] = t[45129] ^ n[45130];
assign t[45131] = t[45130] ^ n[45131];
assign t[45132] = t[45131] ^ n[45132];
assign t[45133] = t[45132] ^ n[45133];
assign t[45134] = t[45133] ^ n[45134];
assign t[45135] = t[45134] ^ n[45135];
assign t[45136] = t[45135] ^ n[45136];
assign t[45137] = t[45136] ^ n[45137];
assign t[45138] = t[45137] ^ n[45138];
assign t[45139] = t[45138] ^ n[45139];
assign t[45140] = t[45139] ^ n[45140];
assign t[45141] = t[45140] ^ n[45141];
assign t[45142] = t[45141] ^ n[45142];
assign t[45143] = t[45142] ^ n[45143];
assign t[45144] = t[45143] ^ n[45144];
assign t[45145] = t[45144] ^ n[45145];
assign t[45146] = t[45145] ^ n[45146];
assign t[45147] = t[45146] ^ n[45147];
assign t[45148] = t[45147] ^ n[45148];
assign t[45149] = t[45148] ^ n[45149];
assign t[45150] = t[45149] ^ n[45150];
assign t[45151] = t[45150] ^ n[45151];
assign t[45152] = t[45151] ^ n[45152];
assign t[45153] = t[45152] ^ n[45153];
assign t[45154] = t[45153] ^ n[45154];
assign t[45155] = t[45154] ^ n[45155];
assign t[45156] = t[45155] ^ n[45156];
assign t[45157] = t[45156] ^ n[45157];
assign t[45158] = t[45157] ^ n[45158];
assign t[45159] = t[45158] ^ n[45159];
assign t[45160] = t[45159] ^ n[45160];
assign t[45161] = t[45160] ^ n[45161];
assign t[45162] = t[45161] ^ n[45162];
assign t[45163] = t[45162] ^ n[45163];
assign t[45164] = t[45163] ^ n[45164];
assign t[45165] = t[45164] ^ n[45165];
assign t[45166] = t[45165] ^ n[45166];
assign t[45167] = t[45166] ^ n[45167];
assign t[45168] = t[45167] ^ n[45168];
assign t[45169] = t[45168] ^ n[45169];
assign t[45170] = t[45169] ^ n[45170];
assign t[45171] = t[45170] ^ n[45171];
assign t[45172] = t[45171] ^ n[45172];
assign t[45173] = t[45172] ^ n[45173];
assign t[45174] = t[45173] ^ n[45174];
assign t[45175] = t[45174] ^ n[45175];
assign t[45176] = t[45175] ^ n[45176];
assign t[45177] = t[45176] ^ n[45177];
assign t[45178] = t[45177] ^ n[45178];
assign t[45179] = t[45178] ^ n[45179];
assign t[45180] = t[45179] ^ n[45180];
assign t[45181] = t[45180] ^ n[45181];
assign t[45182] = t[45181] ^ n[45182];
assign t[45183] = t[45182] ^ n[45183];
assign t[45184] = t[45183] ^ n[45184];
assign t[45185] = t[45184] ^ n[45185];
assign t[45186] = t[45185] ^ n[45186];
assign t[45187] = t[45186] ^ n[45187];
assign t[45188] = t[45187] ^ n[45188];
assign t[45189] = t[45188] ^ n[45189];
assign t[45190] = t[45189] ^ n[45190];
assign t[45191] = t[45190] ^ n[45191];
assign t[45192] = t[45191] ^ n[45192];
assign t[45193] = t[45192] ^ n[45193];
assign t[45194] = t[45193] ^ n[45194];
assign t[45195] = t[45194] ^ n[45195];
assign t[45196] = t[45195] ^ n[45196];
assign t[45197] = t[45196] ^ n[45197];
assign t[45198] = t[45197] ^ n[45198];
assign t[45199] = t[45198] ^ n[45199];
assign t[45200] = t[45199] ^ n[45200];
assign t[45201] = t[45200] ^ n[45201];
assign t[45202] = t[45201] ^ n[45202];
assign t[45203] = t[45202] ^ n[45203];
assign t[45204] = t[45203] ^ n[45204];
assign t[45205] = t[45204] ^ n[45205];
assign t[45206] = t[45205] ^ n[45206];
assign t[45207] = t[45206] ^ n[45207];
assign t[45208] = t[45207] ^ n[45208];
assign t[45209] = t[45208] ^ n[45209];
assign t[45210] = t[45209] ^ n[45210];
assign t[45211] = t[45210] ^ n[45211];
assign t[45212] = t[45211] ^ n[45212];
assign t[45213] = t[45212] ^ n[45213];
assign t[45214] = t[45213] ^ n[45214];
assign t[45215] = t[45214] ^ n[45215];
assign t[45216] = t[45215] ^ n[45216];
assign t[45217] = t[45216] ^ n[45217];
assign t[45218] = t[45217] ^ n[45218];
assign t[45219] = t[45218] ^ n[45219];
assign t[45220] = t[45219] ^ n[45220];
assign t[45221] = t[45220] ^ n[45221];
assign t[45222] = t[45221] ^ n[45222];
assign t[45223] = t[45222] ^ n[45223];
assign t[45224] = t[45223] ^ n[45224];
assign t[45225] = t[45224] ^ n[45225];
assign t[45226] = t[45225] ^ n[45226];
assign t[45227] = t[45226] ^ n[45227];
assign t[45228] = t[45227] ^ n[45228];
assign t[45229] = t[45228] ^ n[45229];
assign t[45230] = t[45229] ^ n[45230];
assign t[45231] = t[45230] ^ n[45231];
assign t[45232] = t[45231] ^ n[45232];
assign t[45233] = t[45232] ^ n[45233];
assign t[45234] = t[45233] ^ n[45234];
assign t[45235] = t[45234] ^ n[45235];
assign t[45236] = t[45235] ^ n[45236];
assign t[45237] = t[45236] ^ n[45237];
assign t[45238] = t[45237] ^ n[45238];
assign t[45239] = t[45238] ^ n[45239];
assign t[45240] = t[45239] ^ n[45240];
assign t[45241] = t[45240] ^ n[45241];
assign t[45242] = t[45241] ^ n[45242];
assign t[45243] = t[45242] ^ n[45243];
assign t[45244] = t[45243] ^ n[45244];
assign t[45245] = t[45244] ^ n[45245];
assign t[45246] = t[45245] ^ n[45246];
assign t[45247] = t[45246] ^ n[45247];
assign t[45248] = t[45247] ^ n[45248];
assign t[45249] = t[45248] ^ n[45249];
assign t[45250] = t[45249] ^ n[45250];
assign t[45251] = t[45250] ^ n[45251];
assign t[45252] = t[45251] ^ n[45252];
assign t[45253] = t[45252] ^ n[45253];
assign t[45254] = t[45253] ^ n[45254];
assign t[45255] = t[45254] ^ n[45255];
assign t[45256] = t[45255] ^ n[45256];
assign t[45257] = t[45256] ^ n[45257];
assign t[45258] = t[45257] ^ n[45258];
assign t[45259] = t[45258] ^ n[45259];
assign t[45260] = t[45259] ^ n[45260];
assign t[45261] = t[45260] ^ n[45261];
assign t[45262] = t[45261] ^ n[45262];
assign t[45263] = t[45262] ^ n[45263];
assign t[45264] = t[45263] ^ n[45264];
assign t[45265] = t[45264] ^ n[45265];
assign t[45266] = t[45265] ^ n[45266];
assign t[45267] = t[45266] ^ n[45267];
assign t[45268] = t[45267] ^ n[45268];
assign t[45269] = t[45268] ^ n[45269];
assign t[45270] = t[45269] ^ n[45270];
assign t[45271] = t[45270] ^ n[45271];
assign t[45272] = t[45271] ^ n[45272];
assign t[45273] = t[45272] ^ n[45273];
assign t[45274] = t[45273] ^ n[45274];
assign t[45275] = t[45274] ^ n[45275];
assign t[45276] = t[45275] ^ n[45276];
assign t[45277] = t[45276] ^ n[45277];
assign t[45278] = t[45277] ^ n[45278];
assign t[45279] = t[45278] ^ n[45279];
assign t[45280] = t[45279] ^ n[45280];
assign t[45281] = t[45280] ^ n[45281];
assign t[45282] = t[45281] ^ n[45282];
assign t[45283] = t[45282] ^ n[45283];
assign t[45284] = t[45283] ^ n[45284];
assign t[45285] = t[45284] ^ n[45285];
assign t[45286] = t[45285] ^ n[45286];
assign t[45287] = t[45286] ^ n[45287];
assign t[45288] = t[45287] ^ n[45288];
assign t[45289] = t[45288] ^ n[45289];
assign t[45290] = t[45289] ^ n[45290];
assign t[45291] = t[45290] ^ n[45291];
assign t[45292] = t[45291] ^ n[45292];
assign t[45293] = t[45292] ^ n[45293];
assign t[45294] = t[45293] ^ n[45294];
assign t[45295] = t[45294] ^ n[45295];
assign t[45296] = t[45295] ^ n[45296];
assign t[45297] = t[45296] ^ n[45297];
assign t[45298] = t[45297] ^ n[45298];
assign t[45299] = t[45298] ^ n[45299];
assign t[45300] = t[45299] ^ n[45300];
assign t[45301] = t[45300] ^ n[45301];
assign t[45302] = t[45301] ^ n[45302];
assign t[45303] = t[45302] ^ n[45303];
assign t[45304] = t[45303] ^ n[45304];
assign t[45305] = t[45304] ^ n[45305];
assign t[45306] = t[45305] ^ n[45306];
assign t[45307] = t[45306] ^ n[45307];
assign t[45308] = t[45307] ^ n[45308];
assign t[45309] = t[45308] ^ n[45309];
assign t[45310] = t[45309] ^ n[45310];
assign t[45311] = t[45310] ^ n[45311];
assign t[45312] = t[45311] ^ n[45312];
assign t[45313] = t[45312] ^ n[45313];
assign t[45314] = t[45313] ^ n[45314];
assign t[45315] = t[45314] ^ n[45315];
assign t[45316] = t[45315] ^ n[45316];
assign t[45317] = t[45316] ^ n[45317];
assign t[45318] = t[45317] ^ n[45318];
assign t[45319] = t[45318] ^ n[45319];
assign t[45320] = t[45319] ^ n[45320];
assign t[45321] = t[45320] ^ n[45321];
assign t[45322] = t[45321] ^ n[45322];
assign t[45323] = t[45322] ^ n[45323];
assign t[45324] = t[45323] ^ n[45324];
assign t[45325] = t[45324] ^ n[45325];
assign t[45326] = t[45325] ^ n[45326];
assign t[45327] = t[45326] ^ n[45327];
assign t[45328] = t[45327] ^ n[45328];
assign t[45329] = t[45328] ^ n[45329];
assign t[45330] = t[45329] ^ n[45330];
assign t[45331] = t[45330] ^ n[45331];
assign t[45332] = t[45331] ^ n[45332];
assign t[45333] = t[45332] ^ n[45333];
assign t[45334] = t[45333] ^ n[45334];
assign t[45335] = t[45334] ^ n[45335];
assign t[45336] = t[45335] ^ n[45336];
assign t[45337] = t[45336] ^ n[45337];
assign t[45338] = t[45337] ^ n[45338];
assign t[45339] = t[45338] ^ n[45339];
assign t[45340] = t[45339] ^ n[45340];
assign t[45341] = t[45340] ^ n[45341];
assign t[45342] = t[45341] ^ n[45342];
assign t[45343] = t[45342] ^ n[45343];
assign t[45344] = t[45343] ^ n[45344];
assign t[45345] = t[45344] ^ n[45345];
assign t[45346] = t[45345] ^ n[45346];
assign t[45347] = t[45346] ^ n[45347];
assign t[45348] = t[45347] ^ n[45348];
assign t[45349] = t[45348] ^ n[45349];
assign t[45350] = t[45349] ^ n[45350];
assign t[45351] = t[45350] ^ n[45351];
assign t[45352] = t[45351] ^ n[45352];
assign t[45353] = t[45352] ^ n[45353];
assign t[45354] = t[45353] ^ n[45354];
assign t[45355] = t[45354] ^ n[45355];
assign t[45356] = t[45355] ^ n[45356];
assign t[45357] = t[45356] ^ n[45357];
assign t[45358] = t[45357] ^ n[45358];
assign t[45359] = t[45358] ^ n[45359];
assign t[45360] = t[45359] ^ n[45360];
assign t[45361] = t[45360] ^ n[45361];
assign t[45362] = t[45361] ^ n[45362];
assign t[45363] = t[45362] ^ n[45363];
assign t[45364] = t[45363] ^ n[45364];
assign t[45365] = t[45364] ^ n[45365];
assign t[45366] = t[45365] ^ n[45366];
assign t[45367] = t[45366] ^ n[45367];
assign t[45368] = t[45367] ^ n[45368];
assign t[45369] = t[45368] ^ n[45369];
assign t[45370] = t[45369] ^ n[45370];
assign t[45371] = t[45370] ^ n[45371];
assign t[45372] = t[45371] ^ n[45372];
assign t[45373] = t[45372] ^ n[45373];
assign t[45374] = t[45373] ^ n[45374];
assign t[45375] = t[45374] ^ n[45375];
assign t[45376] = t[45375] ^ n[45376];
assign t[45377] = t[45376] ^ n[45377];
assign t[45378] = t[45377] ^ n[45378];
assign t[45379] = t[45378] ^ n[45379];
assign t[45380] = t[45379] ^ n[45380];
assign t[45381] = t[45380] ^ n[45381];
assign t[45382] = t[45381] ^ n[45382];
assign t[45383] = t[45382] ^ n[45383];
assign t[45384] = t[45383] ^ n[45384];
assign t[45385] = t[45384] ^ n[45385];
assign t[45386] = t[45385] ^ n[45386];
assign t[45387] = t[45386] ^ n[45387];
assign t[45388] = t[45387] ^ n[45388];
assign t[45389] = t[45388] ^ n[45389];
assign t[45390] = t[45389] ^ n[45390];
assign t[45391] = t[45390] ^ n[45391];
assign t[45392] = t[45391] ^ n[45392];
assign t[45393] = t[45392] ^ n[45393];
assign t[45394] = t[45393] ^ n[45394];
assign t[45395] = t[45394] ^ n[45395];
assign t[45396] = t[45395] ^ n[45396];
assign t[45397] = t[45396] ^ n[45397];
assign t[45398] = t[45397] ^ n[45398];
assign t[45399] = t[45398] ^ n[45399];
assign t[45400] = t[45399] ^ n[45400];
assign t[45401] = t[45400] ^ n[45401];
assign t[45402] = t[45401] ^ n[45402];
assign t[45403] = t[45402] ^ n[45403];
assign t[45404] = t[45403] ^ n[45404];
assign t[45405] = t[45404] ^ n[45405];
assign t[45406] = t[45405] ^ n[45406];
assign t[45407] = t[45406] ^ n[45407];
assign t[45408] = t[45407] ^ n[45408];
assign t[45409] = t[45408] ^ n[45409];
assign t[45410] = t[45409] ^ n[45410];
assign t[45411] = t[45410] ^ n[45411];
assign t[45412] = t[45411] ^ n[45412];
assign t[45413] = t[45412] ^ n[45413];
assign t[45414] = t[45413] ^ n[45414];
assign t[45415] = t[45414] ^ n[45415];
assign t[45416] = t[45415] ^ n[45416];
assign t[45417] = t[45416] ^ n[45417];
assign t[45418] = t[45417] ^ n[45418];
assign t[45419] = t[45418] ^ n[45419];
assign t[45420] = t[45419] ^ n[45420];
assign t[45421] = t[45420] ^ n[45421];
assign t[45422] = t[45421] ^ n[45422];
assign t[45423] = t[45422] ^ n[45423];
assign t[45424] = t[45423] ^ n[45424];
assign t[45425] = t[45424] ^ n[45425];
assign t[45426] = t[45425] ^ n[45426];
assign t[45427] = t[45426] ^ n[45427];
assign t[45428] = t[45427] ^ n[45428];
assign t[45429] = t[45428] ^ n[45429];
assign t[45430] = t[45429] ^ n[45430];
assign t[45431] = t[45430] ^ n[45431];
assign t[45432] = t[45431] ^ n[45432];
assign t[45433] = t[45432] ^ n[45433];
assign t[45434] = t[45433] ^ n[45434];
assign t[45435] = t[45434] ^ n[45435];
assign t[45436] = t[45435] ^ n[45436];
assign t[45437] = t[45436] ^ n[45437];
assign t[45438] = t[45437] ^ n[45438];
assign t[45439] = t[45438] ^ n[45439];
assign t[45440] = t[45439] ^ n[45440];
assign t[45441] = t[45440] ^ n[45441];
assign t[45442] = t[45441] ^ n[45442];
assign t[45443] = t[45442] ^ n[45443];
assign t[45444] = t[45443] ^ n[45444];
assign t[45445] = t[45444] ^ n[45445];
assign t[45446] = t[45445] ^ n[45446];
assign t[45447] = t[45446] ^ n[45447];
assign t[45448] = t[45447] ^ n[45448];
assign t[45449] = t[45448] ^ n[45449];
assign t[45450] = t[45449] ^ n[45450];
assign t[45451] = t[45450] ^ n[45451];
assign t[45452] = t[45451] ^ n[45452];
assign t[45453] = t[45452] ^ n[45453];
assign t[45454] = t[45453] ^ n[45454];
assign t[45455] = t[45454] ^ n[45455];
assign t[45456] = t[45455] ^ n[45456];
assign t[45457] = t[45456] ^ n[45457];
assign t[45458] = t[45457] ^ n[45458];
assign t[45459] = t[45458] ^ n[45459];
assign t[45460] = t[45459] ^ n[45460];
assign t[45461] = t[45460] ^ n[45461];
assign t[45462] = t[45461] ^ n[45462];
assign t[45463] = t[45462] ^ n[45463];
assign t[45464] = t[45463] ^ n[45464];
assign t[45465] = t[45464] ^ n[45465];
assign t[45466] = t[45465] ^ n[45466];
assign t[45467] = t[45466] ^ n[45467];
assign t[45468] = t[45467] ^ n[45468];
assign t[45469] = t[45468] ^ n[45469];
assign t[45470] = t[45469] ^ n[45470];
assign t[45471] = t[45470] ^ n[45471];
assign t[45472] = t[45471] ^ n[45472];
assign t[45473] = t[45472] ^ n[45473];
assign t[45474] = t[45473] ^ n[45474];
assign t[45475] = t[45474] ^ n[45475];
assign t[45476] = t[45475] ^ n[45476];
assign t[45477] = t[45476] ^ n[45477];
assign t[45478] = t[45477] ^ n[45478];
assign t[45479] = t[45478] ^ n[45479];
assign t[45480] = t[45479] ^ n[45480];
assign t[45481] = t[45480] ^ n[45481];
assign t[45482] = t[45481] ^ n[45482];
assign t[45483] = t[45482] ^ n[45483];
assign t[45484] = t[45483] ^ n[45484];
assign t[45485] = t[45484] ^ n[45485];
assign t[45486] = t[45485] ^ n[45486];
assign t[45487] = t[45486] ^ n[45487];
assign t[45488] = t[45487] ^ n[45488];
assign t[45489] = t[45488] ^ n[45489];
assign t[45490] = t[45489] ^ n[45490];
assign t[45491] = t[45490] ^ n[45491];
assign t[45492] = t[45491] ^ n[45492];
assign t[45493] = t[45492] ^ n[45493];
assign t[45494] = t[45493] ^ n[45494];
assign t[45495] = t[45494] ^ n[45495];
assign t[45496] = t[45495] ^ n[45496];
assign t[45497] = t[45496] ^ n[45497];
assign t[45498] = t[45497] ^ n[45498];
assign t[45499] = t[45498] ^ n[45499];
assign t[45500] = t[45499] ^ n[45500];
assign t[45501] = t[45500] ^ n[45501];
assign t[45502] = t[45501] ^ n[45502];
assign t[45503] = t[45502] ^ n[45503];
assign t[45504] = t[45503] ^ n[45504];
assign t[45505] = t[45504] ^ n[45505];
assign t[45506] = t[45505] ^ n[45506];
assign t[45507] = t[45506] ^ n[45507];
assign t[45508] = t[45507] ^ n[45508];
assign t[45509] = t[45508] ^ n[45509];
assign t[45510] = t[45509] ^ n[45510];
assign t[45511] = t[45510] ^ n[45511];
assign t[45512] = t[45511] ^ n[45512];
assign t[45513] = t[45512] ^ n[45513];
assign t[45514] = t[45513] ^ n[45514];
assign t[45515] = t[45514] ^ n[45515];
assign t[45516] = t[45515] ^ n[45516];
assign t[45517] = t[45516] ^ n[45517];
assign t[45518] = t[45517] ^ n[45518];
assign t[45519] = t[45518] ^ n[45519];
assign t[45520] = t[45519] ^ n[45520];
assign t[45521] = t[45520] ^ n[45521];
assign t[45522] = t[45521] ^ n[45522];
assign t[45523] = t[45522] ^ n[45523];
assign t[45524] = t[45523] ^ n[45524];
assign t[45525] = t[45524] ^ n[45525];
assign t[45526] = t[45525] ^ n[45526];
assign t[45527] = t[45526] ^ n[45527];
assign t[45528] = t[45527] ^ n[45528];
assign t[45529] = t[45528] ^ n[45529];
assign t[45530] = t[45529] ^ n[45530];
assign t[45531] = t[45530] ^ n[45531];
assign t[45532] = t[45531] ^ n[45532];
assign t[45533] = t[45532] ^ n[45533];
assign t[45534] = t[45533] ^ n[45534];
assign t[45535] = t[45534] ^ n[45535];
assign t[45536] = t[45535] ^ n[45536];
assign t[45537] = t[45536] ^ n[45537];
assign t[45538] = t[45537] ^ n[45538];
assign t[45539] = t[45538] ^ n[45539];
assign t[45540] = t[45539] ^ n[45540];
assign t[45541] = t[45540] ^ n[45541];
assign t[45542] = t[45541] ^ n[45542];
assign t[45543] = t[45542] ^ n[45543];
assign t[45544] = t[45543] ^ n[45544];
assign t[45545] = t[45544] ^ n[45545];
assign t[45546] = t[45545] ^ n[45546];
assign t[45547] = t[45546] ^ n[45547];
assign t[45548] = t[45547] ^ n[45548];
assign t[45549] = t[45548] ^ n[45549];
assign t[45550] = t[45549] ^ n[45550];
assign t[45551] = t[45550] ^ n[45551];
assign t[45552] = t[45551] ^ n[45552];
assign t[45553] = t[45552] ^ n[45553];
assign t[45554] = t[45553] ^ n[45554];
assign t[45555] = t[45554] ^ n[45555];
assign t[45556] = t[45555] ^ n[45556];
assign t[45557] = t[45556] ^ n[45557];
assign t[45558] = t[45557] ^ n[45558];
assign t[45559] = t[45558] ^ n[45559];
assign t[45560] = t[45559] ^ n[45560];
assign t[45561] = t[45560] ^ n[45561];
assign t[45562] = t[45561] ^ n[45562];
assign t[45563] = t[45562] ^ n[45563];
assign t[45564] = t[45563] ^ n[45564];
assign t[45565] = t[45564] ^ n[45565];
assign t[45566] = t[45565] ^ n[45566];
assign t[45567] = t[45566] ^ n[45567];
assign t[45568] = t[45567] ^ n[45568];
assign t[45569] = t[45568] ^ n[45569];
assign t[45570] = t[45569] ^ n[45570];
assign t[45571] = t[45570] ^ n[45571];
assign t[45572] = t[45571] ^ n[45572];
assign t[45573] = t[45572] ^ n[45573];
assign t[45574] = t[45573] ^ n[45574];
assign t[45575] = t[45574] ^ n[45575];
assign t[45576] = t[45575] ^ n[45576];
assign t[45577] = t[45576] ^ n[45577];
assign t[45578] = t[45577] ^ n[45578];
assign t[45579] = t[45578] ^ n[45579];
assign t[45580] = t[45579] ^ n[45580];
assign t[45581] = t[45580] ^ n[45581];
assign t[45582] = t[45581] ^ n[45582];
assign t[45583] = t[45582] ^ n[45583];
assign t[45584] = t[45583] ^ n[45584];
assign t[45585] = t[45584] ^ n[45585];
assign t[45586] = t[45585] ^ n[45586];
assign t[45587] = t[45586] ^ n[45587];
assign t[45588] = t[45587] ^ n[45588];
assign t[45589] = t[45588] ^ n[45589];
assign t[45590] = t[45589] ^ n[45590];
assign t[45591] = t[45590] ^ n[45591];
assign t[45592] = t[45591] ^ n[45592];
assign t[45593] = t[45592] ^ n[45593];
assign t[45594] = t[45593] ^ n[45594];
assign t[45595] = t[45594] ^ n[45595];
assign t[45596] = t[45595] ^ n[45596];
assign t[45597] = t[45596] ^ n[45597];
assign t[45598] = t[45597] ^ n[45598];
assign t[45599] = t[45598] ^ n[45599];
assign t[45600] = t[45599] ^ n[45600];
assign t[45601] = t[45600] ^ n[45601];
assign t[45602] = t[45601] ^ n[45602];
assign t[45603] = t[45602] ^ n[45603];
assign t[45604] = t[45603] ^ n[45604];
assign t[45605] = t[45604] ^ n[45605];
assign t[45606] = t[45605] ^ n[45606];
assign t[45607] = t[45606] ^ n[45607];
assign t[45608] = t[45607] ^ n[45608];
assign t[45609] = t[45608] ^ n[45609];
assign t[45610] = t[45609] ^ n[45610];
assign t[45611] = t[45610] ^ n[45611];
assign t[45612] = t[45611] ^ n[45612];
assign t[45613] = t[45612] ^ n[45613];
assign t[45614] = t[45613] ^ n[45614];
assign t[45615] = t[45614] ^ n[45615];
assign t[45616] = t[45615] ^ n[45616];
assign t[45617] = t[45616] ^ n[45617];
assign t[45618] = t[45617] ^ n[45618];
assign t[45619] = t[45618] ^ n[45619];
assign t[45620] = t[45619] ^ n[45620];
assign t[45621] = t[45620] ^ n[45621];
assign t[45622] = t[45621] ^ n[45622];
assign t[45623] = t[45622] ^ n[45623];
assign t[45624] = t[45623] ^ n[45624];
assign t[45625] = t[45624] ^ n[45625];
assign t[45626] = t[45625] ^ n[45626];
assign t[45627] = t[45626] ^ n[45627];
assign t[45628] = t[45627] ^ n[45628];
assign t[45629] = t[45628] ^ n[45629];
assign t[45630] = t[45629] ^ n[45630];
assign t[45631] = t[45630] ^ n[45631];
assign t[45632] = t[45631] ^ n[45632];
assign t[45633] = t[45632] ^ n[45633];
assign t[45634] = t[45633] ^ n[45634];
assign t[45635] = t[45634] ^ n[45635];
assign t[45636] = t[45635] ^ n[45636];
assign t[45637] = t[45636] ^ n[45637];
assign t[45638] = t[45637] ^ n[45638];
assign t[45639] = t[45638] ^ n[45639];
assign t[45640] = t[45639] ^ n[45640];
assign t[45641] = t[45640] ^ n[45641];
assign t[45642] = t[45641] ^ n[45642];
assign t[45643] = t[45642] ^ n[45643];
assign t[45644] = t[45643] ^ n[45644];
assign t[45645] = t[45644] ^ n[45645];
assign t[45646] = t[45645] ^ n[45646];
assign t[45647] = t[45646] ^ n[45647];
assign t[45648] = t[45647] ^ n[45648];
assign t[45649] = t[45648] ^ n[45649];
assign t[45650] = t[45649] ^ n[45650];
assign t[45651] = t[45650] ^ n[45651];
assign t[45652] = t[45651] ^ n[45652];
assign t[45653] = t[45652] ^ n[45653];
assign t[45654] = t[45653] ^ n[45654];
assign t[45655] = t[45654] ^ n[45655];
assign t[45656] = t[45655] ^ n[45656];
assign t[45657] = t[45656] ^ n[45657];
assign t[45658] = t[45657] ^ n[45658];
assign t[45659] = t[45658] ^ n[45659];
assign t[45660] = t[45659] ^ n[45660];
assign t[45661] = t[45660] ^ n[45661];
assign t[45662] = t[45661] ^ n[45662];
assign t[45663] = t[45662] ^ n[45663];
assign t[45664] = t[45663] ^ n[45664];
assign t[45665] = t[45664] ^ n[45665];
assign t[45666] = t[45665] ^ n[45666];
assign t[45667] = t[45666] ^ n[45667];
assign t[45668] = t[45667] ^ n[45668];
assign t[45669] = t[45668] ^ n[45669];
assign t[45670] = t[45669] ^ n[45670];
assign t[45671] = t[45670] ^ n[45671];
assign t[45672] = t[45671] ^ n[45672];
assign t[45673] = t[45672] ^ n[45673];
assign t[45674] = t[45673] ^ n[45674];
assign t[45675] = t[45674] ^ n[45675];
assign t[45676] = t[45675] ^ n[45676];
assign t[45677] = t[45676] ^ n[45677];
assign t[45678] = t[45677] ^ n[45678];
assign t[45679] = t[45678] ^ n[45679];
assign t[45680] = t[45679] ^ n[45680];
assign t[45681] = t[45680] ^ n[45681];
assign t[45682] = t[45681] ^ n[45682];
assign t[45683] = t[45682] ^ n[45683];
assign t[45684] = t[45683] ^ n[45684];
assign t[45685] = t[45684] ^ n[45685];
assign t[45686] = t[45685] ^ n[45686];
assign t[45687] = t[45686] ^ n[45687];
assign t[45688] = t[45687] ^ n[45688];
assign t[45689] = t[45688] ^ n[45689];
assign t[45690] = t[45689] ^ n[45690];
assign t[45691] = t[45690] ^ n[45691];
assign t[45692] = t[45691] ^ n[45692];
assign t[45693] = t[45692] ^ n[45693];
assign t[45694] = t[45693] ^ n[45694];
assign t[45695] = t[45694] ^ n[45695];
assign t[45696] = t[45695] ^ n[45696];
assign t[45697] = t[45696] ^ n[45697];
assign t[45698] = t[45697] ^ n[45698];
assign t[45699] = t[45698] ^ n[45699];
assign t[45700] = t[45699] ^ n[45700];
assign t[45701] = t[45700] ^ n[45701];
assign t[45702] = t[45701] ^ n[45702];
assign t[45703] = t[45702] ^ n[45703];
assign t[45704] = t[45703] ^ n[45704];
assign t[45705] = t[45704] ^ n[45705];
assign t[45706] = t[45705] ^ n[45706];
assign t[45707] = t[45706] ^ n[45707];
assign t[45708] = t[45707] ^ n[45708];
assign t[45709] = t[45708] ^ n[45709];
assign t[45710] = t[45709] ^ n[45710];
assign t[45711] = t[45710] ^ n[45711];
assign t[45712] = t[45711] ^ n[45712];
assign t[45713] = t[45712] ^ n[45713];
assign t[45714] = t[45713] ^ n[45714];
assign t[45715] = t[45714] ^ n[45715];
assign t[45716] = t[45715] ^ n[45716];
assign t[45717] = t[45716] ^ n[45717];
assign t[45718] = t[45717] ^ n[45718];
assign t[45719] = t[45718] ^ n[45719];
assign t[45720] = t[45719] ^ n[45720];
assign t[45721] = t[45720] ^ n[45721];
assign t[45722] = t[45721] ^ n[45722];
assign t[45723] = t[45722] ^ n[45723];
assign t[45724] = t[45723] ^ n[45724];
assign t[45725] = t[45724] ^ n[45725];
assign t[45726] = t[45725] ^ n[45726];
assign t[45727] = t[45726] ^ n[45727];
assign t[45728] = t[45727] ^ n[45728];
assign t[45729] = t[45728] ^ n[45729];
assign t[45730] = t[45729] ^ n[45730];
assign t[45731] = t[45730] ^ n[45731];
assign t[45732] = t[45731] ^ n[45732];
assign t[45733] = t[45732] ^ n[45733];
assign t[45734] = t[45733] ^ n[45734];
assign t[45735] = t[45734] ^ n[45735];
assign t[45736] = t[45735] ^ n[45736];
assign t[45737] = t[45736] ^ n[45737];
assign t[45738] = t[45737] ^ n[45738];
assign t[45739] = t[45738] ^ n[45739];
assign t[45740] = t[45739] ^ n[45740];
assign t[45741] = t[45740] ^ n[45741];
assign t[45742] = t[45741] ^ n[45742];
assign t[45743] = t[45742] ^ n[45743];
assign t[45744] = t[45743] ^ n[45744];
assign t[45745] = t[45744] ^ n[45745];
assign t[45746] = t[45745] ^ n[45746];
assign t[45747] = t[45746] ^ n[45747];
assign t[45748] = t[45747] ^ n[45748];
assign t[45749] = t[45748] ^ n[45749];
assign t[45750] = t[45749] ^ n[45750];
assign t[45751] = t[45750] ^ n[45751];
assign t[45752] = t[45751] ^ n[45752];
assign t[45753] = t[45752] ^ n[45753];
assign t[45754] = t[45753] ^ n[45754];
assign t[45755] = t[45754] ^ n[45755];
assign t[45756] = t[45755] ^ n[45756];
assign t[45757] = t[45756] ^ n[45757];
assign t[45758] = t[45757] ^ n[45758];
assign t[45759] = t[45758] ^ n[45759];
assign t[45760] = t[45759] ^ n[45760];
assign t[45761] = t[45760] ^ n[45761];
assign t[45762] = t[45761] ^ n[45762];
assign t[45763] = t[45762] ^ n[45763];
assign t[45764] = t[45763] ^ n[45764];
assign t[45765] = t[45764] ^ n[45765];
assign t[45766] = t[45765] ^ n[45766];
assign t[45767] = t[45766] ^ n[45767];
assign t[45768] = t[45767] ^ n[45768];
assign t[45769] = t[45768] ^ n[45769];
assign t[45770] = t[45769] ^ n[45770];
assign t[45771] = t[45770] ^ n[45771];
assign t[45772] = t[45771] ^ n[45772];
assign t[45773] = t[45772] ^ n[45773];
assign t[45774] = t[45773] ^ n[45774];
assign t[45775] = t[45774] ^ n[45775];
assign t[45776] = t[45775] ^ n[45776];
assign t[45777] = t[45776] ^ n[45777];
assign t[45778] = t[45777] ^ n[45778];
assign t[45779] = t[45778] ^ n[45779];
assign t[45780] = t[45779] ^ n[45780];
assign t[45781] = t[45780] ^ n[45781];
assign t[45782] = t[45781] ^ n[45782];
assign t[45783] = t[45782] ^ n[45783];
assign t[45784] = t[45783] ^ n[45784];
assign t[45785] = t[45784] ^ n[45785];
assign t[45786] = t[45785] ^ n[45786];
assign t[45787] = t[45786] ^ n[45787];
assign t[45788] = t[45787] ^ n[45788];
assign t[45789] = t[45788] ^ n[45789];
assign t[45790] = t[45789] ^ n[45790];
assign t[45791] = t[45790] ^ n[45791];
assign t[45792] = t[45791] ^ n[45792];
assign t[45793] = t[45792] ^ n[45793];
assign t[45794] = t[45793] ^ n[45794];
assign t[45795] = t[45794] ^ n[45795];
assign t[45796] = t[45795] ^ n[45796];
assign t[45797] = t[45796] ^ n[45797];
assign t[45798] = t[45797] ^ n[45798];
assign t[45799] = t[45798] ^ n[45799];
assign t[45800] = t[45799] ^ n[45800];
assign t[45801] = t[45800] ^ n[45801];
assign t[45802] = t[45801] ^ n[45802];
assign t[45803] = t[45802] ^ n[45803];
assign t[45804] = t[45803] ^ n[45804];
assign t[45805] = t[45804] ^ n[45805];
assign t[45806] = t[45805] ^ n[45806];
assign t[45807] = t[45806] ^ n[45807];
assign t[45808] = t[45807] ^ n[45808];
assign t[45809] = t[45808] ^ n[45809];
assign t[45810] = t[45809] ^ n[45810];
assign t[45811] = t[45810] ^ n[45811];
assign t[45812] = t[45811] ^ n[45812];
assign t[45813] = t[45812] ^ n[45813];
assign t[45814] = t[45813] ^ n[45814];
assign t[45815] = t[45814] ^ n[45815];
assign t[45816] = t[45815] ^ n[45816];
assign t[45817] = t[45816] ^ n[45817];
assign t[45818] = t[45817] ^ n[45818];
assign t[45819] = t[45818] ^ n[45819];
assign t[45820] = t[45819] ^ n[45820];
assign t[45821] = t[45820] ^ n[45821];
assign t[45822] = t[45821] ^ n[45822];
assign t[45823] = t[45822] ^ n[45823];
assign t[45824] = t[45823] ^ n[45824];
assign t[45825] = t[45824] ^ n[45825];
assign t[45826] = t[45825] ^ n[45826];
assign t[45827] = t[45826] ^ n[45827];
assign t[45828] = t[45827] ^ n[45828];
assign t[45829] = t[45828] ^ n[45829];
assign t[45830] = t[45829] ^ n[45830];
assign t[45831] = t[45830] ^ n[45831];
assign t[45832] = t[45831] ^ n[45832];
assign t[45833] = t[45832] ^ n[45833];
assign t[45834] = t[45833] ^ n[45834];
assign t[45835] = t[45834] ^ n[45835];
assign t[45836] = t[45835] ^ n[45836];
assign t[45837] = t[45836] ^ n[45837];
assign t[45838] = t[45837] ^ n[45838];
assign t[45839] = t[45838] ^ n[45839];
assign t[45840] = t[45839] ^ n[45840];
assign t[45841] = t[45840] ^ n[45841];
assign t[45842] = t[45841] ^ n[45842];
assign t[45843] = t[45842] ^ n[45843];
assign t[45844] = t[45843] ^ n[45844];
assign t[45845] = t[45844] ^ n[45845];
assign t[45846] = t[45845] ^ n[45846];
assign t[45847] = t[45846] ^ n[45847];
assign t[45848] = t[45847] ^ n[45848];
assign t[45849] = t[45848] ^ n[45849];
assign t[45850] = t[45849] ^ n[45850];
assign t[45851] = t[45850] ^ n[45851];
assign t[45852] = t[45851] ^ n[45852];
assign t[45853] = t[45852] ^ n[45853];
assign t[45854] = t[45853] ^ n[45854];
assign t[45855] = t[45854] ^ n[45855];
assign t[45856] = t[45855] ^ n[45856];
assign t[45857] = t[45856] ^ n[45857];
assign t[45858] = t[45857] ^ n[45858];
assign t[45859] = t[45858] ^ n[45859];
assign t[45860] = t[45859] ^ n[45860];
assign t[45861] = t[45860] ^ n[45861];
assign t[45862] = t[45861] ^ n[45862];
assign t[45863] = t[45862] ^ n[45863];
assign t[45864] = t[45863] ^ n[45864];
assign t[45865] = t[45864] ^ n[45865];
assign t[45866] = t[45865] ^ n[45866];
assign t[45867] = t[45866] ^ n[45867];
assign t[45868] = t[45867] ^ n[45868];
assign t[45869] = t[45868] ^ n[45869];
assign t[45870] = t[45869] ^ n[45870];
assign t[45871] = t[45870] ^ n[45871];
assign t[45872] = t[45871] ^ n[45872];
assign t[45873] = t[45872] ^ n[45873];
assign t[45874] = t[45873] ^ n[45874];
assign t[45875] = t[45874] ^ n[45875];
assign t[45876] = t[45875] ^ n[45876];
assign t[45877] = t[45876] ^ n[45877];
assign t[45878] = t[45877] ^ n[45878];
assign t[45879] = t[45878] ^ n[45879];
assign t[45880] = t[45879] ^ n[45880];
assign t[45881] = t[45880] ^ n[45881];
assign t[45882] = t[45881] ^ n[45882];
assign t[45883] = t[45882] ^ n[45883];
assign t[45884] = t[45883] ^ n[45884];
assign t[45885] = t[45884] ^ n[45885];
assign t[45886] = t[45885] ^ n[45886];
assign t[45887] = t[45886] ^ n[45887];
assign t[45888] = t[45887] ^ n[45888];
assign t[45889] = t[45888] ^ n[45889];
assign t[45890] = t[45889] ^ n[45890];
assign t[45891] = t[45890] ^ n[45891];
assign t[45892] = t[45891] ^ n[45892];
assign t[45893] = t[45892] ^ n[45893];
assign t[45894] = t[45893] ^ n[45894];
assign t[45895] = t[45894] ^ n[45895];
assign t[45896] = t[45895] ^ n[45896];
assign t[45897] = t[45896] ^ n[45897];
assign t[45898] = t[45897] ^ n[45898];
assign t[45899] = t[45898] ^ n[45899];
assign t[45900] = t[45899] ^ n[45900];
assign t[45901] = t[45900] ^ n[45901];
assign t[45902] = t[45901] ^ n[45902];
assign t[45903] = t[45902] ^ n[45903];
assign t[45904] = t[45903] ^ n[45904];
assign t[45905] = t[45904] ^ n[45905];
assign t[45906] = t[45905] ^ n[45906];
assign t[45907] = t[45906] ^ n[45907];
assign t[45908] = t[45907] ^ n[45908];
assign t[45909] = t[45908] ^ n[45909];
assign t[45910] = t[45909] ^ n[45910];
assign t[45911] = t[45910] ^ n[45911];
assign t[45912] = t[45911] ^ n[45912];
assign t[45913] = t[45912] ^ n[45913];
assign t[45914] = t[45913] ^ n[45914];
assign t[45915] = t[45914] ^ n[45915];
assign t[45916] = t[45915] ^ n[45916];
assign t[45917] = t[45916] ^ n[45917];
assign t[45918] = t[45917] ^ n[45918];
assign t[45919] = t[45918] ^ n[45919];
assign t[45920] = t[45919] ^ n[45920];
assign t[45921] = t[45920] ^ n[45921];
assign t[45922] = t[45921] ^ n[45922];
assign t[45923] = t[45922] ^ n[45923];
assign t[45924] = t[45923] ^ n[45924];
assign t[45925] = t[45924] ^ n[45925];
assign t[45926] = t[45925] ^ n[45926];
assign t[45927] = t[45926] ^ n[45927];
assign t[45928] = t[45927] ^ n[45928];
assign t[45929] = t[45928] ^ n[45929];
assign t[45930] = t[45929] ^ n[45930];
assign t[45931] = t[45930] ^ n[45931];
assign t[45932] = t[45931] ^ n[45932];
assign t[45933] = t[45932] ^ n[45933];
assign t[45934] = t[45933] ^ n[45934];
assign t[45935] = t[45934] ^ n[45935];
assign t[45936] = t[45935] ^ n[45936];
assign t[45937] = t[45936] ^ n[45937];
assign t[45938] = t[45937] ^ n[45938];
assign t[45939] = t[45938] ^ n[45939];
assign t[45940] = t[45939] ^ n[45940];
assign t[45941] = t[45940] ^ n[45941];
assign t[45942] = t[45941] ^ n[45942];
assign t[45943] = t[45942] ^ n[45943];
assign t[45944] = t[45943] ^ n[45944];
assign t[45945] = t[45944] ^ n[45945];
assign t[45946] = t[45945] ^ n[45946];
assign t[45947] = t[45946] ^ n[45947];
assign t[45948] = t[45947] ^ n[45948];
assign t[45949] = t[45948] ^ n[45949];
assign t[45950] = t[45949] ^ n[45950];
assign t[45951] = t[45950] ^ n[45951];
assign t[45952] = t[45951] ^ n[45952];
assign t[45953] = t[45952] ^ n[45953];
assign t[45954] = t[45953] ^ n[45954];
assign t[45955] = t[45954] ^ n[45955];
assign t[45956] = t[45955] ^ n[45956];
assign t[45957] = t[45956] ^ n[45957];
assign t[45958] = t[45957] ^ n[45958];
assign t[45959] = t[45958] ^ n[45959];
assign t[45960] = t[45959] ^ n[45960];
assign t[45961] = t[45960] ^ n[45961];
assign t[45962] = t[45961] ^ n[45962];
assign t[45963] = t[45962] ^ n[45963];
assign t[45964] = t[45963] ^ n[45964];
assign t[45965] = t[45964] ^ n[45965];
assign t[45966] = t[45965] ^ n[45966];
assign t[45967] = t[45966] ^ n[45967];
assign t[45968] = t[45967] ^ n[45968];
assign t[45969] = t[45968] ^ n[45969];
assign t[45970] = t[45969] ^ n[45970];
assign t[45971] = t[45970] ^ n[45971];
assign t[45972] = t[45971] ^ n[45972];
assign t[45973] = t[45972] ^ n[45973];
assign t[45974] = t[45973] ^ n[45974];
assign t[45975] = t[45974] ^ n[45975];
assign t[45976] = t[45975] ^ n[45976];
assign t[45977] = t[45976] ^ n[45977];
assign t[45978] = t[45977] ^ n[45978];
assign t[45979] = t[45978] ^ n[45979];
assign t[45980] = t[45979] ^ n[45980];
assign t[45981] = t[45980] ^ n[45981];
assign t[45982] = t[45981] ^ n[45982];
assign t[45983] = t[45982] ^ n[45983];
assign t[45984] = t[45983] ^ n[45984];
assign t[45985] = t[45984] ^ n[45985];
assign t[45986] = t[45985] ^ n[45986];
assign t[45987] = t[45986] ^ n[45987];
assign t[45988] = t[45987] ^ n[45988];
assign t[45989] = t[45988] ^ n[45989];
assign t[45990] = t[45989] ^ n[45990];
assign t[45991] = t[45990] ^ n[45991];
assign t[45992] = t[45991] ^ n[45992];
assign t[45993] = t[45992] ^ n[45993];
assign t[45994] = t[45993] ^ n[45994];
assign t[45995] = t[45994] ^ n[45995];
assign t[45996] = t[45995] ^ n[45996];
assign t[45997] = t[45996] ^ n[45997];
assign t[45998] = t[45997] ^ n[45998];
assign t[45999] = t[45998] ^ n[45999];
assign t[46000] = t[45999] ^ n[46000];
assign t[46001] = t[46000] ^ n[46001];
assign t[46002] = t[46001] ^ n[46002];
assign t[46003] = t[46002] ^ n[46003];
assign t[46004] = t[46003] ^ n[46004];
assign t[46005] = t[46004] ^ n[46005];
assign t[46006] = t[46005] ^ n[46006];
assign t[46007] = t[46006] ^ n[46007];
assign t[46008] = t[46007] ^ n[46008];
assign t[46009] = t[46008] ^ n[46009];
assign t[46010] = t[46009] ^ n[46010];
assign t[46011] = t[46010] ^ n[46011];
assign t[46012] = t[46011] ^ n[46012];
assign t[46013] = t[46012] ^ n[46013];
assign t[46014] = t[46013] ^ n[46014];
assign t[46015] = t[46014] ^ n[46015];
assign t[46016] = t[46015] ^ n[46016];
assign t[46017] = t[46016] ^ n[46017];
assign t[46018] = t[46017] ^ n[46018];
assign t[46019] = t[46018] ^ n[46019];
assign t[46020] = t[46019] ^ n[46020];
assign t[46021] = t[46020] ^ n[46021];
assign t[46022] = t[46021] ^ n[46022];
assign t[46023] = t[46022] ^ n[46023];
assign t[46024] = t[46023] ^ n[46024];
assign t[46025] = t[46024] ^ n[46025];
assign t[46026] = t[46025] ^ n[46026];
assign t[46027] = t[46026] ^ n[46027];
assign t[46028] = t[46027] ^ n[46028];
assign t[46029] = t[46028] ^ n[46029];
assign t[46030] = t[46029] ^ n[46030];
assign t[46031] = t[46030] ^ n[46031];
assign t[46032] = t[46031] ^ n[46032];
assign t[46033] = t[46032] ^ n[46033];
assign t[46034] = t[46033] ^ n[46034];
assign t[46035] = t[46034] ^ n[46035];
assign t[46036] = t[46035] ^ n[46036];
assign t[46037] = t[46036] ^ n[46037];
assign t[46038] = t[46037] ^ n[46038];
assign t[46039] = t[46038] ^ n[46039];
assign t[46040] = t[46039] ^ n[46040];
assign t[46041] = t[46040] ^ n[46041];
assign t[46042] = t[46041] ^ n[46042];
assign t[46043] = t[46042] ^ n[46043];
assign t[46044] = t[46043] ^ n[46044];
assign t[46045] = t[46044] ^ n[46045];
assign t[46046] = t[46045] ^ n[46046];
assign t[46047] = t[46046] ^ n[46047];
assign t[46048] = t[46047] ^ n[46048];
assign t[46049] = t[46048] ^ n[46049];
assign t[46050] = t[46049] ^ n[46050];
assign t[46051] = t[46050] ^ n[46051];
assign t[46052] = t[46051] ^ n[46052];
assign t[46053] = t[46052] ^ n[46053];
assign t[46054] = t[46053] ^ n[46054];
assign t[46055] = t[46054] ^ n[46055];
assign t[46056] = t[46055] ^ n[46056];
assign t[46057] = t[46056] ^ n[46057];
assign t[46058] = t[46057] ^ n[46058];
assign t[46059] = t[46058] ^ n[46059];
assign t[46060] = t[46059] ^ n[46060];
assign t[46061] = t[46060] ^ n[46061];
assign t[46062] = t[46061] ^ n[46062];
assign t[46063] = t[46062] ^ n[46063];
assign t[46064] = t[46063] ^ n[46064];
assign t[46065] = t[46064] ^ n[46065];
assign t[46066] = t[46065] ^ n[46066];
assign t[46067] = t[46066] ^ n[46067];
assign t[46068] = t[46067] ^ n[46068];
assign t[46069] = t[46068] ^ n[46069];
assign t[46070] = t[46069] ^ n[46070];
assign t[46071] = t[46070] ^ n[46071];
assign t[46072] = t[46071] ^ n[46072];
assign t[46073] = t[46072] ^ n[46073];
assign t[46074] = t[46073] ^ n[46074];
assign t[46075] = t[46074] ^ n[46075];
assign t[46076] = t[46075] ^ n[46076];
assign t[46077] = t[46076] ^ n[46077];
assign t[46078] = t[46077] ^ n[46078];
assign t[46079] = t[46078] ^ n[46079];
assign t[46080] = t[46079] ^ n[46080];
assign t[46081] = t[46080] ^ n[46081];
assign t[46082] = t[46081] ^ n[46082];
assign t[46083] = t[46082] ^ n[46083];
assign t[46084] = t[46083] ^ n[46084];
assign t[46085] = t[46084] ^ n[46085];
assign t[46086] = t[46085] ^ n[46086];
assign t[46087] = t[46086] ^ n[46087];
assign t[46088] = t[46087] ^ n[46088];
assign t[46089] = t[46088] ^ n[46089];
assign t[46090] = t[46089] ^ n[46090];
assign t[46091] = t[46090] ^ n[46091];
assign t[46092] = t[46091] ^ n[46092];
assign t[46093] = t[46092] ^ n[46093];
assign t[46094] = t[46093] ^ n[46094];
assign t[46095] = t[46094] ^ n[46095];
assign t[46096] = t[46095] ^ n[46096];
assign t[46097] = t[46096] ^ n[46097];
assign t[46098] = t[46097] ^ n[46098];
assign t[46099] = t[46098] ^ n[46099];
assign t[46100] = t[46099] ^ n[46100];
assign t[46101] = t[46100] ^ n[46101];
assign t[46102] = t[46101] ^ n[46102];
assign t[46103] = t[46102] ^ n[46103];
assign t[46104] = t[46103] ^ n[46104];
assign t[46105] = t[46104] ^ n[46105];
assign t[46106] = t[46105] ^ n[46106];
assign t[46107] = t[46106] ^ n[46107];
assign t[46108] = t[46107] ^ n[46108];
assign t[46109] = t[46108] ^ n[46109];
assign t[46110] = t[46109] ^ n[46110];
assign t[46111] = t[46110] ^ n[46111];
assign t[46112] = t[46111] ^ n[46112];
assign t[46113] = t[46112] ^ n[46113];
assign t[46114] = t[46113] ^ n[46114];
assign t[46115] = t[46114] ^ n[46115];
assign t[46116] = t[46115] ^ n[46116];
assign t[46117] = t[46116] ^ n[46117];
assign t[46118] = t[46117] ^ n[46118];
assign t[46119] = t[46118] ^ n[46119];
assign t[46120] = t[46119] ^ n[46120];
assign t[46121] = t[46120] ^ n[46121];
assign t[46122] = t[46121] ^ n[46122];
assign t[46123] = t[46122] ^ n[46123];
assign t[46124] = t[46123] ^ n[46124];
assign t[46125] = t[46124] ^ n[46125];
assign t[46126] = t[46125] ^ n[46126];
assign t[46127] = t[46126] ^ n[46127];
assign t[46128] = t[46127] ^ n[46128];
assign t[46129] = t[46128] ^ n[46129];
assign t[46130] = t[46129] ^ n[46130];
assign t[46131] = t[46130] ^ n[46131];
assign t[46132] = t[46131] ^ n[46132];
assign t[46133] = t[46132] ^ n[46133];
assign t[46134] = t[46133] ^ n[46134];
assign t[46135] = t[46134] ^ n[46135];
assign t[46136] = t[46135] ^ n[46136];
assign t[46137] = t[46136] ^ n[46137];
assign t[46138] = t[46137] ^ n[46138];
assign t[46139] = t[46138] ^ n[46139];
assign t[46140] = t[46139] ^ n[46140];
assign t[46141] = t[46140] ^ n[46141];
assign t[46142] = t[46141] ^ n[46142];
assign t[46143] = t[46142] ^ n[46143];
assign t[46144] = t[46143] ^ n[46144];
assign t[46145] = t[46144] ^ n[46145];
assign t[46146] = t[46145] ^ n[46146];
assign t[46147] = t[46146] ^ n[46147];
assign t[46148] = t[46147] ^ n[46148];
assign t[46149] = t[46148] ^ n[46149];
assign t[46150] = t[46149] ^ n[46150];
assign t[46151] = t[46150] ^ n[46151];
assign t[46152] = t[46151] ^ n[46152];
assign t[46153] = t[46152] ^ n[46153];
assign t[46154] = t[46153] ^ n[46154];
assign t[46155] = t[46154] ^ n[46155];
assign t[46156] = t[46155] ^ n[46156];
assign t[46157] = t[46156] ^ n[46157];
assign t[46158] = t[46157] ^ n[46158];
assign t[46159] = t[46158] ^ n[46159];
assign t[46160] = t[46159] ^ n[46160];
assign t[46161] = t[46160] ^ n[46161];
assign t[46162] = t[46161] ^ n[46162];
assign t[46163] = t[46162] ^ n[46163];
assign t[46164] = t[46163] ^ n[46164];
assign t[46165] = t[46164] ^ n[46165];
assign t[46166] = t[46165] ^ n[46166];
assign t[46167] = t[46166] ^ n[46167];
assign t[46168] = t[46167] ^ n[46168];
assign t[46169] = t[46168] ^ n[46169];
assign t[46170] = t[46169] ^ n[46170];
assign t[46171] = t[46170] ^ n[46171];
assign t[46172] = t[46171] ^ n[46172];
assign t[46173] = t[46172] ^ n[46173];
assign t[46174] = t[46173] ^ n[46174];
assign t[46175] = t[46174] ^ n[46175];
assign t[46176] = t[46175] ^ n[46176];
assign t[46177] = t[46176] ^ n[46177];
assign t[46178] = t[46177] ^ n[46178];
assign t[46179] = t[46178] ^ n[46179];
assign t[46180] = t[46179] ^ n[46180];
assign t[46181] = t[46180] ^ n[46181];
assign t[46182] = t[46181] ^ n[46182];
assign t[46183] = t[46182] ^ n[46183];
assign t[46184] = t[46183] ^ n[46184];
assign t[46185] = t[46184] ^ n[46185];
assign t[46186] = t[46185] ^ n[46186];
assign t[46187] = t[46186] ^ n[46187];
assign t[46188] = t[46187] ^ n[46188];
assign t[46189] = t[46188] ^ n[46189];
assign t[46190] = t[46189] ^ n[46190];
assign t[46191] = t[46190] ^ n[46191];
assign t[46192] = t[46191] ^ n[46192];
assign t[46193] = t[46192] ^ n[46193];
assign t[46194] = t[46193] ^ n[46194];
assign t[46195] = t[46194] ^ n[46195];
assign t[46196] = t[46195] ^ n[46196];
assign t[46197] = t[46196] ^ n[46197];
assign t[46198] = t[46197] ^ n[46198];
assign t[46199] = t[46198] ^ n[46199];
assign t[46200] = t[46199] ^ n[46200];
assign t[46201] = t[46200] ^ n[46201];
assign t[46202] = t[46201] ^ n[46202];
assign t[46203] = t[46202] ^ n[46203];
assign t[46204] = t[46203] ^ n[46204];
assign t[46205] = t[46204] ^ n[46205];
assign t[46206] = t[46205] ^ n[46206];
assign t[46207] = t[46206] ^ n[46207];
assign t[46208] = t[46207] ^ n[46208];
assign t[46209] = t[46208] ^ n[46209];
assign t[46210] = t[46209] ^ n[46210];
assign t[46211] = t[46210] ^ n[46211];
assign t[46212] = t[46211] ^ n[46212];
assign t[46213] = t[46212] ^ n[46213];
assign t[46214] = t[46213] ^ n[46214];
assign t[46215] = t[46214] ^ n[46215];
assign t[46216] = t[46215] ^ n[46216];
assign t[46217] = t[46216] ^ n[46217];
assign t[46218] = t[46217] ^ n[46218];
assign t[46219] = t[46218] ^ n[46219];
assign t[46220] = t[46219] ^ n[46220];
assign t[46221] = t[46220] ^ n[46221];
assign t[46222] = t[46221] ^ n[46222];
assign t[46223] = t[46222] ^ n[46223];
assign t[46224] = t[46223] ^ n[46224];
assign t[46225] = t[46224] ^ n[46225];
assign t[46226] = t[46225] ^ n[46226];
assign t[46227] = t[46226] ^ n[46227];
assign t[46228] = t[46227] ^ n[46228];
assign t[46229] = t[46228] ^ n[46229];
assign t[46230] = t[46229] ^ n[46230];
assign t[46231] = t[46230] ^ n[46231];
assign t[46232] = t[46231] ^ n[46232];
assign t[46233] = t[46232] ^ n[46233];
assign t[46234] = t[46233] ^ n[46234];
assign t[46235] = t[46234] ^ n[46235];
assign t[46236] = t[46235] ^ n[46236];
assign t[46237] = t[46236] ^ n[46237];
assign t[46238] = t[46237] ^ n[46238];
assign t[46239] = t[46238] ^ n[46239];
assign t[46240] = t[46239] ^ n[46240];
assign t[46241] = t[46240] ^ n[46241];
assign t[46242] = t[46241] ^ n[46242];
assign t[46243] = t[46242] ^ n[46243];
assign t[46244] = t[46243] ^ n[46244];
assign t[46245] = t[46244] ^ n[46245];
assign t[46246] = t[46245] ^ n[46246];
assign t[46247] = t[46246] ^ n[46247];
assign t[46248] = t[46247] ^ n[46248];
assign t[46249] = t[46248] ^ n[46249];
assign t[46250] = t[46249] ^ n[46250];
assign t[46251] = t[46250] ^ n[46251];
assign t[46252] = t[46251] ^ n[46252];
assign t[46253] = t[46252] ^ n[46253];
assign t[46254] = t[46253] ^ n[46254];
assign t[46255] = t[46254] ^ n[46255];
assign t[46256] = t[46255] ^ n[46256];
assign t[46257] = t[46256] ^ n[46257];
assign t[46258] = t[46257] ^ n[46258];
assign t[46259] = t[46258] ^ n[46259];
assign t[46260] = t[46259] ^ n[46260];
assign t[46261] = t[46260] ^ n[46261];
assign t[46262] = t[46261] ^ n[46262];
assign t[46263] = t[46262] ^ n[46263];
assign t[46264] = t[46263] ^ n[46264];
assign t[46265] = t[46264] ^ n[46265];
assign t[46266] = t[46265] ^ n[46266];
assign t[46267] = t[46266] ^ n[46267];
assign t[46268] = t[46267] ^ n[46268];
assign t[46269] = t[46268] ^ n[46269];
assign t[46270] = t[46269] ^ n[46270];
assign t[46271] = t[46270] ^ n[46271];
assign t[46272] = t[46271] ^ n[46272];
assign t[46273] = t[46272] ^ n[46273];
assign t[46274] = t[46273] ^ n[46274];
assign t[46275] = t[46274] ^ n[46275];
assign t[46276] = t[46275] ^ n[46276];
assign t[46277] = t[46276] ^ n[46277];
assign t[46278] = t[46277] ^ n[46278];
assign t[46279] = t[46278] ^ n[46279];
assign t[46280] = t[46279] ^ n[46280];
assign t[46281] = t[46280] ^ n[46281];
assign t[46282] = t[46281] ^ n[46282];
assign t[46283] = t[46282] ^ n[46283];
assign t[46284] = t[46283] ^ n[46284];
assign t[46285] = t[46284] ^ n[46285];
assign t[46286] = t[46285] ^ n[46286];
assign t[46287] = t[46286] ^ n[46287];
assign t[46288] = t[46287] ^ n[46288];
assign t[46289] = t[46288] ^ n[46289];
assign t[46290] = t[46289] ^ n[46290];
assign t[46291] = t[46290] ^ n[46291];
assign t[46292] = t[46291] ^ n[46292];
assign t[46293] = t[46292] ^ n[46293];
assign t[46294] = t[46293] ^ n[46294];
assign t[46295] = t[46294] ^ n[46295];
assign t[46296] = t[46295] ^ n[46296];
assign t[46297] = t[46296] ^ n[46297];
assign t[46298] = t[46297] ^ n[46298];
assign t[46299] = t[46298] ^ n[46299];
assign t[46300] = t[46299] ^ n[46300];
assign t[46301] = t[46300] ^ n[46301];
assign t[46302] = t[46301] ^ n[46302];
assign t[46303] = t[46302] ^ n[46303];
assign t[46304] = t[46303] ^ n[46304];
assign t[46305] = t[46304] ^ n[46305];
assign t[46306] = t[46305] ^ n[46306];
assign t[46307] = t[46306] ^ n[46307];
assign t[46308] = t[46307] ^ n[46308];
assign t[46309] = t[46308] ^ n[46309];
assign t[46310] = t[46309] ^ n[46310];
assign t[46311] = t[46310] ^ n[46311];
assign t[46312] = t[46311] ^ n[46312];
assign t[46313] = t[46312] ^ n[46313];
assign t[46314] = t[46313] ^ n[46314];
assign t[46315] = t[46314] ^ n[46315];
assign t[46316] = t[46315] ^ n[46316];
assign t[46317] = t[46316] ^ n[46317];
assign t[46318] = t[46317] ^ n[46318];
assign t[46319] = t[46318] ^ n[46319];
assign t[46320] = t[46319] ^ n[46320];
assign t[46321] = t[46320] ^ n[46321];
assign t[46322] = t[46321] ^ n[46322];
assign t[46323] = t[46322] ^ n[46323];
assign t[46324] = t[46323] ^ n[46324];
assign t[46325] = t[46324] ^ n[46325];
assign t[46326] = t[46325] ^ n[46326];
assign t[46327] = t[46326] ^ n[46327];
assign t[46328] = t[46327] ^ n[46328];
assign t[46329] = t[46328] ^ n[46329];
assign t[46330] = t[46329] ^ n[46330];
assign t[46331] = t[46330] ^ n[46331];
assign t[46332] = t[46331] ^ n[46332];
assign t[46333] = t[46332] ^ n[46333];
assign t[46334] = t[46333] ^ n[46334];
assign t[46335] = t[46334] ^ n[46335];
assign t[46336] = t[46335] ^ n[46336];
assign t[46337] = t[46336] ^ n[46337];
assign t[46338] = t[46337] ^ n[46338];
assign t[46339] = t[46338] ^ n[46339];
assign t[46340] = t[46339] ^ n[46340];
assign t[46341] = t[46340] ^ n[46341];
assign t[46342] = t[46341] ^ n[46342];
assign t[46343] = t[46342] ^ n[46343];
assign t[46344] = t[46343] ^ n[46344];
assign t[46345] = t[46344] ^ n[46345];
assign t[46346] = t[46345] ^ n[46346];
assign t[46347] = t[46346] ^ n[46347];
assign t[46348] = t[46347] ^ n[46348];
assign t[46349] = t[46348] ^ n[46349];
assign t[46350] = t[46349] ^ n[46350];
assign t[46351] = t[46350] ^ n[46351];
assign t[46352] = t[46351] ^ n[46352];
assign t[46353] = t[46352] ^ n[46353];
assign t[46354] = t[46353] ^ n[46354];
assign t[46355] = t[46354] ^ n[46355];
assign t[46356] = t[46355] ^ n[46356];
assign t[46357] = t[46356] ^ n[46357];
assign t[46358] = t[46357] ^ n[46358];
assign t[46359] = t[46358] ^ n[46359];
assign t[46360] = t[46359] ^ n[46360];
assign t[46361] = t[46360] ^ n[46361];
assign t[46362] = t[46361] ^ n[46362];
assign t[46363] = t[46362] ^ n[46363];
assign t[46364] = t[46363] ^ n[46364];
assign t[46365] = t[46364] ^ n[46365];
assign t[46366] = t[46365] ^ n[46366];
assign t[46367] = t[46366] ^ n[46367];
assign t[46368] = t[46367] ^ n[46368];
assign t[46369] = t[46368] ^ n[46369];
assign t[46370] = t[46369] ^ n[46370];
assign t[46371] = t[46370] ^ n[46371];
assign t[46372] = t[46371] ^ n[46372];
assign t[46373] = t[46372] ^ n[46373];
assign t[46374] = t[46373] ^ n[46374];
assign t[46375] = t[46374] ^ n[46375];
assign t[46376] = t[46375] ^ n[46376];
assign t[46377] = t[46376] ^ n[46377];
assign t[46378] = t[46377] ^ n[46378];
assign t[46379] = t[46378] ^ n[46379];
assign t[46380] = t[46379] ^ n[46380];
assign t[46381] = t[46380] ^ n[46381];
assign t[46382] = t[46381] ^ n[46382];
assign t[46383] = t[46382] ^ n[46383];
assign t[46384] = t[46383] ^ n[46384];
assign t[46385] = t[46384] ^ n[46385];
assign t[46386] = t[46385] ^ n[46386];
assign t[46387] = t[46386] ^ n[46387];
assign t[46388] = t[46387] ^ n[46388];
assign t[46389] = t[46388] ^ n[46389];
assign t[46390] = t[46389] ^ n[46390];
assign t[46391] = t[46390] ^ n[46391];
assign t[46392] = t[46391] ^ n[46392];
assign t[46393] = t[46392] ^ n[46393];
assign t[46394] = t[46393] ^ n[46394];
assign t[46395] = t[46394] ^ n[46395];
assign t[46396] = t[46395] ^ n[46396];
assign t[46397] = t[46396] ^ n[46397];
assign t[46398] = t[46397] ^ n[46398];
assign t[46399] = t[46398] ^ n[46399];
assign t[46400] = t[46399] ^ n[46400];
assign t[46401] = t[46400] ^ n[46401];
assign t[46402] = t[46401] ^ n[46402];
assign t[46403] = t[46402] ^ n[46403];
assign t[46404] = t[46403] ^ n[46404];
assign t[46405] = t[46404] ^ n[46405];
assign t[46406] = t[46405] ^ n[46406];
assign t[46407] = t[46406] ^ n[46407];
assign t[46408] = t[46407] ^ n[46408];
assign t[46409] = t[46408] ^ n[46409];
assign t[46410] = t[46409] ^ n[46410];
assign t[46411] = t[46410] ^ n[46411];
assign t[46412] = t[46411] ^ n[46412];
assign t[46413] = t[46412] ^ n[46413];
assign t[46414] = t[46413] ^ n[46414];
assign t[46415] = t[46414] ^ n[46415];
assign t[46416] = t[46415] ^ n[46416];
assign t[46417] = t[46416] ^ n[46417];
assign t[46418] = t[46417] ^ n[46418];
assign t[46419] = t[46418] ^ n[46419];
assign t[46420] = t[46419] ^ n[46420];
assign t[46421] = t[46420] ^ n[46421];
assign t[46422] = t[46421] ^ n[46422];
assign t[46423] = t[46422] ^ n[46423];
assign t[46424] = t[46423] ^ n[46424];
assign t[46425] = t[46424] ^ n[46425];
assign t[46426] = t[46425] ^ n[46426];
assign t[46427] = t[46426] ^ n[46427];
assign t[46428] = t[46427] ^ n[46428];
assign t[46429] = t[46428] ^ n[46429];
assign t[46430] = t[46429] ^ n[46430];
assign t[46431] = t[46430] ^ n[46431];
assign t[46432] = t[46431] ^ n[46432];
assign t[46433] = t[46432] ^ n[46433];
assign t[46434] = t[46433] ^ n[46434];
assign t[46435] = t[46434] ^ n[46435];
assign t[46436] = t[46435] ^ n[46436];
assign t[46437] = t[46436] ^ n[46437];
assign t[46438] = t[46437] ^ n[46438];
assign t[46439] = t[46438] ^ n[46439];
assign t[46440] = t[46439] ^ n[46440];
assign t[46441] = t[46440] ^ n[46441];
assign t[46442] = t[46441] ^ n[46442];
assign t[46443] = t[46442] ^ n[46443];
assign t[46444] = t[46443] ^ n[46444];
assign t[46445] = t[46444] ^ n[46445];
assign t[46446] = t[46445] ^ n[46446];
assign t[46447] = t[46446] ^ n[46447];
assign t[46448] = t[46447] ^ n[46448];
assign t[46449] = t[46448] ^ n[46449];
assign t[46450] = t[46449] ^ n[46450];
assign t[46451] = t[46450] ^ n[46451];
assign t[46452] = t[46451] ^ n[46452];
assign t[46453] = t[46452] ^ n[46453];
assign t[46454] = t[46453] ^ n[46454];
assign t[46455] = t[46454] ^ n[46455];
assign t[46456] = t[46455] ^ n[46456];
assign t[46457] = t[46456] ^ n[46457];
assign t[46458] = t[46457] ^ n[46458];
assign t[46459] = t[46458] ^ n[46459];
assign t[46460] = t[46459] ^ n[46460];
assign t[46461] = t[46460] ^ n[46461];
assign t[46462] = t[46461] ^ n[46462];
assign t[46463] = t[46462] ^ n[46463];
assign t[46464] = t[46463] ^ n[46464];
assign t[46465] = t[46464] ^ n[46465];
assign t[46466] = t[46465] ^ n[46466];
assign t[46467] = t[46466] ^ n[46467];
assign t[46468] = t[46467] ^ n[46468];
assign t[46469] = t[46468] ^ n[46469];
assign t[46470] = t[46469] ^ n[46470];
assign t[46471] = t[46470] ^ n[46471];
assign t[46472] = t[46471] ^ n[46472];
assign t[46473] = t[46472] ^ n[46473];
assign t[46474] = t[46473] ^ n[46474];
assign t[46475] = t[46474] ^ n[46475];
assign t[46476] = t[46475] ^ n[46476];
assign t[46477] = t[46476] ^ n[46477];
assign t[46478] = t[46477] ^ n[46478];
assign t[46479] = t[46478] ^ n[46479];
assign t[46480] = t[46479] ^ n[46480];
assign t[46481] = t[46480] ^ n[46481];
assign t[46482] = t[46481] ^ n[46482];
assign t[46483] = t[46482] ^ n[46483];
assign t[46484] = t[46483] ^ n[46484];
assign t[46485] = t[46484] ^ n[46485];
assign t[46486] = t[46485] ^ n[46486];
assign t[46487] = t[46486] ^ n[46487];
assign t[46488] = t[46487] ^ n[46488];
assign t[46489] = t[46488] ^ n[46489];
assign t[46490] = t[46489] ^ n[46490];
assign t[46491] = t[46490] ^ n[46491];
assign t[46492] = t[46491] ^ n[46492];
assign t[46493] = t[46492] ^ n[46493];
assign t[46494] = t[46493] ^ n[46494];
assign t[46495] = t[46494] ^ n[46495];
assign t[46496] = t[46495] ^ n[46496];
assign t[46497] = t[46496] ^ n[46497];
assign t[46498] = t[46497] ^ n[46498];
assign t[46499] = t[46498] ^ n[46499];
assign t[46500] = t[46499] ^ n[46500];
assign t[46501] = t[46500] ^ n[46501];
assign t[46502] = t[46501] ^ n[46502];
assign t[46503] = t[46502] ^ n[46503];
assign t[46504] = t[46503] ^ n[46504];
assign t[46505] = t[46504] ^ n[46505];
assign t[46506] = t[46505] ^ n[46506];
assign t[46507] = t[46506] ^ n[46507];
assign t[46508] = t[46507] ^ n[46508];
assign t[46509] = t[46508] ^ n[46509];
assign t[46510] = t[46509] ^ n[46510];
assign t[46511] = t[46510] ^ n[46511];
assign t[46512] = t[46511] ^ n[46512];
assign t[46513] = t[46512] ^ n[46513];
assign t[46514] = t[46513] ^ n[46514];
assign t[46515] = t[46514] ^ n[46515];
assign t[46516] = t[46515] ^ n[46516];
assign t[46517] = t[46516] ^ n[46517];
assign t[46518] = t[46517] ^ n[46518];
assign t[46519] = t[46518] ^ n[46519];
assign t[46520] = t[46519] ^ n[46520];
assign t[46521] = t[46520] ^ n[46521];
assign t[46522] = t[46521] ^ n[46522];
assign t[46523] = t[46522] ^ n[46523];
assign t[46524] = t[46523] ^ n[46524];
assign t[46525] = t[46524] ^ n[46525];
assign t[46526] = t[46525] ^ n[46526];
assign t[46527] = t[46526] ^ n[46527];
assign t[46528] = t[46527] ^ n[46528];
assign t[46529] = t[46528] ^ n[46529];
assign t[46530] = t[46529] ^ n[46530];
assign t[46531] = t[46530] ^ n[46531];
assign t[46532] = t[46531] ^ n[46532];
assign t[46533] = t[46532] ^ n[46533];
assign t[46534] = t[46533] ^ n[46534];
assign t[46535] = t[46534] ^ n[46535];
assign t[46536] = t[46535] ^ n[46536];
assign t[46537] = t[46536] ^ n[46537];
assign t[46538] = t[46537] ^ n[46538];
assign t[46539] = t[46538] ^ n[46539];
assign t[46540] = t[46539] ^ n[46540];
assign t[46541] = t[46540] ^ n[46541];
assign t[46542] = t[46541] ^ n[46542];
assign t[46543] = t[46542] ^ n[46543];
assign t[46544] = t[46543] ^ n[46544];
assign t[46545] = t[46544] ^ n[46545];
assign t[46546] = t[46545] ^ n[46546];
assign t[46547] = t[46546] ^ n[46547];
assign t[46548] = t[46547] ^ n[46548];
assign t[46549] = t[46548] ^ n[46549];
assign t[46550] = t[46549] ^ n[46550];
assign t[46551] = t[46550] ^ n[46551];
assign t[46552] = t[46551] ^ n[46552];
assign t[46553] = t[46552] ^ n[46553];
assign t[46554] = t[46553] ^ n[46554];
assign t[46555] = t[46554] ^ n[46555];
assign t[46556] = t[46555] ^ n[46556];
assign t[46557] = t[46556] ^ n[46557];
assign t[46558] = t[46557] ^ n[46558];
assign t[46559] = t[46558] ^ n[46559];
assign t[46560] = t[46559] ^ n[46560];
assign t[46561] = t[46560] ^ n[46561];
assign t[46562] = t[46561] ^ n[46562];
assign t[46563] = t[46562] ^ n[46563];
assign t[46564] = t[46563] ^ n[46564];
assign t[46565] = t[46564] ^ n[46565];
assign t[46566] = t[46565] ^ n[46566];
assign t[46567] = t[46566] ^ n[46567];
assign t[46568] = t[46567] ^ n[46568];
assign t[46569] = t[46568] ^ n[46569];
assign t[46570] = t[46569] ^ n[46570];
assign t[46571] = t[46570] ^ n[46571];
assign t[46572] = t[46571] ^ n[46572];
assign t[46573] = t[46572] ^ n[46573];
assign t[46574] = t[46573] ^ n[46574];
assign t[46575] = t[46574] ^ n[46575];
assign t[46576] = t[46575] ^ n[46576];
assign t[46577] = t[46576] ^ n[46577];
assign t[46578] = t[46577] ^ n[46578];
assign t[46579] = t[46578] ^ n[46579];
assign t[46580] = t[46579] ^ n[46580];
assign t[46581] = t[46580] ^ n[46581];
assign t[46582] = t[46581] ^ n[46582];
assign t[46583] = t[46582] ^ n[46583];
assign t[46584] = t[46583] ^ n[46584];
assign t[46585] = t[46584] ^ n[46585];
assign t[46586] = t[46585] ^ n[46586];
assign t[46587] = t[46586] ^ n[46587];
assign t[46588] = t[46587] ^ n[46588];
assign t[46589] = t[46588] ^ n[46589];
assign t[46590] = t[46589] ^ n[46590];
assign t[46591] = t[46590] ^ n[46591];
assign t[46592] = t[46591] ^ n[46592];
assign t[46593] = t[46592] ^ n[46593];
assign t[46594] = t[46593] ^ n[46594];
assign t[46595] = t[46594] ^ n[46595];
assign t[46596] = t[46595] ^ n[46596];
assign t[46597] = t[46596] ^ n[46597];
assign t[46598] = t[46597] ^ n[46598];
assign t[46599] = t[46598] ^ n[46599];
assign t[46600] = t[46599] ^ n[46600];
assign t[46601] = t[46600] ^ n[46601];
assign t[46602] = t[46601] ^ n[46602];
assign t[46603] = t[46602] ^ n[46603];
assign t[46604] = t[46603] ^ n[46604];
assign t[46605] = t[46604] ^ n[46605];
assign t[46606] = t[46605] ^ n[46606];
assign t[46607] = t[46606] ^ n[46607];
assign t[46608] = t[46607] ^ n[46608];
assign t[46609] = t[46608] ^ n[46609];
assign t[46610] = t[46609] ^ n[46610];
assign t[46611] = t[46610] ^ n[46611];
assign t[46612] = t[46611] ^ n[46612];
assign t[46613] = t[46612] ^ n[46613];
assign t[46614] = t[46613] ^ n[46614];
assign t[46615] = t[46614] ^ n[46615];
assign t[46616] = t[46615] ^ n[46616];
assign t[46617] = t[46616] ^ n[46617];
assign t[46618] = t[46617] ^ n[46618];
assign t[46619] = t[46618] ^ n[46619];
assign t[46620] = t[46619] ^ n[46620];
assign t[46621] = t[46620] ^ n[46621];
assign t[46622] = t[46621] ^ n[46622];
assign t[46623] = t[46622] ^ n[46623];
assign t[46624] = t[46623] ^ n[46624];
assign t[46625] = t[46624] ^ n[46625];
assign t[46626] = t[46625] ^ n[46626];
assign t[46627] = t[46626] ^ n[46627];
assign t[46628] = t[46627] ^ n[46628];
assign t[46629] = t[46628] ^ n[46629];
assign t[46630] = t[46629] ^ n[46630];
assign t[46631] = t[46630] ^ n[46631];
assign t[46632] = t[46631] ^ n[46632];
assign t[46633] = t[46632] ^ n[46633];
assign t[46634] = t[46633] ^ n[46634];
assign t[46635] = t[46634] ^ n[46635];
assign t[46636] = t[46635] ^ n[46636];
assign t[46637] = t[46636] ^ n[46637];
assign t[46638] = t[46637] ^ n[46638];
assign t[46639] = t[46638] ^ n[46639];
assign t[46640] = t[46639] ^ n[46640];
assign t[46641] = t[46640] ^ n[46641];
assign t[46642] = t[46641] ^ n[46642];
assign t[46643] = t[46642] ^ n[46643];
assign t[46644] = t[46643] ^ n[46644];
assign t[46645] = t[46644] ^ n[46645];
assign t[46646] = t[46645] ^ n[46646];
assign t[46647] = t[46646] ^ n[46647];
assign t[46648] = t[46647] ^ n[46648];
assign t[46649] = t[46648] ^ n[46649];
assign t[46650] = t[46649] ^ n[46650];
assign t[46651] = t[46650] ^ n[46651];
assign t[46652] = t[46651] ^ n[46652];
assign t[46653] = t[46652] ^ n[46653];
assign t[46654] = t[46653] ^ n[46654];
assign t[46655] = t[46654] ^ n[46655];
assign t[46656] = t[46655] ^ n[46656];
assign t[46657] = t[46656] ^ n[46657];
assign t[46658] = t[46657] ^ n[46658];
assign t[46659] = t[46658] ^ n[46659];
assign t[46660] = t[46659] ^ n[46660];
assign t[46661] = t[46660] ^ n[46661];
assign t[46662] = t[46661] ^ n[46662];
assign t[46663] = t[46662] ^ n[46663];
assign t[46664] = t[46663] ^ n[46664];
assign t[46665] = t[46664] ^ n[46665];
assign t[46666] = t[46665] ^ n[46666];
assign t[46667] = t[46666] ^ n[46667];
assign t[46668] = t[46667] ^ n[46668];
assign t[46669] = t[46668] ^ n[46669];
assign t[46670] = t[46669] ^ n[46670];
assign t[46671] = t[46670] ^ n[46671];
assign t[46672] = t[46671] ^ n[46672];
assign t[46673] = t[46672] ^ n[46673];
assign t[46674] = t[46673] ^ n[46674];
assign t[46675] = t[46674] ^ n[46675];
assign t[46676] = t[46675] ^ n[46676];
assign t[46677] = t[46676] ^ n[46677];
assign t[46678] = t[46677] ^ n[46678];
assign t[46679] = t[46678] ^ n[46679];
assign t[46680] = t[46679] ^ n[46680];
assign t[46681] = t[46680] ^ n[46681];
assign t[46682] = t[46681] ^ n[46682];
assign t[46683] = t[46682] ^ n[46683];
assign t[46684] = t[46683] ^ n[46684];
assign t[46685] = t[46684] ^ n[46685];
assign t[46686] = t[46685] ^ n[46686];
assign t[46687] = t[46686] ^ n[46687];
assign t[46688] = t[46687] ^ n[46688];
assign t[46689] = t[46688] ^ n[46689];
assign t[46690] = t[46689] ^ n[46690];
assign t[46691] = t[46690] ^ n[46691];
assign t[46692] = t[46691] ^ n[46692];
assign t[46693] = t[46692] ^ n[46693];
assign t[46694] = t[46693] ^ n[46694];
assign t[46695] = t[46694] ^ n[46695];
assign t[46696] = t[46695] ^ n[46696];
assign t[46697] = t[46696] ^ n[46697];
assign t[46698] = t[46697] ^ n[46698];
assign t[46699] = t[46698] ^ n[46699];
assign t[46700] = t[46699] ^ n[46700];
assign t[46701] = t[46700] ^ n[46701];
assign t[46702] = t[46701] ^ n[46702];
assign t[46703] = t[46702] ^ n[46703];
assign t[46704] = t[46703] ^ n[46704];
assign t[46705] = t[46704] ^ n[46705];
assign t[46706] = t[46705] ^ n[46706];
assign t[46707] = t[46706] ^ n[46707];
assign t[46708] = t[46707] ^ n[46708];
assign t[46709] = t[46708] ^ n[46709];
assign t[46710] = t[46709] ^ n[46710];
assign t[46711] = t[46710] ^ n[46711];
assign t[46712] = t[46711] ^ n[46712];
assign t[46713] = t[46712] ^ n[46713];
assign t[46714] = t[46713] ^ n[46714];
assign t[46715] = t[46714] ^ n[46715];
assign t[46716] = t[46715] ^ n[46716];
assign t[46717] = t[46716] ^ n[46717];
assign t[46718] = t[46717] ^ n[46718];
assign t[46719] = t[46718] ^ n[46719];
assign t[46720] = t[46719] ^ n[46720];
assign t[46721] = t[46720] ^ n[46721];
assign t[46722] = t[46721] ^ n[46722];
assign t[46723] = t[46722] ^ n[46723];
assign t[46724] = t[46723] ^ n[46724];
assign t[46725] = t[46724] ^ n[46725];
assign t[46726] = t[46725] ^ n[46726];
assign t[46727] = t[46726] ^ n[46727];
assign t[46728] = t[46727] ^ n[46728];
assign t[46729] = t[46728] ^ n[46729];
assign t[46730] = t[46729] ^ n[46730];
assign t[46731] = t[46730] ^ n[46731];
assign t[46732] = t[46731] ^ n[46732];
assign t[46733] = t[46732] ^ n[46733];
assign t[46734] = t[46733] ^ n[46734];
assign t[46735] = t[46734] ^ n[46735];
assign t[46736] = t[46735] ^ n[46736];
assign t[46737] = t[46736] ^ n[46737];
assign t[46738] = t[46737] ^ n[46738];
assign t[46739] = t[46738] ^ n[46739];
assign t[46740] = t[46739] ^ n[46740];
assign t[46741] = t[46740] ^ n[46741];
assign t[46742] = t[46741] ^ n[46742];
assign t[46743] = t[46742] ^ n[46743];
assign t[46744] = t[46743] ^ n[46744];
assign t[46745] = t[46744] ^ n[46745];
assign t[46746] = t[46745] ^ n[46746];
assign t[46747] = t[46746] ^ n[46747];
assign t[46748] = t[46747] ^ n[46748];
assign t[46749] = t[46748] ^ n[46749];
assign t[46750] = t[46749] ^ n[46750];
assign t[46751] = t[46750] ^ n[46751];
assign t[46752] = t[46751] ^ n[46752];
assign t[46753] = t[46752] ^ n[46753];
assign t[46754] = t[46753] ^ n[46754];
assign t[46755] = t[46754] ^ n[46755];
assign t[46756] = t[46755] ^ n[46756];
assign t[46757] = t[46756] ^ n[46757];
assign t[46758] = t[46757] ^ n[46758];
assign t[46759] = t[46758] ^ n[46759];
assign t[46760] = t[46759] ^ n[46760];
assign t[46761] = t[46760] ^ n[46761];
assign t[46762] = t[46761] ^ n[46762];
assign t[46763] = t[46762] ^ n[46763];
assign t[46764] = t[46763] ^ n[46764];
assign t[46765] = t[46764] ^ n[46765];
assign t[46766] = t[46765] ^ n[46766];
assign t[46767] = t[46766] ^ n[46767];
assign t[46768] = t[46767] ^ n[46768];
assign t[46769] = t[46768] ^ n[46769];
assign t[46770] = t[46769] ^ n[46770];
assign t[46771] = t[46770] ^ n[46771];
assign t[46772] = t[46771] ^ n[46772];
assign t[46773] = t[46772] ^ n[46773];
assign t[46774] = t[46773] ^ n[46774];
assign t[46775] = t[46774] ^ n[46775];
assign t[46776] = t[46775] ^ n[46776];
assign t[46777] = t[46776] ^ n[46777];
assign t[46778] = t[46777] ^ n[46778];
assign t[46779] = t[46778] ^ n[46779];
assign t[46780] = t[46779] ^ n[46780];
assign t[46781] = t[46780] ^ n[46781];
assign t[46782] = t[46781] ^ n[46782];
assign t[46783] = t[46782] ^ n[46783];
assign t[46784] = t[46783] ^ n[46784];
assign t[46785] = t[46784] ^ n[46785];
assign t[46786] = t[46785] ^ n[46786];
assign t[46787] = t[46786] ^ n[46787];
assign t[46788] = t[46787] ^ n[46788];
assign t[46789] = t[46788] ^ n[46789];
assign t[46790] = t[46789] ^ n[46790];
assign t[46791] = t[46790] ^ n[46791];
assign t[46792] = t[46791] ^ n[46792];
assign t[46793] = t[46792] ^ n[46793];
assign t[46794] = t[46793] ^ n[46794];
assign t[46795] = t[46794] ^ n[46795];
assign t[46796] = t[46795] ^ n[46796];
assign t[46797] = t[46796] ^ n[46797];
assign t[46798] = t[46797] ^ n[46798];
assign t[46799] = t[46798] ^ n[46799];
assign t[46800] = t[46799] ^ n[46800];
assign t[46801] = t[46800] ^ n[46801];
assign t[46802] = t[46801] ^ n[46802];
assign t[46803] = t[46802] ^ n[46803];
assign t[46804] = t[46803] ^ n[46804];
assign t[46805] = t[46804] ^ n[46805];
assign t[46806] = t[46805] ^ n[46806];
assign t[46807] = t[46806] ^ n[46807];
assign t[46808] = t[46807] ^ n[46808];
assign t[46809] = t[46808] ^ n[46809];
assign t[46810] = t[46809] ^ n[46810];
assign t[46811] = t[46810] ^ n[46811];
assign t[46812] = t[46811] ^ n[46812];
assign t[46813] = t[46812] ^ n[46813];
assign t[46814] = t[46813] ^ n[46814];
assign t[46815] = t[46814] ^ n[46815];
assign t[46816] = t[46815] ^ n[46816];
assign t[46817] = t[46816] ^ n[46817];
assign t[46818] = t[46817] ^ n[46818];
assign t[46819] = t[46818] ^ n[46819];
assign t[46820] = t[46819] ^ n[46820];
assign t[46821] = t[46820] ^ n[46821];
assign t[46822] = t[46821] ^ n[46822];
assign t[46823] = t[46822] ^ n[46823];
assign t[46824] = t[46823] ^ n[46824];
assign t[46825] = t[46824] ^ n[46825];
assign t[46826] = t[46825] ^ n[46826];
assign t[46827] = t[46826] ^ n[46827];
assign t[46828] = t[46827] ^ n[46828];
assign t[46829] = t[46828] ^ n[46829];
assign t[46830] = t[46829] ^ n[46830];
assign t[46831] = t[46830] ^ n[46831];
assign t[46832] = t[46831] ^ n[46832];
assign t[46833] = t[46832] ^ n[46833];
assign t[46834] = t[46833] ^ n[46834];
assign t[46835] = t[46834] ^ n[46835];
assign t[46836] = t[46835] ^ n[46836];
assign t[46837] = t[46836] ^ n[46837];
assign t[46838] = t[46837] ^ n[46838];
assign t[46839] = t[46838] ^ n[46839];
assign t[46840] = t[46839] ^ n[46840];
assign t[46841] = t[46840] ^ n[46841];
assign t[46842] = t[46841] ^ n[46842];
assign t[46843] = t[46842] ^ n[46843];
assign t[46844] = t[46843] ^ n[46844];
assign t[46845] = t[46844] ^ n[46845];
assign t[46846] = t[46845] ^ n[46846];
assign t[46847] = t[46846] ^ n[46847];
assign t[46848] = t[46847] ^ n[46848];
assign t[46849] = t[46848] ^ n[46849];
assign t[46850] = t[46849] ^ n[46850];
assign t[46851] = t[46850] ^ n[46851];
assign t[46852] = t[46851] ^ n[46852];
assign t[46853] = t[46852] ^ n[46853];
assign t[46854] = t[46853] ^ n[46854];
assign t[46855] = t[46854] ^ n[46855];
assign t[46856] = t[46855] ^ n[46856];
assign t[46857] = t[46856] ^ n[46857];
assign t[46858] = t[46857] ^ n[46858];
assign t[46859] = t[46858] ^ n[46859];
assign t[46860] = t[46859] ^ n[46860];
assign t[46861] = t[46860] ^ n[46861];
assign t[46862] = t[46861] ^ n[46862];
assign t[46863] = t[46862] ^ n[46863];
assign t[46864] = t[46863] ^ n[46864];
assign t[46865] = t[46864] ^ n[46865];
assign t[46866] = t[46865] ^ n[46866];
assign t[46867] = t[46866] ^ n[46867];
assign t[46868] = t[46867] ^ n[46868];
assign t[46869] = t[46868] ^ n[46869];
assign t[46870] = t[46869] ^ n[46870];
assign t[46871] = t[46870] ^ n[46871];
assign t[46872] = t[46871] ^ n[46872];
assign t[46873] = t[46872] ^ n[46873];
assign t[46874] = t[46873] ^ n[46874];
assign t[46875] = t[46874] ^ n[46875];
assign t[46876] = t[46875] ^ n[46876];
assign t[46877] = t[46876] ^ n[46877];
assign t[46878] = t[46877] ^ n[46878];
assign t[46879] = t[46878] ^ n[46879];
assign t[46880] = t[46879] ^ n[46880];
assign t[46881] = t[46880] ^ n[46881];
assign t[46882] = t[46881] ^ n[46882];
assign t[46883] = t[46882] ^ n[46883];
assign t[46884] = t[46883] ^ n[46884];
assign t[46885] = t[46884] ^ n[46885];
assign t[46886] = t[46885] ^ n[46886];
assign t[46887] = t[46886] ^ n[46887];
assign t[46888] = t[46887] ^ n[46888];
assign t[46889] = t[46888] ^ n[46889];
assign t[46890] = t[46889] ^ n[46890];
assign t[46891] = t[46890] ^ n[46891];
assign t[46892] = t[46891] ^ n[46892];
assign t[46893] = t[46892] ^ n[46893];
assign t[46894] = t[46893] ^ n[46894];
assign t[46895] = t[46894] ^ n[46895];
assign t[46896] = t[46895] ^ n[46896];
assign t[46897] = t[46896] ^ n[46897];
assign t[46898] = t[46897] ^ n[46898];
assign t[46899] = t[46898] ^ n[46899];
assign t[46900] = t[46899] ^ n[46900];
assign t[46901] = t[46900] ^ n[46901];
assign t[46902] = t[46901] ^ n[46902];
assign t[46903] = t[46902] ^ n[46903];
assign t[46904] = t[46903] ^ n[46904];
assign t[46905] = t[46904] ^ n[46905];
assign t[46906] = t[46905] ^ n[46906];
assign t[46907] = t[46906] ^ n[46907];
assign t[46908] = t[46907] ^ n[46908];
assign t[46909] = t[46908] ^ n[46909];
assign t[46910] = t[46909] ^ n[46910];
assign t[46911] = t[46910] ^ n[46911];
assign t[46912] = t[46911] ^ n[46912];
assign t[46913] = t[46912] ^ n[46913];
assign t[46914] = t[46913] ^ n[46914];
assign t[46915] = t[46914] ^ n[46915];
assign t[46916] = t[46915] ^ n[46916];
assign t[46917] = t[46916] ^ n[46917];
assign t[46918] = t[46917] ^ n[46918];
assign t[46919] = t[46918] ^ n[46919];
assign t[46920] = t[46919] ^ n[46920];
assign t[46921] = t[46920] ^ n[46921];
assign t[46922] = t[46921] ^ n[46922];
assign t[46923] = t[46922] ^ n[46923];
assign t[46924] = t[46923] ^ n[46924];
assign t[46925] = t[46924] ^ n[46925];
assign t[46926] = t[46925] ^ n[46926];
assign t[46927] = t[46926] ^ n[46927];
assign t[46928] = t[46927] ^ n[46928];
assign t[46929] = t[46928] ^ n[46929];
assign t[46930] = t[46929] ^ n[46930];
assign t[46931] = t[46930] ^ n[46931];
assign t[46932] = t[46931] ^ n[46932];
assign t[46933] = t[46932] ^ n[46933];
assign t[46934] = t[46933] ^ n[46934];
assign t[46935] = t[46934] ^ n[46935];
assign t[46936] = t[46935] ^ n[46936];
assign t[46937] = t[46936] ^ n[46937];
assign t[46938] = t[46937] ^ n[46938];
assign t[46939] = t[46938] ^ n[46939];
assign t[46940] = t[46939] ^ n[46940];
assign t[46941] = t[46940] ^ n[46941];
assign t[46942] = t[46941] ^ n[46942];
assign t[46943] = t[46942] ^ n[46943];
assign t[46944] = t[46943] ^ n[46944];
assign t[46945] = t[46944] ^ n[46945];
assign t[46946] = t[46945] ^ n[46946];
assign t[46947] = t[46946] ^ n[46947];
assign t[46948] = t[46947] ^ n[46948];
assign t[46949] = t[46948] ^ n[46949];
assign t[46950] = t[46949] ^ n[46950];
assign t[46951] = t[46950] ^ n[46951];
assign t[46952] = t[46951] ^ n[46952];
assign t[46953] = t[46952] ^ n[46953];
assign t[46954] = t[46953] ^ n[46954];
assign t[46955] = t[46954] ^ n[46955];
assign t[46956] = t[46955] ^ n[46956];
assign t[46957] = t[46956] ^ n[46957];
assign t[46958] = t[46957] ^ n[46958];
assign t[46959] = t[46958] ^ n[46959];
assign t[46960] = t[46959] ^ n[46960];
assign t[46961] = t[46960] ^ n[46961];
assign t[46962] = t[46961] ^ n[46962];
assign t[46963] = t[46962] ^ n[46963];
assign t[46964] = t[46963] ^ n[46964];
assign t[46965] = t[46964] ^ n[46965];
assign t[46966] = t[46965] ^ n[46966];
assign t[46967] = t[46966] ^ n[46967];
assign t[46968] = t[46967] ^ n[46968];
assign t[46969] = t[46968] ^ n[46969];
assign t[46970] = t[46969] ^ n[46970];
assign t[46971] = t[46970] ^ n[46971];
assign t[46972] = t[46971] ^ n[46972];
assign t[46973] = t[46972] ^ n[46973];
assign t[46974] = t[46973] ^ n[46974];
assign t[46975] = t[46974] ^ n[46975];
assign t[46976] = t[46975] ^ n[46976];
assign t[46977] = t[46976] ^ n[46977];
assign t[46978] = t[46977] ^ n[46978];
assign t[46979] = t[46978] ^ n[46979];
assign t[46980] = t[46979] ^ n[46980];
assign t[46981] = t[46980] ^ n[46981];
assign t[46982] = t[46981] ^ n[46982];
assign t[46983] = t[46982] ^ n[46983];
assign t[46984] = t[46983] ^ n[46984];
assign t[46985] = t[46984] ^ n[46985];
assign t[46986] = t[46985] ^ n[46986];
assign t[46987] = t[46986] ^ n[46987];
assign t[46988] = t[46987] ^ n[46988];
assign t[46989] = t[46988] ^ n[46989];
assign t[46990] = t[46989] ^ n[46990];
assign t[46991] = t[46990] ^ n[46991];
assign t[46992] = t[46991] ^ n[46992];
assign t[46993] = t[46992] ^ n[46993];
assign t[46994] = t[46993] ^ n[46994];
assign t[46995] = t[46994] ^ n[46995];
assign t[46996] = t[46995] ^ n[46996];
assign t[46997] = t[46996] ^ n[46997];
assign t[46998] = t[46997] ^ n[46998];
assign t[46999] = t[46998] ^ n[46999];
assign t[47000] = t[46999] ^ n[47000];
assign t[47001] = t[47000] ^ n[47001];
assign t[47002] = t[47001] ^ n[47002];
assign t[47003] = t[47002] ^ n[47003];
assign t[47004] = t[47003] ^ n[47004];
assign t[47005] = t[47004] ^ n[47005];
assign t[47006] = t[47005] ^ n[47006];
assign t[47007] = t[47006] ^ n[47007];
assign t[47008] = t[47007] ^ n[47008];
assign t[47009] = t[47008] ^ n[47009];
assign t[47010] = t[47009] ^ n[47010];
assign t[47011] = t[47010] ^ n[47011];
assign t[47012] = t[47011] ^ n[47012];
assign t[47013] = t[47012] ^ n[47013];
assign t[47014] = t[47013] ^ n[47014];
assign t[47015] = t[47014] ^ n[47015];
assign t[47016] = t[47015] ^ n[47016];
assign t[47017] = t[47016] ^ n[47017];
assign t[47018] = t[47017] ^ n[47018];
assign t[47019] = t[47018] ^ n[47019];
assign t[47020] = t[47019] ^ n[47020];
assign t[47021] = t[47020] ^ n[47021];
assign t[47022] = t[47021] ^ n[47022];
assign t[47023] = t[47022] ^ n[47023];
assign t[47024] = t[47023] ^ n[47024];
assign t[47025] = t[47024] ^ n[47025];
assign t[47026] = t[47025] ^ n[47026];
assign t[47027] = t[47026] ^ n[47027];
assign t[47028] = t[47027] ^ n[47028];
assign t[47029] = t[47028] ^ n[47029];
assign t[47030] = t[47029] ^ n[47030];
assign t[47031] = t[47030] ^ n[47031];
assign t[47032] = t[47031] ^ n[47032];
assign t[47033] = t[47032] ^ n[47033];
assign t[47034] = t[47033] ^ n[47034];
assign t[47035] = t[47034] ^ n[47035];
assign t[47036] = t[47035] ^ n[47036];
assign t[47037] = t[47036] ^ n[47037];
assign t[47038] = t[47037] ^ n[47038];
assign t[47039] = t[47038] ^ n[47039];
assign t[47040] = t[47039] ^ n[47040];
assign t[47041] = t[47040] ^ n[47041];
assign t[47042] = t[47041] ^ n[47042];
assign t[47043] = t[47042] ^ n[47043];
assign t[47044] = t[47043] ^ n[47044];
assign t[47045] = t[47044] ^ n[47045];
assign t[47046] = t[47045] ^ n[47046];
assign t[47047] = t[47046] ^ n[47047];
assign t[47048] = t[47047] ^ n[47048];
assign t[47049] = t[47048] ^ n[47049];
assign t[47050] = t[47049] ^ n[47050];
assign t[47051] = t[47050] ^ n[47051];
assign t[47052] = t[47051] ^ n[47052];
assign t[47053] = t[47052] ^ n[47053];
assign t[47054] = t[47053] ^ n[47054];
assign t[47055] = t[47054] ^ n[47055];
assign t[47056] = t[47055] ^ n[47056];
assign t[47057] = t[47056] ^ n[47057];
assign t[47058] = t[47057] ^ n[47058];
assign t[47059] = t[47058] ^ n[47059];
assign t[47060] = t[47059] ^ n[47060];
assign t[47061] = t[47060] ^ n[47061];
assign t[47062] = t[47061] ^ n[47062];
assign t[47063] = t[47062] ^ n[47063];
assign t[47064] = t[47063] ^ n[47064];
assign t[47065] = t[47064] ^ n[47065];
assign t[47066] = t[47065] ^ n[47066];
assign t[47067] = t[47066] ^ n[47067];
assign t[47068] = t[47067] ^ n[47068];
assign t[47069] = t[47068] ^ n[47069];
assign t[47070] = t[47069] ^ n[47070];
assign t[47071] = t[47070] ^ n[47071];
assign t[47072] = t[47071] ^ n[47072];
assign t[47073] = t[47072] ^ n[47073];
assign t[47074] = t[47073] ^ n[47074];
assign t[47075] = t[47074] ^ n[47075];
assign t[47076] = t[47075] ^ n[47076];
assign t[47077] = t[47076] ^ n[47077];
assign t[47078] = t[47077] ^ n[47078];
assign t[47079] = t[47078] ^ n[47079];
assign t[47080] = t[47079] ^ n[47080];
assign t[47081] = t[47080] ^ n[47081];
assign t[47082] = t[47081] ^ n[47082];
assign t[47083] = t[47082] ^ n[47083];
assign t[47084] = t[47083] ^ n[47084];
assign t[47085] = t[47084] ^ n[47085];
assign t[47086] = t[47085] ^ n[47086];
assign t[47087] = t[47086] ^ n[47087];
assign t[47088] = t[47087] ^ n[47088];
assign t[47089] = t[47088] ^ n[47089];
assign t[47090] = t[47089] ^ n[47090];
assign t[47091] = t[47090] ^ n[47091];
assign t[47092] = t[47091] ^ n[47092];
assign t[47093] = t[47092] ^ n[47093];
assign t[47094] = t[47093] ^ n[47094];
assign t[47095] = t[47094] ^ n[47095];
assign t[47096] = t[47095] ^ n[47096];
assign t[47097] = t[47096] ^ n[47097];
assign t[47098] = t[47097] ^ n[47098];
assign t[47099] = t[47098] ^ n[47099];
assign t[47100] = t[47099] ^ n[47100];
assign t[47101] = t[47100] ^ n[47101];
assign t[47102] = t[47101] ^ n[47102];
assign t[47103] = t[47102] ^ n[47103];
assign t[47104] = t[47103] ^ n[47104];
assign t[47105] = t[47104] ^ n[47105];
assign t[47106] = t[47105] ^ n[47106];
assign t[47107] = t[47106] ^ n[47107];
assign t[47108] = t[47107] ^ n[47108];
assign t[47109] = t[47108] ^ n[47109];
assign t[47110] = t[47109] ^ n[47110];
assign t[47111] = t[47110] ^ n[47111];
assign t[47112] = t[47111] ^ n[47112];
assign t[47113] = t[47112] ^ n[47113];
assign t[47114] = t[47113] ^ n[47114];
assign t[47115] = t[47114] ^ n[47115];
assign t[47116] = t[47115] ^ n[47116];
assign t[47117] = t[47116] ^ n[47117];
assign t[47118] = t[47117] ^ n[47118];
assign t[47119] = t[47118] ^ n[47119];
assign t[47120] = t[47119] ^ n[47120];
assign t[47121] = t[47120] ^ n[47121];
assign t[47122] = t[47121] ^ n[47122];
assign t[47123] = t[47122] ^ n[47123];
assign t[47124] = t[47123] ^ n[47124];
assign t[47125] = t[47124] ^ n[47125];
assign t[47126] = t[47125] ^ n[47126];
assign t[47127] = t[47126] ^ n[47127];
assign t[47128] = t[47127] ^ n[47128];
assign t[47129] = t[47128] ^ n[47129];
assign t[47130] = t[47129] ^ n[47130];
assign t[47131] = t[47130] ^ n[47131];
assign t[47132] = t[47131] ^ n[47132];
assign t[47133] = t[47132] ^ n[47133];
assign t[47134] = t[47133] ^ n[47134];
assign t[47135] = t[47134] ^ n[47135];
assign t[47136] = t[47135] ^ n[47136];
assign t[47137] = t[47136] ^ n[47137];
assign t[47138] = t[47137] ^ n[47138];
assign t[47139] = t[47138] ^ n[47139];
assign t[47140] = t[47139] ^ n[47140];
assign t[47141] = t[47140] ^ n[47141];
assign t[47142] = t[47141] ^ n[47142];
assign t[47143] = t[47142] ^ n[47143];
assign t[47144] = t[47143] ^ n[47144];
assign t[47145] = t[47144] ^ n[47145];
assign t[47146] = t[47145] ^ n[47146];
assign t[47147] = t[47146] ^ n[47147];
assign t[47148] = t[47147] ^ n[47148];
assign t[47149] = t[47148] ^ n[47149];
assign t[47150] = t[47149] ^ n[47150];
assign t[47151] = t[47150] ^ n[47151];
assign t[47152] = t[47151] ^ n[47152];
assign t[47153] = t[47152] ^ n[47153];
assign t[47154] = t[47153] ^ n[47154];
assign t[47155] = t[47154] ^ n[47155];
assign t[47156] = t[47155] ^ n[47156];
assign t[47157] = t[47156] ^ n[47157];
assign t[47158] = t[47157] ^ n[47158];
assign t[47159] = t[47158] ^ n[47159];
assign t[47160] = t[47159] ^ n[47160];
assign t[47161] = t[47160] ^ n[47161];
assign t[47162] = t[47161] ^ n[47162];
assign t[47163] = t[47162] ^ n[47163];
assign t[47164] = t[47163] ^ n[47164];
assign t[47165] = t[47164] ^ n[47165];
assign t[47166] = t[47165] ^ n[47166];
assign t[47167] = t[47166] ^ n[47167];
assign t[47168] = t[47167] ^ n[47168];
assign t[47169] = t[47168] ^ n[47169];
assign t[47170] = t[47169] ^ n[47170];
assign t[47171] = t[47170] ^ n[47171];
assign t[47172] = t[47171] ^ n[47172];
assign t[47173] = t[47172] ^ n[47173];
assign t[47174] = t[47173] ^ n[47174];
assign t[47175] = t[47174] ^ n[47175];
assign t[47176] = t[47175] ^ n[47176];
assign t[47177] = t[47176] ^ n[47177];
assign t[47178] = t[47177] ^ n[47178];
assign t[47179] = t[47178] ^ n[47179];
assign t[47180] = t[47179] ^ n[47180];
assign t[47181] = t[47180] ^ n[47181];
assign t[47182] = t[47181] ^ n[47182];
assign t[47183] = t[47182] ^ n[47183];
assign t[47184] = t[47183] ^ n[47184];
assign t[47185] = t[47184] ^ n[47185];
assign t[47186] = t[47185] ^ n[47186];
assign t[47187] = t[47186] ^ n[47187];
assign t[47188] = t[47187] ^ n[47188];
assign t[47189] = t[47188] ^ n[47189];
assign t[47190] = t[47189] ^ n[47190];
assign t[47191] = t[47190] ^ n[47191];
assign t[47192] = t[47191] ^ n[47192];
assign t[47193] = t[47192] ^ n[47193];
assign t[47194] = t[47193] ^ n[47194];
assign t[47195] = t[47194] ^ n[47195];
assign t[47196] = t[47195] ^ n[47196];
assign t[47197] = t[47196] ^ n[47197];
assign t[47198] = t[47197] ^ n[47198];
assign t[47199] = t[47198] ^ n[47199];
assign t[47200] = t[47199] ^ n[47200];
assign t[47201] = t[47200] ^ n[47201];
assign t[47202] = t[47201] ^ n[47202];
assign t[47203] = t[47202] ^ n[47203];
assign t[47204] = t[47203] ^ n[47204];
assign t[47205] = t[47204] ^ n[47205];
assign t[47206] = t[47205] ^ n[47206];
assign t[47207] = t[47206] ^ n[47207];
assign t[47208] = t[47207] ^ n[47208];
assign t[47209] = t[47208] ^ n[47209];
assign t[47210] = t[47209] ^ n[47210];
assign t[47211] = t[47210] ^ n[47211];
assign t[47212] = t[47211] ^ n[47212];
assign t[47213] = t[47212] ^ n[47213];
assign t[47214] = t[47213] ^ n[47214];
assign t[47215] = t[47214] ^ n[47215];
assign t[47216] = t[47215] ^ n[47216];
assign t[47217] = t[47216] ^ n[47217];
assign t[47218] = t[47217] ^ n[47218];
assign t[47219] = t[47218] ^ n[47219];
assign t[47220] = t[47219] ^ n[47220];
assign t[47221] = t[47220] ^ n[47221];
assign t[47222] = t[47221] ^ n[47222];
assign t[47223] = t[47222] ^ n[47223];
assign t[47224] = t[47223] ^ n[47224];
assign t[47225] = t[47224] ^ n[47225];
assign t[47226] = t[47225] ^ n[47226];
assign t[47227] = t[47226] ^ n[47227];
assign t[47228] = t[47227] ^ n[47228];
assign t[47229] = t[47228] ^ n[47229];
assign t[47230] = t[47229] ^ n[47230];
assign t[47231] = t[47230] ^ n[47231];
assign t[47232] = t[47231] ^ n[47232];
assign t[47233] = t[47232] ^ n[47233];
assign t[47234] = t[47233] ^ n[47234];
assign t[47235] = t[47234] ^ n[47235];
assign t[47236] = t[47235] ^ n[47236];
assign t[47237] = t[47236] ^ n[47237];
assign t[47238] = t[47237] ^ n[47238];
assign t[47239] = t[47238] ^ n[47239];
assign t[47240] = t[47239] ^ n[47240];
assign t[47241] = t[47240] ^ n[47241];
assign t[47242] = t[47241] ^ n[47242];
assign t[47243] = t[47242] ^ n[47243];
assign t[47244] = t[47243] ^ n[47244];
assign t[47245] = t[47244] ^ n[47245];
assign t[47246] = t[47245] ^ n[47246];
assign t[47247] = t[47246] ^ n[47247];
assign t[47248] = t[47247] ^ n[47248];
assign t[47249] = t[47248] ^ n[47249];
assign t[47250] = t[47249] ^ n[47250];
assign t[47251] = t[47250] ^ n[47251];
assign t[47252] = t[47251] ^ n[47252];
assign t[47253] = t[47252] ^ n[47253];
assign t[47254] = t[47253] ^ n[47254];
assign t[47255] = t[47254] ^ n[47255];
assign t[47256] = t[47255] ^ n[47256];
assign t[47257] = t[47256] ^ n[47257];
assign t[47258] = t[47257] ^ n[47258];
assign t[47259] = t[47258] ^ n[47259];
assign t[47260] = t[47259] ^ n[47260];
assign t[47261] = t[47260] ^ n[47261];
assign t[47262] = t[47261] ^ n[47262];
assign t[47263] = t[47262] ^ n[47263];
assign t[47264] = t[47263] ^ n[47264];
assign t[47265] = t[47264] ^ n[47265];
assign t[47266] = t[47265] ^ n[47266];
assign t[47267] = t[47266] ^ n[47267];
assign t[47268] = t[47267] ^ n[47268];
assign t[47269] = t[47268] ^ n[47269];
assign t[47270] = t[47269] ^ n[47270];
assign t[47271] = t[47270] ^ n[47271];
assign t[47272] = t[47271] ^ n[47272];
assign t[47273] = t[47272] ^ n[47273];
assign t[47274] = t[47273] ^ n[47274];
assign t[47275] = t[47274] ^ n[47275];
assign t[47276] = t[47275] ^ n[47276];
assign t[47277] = t[47276] ^ n[47277];
assign t[47278] = t[47277] ^ n[47278];
assign t[47279] = t[47278] ^ n[47279];
assign t[47280] = t[47279] ^ n[47280];
assign t[47281] = t[47280] ^ n[47281];
assign t[47282] = t[47281] ^ n[47282];
assign t[47283] = t[47282] ^ n[47283];
assign t[47284] = t[47283] ^ n[47284];
assign t[47285] = t[47284] ^ n[47285];
assign t[47286] = t[47285] ^ n[47286];
assign t[47287] = t[47286] ^ n[47287];
assign t[47288] = t[47287] ^ n[47288];
assign t[47289] = t[47288] ^ n[47289];
assign t[47290] = t[47289] ^ n[47290];
assign t[47291] = t[47290] ^ n[47291];
assign t[47292] = t[47291] ^ n[47292];
assign t[47293] = t[47292] ^ n[47293];
assign t[47294] = t[47293] ^ n[47294];
assign t[47295] = t[47294] ^ n[47295];
assign t[47296] = t[47295] ^ n[47296];
assign t[47297] = t[47296] ^ n[47297];
assign t[47298] = t[47297] ^ n[47298];
assign t[47299] = t[47298] ^ n[47299];
assign t[47300] = t[47299] ^ n[47300];
assign t[47301] = t[47300] ^ n[47301];
assign t[47302] = t[47301] ^ n[47302];
assign t[47303] = t[47302] ^ n[47303];
assign t[47304] = t[47303] ^ n[47304];
assign t[47305] = t[47304] ^ n[47305];
assign t[47306] = t[47305] ^ n[47306];
assign t[47307] = t[47306] ^ n[47307];
assign t[47308] = t[47307] ^ n[47308];
assign t[47309] = t[47308] ^ n[47309];
assign t[47310] = t[47309] ^ n[47310];
assign t[47311] = t[47310] ^ n[47311];
assign t[47312] = t[47311] ^ n[47312];
assign t[47313] = t[47312] ^ n[47313];
assign t[47314] = t[47313] ^ n[47314];
assign t[47315] = t[47314] ^ n[47315];
assign t[47316] = t[47315] ^ n[47316];
assign t[47317] = t[47316] ^ n[47317];
assign t[47318] = t[47317] ^ n[47318];
assign t[47319] = t[47318] ^ n[47319];
assign t[47320] = t[47319] ^ n[47320];
assign t[47321] = t[47320] ^ n[47321];
assign t[47322] = t[47321] ^ n[47322];
assign t[47323] = t[47322] ^ n[47323];
assign t[47324] = t[47323] ^ n[47324];
assign t[47325] = t[47324] ^ n[47325];
assign t[47326] = t[47325] ^ n[47326];
assign t[47327] = t[47326] ^ n[47327];
assign t[47328] = t[47327] ^ n[47328];
assign t[47329] = t[47328] ^ n[47329];
assign t[47330] = t[47329] ^ n[47330];
assign t[47331] = t[47330] ^ n[47331];
assign t[47332] = t[47331] ^ n[47332];
assign t[47333] = t[47332] ^ n[47333];
assign t[47334] = t[47333] ^ n[47334];
assign t[47335] = t[47334] ^ n[47335];
assign t[47336] = t[47335] ^ n[47336];
assign t[47337] = t[47336] ^ n[47337];
assign t[47338] = t[47337] ^ n[47338];
assign t[47339] = t[47338] ^ n[47339];
assign t[47340] = t[47339] ^ n[47340];
assign t[47341] = t[47340] ^ n[47341];
assign t[47342] = t[47341] ^ n[47342];
assign t[47343] = t[47342] ^ n[47343];
assign t[47344] = t[47343] ^ n[47344];
assign t[47345] = t[47344] ^ n[47345];
assign t[47346] = t[47345] ^ n[47346];
assign t[47347] = t[47346] ^ n[47347];
assign t[47348] = t[47347] ^ n[47348];
assign t[47349] = t[47348] ^ n[47349];
assign t[47350] = t[47349] ^ n[47350];
assign t[47351] = t[47350] ^ n[47351];
assign t[47352] = t[47351] ^ n[47352];
assign t[47353] = t[47352] ^ n[47353];
assign t[47354] = t[47353] ^ n[47354];
assign t[47355] = t[47354] ^ n[47355];
assign t[47356] = t[47355] ^ n[47356];
assign t[47357] = t[47356] ^ n[47357];
assign t[47358] = t[47357] ^ n[47358];
assign t[47359] = t[47358] ^ n[47359];
assign t[47360] = t[47359] ^ n[47360];
assign t[47361] = t[47360] ^ n[47361];
assign t[47362] = t[47361] ^ n[47362];
assign t[47363] = t[47362] ^ n[47363];
assign t[47364] = t[47363] ^ n[47364];
assign t[47365] = t[47364] ^ n[47365];
assign t[47366] = t[47365] ^ n[47366];
assign t[47367] = t[47366] ^ n[47367];
assign t[47368] = t[47367] ^ n[47368];
assign t[47369] = t[47368] ^ n[47369];
assign t[47370] = t[47369] ^ n[47370];
assign t[47371] = t[47370] ^ n[47371];
assign t[47372] = t[47371] ^ n[47372];
assign t[47373] = t[47372] ^ n[47373];
assign t[47374] = t[47373] ^ n[47374];
assign t[47375] = t[47374] ^ n[47375];
assign t[47376] = t[47375] ^ n[47376];
assign t[47377] = t[47376] ^ n[47377];
assign t[47378] = t[47377] ^ n[47378];
assign t[47379] = t[47378] ^ n[47379];
assign t[47380] = t[47379] ^ n[47380];
assign t[47381] = t[47380] ^ n[47381];
assign t[47382] = t[47381] ^ n[47382];
assign t[47383] = t[47382] ^ n[47383];
assign t[47384] = t[47383] ^ n[47384];
assign t[47385] = t[47384] ^ n[47385];
assign t[47386] = t[47385] ^ n[47386];
assign t[47387] = t[47386] ^ n[47387];
assign t[47388] = t[47387] ^ n[47388];
assign t[47389] = t[47388] ^ n[47389];
assign t[47390] = t[47389] ^ n[47390];
assign t[47391] = t[47390] ^ n[47391];
assign t[47392] = t[47391] ^ n[47392];
assign t[47393] = t[47392] ^ n[47393];
assign t[47394] = t[47393] ^ n[47394];
assign t[47395] = t[47394] ^ n[47395];
assign t[47396] = t[47395] ^ n[47396];
assign t[47397] = t[47396] ^ n[47397];
assign t[47398] = t[47397] ^ n[47398];
assign t[47399] = t[47398] ^ n[47399];
assign t[47400] = t[47399] ^ n[47400];
assign t[47401] = t[47400] ^ n[47401];
assign t[47402] = t[47401] ^ n[47402];
assign t[47403] = t[47402] ^ n[47403];
assign t[47404] = t[47403] ^ n[47404];
assign t[47405] = t[47404] ^ n[47405];
assign t[47406] = t[47405] ^ n[47406];
assign t[47407] = t[47406] ^ n[47407];
assign t[47408] = t[47407] ^ n[47408];
assign t[47409] = t[47408] ^ n[47409];
assign t[47410] = t[47409] ^ n[47410];
assign t[47411] = t[47410] ^ n[47411];
assign t[47412] = t[47411] ^ n[47412];
assign t[47413] = t[47412] ^ n[47413];
assign t[47414] = t[47413] ^ n[47414];
assign t[47415] = t[47414] ^ n[47415];
assign t[47416] = t[47415] ^ n[47416];
assign t[47417] = t[47416] ^ n[47417];
assign t[47418] = t[47417] ^ n[47418];
assign t[47419] = t[47418] ^ n[47419];
assign t[47420] = t[47419] ^ n[47420];
assign t[47421] = t[47420] ^ n[47421];
assign t[47422] = t[47421] ^ n[47422];
assign t[47423] = t[47422] ^ n[47423];
assign t[47424] = t[47423] ^ n[47424];
assign t[47425] = t[47424] ^ n[47425];
assign t[47426] = t[47425] ^ n[47426];
assign t[47427] = t[47426] ^ n[47427];
assign t[47428] = t[47427] ^ n[47428];
assign t[47429] = t[47428] ^ n[47429];
assign t[47430] = t[47429] ^ n[47430];
assign t[47431] = t[47430] ^ n[47431];
assign t[47432] = t[47431] ^ n[47432];
assign t[47433] = t[47432] ^ n[47433];
assign t[47434] = t[47433] ^ n[47434];
assign t[47435] = t[47434] ^ n[47435];
assign t[47436] = t[47435] ^ n[47436];
assign t[47437] = t[47436] ^ n[47437];
assign t[47438] = t[47437] ^ n[47438];
assign t[47439] = t[47438] ^ n[47439];
assign t[47440] = t[47439] ^ n[47440];
assign t[47441] = t[47440] ^ n[47441];
assign t[47442] = t[47441] ^ n[47442];
assign t[47443] = t[47442] ^ n[47443];
assign t[47444] = t[47443] ^ n[47444];
assign t[47445] = t[47444] ^ n[47445];
assign t[47446] = t[47445] ^ n[47446];
assign t[47447] = t[47446] ^ n[47447];
assign t[47448] = t[47447] ^ n[47448];
assign t[47449] = t[47448] ^ n[47449];
assign t[47450] = t[47449] ^ n[47450];
assign t[47451] = t[47450] ^ n[47451];
assign t[47452] = t[47451] ^ n[47452];
assign t[47453] = t[47452] ^ n[47453];
assign t[47454] = t[47453] ^ n[47454];
assign t[47455] = t[47454] ^ n[47455];
assign t[47456] = t[47455] ^ n[47456];
assign t[47457] = t[47456] ^ n[47457];
assign t[47458] = t[47457] ^ n[47458];
assign t[47459] = t[47458] ^ n[47459];
assign t[47460] = t[47459] ^ n[47460];
assign t[47461] = t[47460] ^ n[47461];
assign t[47462] = t[47461] ^ n[47462];
assign t[47463] = t[47462] ^ n[47463];
assign t[47464] = t[47463] ^ n[47464];
assign t[47465] = t[47464] ^ n[47465];
assign t[47466] = t[47465] ^ n[47466];
assign t[47467] = t[47466] ^ n[47467];
assign t[47468] = t[47467] ^ n[47468];
assign t[47469] = t[47468] ^ n[47469];
assign t[47470] = t[47469] ^ n[47470];
assign t[47471] = t[47470] ^ n[47471];
assign t[47472] = t[47471] ^ n[47472];
assign t[47473] = t[47472] ^ n[47473];
assign t[47474] = t[47473] ^ n[47474];
assign t[47475] = t[47474] ^ n[47475];
assign t[47476] = t[47475] ^ n[47476];
assign t[47477] = t[47476] ^ n[47477];
assign t[47478] = t[47477] ^ n[47478];
assign t[47479] = t[47478] ^ n[47479];
assign t[47480] = t[47479] ^ n[47480];
assign t[47481] = t[47480] ^ n[47481];
assign t[47482] = t[47481] ^ n[47482];
assign t[47483] = t[47482] ^ n[47483];
assign t[47484] = t[47483] ^ n[47484];
assign t[47485] = t[47484] ^ n[47485];
assign t[47486] = t[47485] ^ n[47486];
assign t[47487] = t[47486] ^ n[47487];
assign t[47488] = t[47487] ^ n[47488];
assign t[47489] = t[47488] ^ n[47489];
assign t[47490] = t[47489] ^ n[47490];
assign t[47491] = t[47490] ^ n[47491];
assign t[47492] = t[47491] ^ n[47492];
assign t[47493] = t[47492] ^ n[47493];
assign t[47494] = t[47493] ^ n[47494];
assign t[47495] = t[47494] ^ n[47495];
assign t[47496] = t[47495] ^ n[47496];
assign t[47497] = t[47496] ^ n[47497];
assign t[47498] = t[47497] ^ n[47498];
assign t[47499] = t[47498] ^ n[47499];
assign t[47500] = t[47499] ^ n[47500];
assign t[47501] = t[47500] ^ n[47501];
assign t[47502] = t[47501] ^ n[47502];
assign t[47503] = t[47502] ^ n[47503];
assign t[47504] = t[47503] ^ n[47504];
assign t[47505] = t[47504] ^ n[47505];
assign t[47506] = t[47505] ^ n[47506];
assign t[47507] = t[47506] ^ n[47507];
assign t[47508] = t[47507] ^ n[47508];
assign t[47509] = t[47508] ^ n[47509];
assign t[47510] = t[47509] ^ n[47510];
assign t[47511] = t[47510] ^ n[47511];
assign t[47512] = t[47511] ^ n[47512];
assign t[47513] = t[47512] ^ n[47513];
assign t[47514] = t[47513] ^ n[47514];
assign t[47515] = t[47514] ^ n[47515];
assign t[47516] = t[47515] ^ n[47516];
assign t[47517] = t[47516] ^ n[47517];
assign t[47518] = t[47517] ^ n[47518];
assign t[47519] = t[47518] ^ n[47519];
assign t[47520] = t[47519] ^ n[47520];
assign t[47521] = t[47520] ^ n[47521];
assign t[47522] = t[47521] ^ n[47522];
assign t[47523] = t[47522] ^ n[47523];
assign t[47524] = t[47523] ^ n[47524];
assign t[47525] = t[47524] ^ n[47525];
assign t[47526] = t[47525] ^ n[47526];
assign t[47527] = t[47526] ^ n[47527];
assign t[47528] = t[47527] ^ n[47528];
assign t[47529] = t[47528] ^ n[47529];
assign t[47530] = t[47529] ^ n[47530];
assign t[47531] = t[47530] ^ n[47531];
assign t[47532] = t[47531] ^ n[47532];
assign t[47533] = t[47532] ^ n[47533];
assign t[47534] = t[47533] ^ n[47534];
assign t[47535] = t[47534] ^ n[47535];
assign t[47536] = t[47535] ^ n[47536];
assign t[47537] = t[47536] ^ n[47537];
assign t[47538] = t[47537] ^ n[47538];
assign t[47539] = t[47538] ^ n[47539];
assign t[47540] = t[47539] ^ n[47540];
assign t[47541] = t[47540] ^ n[47541];
assign t[47542] = t[47541] ^ n[47542];
assign t[47543] = t[47542] ^ n[47543];
assign t[47544] = t[47543] ^ n[47544];
assign t[47545] = t[47544] ^ n[47545];
assign t[47546] = t[47545] ^ n[47546];
assign t[47547] = t[47546] ^ n[47547];
assign t[47548] = t[47547] ^ n[47548];
assign t[47549] = t[47548] ^ n[47549];
assign t[47550] = t[47549] ^ n[47550];
assign t[47551] = t[47550] ^ n[47551];
assign t[47552] = t[47551] ^ n[47552];
assign t[47553] = t[47552] ^ n[47553];
assign t[47554] = t[47553] ^ n[47554];
assign t[47555] = t[47554] ^ n[47555];
assign t[47556] = t[47555] ^ n[47556];
assign t[47557] = t[47556] ^ n[47557];
assign t[47558] = t[47557] ^ n[47558];
assign t[47559] = t[47558] ^ n[47559];
assign t[47560] = t[47559] ^ n[47560];
assign t[47561] = t[47560] ^ n[47561];
assign t[47562] = t[47561] ^ n[47562];
assign t[47563] = t[47562] ^ n[47563];
assign t[47564] = t[47563] ^ n[47564];
assign t[47565] = t[47564] ^ n[47565];
assign t[47566] = t[47565] ^ n[47566];
assign t[47567] = t[47566] ^ n[47567];
assign t[47568] = t[47567] ^ n[47568];
assign t[47569] = t[47568] ^ n[47569];
assign t[47570] = t[47569] ^ n[47570];
assign t[47571] = t[47570] ^ n[47571];
assign t[47572] = t[47571] ^ n[47572];
assign t[47573] = t[47572] ^ n[47573];
assign t[47574] = t[47573] ^ n[47574];
assign t[47575] = t[47574] ^ n[47575];
assign t[47576] = t[47575] ^ n[47576];
assign t[47577] = t[47576] ^ n[47577];
assign t[47578] = t[47577] ^ n[47578];
assign t[47579] = t[47578] ^ n[47579];
assign t[47580] = t[47579] ^ n[47580];
assign t[47581] = t[47580] ^ n[47581];
assign t[47582] = t[47581] ^ n[47582];
assign t[47583] = t[47582] ^ n[47583];
assign t[47584] = t[47583] ^ n[47584];
assign t[47585] = t[47584] ^ n[47585];
assign t[47586] = t[47585] ^ n[47586];
assign t[47587] = t[47586] ^ n[47587];
assign t[47588] = t[47587] ^ n[47588];
assign t[47589] = t[47588] ^ n[47589];
assign t[47590] = t[47589] ^ n[47590];
assign t[47591] = t[47590] ^ n[47591];
assign t[47592] = t[47591] ^ n[47592];
assign t[47593] = t[47592] ^ n[47593];
assign t[47594] = t[47593] ^ n[47594];
assign t[47595] = t[47594] ^ n[47595];
assign t[47596] = t[47595] ^ n[47596];
assign t[47597] = t[47596] ^ n[47597];
assign t[47598] = t[47597] ^ n[47598];
assign t[47599] = t[47598] ^ n[47599];
assign t[47600] = t[47599] ^ n[47600];
assign t[47601] = t[47600] ^ n[47601];
assign t[47602] = t[47601] ^ n[47602];
assign t[47603] = t[47602] ^ n[47603];
assign t[47604] = t[47603] ^ n[47604];
assign t[47605] = t[47604] ^ n[47605];
assign t[47606] = t[47605] ^ n[47606];
assign t[47607] = t[47606] ^ n[47607];
assign t[47608] = t[47607] ^ n[47608];
assign t[47609] = t[47608] ^ n[47609];
assign t[47610] = t[47609] ^ n[47610];
assign t[47611] = t[47610] ^ n[47611];
assign t[47612] = t[47611] ^ n[47612];
assign t[47613] = t[47612] ^ n[47613];
assign t[47614] = t[47613] ^ n[47614];
assign t[47615] = t[47614] ^ n[47615];
assign t[47616] = t[47615] ^ n[47616];
assign t[47617] = t[47616] ^ n[47617];
assign t[47618] = t[47617] ^ n[47618];
assign t[47619] = t[47618] ^ n[47619];
assign t[47620] = t[47619] ^ n[47620];
assign t[47621] = t[47620] ^ n[47621];
assign t[47622] = t[47621] ^ n[47622];
assign t[47623] = t[47622] ^ n[47623];
assign t[47624] = t[47623] ^ n[47624];
assign t[47625] = t[47624] ^ n[47625];
assign t[47626] = t[47625] ^ n[47626];
assign t[47627] = t[47626] ^ n[47627];
assign t[47628] = t[47627] ^ n[47628];
assign t[47629] = t[47628] ^ n[47629];
assign t[47630] = t[47629] ^ n[47630];
assign t[47631] = t[47630] ^ n[47631];
assign t[47632] = t[47631] ^ n[47632];
assign t[47633] = t[47632] ^ n[47633];
assign t[47634] = t[47633] ^ n[47634];
assign t[47635] = t[47634] ^ n[47635];
assign t[47636] = t[47635] ^ n[47636];
assign t[47637] = t[47636] ^ n[47637];
assign t[47638] = t[47637] ^ n[47638];
assign t[47639] = t[47638] ^ n[47639];
assign t[47640] = t[47639] ^ n[47640];
assign t[47641] = t[47640] ^ n[47641];
assign t[47642] = t[47641] ^ n[47642];
assign t[47643] = t[47642] ^ n[47643];
assign t[47644] = t[47643] ^ n[47644];
assign t[47645] = t[47644] ^ n[47645];
assign t[47646] = t[47645] ^ n[47646];
assign t[47647] = t[47646] ^ n[47647];
assign t[47648] = t[47647] ^ n[47648];
assign t[47649] = t[47648] ^ n[47649];
assign t[47650] = t[47649] ^ n[47650];
assign t[47651] = t[47650] ^ n[47651];
assign t[47652] = t[47651] ^ n[47652];
assign t[47653] = t[47652] ^ n[47653];
assign t[47654] = t[47653] ^ n[47654];
assign t[47655] = t[47654] ^ n[47655];
assign t[47656] = t[47655] ^ n[47656];
assign t[47657] = t[47656] ^ n[47657];
assign t[47658] = t[47657] ^ n[47658];
assign t[47659] = t[47658] ^ n[47659];
assign t[47660] = t[47659] ^ n[47660];
assign t[47661] = t[47660] ^ n[47661];
assign t[47662] = t[47661] ^ n[47662];
assign t[47663] = t[47662] ^ n[47663];
assign t[47664] = t[47663] ^ n[47664];
assign t[47665] = t[47664] ^ n[47665];
assign t[47666] = t[47665] ^ n[47666];
assign t[47667] = t[47666] ^ n[47667];
assign t[47668] = t[47667] ^ n[47668];
assign t[47669] = t[47668] ^ n[47669];
assign t[47670] = t[47669] ^ n[47670];
assign t[47671] = t[47670] ^ n[47671];
assign t[47672] = t[47671] ^ n[47672];
assign t[47673] = t[47672] ^ n[47673];
assign t[47674] = t[47673] ^ n[47674];
assign t[47675] = t[47674] ^ n[47675];
assign t[47676] = t[47675] ^ n[47676];
assign t[47677] = t[47676] ^ n[47677];
assign t[47678] = t[47677] ^ n[47678];
assign t[47679] = t[47678] ^ n[47679];
assign t[47680] = t[47679] ^ n[47680];
assign t[47681] = t[47680] ^ n[47681];
assign t[47682] = t[47681] ^ n[47682];
assign t[47683] = t[47682] ^ n[47683];
assign t[47684] = t[47683] ^ n[47684];
assign t[47685] = t[47684] ^ n[47685];
assign t[47686] = t[47685] ^ n[47686];
assign t[47687] = t[47686] ^ n[47687];
assign t[47688] = t[47687] ^ n[47688];
assign t[47689] = t[47688] ^ n[47689];
assign t[47690] = t[47689] ^ n[47690];
assign t[47691] = t[47690] ^ n[47691];
assign t[47692] = t[47691] ^ n[47692];
assign t[47693] = t[47692] ^ n[47693];
assign t[47694] = t[47693] ^ n[47694];
assign t[47695] = t[47694] ^ n[47695];
assign t[47696] = t[47695] ^ n[47696];
assign t[47697] = t[47696] ^ n[47697];
assign t[47698] = t[47697] ^ n[47698];
assign t[47699] = t[47698] ^ n[47699];
assign t[47700] = t[47699] ^ n[47700];
assign t[47701] = t[47700] ^ n[47701];
assign t[47702] = t[47701] ^ n[47702];
assign t[47703] = t[47702] ^ n[47703];
assign t[47704] = t[47703] ^ n[47704];
assign t[47705] = t[47704] ^ n[47705];
assign t[47706] = t[47705] ^ n[47706];
assign t[47707] = t[47706] ^ n[47707];
assign t[47708] = t[47707] ^ n[47708];
assign t[47709] = t[47708] ^ n[47709];
assign t[47710] = t[47709] ^ n[47710];
assign t[47711] = t[47710] ^ n[47711];
assign t[47712] = t[47711] ^ n[47712];
assign t[47713] = t[47712] ^ n[47713];
assign t[47714] = t[47713] ^ n[47714];
assign t[47715] = t[47714] ^ n[47715];
assign t[47716] = t[47715] ^ n[47716];
assign t[47717] = t[47716] ^ n[47717];
assign t[47718] = t[47717] ^ n[47718];
assign t[47719] = t[47718] ^ n[47719];
assign t[47720] = t[47719] ^ n[47720];
assign t[47721] = t[47720] ^ n[47721];
assign t[47722] = t[47721] ^ n[47722];
assign t[47723] = t[47722] ^ n[47723];
assign t[47724] = t[47723] ^ n[47724];
assign t[47725] = t[47724] ^ n[47725];
assign t[47726] = t[47725] ^ n[47726];
assign t[47727] = t[47726] ^ n[47727];
assign t[47728] = t[47727] ^ n[47728];
assign t[47729] = t[47728] ^ n[47729];
assign t[47730] = t[47729] ^ n[47730];
assign t[47731] = t[47730] ^ n[47731];
assign t[47732] = t[47731] ^ n[47732];
assign t[47733] = t[47732] ^ n[47733];
assign t[47734] = t[47733] ^ n[47734];
assign t[47735] = t[47734] ^ n[47735];
assign t[47736] = t[47735] ^ n[47736];
assign t[47737] = t[47736] ^ n[47737];
assign t[47738] = t[47737] ^ n[47738];
assign t[47739] = t[47738] ^ n[47739];
assign t[47740] = t[47739] ^ n[47740];
assign t[47741] = t[47740] ^ n[47741];
assign t[47742] = t[47741] ^ n[47742];
assign t[47743] = t[47742] ^ n[47743];
assign t[47744] = t[47743] ^ n[47744];
assign t[47745] = t[47744] ^ n[47745];
assign t[47746] = t[47745] ^ n[47746];
assign t[47747] = t[47746] ^ n[47747];
assign t[47748] = t[47747] ^ n[47748];
assign t[47749] = t[47748] ^ n[47749];
assign t[47750] = t[47749] ^ n[47750];
assign t[47751] = t[47750] ^ n[47751];
assign t[47752] = t[47751] ^ n[47752];
assign t[47753] = t[47752] ^ n[47753];
assign t[47754] = t[47753] ^ n[47754];
assign t[47755] = t[47754] ^ n[47755];
assign t[47756] = t[47755] ^ n[47756];
assign t[47757] = t[47756] ^ n[47757];
assign t[47758] = t[47757] ^ n[47758];
assign t[47759] = t[47758] ^ n[47759];
assign t[47760] = t[47759] ^ n[47760];
assign t[47761] = t[47760] ^ n[47761];
assign t[47762] = t[47761] ^ n[47762];
assign t[47763] = t[47762] ^ n[47763];
assign t[47764] = t[47763] ^ n[47764];
assign t[47765] = t[47764] ^ n[47765];
assign t[47766] = t[47765] ^ n[47766];
assign t[47767] = t[47766] ^ n[47767];
assign t[47768] = t[47767] ^ n[47768];
assign t[47769] = t[47768] ^ n[47769];
assign t[47770] = t[47769] ^ n[47770];
assign t[47771] = t[47770] ^ n[47771];
assign t[47772] = t[47771] ^ n[47772];
assign t[47773] = t[47772] ^ n[47773];
assign t[47774] = t[47773] ^ n[47774];
assign t[47775] = t[47774] ^ n[47775];
assign t[47776] = t[47775] ^ n[47776];
assign t[47777] = t[47776] ^ n[47777];
assign t[47778] = t[47777] ^ n[47778];
assign t[47779] = t[47778] ^ n[47779];
assign t[47780] = t[47779] ^ n[47780];
assign t[47781] = t[47780] ^ n[47781];
assign t[47782] = t[47781] ^ n[47782];
assign t[47783] = t[47782] ^ n[47783];
assign t[47784] = t[47783] ^ n[47784];
assign t[47785] = t[47784] ^ n[47785];
assign t[47786] = t[47785] ^ n[47786];
assign t[47787] = t[47786] ^ n[47787];
assign t[47788] = t[47787] ^ n[47788];
assign t[47789] = t[47788] ^ n[47789];
assign t[47790] = t[47789] ^ n[47790];
assign t[47791] = t[47790] ^ n[47791];
assign t[47792] = t[47791] ^ n[47792];
assign t[47793] = t[47792] ^ n[47793];
assign t[47794] = t[47793] ^ n[47794];
assign t[47795] = t[47794] ^ n[47795];
assign t[47796] = t[47795] ^ n[47796];
assign t[47797] = t[47796] ^ n[47797];
assign t[47798] = t[47797] ^ n[47798];
assign t[47799] = t[47798] ^ n[47799];
assign t[47800] = t[47799] ^ n[47800];
assign t[47801] = t[47800] ^ n[47801];
assign t[47802] = t[47801] ^ n[47802];
assign t[47803] = t[47802] ^ n[47803];
assign t[47804] = t[47803] ^ n[47804];
assign t[47805] = t[47804] ^ n[47805];
assign t[47806] = t[47805] ^ n[47806];
assign t[47807] = t[47806] ^ n[47807];
assign t[47808] = t[47807] ^ n[47808];
assign t[47809] = t[47808] ^ n[47809];
assign t[47810] = t[47809] ^ n[47810];
assign t[47811] = t[47810] ^ n[47811];
assign t[47812] = t[47811] ^ n[47812];
assign t[47813] = t[47812] ^ n[47813];
assign t[47814] = t[47813] ^ n[47814];
assign t[47815] = t[47814] ^ n[47815];
assign t[47816] = t[47815] ^ n[47816];
assign t[47817] = t[47816] ^ n[47817];
assign t[47818] = t[47817] ^ n[47818];
assign t[47819] = t[47818] ^ n[47819];
assign t[47820] = t[47819] ^ n[47820];
assign t[47821] = t[47820] ^ n[47821];
assign t[47822] = t[47821] ^ n[47822];
assign t[47823] = t[47822] ^ n[47823];
assign t[47824] = t[47823] ^ n[47824];
assign t[47825] = t[47824] ^ n[47825];
assign t[47826] = t[47825] ^ n[47826];
assign t[47827] = t[47826] ^ n[47827];
assign t[47828] = t[47827] ^ n[47828];
assign t[47829] = t[47828] ^ n[47829];
assign t[47830] = t[47829] ^ n[47830];
assign t[47831] = t[47830] ^ n[47831];
assign t[47832] = t[47831] ^ n[47832];
assign t[47833] = t[47832] ^ n[47833];
assign t[47834] = t[47833] ^ n[47834];
assign t[47835] = t[47834] ^ n[47835];
assign t[47836] = t[47835] ^ n[47836];
assign t[47837] = t[47836] ^ n[47837];
assign t[47838] = t[47837] ^ n[47838];
assign t[47839] = t[47838] ^ n[47839];
assign t[47840] = t[47839] ^ n[47840];
assign t[47841] = t[47840] ^ n[47841];
assign t[47842] = t[47841] ^ n[47842];
assign t[47843] = t[47842] ^ n[47843];
assign t[47844] = t[47843] ^ n[47844];
assign t[47845] = t[47844] ^ n[47845];
assign t[47846] = t[47845] ^ n[47846];
assign t[47847] = t[47846] ^ n[47847];
assign t[47848] = t[47847] ^ n[47848];
assign t[47849] = t[47848] ^ n[47849];
assign t[47850] = t[47849] ^ n[47850];
assign t[47851] = t[47850] ^ n[47851];
assign t[47852] = t[47851] ^ n[47852];
assign t[47853] = t[47852] ^ n[47853];
assign t[47854] = t[47853] ^ n[47854];
assign t[47855] = t[47854] ^ n[47855];
assign t[47856] = t[47855] ^ n[47856];
assign t[47857] = t[47856] ^ n[47857];
assign t[47858] = t[47857] ^ n[47858];
assign t[47859] = t[47858] ^ n[47859];
assign t[47860] = t[47859] ^ n[47860];
assign t[47861] = t[47860] ^ n[47861];
assign t[47862] = t[47861] ^ n[47862];
assign t[47863] = t[47862] ^ n[47863];
assign t[47864] = t[47863] ^ n[47864];
assign t[47865] = t[47864] ^ n[47865];
assign t[47866] = t[47865] ^ n[47866];
assign t[47867] = t[47866] ^ n[47867];
assign t[47868] = t[47867] ^ n[47868];
assign t[47869] = t[47868] ^ n[47869];
assign t[47870] = t[47869] ^ n[47870];
assign t[47871] = t[47870] ^ n[47871];
assign t[47872] = t[47871] ^ n[47872];
assign t[47873] = t[47872] ^ n[47873];
assign t[47874] = t[47873] ^ n[47874];
assign t[47875] = t[47874] ^ n[47875];
assign t[47876] = t[47875] ^ n[47876];
assign t[47877] = t[47876] ^ n[47877];
assign t[47878] = t[47877] ^ n[47878];
assign t[47879] = t[47878] ^ n[47879];
assign t[47880] = t[47879] ^ n[47880];
assign t[47881] = t[47880] ^ n[47881];
assign t[47882] = t[47881] ^ n[47882];
assign t[47883] = t[47882] ^ n[47883];
assign t[47884] = t[47883] ^ n[47884];
assign t[47885] = t[47884] ^ n[47885];
assign t[47886] = t[47885] ^ n[47886];
assign t[47887] = t[47886] ^ n[47887];
assign t[47888] = t[47887] ^ n[47888];
assign t[47889] = t[47888] ^ n[47889];
assign t[47890] = t[47889] ^ n[47890];
assign t[47891] = t[47890] ^ n[47891];
assign t[47892] = t[47891] ^ n[47892];
assign t[47893] = t[47892] ^ n[47893];
assign t[47894] = t[47893] ^ n[47894];
assign t[47895] = t[47894] ^ n[47895];
assign t[47896] = t[47895] ^ n[47896];
assign t[47897] = t[47896] ^ n[47897];
assign t[47898] = t[47897] ^ n[47898];
assign t[47899] = t[47898] ^ n[47899];
assign t[47900] = t[47899] ^ n[47900];
assign t[47901] = t[47900] ^ n[47901];
assign t[47902] = t[47901] ^ n[47902];
assign t[47903] = t[47902] ^ n[47903];
assign t[47904] = t[47903] ^ n[47904];
assign t[47905] = t[47904] ^ n[47905];
assign t[47906] = t[47905] ^ n[47906];
assign t[47907] = t[47906] ^ n[47907];
assign t[47908] = t[47907] ^ n[47908];
assign t[47909] = t[47908] ^ n[47909];
assign t[47910] = t[47909] ^ n[47910];
assign t[47911] = t[47910] ^ n[47911];
assign t[47912] = t[47911] ^ n[47912];
assign t[47913] = t[47912] ^ n[47913];
assign t[47914] = t[47913] ^ n[47914];
assign t[47915] = t[47914] ^ n[47915];
assign t[47916] = t[47915] ^ n[47916];
assign t[47917] = t[47916] ^ n[47917];
assign t[47918] = t[47917] ^ n[47918];
assign t[47919] = t[47918] ^ n[47919];
assign t[47920] = t[47919] ^ n[47920];
assign t[47921] = t[47920] ^ n[47921];
assign t[47922] = t[47921] ^ n[47922];
assign t[47923] = t[47922] ^ n[47923];
assign t[47924] = t[47923] ^ n[47924];
assign t[47925] = t[47924] ^ n[47925];
assign t[47926] = t[47925] ^ n[47926];
assign t[47927] = t[47926] ^ n[47927];
assign t[47928] = t[47927] ^ n[47928];
assign t[47929] = t[47928] ^ n[47929];
assign t[47930] = t[47929] ^ n[47930];
assign t[47931] = t[47930] ^ n[47931];
assign t[47932] = t[47931] ^ n[47932];
assign t[47933] = t[47932] ^ n[47933];
assign t[47934] = t[47933] ^ n[47934];
assign t[47935] = t[47934] ^ n[47935];
assign t[47936] = t[47935] ^ n[47936];
assign t[47937] = t[47936] ^ n[47937];
assign t[47938] = t[47937] ^ n[47938];
assign t[47939] = t[47938] ^ n[47939];
assign t[47940] = t[47939] ^ n[47940];
assign t[47941] = t[47940] ^ n[47941];
assign t[47942] = t[47941] ^ n[47942];
assign t[47943] = t[47942] ^ n[47943];
assign t[47944] = t[47943] ^ n[47944];
assign t[47945] = t[47944] ^ n[47945];
assign t[47946] = t[47945] ^ n[47946];
assign t[47947] = t[47946] ^ n[47947];
assign t[47948] = t[47947] ^ n[47948];
assign t[47949] = t[47948] ^ n[47949];
assign t[47950] = t[47949] ^ n[47950];
assign t[47951] = t[47950] ^ n[47951];
assign t[47952] = t[47951] ^ n[47952];
assign t[47953] = t[47952] ^ n[47953];
assign t[47954] = t[47953] ^ n[47954];
assign t[47955] = t[47954] ^ n[47955];
assign t[47956] = t[47955] ^ n[47956];
assign t[47957] = t[47956] ^ n[47957];
assign t[47958] = t[47957] ^ n[47958];
assign t[47959] = t[47958] ^ n[47959];
assign t[47960] = t[47959] ^ n[47960];
assign t[47961] = t[47960] ^ n[47961];
assign t[47962] = t[47961] ^ n[47962];
assign t[47963] = t[47962] ^ n[47963];
assign t[47964] = t[47963] ^ n[47964];
assign t[47965] = t[47964] ^ n[47965];
assign t[47966] = t[47965] ^ n[47966];
assign t[47967] = t[47966] ^ n[47967];
assign t[47968] = t[47967] ^ n[47968];
assign t[47969] = t[47968] ^ n[47969];
assign t[47970] = t[47969] ^ n[47970];
assign t[47971] = t[47970] ^ n[47971];
assign t[47972] = t[47971] ^ n[47972];
assign t[47973] = t[47972] ^ n[47973];
assign t[47974] = t[47973] ^ n[47974];
assign t[47975] = t[47974] ^ n[47975];
assign t[47976] = t[47975] ^ n[47976];
assign t[47977] = t[47976] ^ n[47977];
assign t[47978] = t[47977] ^ n[47978];
assign t[47979] = t[47978] ^ n[47979];
assign t[47980] = t[47979] ^ n[47980];
assign t[47981] = t[47980] ^ n[47981];
assign t[47982] = t[47981] ^ n[47982];
assign t[47983] = t[47982] ^ n[47983];
assign t[47984] = t[47983] ^ n[47984];
assign t[47985] = t[47984] ^ n[47985];
assign t[47986] = t[47985] ^ n[47986];
assign t[47987] = t[47986] ^ n[47987];
assign t[47988] = t[47987] ^ n[47988];
assign t[47989] = t[47988] ^ n[47989];
assign t[47990] = t[47989] ^ n[47990];
assign t[47991] = t[47990] ^ n[47991];
assign t[47992] = t[47991] ^ n[47992];
assign t[47993] = t[47992] ^ n[47993];
assign t[47994] = t[47993] ^ n[47994];
assign t[47995] = t[47994] ^ n[47995];
assign t[47996] = t[47995] ^ n[47996];
assign t[47997] = t[47996] ^ n[47997];
assign t[47998] = t[47997] ^ n[47998];
assign t[47999] = t[47998] ^ n[47999];
assign t[48000] = t[47999] ^ n[48000];
assign t[48001] = t[48000] ^ n[48001];
assign t[48002] = t[48001] ^ n[48002];
assign t[48003] = t[48002] ^ n[48003];
assign t[48004] = t[48003] ^ n[48004];
assign t[48005] = t[48004] ^ n[48005];
assign t[48006] = t[48005] ^ n[48006];
assign t[48007] = t[48006] ^ n[48007];
assign t[48008] = t[48007] ^ n[48008];
assign t[48009] = t[48008] ^ n[48009];
assign t[48010] = t[48009] ^ n[48010];
assign t[48011] = t[48010] ^ n[48011];
assign t[48012] = t[48011] ^ n[48012];
assign t[48013] = t[48012] ^ n[48013];
assign t[48014] = t[48013] ^ n[48014];
assign t[48015] = t[48014] ^ n[48015];
assign t[48016] = t[48015] ^ n[48016];
assign t[48017] = t[48016] ^ n[48017];
assign t[48018] = t[48017] ^ n[48018];
assign t[48019] = t[48018] ^ n[48019];
assign t[48020] = t[48019] ^ n[48020];
assign t[48021] = t[48020] ^ n[48021];
assign t[48022] = t[48021] ^ n[48022];
assign t[48023] = t[48022] ^ n[48023];
assign t[48024] = t[48023] ^ n[48024];
assign t[48025] = t[48024] ^ n[48025];
assign t[48026] = t[48025] ^ n[48026];
assign t[48027] = t[48026] ^ n[48027];
assign t[48028] = t[48027] ^ n[48028];
assign t[48029] = t[48028] ^ n[48029];
assign t[48030] = t[48029] ^ n[48030];
assign t[48031] = t[48030] ^ n[48031];
assign t[48032] = t[48031] ^ n[48032];
assign t[48033] = t[48032] ^ n[48033];
assign t[48034] = t[48033] ^ n[48034];
assign t[48035] = t[48034] ^ n[48035];
assign t[48036] = t[48035] ^ n[48036];
assign t[48037] = t[48036] ^ n[48037];
assign t[48038] = t[48037] ^ n[48038];
assign t[48039] = t[48038] ^ n[48039];
assign t[48040] = t[48039] ^ n[48040];
assign t[48041] = t[48040] ^ n[48041];
assign t[48042] = t[48041] ^ n[48042];
assign t[48043] = t[48042] ^ n[48043];
assign t[48044] = t[48043] ^ n[48044];
assign t[48045] = t[48044] ^ n[48045];
assign t[48046] = t[48045] ^ n[48046];
assign t[48047] = t[48046] ^ n[48047];
assign t[48048] = t[48047] ^ n[48048];
assign t[48049] = t[48048] ^ n[48049];
assign t[48050] = t[48049] ^ n[48050];
assign t[48051] = t[48050] ^ n[48051];
assign t[48052] = t[48051] ^ n[48052];
assign t[48053] = t[48052] ^ n[48053];
assign t[48054] = t[48053] ^ n[48054];
assign t[48055] = t[48054] ^ n[48055];
assign t[48056] = t[48055] ^ n[48056];
assign t[48057] = t[48056] ^ n[48057];
assign t[48058] = t[48057] ^ n[48058];
assign t[48059] = t[48058] ^ n[48059];
assign t[48060] = t[48059] ^ n[48060];
assign t[48061] = t[48060] ^ n[48061];
assign t[48062] = t[48061] ^ n[48062];
assign t[48063] = t[48062] ^ n[48063];
assign t[48064] = t[48063] ^ n[48064];
assign t[48065] = t[48064] ^ n[48065];
assign t[48066] = t[48065] ^ n[48066];
assign t[48067] = t[48066] ^ n[48067];
assign t[48068] = t[48067] ^ n[48068];
assign t[48069] = t[48068] ^ n[48069];
assign t[48070] = t[48069] ^ n[48070];
assign t[48071] = t[48070] ^ n[48071];
assign t[48072] = t[48071] ^ n[48072];
assign t[48073] = t[48072] ^ n[48073];
assign t[48074] = t[48073] ^ n[48074];
assign t[48075] = t[48074] ^ n[48075];
assign t[48076] = t[48075] ^ n[48076];
assign t[48077] = t[48076] ^ n[48077];
assign t[48078] = t[48077] ^ n[48078];
assign t[48079] = t[48078] ^ n[48079];
assign t[48080] = t[48079] ^ n[48080];
assign t[48081] = t[48080] ^ n[48081];
assign t[48082] = t[48081] ^ n[48082];
assign t[48083] = t[48082] ^ n[48083];
assign t[48084] = t[48083] ^ n[48084];
assign t[48085] = t[48084] ^ n[48085];
assign t[48086] = t[48085] ^ n[48086];
assign t[48087] = t[48086] ^ n[48087];
assign t[48088] = t[48087] ^ n[48088];
assign t[48089] = t[48088] ^ n[48089];
assign t[48090] = t[48089] ^ n[48090];
assign t[48091] = t[48090] ^ n[48091];
assign t[48092] = t[48091] ^ n[48092];
assign t[48093] = t[48092] ^ n[48093];
assign t[48094] = t[48093] ^ n[48094];
assign t[48095] = t[48094] ^ n[48095];
assign t[48096] = t[48095] ^ n[48096];
assign t[48097] = t[48096] ^ n[48097];
assign t[48098] = t[48097] ^ n[48098];
assign t[48099] = t[48098] ^ n[48099];
assign t[48100] = t[48099] ^ n[48100];
assign t[48101] = t[48100] ^ n[48101];
assign t[48102] = t[48101] ^ n[48102];
assign t[48103] = t[48102] ^ n[48103];
assign t[48104] = t[48103] ^ n[48104];
assign t[48105] = t[48104] ^ n[48105];
assign t[48106] = t[48105] ^ n[48106];
assign t[48107] = t[48106] ^ n[48107];
assign t[48108] = t[48107] ^ n[48108];
assign t[48109] = t[48108] ^ n[48109];
assign t[48110] = t[48109] ^ n[48110];
assign t[48111] = t[48110] ^ n[48111];
assign t[48112] = t[48111] ^ n[48112];
assign t[48113] = t[48112] ^ n[48113];
assign t[48114] = t[48113] ^ n[48114];
assign t[48115] = t[48114] ^ n[48115];
assign t[48116] = t[48115] ^ n[48116];
assign t[48117] = t[48116] ^ n[48117];
assign t[48118] = t[48117] ^ n[48118];
assign t[48119] = t[48118] ^ n[48119];
assign t[48120] = t[48119] ^ n[48120];
assign t[48121] = t[48120] ^ n[48121];
assign t[48122] = t[48121] ^ n[48122];
assign t[48123] = t[48122] ^ n[48123];
assign t[48124] = t[48123] ^ n[48124];
assign t[48125] = t[48124] ^ n[48125];
assign t[48126] = t[48125] ^ n[48126];
assign t[48127] = t[48126] ^ n[48127];
assign t[48128] = t[48127] ^ n[48128];
assign t[48129] = t[48128] ^ n[48129];
assign t[48130] = t[48129] ^ n[48130];
assign t[48131] = t[48130] ^ n[48131];
assign t[48132] = t[48131] ^ n[48132];
assign t[48133] = t[48132] ^ n[48133];
assign t[48134] = t[48133] ^ n[48134];
assign t[48135] = t[48134] ^ n[48135];
assign t[48136] = t[48135] ^ n[48136];
assign t[48137] = t[48136] ^ n[48137];
assign t[48138] = t[48137] ^ n[48138];
assign t[48139] = t[48138] ^ n[48139];
assign t[48140] = t[48139] ^ n[48140];
assign t[48141] = t[48140] ^ n[48141];
assign t[48142] = t[48141] ^ n[48142];
assign t[48143] = t[48142] ^ n[48143];
assign t[48144] = t[48143] ^ n[48144];
assign t[48145] = t[48144] ^ n[48145];
assign t[48146] = t[48145] ^ n[48146];
assign t[48147] = t[48146] ^ n[48147];
assign t[48148] = t[48147] ^ n[48148];
assign t[48149] = t[48148] ^ n[48149];
assign t[48150] = t[48149] ^ n[48150];
assign t[48151] = t[48150] ^ n[48151];
assign t[48152] = t[48151] ^ n[48152];
assign t[48153] = t[48152] ^ n[48153];
assign t[48154] = t[48153] ^ n[48154];
assign t[48155] = t[48154] ^ n[48155];
assign t[48156] = t[48155] ^ n[48156];
assign t[48157] = t[48156] ^ n[48157];
assign t[48158] = t[48157] ^ n[48158];
assign t[48159] = t[48158] ^ n[48159];
assign t[48160] = t[48159] ^ n[48160];
assign t[48161] = t[48160] ^ n[48161];
assign t[48162] = t[48161] ^ n[48162];
assign t[48163] = t[48162] ^ n[48163];
assign t[48164] = t[48163] ^ n[48164];
assign t[48165] = t[48164] ^ n[48165];
assign t[48166] = t[48165] ^ n[48166];
assign t[48167] = t[48166] ^ n[48167];
assign t[48168] = t[48167] ^ n[48168];
assign t[48169] = t[48168] ^ n[48169];
assign t[48170] = t[48169] ^ n[48170];
assign t[48171] = t[48170] ^ n[48171];
assign t[48172] = t[48171] ^ n[48172];
assign t[48173] = t[48172] ^ n[48173];
assign t[48174] = t[48173] ^ n[48174];
assign t[48175] = t[48174] ^ n[48175];
assign t[48176] = t[48175] ^ n[48176];
assign t[48177] = t[48176] ^ n[48177];
assign t[48178] = t[48177] ^ n[48178];
assign t[48179] = t[48178] ^ n[48179];
assign t[48180] = t[48179] ^ n[48180];
assign t[48181] = t[48180] ^ n[48181];
assign t[48182] = t[48181] ^ n[48182];
assign t[48183] = t[48182] ^ n[48183];
assign t[48184] = t[48183] ^ n[48184];
assign t[48185] = t[48184] ^ n[48185];
assign t[48186] = t[48185] ^ n[48186];
assign t[48187] = t[48186] ^ n[48187];
assign t[48188] = t[48187] ^ n[48188];
assign t[48189] = t[48188] ^ n[48189];
assign t[48190] = t[48189] ^ n[48190];
assign t[48191] = t[48190] ^ n[48191];
assign t[48192] = t[48191] ^ n[48192];
assign t[48193] = t[48192] ^ n[48193];
assign t[48194] = t[48193] ^ n[48194];
assign t[48195] = t[48194] ^ n[48195];
assign t[48196] = t[48195] ^ n[48196];
assign t[48197] = t[48196] ^ n[48197];
assign t[48198] = t[48197] ^ n[48198];
assign t[48199] = t[48198] ^ n[48199];
assign t[48200] = t[48199] ^ n[48200];
assign t[48201] = t[48200] ^ n[48201];
assign t[48202] = t[48201] ^ n[48202];
assign t[48203] = t[48202] ^ n[48203];
assign t[48204] = t[48203] ^ n[48204];
assign t[48205] = t[48204] ^ n[48205];
assign t[48206] = t[48205] ^ n[48206];
assign t[48207] = t[48206] ^ n[48207];
assign t[48208] = t[48207] ^ n[48208];
assign t[48209] = t[48208] ^ n[48209];
assign t[48210] = t[48209] ^ n[48210];
assign t[48211] = t[48210] ^ n[48211];
assign t[48212] = t[48211] ^ n[48212];
assign t[48213] = t[48212] ^ n[48213];
assign t[48214] = t[48213] ^ n[48214];
assign t[48215] = t[48214] ^ n[48215];
assign t[48216] = t[48215] ^ n[48216];
assign t[48217] = t[48216] ^ n[48217];
assign t[48218] = t[48217] ^ n[48218];
assign t[48219] = t[48218] ^ n[48219];
assign t[48220] = t[48219] ^ n[48220];
assign t[48221] = t[48220] ^ n[48221];
assign t[48222] = t[48221] ^ n[48222];
assign t[48223] = t[48222] ^ n[48223];
assign t[48224] = t[48223] ^ n[48224];
assign t[48225] = t[48224] ^ n[48225];
assign t[48226] = t[48225] ^ n[48226];
assign t[48227] = t[48226] ^ n[48227];
assign t[48228] = t[48227] ^ n[48228];
assign t[48229] = t[48228] ^ n[48229];
assign t[48230] = t[48229] ^ n[48230];
assign t[48231] = t[48230] ^ n[48231];
assign t[48232] = t[48231] ^ n[48232];
assign t[48233] = t[48232] ^ n[48233];
assign t[48234] = t[48233] ^ n[48234];
assign t[48235] = t[48234] ^ n[48235];
assign t[48236] = t[48235] ^ n[48236];
assign t[48237] = t[48236] ^ n[48237];
assign t[48238] = t[48237] ^ n[48238];
assign t[48239] = t[48238] ^ n[48239];
assign t[48240] = t[48239] ^ n[48240];
assign t[48241] = t[48240] ^ n[48241];
assign t[48242] = t[48241] ^ n[48242];
assign t[48243] = t[48242] ^ n[48243];
assign t[48244] = t[48243] ^ n[48244];
assign t[48245] = t[48244] ^ n[48245];
assign t[48246] = t[48245] ^ n[48246];
assign t[48247] = t[48246] ^ n[48247];
assign t[48248] = t[48247] ^ n[48248];
assign t[48249] = t[48248] ^ n[48249];
assign t[48250] = t[48249] ^ n[48250];
assign t[48251] = t[48250] ^ n[48251];
assign t[48252] = t[48251] ^ n[48252];
assign t[48253] = t[48252] ^ n[48253];
assign t[48254] = t[48253] ^ n[48254];
assign t[48255] = t[48254] ^ n[48255];
assign t[48256] = t[48255] ^ n[48256];
assign t[48257] = t[48256] ^ n[48257];
assign t[48258] = t[48257] ^ n[48258];
assign t[48259] = t[48258] ^ n[48259];
assign t[48260] = t[48259] ^ n[48260];
assign t[48261] = t[48260] ^ n[48261];
assign t[48262] = t[48261] ^ n[48262];
assign t[48263] = t[48262] ^ n[48263];
assign t[48264] = t[48263] ^ n[48264];
assign t[48265] = t[48264] ^ n[48265];
assign t[48266] = t[48265] ^ n[48266];
assign t[48267] = t[48266] ^ n[48267];
assign t[48268] = t[48267] ^ n[48268];
assign t[48269] = t[48268] ^ n[48269];
assign t[48270] = t[48269] ^ n[48270];
assign t[48271] = t[48270] ^ n[48271];
assign t[48272] = t[48271] ^ n[48272];
assign t[48273] = t[48272] ^ n[48273];
assign t[48274] = t[48273] ^ n[48274];
assign t[48275] = t[48274] ^ n[48275];
assign t[48276] = t[48275] ^ n[48276];
assign t[48277] = t[48276] ^ n[48277];
assign t[48278] = t[48277] ^ n[48278];
assign t[48279] = t[48278] ^ n[48279];
assign t[48280] = t[48279] ^ n[48280];
assign t[48281] = t[48280] ^ n[48281];
assign t[48282] = t[48281] ^ n[48282];
assign t[48283] = t[48282] ^ n[48283];
assign t[48284] = t[48283] ^ n[48284];
assign t[48285] = t[48284] ^ n[48285];
assign t[48286] = t[48285] ^ n[48286];
assign t[48287] = t[48286] ^ n[48287];
assign t[48288] = t[48287] ^ n[48288];
assign t[48289] = t[48288] ^ n[48289];
assign t[48290] = t[48289] ^ n[48290];
assign t[48291] = t[48290] ^ n[48291];
assign t[48292] = t[48291] ^ n[48292];
assign t[48293] = t[48292] ^ n[48293];
assign t[48294] = t[48293] ^ n[48294];
assign t[48295] = t[48294] ^ n[48295];
assign t[48296] = t[48295] ^ n[48296];
assign t[48297] = t[48296] ^ n[48297];
assign t[48298] = t[48297] ^ n[48298];
assign t[48299] = t[48298] ^ n[48299];
assign t[48300] = t[48299] ^ n[48300];
assign t[48301] = t[48300] ^ n[48301];
assign t[48302] = t[48301] ^ n[48302];
assign t[48303] = t[48302] ^ n[48303];
assign t[48304] = t[48303] ^ n[48304];
assign t[48305] = t[48304] ^ n[48305];
assign t[48306] = t[48305] ^ n[48306];
assign t[48307] = t[48306] ^ n[48307];
assign t[48308] = t[48307] ^ n[48308];
assign t[48309] = t[48308] ^ n[48309];
assign t[48310] = t[48309] ^ n[48310];
assign t[48311] = t[48310] ^ n[48311];
assign t[48312] = t[48311] ^ n[48312];
assign t[48313] = t[48312] ^ n[48313];
assign t[48314] = t[48313] ^ n[48314];
assign t[48315] = t[48314] ^ n[48315];
assign t[48316] = t[48315] ^ n[48316];
assign t[48317] = t[48316] ^ n[48317];
assign t[48318] = t[48317] ^ n[48318];
assign t[48319] = t[48318] ^ n[48319];
assign t[48320] = t[48319] ^ n[48320];
assign t[48321] = t[48320] ^ n[48321];
assign t[48322] = t[48321] ^ n[48322];
assign t[48323] = t[48322] ^ n[48323];
assign t[48324] = t[48323] ^ n[48324];
assign t[48325] = t[48324] ^ n[48325];
assign t[48326] = t[48325] ^ n[48326];
assign t[48327] = t[48326] ^ n[48327];
assign t[48328] = t[48327] ^ n[48328];
assign t[48329] = t[48328] ^ n[48329];
assign t[48330] = t[48329] ^ n[48330];
assign t[48331] = t[48330] ^ n[48331];
assign t[48332] = t[48331] ^ n[48332];
assign t[48333] = t[48332] ^ n[48333];
assign t[48334] = t[48333] ^ n[48334];
assign t[48335] = t[48334] ^ n[48335];
assign t[48336] = t[48335] ^ n[48336];
assign t[48337] = t[48336] ^ n[48337];
assign t[48338] = t[48337] ^ n[48338];
assign t[48339] = t[48338] ^ n[48339];
assign t[48340] = t[48339] ^ n[48340];
assign t[48341] = t[48340] ^ n[48341];
assign t[48342] = t[48341] ^ n[48342];
assign t[48343] = t[48342] ^ n[48343];
assign t[48344] = t[48343] ^ n[48344];
assign t[48345] = t[48344] ^ n[48345];
assign t[48346] = t[48345] ^ n[48346];
assign t[48347] = t[48346] ^ n[48347];
assign t[48348] = t[48347] ^ n[48348];
assign t[48349] = t[48348] ^ n[48349];
assign t[48350] = t[48349] ^ n[48350];
assign t[48351] = t[48350] ^ n[48351];
assign t[48352] = t[48351] ^ n[48352];
assign t[48353] = t[48352] ^ n[48353];
assign t[48354] = t[48353] ^ n[48354];
assign t[48355] = t[48354] ^ n[48355];
assign t[48356] = t[48355] ^ n[48356];
assign t[48357] = t[48356] ^ n[48357];
assign t[48358] = t[48357] ^ n[48358];
assign t[48359] = t[48358] ^ n[48359];
assign t[48360] = t[48359] ^ n[48360];
assign t[48361] = t[48360] ^ n[48361];
assign t[48362] = t[48361] ^ n[48362];
assign t[48363] = t[48362] ^ n[48363];
assign t[48364] = t[48363] ^ n[48364];
assign t[48365] = t[48364] ^ n[48365];
assign t[48366] = t[48365] ^ n[48366];
assign t[48367] = t[48366] ^ n[48367];
assign t[48368] = t[48367] ^ n[48368];
assign t[48369] = t[48368] ^ n[48369];
assign t[48370] = t[48369] ^ n[48370];
assign t[48371] = t[48370] ^ n[48371];
assign t[48372] = t[48371] ^ n[48372];
assign t[48373] = t[48372] ^ n[48373];
assign t[48374] = t[48373] ^ n[48374];
assign t[48375] = t[48374] ^ n[48375];
assign t[48376] = t[48375] ^ n[48376];
assign t[48377] = t[48376] ^ n[48377];
assign t[48378] = t[48377] ^ n[48378];
assign t[48379] = t[48378] ^ n[48379];
assign t[48380] = t[48379] ^ n[48380];
assign t[48381] = t[48380] ^ n[48381];
assign t[48382] = t[48381] ^ n[48382];
assign t[48383] = t[48382] ^ n[48383];
assign t[48384] = t[48383] ^ n[48384];
assign t[48385] = t[48384] ^ n[48385];
assign t[48386] = t[48385] ^ n[48386];
assign t[48387] = t[48386] ^ n[48387];
assign t[48388] = t[48387] ^ n[48388];
assign t[48389] = t[48388] ^ n[48389];
assign t[48390] = t[48389] ^ n[48390];
assign t[48391] = t[48390] ^ n[48391];
assign t[48392] = t[48391] ^ n[48392];
assign t[48393] = t[48392] ^ n[48393];
assign t[48394] = t[48393] ^ n[48394];
assign t[48395] = t[48394] ^ n[48395];
assign t[48396] = t[48395] ^ n[48396];
assign t[48397] = t[48396] ^ n[48397];
assign t[48398] = t[48397] ^ n[48398];
assign t[48399] = t[48398] ^ n[48399];
assign t[48400] = t[48399] ^ n[48400];
assign t[48401] = t[48400] ^ n[48401];
assign t[48402] = t[48401] ^ n[48402];
assign t[48403] = t[48402] ^ n[48403];
assign t[48404] = t[48403] ^ n[48404];
assign t[48405] = t[48404] ^ n[48405];
assign t[48406] = t[48405] ^ n[48406];
assign t[48407] = t[48406] ^ n[48407];
assign t[48408] = t[48407] ^ n[48408];
assign t[48409] = t[48408] ^ n[48409];
assign t[48410] = t[48409] ^ n[48410];
assign t[48411] = t[48410] ^ n[48411];
assign t[48412] = t[48411] ^ n[48412];
assign t[48413] = t[48412] ^ n[48413];
assign t[48414] = t[48413] ^ n[48414];
assign t[48415] = t[48414] ^ n[48415];
assign t[48416] = t[48415] ^ n[48416];
assign t[48417] = t[48416] ^ n[48417];
assign t[48418] = t[48417] ^ n[48418];
assign t[48419] = t[48418] ^ n[48419];
assign t[48420] = t[48419] ^ n[48420];
assign t[48421] = t[48420] ^ n[48421];
assign t[48422] = t[48421] ^ n[48422];
assign t[48423] = t[48422] ^ n[48423];
assign t[48424] = t[48423] ^ n[48424];
assign t[48425] = t[48424] ^ n[48425];
assign t[48426] = t[48425] ^ n[48426];
assign t[48427] = t[48426] ^ n[48427];
assign t[48428] = t[48427] ^ n[48428];
assign t[48429] = t[48428] ^ n[48429];
assign t[48430] = t[48429] ^ n[48430];
assign t[48431] = t[48430] ^ n[48431];
assign t[48432] = t[48431] ^ n[48432];
assign t[48433] = t[48432] ^ n[48433];
assign t[48434] = t[48433] ^ n[48434];
assign t[48435] = t[48434] ^ n[48435];
assign t[48436] = t[48435] ^ n[48436];
assign t[48437] = t[48436] ^ n[48437];
assign t[48438] = t[48437] ^ n[48438];
assign t[48439] = t[48438] ^ n[48439];
assign t[48440] = t[48439] ^ n[48440];
assign t[48441] = t[48440] ^ n[48441];
assign t[48442] = t[48441] ^ n[48442];
assign t[48443] = t[48442] ^ n[48443];
assign t[48444] = t[48443] ^ n[48444];
assign t[48445] = t[48444] ^ n[48445];
assign t[48446] = t[48445] ^ n[48446];
assign t[48447] = t[48446] ^ n[48447];
assign t[48448] = t[48447] ^ n[48448];
assign t[48449] = t[48448] ^ n[48449];
assign t[48450] = t[48449] ^ n[48450];
assign t[48451] = t[48450] ^ n[48451];
assign t[48452] = t[48451] ^ n[48452];
assign t[48453] = t[48452] ^ n[48453];
assign t[48454] = t[48453] ^ n[48454];
assign t[48455] = t[48454] ^ n[48455];
assign t[48456] = t[48455] ^ n[48456];
assign t[48457] = t[48456] ^ n[48457];
assign t[48458] = t[48457] ^ n[48458];
assign t[48459] = t[48458] ^ n[48459];
assign t[48460] = t[48459] ^ n[48460];
assign t[48461] = t[48460] ^ n[48461];
assign t[48462] = t[48461] ^ n[48462];
assign t[48463] = t[48462] ^ n[48463];
assign t[48464] = t[48463] ^ n[48464];
assign t[48465] = t[48464] ^ n[48465];
assign t[48466] = t[48465] ^ n[48466];
assign t[48467] = t[48466] ^ n[48467];
assign t[48468] = t[48467] ^ n[48468];
assign t[48469] = t[48468] ^ n[48469];
assign t[48470] = t[48469] ^ n[48470];
assign t[48471] = t[48470] ^ n[48471];
assign t[48472] = t[48471] ^ n[48472];
assign t[48473] = t[48472] ^ n[48473];
assign t[48474] = t[48473] ^ n[48474];
assign t[48475] = t[48474] ^ n[48475];
assign t[48476] = t[48475] ^ n[48476];
assign t[48477] = t[48476] ^ n[48477];
assign t[48478] = t[48477] ^ n[48478];
assign t[48479] = t[48478] ^ n[48479];
assign t[48480] = t[48479] ^ n[48480];
assign t[48481] = t[48480] ^ n[48481];
assign t[48482] = t[48481] ^ n[48482];
assign t[48483] = t[48482] ^ n[48483];
assign t[48484] = t[48483] ^ n[48484];
assign t[48485] = t[48484] ^ n[48485];
assign t[48486] = t[48485] ^ n[48486];
assign t[48487] = t[48486] ^ n[48487];
assign t[48488] = t[48487] ^ n[48488];
assign t[48489] = t[48488] ^ n[48489];
assign t[48490] = t[48489] ^ n[48490];
assign t[48491] = t[48490] ^ n[48491];
assign t[48492] = t[48491] ^ n[48492];
assign t[48493] = t[48492] ^ n[48493];
assign t[48494] = t[48493] ^ n[48494];
assign t[48495] = t[48494] ^ n[48495];
assign t[48496] = t[48495] ^ n[48496];
assign t[48497] = t[48496] ^ n[48497];
assign t[48498] = t[48497] ^ n[48498];
assign t[48499] = t[48498] ^ n[48499];
assign t[48500] = t[48499] ^ n[48500];
assign t[48501] = t[48500] ^ n[48501];
assign t[48502] = t[48501] ^ n[48502];
assign t[48503] = t[48502] ^ n[48503];
assign t[48504] = t[48503] ^ n[48504];
assign t[48505] = t[48504] ^ n[48505];
assign t[48506] = t[48505] ^ n[48506];
assign t[48507] = t[48506] ^ n[48507];
assign t[48508] = t[48507] ^ n[48508];
assign t[48509] = t[48508] ^ n[48509];
assign t[48510] = t[48509] ^ n[48510];
assign t[48511] = t[48510] ^ n[48511];
assign t[48512] = t[48511] ^ n[48512];
assign t[48513] = t[48512] ^ n[48513];
assign t[48514] = t[48513] ^ n[48514];
assign t[48515] = t[48514] ^ n[48515];
assign t[48516] = t[48515] ^ n[48516];
assign t[48517] = t[48516] ^ n[48517];
assign t[48518] = t[48517] ^ n[48518];
assign t[48519] = t[48518] ^ n[48519];
assign t[48520] = t[48519] ^ n[48520];
assign t[48521] = t[48520] ^ n[48521];
assign t[48522] = t[48521] ^ n[48522];
assign t[48523] = t[48522] ^ n[48523];
assign t[48524] = t[48523] ^ n[48524];
assign t[48525] = t[48524] ^ n[48525];
assign t[48526] = t[48525] ^ n[48526];
assign t[48527] = t[48526] ^ n[48527];
assign t[48528] = t[48527] ^ n[48528];
assign t[48529] = t[48528] ^ n[48529];
assign t[48530] = t[48529] ^ n[48530];
assign t[48531] = t[48530] ^ n[48531];
assign t[48532] = t[48531] ^ n[48532];
assign t[48533] = t[48532] ^ n[48533];
assign t[48534] = t[48533] ^ n[48534];
assign t[48535] = t[48534] ^ n[48535];
assign t[48536] = t[48535] ^ n[48536];
assign t[48537] = t[48536] ^ n[48537];
assign t[48538] = t[48537] ^ n[48538];
assign t[48539] = t[48538] ^ n[48539];
assign t[48540] = t[48539] ^ n[48540];
assign t[48541] = t[48540] ^ n[48541];
assign t[48542] = t[48541] ^ n[48542];
assign t[48543] = t[48542] ^ n[48543];
assign t[48544] = t[48543] ^ n[48544];
assign t[48545] = t[48544] ^ n[48545];
assign t[48546] = t[48545] ^ n[48546];
assign t[48547] = t[48546] ^ n[48547];
assign t[48548] = t[48547] ^ n[48548];
assign t[48549] = t[48548] ^ n[48549];
assign t[48550] = t[48549] ^ n[48550];
assign t[48551] = t[48550] ^ n[48551];
assign t[48552] = t[48551] ^ n[48552];
assign t[48553] = t[48552] ^ n[48553];
assign t[48554] = t[48553] ^ n[48554];
assign t[48555] = t[48554] ^ n[48555];
assign t[48556] = t[48555] ^ n[48556];
assign t[48557] = t[48556] ^ n[48557];
assign t[48558] = t[48557] ^ n[48558];
assign t[48559] = t[48558] ^ n[48559];
assign t[48560] = t[48559] ^ n[48560];
assign t[48561] = t[48560] ^ n[48561];
assign t[48562] = t[48561] ^ n[48562];
assign t[48563] = t[48562] ^ n[48563];
assign t[48564] = t[48563] ^ n[48564];
assign t[48565] = t[48564] ^ n[48565];
assign t[48566] = t[48565] ^ n[48566];
assign t[48567] = t[48566] ^ n[48567];
assign t[48568] = t[48567] ^ n[48568];
assign t[48569] = t[48568] ^ n[48569];
assign t[48570] = t[48569] ^ n[48570];
assign t[48571] = t[48570] ^ n[48571];
assign t[48572] = t[48571] ^ n[48572];
assign t[48573] = t[48572] ^ n[48573];
assign t[48574] = t[48573] ^ n[48574];
assign t[48575] = t[48574] ^ n[48575];
assign t[48576] = t[48575] ^ n[48576];
assign t[48577] = t[48576] ^ n[48577];
assign t[48578] = t[48577] ^ n[48578];
assign t[48579] = t[48578] ^ n[48579];
assign t[48580] = t[48579] ^ n[48580];
assign t[48581] = t[48580] ^ n[48581];
assign t[48582] = t[48581] ^ n[48582];
assign t[48583] = t[48582] ^ n[48583];
assign t[48584] = t[48583] ^ n[48584];
assign t[48585] = t[48584] ^ n[48585];
assign t[48586] = t[48585] ^ n[48586];
assign t[48587] = t[48586] ^ n[48587];
assign t[48588] = t[48587] ^ n[48588];
assign t[48589] = t[48588] ^ n[48589];
assign t[48590] = t[48589] ^ n[48590];
assign t[48591] = t[48590] ^ n[48591];
assign t[48592] = t[48591] ^ n[48592];
assign t[48593] = t[48592] ^ n[48593];
assign t[48594] = t[48593] ^ n[48594];
assign t[48595] = t[48594] ^ n[48595];
assign t[48596] = t[48595] ^ n[48596];
assign t[48597] = t[48596] ^ n[48597];
assign t[48598] = t[48597] ^ n[48598];
assign t[48599] = t[48598] ^ n[48599];
assign t[48600] = t[48599] ^ n[48600];
assign t[48601] = t[48600] ^ n[48601];
assign t[48602] = t[48601] ^ n[48602];
assign t[48603] = t[48602] ^ n[48603];
assign t[48604] = t[48603] ^ n[48604];
assign t[48605] = t[48604] ^ n[48605];
assign t[48606] = t[48605] ^ n[48606];
assign t[48607] = t[48606] ^ n[48607];
assign t[48608] = t[48607] ^ n[48608];
assign t[48609] = t[48608] ^ n[48609];
assign t[48610] = t[48609] ^ n[48610];
assign t[48611] = t[48610] ^ n[48611];
assign t[48612] = t[48611] ^ n[48612];
assign t[48613] = t[48612] ^ n[48613];
assign t[48614] = t[48613] ^ n[48614];
assign t[48615] = t[48614] ^ n[48615];
assign t[48616] = t[48615] ^ n[48616];
assign t[48617] = t[48616] ^ n[48617];
assign t[48618] = t[48617] ^ n[48618];
assign t[48619] = t[48618] ^ n[48619];
assign t[48620] = t[48619] ^ n[48620];
assign t[48621] = t[48620] ^ n[48621];
assign t[48622] = t[48621] ^ n[48622];
assign t[48623] = t[48622] ^ n[48623];
assign t[48624] = t[48623] ^ n[48624];
assign t[48625] = t[48624] ^ n[48625];
assign t[48626] = t[48625] ^ n[48626];
assign t[48627] = t[48626] ^ n[48627];
assign t[48628] = t[48627] ^ n[48628];
assign t[48629] = t[48628] ^ n[48629];
assign t[48630] = t[48629] ^ n[48630];
assign t[48631] = t[48630] ^ n[48631];
assign t[48632] = t[48631] ^ n[48632];
assign t[48633] = t[48632] ^ n[48633];
assign t[48634] = t[48633] ^ n[48634];
assign t[48635] = t[48634] ^ n[48635];
assign t[48636] = t[48635] ^ n[48636];
assign t[48637] = t[48636] ^ n[48637];
assign t[48638] = t[48637] ^ n[48638];
assign t[48639] = t[48638] ^ n[48639];
assign t[48640] = t[48639] ^ n[48640];
assign t[48641] = t[48640] ^ n[48641];
assign t[48642] = t[48641] ^ n[48642];
assign t[48643] = t[48642] ^ n[48643];
assign t[48644] = t[48643] ^ n[48644];
assign t[48645] = t[48644] ^ n[48645];
assign t[48646] = t[48645] ^ n[48646];
assign t[48647] = t[48646] ^ n[48647];
assign t[48648] = t[48647] ^ n[48648];
assign t[48649] = t[48648] ^ n[48649];
assign t[48650] = t[48649] ^ n[48650];
assign t[48651] = t[48650] ^ n[48651];
assign t[48652] = t[48651] ^ n[48652];
assign t[48653] = t[48652] ^ n[48653];
assign t[48654] = t[48653] ^ n[48654];
assign t[48655] = t[48654] ^ n[48655];
assign t[48656] = t[48655] ^ n[48656];
assign t[48657] = t[48656] ^ n[48657];
assign t[48658] = t[48657] ^ n[48658];
assign t[48659] = t[48658] ^ n[48659];
assign t[48660] = t[48659] ^ n[48660];
assign t[48661] = t[48660] ^ n[48661];
assign t[48662] = t[48661] ^ n[48662];
assign t[48663] = t[48662] ^ n[48663];
assign t[48664] = t[48663] ^ n[48664];
assign t[48665] = t[48664] ^ n[48665];
assign t[48666] = t[48665] ^ n[48666];
assign t[48667] = t[48666] ^ n[48667];
assign t[48668] = t[48667] ^ n[48668];
assign t[48669] = t[48668] ^ n[48669];
assign t[48670] = t[48669] ^ n[48670];
assign t[48671] = t[48670] ^ n[48671];
assign t[48672] = t[48671] ^ n[48672];
assign t[48673] = t[48672] ^ n[48673];
assign t[48674] = t[48673] ^ n[48674];
assign t[48675] = t[48674] ^ n[48675];
assign t[48676] = t[48675] ^ n[48676];
assign t[48677] = t[48676] ^ n[48677];
assign t[48678] = t[48677] ^ n[48678];
assign t[48679] = t[48678] ^ n[48679];
assign t[48680] = t[48679] ^ n[48680];
assign t[48681] = t[48680] ^ n[48681];
assign t[48682] = t[48681] ^ n[48682];
assign t[48683] = t[48682] ^ n[48683];
assign t[48684] = t[48683] ^ n[48684];
assign t[48685] = t[48684] ^ n[48685];
assign t[48686] = t[48685] ^ n[48686];
assign t[48687] = t[48686] ^ n[48687];
assign t[48688] = t[48687] ^ n[48688];
assign t[48689] = t[48688] ^ n[48689];
assign t[48690] = t[48689] ^ n[48690];
assign t[48691] = t[48690] ^ n[48691];
assign t[48692] = t[48691] ^ n[48692];
assign t[48693] = t[48692] ^ n[48693];
assign t[48694] = t[48693] ^ n[48694];
assign t[48695] = t[48694] ^ n[48695];
assign t[48696] = t[48695] ^ n[48696];
assign t[48697] = t[48696] ^ n[48697];
assign t[48698] = t[48697] ^ n[48698];
assign t[48699] = t[48698] ^ n[48699];
assign t[48700] = t[48699] ^ n[48700];
assign t[48701] = t[48700] ^ n[48701];
assign t[48702] = t[48701] ^ n[48702];
assign t[48703] = t[48702] ^ n[48703];
assign t[48704] = t[48703] ^ n[48704];
assign t[48705] = t[48704] ^ n[48705];
assign t[48706] = t[48705] ^ n[48706];
assign t[48707] = t[48706] ^ n[48707];
assign t[48708] = t[48707] ^ n[48708];
assign t[48709] = t[48708] ^ n[48709];
assign t[48710] = t[48709] ^ n[48710];
assign t[48711] = t[48710] ^ n[48711];
assign t[48712] = t[48711] ^ n[48712];
assign t[48713] = t[48712] ^ n[48713];
assign t[48714] = t[48713] ^ n[48714];
assign t[48715] = t[48714] ^ n[48715];
assign t[48716] = t[48715] ^ n[48716];
assign t[48717] = t[48716] ^ n[48717];
assign t[48718] = t[48717] ^ n[48718];
assign t[48719] = t[48718] ^ n[48719];
assign t[48720] = t[48719] ^ n[48720];
assign t[48721] = t[48720] ^ n[48721];
assign t[48722] = t[48721] ^ n[48722];
assign t[48723] = t[48722] ^ n[48723];
assign t[48724] = t[48723] ^ n[48724];
assign t[48725] = t[48724] ^ n[48725];
assign t[48726] = t[48725] ^ n[48726];
assign t[48727] = t[48726] ^ n[48727];
assign t[48728] = t[48727] ^ n[48728];
assign t[48729] = t[48728] ^ n[48729];
assign t[48730] = t[48729] ^ n[48730];
assign t[48731] = t[48730] ^ n[48731];
assign t[48732] = t[48731] ^ n[48732];
assign t[48733] = t[48732] ^ n[48733];
assign t[48734] = t[48733] ^ n[48734];
assign t[48735] = t[48734] ^ n[48735];
assign t[48736] = t[48735] ^ n[48736];
assign t[48737] = t[48736] ^ n[48737];
assign t[48738] = t[48737] ^ n[48738];
assign t[48739] = t[48738] ^ n[48739];
assign t[48740] = t[48739] ^ n[48740];
assign t[48741] = t[48740] ^ n[48741];
assign t[48742] = t[48741] ^ n[48742];
assign t[48743] = t[48742] ^ n[48743];
assign t[48744] = t[48743] ^ n[48744];
assign t[48745] = t[48744] ^ n[48745];
assign t[48746] = t[48745] ^ n[48746];
assign t[48747] = t[48746] ^ n[48747];
assign t[48748] = t[48747] ^ n[48748];
assign t[48749] = t[48748] ^ n[48749];
assign t[48750] = t[48749] ^ n[48750];
assign t[48751] = t[48750] ^ n[48751];
assign t[48752] = t[48751] ^ n[48752];
assign t[48753] = t[48752] ^ n[48753];
assign t[48754] = t[48753] ^ n[48754];
assign t[48755] = t[48754] ^ n[48755];
assign t[48756] = t[48755] ^ n[48756];
assign t[48757] = t[48756] ^ n[48757];
assign t[48758] = t[48757] ^ n[48758];
assign t[48759] = t[48758] ^ n[48759];
assign t[48760] = t[48759] ^ n[48760];
assign t[48761] = t[48760] ^ n[48761];
assign t[48762] = t[48761] ^ n[48762];
assign t[48763] = t[48762] ^ n[48763];
assign t[48764] = t[48763] ^ n[48764];
assign t[48765] = t[48764] ^ n[48765];
assign t[48766] = t[48765] ^ n[48766];
assign t[48767] = t[48766] ^ n[48767];
assign t[48768] = t[48767] ^ n[48768];
assign t[48769] = t[48768] ^ n[48769];
assign t[48770] = t[48769] ^ n[48770];
assign t[48771] = t[48770] ^ n[48771];
assign t[48772] = t[48771] ^ n[48772];
assign t[48773] = t[48772] ^ n[48773];
assign t[48774] = t[48773] ^ n[48774];
assign t[48775] = t[48774] ^ n[48775];
assign t[48776] = t[48775] ^ n[48776];
assign t[48777] = t[48776] ^ n[48777];
assign t[48778] = t[48777] ^ n[48778];
assign t[48779] = t[48778] ^ n[48779];
assign t[48780] = t[48779] ^ n[48780];
assign t[48781] = t[48780] ^ n[48781];
assign t[48782] = t[48781] ^ n[48782];
assign t[48783] = t[48782] ^ n[48783];
assign t[48784] = t[48783] ^ n[48784];
assign t[48785] = t[48784] ^ n[48785];
assign t[48786] = t[48785] ^ n[48786];
assign t[48787] = t[48786] ^ n[48787];
assign t[48788] = t[48787] ^ n[48788];
assign t[48789] = t[48788] ^ n[48789];
assign t[48790] = t[48789] ^ n[48790];
assign t[48791] = t[48790] ^ n[48791];
assign t[48792] = t[48791] ^ n[48792];
assign t[48793] = t[48792] ^ n[48793];
assign t[48794] = t[48793] ^ n[48794];
assign t[48795] = t[48794] ^ n[48795];
assign t[48796] = t[48795] ^ n[48796];
assign t[48797] = t[48796] ^ n[48797];
assign t[48798] = t[48797] ^ n[48798];
assign t[48799] = t[48798] ^ n[48799];
assign t[48800] = t[48799] ^ n[48800];
assign t[48801] = t[48800] ^ n[48801];
assign t[48802] = t[48801] ^ n[48802];
assign t[48803] = t[48802] ^ n[48803];
assign t[48804] = t[48803] ^ n[48804];
assign t[48805] = t[48804] ^ n[48805];
assign t[48806] = t[48805] ^ n[48806];
assign t[48807] = t[48806] ^ n[48807];
assign t[48808] = t[48807] ^ n[48808];
assign t[48809] = t[48808] ^ n[48809];
assign t[48810] = t[48809] ^ n[48810];
assign t[48811] = t[48810] ^ n[48811];
assign t[48812] = t[48811] ^ n[48812];
assign t[48813] = t[48812] ^ n[48813];
assign t[48814] = t[48813] ^ n[48814];
assign t[48815] = t[48814] ^ n[48815];
assign t[48816] = t[48815] ^ n[48816];
assign t[48817] = t[48816] ^ n[48817];
assign t[48818] = t[48817] ^ n[48818];
assign t[48819] = t[48818] ^ n[48819];
assign t[48820] = t[48819] ^ n[48820];
assign t[48821] = t[48820] ^ n[48821];
assign t[48822] = t[48821] ^ n[48822];
assign t[48823] = t[48822] ^ n[48823];
assign t[48824] = t[48823] ^ n[48824];
assign t[48825] = t[48824] ^ n[48825];
assign t[48826] = t[48825] ^ n[48826];
assign t[48827] = t[48826] ^ n[48827];
assign t[48828] = t[48827] ^ n[48828];
assign t[48829] = t[48828] ^ n[48829];
assign t[48830] = t[48829] ^ n[48830];
assign t[48831] = t[48830] ^ n[48831];
assign t[48832] = t[48831] ^ n[48832];
assign t[48833] = t[48832] ^ n[48833];
assign t[48834] = t[48833] ^ n[48834];
assign t[48835] = t[48834] ^ n[48835];
assign t[48836] = t[48835] ^ n[48836];
assign t[48837] = t[48836] ^ n[48837];
assign t[48838] = t[48837] ^ n[48838];
assign t[48839] = t[48838] ^ n[48839];
assign t[48840] = t[48839] ^ n[48840];
assign t[48841] = t[48840] ^ n[48841];
assign t[48842] = t[48841] ^ n[48842];
assign t[48843] = t[48842] ^ n[48843];
assign t[48844] = t[48843] ^ n[48844];
assign t[48845] = t[48844] ^ n[48845];
assign t[48846] = t[48845] ^ n[48846];
assign t[48847] = t[48846] ^ n[48847];
assign t[48848] = t[48847] ^ n[48848];
assign t[48849] = t[48848] ^ n[48849];
assign t[48850] = t[48849] ^ n[48850];
assign t[48851] = t[48850] ^ n[48851];
assign t[48852] = t[48851] ^ n[48852];
assign t[48853] = t[48852] ^ n[48853];
assign t[48854] = t[48853] ^ n[48854];
assign t[48855] = t[48854] ^ n[48855];
assign t[48856] = t[48855] ^ n[48856];
assign t[48857] = t[48856] ^ n[48857];
assign t[48858] = t[48857] ^ n[48858];
assign t[48859] = t[48858] ^ n[48859];
assign t[48860] = t[48859] ^ n[48860];
assign t[48861] = t[48860] ^ n[48861];
assign t[48862] = t[48861] ^ n[48862];
assign t[48863] = t[48862] ^ n[48863];
assign t[48864] = t[48863] ^ n[48864];
assign t[48865] = t[48864] ^ n[48865];
assign t[48866] = t[48865] ^ n[48866];
assign t[48867] = t[48866] ^ n[48867];
assign t[48868] = t[48867] ^ n[48868];
assign t[48869] = t[48868] ^ n[48869];
assign t[48870] = t[48869] ^ n[48870];
assign t[48871] = t[48870] ^ n[48871];
assign t[48872] = t[48871] ^ n[48872];
assign t[48873] = t[48872] ^ n[48873];
assign t[48874] = t[48873] ^ n[48874];
assign t[48875] = t[48874] ^ n[48875];
assign t[48876] = t[48875] ^ n[48876];
assign t[48877] = t[48876] ^ n[48877];
assign t[48878] = t[48877] ^ n[48878];
assign t[48879] = t[48878] ^ n[48879];
assign t[48880] = t[48879] ^ n[48880];
assign t[48881] = t[48880] ^ n[48881];
assign t[48882] = t[48881] ^ n[48882];
assign t[48883] = t[48882] ^ n[48883];
assign t[48884] = t[48883] ^ n[48884];
assign t[48885] = t[48884] ^ n[48885];
assign t[48886] = t[48885] ^ n[48886];
assign t[48887] = t[48886] ^ n[48887];
assign t[48888] = t[48887] ^ n[48888];
assign t[48889] = t[48888] ^ n[48889];
assign t[48890] = t[48889] ^ n[48890];
assign t[48891] = t[48890] ^ n[48891];
assign t[48892] = t[48891] ^ n[48892];
assign t[48893] = t[48892] ^ n[48893];
assign t[48894] = t[48893] ^ n[48894];
assign t[48895] = t[48894] ^ n[48895];
assign t[48896] = t[48895] ^ n[48896];
assign t[48897] = t[48896] ^ n[48897];
assign t[48898] = t[48897] ^ n[48898];
assign t[48899] = t[48898] ^ n[48899];
assign t[48900] = t[48899] ^ n[48900];
assign t[48901] = t[48900] ^ n[48901];
assign t[48902] = t[48901] ^ n[48902];
assign t[48903] = t[48902] ^ n[48903];
assign t[48904] = t[48903] ^ n[48904];
assign t[48905] = t[48904] ^ n[48905];
assign t[48906] = t[48905] ^ n[48906];
assign t[48907] = t[48906] ^ n[48907];
assign t[48908] = t[48907] ^ n[48908];
assign t[48909] = t[48908] ^ n[48909];
assign t[48910] = t[48909] ^ n[48910];
assign t[48911] = t[48910] ^ n[48911];
assign t[48912] = t[48911] ^ n[48912];
assign t[48913] = t[48912] ^ n[48913];
assign t[48914] = t[48913] ^ n[48914];
assign t[48915] = t[48914] ^ n[48915];
assign t[48916] = t[48915] ^ n[48916];
assign t[48917] = t[48916] ^ n[48917];
assign t[48918] = t[48917] ^ n[48918];
assign t[48919] = t[48918] ^ n[48919];
assign t[48920] = t[48919] ^ n[48920];
assign t[48921] = t[48920] ^ n[48921];
assign t[48922] = t[48921] ^ n[48922];
assign t[48923] = t[48922] ^ n[48923];
assign t[48924] = t[48923] ^ n[48924];
assign t[48925] = t[48924] ^ n[48925];
assign t[48926] = t[48925] ^ n[48926];
assign t[48927] = t[48926] ^ n[48927];
assign t[48928] = t[48927] ^ n[48928];
assign t[48929] = t[48928] ^ n[48929];
assign t[48930] = t[48929] ^ n[48930];
assign t[48931] = t[48930] ^ n[48931];
assign t[48932] = t[48931] ^ n[48932];
assign t[48933] = t[48932] ^ n[48933];
assign t[48934] = t[48933] ^ n[48934];
assign t[48935] = t[48934] ^ n[48935];
assign t[48936] = t[48935] ^ n[48936];
assign t[48937] = t[48936] ^ n[48937];
assign t[48938] = t[48937] ^ n[48938];
assign t[48939] = t[48938] ^ n[48939];
assign t[48940] = t[48939] ^ n[48940];
assign t[48941] = t[48940] ^ n[48941];
assign t[48942] = t[48941] ^ n[48942];
assign t[48943] = t[48942] ^ n[48943];
assign t[48944] = t[48943] ^ n[48944];
assign t[48945] = t[48944] ^ n[48945];
assign t[48946] = t[48945] ^ n[48946];
assign t[48947] = t[48946] ^ n[48947];
assign t[48948] = t[48947] ^ n[48948];
assign t[48949] = t[48948] ^ n[48949];
assign t[48950] = t[48949] ^ n[48950];
assign t[48951] = t[48950] ^ n[48951];
assign t[48952] = t[48951] ^ n[48952];
assign t[48953] = t[48952] ^ n[48953];
assign t[48954] = t[48953] ^ n[48954];
assign t[48955] = t[48954] ^ n[48955];
assign t[48956] = t[48955] ^ n[48956];
assign t[48957] = t[48956] ^ n[48957];
assign t[48958] = t[48957] ^ n[48958];
assign t[48959] = t[48958] ^ n[48959];
assign t[48960] = t[48959] ^ n[48960];
assign t[48961] = t[48960] ^ n[48961];
assign t[48962] = t[48961] ^ n[48962];
assign t[48963] = t[48962] ^ n[48963];
assign t[48964] = t[48963] ^ n[48964];
assign t[48965] = t[48964] ^ n[48965];
assign t[48966] = t[48965] ^ n[48966];
assign t[48967] = t[48966] ^ n[48967];
assign t[48968] = t[48967] ^ n[48968];
assign t[48969] = t[48968] ^ n[48969];
assign t[48970] = t[48969] ^ n[48970];
assign t[48971] = t[48970] ^ n[48971];
assign t[48972] = t[48971] ^ n[48972];
assign t[48973] = t[48972] ^ n[48973];
assign t[48974] = t[48973] ^ n[48974];
assign t[48975] = t[48974] ^ n[48975];
assign t[48976] = t[48975] ^ n[48976];
assign t[48977] = t[48976] ^ n[48977];
assign t[48978] = t[48977] ^ n[48978];
assign t[48979] = t[48978] ^ n[48979];
assign t[48980] = t[48979] ^ n[48980];
assign t[48981] = t[48980] ^ n[48981];
assign t[48982] = t[48981] ^ n[48982];
assign t[48983] = t[48982] ^ n[48983];
assign t[48984] = t[48983] ^ n[48984];
assign t[48985] = t[48984] ^ n[48985];
assign t[48986] = t[48985] ^ n[48986];
assign t[48987] = t[48986] ^ n[48987];
assign t[48988] = t[48987] ^ n[48988];
assign t[48989] = t[48988] ^ n[48989];
assign t[48990] = t[48989] ^ n[48990];
assign t[48991] = t[48990] ^ n[48991];
assign t[48992] = t[48991] ^ n[48992];
assign t[48993] = t[48992] ^ n[48993];
assign t[48994] = t[48993] ^ n[48994];
assign t[48995] = t[48994] ^ n[48995];
assign t[48996] = t[48995] ^ n[48996];
assign t[48997] = t[48996] ^ n[48997];
assign t[48998] = t[48997] ^ n[48998];
assign t[48999] = t[48998] ^ n[48999];
assign t[49000] = t[48999] ^ n[49000];
assign t[49001] = t[49000] ^ n[49001];
assign t[49002] = t[49001] ^ n[49002];
assign t[49003] = t[49002] ^ n[49003];
assign t[49004] = t[49003] ^ n[49004];
assign t[49005] = t[49004] ^ n[49005];
assign t[49006] = t[49005] ^ n[49006];
assign t[49007] = t[49006] ^ n[49007];
assign t[49008] = t[49007] ^ n[49008];
assign t[49009] = t[49008] ^ n[49009];
assign t[49010] = t[49009] ^ n[49010];
assign t[49011] = t[49010] ^ n[49011];
assign t[49012] = t[49011] ^ n[49012];
assign t[49013] = t[49012] ^ n[49013];
assign t[49014] = t[49013] ^ n[49014];
assign t[49015] = t[49014] ^ n[49015];
assign t[49016] = t[49015] ^ n[49016];
assign t[49017] = t[49016] ^ n[49017];
assign t[49018] = t[49017] ^ n[49018];
assign t[49019] = t[49018] ^ n[49019];
assign t[49020] = t[49019] ^ n[49020];
assign t[49021] = t[49020] ^ n[49021];
assign t[49022] = t[49021] ^ n[49022];
assign t[49023] = t[49022] ^ n[49023];
assign t[49024] = t[49023] ^ n[49024];
assign t[49025] = t[49024] ^ n[49025];
assign t[49026] = t[49025] ^ n[49026];
assign t[49027] = t[49026] ^ n[49027];
assign t[49028] = t[49027] ^ n[49028];
assign t[49029] = t[49028] ^ n[49029];
assign t[49030] = t[49029] ^ n[49030];
assign t[49031] = t[49030] ^ n[49031];
assign t[49032] = t[49031] ^ n[49032];
assign t[49033] = t[49032] ^ n[49033];
assign t[49034] = t[49033] ^ n[49034];
assign t[49035] = t[49034] ^ n[49035];
assign t[49036] = t[49035] ^ n[49036];
assign t[49037] = t[49036] ^ n[49037];
assign t[49038] = t[49037] ^ n[49038];
assign t[49039] = t[49038] ^ n[49039];
assign t[49040] = t[49039] ^ n[49040];
assign t[49041] = t[49040] ^ n[49041];
assign t[49042] = t[49041] ^ n[49042];
assign t[49043] = t[49042] ^ n[49043];
assign t[49044] = t[49043] ^ n[49044];
assign t[49045] = t[49044] ^ n[49045];
assign t[49046] = t[49045] ^ n[49046];
assign t[49047] = t[49046] ^ n[49047];
assign t[49048] = t[49047] ^ n[49048];
assign t[49049] = t[49048] ^ n[49049];
assign t[49050] = t[49049] ^ n[49050];
assign t[49051] = t[49050] ^ n[49051];
assign t[49052] = t[49051] ^ n[49052];
assign t[49053] = t[49052] ^ n[49053];
assign t[49054] = t[49053] ^ n[49054];
assign t[49055] = t[49054] ^ n[49055];
assign t[49056] = t[49055] ^ n[49056];
assign t[49057] = t[49056] ^ n[49057];
assign t[49058] = t[49057] ^ n[49058];
assign t[49059] = t[49058] ^ n[49059];
assign t[49060] = t[49059] ^ n[49060];
assign t[49061] = t[49060] ^ n[49061];
assign t[49062] = t[49061] ^ n[49062];
assign t[49063] = t[49062] ^ n[49063];
assign t[49064] = t[49063] ^ n[49064];
assign t[49065] = t[49064] ^ n[49065];
assign t[49066] = t[49065] ^ n[49066];
assign t[49067] = t[49066] ^ n[49067];
assign t[49068] = t[49067] ^ n[49068];
assign t[49069] = t[49068] ^ n[49069];
assign t[49070] = t[49069] ^ n[49070];
assign t[49071] = t[49070] ^ n[49071];
assign t[49072] = t[49071] ^ n[49072];
assign t[49073] = t[49072] ^ n[49073];
assign t[49074] = t[49073] ^ n[49074];
assign t[49075] = t[49074] ^ n[49075];
assign t[49076] = t[49075] ^ n[49076];
assign t[49077] = t[49076] ^ n[49077];
assign t[49078] = t[49077] ^ n[49078];
assign t[49079] = t[49078] ^ n[49079];
assign t[49080] = t[49079] ^ n[49080];
assign t[49081] = t[49080] ^ n[49081];
assign t[49082] = t[49081] ^ n[49082];
assign t[49083] = t[49082] ^ n[49083];
assign t[49084] = t[49083] ^ n[49084];
assign t[49085] = t[49084] ^ n[49085];
assign t[49086] = t[49085] ^ n[49086];
assign t[49087] = t[49086] ^ n[49087];
assign t[49088] = t[49087] ^ n[49088];
assign t[49089] = t[49088] ^ n[49089];
assign t[49090] = t[49089] ^ n[49090];
assign t[49091] = t[49090] ^ n[49091];
assign t[49092] = t[49091] ^ n[49092];
assign t[49093] = t[49092] ^ n[49093];
assign t[49094] = t[49093] ^ n[49094];
assign t[49095] = t[49094] ^ n[49095];
assign t[49096] = t[49095] ^ n[49096];
assign t[49097] = t[49096] ^ n[49097];
assign t[49098] = t[49097] ^ n[49098];
assign t[49099] = t[49098] ^ n[49099];
assign t[49100] = t[49099] ^ n[49100];
assign t[49101] = t[49100] ^ n[49101];
assign t[49102] = t[49101] ^ n[49102];
assign t[49103] = t[49102] ^ n[49103];
assign t[49104] = t[49103] ^ n[49104];
assign t[49105] = t[49104] ^ n[49105];
assign t[49106] = t[49105] ^ n[49106];
assign t[49107] = t[49106] ^ n[49107];
assign t[49108] = t[49107] ^ n[49108];
assign t[49109] = t[49108] ^ n[49109];
assign t[49110] = t[49109] ^ n[49110];
assign t[49111] = t[49110] ^ n[49111];
assign t[49112] = t[49111] ^ n[49112];
assign t[49113] = t[49112] ^ n[49113];
assign t[49114] = t[49113] ^ n[49114];
assign t[49115] = t[49114] ^ n[49115];
assign t[49116] = t[49115] ^ n[49116];
assign t[49117] = t[49116] ^ n[49117];
assign t[49118] = t[49117] ^ n[49118];
assign t[49119] = t[49118] ^ n[49119];
assign t[49120] = t[49119] ^ n[49120];
assign t[49121] = t[49120] ^ n[49121];
assign t[49122] = t[49121] ^ n[49122];
assign t[49123] = t[49122] ^ n[49123];
assign t[49124] = t[49123] ^ n[49124];
assign t[49125] = t[49124] ^ n[49125];
assign t[49126] = t[49125] ^ n[49126];
assign t[49127] = t[49126] ^ n[49127];
assign t[49128] = t[49127] ^ n[49128];
assign t[49129] = t[49128] ^ n[49129];
assign t[49130] = t[49129] ^ n[49130];
assign t[49131] = t[49130] ^ n[49131];
assign t[49132] = t[49131] ^ n[49132];
assign t[49133] = t[49132] ^ n[49133];
assign t[49134] = t[49133] ^ n[49134];
assign t[49135] = t[49134] ^ n[49135];
assign t[49136] = t[49135] ^ n[49136];
assign t[49137] = t[49136] ^ n[49137];
assign t[49138] = t[49137] ^ n[49138];
assign t[49139] = t[49138] ^ n[49139];
assign t[49140] = t[49139] ^ n[49140];
assign t[49141] = t[49140] ^ n[49141];
assign t[49142] = t[49141] ^ n[49142];
assign t[49143] = t[49142] ^ n[49143];
assign t[49144] = t[49143] ^ n[49144];
assign t[49145] = t[49144] ^ n[49145];
assign t[49146] = t[49145] ^ n[49146];
assign t[49147] = t[49146] ^ n[49147];
assign t[49148] = t[49147] ^ n[49148];
assign t[49149] = t[49148] ^ n[49149];
assign t[49150] = t[49149] ^ n[49150];
assign t[49151] = t[49150] ^ n[49151];
assign t[49152] = t[49151] ^ n[49152];
assign t[49153] = t[49152] ^ n[49153];
assign t[49154] = t[49153] ^ n[49154];
assign t[49155] = t[49154] ^ n[49155];
assign t[49156] = t[49155] ^ n[49156];
assign t[49157] = t[49156] ^ n[49157];
assign t[49158] = t[49157] ^ n[49158];
assign t[49159] = t[49158] ^ n[49159];
assign t[49160] = t[49159] ^ n[49160];
assign t[49161] = t[49160] ^ n[49161];
assign t[49162] = t[49161] ^ n[49162];
assign t[49163] = t[49162] ^ n[49163];
assign t[49164] = t[49163] ^ n[49164];
assign t[49165] = t[49164] ^ n[49165];
assign t[49166] = t[49165] ^ n[49166];
assign t[49167] = t[49166] ^ n[49167];
assign t[49168] = t[49167] ^ n[49168];
assign t[49169] = t[49168] ^ n[49169];
assign t[49170] = t[49169] ^ n[49170];
assign t[49171] = t[49170] ^ n[49171];
assign t[49172] = t[49171] ^ n[49172];
assign t[49173] = t[49172] ^ n[49173];
assign t[49174] = t[49173] ^ n[49174];
assign t[49175] = t[49174] ^ n[49175];
assign t[49176] = t[49175] ^ n[49176];
assign t[49177] = t[49176] ^ n[49177];
assign t[49178] = t[49177] ^ n[49178];
assign t[49179] = t[49178] ^ n[49179];
assign t[49180] = t[49179] ^ n[49180];
assign t[49181] = t[49180] ^ n[49181];
assign t[49182] = t[49181] ^ n[49182];
assign t[49183] = t[49182] ^ n[49183];
assign t[49184] = t[49183] ^ n[49184];
assign t[49185] = t[49184] ^ n[49185];
assign t[49186] = t[49185] ^ n[49186];
assign t[49187] = t[49186] ^ n[49187];
assign t[49188] = t[49187] ^ n[49188];
assign t[49189] = t[49188] ^ n[49189];
assign t[49190] = t[49189] ^ n[49190];
assign t[49191] = t[49190] ^ n[49191];
assign t[49192] = t[49191] ^ n[49192];
assign t[49193] = t[49192] ^ n[49193];
assign t[49194] = t[49193] ^ n[49194];
assign t[49195] = t[49194] ^ n[49195];
assign t[49196] = t[49195] ^ n[49196];
assign t[49197] = t[49196] ^ n[49197];
assign t[49198] = t[49197] ^ n[49198];
assign t[49199] = t[49198] ^ n[49199];
assign t[49200] = t[49199] ^ n[49200];
assign t[49201] = t[49200] ^ n[49201];
assign t[49202] = t[49201] ^ n[49202];
assign t[49203] = t[49202] ^ n[49203];
assign t[49204] = t[49203] ^ n[49204];
assign t[49205] = t[49204] ^ n[49205];
assign t[49206] = t[49205] ^ n[49206];
assign t[49207] = t[49206] ^ n[49207];
assign t[49208] = t[49207] ^ n[49208];
assign t[49209] = t[49208] ^ n[49209];
assign t[49210] = t[49209] ^ n[49210];
assign t[49211] = t[49210] ^ n[49211];
assign t[49212] = t[49211] ^ n[49212];
assign t[49213] = t[49212] ^ n[49213];
assign t[49214] = t[49213] ^ n[49214];
assign t[49215] = t[49214] ^ n[49215];
assign t[49216] = t[49215] ^ n[49216];
assign t[49217] = t[49216] ^ n[49217];
assign t[49218] = t[49217] ^ n[49218];
assign t[49219] = t[49218] ^ n[49219];
assign t[49220] = t[49219] ^ n[49220];
assign t[49221] = t[49220] ^ n[49221];
assign t[49222] = t[49221] ^ n[49222];
assign t[49223] = t[49222] ^ n[49223];
assign t[49224] = t[49223] ^ n[49224];
assign t[49225] = t[49224] ^ n[49225];
assign t[49226] = t[49225] ^ n[49226];
assign t[49227] = t[49226] ^ n[49227];
assign t[49228] = t[49227] ^ n[49228];
assign t[49229] = t[49228] ^ n[49229];
assign t[49230] = t[49229] ^ n[49230];
assign t[49231] = t[49230] ^ n[49231];
assign t[49232] = t[49231] ^ n[49232];
assign t[49233] = t[49232] ^ n[49233];
assign t[49234] = t[49233] ^ n[49234];
assign t[49235] = t[49234] ^ n[49235];
assign t[49236] = t[49235] ^ n[49236];
assign t[49237] = t[49236] ^ n[49237];
assign t[49238] = t[49237] ^ n[49238];
assign t[49239] = t[49238] ^ n[49239];
assign t[49240] = t[49239] ^ n[49240];
assign t[49241] = t[49240] ^ n[49241];
assign t[49242] = t[49241] ^ n[49242];
assign t[49243] = t[49242] ^ n[49243];
assign t[49244] = t[49243] ^ n[49244];
assign t[49245] = t[49244] ^ n[49245];
assign t[49246] = t[49245] ^ n[49246];
assign t[49247] = t[49246] ^ n[49247];
assign t[49248] = t[49247] ^ n[49248];
assign t[49249] = t[49248] ^ n[49249];
assign t[49250] = t[49249] ^ n[49250];
assign t[49251] = t[49250] ^ n[49251];
assign t[49252] = t[49251] ^ n[49252];
assign t[49253] = t[49252] ^ n[49253];
assign t[49254] = t[49253] ^ n[49254];
assign t[49255] = t[49254] ^ n[49255];
assign t[49256] = t[49255] ^ n[49256];
assign t[49257] = t[49256] ^ n[49257];
assign t[49258] = t[49257] ^ n[49258];
assign t[49259] = t[49258] ^ n[49259];
assign t[49260] = t[49259] ^ n[49260];
assign t[49261] = t[49260] ^ n[49261];
assign t[49262] = t[49261] ^ n[49262];
assign t[49263] = t[49262] ^ n[49263];
assign t[49264] = t[49263] ^ n[49264];
assign t[49265] = t[49264] ^ n[49265];
assign t[49266] = t[49265] ^ n[49266];
assign t[49267] = t[49266] ^ n[49267];
assign t[49268] = t[49267] ^ n[49268];
assign t[49269] = t[49268] ^ n[49269];
assign t[49270] = t[49269] ^ n[49270];
assign t[49271] = t[49270] ^ n[49271];
assign t[49272] = t[49271] ^ n[49272];
assign t[49273] = t[49272] ^ n[49273];
assign t[49274] = t[49273] ^ n[49274];
assign t[49275] = t[49274] ^ n[49275];
assign t[49276] = t[49275] ^ n[49276];
assign t[49277] = t[49276] ^ n[49277];
assign t[49278] = t[49277] ^ n[49278];
assign t[49279] = t[49278] ^ n[49279];
assign t[49280] = t[49279] ^ n[49280];
assign t[49281] = t[49280] ^ n[49281];
assign t[49282] = t[49281] ^ n[49282];
assign t[49283] = t[49282] ^ n[49283];
assign t[49284] = t[49283] ^ n[49284];
assign t[49285] = t[49284] ^ n[49285];
assign t[49286] = t[49285] ^ n[49286];
assign t[49287] = t[49286] ^ n[49287];
assign t[49288] = t[49287] ^ n[49288];
assign t[49289] = t[49288] ^ n[49289];
assign t[49290] = t[49289] ^ n[49290];
assign t[49291] = t[49290] ^ n[49291];
assign t[49292] = t[49291] ^ n[49292];
assign t[49293] = t[49292] ^ n[49293];
assign t[49294] = t[49293] ^ n[49294];
assign t[49295] = t[49294] ^ n[49295];
assign t[49296] = t[49295] ^ n[49296];
assign t[49297] = t[49296] ^ n[49297];
assign t[49298] = t[49297] ^ n[49298];
assign t[49299] = t[49298] ^ n[49299];
assign t[49300] = t[49299] ^ n[49300];
assign t[49301] = t[49300] ^ n[49301];
assign t[49302] = t[49301] ^ n[49302];
assign t[49303] = t[49302] ^ n[49303];
assign t[49304] = t[49303] ^ n[49304];
assign t[49305] = t[49304] ^ n[49305];
assign t[49306] = t[49305] ^ n[49306];
assign t[49307] = t[49306] ^ n[49307];
assign t[49308] = t[49307] ^ n[49308];
assign t[49309] = t[49308] ^ n[49309];
assign t[49310] = t[49309] ^ n[49310];
assign t[49311] = t[49310] ^ n[49311];
assign t[49312] = t[49311] ^ n[49312];
assign t[49313] = t[49312] ^ n[49313];
assign t[49314] = t[49313] ^ n[49314];
assign t[49315] = t[49314] ^ n[49315];
assign t[49316] = t[49315] ^ n[49316];
assign t[49317] = t[49316] ^ n[49317];
assign t[49318] = t[49317] ^ n[49318];
assign t[49319] = t[49318] ^ n[49319];
assign t[49320] = t[49319] ^ n[49320];
assign t[49321] = t[49320] ^ n[49321];
assign t[49322] = t[49321] ^ n[49322];
assign t[49323] = t[49322] ^ n[49323];
assign t[49324] = t[49323] ^ n[49324];
assign t[49325] = t[49324] ^ n[49325];
assign t[49326] = t[49325] ^ n[49326];
assign t[49327] = t[49326] ^ n[49327];
assign t[49328] = t[49327] ^ n[49328];
assign t[49329] = t[49328] ^ n[49329];
assign t[49330] = t[49329] ^ n[49330];
assign t[49331] = t[49330] ^ n[49331];
assign t[49332] = t[49331] ^ n[49332];
assign t[49333] = t[49332] ^ n[49333];
assign t[49334] = t[49333] ^ n[49334];
assign t[49335] = t[49334] ^ n[49335];
assign t[49336] = t[49335] ^ n[49336];
assign t[49337] = t[49336] ^ n[49337];
assign t[49338] = t[49337] ^ n[49338];
assign t[49339] = t[49338] ^ n[49339];
assign t[49340] = t[49339] ^ n[49340];
assign t[49341] = t[49340] ^ n[49341];
assign t[49342] = t[49341] ^ n[49342];
assign t[49343] = t[49342] ^ n[49343];
assign t[49344] = t[49343] ^ n[49344];
assign t[49345] = t[49344] ^ n[49345];
assign t[49346] = t[49345] ^ n[49346];
assign t[49347] = t[49346] ^ n[49347];
assign t[49348] = t[49347] ^ n[49348];
assign t[49349] = t[49348] ^ n[49349];
assign t[49350] = t[49349] ^ n[49350];
assign t[49351] = t[49350] ^ n[49351];
assign t[49352] = t[49351] ^ n[49352];
assign t[49353] = t[49352] ^ n[49353];
assign t[49354] = t[49353] ^ n[49354];
assign t[49355] = t[49354] ^ n[49355];
assign t[49356] = t[49355] ^ n[49356];
assign t[49357] = t[49356] ^ n[49357];
assign t[49358] = t[49357] ^ n[49358];
assign t[49359] = t[49358] ^ n[49359];
assign t[49360] = t[49359] ^ n[49360];
assign t[49361] = t[49360] ^ n[49361];
assign t[49362] = t[49361] ^ n[49362];
assign t[49363] = t[49362] ^ n[49363];
assign t[49364] = t[49363] ^ n[49364];
assign t[49365] = t[49364] ^ n[49365];
assign t[49366] = t[49365] ^ n[49366];
assign t[49367] = t[49366] ^ n[49367];
assign t[49368] = t[49367] ^ n[49368];
assign t[49369] = t[49368] ^ n[49369];
assign t[49370] = t[49369] ^ n[49370];
assign t[49371] = t[49370] ^ n[49371];
assign t[49372] = t[49371] ^ n[49372];
assign t[49373] = t[49372] ^ n[49373];
assign t[49374] = t[49373] ^ n[49374];
assign t[49375] = t[49374] ^ n[49375];
assign t[49376] = t[49375] ^ n[49376];
assign t[49377] = t[49376] ^ n[49377];
assign t[49378] = t[49377] ^ n[49378];
assign t[49379] = t[49378] ^ n[49379];
assign t[49380] = t[49379] ^ n[49380];
assign t[49381] = t[49380] ^ n[49381];
assign t[49382] = t[49381] ^ n[49382];
assign t[49383] = t[49382] ^ n[49383];
assign t[49384] = t[49383] ^ n[49384];
assign t[49385] = t[49384] ^ n[49385];
assign t[49386] = t[49385] ^ n[49386];
assign t[49387] = t[49386] ^ n[49387];
assign t[49388] = t[49387] ^ n[49388];
assign t[49389] = t[49388] ^ n[49389];
assign t[49390] = t[49389] ^ n[49390];
assign t[49391] = t[49390] ^ n[49391];
assign t[49392] = t[49391] ^ n[49392];
assign t[49393] = t[49392] ^ n[49393];
assign t[49394] = t[49393] ^ n[49394];
assign t[49395] = t[49394] ^ n[49395];
assign t[49396] = t[49395] ^ n[49396];
assign t[49397] = t[49396] ^ n[49397];
assign t[49398] = t[49397] ^ n[49398];
assign t[49399] = t[49398] ^ n[49399];
assign t[49400] = t[49399] ^ n[49400];
assign t[49401] = t[49400] ^ n[49401];
assign t[49402] = t[49401] ^ n[49402];
assign t[49403] = t[49402] ^ n[49403];
assign t[49404] = t[49403] ^ n[49404];
assign t[49405] = t[49404] ^ n[49405];
assign t[49406] = t[49405] ^ n[49406];
assign t[49407] = t[49406] ^ n[49407];
assign t[49408] = t[49407] ^ n[49408];
assign t[49409] = t[49408] ^ n[49409];
assign t[49410] = t[49409] ^ n[49410];
assign t[49411] = t[49410] ^ n[49411];
assign t[49412] = t[49411] ^ n[49412];
assign t[49413] = t[49412] ^ n[49413];
assign t[49414] = t[49413] ^ n[49414];
assign t[49415] = t[49414] ^ n[49415];
assign t[49416] = t[49415] ^ n[49416];
assign t[49417] = t[49416] ^ n[49417];
assign t[49418] = t[49417] ^ n[49418];
assign t[49419] = t[49418] ^ n[49419];
assign t[49420] = t[49419] ^ n[49420];
assign t[49421] = t[49420] ^ n[49421];
assign t[49422] = t[49421] ^ n[49422];
assign t[49423] = t[49422] ^ n[49423];
assign t[49424] = t[49423] ^ n[49424];
assign t[49425] = t[49424] ^ n[49425];
assign t[49426] = t[49425] ^ n[49426];
assign t[49427] = t[49426] ^ n[49427];
assign t[49428] = t[49427] ^ n[49428];
assign t[49429] = t[49428] ^ n[49429];
assign t[49430] = t[49429] ^ n[49430];
assign t[49431] = t[49430] ^ n[49431];
assign t[49432] = t[49431] ^ n[49432];
assign t[49433] = t[49432] ^ n[49433];
assign t[49434] = t[49433] ^ n[49434];
assign t[49435] = t[49434] ^ n[49435];
assign t[49436] = t[49435] ^ n[49436];
assign t[49437] = t[49436] ^ n[49437];
assign t[49438] = t[49437] ^ n[49438];
assign t[49439] = t[49438] ^ n[49439];
assign t[49440] = t[49439] ^ n[49440];
assign t[49441] = t[49440] ^ n[49441];
assign t[49442] = t[49441] ^ n[49442];
assign t[49443] = t[49442] ^ n[49443];
assign t[49444] = t[49443] ^ n[49444];
assign t[49445] = t[49444] ^ n[49445];
assign t[49446] = t[49445] ^ n[49446];
assign t[49447] = t[49446] ^ n[49447];
assign t[49448] = t[49447] ^ n[49448];
assign t[49449] = t[49448] ^ n[49449];
assign t[49450] = t[49449] ^ n[49450];
assign t[49451] = t[49450] ^ n[49451];
assign t[49452] = t[49451] ^ n[49452];
assign t[49453] = t[49452] ^ n[49453];
assign t[49454] = t[49453] ^ n[49454];
assign t[49455] = t[49454] ^ n[49455];
assign t[49456] = t[49455] ^ n[49456];
assign t[49457] = t[49456] ^ n[49457];
assign t[49458] = t[49457] ^ n[49458];
assign t[49459] = t[49458] ^ n[49459];
assign t[49460] = t[49459] ^ n[49460];
assign t[49461] = t[49460] ^ n[49461];
assign t[49462] = t[49461] ^ n[49462];
assign t[49463] = t[49462] ^ n[49463];
assign t[49464] = t[49463] ^ n[49464];
assign t[49465] = t[49464] ^ n[49465];
assign t[49466] = t[49465] ^ n[49466];
assign t[49467] = t[49466] ^ n[49467];
assign t[49468] = t[49467] ^ n[49468];
assign t[49469] = t[49468] ^ n[49469];
assign t[49470] = t[49469] ^ n[49470];
assign t[49471] = t[49470] ^ n[49471];
assign t[49472] = t[49471] ^ n[49472];
assign t[49473] = t[49472] ^ n[49473];
assign t[49474] = t[49473] ^ n[49474];
assign t[49475] = t[49474] ^ n[49475];
assign t[49476] = t[49475] ^ n[49476];
assign t[49477] = t[49476] ^ n[49477];
assign t[49478] = t[49477] ^ n[49478];
assign t[49479] = t[49478] ^ n[49479];
assign t[49480] = t[49479] ^ n[49480];
assign t[49481] = t[49480] ^ n[49481];
assign t[49482] = t[49481] ^ n[49482];
assign t[49483] = t[49482] ^ n[49483];
assign t[49484] = t[49483] ^ n[49484];
assign t[49485] = t[49484] ^ n[49485];
assign t[49486] = t[49485] ^ n[49486];
assign t[49487] = t[49486] ^ n[49487];
assign t[49488] = t[49487] ^ n[49488];
assign t[49489] = t[49488] ^ n[49489];
assign t[49490] = t[49489] ^ n[49490];
assign t[49491] = t[49490] ^ n[49491];
assign t[49492] = t[49491] ^ n[49492];
assign t[49493] = t[49492] ^ n[49493];
assign t[49494] = t[49493] ^ n[49494];
assign t[49495] = t[49494] ^ n[49495];
assign t[49496] = t[49495] ^ n[49496];
assign t[49497] = t[49496] ^ n[49497];
assign t[49498] = t[49497] ^ n[49498];
assign t[49499] = t[49498] ^ n[49499];
assign t[49500] = t[49499] ^ n[49500];
assign t[49501] = t[49500] ^ n[49501];
assign t[49502] = t[49501] ^ n[49502];
assign t[49503] = t[49502] ^ n[49503];
assign t[49504] = t[49503] ^ n[49504];
assign t[49505] = t[49504] ^ n[49505];
assign t[49506] = t[49505] ^ n[49506];
assign t[49507] = t[49506] ^ n[49507];
assign t[49508] = t[49507] ^ n[49508];
assign t[49509] = t[49508] ^ n[49509];
assign t[49510] = t[49509] ^ n[49510];
assign t[49511] = t[49510] ^ n[49511];
assign t[49512] = t[49511] ^ n[49512];
assign t[49513] = t[49512] ^ n[49513];
assign t[49514] = t[49513] ^ n[49514];
assign t[49515] = t[49514] ^ n[49515];
assign t[49516] = t[49515] ^ n[49516];
assign t[49517] = t[49516] ^ n[49517];
assign t[49518] = t[49517] ^ n[49518];
assign t[49519] = t[49518] ^ n[49519];
assign t[49520] = t[49519] ^ n[49520];
assign t[49521] = t[49520] ^ n[49521];
assign t[49522] = t[49521] ^ n[49522];
assign t[49523] = t[49522] ^ n[49523];
assign t[49524] = t[49523] ^ n[49524];
assign t[49525] = t[49524] ^ n[49525];
assign t[49526] = t[49525] ^ n[49526];
assign t[49527] = t[49526] ^ n[49527];
assign t[49528] = t[49527] ^ n[49528];
assign t[49529] = t[49528] ^ n[49529];
assign t[49530] = t[49529] ^ n[49530];
assign t[49531] = t[49530] ^ n[49531];
assign t[49532] = t[49531] ^ n[49532];
assign t[49533] = t[49532] ^ n[49533];
assign t[49534] = t[49533] ^ n[49534];
assign t[49535] = t[49534] ^ n[49535];
assign t[49536] = t[49535] ^ n[49536];
assign t[49537] = t[49536] ^ n[49537];
assign t[49538] = t[49537] ^ n[49538];
assign t[49539] = t[49538] ^ n[49539];
assign t[49540] = t[49539] ^ n[49540];
assign t[49541] = t[49540] ^ n[49541];
assign t[49542] = t[49541] ^ n[49542];
assign t[49543] = t[49542] ^ n[49543];
assign t[49544] = t[49543] ^ n[49544];
assign t[49545] = t[49544] ^ n[49545];
assign t[49546] = t[49545] ^ n[49546];
assign t[49547] = t[49546] ^ n[49547];
assign t[49548] = t[49547] ^ n[49548];
assign t[49549] = t[49548] ^ n[49549];
assign t[49550] = t[49549] ^ n[49550];
assign t[49551] = t[49550] ^ n[49551];
assign t[49552] = t[49551] ^ n[49552];
assign t[49553] = t[49552] ^ n[49553];
assign t[49554] = t[49553] ^ n[49554];
assign t[49555] = t[49554] ^ n[49555];
assign t[49556] = t[49555] ^ n[49556];
assign t[49557] = t[49556] ^ n[49557];
assign t[49558] = t[49557] ^ n[49558];
assign t[49559] = t[49558] ^ n[49559];
assign t[49560] = t[49559] ^ n[49560];
assign t[49561] = t[49560] ^ n[49561];
assign t[49562] = t[49561] ^ n[49562];
assign t[49563] = t[49562] ^ n[49563];
assign t[49564] = t[49563] ^ n[49564];
assign t[49565] = t[49564] ^ n[49565];
assign t[49566] = t[49565] ^ n[49566];
assign t[49567] = t[49566] ^ n[49567];
assign t[49568] = t[49567] ^ n[49568];
assign t[49569] = t[49568] ^ n[49569];
assign t[49570] = t[49569] ^ n[49570];
assign t[49571] = t[49570] ^ n[49571];
assign t[49572] = t[49571] ^ n[49572];
assign t[49573] = t[49572] ^ n[49573];
assign t[49574] = t[49573] ^ n[49574];
assign t[49575] = t[49574] ^ n[49575];
assign t[49576] = t[49575] ^ n[49576];
assign t[49577] = t[49576] ^ n[49577];
assign t[49578] = t[49577] ^ n[49578];
assign t[49579] = t[49578] ^ n[49579];
assign t[49580] = t[49579] ^ n[49580];
assign t[49581] = t[49580] ^ n[49581];
assign t[49582] = t[49581] ^ n[49582];
assign t[49583] = t[49582] ^ n[49583];
assign t[49584] = t[49583] ^ n[49584];
assign t[49585] = t[49584] ^ n[49585];
assign t[49586] = t[49585] ^ n[49586];
assign t[49587] = t[49586] ^ n[49587];
assign t[49588] = t[49587] ^ n[49588];
assign t[49589] = t[49588] ^ n[49589];
assign t[49590] = t[49589] ^ n[49590];
assign t[49591] = t[49590] ^ n[49591];
assign t[49592] = t[49591] ^ n[49592];
assign t[49593] = t[49592] ^ n[49593];
assign t[49594] = t[49593] ^ n[49594];
assign t[49595] = t[49594] ^ n[49595];
assign t[49596] = t[49595] ^ n[49596];
assign t[49597] = t[49596] ^ n[49597];
assign t[49598] = t[49597] ^ n[49598];
assign t[49599] = t[49598] ^ n[49599];
assign t[49600] = t[49599] ^ n[49600];
assign t[49601] = t[49600] ^ n[49601];
assign t[49602] = t[49601] ^ n[49602];
assign t[49603] = t[49602] ^ n[49603];
assign t[49604] = t[49603] ^ n[49604];
assign t[49605] = t[49604] ^ n[49605];
assign t[49606] = t[49605] ^ n[49606];
assign t[49607] = t[49606] ^ n[49607];
assign t[49608] = t[49607] ^ n[49608];
assign t[49609] = t[49608] ^ n[49609];
assign t[49610] = t[49609] ^ n[49610];
assign t[49611] = t[49610] ^ n[49611];
assign t[49612] = t[49611] ^ n[49612];
assign t[49613] = t[49612] ^ n[49613];
assign t[49614] = t[49613] ^ n[49614];
assign t[49615] = t[49614] ^ n[49615];
assign t[49616] = t[49615] ^ n[49616];
assign t[49617] = t[49616] ^ n[49617];
assign t[49618] = t[49617] ^ n[49618];
assign t[49619] = t[49618] ^ n[49619];
assign t[49620] = t[49619] ^ n[49620];
assign t[49621] = t[49620] ^ n[49621];
assign t[49622] = t[49621] ^ n[49622];
assign t[49623] = t[49622] ^ n[49623];
assign t[49624] = t[49623] ^ n[49624];
assign t[49625] = t[49624] ^ n[49625];
assign t[49626] = t[49625] ^ n[49626];
assign t[49627] = t[49626] ^ n[49627];
assign t[49628] = t[49627] ^ n[49628];
assign t[49629] = t[49628] ^ n[49629];
assign t[49630] = t[49629] ^ n[49630];
assign t[49631] = t[49630] ^ n[49631];
assign t[49632] = t[49631] ^ n[49632];
assign t[49633] = t[49632] ^ n[49633];
assign t[49634] = t[49633] ^ n[49634];
assign t[49635] = t[49634] ^ n[49635];
assign t[49636] = t[49635] ^ n[49636];
assign t[49637] = t[49636] ^ n[49637];
assign t[49638] = t[49637] ^ n[49638];
assign t[49639] = t[49638] ^ n[49639];
assign t[49640] = t[49639] ^ n[49640];
assign t[49641] = t[49640] ^ n[49641];
assign t[49642] = t[49641] ^ n[49642];
assign t[49643] = t[49642] ^ n[49643];
assign t[49644] = t[49643] ^ n[49644];
assign t[49645] = t[49644] ^ n[49645];
assign t[49646] = t[49645] ^ n[49646];
assign t[49647] = t[49646] ^ n[49647];
assign t[49648] = t[49647] ^ n[49648];
assign t[49649] = t[49648] ^ n[49649];
assign t[49650] = t[49649] ^ n[49650];
assign t[49651] = t[49650] ^ n[49651];
assign t[49652] = t[49651] ^ n[49652];
assign t[49653] = t[49652] ^ n[49653];
assign t[49654] = t[49653] ^ n[49654];
assign t[49655] = t[49654] ^ n[49655];
assign t[49656] = t[49655] ^ n[49656];
assign t[49657] = t[49656] ^ n[49657];
assign t[49658] = t[49657] ^ n[49658];
assign t[49659] = t[49658] ^ n[49659];
assign t[49660] = t[49659] ^ n[49660];
assign t[49661] = t[49660] ^ n[49661];
assign t[49662] = t[49661] ^ n[49662];
assign t[49663] = t[49662] ^ n[49663];
assign t[49664] = t[49663] ^ n[49664];
assign t[49665] = t[49664] ^ n[49665];
assign t[49666] = t[49665] ^ n[49666];
assign t[49667] = t[49666] ^ n[49667];
assign t[49668] = t[49667] ^ n[49668];
assign t[49669] = t[49668] ^ n[49669];
assign t[49670] = t[49669] ^ n[49670];
assign t[49671] = t[49670] ^ n[49671];
assign t[49672] = t[49671] ^ n[49672];
assign t[49673] = t[49672] ^ n[49673];
assign t[49674] = t[49673] ^ n[49674];
assign t[49675] = t[49674] ^ n[49675];
assign t[49676] = t[49675] ^ n[49676];
assign t[49677] = t[49676] ^ n[49677];
assign t[49678] = t[49677] ^ n[49678];
assign t[49679] = t[49678] ^ n[49679];
assign t[49680] = t[49679] ^ n[49680];
assign t[49681] = t[49680] ^ n[49681];
assign t[49682] = t[49681] ^ n[49682];
assign t[49683] = t[49682] ^ n[49683];
assign t[49684] = t[49683] ^ n[49684];
assign t[49685] = t[49684] ^ n[49685];
assign t[49686] = t[49685] ^ n[49686];
assign t[49687] = t[49686] ^ n[49687];
assign t[49688] = t[49687] ^ n[49688];
assign t[49689] = t[49688] ^ n[49689];
assign t[49690] = t[49689] ^ n[49690];
assign t[49691] = t[49690] ^ n[49691];
assign t[49692] = t[49691] ^ n[49692];
assign t[49693] = t[49692] ^ n[49693];
assign t[49694] = t[49693] ^ n[49694];
assign t[49695] = t[49694] ^ n[49695];
assign t[49696] = t[49695] ^ n[49696];
assign t[49697] = t[49696] ^ n[49697];
assign t[49698] = t[49697] ^ n[49698];
assign t[49699] = t[49698] ^ n[49699];
assign t[49700] = t[49699] ^ n[49700];
assign t[49701] = t[49700] ^ n[49701];
assign t[49702] = t[49701] ^ n[49702];
assign t[49703] = t[49702] ^ n[49703];
assign t[49704] = t[49703] ^ n[49704];
assign t[49705] = t[49704] ^ n[49705];
assign t[49706] = t[49705] ^ n[49706];
assign t[49707] = t[49706] ^ n[49707];
assign t[49708] = t[49707] ^ n[49708];
assign t[49709] = t[49708] ^ n[49709];
assign t[49710] = t[49709] ^ n[49710];
assign t[49711] = t[49710] ^ n[49711];
assign t[49712] = t[49711] ^ n[49712];
assign t[49713] = t[49712] ^ n[49713];
assign t[49714] = t[49713] ^ n[49714];
assign t[49715] = t[49714] ^ n[49715];
assign t[49716] = t[49715] ^ n[49716];
assign t[49717] = t[49716] ^ n[49717];
assign t[49718] = t[49717] ^ n[49718];
assign t[49719] = t[49718] ^ n[49719];
assign t[49720] = t[49719] ^ n[49720];
assign t[49721] = t[49720] ^ n[49721];
assign t[49722] = t[49721] ^ n[49722];
assign t[49723] = t[49722] ^ n[49723];
assign t[49724] = t[49723] ^ n[49724];
assign t[49725] = t[49724] ^ n[49725];
assign t[49726] = t[49725] ^ n[49726];
assign t[49727] = t[49726] ^ n[49727];
assign t[49728] = t[49727] ^ n[49728];
assign t[49729] = t[49728] ^ n[49729];
assign t[49730] = t[49729] ^ n[49730];
assign t[49731] = t[49730] ^ n[49731];
assign t[49732] = t[49731] ^ n[49732];
assign t[49733] = t[49732] ^ n[49733];
assign t[49734] = t[49733] ^ n[49734];
assign t[49735] = t[49734] ^ n[49735];
assign t[49736] = t[49735] ^ n[49736];
assign t[49737] = t[49736] ^ n[49737];
assign t[49738] = t[49737] ^ n[49738];
assign t[49739] = t[49738] ^ n[49739];
assign t[49740] = t[49739] ^ n[49740];
assign t[49741] = t[49740] ^ n[49741];
assign t[49742] = t[49741] ^ n[49742];
assign t[49743] = t[49742] ^ n[49743];
assign t[49744] = t[49743] ^ n[49744];
assign t[49745] = t[49744] ^ n[49745];
assign t[49746] = t[49745] ^ n[49746];
assign t[49747] = t[49746] ^ n[49747];
assign t[49748] = t[49747] ^ n[49748];
assign t[49749] = t[49748] ^ n[49749];
assign t[49750] = t[49749] ^ n[49750];
assign t[49751] = t[49750] ^ n[49751];
assign t[49752] = t[49751] ^ n[49752];
assign t[49753] = t[49752] ^ n[49753];
assign t[49754] = t[49753] ^ n[49754];
assign t[49755] = t[49754] ^ n[49755];
assign t[49756] = t[49755] ^ n[49756];
assign t[49757] = t[49756] ^ n[49757];
assign t[49758] = t[49757] ^ n[49758];
assign t[49759] = t[49758] ^ n[49759];
assign t[49760] = t[49759] ^ n[49760];
assign t[49761] = t[49760] ^ n[49761];
assign t[49762] = t[49761] ^ n[49762];
assign t[49763] = t[49762] ^ n[49763];
assign t[49764] = t[49763] ^ n[49764];
assign t[49765] = t[49764] ^ n[49765];
assign t[49766] = t[49765] ^ n[49766];
assign t[49767] = t[49766] ^ n[49767];
assign t[49768] = t[49767] ^ n[49768];
assign t[49769] = t[49768] ^ n[49769];
assign t[49770] = t[49769] ^ n[49770];
assign t[49771] = t[49770] ^ n[49771];
assign t[49772] = t[49771] ^ n[49772];
assign t[49773] = t[49772] ^ n[49773];
assign t[49774] = t[49773] ^ n[49774];
assign t[49775] = t[49774] ^ n[49775];
assign t[49776] = t[49775] ^ n[49776];
assign t[49777] = t[49776] ^ n[49777];
assign t[49778] = t[49777] ^ n[49778];
assign t[49779] = t[49778] ^ n[49779];
assign t[49780] = t[49779] ^ n[49780];
assign t[49781] = t[49780] ^ n[49781];
assign t[49782] = t[49781] ^ n[49782];
assign t[49783] = t[49782] ^ n[49783];
assign t[49784] = t[49783] ^ n[49784];
assign t[49785] = t[49784] ^ n[49785];
assign t[49786] = t[49785] ^ n[49786];
assign t[49787] = t[49786] ^ n[49787];
assign t[49788] = t[49787] ^ n[49788];
assign t[49789] = t[49788] ^ n[49789];
assign t[49790] = t[49789] ^ n[49790];
assign t[49791] = t[49790] ^ n[49791];
assign t[49792] = t[49791] ^ n[49792];
assign t[49793] = t[49792] ^ n[49793];
assign t[49794] = t[49793] ^ n[49794];
assign t[49795] = t[49794] ^ n[49795];
assign t[49796] = t[49795] ^ n[49796];
assign t[49797] = t[49796] ^ n[49797];
assign t[49798] = t[49797] ^ n[49798];
assign t[49799] = t[49798] ^ n[49799];
assign t[49800] = t[49799] ^ n[49800];
assign t[49801] = t[49800] ^ n[49801];
assign t[49802] = t[49801] ^ n[49802];
assign t[49803] = t[49802] ^ n[49803];
assign t[49804] = t[49803] ^ n[49804];
assign t[49805] = t[49804] ^ n[49805];
assign t[49806] = t[49805] ^ n[49806];
assign t[49807] = t[49806] ^ n[49807];
assign t[49808] = t[49807] ^ n[49808];
assign t[49809] = t[49808] ^ n[49809];
assign t[49810] = t[49809] ^ n[49810];
assign t[49811] = t[49810] ^ n[49811];
assign t[49812] = t[49811] ^ n[49812];
assign t[49813] = t[49812] ^ n[49813];
assign t[49814] = t[49813] ^ n[49814];
assign t[49815] = t[49814] ^ n[49815];
assign t[49816] = t[49815] ^ n[49816];
assign t[49817] = t[49816] ^ n[49817];
assign t[49818] = t[49817] ^ n[49818];
assign t[49819] = t[49818] ^ n[49819];
assign t[49820] = t[49819] ^ n[49820];
assign t[49821] = t[49820] ^ n[49821];
assign t[49822] = t[49821] ^ n[49822];
assign t[49823] = t[49822] ^ n[49823];
assign t[49824] = t[49823] ^ n[49824];
assign t[49825] = t[49824] ^ n[49825];
assign t[49826] = t[49825] ^ n[49826];
assign t[49827] = t[49826] ^ n[49827];
assign t[49828] = t[49827] ^ n[49828];
assign t[49829] = t[49828] ^ n[49829];
assign t[49830] = t[49829] ^ n[49830];
assign t[49831] = t[49830] ^ n[49831];
assign t[49832] = t[49831] ^ n[49832];
assign t[49833] = t[49832] ^ n[49833];
assign t[49834] = t[49833] ^ n[49834];
assign t[49835] = t[49834] ^ n[49835];
assign t[49836] = t[49835] ^ n[49836];
assign t[49837] = t[49836] ^ n[49837];
assign t[49838] = t[49837] ^ n[49838];
assign t[49839] = t[49838] ^ n[49839];
assign t[49840] = t[49839] ^ n[49840];
assign t[49841] = t[49840] ^ n[49841];
assign t[49842] = t[49841] ^ n[49842];
assign t[49843] = t[49842] ^ n[49843];
assign t[49844] = t[49843] ^ n[49844];
assign t[49845] = t[49844] ^ n[49845];
assign t[49846] = t[49845] ^ n[49846];
assign t[49847] = t[49846] ^ n[49847];
assign t[49848] = t[49847] ^ n[49848];
assign t[49849] = t[49848] ^ n[49849];
assign t[49850] = t[49849] ^ n[49850];
assign t[49851] = t[49850] ^ n[49851];
assign t[49852] = t[49851] ^ n[49852];
assign t[49853] = t[49852] ^ n[49853];
assign t[49854] = t[49853] ^ n[49854];
assign t[49855] = t[49854] ^ n[49855];
assign t[49856] = t[49855] ^ n[49856];
assign t[49857] = t[49856] ^ n[49857];
assign t[49858] = t[49857] ^ n[49858];
assign t[49859] = t[49858] ^ n[49859];
assign t[49860] = t[49859] ^ n[49860];
assign t[49861] = t[49860] ^ n[49861];
assign t[49862] = t[49861] ^ n[49862];
assign t[49863] = t[49862] ^ n[49863];
assign t[49864] = t[49863] ^ n[49864];
assign t[49865] = t[49864] ^ n[49865];
assign t[49866] = t[49865] ^ n[49866];
assign t[49867] = t[49866] ^ n[49867];
assign t[49868] = t[49867] ^ n[49868];
assign t[49869] = t[49868] ^ n[49869];
assign t[49870] = t[49869] ^ n[49870];
assign t[49871] = t[49870] ^ n[49871];
assign t[49872] = t[49871] ^ n[49872];
assign t[49873] = t[49872] ^ n[49873];
assign t[49874] = t[49873] ^ n[49874];
assign t[49875] = t[49874] ^ n[49875];
assign t[49876] = t[49875] ^ n[49876];
assign t[49877] = t[49876] ^ n[49877];
assign t[49878] = t[49877] ^ n[49878];
assign t[49879] = t[49878] ^ n[49879];
assign t[49880] = t[49879] ^ n[49880];
assign t[49881] = t[49880] ^ n[49881];
assign t[49882] = t[49881] ^ n[49882];
assign t[49883] = t[49882] ^ n[49883];
assign t[49884] = t[49883] ^ n[49884];
assign t[49885] = t[49884] ^ n[49885];
assign t[49886] = t[49885] ^ n[49886];
assign t[49887] = t[49886] ^ n[49887];
assign t[49888] = t[49887] ^ n[49888];
assign t[49889] = t[49888] ^ n[49889];
assign t[49890] = t[49889] ^ n[49890];
assign t[49891] = t[49890] ^ n[49891];
assign t[49892] = t[49891] ^ n[49892];
assign t[49893] = t[49892] ^ n[49893];
assign t[49894] = t[49893] ^ n[49894];
assign t[49895] = t[49894] ^ n[49895];
assign t[49896] = t[49895] ^ n[49896];
assign t[49897] = t[49896] ^ n[49897];
assign t[49898] = t[49897] ^ n[49898];
assign t[49899] = t[49898] ^ n[49899];
assign t[49900] = t[49899] ^ n[49900];
assign t[49901] = t[49900] ^ n[49901];
assign t[49902] = t[49901] ^ n[49902];
assign t[49903] = t[49902] ^ n[49903];
assign t[49904] = t[49903] ^ n[49904];
assign t[49905] = t[49904] ^ n[49905];
assign t[49906] = t[49905] ^ n[49906];
assign t[49907] = t[49906] ^ n[49907];
assign t[49908] = t[49907] ^ n[49908];
assign t[49909] = t[49908] ^ n[49909];
assign t[49910] = t[49909] ^ n[49910];
assign t[49911] = t[49910] ^ n[49911];
assign t[49912] = t[49911] ^ n[49912];
assign t[49913] = t[49912] ^ n[49913];
assign t[49914] = t[49913] ^ n[49914];
assign t[49915] = t[49914] ^ n[49915];
assign t[49916] = t[49915] ^ n[49916];
assign t[49917] = t[49916] ^ n[49917];
assign t[49918] = t[49917] ^ n[49918];
assign t[49919] = t[49918] ^ n[49919];
assign t[49920] = t[49919] ^ n[49920];
assign t[49921] = t[49920] ^ n[49921];
assign t[49922] = t[49921] ^ n[49922];
assign t[49923] = t[49922] ^ n[49923];
assign t[49924] = t[49923] ^ n[49924];
assign t[49925] = t[49924] ^ n[49925];
assign t[49926] = t[49925] ^ n[49926];
assign t[49927] = t[49926] ^ n[49927];
assign t[49928] = t[49927] ^ n[49928];
assign t[49929] = t[49928] ^ n[49929];
assign t[49930] = t[49929] ^ n[49930];
assign t[49931] = t[49930] ^ n[49931];
assign t[49932] = t[49931] ^ n[49932];
assign t[49933] = t[49932] ^ n[49933];
assign t[49934] = t[49933] ^ n[49934];
assign t[49935] = t[49934] ^ n[49935];
assign t[49936] = t[49935] ^ n[49936];
assign t[49937] = t[49936] ^ n[49937];
assign t[49938] = t[49937] ^ n[49938];
assign t[49939] = t[49938] ^ n[49939];
assign t[49940] = t[49939] ^ n[49940];
assign t[49941] = t[49940] ^ n[49941];
assign t[49942] = t[49941] ^ n[49942];
assign t[49943] = t[49942] ^ n[49943];
assign t[49944] = t[49943] ^ n[49944];
assign t[49945] = t[49944] ^ n[49945];
assign t[49946] = t[49945] ^ n[49946];
assign t[49947] = t[49946] ^ n[49947];
assign t[49948] = t[49947] ^ n[49948];
assign t[49949] = t[49948] ^ n[49949];
assign t[49950] = t[49949] ^ n[49950];
assign t[49951] = t[49950] ^ n[49951];
assign t[49952] = t[49951] ^ n[49952];
assign t[49953] = t[49952] ^ n[49953];
assign t[49954] = t[49953] ^ n[49954];
assign t[49955] = t[49954] ^ n[49955];
assign t[49956] = t[49955] ^ n[49956];
assign t[49957] = t[49956] ^ n[49957];
assign t[49958] = t[49957] ^ n[49958];
assign t[49959] = t[49958] ^ n[49959];
assign t[49960] = t[49959] ^ n[49960];
assign t[49961] = t[49960] ^ n[49961];
assign t[49962] = t[49961] ^ n[49962];
assign t[49963] = t[49962] ^ n[49963];
assign t[49964] = t[49963] ^ n[49964];
assign t[49965] = t[49964] ^ n[49965];
assign t[49966] = t[49965] ^ n[49966];
assign t[49967] = t[49966] ^ n[49967];
assign t[49968] = t[49967] ^ n[49968];
assign t[49969] = t[49968] ^ n[49969];
assign t[49970] = t[49969] ^ n[49970];
assign t[49971] = t[49970] ^ n[49971];
assign t[49972] = t[49971] ^ n[49972];
assign t[49973] = t[49972] ^ n[49973];
assign t[49974] = t[49973] ^ n[49974];
assign t[49975] = t[49974] ^ n[49975];
assign t[49976] = t[49975] ^ n[49976];
assign t[49977] = t[49976] ^ n[49977];
assign t[49978] = t[49977] ^ n[49978];
assign t[49979] = t[49978] ^ n[49979];
assign t[49980] = t[49979] ^ n[49980];
assign t[49981] = t[49980] ^ n[49981];
assign t[49982] = t[49981] ^ n[49982];
assign t[49983] = t[49982] ^ n[49983];
assign t[49984] = t[49983] ^ n[49984];
assign t[49985] = t[49984] ^ n[49985];
assign t[49986] = t[49985] ^ n[49986];
assign t[49987] = t[49986] ^ n[49987];
assign t[49988] = t[49987] ^ n[49988];
assign t[49989] = t[49988] ^ n[49989];
assign t[49990] = t[49989] ^ n[49990];
assign t[49991] = t[49990] ^ n[49991];
assign t[49992] = t[49991] ^ n[49992];
assign t[49993] = t[49992] ^ n[49993];
assign t[49994] = t[49993] ^ n[49994];
assign t[49995] = t[49994] ^ n[49995];
assign t[49996] = t[49995] ^ n[49996];
assign t[49997] = t[49996] ^ n[49997];
assign t[49998] = t[49997] ^ n[49998];
assign t[49999] = t[49998] ^ n[49999];
assign t[50000] = t[49999] ^ n[50000];
assign t[50001] = t[50000] ^ n[50001];
assign t[50002] = t[50001] ^ n[50002];
assign t[50003] = t[50002] ^ n[50003];
assign t[50004] = t[50003] ^ n[50004];
assign t[50005] = t[50004] ^ n[50005];
assign t[50006] = t[50005] ^ n[50006];
assign t[50007] = t[50006] ^ n[50007];
assign t[50008] = t[50007] ^ n[50008];
assign t[50009] = t[50008] ^ n[50009];
assign t[50010] = t[50009] ^ n[50010];
assign t[50011] = t[50010] ^ n[50011];
assign t[50012] = t[50011] ^ n[50012];
assign t[50013] = t[50012] ^ n[50013];
assign t[50014] = t[50013] ^ n[50014];
assign t[50015] = t[50014] ^ n[50015];
assign t[50016] = t[50015] ^ n[50016];
assign t[50017] = t[50016] ^ n[50017];
assign t[50018] = t[50017] ^ n[50018];
assign t[50019] = t[50018] ^ n[50019];
assign t[50020] = t[50019] ^ n[50020];
assign t[50021] = t[50020] ^ n[50021];
assign t[50022] = t[50021] ^ n[50022];
assign t[50023] = t[50022] ^ n[50023];
assign t[50024] = t[50023] ^ n[50024];
assign t[50025] = t[50024] ^ n[50025];
assign t[50026] = t[50025] ^ n[50026];
assign t[50027] = t[50026] ^ n[50027];
assign t[50028] = t[50027] ^ n[50028];
assign t[50029] = t[50028] ^ n[50029];
assign t[50030] = t[50029] ^ n[50030];
assign t[50031] = t[50030] ^ n[50031];
assign t[50032] = t[50031] ^ n[50032];
assign t[50033] = t[50032] ^ n[50033];
assign t[50034] = t[50033] ^ n[50034];
assign t[50035] = t[50034] ^ n[50035];
assign t[50036] = t[50035] ^ n[50036];
assign t[50037] = t[50036] ^ n[50037];
assign t[50038] = t[50037] ^ n[50038];
assign t[50039] = t[50038] ^ n[50039];
assign t[50040] = t[50039] ^ n[50040];
assign t[50041] = t[50040] ^ n[50041];
assign t[50042] = t[50041] ^ n[50042];
assign t[50043] = t[50042] ^ n[50043];
assign t[50044] = t[50043] ^ n[50044];
assign t[50045] = t[50044] ^ n[50045];
assign t[50046] = t[50045] ^ n[50046];
assign t[50047] = t[50046] ^ n[50047];
assign t[50048] = t[50047] ^ n[50048];
assign t[50049] = t[50048] ^ n[50049];
assign t[50050] = t[50049] ^ n[50050];
assign t[50051] = t[50050] ^ n[50051];
assign t[50052] = t[50051] ^ n[50052];
assign t[50053] = t[50052] ^ n[50053];
assign t[50054] = t[50053] ^ n[50054];
assign t[50055] = t[50054] ^ n[50055];
assign t[50056] = t[50055] ^ n[50056];
assign t[50057] = t[50056] ^ n[50057];
assign t[50058] = t[50057] ^ n[50058];
assign t[50059] = t[50058] ^ n[50059];
assign t[50060] = t[50059] ^ n[50060];
assign t[50061] = t[50060] ^ n[50061];
assign t[50062] = t[50061] ^ n[50062];
assign t[50063] = t[50062] ^ n[50063];
assign t[50064] = t[50063] ^ n[50064];
assign t[50065] = t[50064] ^ n[50065];
assign t[50066] = t[50065] ^ n[50066];
assign t[50067] = t[50066] ^ n[50067];
assign t[50068] = t[50067] ^ n[50068];
assign t[50069] = t[50068] ^ n[50069];
assign t[50070] = t[50069] ^ n[50070];
assign t[50071] = t[50070] ^ n[50071];
assign t[50072] = t[50071] ^ n[50072];
assign t[50073] = t[50072] ^ n[50073];
assign t[50074] = t[50073] ^ n[50074];
assign t[50075] = t[50074] ^ n[50075];
assign t[50076] = t[50075] ^ n[50076];
assign t[50077] = t[50076] ^ n[50077];
assign t[50078] = t[50077] ^ n[50078];
assign t[50079] = t[50078] ^ n[50079];
assign t[50080] = t[50079] ^ n[50080];
assign t[50081] = t[50080] ^ n[50081];
assign t[50082] = t[50081] ^ n[50082];
assign t[50083] = t[50082] ^ n[50083];
assign t[50084] = t[50083] ^ n[50084];
assign t[50085] = t[50084] ^ n[50085];
assign t[50086] = t[50085] ^ n[50086];
assign t[50087] = t[50086] ^ n[50087];
assign t[50088] = t[50087] ^ n[50088];
assign t[50089] = t[50088] ^ n[50089];
assign t[50090] = t[50089] ^ n[50090];
assign t[50091] = t[50090] ^ n[50091];
assign t[50092] = t[50091] ^ n[50092];
assign t[50093] = t[50092] ^ n[50093];
assign t[50094] = t[50093] ^ n[50094];
assign t[50095] = t[50094] ^ n[50095];
assign t[50096] = t[50095] ^ n[50096];
assign t[50097] = t[50096] ^ n[50097];
assign t[50098] = t[50097] ^ n[50098];
assign t[50099] = t[50098] ^ n[50099];
assign t[50100] = t[50099] ^ n[50100];
assign t[50101] = t[50100] ^ n[50101];
assign t[50102] = t[50101] ^ n[50102];
assign t[50103] = t[50102] ^ n[50103];
assign t[50104] = t[50103] ^ n[50104];
assign t[50105] = t[50104] ^ n[50105];
assign t[50106] = t[50105] ^ n[50106];
assign t[50107] = t[50106] ^ n[50107];
assign t[50108] = t[50107] ^ n[50108];
assign t[50109] = t[50108] ^ n[50109];
assign t[50110] = t[50109] ^ n[50110];
assign t[50111] = t[50110] ^ n[50111];
assign t[50112] = t[50111] ^ n[50112];
assign t[50113] = t[50112] ^ n[50113];
assign t[50114] = t[50113] ^ n[50114];
assign t[50115] = t[50114] ^ n[50115];
assign t[50116] = t[50115] ^ n[50116];
assign t[50117] = t[50116] ^ n[50117];
assign t[50118] = t[50117] ^ n[50118];
assign t[50119] = t[50118] ^ n[50119];
assign t[50120] = t[50119] ^ n[50120];
assign t[50121] = t[50120] ^ n[50121];
assign t[50122] = t[50121] ^ n[50122];
assign t[50123] = t[50122] ^ n[50123];
assign t[50124] = t[50123] ^ n[50124];
assign t[50125] = t[50124] ^ n[50125];
assign t[50126] = t[50125] ^ n[50126];
assign t[50127] = t[50126] ^ n[50127];
assign t[50128] = t[50127] ^ n[50128];
assign t[50129] = t[50128] ^ n[50129];
assign t[50130] = t[50129] ^ n[50130];
assign t[50131] = t[50130] ^ n[50131];
assign t[50132] = t[50131] ^ n[50132];
assign t[50133] = t[50132] ^ n[50133];
assign t[50134] = t[50133] ^ n[50134];
assign t[50135] = t[50134] ^ n[50135];
assign t[50136] = t[50135] ^ n[50136];
assign t[50137] = t[50136] ^ n[50137];
assign t[50138] = t[50137] ^ n[50138];
assign t[50139] = t[50138] ^ n[50139];
assign t[50140] = t[50139] ^ n[50140];
assign t[50141] = t[50140] ^ n[50141];
assign t[50142] = t[50141] ^ n[50142];
assign t[50143] = t[50142] ^ n[50143];
assign t[50144] = t[50143] ^ n[50144];
assign t[50145] = t[50144] ^ n[50145];
assign t[50146] = t[50145] ^ n[50146];
assign t[50147] = t[50146] ^ n[50147];
assign t[50148] = t[50147] ^ n[50148];
assign t[50149] = t[50148] ^ n[50149];
assign t[50150] = t[50149] ^ n[50150];
assign t[50151] = t[50150] ^ n[50151];
assign t[50152] = t[50151] ^ n[50152];
assign t[50153] = t[50152] ^ n[50153];
assign t[50154] = t[50153] ^ n[50154];
assign t[50155] = t[50154] ^ n[50155];
assign t[50156] = t[50155] ^ n[50156];
assign t[50157] = t[50156] ^ n[50157];
assign t[50158] = t[50157] ^ n[50158];
assign t[50159] = t[50158] ^ n[50159];
assign t[50160] = t[50159] ^ n[50160];
assign t[50161] = t[50160] ^ n[50161];
assign t[50162] = t[50161] ^ n[50162];
assign t[50163] = t[50162] ^ n[50163];
assign t[50164] = t[50163] ^ n[50164];
assign t[50165] = t[50164] ^ n[50165];
assign t[50166] = t[50165] ^ n[50166];
assign t[50167] = t[50166] ^ n[50167];
assign t[50168] = t[50167] ^ n[50168];
assign t[50169] = t[50168] ^ n[50169];
assign t[50170] = t[50169] ^ n[50170];
assign t[50171] = t[50170] ^ n[50171];
assign t[50172] = t[50171] ^ n[50172];
assign t[50173] = t[50172] ^ n[50173];
assign t[50174] = t[50173] ^ n[50174];
assign t[50175] = t[50174] ^ n[50175];
assign t[50176] = t[50175] ^ n[50176];
assign t[50177] = t[50176] ^ n[50177];
assign t[50178] = t[50177] ^ n[50178];
assign t[50179] = t[50178] ^ n[50179];
assign t[50180] = t[50179] ^ n[50180];
assign t[50181] = t[50180] ^ n[50181];
assign t[50182] = t[50181] ^ n[50182];
assign t[50183] = t[50182] ^ n[50183];
assign t[50184] = t[50183] ^ n[50184];
assign t[50185] = t[50184] ^ n[50185];
assign t[50186] = t[50185] ^ n[50186];
assign t[50187] = t[50186] ^ n[50187];
assign t[50188] = t[50187] ^ n[50188];
assign t[50189] = t[50188] ^ n[50189];
assign t[50190] = t[50189] ^ n[50190];
assign t[50191] = t[50190] ^ n[50191];
assign t[50192] = t[50191] ^ n[50192];
assign t[50193] = t[50192] ^ n[50193];
assign t[50194] = t[50193] ^ n[50194];
assign t[50195] = t[50194] ^ n[50195];
assign t[50196] = t[50195] ^ n[50196];
assign t[50197] = t[50196] ^ n[50197];
assign t[50198] = t[50197] ^ n[50198];
assign t[50199] = t[50198] ^ n[50199];
assign t[50200] = t[50199] ^ n[50200];
assign t[50201] = t[50200] ^ n[50201];
assign t[50202] = t[50201] ^ n[50202];
assign t[50203] = t[50202] ^ n[50203];
assign t[50204] = t[50203] ^ n[50204];
assign t[50205] = t[50204] ^ n[50205];
assign t[50206] = t[50205] ^ n[50206];
assign t[50207] = t[50206] ^ n[50207];
assign t[50208] = t[50207] ^ n[50208];
assign t[50209] = t[50208] ^ n[50209];
assign t[50210] = t[50209] ^ n[50210];
assign t[50211] = t[50210] ^ n[50211];
assign t[50212] = t[50211] ^ n[50212];
assign t[50213] = t[50212] ^ n[50213];
assign t[50214] = t[50213] ^ n[50214];
assign t[50215] = t[50214] ^ n[50215];
assign t[50216] = t[50215] ^ n[50216];
assign t[50217] = t[50216] ^ n[50217];
assign t[50218] = t[50217] ^ n[50218];
assign t[50219] = t[50218] ^ n[50219];
assign t[50220] = t[50219] ^ n[50220];
assign t[50221] = t[50220] ^ n[50221];
assign t[50222] = t[50221] ^ n[50222];
assign t[50223] = t[50222] ^ n[50223];
assign t[50224] = t[50223] ^ n[50224];
assign t[50225] = t[50224] ^ n[50225];
assign t[50226] = t[50225] ^ n[50226];
assign t[50227] = t[50226] ^ n[50227];
assign t[50228] = t[50227] ^ n[50228];
assign t[50229] = t[50228] ^ n[50229];
assign t[50230] = t[50229] ^ n[50230];
assign t[50231] = t[50230] ^ n[50231];
assign t[50232] = t[50231] ^ n[50232];
assign t[50233] = t[50232] ^ n[50233];
assign t[50234] = t[50233] ^ n[50234];
assign t[50235] = t[50234] ^ n[50235];
assign t[50236] = t[50235] ^ n[50236];
assign t[50237] = t[50236] ^ n[50237];
assign t[50238] = t[50237] ^ n[50238];
assign t[50239] = t[50238] ^ n[50239];
assign t[50240] = t[50239] ^ n[50240];
assign t[50241] = t[50240] ^ n[50241];
assign t[50242] = t[50241] ^ n[50242];
assign t[50243] = t[50242] ^ n[50243];
assign t[50244] = t[50243] ^ n[50244];
assign t[50245] = t[50244] ^ n[50245];
assign t[50246] = t[50245] ^ n[50246];
assign t[50247] = t[50246] ^ n[50247];
assign t[50248] = t[50247] ^ n[50248];
assign t[50249] = t[50248] ^ n[50249];
assign t[50250] = t[50249] ^ n[50250];
assign t[50251] = t[50250] ^ n[50251];
assign t[50252] = t[50251] ^ n[50252];
assign t[50253] = t[50252] ^ n[50253];
assign t[50254] = t[50253] ^ n[50254];
assign t[50255] = t[50254] ^ n[50255];
assign t[50256] = t[50255] ^ n[50256];
assign t[50257] = t[50256] ^ n[50257];
assign t[50258] = t[50257] ^ n[50258];
assign t[50259] = t[50258] ^ n[50259];
assign t[50260] = t[50259] ^ n[50260];
assign t[50261] = t[50260] ^ n[50261];
assign t[50262] = t[50261] ^ n[50262];
assign t[50263] = t[50262] ^ n[50263];
assign t[50264] = t[50263] ^ n[50264];
assign t[50265] = t[50264] ^ n[50265];
assign t[50266] = t[50265] ^ n[50266];
assign t[50267] = t[50266] ^ n[50267];
assign t[50268] = t[50267] ^ n[50268];
assign t[50269] = t[50268] ^ n[50269];
assign t[50270] = t[50269] ^ n[50270];
assign t[50271] = t[50270] ^ n[50271];
assign t[50272] = t[50271] ^ n[50272];
assign t[50273] = t[50272] ^ n[50273];
assign t[50274] = t[50273] ^ n[50274];
assign t[50275] = t[50274] ^ n[50275];
assign t[50276] = t[50275] ^ n[50276];
assign t[50277] = t[50276] ^ n[50277];
assign t[50278] = t[50277] ^ n[50278];
assign t[50279] = t[50278] ^ n[50279];
assign t[50280] = t[50279] ^ n[50280];
assign t[50281] = t[50280] ^ n[50281];
assign t[50282] = t[50281] ^ n[50282];
assign t[50283] = t[50282] ^ n[50283];
assign t[50284] = t[50283] ^ n[50284];
assign t[50285] = t[50284] ^ n[50285];
assign t[50286] = t[50285] ^ n[50286];
assign t[50287] = t[50286] ^ n[50287];
assign t[50288] = t[50287] ^ n[50288];
assign t[50289] = t[50288] ^ n[50289];
assign t[50290] = t[50289] ^ n[50290];
assign t[50291] = t[50290] ^ n[50291];
assign t[50292] = t[50291] ^ n[50292];
assign t[50293] = t[50292] ^ n[50293];
assign t[50294] = t[50293] ^ n[50294];
assign t[50295] = t[50294] ^ n[50295];
assign t[50296] = t[50295] ^ n[50296];
assign t[50297] = t[50296] ^ n[50297];
assign t[50298] = t[50297] ^ n[50298];
assign t[50299] = t[50298] ^ n[50299];
assign t[50300] = t[50299] ^ n[50300];
assign t[50301] = t[50300] ^ n[50301];
assign t[50302] = t[50301] ^ n[50302];
assign t[50303] = t[50302] ^ n[50303];
assign t[50304] = t[50303] ^ n[50304];
assign t[50305] = t[50304] ^ n[50305];
assign t[50306] = t[50305] ^ n[50306];
assign t[50307] = t[50306] ^ n[50307];
assign t[50308] = t[50307] ^ n[50308];
assign t[50309] = t[50308] ^ n[50309];
assign t[50310] = t[50309] ^ n[50310];
assign t[50311] = t[50310] ^ n[50311];
assign t[50312] = t[50311] ^ n[50312];
assign t[50313] = t[50312] ^ n[50313];
assign t[50314] = t[50313] ^ n[50314];
assign t[50315] = t[50314] ^ n[50315];
assign t[50316] = t[50315] ^ n[50316];
assign t[50317] = t[50316] ^ n[50317];
assign t[50318] = t[50317] ^ n[50318];
assign t[50319] = t[50318] ^ n[50319];
assign t[50320] = t[50319] ^ n[50320];
assign t[50321] = t[50320] ^ n[50321];
assign t[50322] = t[50321] ^ n[50322];
assign t[50323] = t[50322] ^ n[50323];
assign t[50324] = t[50323] ^ n[50324];
assign t[50325] = t[50324] ^ n[50325];
assign t[50326] = t[50325] ^ n[50326];
assign t[50327] = t[50326] ^ n[50327];
assign t[50328] = t[50327] ^ n[50328];
assign t[50329] = t[50328] ^ n[50329];
assign t[50330] = t[50329] ^ n[50330];
assign t[50331] = t[50330] ^ n[50331];
assign t[50332] = t[50331] ^ n[50332];
assign t[50333] = t[50332] ^ n[50333];
assign t[50334] = t[50333] ^ n[50334];
assign t[50335] = t[50334] ^ n[50335];
assign t[50336] = t[50335] ^ n[50336];
assign t[50337] = t[50336] ^ n[50337];
assign t[50338] = t[50337] ^ n[50338];
assign t[50339] = t[50338] ^ n[50339];
assign t[50340] = t[50339] ^ n[50340];
assign t[50341] = t[50340] ^ n[50341];
assign t[50342] = t[50341] ^ n[50342];
assign t[50343] = t[50342] ^ n[50343];
assign t[50344] = t[50343] ^ n[50344];
assign t[50345] = t[50344] ^ n[50345];
assign t[50346] = t[50345] ^ n[50346];
assign t[50347] = t[50346] ^ n[50347];
assign t[50348] = t[50347] ^ n[50348];
assign t[50349] = t[50348] ^ n[50349];
assign t[50350] = t[50349] ^ n[50350];
assign t[50351] = t[50350] ^ n[50351];
assign t[50352] = t[50351] ^ n[50352];
assign t[50353] = t[50352] ^ n[50353];
assign t[50354] = t[50353] ^ n[50354];
assign t[50355] = t[50354] ^ n[50355];
assign t[50356] = t[50355] ^ n[50356];
assign t[50357] = t[50356] ^ n[50357];
assign t[50358] = t[50357] ^ n[50358];
assign t[50359] = t[50358] ^ n[50359];
assign t[50360] = t[50359] ^ n[50360];
assign t[50361] = t[50360] ^ n[50361];
assign t[50362] = t[50361] ^ n[50362];
assign t[50363] = t[50362] ^ n[50363];
assign t[50364] = t[50363] ^ n[50364];
assign t[50365] = t[50364] ^ n[50365];
assign t[50366] = t[50365] ^ n[50366];
assign t[50367] = t[50366] ^ n[50367];
assign t[50368] = t[50367] ^ n[50368];
assign t[50369] = t[50368] ^ n[50369];
assign t[50370] = t[50369] ^ n[50370];
assign t[50371] = t[50370] ^ n[50371];
assign t[50372] = t[50371] ^ n[50372];
assign t[50373] = t[50372] ^ n[50373];
assign t[50374] = t[50373] ^ n[50374];
assign t[50375] = t[50374] ^ n[50375];
assign t[50376] = t[50375] ^ n[50376];
assign t[50377] = t[50376] ^ n[50377];
assign t[50378] = t[50377] ^ n[50378];
assign t[50379] = t[50378] ^ n[50379];
assign t[50380] = t[50379] ^ n[50380];
assign t[50381] = t[50380] ^ n[50381];
assign t[50382] = t[50381] ^ n[50382];
assign t[50383] = t[50382] ^ n[50383];
assign t[50384] = t[50383] ^ n[50384];
assign t[50385] = t[50384] ^ n[50385];
assign t[50386] = t[50385] ^ n[50386];
assign t[50387] = t[50386] ^ n[50387];
assign t[50388] = t[50387] ^ n[50388];
assign t[50389] = t[50388] ^ n[50389];
assign t[50390] = t[50389] ^ n[50390];
assign t[50391] = t[50390] ^ n[50391];
assign t[50392] = t[50391] ^ n[50392];
assign t[50393] = t[50392] ^ n[50393];
assign t[50394] = t[50393] ^ n[50394];
assign t[50395] = t[50394] ^ n[50395];
assign t[50396] = t[50395] ^ n[50396];
assign t[50397] = t[50396] ^ n[50397];
assign t[50398] = t[50397] ^ n[50398];
assign t[50399] = t[50398] ^ n[50399];
assign t[50400] = t[50399] ^ n[50400];
assign t[50401] = t[50400] ^ n[50401];
assign t[50402] = t[50401] ^ n[50402];
assign t[50403] = t[50402] ^ n[50403];
assign t[50404] = t[50403] ^ n[50404];
assign t[50405] = t[50404] ^ n[50405];
assign t[50406] = t[50405] ^ n[50406];
assign t[50407] = t[50406] ^ n[50407];
assign t[50408] = t[50407] ^ n[50408];
assign t[50409] = t[50408] ^ n[50409];
assign t[50410] = t[50409] ^ n[50410];
assign t[50411] = t[50410] ^ n[50411];
assign t[50412] = t[50411] ^ n[50412];
assign t[50413] = t[50412] ^ n[50413];
assign t[50414] = t[50413] ^ n[50414];
assign t[50415] = t[50414] ^ n[50415];
assign t[50416] = t[50415] ^ n[50416];
assign t[50417] = t[50416] ^ n[50417];
assign t[50418] = t[50417] ^ n[50418];
assign t[50419] = t[50418] ^ n[50419];
assign t[50420] = t[50419] ^ n[50420];
assign t[50421] = t[50420] ^ n[50421];
assign t[50422] = t[50421] ^ n[50422];
assign t[50423] = t[50422] ^ n[50423];
assign t[50424] = t[50423] ^ n[50424];
assign t[50425] = t[50424] ^ n[50425];
assign t[50426] = t[50425] ^ n[50426];
assign t[50427] = t[50426] ^ n[50427];
assign t[50428] = t[50427] ^ n[50428];
assign t[50429] = t[50428] ^ n[50429];
assign t[50430] = t[50429] ^ n[50430];
assign t[50431] = t[50430] ^ n[50431];
assign t[50432] = t[50431] ^ n[50432];
assign t[50433] = t[50432] ^ n[50433];
assign t[50434] = t[50433] ^ n[50434];
assign t[50435] = t[50434] ^ n[50435];
assign t[50436] = t[50435] ^ n[50436];
assign t[50437] = t[50436] ^ n[50437];
assign t[50438] = t[50437] ^ n[50438];
assign t[50439] = t[50438] ^ n[50439];
assign t[50440] = t[50439] ^ n[50440];
assign t[50441] = t[50440] ^ n[50441];
assign t[50442] = t[50441] ^ n[50442];
assign t[50443] = t[50442] ^ n[50443];
assign t[50444] = t[50443] ^ n[50444];
assign t[50445] = t[50444] ^ n[50445];
assign t[50446] = t[50445] ^ n[50446];
assign t[50447] = t[50446] ^ n[50447];
assign t[50448] = t[50447] ^ n[50448];
assign t[50449] = t[50448] ^ n[50449];
assign t[50450] = t[50449] ^ n[50450];
assign t[50451] = t[50450] ^ n[50451];
assign t[50452] = t[50451] ^ n[50452];
assign t[50453] = t[50452] ^ n[50453];
assign t[50454] = t[50453] ^ n[50454];
assign t[50455] = t[50454] ^ n[50455];
assign t[50456] = t[50455] ^ n[50456];
assign t[50457] = t[50456] ^ n[50457];
assign t[50458] = t[50457] ^ n[50458];
assign t[50459] = t[50458] ^ n[50459];
assign t[50460] = t[50459] ^ n[50460];
assign t[50461] = t[50460] ^ n[50461];
assign t[50462] = t[50461] ^ n[50462];
assign t[50463] = t[50462] ^ n[50463];
assign t[50464] = t[50463] ^ n[50464];
assign t[50465] = t[50464] ^ n[50465];
assign t[50466] = t[50465] ^ n[50466];
assign t[50467] = t[50466] ^ n[50467];
assign t[50468] = t[50467] ^ n[50468];
assign t[50469] = t[50468] ^ n[50469];
assign t[50470] = t[50469] ^ n[50470];
assign t[50471] = t[50470] ^ n[50471];
assign t[50472] = t[50471] ^ n[50472];
assign t[50473] = t[50472] ^ n[50473];
assign t[50474] = t[50473] ^ n[50474];
assign t[50475] = t[50474] ^ n[50475];
assign t[50476] = t[50475] ^ n[50476];
assign t[50477] = t[50476] ^ n[50477];
assign t[50478] = t[50477] ^ n[50478];
assign t[50479] = t[50478] ^ n[50479];
assign t[50480] = t[50479] ^ n[50480];
assign t[50481] = t[50480] ^ n[50481];
assign t[50482] = t[50481] ^ n[50482];
assign t[50483] = t[50482] ^ n[50483];
assign t[50484] = t[50483] ^ n[50484];
assign t[50485] = t[50484] ^ n[50485];
assign t[50486] = t[50485] ^ n[50486];
assign t[50487] = t[50486] ^ n[50487];
assign t[50488] = t[50487] ^ n[50488];
assign t[50489] = t[50488] ^ n[50489];
assign t[50490] = t[50489] ^ n[50490];
assign t[50491] = t[50490] ^ n[50491];
assign t[50492] = t[50491] ^ n[50492];
assign t[50493] = t[50492] ^ n[50493];
assign t[50494] = t[50493] ^ n[50494];
assign t[50495] = t[50494] ^ n[50495];
assign t[50496] = t[50495] ^ n[50496];
assign t[50497] = t[50496] ^ n[50497];
assign t[50498] = t[50497] ^ n[50498];
assign t[50499] = t[50498] ^ n[50499];
assign t[50500] = t[50499] ^ n[50500];
assign t[50501] = t[50500] ^ n[50501];
assign t[50502] = t[50501] ^ n[50502];
assign t[50503] = t[50502] ^ n[50503];
assign t[50504] = t[50503] ^ n[50504];
assign t[50505] = t[50504] ^ n[50505];
assign t[50506] = t[50505] ^ n[50506];
assign t[50507] = t[50506] ^ n[50507];
assign t[50508] = t[50507] ^ n[50508];
assign t[50509] = t[50508] ^ n[50509];
assign t[50510] = t[50509] ^ n[50510];
assign t[50511] = t[50510] ^ n[50511];
assign t[50512] = t[50511] ^ n[50512];
assign t[50513] = t[50512] ^ n[50513];
assign t[50514] = t[50513] ^ n[50514];
assign t[50515] = t[50514] ^ n[50515];
assign t[50516] = t[50515] ^ n[50516];
assign t[50517] = t[50516] ^ n[50517];
assign t[50518] = t[50517] ^ n[50518];
assign t[50519] = t[50518] ^ n[50519];
assign t[50520] = t[50519] ^ n[50520];
assign t[50521] = t[50520] ^ n[50521];
assign t[50522] = t[50521] ^ n[50522];
assign t[50523] = t[50522] ^ n[50523];
assign t[50524] = t[50523] ^ n[50524];
assign t[50525] = t[50524] ^ n[50525];
assign t[50526] = t[50525] ^ n[50526];
assign t[50527] = t[50526] ^ n[50527];
assign t[50528] = t[50527] ^ n[50528];
assign t[50529] = t[50528] ^ n[50529];
assign t[50530] = t[50529] ^ n[50530];
assign t[50531] = t[50530] ^ n[50531];
assign t[50532] = t[50531] ^ n[50532];
assign t[50533] = t[50532] ^ n[50533];
assign t[50534] = t[50533] ^ n[50534];
assign t[50535] = t[50534] ^ n[50535];
assign t[50536] = t[50535] ^ n[50536];
assign t[50537] = t[50536] ^ n[50537];
assign t[50538] = t[50537] ^ n[50538];
assign t[50539] = t[50538] ^ n[50539];
assign t[50540] = t[50539] ^ n[50540];
assign t[50541] = t[50540] ^ n[50541];
assign t[50542] = t[50541] ^ n[50542];
assign t[50543] = t[50542] ^ n[50543];
assign t[50544] = t[50543] ^ n[50544];
assign t[50545] = t[50544] ^ n[50545];
assign t[50546] = t[50545] ^ n[50546];
assign t[50547] = t[50546] ^ n[50547];
assign t[50548] = t[50547] ^ n[50548];
assign t[50549] = t[50548] ^ n[50549];
assign t[50550] = t[50549] ^ n[50550];
assign t[50551] = t[50550] ^ n[50551];
assign t[50552] = t[50551] ^ n[50552];
assign t[50553] = t[50552] ^ n[50553];
assign t[50554] = t[50553] ^ n[50554];
assign t[50555] = t[50554] ^ n[50555];
assign t[50556] = t[50555] ^ n[50556];
assign t[50557] = t[50556] ^ n[50557];
assign t[50558] = t[50557] ^ n[50558];
assign t[50559] = t[50558] ^ n[50559];
assign t[50560] = t[50559] ^ n[50560];
assign t[50561] = t[50560] ^ n[50561];
assign t[50562] = t[50561] ^ n[50562];
assign t[50563] = t[50562] ^ n[50563];
assign t[50564] = t[50563] ^ n[50564];
assign t[50565] = t[50564] ^ n[50565];
assign t[50566] = t[50565] ^ n[50566];
assign t[50567] = t[50566] ^ n[50567];
assign t[50568] = t[50567] ^ n[50568];
assign t[50569] = t[50568] ^ n[50569];
assign t[50570] = t[50569] ^ n[50570];
assign t[50571] = t[50570] ^ n[50571];
assign t[50572] = t[50571] ^ n[50572];
assign t[50573] = t[50572] ^ n[50573];
assign t[50574] = t[50573] ^ n[50574];
assign t[50575] = t[50574] ^ n[50575];
assign t[50576] = t[50575] ^ n[50576];
assign t[50577] = t[50576] ^ n[50577];
assign t[50578] = t[50577] ^ n[50578];
assign t[50579] = t[50578] ^ n[50579];
assign t[50580] = t[50579] ^ n[50580];
assign t[50581] = t[50580] ^ n[50581];
assign t[50582] = t[50581] ^ n[50582];
assign t[50583] = t[50582] ^ n[50583];
assign t[50584] = t[50583] ^ n[50584];
assign t[50585] = t[50584] ^ n[50585];
assign t[50586] = t[50585] ^ n[50586];
assign t[50587] = t[50586] ^ n[50587];
assign t[50588] = t[50587] ^ n[50588];
assign t[50589] = t[50588] ^ n[50589];
assign t[50590] = t[50589] ^ n[50590];
assign t[50591] = t[50590] ^ n[50591];
assign t[50592] = t[50591] ^ n[50592];
assign t[50593] = t[50592] ^ n[50593];
assign t[50594] = t[50593] ^ n[50594];
assign t[50595] = t[50594] ^ n[50595];
assign t[50596] = t[50595] ^ n[50596];
assign t[50597] = t[50596] ^ n[50597];
assign t[50598] = t[50597] ^ n[50598];
assign t[50599] = t[50598] ^ n[50599];
assign t[50600] = t[50599] ^ n[50600];
assign t[50601] = t[50600] ^ n[50601];
assign t[50602] = t[50601] ^ n[50602];
assign t[50603] = t[50602] ^ n[50603];
assign t[50604] = t[50603] ^ n[50604];
assign t[50605] = t[50604] ^ n[50605];
assign t[50606] = t[50605] ^ n[50606];
assign t[50607] = t[50606] ^ n[50607];
assign t[50608] = t[50607] ^ n[50608];
assign t[50609] = t[50608] ^ n[50609];
assign t[50610] = t[50609] ^ n[50610];
assign t[50611] = t[50610] ^ n[50611];
assign t[50612] = t[50611] ^ n[50612];
assign t[50613] = t[50612] ^ n[50613];
assign t[50614] = t[50613] ^ n[50614];
assign t[50615] = t[50614] ^ n[50615];
assign t[50616] = t[50615] ^ n[50616];
assign t[50617] = t[50616] ^ n[50617];
assign t[50618] = t[50617] ^ n[50618];
assign t[50619] = t[50618] ^ n[50619];
assign t[50620] = t[50619] ^ n[50620];
assign t[50621] = t[50620] ^ n[50621];
assign t[50622] = t[50621] ^ n[50622];
assign t[50623] = t[50622] ^ n[50623];
assign t[50624] = t[50623] ^ n[50624];
assign t[50625] = t[50624] ^ n[50625];
assign t[50626] = t[50625] ^ n[50626];
assign t[50627] = t[50626] ^ n[50627];
assign t[50628] = t[50627] ^ n[50628];
assign t[50629] = t[50628] ^ n[50629];
assign t[50630] = t[50629] ^ n[50630];
assign t[50631] = t[50630] ^ n[50631];
assign t[50632] = t[50631] ^ n[50632];
assign t[50633] = t[50632] ^ n[50633];
assign t[50634] = t[50633] ^ n[50634];
assign t[50635] = t[50634] ^ n[50635];
assign t[50636] = t[50635] ^ n[50636];
assign t[50637] = t[50636] ^ n[50637];
assign t[50638] = t[50637] ^ n[50638];
assign t[50639] = t[50638] ^ n[50639];
assign t[50640] = t[50639] ^ n[50640];
assign t[50641] = t[50640] ^ n[50641];
assign t[50642] = t[50641] ^ n[50642];
assign t[50643] = t[50642] ^ n[50643];
assign t[50644] = t[50643] ^ n[50644];
assign t[50645] = t[50644] ^ n[50645];
assign t[50646] = t[50645] ^ n[50646];
assign t[50647] = t[50646] ^ n[50647];
assign t[50648] = t[50647] ^ n[50648];
assign t[50649] = t[50648] ^ n[50649];
assign t[50650] = t[50649] ^ n[50650];
assign t[50651] = t[50650] ^ n[50651];
assign t[50652] = t[50651] ^ n[50652];
assign t[50653] = t[50652] ^ n[50653];
assign t[50654] = t[50653] ^ n[50654];
assign t[50655] = t[50654] ^ n[50655];
assign t[50656] = t[50655] ^ n[50656];
assign t[50657] = t[50656] ^ n[50657];
assign t[50658] = t[50657] ^ n[50658];
assign t[50659] = t[50658] ^ n[50659];
assign t[50660] = t[50659] ^ n[50660];
assign t[50661] = t[50660] ^ n[50661];
assign t[50662] = t[50661] ^ n[50662];
assign t[50663] = t[50662] ^ n[50663];
assign t[50664] = t[50663] ^ n[50664];
assign t[50665] = t[50664] ^ n[50665];
assign t[50666] = t[50665] ^ n[50666];
assign t[50667] = t[50666] ^ n[50667];
assign t[50668] = t[50667] ^ n[50668];
assign t[50669] = t[50668] ^ n[50669];
assign t[50670] = t[50669] ^ n[50670];
assign t[50671] = t[50670] ^ n[50671];
assign t[50672] = t[50671] ^ n[50672];
assign t[50673] = t[50672] ^ n[50673];
assign t[50674] = t[50673] ^ n[50674];
assign t[50675] = t[50674] ^ n[50675];
assign t[50676] = t[50675] ^ n[50676];
assign t[50677] = t[50676] ^ n[50677];
assign t[50678] = t[50677] ^ n[50678];
assign t[50679] = t[50678] ^ n[50679];
assign t[50680] = t[50679] ^ n[50680];
assign t[50681] = t[50680] ^ n[50681];
assign t[50682] = t[50681] ^ n[50682];
assign t[50683] = t[50682] ^ n[50683];
assign t[50684] = t[50683] ^ n[50684];
assign t[50685] = t[50684] ^ n[50685];
assign t[50686] = t[50685] ^ n[50686];
assign t[50687] = t[50686] ^ n[50687];
assign t[50688] = t[50687] ^ n[50688];
assign t[50689] = t[50688] ^ n[50689];
assign t[50690] = t[50689] ^ n[50690];
assign t[50691] = t[50690] ^ n[50691];
assign t[50692] = t[50691] ^ n[50692];
assign t[50693] = t[50692] ^ n[50693];
assign t[50694] = t[50693] ^ n[50694];
assign t[50695] = t[50694] ^ n[50695];
assign t[50696] = t[50695] ^ n[50696];
assign t[50697] = t[50696] ^ n[50697];
assign t[50698] = t[50697] ^ n[50698];
assign t[50699] = t[50698] ^ n[50699];
assign t[50700] = t[50699] ^ n[50700];
assign t[50701] = t[50700] ^ n[50701];
assign t[50702] = t[50701] ^ n[50702];
assign t[50703] = t[50702] ^ n[50703];
assign t[50704] = t[50703] ^ n[50704];
assign t[50705] = t[50704] ^ n[50705];
assign t[50706] = t[50705] ^ n[50706];
assign t[50707] = t[50706] ^ n[50707];
assign t[50708] = t[50707] ^ n[50708];
assign t[50709] = t[50708] ^ n[50709];
assign t[50710] = t[50709] ^ n[50710];
assign t[50711] = t[50710] ^ n[50711];
assign t[50712] = t[50711] ^ n[50712];
assign t[50713] = t[50712] ^ n[50713];
assign t[50714] = t[50713] ^ n[50714];
assign t[50715] = t[50714] ^ n[50715];
assign t[50716] = t[50715] ^ n[50716];
assign t[50717] = t[50716] ^ n[50717];
assign t[50718] = t[50717] ^ n[50718];
assign t[50719] = t[50718] ^ n[50719];
assign t[50720] = t[50719] ^ n[50720];
assign t[50721] = t[50720] ^ n[50721];
assign t[50722] = t[50721] ^ n[50722];
assign t[50723] = t[50722] ^ n[50723];
assign t[50724] = t[50723] ^ n[50724];
assign t[50725] = t[50724] ^ n[50725];
assign t[50726] = t[50725] ^ n[50726];
assign t[50727] = t[50726] ^ n[50727];
assign t[50728] = t[50727] ^ n[50728];
assign t[50729] = t[50728] ^ n[50729];
assign t[50730] = t[50729] ^ n[50730];
assign t[50731] = t[50730] ^ n[50731];
assign t[50732] = t[50731] ^ n[50732];
assign t[50733] = t[50732] ^ n[50733];
assign t[50734] = t[50733] ^ n[50734];
assign t[50735] = t[50734] ^ n[50735];
assign t[50736] = t[50735] ^ n[50736];
assign t[50737] = t[50736] ^ n[50737];
assign t[50738] = t[50737] ^ n[50738];
assign t[50739] = t[50738] ^ n[50739];
assign t[50740] = t[50739] ^ n[50740];
assign t[50741] = t[50740] ^ n[50741];
assign t[50742] = t[50741] ^ n[50742];
assign t[50743] = t[50742] ^ n[50743];
assign t[50744] = t[50743] ^ n[50744];
assign t[50745] = t[50744] ^ n[50745];
assign t[50746] = t[50745] ^ n[50746];
assign t[50747] = t[50746] ^ n[50747];
assign t[50748] = t[50747] ^ n[50748];
assign t[50749] = t[50748] ^ n[50749];
assign t[50750] = t[50749] ^ n[50750];
assign t[50751] = t[50750] ^ n[50751];
assign t[50752] = t[50751] ^ n[50752];
assign t[50753] = t[50752] ^ n[50753];
assign t[50754] = t[50753] ^ n[50754];
assign t[50755] = t[50754] ^ n[50755];
assign t[50756] = t[50755] ^ n[50756];
assign t[50757] = t[50756] ^ n[50757];
assign t[50758] = t[50757] ^ n[50758];
assign t[50759] = t[50758] ^ n[50759];
assign t[50760] = t[50759] ^ n[50760];
assign t[50761] = t[50760] ^ n[50761];
assign t[50762] = t[50761] ^ n[50762];
assign t[50763] = t[50762] ^ n[50763];
assign t[50764] = t[50763] ^ n[50764];
assign t[50765] = t[50764] ^ n[50765];
assign t[50766] = t[50765] ^ n[50766];
assign t[50767] = t[50766] ^ n[50767];
assign t[50768] = t[50767] ^ n[50768];
assign t[50769] = t[50768] ^ n[50769];
assign t[50770] = t[50769] ^ n[50770];
assign t[50771] = t[50770] ^ n[50771];
assign t[50772] = t[50771] ^ n[50772];
assign t[50773] = t[50772] ^ n[50773];
assign t[50774] = t[50773] ^ n[50774];
assign t[50775] = t[50774] ^ n[50775];
assign t[50776] = t[50775] ^ n[50776];
assign t[50777] = t[50776] ^ n[50777];
assign t[50778] = t[50777] ^ n[50778];
assign t[50779] = t[50778] ^ n[50779];
assign t[50780] = t[50779] ^ n[50780];
assign t[50781] = t[50780] ^ n[50781];
assign t[50782] = t[50781] ^ n[50782];
assign t[50783] = t[50782] ^ n[50783];
assign t[50784] = t[50783] ^ n[50784];
assign t[50785] = t[50784] ^ n[50785];
assign t[50786] = t[50785] ^ n[50786];
assign t[50787] = t[50786] ^ n[50787];
assign t[50788] = t[50787] ^ n[50788];
assign t[50789] = t[50788] ^ n[50789];
assign t[50790] = t[50789] ^ n[50790];
assign t[50791] = t[50790] ^ n[50791];
assign t[50792] = t[50791] ^ n[50792];
assign t[50793] = t[50792] ^ n[50793];
assign t[50794] = t[50793] ^ n[50794];
assign t[50795] = t[50794] ^ n[50795];
assign t[50796] = t[50795] ^ n[50796];
assign t[50797] = t[50796] ^ n[50797];
assign t[50798] = t[50797] ^ n[50798];
assign t[50799] = t[50798] ^ n[50799];
assign t[50800] = t[50799] ^ n[50800];
assign t[50801] = t[50800] ^ n[50801];
assign t[50802] = t[50801] ^ n[50802];
assign t[50803] = t[50802] ^ n[50803];
assign t[50804] = t[50803] ^ n[50804];
assign t[50805] = t[50804] ^ n[50805];
assign t[50806] = t[50805] ^ n[50806];
assign t[50807] = t[50806] ^ n[50807];
assign t[50808] = t[50807] ^ n[50808];
assign t[50809] = t[50808] ^ n[50809];
assign t[50810] = t[50809] ^ n[50810];
assign t[50811] = t[50810] ^ n[50811];
assign t[50812] = t[50811] ^ n[50812];
assign t[50813] = t[50812] ^ n[50813];
assign t[50814] = t[50813] ^ n[50814];
assign t[50815] = t[50814] ^ n[50815];
assign t[50816] = t[50815] ^ n[50816];
assign t[50817] = t[50816] ^ n[50817];
assign t[50818] = t[50817] ^ n[50818];
assign t[50819] = t[50818] ^ n[50819];
assign t[50820] = t[50819] ^ n[50820];
assign t[50821] = t[50820] ^ n[50821];
assign t[50822] = t[50821] ^ n[50822];
assign t[50823] = t[50822] ^ n[50823];
assign t[50824] = t[50823] ^ n[50824];
assign t[50825] = t[50824] ^ n[50825];
assign t[50826] = t[50825] ^ n[50826];
assign t[50827] = t[50826] ^ n[50827];
assign t[50828] = t[50827] ^ n[50828];
assign t[50829] = t[50828] ^ n[50829];
assign t[50830] = t[50829] ^ n[50830];
assign t[50831] = t[50830] ^ n[50831];
assign t[50832] = t[50831] ^ n[50832];
assign t[50833] = t[50832] ^ n[50833];
assign t[50834] = t[50833] ^ n[50834];
assign t[50835] = t[50834] ^ n[50835];
assign t[50836] = t[50835] ^ n[50836];
assign t[50837] = t[50836] ^ n[50837];
assign t[50838] = t[50837] ^ n[50838];
assign t[50839] = t[50838] ^ n[50839];
assign t[50840] = t[50839] ^ n[50840];
assign t[50841] = t[50840] ^ n[50841];
assign t[50842] = t[50841] ^ n[50842];
assign t[50843] = t[50842] ^ n[50843];
assign t[50844] = t[50843] ^ n[50844];
assign t[50845] = t[50844] ^ n[50845];
assign t[50846] = t[50845] ^ n[50846];
assign t[50847] = t[50846] ^ n[50847];
assign t[50848] = t[50847] ^ n[50848];
assign t[50849] = t[50848] ^ n[50849];
assign t[50850] = t[50849] ^ n[50850];
assign t[50851] = t[50850] ^ n[50851];
assign t[50852] = t[50851] ^ n[50852];
assign t[50853] = t[50852] ^ n[50853];
assign t[50854] = t[50853] ^ n[50854];
assign t[50855] = t[50854] ^ n[50855];
assign t[50856] = t[50855] ^ n[50856];
assign t[50857] = t[50856] ^ n[50857];
assign t[50858] = t[50857] ^ n[50858];
assign t[50859] = t[50858] ^ n[50859];
assign t[50860] = t[50859] ^ n[50860];
assign t[50861] = t[50860] ^ n[50861];
assign t[50862] = t[50861] ^ n[50862];
assign t[50863] = t[50862] ^ n[50863];
assign t[50864] = t[50863] ^ n[50864];
assign t[50865] = t[50864] ^ n[50865];
assign t[50866] = t[50865] ^ n[50866];
assign t[50867] = t[50866] ^ n[50867];
assign t[50868] = t[50867] ^ n[50868];
assign t[50869] = t[50868] ^ n[50869];
assign t[50870] = t[50869] ^ n[50870];
assign t[50871] = t[50870] ^ n[50871];
assign t[50872] = t[50871] ^ n[50872];
assign t[50873] = t[50872] ^ n[50873];
assign t[50874] = t[50873] ^ n[50874];
assign t[50875] = t[50874] ^ n[50875];
assign t[50876] = t[50875] ^ n[50876];
assign t[50877] = t[50876] ^ n[50877];
assign t[50878] = t[50877] ^ n[50878];
assign t[50879] = t[50878] ^ n[50879];
assign t[50880] = t[50879] ^ n[50880];
assign t[50881] = t[50880] ^ n[50881];
assign t[50882] = t[50881] ^ n[50882];
assign t[50883] = t[50882] ^ n[50883];
assign t[50884] = t[50883] ^ n[50884];
assign t[50885] = t[50884] ^ n[50885];
assign t[50886] = t[50885] ^ n[50886];
assign t[50887] = t[50886] ^ n[50887];
assign t[50888] = t[50887] ^ n[50888];
assign t[50889] = t[50888] ^ n[50889];
assign t[50890] = t[50889] ^ n[50890];
assign t[50891] = t[50890] ^ n[50891];
assign t[50892] = t[50891] ^ n[50892];
assign t[50893] = t[50892] ^ n[50893];
assign t[50894] = t[50893] ^ n[50894];
assign t[50895] = t[50894] ^ n[50895];
assign t[50896] = t[50895] ^ n[50896];
assign t[50897] = t[50896] ^ n[50897];
assign t[50898] = t[50897] ^ n[50898];
assign t[50899] = t[50898] ^ n[50899];
assign t[50900] = t[50899] ^ n[50900];
assign t[50901] = t[50900] ^ n[50901];
assign t[50902] = t[50901] ^ n[50902];
assign t[50903] = t[50902] ^ n[50903];
assign t[50904] = t[50903] ^ n[50904];
assign t[50905] = t[50904] ^ n[50905];
assign t[50906] = t[50905] ^ n[50906];
assign t[50907] = t[50906] ^ n[50907];
assign t[50908] = t[50907] ^ n[50908];
assign t[50909] = t[50908] ^ n[50909];
assign t[50910] = t[50909] ^ n[50910];
assign t[50911] = t[50910] ^ n[50911];
assign t[50912] = t[50911] ^ n[50912];
assign t[50913] = t[50912] ^ n[50913];
assign t[50914] = t[50913] ^ n[50914];
assign t[50915] = t[50914] ^ n[50915];
assign t[50916] = t[50915] ^ n[50916];
assign t[50917] = t[50916] ^ n[50917];
assign t[50918] = t[50917] ^ n[50918];
assign t[50919] = t[50918] ^ n[50919];
assign t[50920] = t[50919] ^ n[50920];
assign t[50921] = t[50920] ^ n[50921];
assign t[50922] = t[50921] ^ n[50922];
assign t[50923] = t[50922] ^ n[50923];
assign t[50924] = t[50923] ^ n[50924];
assign t[50925] = t[50924] ^ n[50925];
assign t[50926] = t[50925] ^ n[50926];
assign t[50927] = t[50926] ^ n[50927];
assign t[50928] = t[50927] ^ n[50928];
assign t[50929] = t[50928] ^ n[50929];
assign t[50930] = t[50929] ^ n[50930];
assign t[50931] = t[50930] ^ n[50931];
assign t[50932] = t[50931] ^ n[50932];
assign t[50933] = t[50932] ^ n[50933];
assign t[50934] = t[50933] ^ n[50934];
assign t[50935] = t[50934] ^ n[50935];
assign t[50936] = t[50935] ^ n[50936];
assign t[50937] = t[50936] ^ n[50937];
assign t[50938] = t[50937] ^ n[50938];
assign t[50939] = t[50938] ^ n[50939];
assign t[50940] = t[50939] ^ n[50940];
assign t[50941] = t[50940] ^ n[50941];
assign t[50942] = t[50941] ^ n[50942];
assign t[50943] = t[50942] ^ n[50943];
assign t[50944] = t[50943] ^ n[50944];
assign t[50945] = t[50944] ^ n[50945];
assign t[50946] = t[50945] ^ n[50946];
assign t[50947] = t[50946] ^ n[50947];
assign t[50948] = t[50947] ^ n[50948];
assign t[50949] = t[50948] ^ n[50949];
assign t[50950] = t[50949] ^ n[50950];
assign t[50951] = t[50950] ^ n[50951];
assign t[50952] = t[50951] ^ n[50952];
assign t[50953] = t[50952] ^ n[50953];
assign t[50954] = t[50953] ^ n[50954];
assign t[50955] = t[50954] ^ n[50955];
assign t[50956] = t[50955] ^ n[50956];
assign t[50957] = t[50956] ^ n[50957];
assign t[50958] = t[50957] ^ n[50958];
assign t[50959] = t[50958] ^ n[50959];
assign t[50960] = t[50959] ^ n[50960];
assign t[50961] = t[50960] ^ n[50961];
assign t[50962] = t[50961] ^ n[50962];
assign t[50963] = t[50962] ^ n[50963];
assign t[50964] = t[50963] ^ n[50964];
assign t[50965] = t[50964] ^ n[50965];
assign t[50966] = t[50965] ^ n[50966];
assign t[50967] = t[50966] ^ n[50967];
assign t[50968] = t[50967] ^ n[50968];
assign t[50969] = t[50968] ^ n[50969];
assign t[50970] = t[50969] ^ n[50970];
assign t[50971] = t[50970] ^ n[50971];
assign t[50972] = t[50971] ^ n[50972];
assign t[50973] = t[50972] ^ n[50973];
assign t[50974] = t[50973] ^ n[50974];
assign t[50975] = t[50974] ^ n[50975];
assign t[50976] = t[50975] ^ n[50976];
assign t[50977] = t[50976] ^ n[50977];
assign t[50978] = t[50977] ^ n[50978];
assign t[50979] = t[50978] ^ n[50979];
assign t[50980] = t[50979] ^ n[50980];
assign t[50981] = t[50980] ^ n[50981];
assign t[50982] = t[50981] ^ n[50982];
assign t[50983] = t[50982] ^ n[50983];
assign t[50984] = t[50983] ^ n[50984];
assign t[50985] = t[50984] ^ n[50985];
assign t[50986] = t[50985] ^ n[50986];
assign t[50987] = t[50986] ^ n[50987];
assign t[50988] = t[50987] ^ n[50988];
assign t[50989] = t[50988] ^ n[50989];
assign t[50990] = t[50989] ^ n[50990];
assign t[50991] = t[50990] ^ n[50991];
assign t[50992] = t[50991] ^ n[50992];
assign t[50993] = t[50992] ^ n[50993];
assign t[50994] = t[50993] ^ n[50994];
assign t[50995] = t[50994] ^ n[50995];
assign t[50996] = t[50995] ^ n[50996];
assign t[50997] = t[50996] ^ n[50997];
assign t[50998] = t[50997] ^ n[50998];
assign t[50999] = t[50998] ^ n[50999];
assign t[51000] = t[50999] ^ n[51000];
assign t[51001] = t[51000] ^ n[51001];
assign t[51002] = t[51001] ^ n[51002];
assign t[51003] = t[51002] ^ n[51003];
assign t[51004] = t[51003] ^ n[51004];
assign t[51005] = t[51004] ^ n[51005];
assign t[51006] = t[51005] ^ n[51006];
assign t[51007] = t[51006] ^ n[51007];
assign t[51008] = t[51007] ^ n[51008];
assign t[51009] = t[51008] ^ n[51009];
assign t[51010] = t[51009] ^ n[51010];
assign t[51011] = t[51010] ^ n[51011];
assign t[51012] = t[51011] ^ n[51012];
assign t[51013] = t[51012] ^ n[51013];
assign t[51014] = t[51013] ^ n[51014];
assign t[51015] = t[51014] ^ n[51015];
assign t[51016] = t[51015] ^ n[51016];
assign t[51017] = t[51016] ^ n[51017];
assign t[51018] = t[51017] ^ n[51018];
assign t[51019] = t[51018] ^ n[51019];
assign t[51020] = t[51019] ^ n[51020];
assign t[51021] = t[51020] ^ n[51021];
assign t[51022] = t[51021] ^ n[51022];
assign t[51023] = t[51022] ^ n[51023];
assign t[51024] = t[51023] ^ n[51024];
assign t[51025] = t[51024] ^ n[51025];
assign t[51026] = t[51025] ^ n[51026];
assign t[51027] = t[51026] ^ n[51027];
assign t[51028] = t[51027] ^ n[51028];
assign t[51029] = t[51028] ^ n[51029];
assign t[51030] = t[51029] ^ n[51030];
assign t[51031] = t[51030] ^ n[51031];
assign t[51032] = t[51031] ^ n[51032];
assign t[51033] = t[51032] ^ n[51033];
assign t[51034] = t[51033] ^ n[51034];
assign t[51035] = t[51034] ^ n[51035];
assign t[51036] = t[51035] ^ n[51036];
assign t[51037] = t[51036] ^ n[51037];
assign t[51038] = t[51037] ^ n[51038];
assign t[51039] = t[51038] ^ n[51039];
assign t[51040] = t[51039] ^ n[51040];
assign t[51041] = t[51040] ^ n[51041];
assign t[51042] = t[51041] ^ n[51042];
assign t[51043] = t[51042] ^ n[51043];
assign t[51044] = t[51043] ^ n[51044];
assign t[51045] = t[51044] ^ n[51045];
assign t[51046] = t[51045] ^ n[51046];
assign t[51047] = t[51046] ^ n[51047];
assign t[51048] = t[51047] ^ n[51048];
assign t[51049] = t[51048] ^ n[51049];
assign t[51050] = t[51049] ^ n[51050];
assign t[51051] = t[51050] ^ n[51051];
assign t[51052] = t[51051] ^ n[51052];
assign t[51053] = t[51052] ^ n[51053];
assign t[51054] = t[51053] ^ n[51054];
assign t[51055] = t[51054] ^ n[51055];
assign t[51056] = t[51055] ^ n[51056];
assign t[51057] = t[51056] ^ n[51057];
assign t[51058] = t[51057] ^ n[51058];
assign t[51059] = t[51058] ^ n[51059];
assign t[51060] = t[51059] ^ n[51060];
assign t[51061] = t[51060] ^ n[51061];
assign t[51062] = t[51061] ^ n[51062];
assign t[51063] = t[51062] ^ n[51063];
assign t[51064] = t[51063] ^ n[51064];
assign t[51065] = t[51064] ^ n[51065];
assign t[51066] = t[51065] ^ n[51066];
assign t[51067] = t[51066] ^ n[51067];
assign t[51068] = t[51067] ^ n[51068];
assign t[51069] = t[51068] ^ n[51069];
assign t[51070] = t[51069] ^ n[51070];
assign t[51071] = t[51070] ^ n[51071];
assign t[51072] = t[51071] ^ n[51072];
assign t[51073] = t[51072] ^ n[51073];
assign t[51074] = t[51073] ^ n[51074];
assign t[51075] = t[51074] ^ n[51075];
assign t[51076] = t[51075] ^ n[51076];
assign t[51077] = t[51076] ^ n[51077];
assign t[51078] = t[51077] ^ n[51078];
assign t[51079] = t[51078] ^ n[51079];
assign t[51080] = t[51079] ^ n[51080];
assign t[51081] = t[51080] ^ n[51081];
assign t[51082] = t[51081] ^ n[51082];
assign t[51083] = t[51082] ^ n[51083];
assign t[51084] = t[51083] ^ n[51084];
assign t[51085] = t[51084] ^ n[51085];
assign t[51086] = t[51085] ^ n[51086];
assign t[51087] = t[51086] ^ n[51087];
assign t[51088] = t[51087] ^ n[51088];
assign t[51089] = t[51088] ^ n[51089];
assign t[51090] = t[51089] ^ n[51090];
assign t[51091] = t[51090] ^ n[51091];
assign t[51092] = t[51091] ^ n[51092];
assign t[51093] = t[51092] ^ n[51093];
assign t[51094] = t[51093] ^ n[51094];
assign t[51095] = t[51094] ^ n[51095];
assign t[51096] = t[51095] ^ n[51096];
assign t[51097] = t[51096] ^ n[51097];
assign t[51098] = t[51097] ^ n[51098];
assign t[51099] = t[51098] ^ n[51099];
assign t[51100] = t[51099] ^ n[51100];
assign t[51101] = t[51100] ^ n[51101];
assign t[51102] = t[51101] ^ n[51102];
assign t[51103] = t[51102] ^ n[51103];
assign t[51104] = t[51103] ^ n[51104];
assign t[51105] = t[51104] ^ n[51105];
assign t[51106] = t[51105] ^ n[51106];
assign t[51107] = t[51106] ^ n[51107];
assign t[51108] = t[51107] ^ n[51108];
assign t[51109] = t[51108] ^ n[51109];
assign t[51110] = t[51109] ^ n[51110];
assign t[51111] = t[51110] ^ n[51111];
assign t[51112] = t[51111] ^ n[51112];
assign t[51113] = t[51112] ^ n[51113];
assign t[51114] = t[51113] ^ n[51114];
assign t[51115] = t[51114] ^ n[51115];
assign t[51116] = t[51115] ^ n[51116];
assign t[51117] = t[51116] ^ n[51117];
assign t[51118] = t[51117] ^ n[51118];
assign t[51119] = t[51118] ^ n[51119];
assign t[51120] = t[51119] ^ n[51120];
assign t[51121] = t[51120] ^ n[51121];
assign t[51122] = t[51121] ^ n[51122];
assign t[51123] = t[51122] ^ n[51123];
assign t[51124] = t[51123] ^ n[51124];
assign t[51125] = t[51124] ^ n[51125];
assign t[51126] = t[51125] ^ n[51126];
assign t[51127] = t[51126] ^ n[51127];
assign t[51128] = t[51127] ^ n[51128];
assign t[51129] = t[51128] ^ n[51129];
assign t[51130] = t[51129] ^ n[51130];
assign t[51131] = t[51130] ^ n[51131];
assign t[51132] = t[51131] ^ n[51132];
assign t[51133] = t[51132] ^ n[51133];
assign t[51134] = t[51133] ^ n[51134];
assign t[51135] = t[51134] ^ n[51135];
assign t[51136] = t[51135] ^ n[51136];
assign t[51137] = t[51136] ^ n[51137];
assign t[51138] = t[51137] ^ n[51138];
assign t[51139] = t[51138] ^ n[51139];
assign t[51140] = t[51139] ^ n[51140];
assign t[51141] = t[51140] ^ n[51141];
assign t[51142] = t[51141] ^ n[51142];
assign t[51143] = t[51142] ^ n[51143];
assign t[51144] = t[51143] ^ n[51144];
assign t[51145] = t[51144] ^ n[51145];
assign t[51146] = t[51145] ^ n[51146];
assign t[51147] = t[51146] ^ n[51147];
assign t[51148] = t[51147] ^ n[51148];
assign t[51149] = t[51148] ^ n[51149];
assign t[51150] = t[51149] ^ n[51150];
assign t[51151] = t[51150] ^ n[51151];
assign t[51152] = t[51151] ^ n[51152];
assign t[51153] = t[51152] ^ n[51153];
assign t[51154] = t[51153] ^ n[51154];
assign t[51155] = t[51154] ^ n[51155];
assign t[51156] = t[51155] ^ n[51156];
assign t[51157] = t[51156] ^ n[51157];
assign t[51158] = t[51157] ^ n[51158];
assign t[51159] = t[51158] ^ n[51159];
assign t[51160] = t[51159] ^ n[51160];
assign t[51161] = t[51160] ^ n[51161];
assign t[51162] = t[51161] ^ n[51162];
assign t[51163] = t[51162] ^ n[51163];
assign t[51164] = t[51163] ^ n[51164];
assign t[51165] = t[51164] ^ n[51165];
assign t[51166] = t[51165] ^ n[51166];
assign t[51167] = t[51166] ^ n[51167];
assign t[51168] = t[51167] ^ n[51168];
assign t[51169] = t[51168] ^ n[51169];
assign t[51170] = t[51169] ^ n[51170];
assign t[51171] = t[51170] ^ n[51171];
assign t[51172] = t[51171] ^ n[51172];
assign t[51173] = t[51172] ^ n[51173];
assign t[51174] = t[51173] ^ n[51174];
assign t[51175] = t[51174] ^ n[51175];
assign t[51176] = t[51175] ^ n[51176];
assign t[51177] = t[51176] ^ n[51177];
assign t[51178] = t[51177] ^ n[51178];
assign t[51179] = t[51178] ^ n[51179];
assign t[51180] = t[51179] ^ n[51180];
assign t[51181] = t[51180] ^ n[51181];
assign t[51182] = t[51181] ^ n[51182];
assign t[51183] = t[51182] ^ n[51183];
assign t[51184] = t[51183] ^ n[51184];
assign t[51185] = t[51184] ^ n[51185];
assign t[51186] = t[51185] ^ n[51186];
assign t[51187] = t[51186] ^ n[51187];
assign t[51188] = t[51187] ^ n[51188];
assign t[51189] = t[51188] ^ n[51189];
assign t[51190] = t[51189] ^ n[51190];
assign t[51191] = t[51190] ^ n[51191];
assign t[51192] = t[51191] ^ n[51192];
assign t[51193] = t[51192] ^ n[51193];
assign t[51194] = t[51193] ^ n[51194];
assign t[51195] = t[51194] ^ n[51195];
assign t[51196] = t[51195] ^ n[51196];
assign t[51197] = t[51196] ^ n[51197];
assign t[51198] = t[51197] ^ n[51198];
assign t[51199] = t[51198] ^ n[51199];
assign t[51200] = t[51199] ^ n[51200];
assign t[51201] = t[51200] ^ n[51201];
assign t[51202] = t[51201] ^ n[51202];
assign t[51203] = t[51202] ^ n[51203];
assign t[51204] = t[51203] ^ n[51204];
assign t[51205] = t[51204] ^ n[51205];
assign t[51206] = t[51205] ^ n[51206];
assign t[51207] = t[51206] ^ n[51207];
assign t[51208] = t[51207] ^ n[51208];
assign t[51209] = t[51208] ^ n[51209];
assign t[51210] = t[51209] ^ n[51210];
assign t[51211] = t[51210] ^ n[51211];
assign t[51212] = t[51211] ^ n[51212];
assign t[51213] = t[51212] ^ n[51213];
assign t[51214] = t[51213] ^ n[51214];
assign t[51215] = t[51214] ^ n[51215];
assign t[51216] = t[51215] ^ n[51216];
assign t[51217] = t[51216] ^ n[51217];
assign t[51218] = t[51217] ^ n[51218];
assign t[51219] = t[51218] ^ n[51219];
assign t[51220] = t[51219] ^ n[51220];
assign t[51221] = t[51220] ^ n[51221];
assign t[51222] = t[51221] ^ n[51222];
assign t[51223] = t[51222] ^ n[51223];
assign t[51224] = t[51223] ^ n[51224];
assign t[51225] = t[51224] ^ n[51225];
assign t[51226] = t[51225] ^ n[51226];
assign t[51227] = t[51226] ^ n[51227];
assign t[51228] = t[51227] ^ n[51228];
assign t[51229] = t[51228] ^ n[51229];
assign t[51230] = t[51229] ^ n[51230];
assign t[51231] = t[51230] ^ n[51231];
assign t[51232] = t[51231] ^ n[51232];
assign t[51233] = t[51232] ^ n[51233];
assign t[51234] = t[51233] ^ n[51234];
assign t[51235] = t[51234] ^ n[51235];
assign t[51236] = t[51235] ^ n[51236];
assign t[51237] = t[51236] ^ n[51237];
assign t[51238] = t[51237] ^ n[51238];
assign t[51239] = t[51238] ^ n[51239];
assign t[51240] = t[51239] ^ n[51240];
assign t[51241] = t[51240] ^ n[51241];
assign t[51242] = t[51241] ^ n[51242];
assign t[51243] = t[51242] ^ n[51243];
assign t[51244] = t[51243] ^ n[51244];
assign t[51245] = t[51244] ^ n[51245];
assign t[51246] = t[51245] ^ n[51246];
assign t[51247] = t[51246] ^ n[51247];
assign t[51248] = t[51247] ^ n[51248];
assign t[51249] = t[51248] ^ n[51249];
assign t[51250] = t[51249] ^ n[51250];
assign t[51251] = t[51250] ^ n[51251];
assign t[51252] = t[51251] ^ n[51252];
assign t[51253] = t[51252] ^ n[51253];
assign t[51254] = t[51253] ^ n[51254];
assign t[51255] = t[51254] ^ n[51255];
assign t[51256] = t[51255] ^ n[51256];
assign t[51257] = t[51256] ^ n[51257];
assign t[51258] = t[51257] ^ n[51258];
assign t[51259] = t[51258] ^ n[51259];
assign t[51260] = t[51259] ^ n[51260];
assign t[51261] = t[51260] ^ n[51261];
assign t[51262] = t[51261] ^ n[51262];
assign t[51263] = t[51262] ^ n[51263];
assign t[51264] = t[51263] ^ n[51264];
assign t[51265] = t[51264] ^ n[51265];
assign t[51266] = t[51265] ^ n[51266];
assign t[51267] = t[51266] ^ n[51267];
assign t[51268] = t[51267] ^ n[51268];
assign t[51269] = t[51268] ^ n[51269];
assign t[51270] = t[51269] ^ n[51270];
assign t[51271] = t[51270] ^ n[51271];
assign t[51272] = t[51271] ^ n[51272];
assign t[51273] = t[51272] ^ n[51273];
assign t[51274] = t[51273] ^ n[51274];
assign t[51275] = t[51274] ^ n[51275];
assign t[51276] = t[51275] ^ n[51276];
assign t[51277] = t[51276] ^ n[51277];
assign t[51278] = t[51277] ^ n[51278];
assign t[51279] = t[51278] ^ n[51279];
assign t[51280] = t[51279] ^ n[51280];
assign t[51281] = t[51280] ^ n[51281];
assign t[51282] = t[51281] ^ n[51282];
assign t[51283] = t[51282] ^ n[51283];
assign t[51284] = t[51283] ^ n[51284];
assign t[51285] = t[51284] ^ n[51285];
assign t[51286] = t[51285] ^ n[51286];
assign t[51287] = t[51286] ^ n[51287];
assign t[51288] = t[51287] ^ n[51288];
assign t[51289] = t[51288] ^ n[51289];
assign t[51290] = t[51289] ^ n[51290];
assign t[51291] = t[51290] ^ n[51291];
assign t[51292] = t[51291] ^ n[51292];
assign t[51293] = t[51292] ^ n[51293];
assign t[51294] = t[51293] ^ n[51294];
assign t[51295] = t[51294] ^ n[51295];
assign t[51296] = t[51295] ^ n[51296];
assign t[51297] = t[51296] ^ n[51297];
assign t[51298] = t[51297] ^ n[51298];
assign t[51299] = t[51298] ^ n[51299];
assign t[51300] = t[51299] ^ n[51300];
assign t[51301] = t[51300] ^ n[51301];
assign t[51302] = t[51301] ^ n[51302];
assign t[51303] = t[51302] ^ n[51303];
assign t[51304] = t[51303] ^ n[51304];
assign t[51305] = t[51304] ^ n[51305];
assign t[51306] = t[51305] ^ n[51306];
assign t[51307] = t[51306] ^ n[51307];
assign t[51308] = t[51307] ^ n[51308];
assign t[51309] = t[51308] ^ n[51309];
assign t[51310] = t[51309] ^ n[51310];
assign t[51311] = t[51310] ^ n[51311];
assign t[51312] = t[51311] ^ n[51312];
assign t[51313] = t[51312] ^ n[51313];
assign t[51314] = t[51313] ^ n[51314];
assign t[51315] = t[51314] ^ n[51315];
assign t[51316] = t[51315] ^ n[51316];
assign t[51317] = t[51316] ^ n[51317];
assign t[51318] = t[51317] ^ n[51318];
assign t[51319] = t[51318] ^ n[51319];
assign t[51320] = t[51319] ^ n[51320];
assign t[51321] = t[51320] ^ n[51321];
assign t[51322] = t[51321] ^ n[51322];
assign t[51323] = t[51322] ^ n[51323];
assign t[51324] = t[51323] ^ n[51324];
assign t[51325] = t[51324] ^ n[51325];
assign t[51326] = t[51325] ^ n[51326];
assign t[51327] = t[51326] ^ n[51327];
assign t[51328] = t[51327] ^ n[51328];
assign t[51329] = t[51328] ^ n[51329];
assign t[51330] = t[51329] ^ n[51330];
assign t[51331] = t[51330] ^ n[51331];
assign t[51332] = t[51331] ^ n[51332];
assign t[51333] = t[51332] ^ n[51333];
assign t[51334] = t[51333] ^ n[51334];
assign t[51335] = t[51334] ^ n[51335];
assign t[51336] = t[51335] ^ n[51336];
assign t[51337] = t[51336] ^ n[51337];
assign t[51338] = t[51337] ^ n[51338];
assign t[51339] = t[51338] ^ n[51339];
assign t[51340] = t[51339] ^ n[51340];
assign t[51341] = t[51340] ^ n[51341];
assign t[51342] = t[51341] ^ n[51342];
assign t[51343] = t[51342] ^ n[51343];
assign t[51344] = t[51343] ^ n[51344];
assign t[51345] = t[51344] ^ n[51345];
assign t[51346] = t[51345] ^ n[51346];
assign t[51347] = t[51346] ^ n[51347];
assign t[51348] = t[51347] ^ n[51348];
assign t[51349] = t[51348] ^ n[51349];
assign t[51350] = t[51349] ^ n[51350];
assign t[51351] = t[51350] ^ n[51351];
assign t[51352] = t[51351] ^ n[51352];
assign t[51353] = t[51352] ^ n[51353];
assign t[51354] = t[51353] ^ n[51354];
assign t[51355] = t[51354] ^ n[51355];
assign t[51356] = t[51355] ^ n[51356];
assign t[51357] = t[51356] ^ n[51357];
assign t[51358] = t[51357] ^ n[51358];
assign t[51359] = t[51358] ^ n[51359];
assign t[51360] = t[51359] ^ n[51360];
assign t[51361] = t[51360] ^ n[51361];
assign t[51362] = t[51361] ^ n[51362];
assign t[51363] = t[51362] ^ n[51363];
assign t[51364] = t[51363] ^ n[51364];
assign t[51365] = t[51364] ^ n[51365];
assign t[51366] = t[51365] ^ n[51366];
assign t[51367] = t[51366] ^ n[51367];
assign t[51368] = t[51367] ^ n[51368];
assign t[51369] = t[51368] ^ n[51369];
assign t[51370] = t[51369] ^ n[51370];
assign t[51371] = t[51370] ^ n[51371];
assign t[51372] = t[51371] ^ n[51372];
assign t[51373] = t[51372] ^ n[51373];
assign t[51374] = t[51373] ^ n[51374];
assign t[51375] = t[51374] ^ n[51375];
assign t[51376] = t[51375] ^ n[51376];
assign t[51377] = t[51376] ^ n[51377];
assign t[51378] = t[51377] ^ n[51378];
assign t[51379] = t[51378] ^ n[51379];
assign t[51380] = t[51379] ^ n[51380];
assign t[51381] = t[51380] ^ n[51381];
assign t[51382] = t[51381] ^ n[51382];
assign t[51383] = t[51382] ^ n[51383];
assign t[51384] = t[51383] ^ n[51384];
assign t[51385] = t[51384] ^ n[51385];
assign t[51386] = t[51385] ^ n[51386];
assign t[51387] = t[51386] ^ n[51387];
assign t[51388] = t[51387] ^ n[51388];
assign t[51389] = t[51388] ^ n[51389];
assign t[51390] = t[51389] ^ n[51390];
assign t[51391] = t[51390] ^ n[51391];
assign t[51392] = t[51391] ^ n[51392];
assign t[51393] = t[51392] ^ n[51393];
assign t[51394] = t[51393] ^ n[51394];
assign t[51395] = t[51394] ^ n[51395];
assign t[51396] = t[51395] ^ n[51396];
assign t[51397] = t[51396] ^ n[51397];
assign t[51398] = t[51397] ^ n[51398];
assign t[51399] = t[51398] ^ n[51399];
assign t[51400] = t[51399] ^ n[51400];
assign t[51401] = t[51400] ^ n[51401];
assign t[51402] = t[51401] ^ n[51402];
assign t[51403] = t[51402] ^ n[51403];
assign t[51404] = t[51403] ^ n[51404];
assign t[51405] = t[51404] ^ n[51405];
assign t[51406] = t[51405] ^ n[51406];
assign t[51407] = t[51406] ^ n[51407];
assign t[51408] = t[51407] ^ n[51408];
assign t[51409] = t[51408] ^ n[51409];
assign t[51410] = t[51409] ^ n[51410];
assign t[51411] = t[51410] ^ n[51411];
assign t[51412] = t[51411] ^ n[51412];
assign t[51413] = t[51412] ^ n[51413];
assign t[51414] = t[51413] ^ n[51414];
assign t[51415] = t[51414] ^ n[51415];
assign t[51416] = t[51415] ^ n[51416];
assign t[51417] = t[51416] ^ n[51417];
assign t[51418] = t[51417] ^ n[51418];
assign t[51419] = t[51418] ^ n[51419];
assign t[51420] = t[51419] ^ n[51420];
assign t[51421] = t[51420] ^ n[51421];
assign t[51422] = t[51421] ^ n[51422];
assign t[51423] = t[51422] ^ n[51423];
assign t[51424] = t[51423] ^ n[51424];
assign t[51425] = t[51424] ^ n[51425];
assign t[51426] = t[51425] ^ n[51426];
assign t[51427] = t[51426] ^ n[51427];
assign t[51428] = t[51427] ^ n[51428];
assign t[51429] = t[51428] ^ n[51429];
assign t[51430] = t[51429] ^ n[51430];
assign t[51431] = t[51430] ^ n[51431];
assign t[51432] = t[51431] ^ n[51432];
assign t[51433] = t[51432] ^ n[51433];
assign t[51434] = t[51433] ^ n[51434];
assign t[51435] = t[51434] ^ n[51435];
assign t[51436] = t[51435] ^ n[51436];
assign t[51437] = t[51436] ^ n[51437];
assign t[51438] = t[51437] ^ n[51438];
assign t[51439] = t[51438] ^ n[51439];
assign t[51440] = t[51439] ^ n[51440];
assign t[51441] = t[51440] ^ n[51441];
assign t[51442] = t[51441] ^ n[51442];
assign t[51443] = t[51442] ^ n[51443];
assign t[51444] = t[51443] ^ n[51444];
assign t[51445] = t[51444] ^ n[51445];
assign t[51446] = t[51445] ^ n[51446];
assign t[51447] = t[51446] ^ n[51447];
assign t[51448] = t[51447] ^ n[51448];
assign t[51449] = t[51448] ^ n[51449];
assign t[51450] = t[51449] ^ n[51450];
assign t[51451] = t[51450] ^ n[51451];
assign t[51452] = t[51451] ^ n[51452];
assign t[51453] = t[51452] ^ n[51453];
assign t[51454] = t[51453] ^ n[51454];
assign t[51455] = t[51454] ^ n[51455];
assign t[51456] = t[51455] ^ n[51456];
assign t[51457] = t[51456] ^ n[51457];
assign t[51458] = t[51457] ^ n[51458];
assign t[51459] = t[51458] ^ n[51459];
assign t[51460] = t[51459] ^ n[51460];
assign t[51461] = t[51460] ^ n[51461];
assign t[51462] = t[51461] ^ n[51462];
assign t[51463] = t[51462] ^ n[51463];
assign t[51464] = t[51463] ^ n[51464];
assign t[51465] = t[51464] ^ n[51465];
assign t[51466] = t[51465] ^ n[51466];
assign t[51467] = t[51466] ^ n[51467];
assign t[51468] = t[51467] ^ n[51468];
assign t[51469] = t[51468] ^ n[51469];
assign t[51470] = t[51469] ^ n[51470];
assign t[51471] = t[51470] ^ n[51471];
assign t[51472] = t[51471] ^ n[51472];
assign t[51473] = t[51472] ^ n[51473];
assign t[51474] = t[51473] ^ n[51474];
assign t[51475] = t[51474] ^ n[51475];
assign t[51476] = t[51475] ^ n[51476];
assign t[51477] = t[51476] ^ n[51477];
assign t[51478] = t[51477] ^ n[51478];
assign t[51479] = t[51478] ^ n[51479];
assign t[51480] = t[51479] ^ n[51480];
assign t[51481] = t[51480] ^ n[51481];
assign t[51482] = t[51481] ^ n[51482];
assign t[51483] = t[51482] ^ n[51483];
assign t[51484] = t[51483] ^ n[51484];
assign t[51485] = t[51484] ^ n[51485];
assign t[51486] = t[51485] ^ n[51486];
assign t[51487] = t[51486] ^ n[51487];
assign t[51488] = t[51487] ^ n[51488];
assign t[51489] = t[51488] ^ n[51489];
assign t[51490] = t[51489] ^ n[51490];
assign t[51491] = t[51490] ^ n[51491];
assign t[51492] = t[51491] ^ n[51492];
assign t[51493] = t[51492] ^ n[51493];
assign t[51494] = t[51493] ^ n[51494];
assign t[51495] = t[51494] ^ n[51495];
assign t[51496] = t[51495] ^ n[51496];
assign t[51497] = t[51496] ^ n[51497];
assign t[51498] = t[51497] ^ n[51498];
assign t[51499] = t[51498] ^ n[51499];
assign t[51500] = t[51499] ^ n[51500];
assign t[51501] = t[51500] ^ n[51501];
assign t[51502] = t[51501] ^ n[51502];
assign t[51503] = t[51502] ^ n[51503];
assign t[51504] = t[51503] ^ n[51504];
assign t[51505] = t[51504] ^ n[51505];
assign t[51506] = t[51505] ^ n[51506];
assign t[51507] = t[51506] ^ n[51507];
assign t[51508] = t[51507] ^ n[51508];
assign t[51509] = t[51508] ^ n[51509];
assign t[51510] = t[51509] ^ n[51510];
assign t[51511] = t[51510] ^ n[51511];
assign t[51512] = t[51511] ^ n[51512];
assign t[51513] = t[51512] ^ n[51513];
assign t[51514] = t[51513] ^ n[51514];
assign t[51515] = t[51514] ^ n[51515];
assign t[51516] = t[51515] ^ n[51516];
assign t[51517] = t[51516] ^ n[51517];
assign t[51518] = t[51517] ^ n[51518];
assign t[51519] = t[51518] ^ n[51519];
assign t[51520] = t[51519] ^ n[51520];
assign t[51521] = t[51520] ^ n[51521];
assign t[51522] = t[51521] ^ n[51522];
assign t[51523] = t[51522] ^ n[51523];
assign t[51524] = t[51523] ^ n[51524];
assign t[51525] = t[51524] ^ n[51525];
assign t[51526] = t[51525] ^ n[51526];
assign t[51527] = t[51526] ^ n[51527];
assign t[51528] = t[51527] ^ n[51528];
assign t[51529] = t[51528] ^ n[51529];
assign t[51530] = t[51529] ^ n[51530];
assign t[51531] = t[51530] ^ n[51531];
assign t[51532] = t[51531] ^ n[51532];
assign t[51533] = t[51532] ^ n[51533];
assign t[51534] = t[51533] ^ n[51534];
assign t[51535] = t[51534] ^ n[51535];
assign t[51536] = t[51535] ^ n[51536];
assign t[51537] = t[51536] ^ n[51537];
assign t[51538] = t[51537] ^ n[51538];
assign t[51539] = t[51538] ^ n[51539];
assign t[51540] = t[51539] ^ n[51540];
assign t[51541] = t[51540] ^ n[51541];
assign t[51542] = t[51541] ^ n[51542];
assign t[51543] = t[51542] ^ n[51543];
assign t[51544] = t[51543] ^ n[51544];
assign t[51545] = t[51544] ^ n[51545];
assign t[51546] = t[51545] ^ n[51546];
assign t[51547] = t[51546] ^ n[51547];
assign t[51548] = t[51547] ^ n[51548];
assign t[51549] = t[51548] ^ n[51549];
assign t[51550] = t[51549] ^ n[51550];
assign t[51551] = t[51550] ^ n[51551];
assign t[51552] = t[51551] ^ n[51552];
assign t[51553] = t[51552] ^ n[51553];
assign t[51554] = t[51553] ^ n[51554];
assign t[51555] = t[51554] ^ n[51555];
assign t[51556] = t[51555] ^ n[51556];
assign t[51557] = t[51556] ^ n[51557];
assign t[51558] = t[51557] ^ n[51558];
assign t[51559] = t[51558] ^ n[51559];
assign t[51560] = t[51559] ^ n[51560];
assign t[51561] = t[51560] ^ n[51561];
assign t[51562] = t[51561] ^ n[51562];
assign t[51563] = t[51562] ^ n[51563];
assign t[51564] = t[51563] ^ n[51564];
assign t[51565] = t[51564] ^ n[51565];
assign t[51566] = t[51565] ^ n[51566];
assign t[51567] = t[51566] ^ n[51567];
assign t[51568] = t[51567] ^ n[51568];
assign t[51569] = t[51568] ^ n[51569];
assign t[51570] = t[51569] ^ n[51570];
assign t[51571] = t[51570] ^ n[51571];
assign t[51572] = t[51571] ^ n[51572];
assign t[51573] = t[51572] ^ n[51573];
assign t[51574] = t[51573] ^ n[51574];
assign t[51575] = t[51574] ^ n[51575];
assign t[51576] = t[51575] ^ n[51576];
assign t[51577] = t[51576] ^ n[51577];
assign t[51578] = t[51577] ^ n[51578];
assign t[51579] = t[51578] ^ n[51579];
assign t[51580] = t[51579] ^ n[51580];
assign t[51581] = t[51580] ^ n[51581];
assign t[51582] = t[51581] ^ n[51582];
assign t[51583] = t[51582] ^ n[51583];
assign t[51584] = t[51583] ^ n[51584];
assign t[51585] = t[51584] ^ n[51585];
assign t[51586] = t[51585] ^ n[51586];
assign t[51587] = t[51586] ^ n[51587];
assign t[51588] = t[51587] ^ n[51588];
assign t[51589] = t[51588] ^ n[51589];
assign t[51590] = t[51589] ^ n[51590];
assign t[51591] = t[51590] ^ n[51591];
assign t[51592] = t[51591] ^ n[51592];
assign t[51593] = t[51592] ^ n[51593];
assign t[51594] = t[51593] ^ n[51594];
assign t[51595] = t[51594] ^ n[51595];
assign t[51596] = t[51595] ^ n[51596];
assign t[51597] = t[51596] ^ n[51597];
assign t[51598] = t[51597] ^ n[51598];
assign t[51599] = t[51598] ^ n[51599];
assign t[51600] = t[51599] ^ n[51600];
assign t[51601] = t[51600] ^ n[51601];
assign t[51602] = t[51601] ^ n[51602];
assign t[51603] = t[51602] ^ n[51603];
assign t[51604] = t[51603] ^ n[51604];
assign t[51605] = t[51604] ^ n[51605];
assign t[51606] = t[51605] ^ n[51606];
assign t[51607] = t[51606] ^ n[51607];
assign t[51608] = t[51607] ^ n[51608];
assign t[51609] = t[51608] ^ n[51609];
assign t[51610] = t[51609] ^ n[51610];
assign t[51611] = t[51610] ^ n[51611];
assign t[51612] = t[51611] ^ n[51612];
assign t[51613] = t[51612] ^ n[51613];
assign t[51614] = t[51613] ^ n[51614];
assign t[51615] = t[51614] ^ n[51615];
assign t[51616] = t[51615] ^ n[51616];
assign t[51617] = t[51616] ^ n[51617];
assign t[51618] = t[51617] ^ n[51618];
assign t[51619] = t[51618] ^ n[51619];
assign t[51620] = t[51619] ^ n[51620];
assign t[51621] = t[51620] ^ n[51621];
assign t[51622] = t[51621] ^ n[51622];
assign t[51623] = t[51622] ^ n[51623];
assign t[51624] = t[51623] ^ n[51624];
assign t[51625] = t[51624] ^ n[51625];
assign t[51626] = t[51625] ^ n[51626];
assign t[51627] = t[51626] ^ n[51627];
assign t[51628] = t[51627] ^ n[51628];
assign t[51629] = t[51628] ^ n[51629];
assign t[51630] = t[51629] ^ n[51630];
assign t[51631] = t[51630] ^ n[51631];
assign t[51632] = t[51631] ^ n[51632];
assign t[51633] = t[51632] ^ n[51633];
assign t[51634] = t[51633] ^ n[51634];
assign t[51635] = t[51634] ^ n[51635];
assign t[51636] = t[51635] ^ n[51636];
assign t[51637] = t[51636] ^ n[51637];
assign t[51638] = t[51637] ^ n[51638];
assign t[51639] = t[51638] ^ n[51639];
assign t[51640] = t[51639] ^ n[51640];
assign t[51641] = t[51640] ^ n[51641];
assign t[51642] = t[51641] ^ n[51642];
assign t[51643] = t[51642] ^ n[51643];
assign t[51644] = t[51643] ^ n[51644];
assign t[51645] = t[51644] ^ n[51645];
assign t[51646] = t[51645] ^ n[51646];
assign t[51647] = t[51646] ^ n[51647];
assign t[51648] = t[51647] ^ n[51648];
assign t[51649] = t[51648] ^ n[51649];
assign t[51650] = t[51649] ^ n[51650];
assign t[51651] = t[51650] ^ n[51651];
assign t[51652] = t[51651] ^ n[51652];
assign t[51653] = t[51652] ^ n[51653];
assign t[51654] = t[51653] ^ n[51654];
assign t[51655] = t[51654] ^ n[51655];
assign t[51656] = t[51655] ^ n[51656];
assign t[51657] = t[51656] ^ n[51657];
assign t[51658] = t[51657] ^ n[51658];
assign t[51659] = t[51658] ^ n[51659];
assign t[51660] = t[51659] ^ n[51660];
assign t[51661] = t[51660] ^ n[51661];
assign t[51662] = t[51661] ^ n[51662];
assign t[51663] = t[51662] ^ n[51663];
assign t[51664] = t[51663] ^ n[51664];
assign t[51665] = t[51664] ^ n[51665];
assign t[51666] = t[51665] ^ n[51666];
assign t[51667] = t[51666] ^ n[51667];
assign t[51668] = t[51667] ^ n[51668];
assign t[51669] = t[51668] ^ n[51669];
assign t[51670] = t[51669] ^ n[51670];
assign t[51671] = t[51670] ^ n[51671];
assign t[51672] = t[51671] ^ n[51672];
assign t[51673] = t[51672] ^ n[51673];
assign t[51674] = t[51673] ^ n[51674];
assign t[51675] = t[51674] ^ n[51675];
assign t[51676] = t[51675] ^ n[51676];
assign t[51677] = t[51676] ^ n[51677];
assign t[51678] = t[51677] ^ n[51678];
assign t[51679] = t[51678] ^ n[51679];
assign t[51680] = t[51679] ^ n[51680];
assign t[51681] = t[51680] ^ n[51681];
assign t[51682] = t[51681] ^ n[51682];
assign t[51683] = t[51682] ^ n[51683];
assign t[51684] = t[51683] ^ n[51684];
assign t[51685] = t[51684] ^ n[51685];
assign t[51686] = t[51685] ^ n[51686];
assign t[51687] = t[51686] ^ n[51687];
assign t[51688] = t[51687] ^ n[51688];
assign t[51689] = t[51688] ^ n[51689];
assign t[51690] = t[51689] ^ n[51690];
assign t[51691] = t[51690] ^ n[51691];
assign t[51692] = t[51691] ^ n[51692];
assign t[51693] = t[51692] ^ n[51693];
assign t[51694] = t[51693] ^ n[51694];
assign t[51695] = t[51694] ^ n[51695];
assign t[51696] = t[51695] ^ n[51696];
assign t[51697] = t[51696] ^ n[51697];
assign t[51698] = t[51697] ^ n[51698];
assign t[51699] = t[51698] ^ n[51699];
assign t[51700] = t[51699] ^ n[51700];
assign t[51701] = t[51700] ^ n[51701];
assign t[51702] = t[51701] ^ n[51702];
assign t[51703] = t[51702] ^ n[51703];
assign t[51704] = t[51703] ^ n[51704];
assign t[51705] = t[51704] ^ n[51705];
assign t[51706] = t[51705] ^ n[51706];
assign t[51707] = t[51706] ^ n[51707];
assign t[51708] = t[51707] ^ n[51708];
assign t[51709] = t[51708] ^ n[51709];
assign t[51710] = t[51709] ^ n[51710];
assign t[51711] = t[51710] ^ n[51711];
assign t[51712] = t[51711] ^ n[51712];
assign t[51713] = t[51712] ^ n[51713];
assign t[51714] = t[51713] ^ n[51714];
assign t[51715] = t[51714] ^ n[51715];
assign t[51716] = t[51715] ^ n[51716];
assign t[51717] = t[51716] ^ n[51717];
assign t[51718] = t[51717] ^ n[51718];
assign t[51719] = t[51718] ^ n[51719];
assign t[51720] = t[51719] ^ n[51720];
assign t[51721] = t[51720] ^ n[51721];
assign t[51722] = t[51721] ^ n[51722];
assign t[51723] = t[51722] ^ n[51723];
assign t[51724] = t[51723] ^ n[51724];
assign t[51725] = t[51724] ^ n[51725];
assign t[51726] = t[51725] ^ n[51726];
assign t[51727] = t[51726] ^ n[51727];
assign t[51728] = t[51727] ^ n[51728];
assign t[51729] = t[51728] ^ n[51729];
assign t[51730] = t[51729] ^ n[51730];
assign t[51731] = t[51730] ^ n[51731];
assign t[51732] = t[51731] ^ n[51732];
assign t[51733] = t[51732] ^ n[51733];
assign t[51734] = t[51733] ^ n[51734];
assign t[51735] = t[51734] ^ n[51735];
assign t[51736] = t[51735] ^ n[51736];
assign t[51737] = t[51736] ^ n[51737];
assign t[51738] = t[51737] ^ n[51738];
assign t[51739] = t[51738] ^ n[51739];
assign t[51740] = t[51739] ^ n[51740];
assign t[51741] = t[51740] ^ n[51741];
assign t[51742] = t[51741] ^ n[51742];
assign t[51743] = t[51742] ^ n[51743];
assign t[51744] = t[51743] ^ n[51744];
assign t[51745] = t[51744] ^ n[51745];
assign t[51746] = t[51745] ^ n[51746];
assign t[51747] = t[51746] ^ n[51747];
assign t[51748] = t[51747] ^ n[51748];
assign t[51749] = t[51748] ^ n[51749];
assign t[51750] = t[51749] ^ n[51750];
assign t[51751] = t[51750] ^ n[51751];
assign t[51752] = t[51751] ^ n[51752];
assign t[51753] = t[51752] ^ n[51753];
assign t[51754] = t[51753] ^ n[51754];
assign t[51755] = t[51754] ^ n[51755];
assign t[51756] = t[51755] ^ n[51756];
assign t[51757] = t[51756] ^ n[51757];
assign t[51758] = t[51757] ^ n[51758];
assign t[51759] = t[51758] ^ n[51759];
assign t[51760] = t[51759] ^ n[51760];
assign t[51761] = t[51760] ^ n[51761];
assign t[51762] = t[51761] ^ n[51762];
assign t[51763] = t[51762] ^ n[51763];
assign t[51764] = t[51763] ^ n[51764];
assign t[51765] = t[51764] ^ n[51765];
assign t[51766] = t[51765] ^ n[51766];
assign t[51767] = t[51766] ^ n[51767];
assign t[51768] = t[51767] ^ n[51768];
assign t[51769] = t[51768] ^ n[51769];
assign t[51770] = t[51769] ^ n[51770];
assign t[51771] = t[51770] ^ n[51771];
assign t[51772] = t[51771] ^ n[51772];
assign t[51773] = t[51772] ^ n[51773];
assign t[51774] = t[51773] ^ n[51774];
assign t[51775] = t[51774] ^ n[51775];
assign t[51776] = t[51775] ^ n[51776];
assign t[51777] = t[51776] ^ n[51777];
assign t[51778] = t[51777] ^ n[51778];
assign t[51779] = t[51778] ^ n[51779];
assign t[51780] = t[51779] ^ n[51780];
assign t[51781] = t[51780] ^ n[51781];
assign t[51782] = t[51781] ^ n[51782];
assign t[51783] = t[51782] ^ n[51783];
assign t[51784] = t[51783] ^ n[51784];
assign t[51785] = t[51784] ^ n[51785];
assign t[51786] = t[51785] ^ n[51786];
assign t[51787] = t[51786] ^ n[51787];
assign t[51788] = t[51787] ^ n[51788];
assign t[51789] = t[51788] ^ n[51789];
assign t[51790] = t[51789] ^ n[51790];
assign t[51791] = t[51790] ^ n[51791];
assign t[51792] = t[51791] ^ n[51792];
assign t[51793] = t[51792] ^ n[51793];
assign t[51794] = t[51793] ^ n[51794];
assign t[51795] = t[51794] ^ n[51795];
assign t[51796] = t[51795] ^ n[51796];
assign t[51797] = t[51796] ^ n[51797];
assign t[51798] = t[51797] ^ n[51798];
assign t[51799] = t[51798] ^ n[51799];
assign t[51800] = t[51799] ^ n[51800];
assign t[51801] = t[51800] ^ n[51801];
assign t[51802] = t[51801] ^ n[51802];
assign t[51803] = t[51802] ^ n[51803];
assign t[51804] = t[51803] ^ n[51804];
assign t[51805] = t[51804] ^ n[51805];
assign t[51806] = t[51805] ^ n[51806];
assign t[51807] = t[51806] ^ n[51807];
assign t[51808] = t[51807] ^ n[51808];
assign t[51809] = t[51808] ^ n[51809];
assign t[51810] = t[51809] ^ n[51810];
assign t[51811] = t[51810] ^ n[51811];
assign t[51812] = t[51811] ^ n[51812];
assign t[51813] = t[51812] ^ n[51813];
assign t[51814] = t[51813] ^ n[51814];
assign t[51815] = t[51814] ^ n[51815];
assign t[51816] = t[51815] ^ n[51816];
assign t[51817] = t[51816] ^ n[51817];
assign t[51818] = t[51817] ^ n[51818];
assign t[51819] = t[51818] ^ n[51819];
assign t[51820] = t[51819] ^ n[51820];
assign t[51821] = t[51820] ^ n[51821];
assign t[51822] = t[51821] ^ n[51822];
assign t[51823] = t[51822] ^ n[51823];
assign t[51824] = t[51823] ^ n[51824];
assign t[51825] = t[51824] ^ n[51825];
assign t[51826] = t[51825] ^ n[51826];
assign t[51827] = t[51826] ^ n[51827];
assign t[51828] = t[51827] ^ n[51828];
assign t[51829] = t[51828] ^ n[51829];
assign t[51830] = t[51829] ^ n[51830];
assign t[51831] = t[51830] ^ n[51831];
assign t[51832] = t[51831] ^ n[51832];
assign t[51833] = t[51832] ^ n[51833];
assign t[51834] = t[51833] ^ n[51834];
assign t[51835] = t[51834] ^ n[51835];
assign t[51836] = t[51835] ^ n[51836];
assign t[51837] = t[51836] ^ n[51837];
assign t[51838] = t[51837] ^ n[51838];
assign t[51839] = t[51838] ^ n[51839];
assign t[51840] = t[51839] ^ n[51840];
assign t[51841] = t[51840] ^ n[51841];
assign t[51842] = t[51841] ^ n[51842];
assign t[51843] = t[51842] ^ n[51843];
assign t[51844] = t[51843] ^ n[51844];
assign t[51845] = t[51844] ^ n[51845];
assign t[51846] = t[51845] ^ n[51846];
assign t[51847] = t[51846] ^ n[51847];
assign t[51848] = t[51847] ^ n[51848];
assign t[51849] = t[51848] ^ n[51849];
assign t[51850] = t[51849] ^ n[51850];
assign t[51851] = t[51850] ^ n[51851];
assign t[51852] = t[51851] ^ n[51852];
assign t[51853] = t[51852] ^ n[51853];
assign t[51854] = t[51853] ^ n[51854];
assign t[51855] = t[51854] ^ n[51855];
assign t[51856] = t[51855] ^ n[51856];
assign t[51857] = t[51856] ^ n[51857];
assign t[51858] = t[51857] ^ n[51858];
assign t[51859] = t[51858] ^ n[51859];
assign t[51860] = t[51859] ^ n[51860];
assign t[51861] = t[51860] ^ n[51861];
assign t[51862] = t[51861] ^ n[51862];
assign t[51863] = t[51862] ^ n[51863];
assign t[51864] = t[51863] ^ n[51864];
assign t[51865] = t[51864] ^ n[51865];
assign t[51866] = t[51865] ^ n[51866];
assign t[51867] = t[51866] ^ n[51867];
assign t[51868] = t[51867] ^ n[51868];
assign t[51869] = t[51868] ^ n[51869];
assign t[51870] = t[51869] ^ n[51870];
assign t[51871] = t[51870] ^ n[51871];
assign t[51872] = t[51871] ^ n[51872];
assign t[51873] = t[51872] ^ n[51873];
assign t[51874] = t[51873] ^ n[51874];
assign t[51875] = t[51874] ^ n[51875];
assign t[51876] = t[51875] ^ n[51876];
assign t[51877] = t[51876] ^ n[51877];
assign t[51878] = t[51877] ^ n[51878];
assign t[51879] = t[51878] ^ n[51879];
assign t[51880] = t[51879] ^ n[51880];
assign t[51881] = t[51880] ^ n[51881];
assign t[51882] = t[51881] ^ n[51882];
assign t[51883] = t[51882] ^ n[51883];
assign t[51884] = t[51883] ^ n[51884];
assign t[51885] = t[51884] ^ n[51885];
assign t[51886] = t[51885] ^ n[51886];
assign t[51887] = t[51886] ^ n[51887];
assign t[51888] = t[51887] ^ n[51888];
assign t[51889] = t[51888] ^ n[51889];
assign t[51890] = t[51889] ^ n[51890];
assign t[51891] = t[51890] ^ n[51891];
assign t[51892] = t[51891] ^ n[51892];
assign t[51893] = t[51892] ^ n[51893];
assign t[51894] = t[51893] ^ n[51894];
assign t[51895] = t[51894] ^ n[51895];
assign t[51896] = t[51895] ^ n[51896];
assign t[51897] = t[51896] ^ n[51897];
assign t[51898] = t[51897] ^ n[51898];
assign t[51899] = t[51898] ^ n[51899];
assign t[51900] = t[51899] ^ n[51900];
assign t[51901] = t[51900] ^ n[51901];
assign t[51902] = t[51901] ^ n[51902];
assign t[51903] = t[51902] ^ n[51903];
assign t[51904] = t[51903] ^ n[51904];
assign t[51905] = t[51904] ^ n[51905];
assign t[51906] = t[51905] ^ n[51906];
assign t[51907] = t[51906] ^ n[51907];
assign t[51908] = t[51907] ^ n[51908];
assign t[51909] = t[51908] ^ n[51909];
assign t[51910] = t[51909] ^ n[51910];
assign t[51911] = t[51910] ^ n[51911];
assign t[51912] = t[51911] ^ n[51912];
assign t[51913] = t[51912] ^ n[51913];
assign t[51914] = t[51913] ^ n[51914];
assign t[51915] = t[51914] ^ n[51915];
assign t[51916] = t[51915] ^ n[51916];
assign t[51917] = t[51916] ^ n[51917];
assign t[51918] = t[51917] ^ n[51918];
assign t[51919] = t[51918] ^ n[51919];
assign t[51920] = t[51919] ^ n[51920];
assign t[51921] = t[51920] ^ n[51921];
assign t[51922] = t[51921] ^ n[51922];
assign t[51923] = t[51922] ^ n[51923];
assign t[51924] = t[51923] ^ n[51924];
assign t[51925] = t[51924] ^ n[51925];
assign t[51926] = t[51925] ^ n[51926];
assign t[51927] = t[51926] ^ n[51927];
assign t[51928] = t[51927] ^ n[51928];
assign t[51929] = t[51928] ^ n[51929];
assign t[51930] = t[51929] ^ n[51930];
assign t[51931] = t[51930] ^ n[51931];
assign t[51932] = t[51931] ^ n[51932];
assign t[51933] = t[51932] ^ n[51933];
assign t[51934] = t[51933] ^ n[51934];
assign t[51935] = t[51934] ^ n[51935];
assign t[51936] = t[51935] ^ n[51936];
assign t[51937] = t[51936] ^ n[51937];
assign t[51938] = t[51937] ^ n[51938];
assign t[51939] = t[51938] ^ n[51939];
assign t[51940] = t[51939] ^ n[51940];
assign t[51941] = t[51940] ^ n[51941];
assign t[51942] = t[51941] ^ n[51942];
assign t[51943] = t[51942] ^ n[51943];
assign t[51944] = t[51943] ^ n[51944];
assign t[51945] = t[51944] ^ n[51945];
assign t[51946] = t[51945] ^ n[51946];
assign t[51947] = t[51946] ^ n[51947];
assign t[51948] = t[51947] ^ n[51948];
assign t[51949] = t[51948] ^ n[51949];
assign t[51950] = t[51949] ^ n[51950];
assign t[51951] = t[51950] ^ n[51951];
assign t[51952] = t[51951] ^ n[51952];
assign t[51953] = t[51952] ^ n[51953];
assign t[51954] = t[51953] ^ n[51954];
assign t[51955] = t[51954] ^ n[51955];
assign t[51956] = t[51955] ^ n[51956];
assign t[51957] = t[51956] ^ n[51957];
assign t[51958] = t[51957] ^ n[51958];
assign t[51959] = t[51958] ^ n[51959];
assign t[51960] = t[51959] ^ n[51960];
assign t[51961] = t[51960] ^ n[51961];
assign t[51962] = t[51961] ^ n[51962];
assign t[51963] = t[51962] ^ n[51963];
assign t[51964] = t[51963] ^ n[51964];
assign t[51965] = t[51964] ^ n[51965];
assign t[51966] = t[51965] ^ n[51966];
assign t[51967] = t[51966] ^ n[51967];
assign t[51968] = t[51967] ^ n[51968];
assign t[51969] = t[51968] ^ n[51969];
assign t[51970] = t[51969] ^ n[51970];
assign t[51971] = t[51970] ^ n[51971];
assign t[51972] = t[51971] ^ n[51972];
assign t[51973] = t[51972] ^ n[51973];
assign t[51974] = t[51973] ^ n[51974];
assign t[51975] = t[51974] ^ n[51975];
assign t[51976] = t[51975] ^ n[51976];
assign t[51977] = t[51976] ^ n[51977];
assign t[51978] = t[51977] ^ n[51978];
assign t[51979] = t[51978] ^ n[51979];
assign t[51980] = t[51979] ^ n[51980];
assign t[51981] = t[51980] ^ n[51981];
assign t[51982] = t[51981] ^ n[51982];
assign t[51983] = t[51982] ^ n[51983];
assign t[51984] = t[51983] ^ n[51984];
assign t[51985] = t[51984] ^ n[51985];
assign t[51986] = t[51985] ^ n[51986];
assign t[51987] = t[51986] ^ n[51987];
assign t[51988] = t[51987] ^ n[51988];
assign t[51989] = t[51988] ^ n[51989];
assign t[51990] = t[51989] ^ n[51990];
assign t[51991] = t[51990] ^ n[51991];
assign t[51992] = t[51991] ^ n[51992];
assign t[51993] = t[51992] ^ n[51993];
assign t[51994] = t[51993] ^ n[51994];
assign t[51995] = t[51994] ^ n[51995];
assign t[51996] = t[51995] ^ n[51996];
assign t[51997] = t[51996] ^ n[51997];
assign t[51998] = t[51997] ^ n[51998];
assign t[51999] = t[51998] ^ n[51999];
assign t[52000] = t[51999] ^ n[52000];
assign t[52001] = t[52000] ^ n[52001];
assign t[52002] = t[52001] ^ n[52002];
assign t[52003] = t[52002] ^ n[52003];
assign t[52004] = t[52003] ^ n[52004];
assign t[52005] = t[52004] ^ n[52005];
assign t[52006] = t[52005] ^ n[52006];
assign t[52007] = t[52006] ^ n[52007];
assign t[52008] = t[52007] ^ n[52008];
assign t[52009] = t[52008] ^ n[52009];
assign t[52010] = t[52009] ^ n[52010];
assign t[52011] = t[52010] ^ n[52011];
assign t[52012] = t[52011] ^ n[52012];
assign t[52013] = t[52012] ^ n[52013];
assign t[52014] = t[52013] ^ n[52014];
assign t[52015] = t[52014] ^ n[52015];
assign t[52016] = t[52015] ^ n[52016];
assign t[52017] = t[52016] ^ n[52017];
assign t[52018] = t[52017] ^ n[52018];
assign t[52019] = t[52018] ^ n[52019];
assign t[52020] = t[52019] ^ n[52020];
assign t[52021] = t[52020] ^ n[52021];
assign t[52022] = t[52021] ^ n[52022];
assign t[52023] = t[52022] ^ n[52023];
assign t[52024] = t[52023] ^ n[52024];
assign t[52025] = t[52024] ^ n[52025];
assign t[52026] = t[52025] ^ n[52026];
assign t[52027] = t[52026] ^ n[52027];
assign t[52028] = t[52027] ^ n[52028];
assign t[52029] = t[52028] ^ n[52029];
assign t[52030] = t[52029] ^ n[52030];
assign t[52031] = t[52030] ^ n[52031];
assign t[52032] = t[52031] ^ n[52032];
assign t[52033] = t[52032] ^ n[52033];
assign t[52034] = t[52033] ^ n[52034];
assign t[52035] = t[52034] ^ n[52035];
assign t[52036] = t[52035] ^ n[52036];
assign t[52037] = t[52036] ^ n[52037];
assign t[52038] = t[52037] ^ n[52038];
assign t[52039] = t[52038] ^ n[52039];
assign t[52040] = t[52039] ^ n[52040];
assign t[52041] = t[52040] ^ n[52041];
assign t[52042] = t[52041] ^ n[52042];
assign t[52043] = t[52042] ^ n[52043];
assign t[52044] = t[52043] ^ n[52044];
assign t[52045] = t[52044] ^ n[52045];
assign t[52046] = t[52045] ^ n[52046];
assign t[52047] = t[52046] ^ n[52047];
assign t[52048] = t[52047] ^ n[52048];
assign t[52049] = t[52048] ^ n[52049];
assign t[52050] = t[52049] ^ n[52050];
assign t[52051] = t[52050] ^ n[52051];
assign t[52052] = t[52051] ^ n[52052];
assign t[52053] = t[52052] ^ n[52053];
assign t[52054] = t[52053] ^ n[52054];
assign t[52055] = t[52054] ^ n[52055];
assign t[52056] = t[52055] ^ n[52056];
assign t[52057] = t[52056] ^ n[52057];
assign t[52058] = t[52057] ^ n[52058];
assign t[52059] = t[52058] ^ n[52059];
assign t[52060] = t[52059] ^ n[52060];
assign t[52061] = t[52060] ^ n[52061];
assign t[52062] = t[52061] ^ n[52062];
assign t[52063] = t[52062] ^ n[52063];
assign t[52064] = t[52063] ^ n[52064];
assign t[52065] = t[52064] ^ n[52065];
assign t[52066] = t[52065] ^ n[52066];
assign t[52067] = t[52066] ^ n[52067];
assign t[52068] = t[52067] ^ n[52068];
assign t[52069] = t[52068] ^ n[52069];
assign t[52070] = t[52069] ^ n[52070];
assign t[52071] = t[52070] ^ n[52071];
assign t[52072] = t[52071] ^ n[52072];
assign t[52073] = t[52072] ^ n[52073];
assign t[52074] = t[52073] ^ n[52074];
assign t[52075] = t[52074] ^ n[52075];
assign t[52076] = t[52075] ^ n[52076];
assign t[52077] = t[52076] ^ n[52077];
assign t[52078] = t[52077] ^ n[52078];
assign t[52079] = t[52078] ^ n[52079];
assign t[52080] = t[52079] ^ n[52080];
assign t[52081] = t[52080] ^ n[52081];
assign t[52082] = t[52081] ^ n[52082];
assign t[52083] = t[52082] ^ n[52083];
assign t[52084] = t[52083] ^ n[52084];
assign t[52085] = t[52084] ^ n[52085];
assign t[52086] = t[52085] ^ n[52086];
assign t[52087] = t[52086] ^ n[52087];
assign t[52088] = t[52087] ^ n[52088];
assign t[52089] = t[52088] ^ n[52089];
assign t[52090] = t[52089] ^ n[52090];
assign t[52091] = t[52090] ^ n[52091];
assign t[52092] = t[52091] ^ n[52092];
assign t[52093] = t[52092] ^ n[52093];
assign t[52094] = t[52093] ^ n[52094];
assign t[52095] = t[52094] ^ n[52095];
assign t[52096] = t[52095] ^ n[52096];
assign t[52097] = t[52096] ^ n[52097];
assign t[52098] = t[52097] ^ n[52098];
assign t[52099] = t[52098] ^ n[52099];
assign t[52100] = t[52099] ^ n[52100];
assign t[52101] = t[52100] ^ n[52101];
assign t[52102] = t[52101] ^ n[52102];
assign t[52103] = t[52102] ^ n[52103];
assign t[52104] = t[52103] ^ n[52104];
assign t[52105] = t[52104] ^ n[52105];
assign t[52106] = t[52105] ^ n[52106];
assign t[52107] = t[52106] ^ n[52107];
assign t[52108] = t[52107] ^ n[52108];
assign t[52109] = t[52108] ^ n[52109];
assign t[52110] = t[52109] ^ n[52110];
assign t[52111] = t[52110] ^ n[52111];
assign t[52112] = t[52111] ^ n[52112];
assign t[52113] = t[52112] ^ n[52113];
assign t[52114] = t[52113] ^ n[52114];
assign t[52115] = t[52114] ^ n[52115];
assign t[52116] = t[52115] ^ n[52116];
assign t[52117] = t[52116] ^ n[52117];
assign t[52118] = t[52117] ^ n[52118];
assign t[52119] = t[52118] ^ n[52119];
assign t[52120] = t[52119] ^ n[52120];
assign t[52121] = t[52120] ^ n[52121];
assign t[52122] = t[52121] ^ n[52122];
assign t[52123] = t[52122] ^ n[52123];
assign t[52124] = t[52123] ^ n[52124];
assign t[52125] = t[52124] ^ n[52125];
assign t[52126] = t[52125] ^ n[52126];
assign t[52127] = t[52126] ^ n[52127];
assign t[52128] = t[52127] ^ n[52128];
assign t[52129] = t[52128] ^ n[52129];
assign t[52130] = t[52129] ^ n[52130];
assign t[52131] = t[52130] ^ n[52131];
assign t[52132] = t[52131] ^ n[52132];
assign t[52133] = t[52132] ^ n[52133];
assign t[52134] = t[52133] ^ n[52134];
assign t[52135] = t[52134] ^ n[52135];
assign t[52136] = t[52135] ^ n[52136];
assign t[52137] = t[52136] ^ n[52137];
assign t[52138] = t[52137] ^ n[52138];
assign t[52139] = t[52138] ^ n[52139];
assign t[52140] = t[52139] ^ n[52140];
assign t[52141] = t[52140] ^ n[52141];
assign t[52142] = t[52141] ^ n[52142];
assign t[52143] = t[52142] ^ n[52143];
assign t[52144] = t[52143] ^ n[52144];
assign t[52145] = t[52144] ^ n[52145];
assign t[52146] = t[52145] ^ n[52146];
assign t[52147] = t[52146] ^ n[52147];
assign t[52148] = t[52147] ^ n[52148];
assign t[52149] = t[52148] ^ n[52149];
assign t[52150] = t[52149] ^ n[52150];
assign t[52151] = t[52150] ^ n[52151];
assign t[52152] = t[52151] ^ n[52152];
assign t[52153] = t[52152] ^ n[52153];
assign t[52154] = t[52153] ^ n[52154];
assign t[52155] = t[52154] ^ n[52155];
assign t[52156] = t[52155] ^ n[52156];
assign t[52157] = t[52156] ^ n[52157];
assign t[52158] = t[52157] ^ n[52158];
assign t[52159] = t[52158] ^ n[52159];
assign t[52160] = t[52159] ^ n[52160];
assign t[52161] = t[52160] ^ n[52161];
assign t[52162] = t[52161] ^ n[52162];
assign t[52163] = t[52162] ^ n[52163];
assign t[52164] = t[52163] ^ n[52164];
assign t[52165] = t[52164] ^ n[52165];
assign t[52166] = t[52165] ^ n[52166];
assign t[52167] = t[52166] ^ n[52167];
assign t[52168] = t[52167] ^ n[52168];
assign t[52169] = t[52168] ^ n[52169];
assign t[52170] = t[52169] ^ n[52170];
assign t[52171] = t[52170] ^ n[52171];
assign t[52172] = t[52171] ^ n[52172];
assign t[52173] = t[52172] ^ n[52173];
assign t[52174] = t[52173] ^ n[52174];
assign t[52175] = t[52174] ^ n[52175];
assign t[52176] = t[52175] ^ n[52176];
assign t[52177] = t[52176] ^ n[52177];
assign t[52178] = t[52177] ^ n[52178];
assign t[52179] = t[52178] ^ n[52179];
assign t[52180] = t[52179] ^ n[52180];
assign t[52181] = t[52180] ^ n[52181];
assign t[52182] = t[52181] ^ n[52182];
assign t[52183] = t[52182] ^ n[52183];
assign t[52184] = t[52183] ^ n[52184];
assign t[52185] = t[52184] ^ n[52185];
assign t[52186] = t[52185] ^ n[52186];
assign t[52187] = t[52186] ^ n[52187];
assign t[52188] = t[52187] ^ n[52188];
assign t[52189] = t[52188] ^ n[52189];
assign t[52190] = t[52189] ^ n[52190];
assign t[52191] = t[52190] ^ n[52191];
assign t[52192] = t[52191] ^ n[52192];
assign t[52193] = t[52192] ^ n[52193];
assign t[52194] = t[52193] ^ n[52194];
assign t[52195] = t[52194] ^ n[52195];
assign t[52196] = t[52195] ^ n[52196];
assign t[52197] = t[52196] ^ n[52197];
assign t[52198] = t[52197] ^ n[52198];
assign t[52199] = t[52198] ^ n[52199];
assign t[52200] = t[52199] ^ n[52200];
assign t[52201] = t[52200] ^ n[52201];
assign t[52202] = t[52201] ^ n[52202];
assign t[52203] = t[52202] ^ n[52203];
assign t[52204] = t[52203] ^ n[52204];
assign t[52205] = t[52204] ^ n[52205];
assign t[52206] = t[52205] ^ n[52206];
assign t[52207] = t[52206] ^ n[52207];
assign t[52208] = t[52207] ^ n[52208];
assign t[52209] = t[52208] ^ n[52209];
assign t[52210] = t[52209] ^ n[52210];
assign t[52211] = t[52210] ^ n[52211];
assign t[52212] = t[52211] ^ n[52212];
assign t[52213] = t[52212] ^ n[52213];
assign t[52214] = t[52213] ^ n[52214];
assign t[52215] = t[52214] ^ n[52215];
assign t[52216] = t[52215] ^ n[52216];
assign t[52217] = t[52216] ^ n[52217];
assign t[52218] = t[52217] ^ n[52218];
assign t[52219] = t[52218] ^ n[52219];
assign t[52220] = t[52219] ^ n[52220];
assign t[52221] = t[52220] ^ n[52221];
assign t[52222] = t[52221] ^ n[52222];
assign t[52223] = t[52222] ^ n[52223];
assign t[52224] = t[52223] ^ n[52224];
assign t[52225] = t[52224] ^ n[52225];
assign t[52226] = t[52225] ^ n[52226];
assign t[52227] = t[52226] ^ n[52227];
assign t[52228] = t[52227] ^ n[52228];
assign t[52229] = t[52228] ^ n[52229];
assign t[52230] = t[52229] ^ n[52230];
assign t[52231] = t[52230] ^ n[52231];
assign t[52232] = t[52231] ^ n[52232];
assign t[52233] = t[52232] ^ n[52233];
assign t[52234] = t[52233] ^ n[52234];
assign t[52235] = t[52234] ^ n[52235];
assign t[52236] = t[52235] ^ n[52236];
assign t[52237] = t[52236] ^ n[52237];
assign t[52238] = t[52237] ^ n[52238];
assign t[52239] = t[52238] ^ n[52239];
assign t[52240] = t[52239] ^ n[52240];
assign t[52241] = t[52240] ^ n[52241];
assign t[52242] = t[52241] ^ n[52242];
assign t[52243] = t[52242] ^ n[52243];
assign t[52244] = t[52243] ^ n[52244];
assign t[52245] = t[52244] ^ n[52245];
assign t[52246] = t[52245] ^ n[52246];
assign t[52247] = t[52246] ^ n[52247];
assign t[52248] = t[52247] ^ n[52248];
assign t[52249] = t[52248] ^ n[52249];
assign t[52250] = t[52249] ^ n[52250];
assign t[52251] = t[52250] ^ n[52251];
assign t[52252] = t[52251] ^ n[52252];
assign t[52253] = t[52252] ^ n[52253];
assign t[52254] = t[52253] ^ n[52254];
assign t[52255] = t[52254] ^ n[52255];
assign t[52256] = t[52255] ^ n[52256];
assign t[52257] = t[52256] ^ n[52257];
assign t[52258] = t[52257] ^ n[52258];
assign t[52259] = t[52258] ^ n[52259];
assign t[52260] = t[52259] ^ n[52260];
assign t[52261] = t[52260] ^ n[52261];
assign t[52262] = t[52261] ^ n[52262];
assign t[52263] = t[52262] ^ n[52263];
assign t[52264] = t[52263] ^ n[52264];
assign t[52265] = t[52264] ^ n[52265];
assign t[52266] = t[52265] ^ n[52266];
assign t[52267] = t[52266] ^ n[52267];
assign t[52268] = t[52267] ^ n[52268];
assign t[52269] = t[52268] ^ n[52269];
assign t[52270] = t[52269] ^ n[52270];
assign t[52271] = t[52270] ^ n[52271];
assign t[52272] = t[52271] ^ n[52272];
assign t[52273] = t[52272] ^ n[52273];
assign t[52274] = t[52273] ^ n[52274];
assign t[52275] = t[52274] ^ n[52275];
assign t[52276] = t[52275] ^ n[52276];
assign t[52277] = t[52276] ^ n[52277];
assign t[52278] = t[52277] ^ n[52278];
assign t[52279] = t[52278] ^ n[52279];
assign t[52280] = t[52279] ^ n[52280];
assign t[52281] = t[52280] ^ n[52281];
assign t[52282] = t[52281] ^ n[52282];
assign t[52283] = t[52282] ^ n[52283];
assign t[52284] = t[52283] ^ n[52284];
assign t[52285] = t[52284] ^ n[52285];
assign t[52286] = t[52285] ^ n[52286];
assign t[52287] = t[52286] ^ n[52287];
assign t[52288] = t[52287] ^ n[52288];
assign t[52289] = t[52288] ^ n[52289];
assign t[52290] = t[52289] ^ n[52290];
assign t[52291] = t[52290] ^ n[52291];
assign t[52292] = t[52291] ^ n[52292];
assign t[52293] = t[52292] ^ n[52293];
assign t[52294] = t[52293] ^ n[52294];
assign t[52295] = t[52294] ^ n[52295];
assign t[52296] = t[52295] ^ n[52296];
assign t[52297] = t[52296] ^ n[52297];
assign t[52298] = t[52297] ^ n[52298];
assign t[52299] = t[52298] ^ n[52299];
assign t[52300] = t[52299] ^ n[52300];
assign t[52301] = t[52300] ^ n[52301];
assign t[52302] = t[52301] ^ n[52302];
assign t[52303] = t[52302] ^ n[52303];
assign t[52304] = t[52303] ^ n[52304];
assign t[52305] = t[52304] ^ n[52305];
assign t[52306] = t[52305] ^ n[52306];
assign t[52307] = t[52306] ^ n[52307];
assign t[52308] = t[52307] ^ n[52308];
assign t[52309] = t[52308] ^ n[52309];
assign t[52310] = t[52309] ^ n[52310];
assign t[52311] = t[52310] ^ n[52311];
assign t[52312] = t[52311] ^ n[52312];
assign t[52313] = t[52312] ^ n[52313];
assign t[52314] = t[52313] ^ n[52314];
assign t[52315] = t[52314] ^ n[52315];
assign t[52316] = t[52315] ^ n[52316];
assign t[52317] = t[52316] ^ n[52317];
assign t[52318] = t[52317] ^ n[52318];
assign t[52319] = t[52318] ^ n[52319];
assign t[52320] = t[52319] ^ n[52320];
assign t[52321] = t[52320] ^ n[52321];
assign t[52322] = t[52321] ^ n[52322];
assign t[52323] = t[52322] ^ n[52323];
assign t[52324] = t[52323] ^ n[52324];
assign t[52325] = t[52324] ^ n[52325];
assign t[52326] = t[52325] ^ n[52326];
assign t[52327] = t[52326] ^ n[52327];
assign t[52328] = t[52327] ^ n[52328];
assign t[52329] = t[52328] ^ n[52329];
assign t[52330] = t[52329] ^ n[52330];
assign t[52331] = t[52330] ^ n[52331];
assign t[52332] = t[52331] ^ n[52332];
assign t[52333] = t[52332] ^ n[52333];
assign t[52334] = t[52333] ^ n[52334];
assign t[52335] = t[52334] ^ n[52335];
assign t[52336] = t[52335] ^ n[52336];
assign t[52337] = t[52336] ^ n[52337];
assign t[52338] = t[52337] ^ n[52338];
assign t[52339] = t[52338] ^ n[52339];
assign t[52340] = t[52339] ^ n[52340];
assign t[52341] = t[52340] ^ n[52341];
assign t[52342] = t[52341] ^ n[52342];
assign t[52343] = t[52342] ^ n[52343];
assign t[52344] = t[52343] ^ n[52344];
assign t[52345] = t[52344] ^ n[52345];
assign t[52346] = t[52345] ^ n[52346];
assign t[52347] = t[52346] ^ n[52347];
assign t[52348] = t[52347] ^ n[52348];
assign t[52349] = t[52348] ^ n[52349];
assign t[52350] = t[52349] ^ n[52350];
assign t[52351] = t[52350] ^ n[52351];
assign t[52352] = t[52351] ^ n[52352];
assign t[52353] = t[52352] ^ n[52353];
assign t[52354] = t[52353] ^ n[52354];
assign t[52355] = t[52354] ^ n[52355];
assign t[52356] = t[52355] ^ n[52356];
assign t[52357] = t[52356] ^ n[52357];
assign t[52358] = t[52357] ^ n[52358];
assign t[52359] = t[52358] ^ n[52359];
assign t[52360] = t[52359] ^ n[52360];
assign t[52361] = t[52360] ^ n[52361];
assign t[52362] = t[52361] ^ n[52362];
assign t[52363] = t[52362] ^ n[52363];
assign t[52364] = t[52363] ^ n[52364];
assign t[52365] = t[52364] ^ n[52365];
assign t[52366] = t[52365] ^ n[52366];
assign t[52367] = t[52366] ^ n[52367];
assign t[52368] = t[52367] ^ n[52368];
assign t[52369] = t[52368] ^ n[52369];
assign t[52370] = t[52369] ^ n[52370];
assign t[52371] = t[52370] ^ n[52371];
assign t[52372] = t[52371] ^ n[52372];
assign t[52373] = t[52372] ^ n[52373];
assign t[52374] = t[52373] ^ n[52374];
assign t[52375] = t[52374] ^ n[52375];
assign t[52376] = t[52375] ^ n[52376];
assign t[52377] = t[52376] ^ n[52377];
assign t[52378] = t[52377] ^ n[52378];
assign t[52379] = t[52378] ^ n[52379];
assign t[52380] = t[52379] ^ n[52380];
assign t[52381] = t[52380] ^ n[52381];
assign t[52382] = t[52381] ^ n[52382];
assign t[52383] = t[52382] ^ n[52383];
assign t[52384] = t[52383] ^ n[52384];
assign t[52385] = t[52384] ^ n[52385];
assign t[52386] = t[52385] ^ n[52386];
assign t[52387] = t[52386] ^ n[52387];
assign t[52388] = t[52387] ^ n[52388];
assign t[52389] = t[52388] ^ n[52389];
assign t[52390] = t[52389] ^ n[52390];
assign t[52391] = t[52390] ^ n[52391];
assign t[52392] = t[52391] ^ n[52392];
assign t[52393] = t[52392] ^ n[52393];
assign t[52394] = t[52393] ^ n[52394];
assign t[52395] = t[52394] ^ n[52395];
assign t[52396] = t[52395] ^ n[52396];
assign t[52397] = t[52396] ^ n[52397];
assign t[52398] = t[52397] ^ n[52398];
assign t[52399] = t[52398] ^ n[52399];
assign t[52400] = t[52399] ^ n[52400];
assign t[52401] = t[52400] ^ n[52401];
assign t[52402] = t[52401] ^ n[52402];
assign t[52403] = t[52402] ^ n[52403];
assign t[52404] = t[52403] ^ n[52404];
assign t[52405] = t[52404] ^ n[52405];
assign t[52406] = t[52405] ^ n[52406];
assign t[52407] = t[52406] ^ n[52407];
assign t[52408] = t[52407] ^ n[52408];
assign t[52409] = t[52408] ^ n[52409];
assign t[52410] = t[52409] ^ n[52410];
assign t[52411] = t[52410] ^ n[52411];
assign t[52412] = t[52411] ^ n[52412];
assign t[52413] = t[52412] ^ n[52413];
assign t[52414] = t[52413] ^ n[52414];
assign t[52415] = t[52414] ^ n[52415];
assign t[52416] = t[52415] ^ n[52416];
assign t[52417] = t[52416] ^ n[52417];
assign t[52418] = t[52417] ^ n[52418];
assign t[52419] = t[52418] ^ n[52419];
assign t[52420] = t[52419] ^ n[52420];
assign t[52421] = t[52420] ^ n[52421];
assign t[52422] = t[52421] ^ n[52422];
assign t[52423] = t[52422] ^ n[52423];
assign t[52424] = t[52423] ^ n[52424];
assign t[52425] = t[52424] ^ n[52425];
assign t[52426] = t[52425] ^ n[52426];
assign t[52427] = t[52426] ^ n[52427];
assign t[52428] = t[52427] ^ n[52428];
assign t[52429] = t[52428] ^ n[52429];
assign t[52430] = t[52429] ^ n[52430];
assign t[52431] = t[52430] ^ n[52431];
assign t[52432] = t[52431] ^ n[52432];
assign t[52433] = t[52432] ^ n[52433];
assign t[52434] = t[52433] ^ n[52434];
assign t[52435] = t[52434] ^ n[52435];
assign t[52436] = t[52435] ^ n[52436];
assign t[52437] = t[52436] ^ n[52437];
assign t[52438] = t[52437] ^ n[52438];
assign t[52439] = t[52438] ^ n[52439];
assign t[52440] = t[52439] ^ n[52440];
assign t[52441] = t[52440] ^ n[52441];
assign t[52442] = t[52441] ^ n[52442];
assign t[52443] = t[52442] ^ n[52443];
assign t[52444] = t[52443] ^ n[52444];
assign t[52445] = t[52444] ^ n[52445];
assign t[52446] = t[52445] ^ n[52446];
assign t[52447] = t[52446] ^ n[52447];
assign t[52448] = t[52447] ^ n[52448];
assign t[52449] = t[52448] ^ n[52449];
assign t[52450] = t[52449] ^ n[52450];
assign t[52451] = t[52450] ^ n[52451];
assign t[52452] = t[52451] ^ n[52452];
assign t[52453] = t[52452] ^ n[52453];
assign t[52454] = t[52453] ^ n[52454];
assign t[52455] = t[52454] ^ n[52455];
assign t[52456] = t[52455] ^ n[52456];
assign t[52457] = t[52456] ^ n[52457];
assign t[52458] = t[52457] ^ n[52458];
assign t[52459] = t[52458] ^ n[52459];
assign t[52460] = t[52459] ^ n[52460];
assign t[52461] = t[52460] ^ n[52461];
assign t[52462] = t[52461] ^ n[52462];
assign t[52463] = t[52462] ^ n[52463];
assign t[52464] = t[52463] ^ n[52464];
assign t[52465] = t[52464] ^ n[52465];
assign t[52466] = t[52465] ^ n[52466];
assign t[52467] = t[52466] ^ n[52467];
assign t[52468] = t[52467] ^ n[52468];
assign t[52469] = t[52468] ^ n[52469];
assign t[52470] = t[52469] ^ n[52470];
assign t[52471] = t[52470] ^ n[52471];
assign t[52472] = t[52471] ^ n[52472];
assign t[52473] = t[52472] ^ n[52473];
assign t[52474] = t[52473] ^ n[52474];
assign t[52475] = t[52474] ^ n[52475];
assign t[52476] = t[52475] ^ n[52476];
assign t[52477] = t[52476] ^ n[52477];
assign t[52478] = t[52477] ^ n[52478];
assign t[52479] = t[52478] ^ n[52479];
assign t[52480] = t[52479] ^ n[52480];
assign t[52481] = t[52480] ^ n[52481];
assign t[52482] = t[52481] ^ n[52482];
assign t[52483] = t[52482] ^ n[52483];
assign t[52484] = t[52483] ^ n[52484];
assign t[52485] = t[52484] ^ n[52485];
assign t[52486] = t[52485] ^ n[52486];
assign t[52487] = t[52486] ^ n[52487];
assign t[52488] = t[52487] ^ n[52488];
assign t[52489] = t[52488] ^ n[52489];
assign t[52490] = t[52489] ^ n[52490];
assign t[52491] = t[52490] ^ n[52491];
assign t[52492] = t[52491] ^ n[52492];
assign t[52493] = t[52492] ^ n[52493];
assign t[52494] = t[52493] ^ n[52494];
assign t[52495] = t[52494] ^ n[52495];
assign t[52496] = t[52495] ^ n[52496];
assign t[52497] = t[52496] ^ n[52497];
assign t[52498] = t[52497] ^ n[52498];
assign t[52499] = t[52498] ^ n[52499];
assign t[52500] = t[52499] ^ n[52500];
assign t[52501] = t[52500] ^ n[52501];
assign t[52502] = t[52501] ^ n[52502];
assign t[52503] = t[52502] ^ n[52503];
assign t[52504] = t[52503] ^ n[52504];
assign t[52505] = t[52504] ^ n[52505];
assign t[52506] = t[52505] ^ n[52506];
assign t[52507] = t[52506] ^ n[52507];
assign t[52508] = t[52507] ^ n[52508];
assign t[52509] = t[52508] ^ n[52509];
assign t[52510] = t[52509] ^ n[52510];
assign t[52511] = t[52510] ^ n[52511];
assign t[52512] = t[52511] ^ n[52512];
assign t[52513] = t[52512] ^ n[52513];
assign t[52514] = t[52513] ^ n[52514];
assign t[52515] = t[52514] ^ n[52515];
assign t[52516] = t[52515] ^ n[52516];
assign t[52517] = t[52516] ^ n[52517];
assign t[52518] = t[52517] ^ n[52518];
assign t[52519] = t[52518] ^ n[52519];
assign t[52520] = t[52519] ^ n[52520];
assign t[52521] = t[52520] ^ n[52521];
assign t[52522] = t[52521] ^ n[52522];
assign t[52523] = t[52522] ^ n[52523];
assign t[52524] = t[52523] ^ n[52524];
assign t[52525] = t[52524] ^ n[52525];
assign t[52526] = t[52525] ^ n[52526];
assign t[52527] = t[52526] ^ n[52527];
assign t[52528] = t[52527] ^ n[52528];
assign t[52529] = t[52528] ^ n[52529];
assign t[52530] = t[52529] ^ n[52530];
assign t[52531] = t[52530] ^ n[52531];
assign t[52532] = t[52531] ^ n[52532];
assign t[52533] = t[52532] ^ n[52533];
assign t[52534] = t[52533] ^ n[52534];
assign t[52535] = t[52534] ^ n[52535];
assign t[52536] = t[52535] ^ n[52536];
assign t[52537] = t[52536] ^ n[52537];
assign t[52538] = t[52537] ^ n[52538];
assign t[52539] = t[52538] ^ n[52539];
assign t[52540] = t[52539] ^ n[52540];
assign t[52541] = t[52540] ^ n[52541];
assign t[52542] = t[52541] ^ n[52542];
assign t[52543] = t[52542] ^ n[52543];
assign t[52544] = t[52543] ^ n[52544];
assign t[52545] = t[52544] ^ n[52545];
assign t[52546] = t[52545] ^ n[52546];
assign t[52547] = t[52546] ^ n[52547];
assign t[52548] = t[52547] ^ n[52548];
assign t[52549] = t[52548] ^ n[52549];
assign t[52550] = t[52549] ^ n[52550];
assign t[52551] = t[52550] ^ n[52551];
assign t[52552] = t[52551] ^ n[52552];
assign t[52553] = t[52552] ^ n[52553];
assign t[52554] = t[52553] ^ n[52554];
assign t[52555] = t[52554] ^ n[52555];
assign t[52556] = t[52555] ^ n[52556];
assign t[52557] = t[52556] ^ n[52557];
assign t[52558] = t[52557] ^ n[52558];
assign t[52559] = t[52558] ^ n[52559];
assign t[52560] = t[52559] ^ n[52560];
assign t[52561] = t[52560] ^ n[52561];
assign t[52562] = t[52561] ^ n[52562];
assign t[52563] = t[52562] ^ n[52563];
assign t[52564] = t[52563] ^ n[52564];
assign t[52565] = t[52564] ^ n[52565];
assign t[52566] = t[52565] ^ n[52566];
assign t[52567] = t[52566] ^ n[52567];
assign t[52568] = t[52567] ^ n[52568];
assign t[52569] = t[52568] ^ n[52569];
assign t[52570] = t[52569] ^ n[52570];
assign t[52571] = t[52570] ^ n[52571];
assign t[52572] = t[52571] ^ n[52572];
assign t[52573] = t[52572] ^ n[52573];
assign t[52574] = t[52573] ^ n[52574];
assign t[52575] = t[52574] ^ n[52575];
assign t[52576] = t[52575] ^ n[52576];
assign t[52577] = t[52576] ^ n[52577];
assign t[52578] = t[52577] ^ n[52578];
assign t[52579] = t[52578] ^ n[52579];
assign t[52580] = t[52579] ^ n[52580];
assign t[52581] = t[52580] ^ n[52581];
assign t[52582] = t[52581] ^ n[52582];
assign t[52583] = t[52582] ^ n[52583];
assign t[52584] = t[52583] ^ n[52584];
assign t[52585] = t[52584] ^ n[52585];
assign t[52586] = t[52585] ^ n[52586];
assign t[52587] = t[52586] ^ n[52587];
assign t[52588] = t[52587] ^ n[52588];
assign t[52589] = t[52588] ^ n[52589];
assign t[52590] = t[52589] ^ n[52590];
assign t[52591] = t[52590] ^ n[52591];
assign t[52592] = t[52591] ^ n[52592];
assign t[52593] = t[52592] ^ n[52593];
assign t[52594] = t[52593] ^ n[52594];
assign t[52595] = t[52594] ^ n[52595];
assign t[52596] = t[52595] ^ n[52596];
assign t[52597] = t[52596] ^ n[52597];
assign t[52598] = t[52597] ^ n[52598];
assign t[52599] = t[52598] ^ n[52599];
assign t[52600] = t[52599] ^ n[52600];
assign t[52601] = t[52600] ^ n[52601];
assign t[52602] = t[52601] ^ n[52602];
assign t[52603] = t[52602] ^ n[52603];
assign t[52604] = t[52603] ^ n[52604];
assign t[52605] = t[52604] ^ n[52605];
assign t[52606] = t[52605] ^ n[52606];
assign t[52607] = t[52606] ^ n[52607];
assign t[52608] = t[52607] ^ n[52608];
assign t[52609] = t[52608] ^ n[52609];
assign t[52610] = t[52609] ^ n[52610];
assign t[52611] = t[52610] ^ n[52611];
assign t[52612] = t[52611] ^ n[52612];
assign t[52613] = t[52612] ^ n[52613];
assign t[52614] = t[52613] ^ n[52614];
assign t[52615] = t[52614] ^ n[52615];
assign t[52616] = t[52615] ^ n[52616];
assign t[52617] = t[52616] ^ n[52617];
assign t[52618] = t[52617] ^ n[52618];
assign t[52619] = t[52618] ^ n[52619];
assign t[52620] = t[52619] ^ n[52620];
assign t[52621] = t[52620] ^ n[52621];
assign t[52622] = t[52621] ^ n[52622];
assign t[52623] = t[52622] ^ n[52623];
assign t[52624] = t[52623] ^ n[52624];
assign t[52625] = t[52624] ^ n[52625];
assign t[52626] = t[52625] ^ n[52626];
assign t[52627] = t[52626] ^ n[52627];
assign t[52628] = t[52627] ^ n[52628];
assign t[52629] = t[52628] ^ n[52629];
assign t[52630] = t[52629] ^ n[52630];
assign t[52631] = t[52630] ^ n[52631];
assign t[52632] = t[52631] ^ n[52632];
assign t[52633] = t[52632] ^ n[52633];
assign t[52634] = t[52633] ^ n[52634];
assign t[52635] = t[52634] ^ n[52635];
assign t[52636] = t[52635] ^ n[52636];
assign t[52637] = t[52636] ^ n[52637];
assign t[52638] = t[52637] ^ n[52638];
assign t[52639] = t[52638] ^ n[52639];
assign t[52640] = t[52639] ^ n[52640];
assign t[52641] = t[52640] ^ n[52641];
assign t[52642] = t[52641] ^ n[52642];
assign t[52643] = t[52642] ^ n[52643];
assign t[52644] = t[52643] ^ n[52644];
assign t[52645] = t[52644] ^ n[52645];
assign t[52646] = t[52645] ^ n[52646];
assign t[52647] = t[52646] ^ n[52647];
assign t[52648] = t[52647] ^ n[52648];
assign t[52649] = t[52648] ^ n[52649];
assign t[52650] = t[52649] ^ n[52650];
assign t[52651] = t[52650] ^ n[52651];
assign t[52652] = t[52651] ^ n[52652];
assign t[52653] = t[52652] ^ n[52653];
assign t[52654] = t[52653] ^ n[52654];
assign t[52655] = t[52654] ^ n[52655];
assign t[52656] = t[52655] ^ n[52656];
assign t[52657] = t[52656] ^ n[52657];
assign t[52658] = t[52657] ^ n[52658];
assign t[52659] = t[52658] ^ n[52659];
assign t[52660] = t[52659] ^ n[52660];
assign t[52661] = t[52660] ^ n[52661];
assign t[52662] = t[52661] ^ n[52662];
assign t[52663] = t[52662] ^ n[52663];
assign t[52664] = t[52663] ^ n[52664];
assign t[52665] = t[52664] ^ n[52665];
assign t[52666] = t[52665] ^ n[52666];
assign t[52667] = t[52666] ^ n[52667];
assign t[52668] = t[52667] ^ n[52668];
assign t[52669] = t[52668] ^ n[52669];
assign t[52670] = t[52669] ^ n[52670];
assign t[52671] = t[52670] ^ n[52671];
assign t[52672] = t[52671] ^ n[52672];
assign t[52673] = t[52672] ^ n[52673];
assign t[52674] = t[52673] ^ n[52674];
assign t[52675] = t[52674] ^ n[52675];
assign t[52676] = t[52675] ^ n[52676];
assign t[52677] = t[52676] ^ n[52677];
assign t[52678] = t[52677] ^ n[52678];
assign t[52679] = t[52678] ^ n[52679];
assign t[52680] = t[52679] ^ n[52680];
assign t[52681] = t[52680] ^ n[52681];
assign t[52682] = t[52681] ^ n[52682];
assign t[52683] = t[52682] ^ n[52683];
assign t[52684] = t[52683] ^ n[52684];
assign t[52685] = t[52684] ^ n[52685];
assign t[52686] = t[52685] ^ n[52686];
assign t[52687] = t[52686] ^ n[52687];
assign t[52688] = t[52687] ^ n[52688];
assign t[52689] = t[52688] ^ n[52689];
assign t[52690] = t[52689] ^ n[52690];
assign t[52691] = t[52690] ^ n[52691];
assign t[52692] = t[52691] ^ n[52692];
assign t[52693] = t[52692] ^ n[52693];
assign t[52694] = t[52693] ^ n[52694];
assign t[52695] = t[52694] ^ n[52695];
assign t[52696] = t[52695] ^ n[52696];
assign t[52697] = t[52696] ^ n[52697];
assign t[52698] = t[52697] ^ n[52698];
assign t[52699] = t[52698] ^ n[52699];
assign t[52700] = t[52699] ^ n[52700];
assign t[52701] = t[52700] ^ n[52701];
assign t[52702] = t[52701] ^ n[52702];
assign t[52703] = t[52702] ^ n[52703];
assign t[52704] = t[52703] ^ n[52704];
assign t[52705] = t[52704] ^ n[52705];
assign t[52706] = t[52705] ^ n[52706];
assign t[52707] = t[52706] ^ n[52707];
assign t[52708] = t[52707] ^ n[52708];
assign t[52709] = t[52708] ^ n[52709];
assign t[52710] = t[52709] ^ n[52710];
assign t[52711] = t[52710] ^ n[52711];
assign t[52712] = t[52711] ^ n[52712];
assign t[52713] = t[52712] ^ n[52713];
assign t[52714] = t[52713] ^ n[52714];
assign t[52715] = t[52714] ^ n[52715];
assign t[52716] = t[52715] ^ n[52716];
assign t[52717] = t[52716] ^ n[52717];
assign t[52718] = t[52717] ^ n[52718];
assign t[52719] = t[52718] ^ n[52719];
assign t[52720] = t[52719] ^ n[52720];
assign t[52721] = t[52720] ^ n[52721];
assign t[52722] = t[52721] ^ n[52722];
assign t[52723] = t[52722] ^ n[52723];
assign t[52724] = t[52723] ^ n[52724];
assign t[52725] = t[52724] ^ n[52725];
assign t[52726] = t[52725] ^ n[52726];
assign t[52727] = t[52726] ^ n[52727];
assign t[52728] = t[52727] ^ n[52728];
assign t[52729] = t[52728] ^ n[52729];
assign t[52730] = t[52729] ^ n[52730];
assign t[52731] = t[52730] ^ n[52731];
assign t[52732] = t[52731] ^ n[52732];
assign t[52733] = t[52732] ^ n[52733];
assign t[52734] = t[52733] ^ n[52734];
assign t[52735] = t[52734] ^ n[52735];
assign t[52736] = t[52735] ^ n[52736];
assign t[52737] = t[52736] ^ n[52737];
assign t[52738] = t[52737] ^ n[52738];
assign t[52739] = t[52738] ^ n[52739];
assign t[52740] = t[52739] ^ n[52740];
assign t[52741] = t[52740] ^ n[52741];
assign t[52742] = t[52741] ^ n[52742];
assign t[52743] = t[52742] ^ n[52743];
assign t[52744] = t[52743] ^ n[52744];
assign t[52745] = t[52744] ^ n[52745];
assign t[52746] = t[52745] ^ n[52746];
assign t[52747] = t[52746] ^ n[52747];
assign t[52748] = t[52747] ^ n[52748];
assign t[52749] = t[52748] ^ n[52749];
assign t[52750] = t[52749] ^ n[52750];
assign t[52751] = t[52750] ^ n[52751];
assign t[52752] = t[52751] ^ n[52752];
assign t[52753] = t[52752] ^ n[52753];
assign t[52754] = t[52753] ^ n[52754];
assign t[52755] = t[52754] ^ n[52755];
assign t[52756] = t[52755] ^ n[52756];
assign t[52757] = t[52756] ^ n[52757];
assign t[52758] = t[52757] ^ n[52758];
assign t[52759] = t[52758] ^ n[52759];
assign t[52760] = t[52759] ^ n[52760];
assign t[52761] = t[52760] ^ n[52761];
assign t[52762] = t[52761] ^ n[52762];
assign t[52763] = t[52762] ^ n[52763];
assign t[52764] = t[52763] ^ n[52764];
assign t[52765] = t[52764] ^ n[52765];
assign t[52766] = t[52765] ^ n[52766];
assign t[52767] = t[52766] ^ n[52767];
assign t[52768] = t[52767] ^ n[52768];
assign t[52769] = t[52768] ^ n[52769];
assign t[52770] = t[52769] ^ n[52770];
assign t[52771] = t[52770] ^ n[52771];
assign t[52772] = t[52771] ^ n[52772];
assign t[52773] = t[52772] ^ n[52773];
assign t[52774] = t[52773] ^ n[52774];
assign t[52775] = t[52774] ^ n[52775];
assign t[52776] = t[52775] ^ n[52776];
assign t[52777] = t[52776] ^ n[52777];
assign t[52778] = t[52777] ^ n[52778];
assign t[52779] = t[52778] ^ n[52779];
assign t[52780] = t[52779] ^ n[52780];
assign t[52781] = t[52780] ^ n[52781];
assign t[52782] = t[52781] ^ n[52782];
assign t[52783] = t[52782] ^ n[52783];
assign t[52784] = t[52783] ^ n[52784];
assign t[52785] = t[52784] ^ n[52785];
assign t[52786] = t[52785] ^ n[52786];
assign t[52787] = t[52786] ^ n[52787];
assign t[52788] = t[52787] ^ n[52788];
assign t[52789] = t[52788] ^ n[52789];
assign t[52790] = t[52789] ^ n[52790];
assign t[52791] = t[52790] ^ n[52791];
assign t[52792] = t[52791] ^ n[52792];
assign t[52793] = t[52792] ^ n[52793];
assign t[52794] = t[52793] ^ n[52794];
assign t[52795] = t[52794] ^ n[52795];
assign t[52796] = t[52795] ^ n[52796];
assign t[52797] = t[52796] ^ n[52797];
assign t[52798] = t[52797] ^ n[52798];
assign t[52799] = t[52798] ^ n[52799];
assign t[52800] = t[52799] ^ n[52800];
assign t[52801] = t[52800] ^ n[52801];
assign t[52802] = t[52801] ^ n[52802];
assign t[52803] = t[52802] ^ n[52803];
assign t[52804] = t[52803] ^ n[52804];
assign t[52805] = t[52804] ^ n[52805];
assign t[52806] = t[52805] ^ n[52806];
assign t[52807] = t[52806] ^ n[52807];
assign t[52808] = t[52807] ^ n[52808];
assign t[52809] = t[52808] ^ n[52809];
assign t[52810] = t[52809] ^ n[52810];
assign t[52811] = t[52810] ^ n[52811];
assign t[52812] = t[52811] ^ n[52812];
assign t[52813] = t[52812] ^ n[52813];
assign t[52814] = t[52813] ^ n[52814];
assign t[52815] = t[52814] ^ n[52815];
assign t[52816] = t[52815] ^ n[52816];
assign t[52817] = t[52816] ^ n[52817];
assign t[52818] = t[52817] ^ n[52818];
assign t[52819] = t[52818] ^ n[52819];
assign t[52820] = t[52819] ^ n[52820];
assign t[52821] = t[52820] ^ n[52821];
assign t[52822] = t[52821] ^ n[52822];
assign t[52823] = t[52822] ^ n[52823];
assign t[52824] = t[52823] ^ n[52824];
assign t[52825] = t[52824] ^ n[52825];
assign t[52826] = t[52825] ^ n[52826];
assign t[52827] = t[52826] ^ n[52827];
assign t[52828] = t[52827] ^ n[52828];
assign t[52829] = t[52828] ^ n[52829];
assign t[52830] = t[52829] ^ n[52830];
assign t[52831] = t[52830] ^ n[52831];
assign t[52832] = t[52831] ^ n[52832];
assign t[52833] = t[52832] ^ n[52833];
assign t[52834] = t[52833] ^ n[52834];
assign t[52835] = t[52834] ^ n[52835];
assign t[52836] = t[52835] ^ n[52836];
assign t[52837] = t[52836] ^ n[52837];
assign t[52838] = t[52837] ^ n[52838];
assign t[52839] = t[52838] ^ n[52839];
assign t[52840] = t[52839] ^ n[52840];
assign t[52841] = t[52840] ^ n[52841];
assign t[52842] = t[52841] ^ n[52842];
assign t[52843] = t[52842] ^ n[52843];
assign t[52844] = t[52843] ^ n[52844];
assign t[52845] = t[52844] ^ n[52845];
assign t[52846] = t[52845] ^ n[52846];
assign t[52847] = t[52846] ^ n[52847];
assign t[52848] = t[52847] ^ n[52848];
assign t[52849] = t[52848] ^ n[52849];
assign t[52850] = t[52849] ^ n[52850];
assign t[52851] = t[52850] ^ n[52851];
assign t[52852] = t[52851] ^ n[52852];
assign t[52853] = t[52852] ^ n[52853];
assign t[52854] = t[52853] ^ n[52854];
assign t[52855] = t[52854] ^ n[52855];
assign t[52856] = t[52855] ^ n[52856];
assign t[52857] = t[52856] ^ n[52857];
assign t[52858] = t[52857] ^ n[52858];
assign t[52859] = t[52858] ^ n[52859];
assign t[52860] = t[52859] ^ n[52860];
assign t[52861] = t[52860] ^ n[52861];
assign t[52862] = t[52861] ^ n[52862];
assign t[52863] = t[52862] ^ n[52863];
assign t[52864] = t[52863] ^ n[52864];
assign t[52865] = t[52864] ^ n[52865];
assign t[52866] = t[52865] ^ n[52866];
assign t[52867] = t[52866] ^ n[52867];
assign t[52868] = t[52867] ^ n[52868];
assign t[52869] = t[52868] ^ n[52869];
assign t[52870] = t[52869] ^ n[52870];
assign t[52871] = t[52870] ^ n[52871];
assign t[52872] = t[52871] ^ n[52872];
assign t[52873] = t[52872] ^ n[52873];
assign t[52874] = t[52873] ^ n[52874];
assign t[52875] = t[52874] ^ n[52875];
assign t[52876] = t[52875] ^ n[52876];
assign t[52877] = t[52876] ^ n[52877];
assign t[52878] = t[52877] ^ n[52878];
assign t[52879] = t[52878] ^ n[52879];
assign t[52880] = t[52879] ^ n[52880];
assign t[52881] = t[52880] ^ n[52881];
assign t[52882] = t[52881] ^ n[52882];
assign t[52883] = t[52882] ^ n[52883];
assign t[52884] = t[52883] ^ n[52884];
assign t[52885] = t[52884] ^ n[52885];
assign t[52886] = t[52885] ^ n[52886];
assign t[52887] = t[52886] ^ n[52887];
assign t[52888] = t[52887] ^ n[52888];
assign t[52889] = t[52888] ^ n[52889];
assign t[52890] = t[52889] ^ n[52890];
assign t[52891] = t[52890] ^ n[52891];
assign t[52892] = t[52891] ^ n[52892];
assign t[52893] = t[52892] ^ n[52893];
assign t[52894] = t[52893] ^ n[52894];
assign t[52895] = t[52894] ^ n[52895];
assign t[52896] = t[52895] ^ n[52896];
assign t[52897] = t[52896] ^ n[52897];
assign t[52898] = t[52897] ^ n[52898];
assign t[52899] = t[52898] ^ n[52899];
assign t[52900] = t[52899] ^ n[52900];
assign t[52901] = t[52900] ^ n[52901];
assign t[52902] = t[52901] ^ n[52902];
assign t[52903] = t[52902] ^ n[52903];
assign t[52904] = t[52903] ^ n[52904];
assign t[52905] = t[52904] ^ n[52905];
assign t[52906] = t[52905] ^ n[52906];
assign t[52907] = t[52906] ^ n[52907];
assign t[52908] = t[52907] ^ n[52908];
assign t[52909] = t[52908] ^ n[52909];
assign t[52910] = t[52909] ^ n[52910];
assign t[52911] = t[52910] ^ n[52911];
assign t[52912] = t[52911] ^ n[52912];
assign t[52913] = t[52912] ^ n[52913];
assign t[52914] = t[52913] ^ n[52914];
assign t[52915] = t[52914] ^ n[52915];
assign t[52916] = t[52915] ^ n[52916];
assign t[52917] = t[52916] ^ n[52917];
assign t[52918] = t[52917] ^ n[52918];
assign t[52919] = t[52918] ^ n[52919];
assign t[52920] = t[52919] ^ n[52920];
assign t[52921] = t[52920] ^ n[52921];
assign t[52922] = t[52921] ^ n[52922];
assign t[52923] = t[52922] ^ n[52923];
assign t[52924] = t[52923] ^ n[52924];
assign t[52925] = t[52924] ^ n[52925];
assign t[52926] = t[52925] ^ n[52926];
assign t[52927] = t[52926] ^ n[52927];
assign t[52928] = t[52927] ^ n[52928];
assign t[52929] = t[52928] ^ n[52929];
assign t[52930] = t[52929] ^ n[52930];
assign t[52931] = t[52930] ^ n[52931];
assign t[52932] = t[52931] ^ n[52932];
assign t[52933] = t[52932] ^ n[52933];
assign t[52934] = t[52933] ^ n[52934];
assign t[52935] = t[52934] ^ n[52935];
assign t[52936] = t[52935] ^ n[52936];
assign t[52937] = t[52936] ^ n[52937];
assign t[52938] = t[52937] ^ n[52938];
assign t[52939] = t[52938] ^ n[52939];
assign t[52940] = t[52939] ^ n[52940];
assign t[52941] = t[52940] ^ n[52941];
assign t[52942] = t[52941] ^ n[52942];
assign t[52943] = t[52942] ^ n[52943];
assign t[52944] = t[52943] ^ n[52944];
assign t[52945] = t[52944] ^ n[52945];
assign t[52946] = t[52945] ^ n[52946];
assign t[52947] = t[52946] ^ n[52947];
assign t[52948] = t[52947] ^ n[52948];
assign t[52949] = t[52948] ^ n[52949];
assign t[52950] = t[52949] ^ n[52950];
assign t[52951] = t[52950] ^ n[52951];
assign t[52952] = t[52951] ^ n[52952];
assign t[52953] = t[52952] ^ n[52953];
assign t[52954] = t[52953] ^ n[52954];
assign t[52955] = t[52954] ^ n[52955];
assign t[52956] = t[52955] ^ n[52956];
assign t[52957] = t[52956] ^ n[52957];
assign t[52958] = t[52957] ^ n[52958];
assign t[52959] = t[52958] ^ n[52959];
assign t[52960] = t[52959] ^ n[52960];
assign t[52961] = t[52960] ^ n[52961];
assign t[52962] = t[52961] ^ n[52962];
assign t[52963] = t[52962] ^ n[52963];
assign t[52964] = t[52963] ^ n[52964];
assign t[52965] = t[52964] ^ n[52965];
assign t[52966] = t[52965] ^ n[52966];
assign t[52967] = t[52966] ^ n[52967];
assign t[52968] = t[52967] ^ n[52968];
assign t[52969] = t[52968] ^ n[52969];
assign t[52970] = t[52969] ^ n[52970];
assign t[52971] = t[52970] ^ n[52971];
assign t[52972] = t[52971] ^ n[52972];
assign t[52973] = t[52972] ^ n[52973];
assign t[52974] = t[52973] ^ n[52974];
assign t[52975] = t[52974] ^ n[52975];
assign t[52976] = t[52975] ^ n[52976];
assign t[52977] = t[52976] ^ n[52977];
assign t[52978] = t[52977] ^ n[52978];
assign t[52979] = t[52978] ^ n[52979];
assign t[52980] = t[52979] ^ n[52980];
assign t[52981] = t[52980] ^ n[52981];
assign t[52982] = t[52981] ^ n[52982];
assign t[52983] = t[52982] ^ n[52983];
assign t[52984] = t[52983] ^ n[52984];
assign t[52985] = t[52984] ^ n[52985];
assign t[52986] = t[52985] ^ n[52986];
assign t[52987] = t[52986] ^ n[52987];
assign t[52988] = t[52987] ^ n[52988];
assign t[52989] = t[52988] ^ n[52989];
assign t[52990] = t[52989] ^ n[52990];
assign t[52991] = t[52990] ^ n[52991];
assign t[52992] = t[52991] ^ n[52992];
assign t[52993] = t[52992] ^ n[52993];
assign t[52994] = t[52993] ^ n[52994];
assign t[52995] = t[52994] ^ n[52995];
assign t[52996] = t[52995] ^ n[52996];
assign t[52997] = t[52996] ^ n[52997];
assign t[52998] = t[52997] ^ n[52998];
assign t[52999] = t[52998] ^ n[52999];
assign t[53000] = t[52999] ^ n[53000];
assign t[53001] = t[53000] ^ n[53001];
assign t[53002] = t[53001] ^ n[53002];
assign t[53003] = t[53002] ^ n[53003];
assign t[53004] = t[53003] ^ n[53004];
assign t[53005] = t[53004] ^ n[53005];
assign t[53006] = t[53005] ^ n[53006];
assign t[53007] = t[53006] ^ n[53007];
assign t[53008] = t[53007] ^ n[53008];
assign t[53009] = t[53008] ^ n[53009];
assign t[53010] = t[53009] ^ n[53010];
assign t[53011] = t[53010] ^ n[53011];
assign t[53012] = t[53011] ^ n[53012];
assign t[53013] = t[53012] ^ n[53013];
assign t[53014] = t[53013] ^ n[53014];
assign t[53015] = t[53014] ^ n[53015];
assign t[53016] = t[53015] ^ n[53016];
assign t[53017] = t[53016] ^ n[53017];
assign t[53018] = t[53017] ^ n[53018];
assign t[53019] = t[53018] ^ n[53019];
assign t[53020] = t[53019] ^ n[53020];
assign t[53021] = t[53020] ^ n[53021];
assign t[53022] = t[53021] ^ n[53022];
assign t[53023] = t[53022] ^ n[53023];
assign t[53024] = t[53023] ^ n[53024];
assign t[53025] = t[53024] ^ n[53025];
assign t[53026] = t[53025] ^ n[53026];
assign t[53027] = t[53026] ^ n[53027];
assign t[53028] = t[53027] ^ n[53028];
assign t[53029] = t[53028] ^ n[53029];
assign t[53030] = t[53029] ^ n[53030];
assign t[53031] = t[53030] ^ n[53031];
assign t[53032] = t[53031] ^ n[53032];
assign t[53033] = t[53032] ^ n[53033];
assign t[53034] = t[53033] ^ n[53034];
assign t[53035] = t[53034] ^ n[53035];
assign t[53036] = t[53035] ^ n[53036];
assign t[53037] = t[53036] ^ n[53037];
assign t[53038] = t[53037] ^ n[53038];
assign t[53039] = t[53038] ^ n[53039];
assign t[53040] = t[53039] ^ n[53040];
assign t[53041] = t[53040] ^ n[53041];
assign t[53042] = t[53041] ^ n[53042];
assign t[53043] = t[53042] ^ n[53043];
assign t[53044] = t[53043] ^ n[53044];
assign t[53045] = t[53044] ^ n[53045];
assign t[53046] = t[53045] ^ n[53046];
assign t[53047] = t[53046] ^ n[53047];
assign t[53048] = t[53047] ^ n[53048];
assign t[53049] = t[53048] ^ n[53049];
assign t[53050] = t[53049] ^ n[53050];
assign t[53051] = t[53050] ^ n[53051];
assign t[53052] = t[53051] ^ n[53052];
assign t[53053] = t[53052] ^ n[53053];
assign t[53054] = t[53053] ^ n[53054];
assign t[53055] = t[53054] ^ n[53055];
assign t[53056] = t[53055] ^ n[53056];
assign t[53057] = t[53056] ^ n[53057];
assign t[53058] = t[53057] ^ n[53058];
assign t[53059] = t[53058] ^ n[53059];
assign t[53060] = t[53059] ^ n[53060];
assign t[53061] = t[53060] ^ n[53061];
assign t[53062] = t[53061] ^ n[53062];
assign t[53063] = t[53062] ^ n[53063];
assign t[53064] = t[53063] ^ n[53064];
assign t[53065] = t[53064] ^ n[53065];
assign t[53066] = t[53065] ^ n[53066];
assign t[53067] = t[53066] ^ n[53067];
assign t[53068] = t[53067] ^ n[53068];
assign t[53069] = t[53068] ^ n[53069];
assign t[53070] = t[53069] ^ n[53070];
assign t[53071] = t[53070] ^ n[53071];
assign t[53072] = t[53071] ^ n[53072];
assign t[53073] = t[53072] ^ n[53073];
assign t[53074] = t[53073] ^ n[53074];
assign t[53075] = t[53074] ^ n[53075];
assign t[53076] = t[53075] ^ n[53076];
assign t[53077] = t[53076] ^ n[53077];
assign t[53078] = t[53077] ^ n[53078];
assign t[53079] = t[53078] ^ n[53079];
assign t[53080] = t[53079] ^ n[53080];
assign t[53081] = t[53080] ^ n[53081];
assign t[53082] = t[53081] ^ n[53082];
assign t[53083] = t[53082] ^ n[53083];
assign t[53084] = t[53083] ^ n[53084];
assign t[53085] = t[53084] ^ n[53085];
assign t[53086] = t[53085] ^ n[53086];
assign t[53087] = t[53086] ^ n[53087];
assign t[53088] = t[53087] ^ n[53088];
assign t[53089] = t[53088] ^ n[53089];
assign t[53090] = t[53089] ^ n[53090];
assign t[53091] = t[53090] ^ n[53091];
assign t[53092] = t[53091] ^ n[53092];
assign t[53093] = t[53092] ^ n[53093];
assign t[53094] = t[53093] ^ n[53094];
assign t[53095] = t[53094] ^ n[53095];
assign t[53096] = t[53095] ^ n[53096];
assign t[53097] = t[53096] ^ n[53097];
assign t[53098] = t[53097] ^ n[53098];
assign t[53099] = t[53098] ^ n[53099];
assign t[53100] = t[53099] ^ n[53100];
assign t[53101] = t[53100] ^ n[53101];
assign t[53102] = t[53101] ^ n[53102];
assign t[53103] = t[53102] ^ n[53103];
assign t[53104] = t[53103] ^ n[53104];
assign t[53105] = t[53104] ^ n[53105];
assign t[53106] = t[53105] ^ n[53106];
assign t[53107] = t[53106] ^ n[53107];
assign t[53108] = t[53107] ^ n[53108];
assign t[53109] = t[53108] ^ n[53109];
assign t[53110] = t[53109] ^ n[53110];
assign t[53111] = t[53110] ^ n[53111];
assign t[53112] = t[53111] ^ n[53112];
assign t[53113] = t[53112] ^ n[53113];
assign t[53114] = t[53113] ^ n[53114];
assign t[53115] = t[53114] ^ n[53115];
assign t[53116] = t[53115] ^ n[53116];
assign t[53117] = t[53116] ^ n[53117];
assign t[53118] = t[53117] ^ n[53118];
assign t[53119] = t[53118] ^ n[53119];
assign t[53120] = t[53119] ^ n[53120];
assign t[53121] = t[53120] ^ n[53121];
assign t[53122] = t[53121] ^ n[53122];
assign t[53123] = t[53122] ^ n[53123];
assign t[53124] = t[53123] ^ n[53124];
assign t[53125] = t[53124] ^ n[53125];
assign t[53126] = t[53125] ^ n[53126];
assign t[53127] = t[53126] ^ n[53127];
assign t[53128] = t[53127] ^ n[53128];
assign t[53129] = t[53128] ^ n[53129];
assign t[53130] = t[53129] ^ n[53130];
assign t[53131] = t[53130] ^ n[53131];
assign t[53132] = t[53131] ^ n[53132];
assign t[53133] = t[53132] ^ n[53133];
assign t[53134] = t[53133] ^ n[53134];
assign t[53135] = t[53134] ^ n[53135];
assign t[53136] = t[53135] ^ n[53136];
assign t[53137] = t[53136] ^ n[53137];
assign t[53138] = t[53137] ^ n[53138];
assign t[53139] = t[53138] ^ n[53139];
assign t[53140] = t[53139] ^ n[53140];
assign t[53141] = t[53140] ^ n[53141];
assign t[53142] = t[53141] ^ n[53142];
assign t[53143] = t[53142] ^ n[53143];
assign t[53144] = t[53143] ^ n[53144];
assign t[53145] = t[53144] ^ n[53145];
assign t[53146] = t[53145] ^ n[53146];
assign t[53147] = t[53146] ^ n[53147];
assign t[53148] = t[53147] ^ n[53148];
assign t[53149] = t[53148] ^ n[53149];
assign t[53150] = t[53149] ^ n[53150];
assign t[53151] = t[53150] ^ n[53151];
assign t[53152] = t[53151] ^ n[53152];
assign t[53153] = t[53152] ^ n[53153];
assign t[53154] = t[53153] ^ n[53154];
assign t[53155] = t[53154] ^ n[53155];
assign t[53156] = t[53155] ^ n[53156];
assign t[53157] = t[53156] ^ n[53157];
assign t[53158] = t[53157] ^ n[53158];
assign t[53159] = t[53158] ^ n[53159];
assign t[53160] = t[53159] ^ n[53160];
assign t[53161] = t[53160] ^ n[53161];
assign t[53162] = t[53161] ^ n[53162];
assign t[53163] = t[53162] ^ n[53163];
assign t[53164] = t[53163] ^ n[53164];
assign t[53165] = t[53164] ^ n[53165];
assign t[53166] = t[53165] ^ n[53166];
assign t[53167] = t[53166] ^ n[53167];
assign t[53168] = t[53167] ^ n[53168];
assign t[53169] = t[53168] ^ n[53169];
assign t[53170] = t[53169] ^ n[53170];
assign t[53171] = t[53170] ^ n[53171];
assign t[53172] = t[53171] ^ n[53172];
assign t[53173] = t[53172] ^ n[53173];
assign t[53174] = t[53173] ^ n[53174];
assign t[53175] = t[53174] ^ n[53175];
assign t[53176] = t[53175] ^ n[53176];
assign t[53177] = t[53176] ^ n[53177];
assign t[53178] = t[53177] ^ n[53178];
assign t[53179] = t[53178] ^ n[53179];
assign t[53180] = t[53179] ^ n[53180];
assign t[53181] = t[53180] ^ n[53181];
assign t[53182] = t[53181] ^ n[53182];
assign t[53183] = t[53182] ^ n[53183];
assign t[53184] = t[53183] ^ n[53184];
assign t[53185] = t[53184] ^ n[53185];
assign t[53186] = t[53185] ^ n[53186];
assign t[53187] = t[53186] ^ n[53187];
assign t[53188] = t[53187] ^ n[53188];
assign t[53189] = t[53188] ^ n[53189];
assign t[53190] = t[53189] ^ n[53190];
assign t[53191] = t[53190] ^ n[53191];
assign t[53192] = t[53191] ^ n[53192];
assign t[53193] = t[53192] ^ n[53193];
assign t[53194] = t[53193] ^ n[53194];
assign t[53195] = t[53194] ^ n[53195];
assign t[53196] = t[53195] ^ n[53196];
assign t[53197] = t[53196] ^ n[53197];
assign t[53198] = t[53197] ^ n[53198];
assign t[53199] = t[53198] ^ n[53199];
assign t[53200] = t[53199] ^ n[53200];
assign t[53201] = t[53200] ^ n[53201];
assign t[53202] = t[53201] ^ n[53202];
assign t[53203] = t[53202] ^ n[53203];
assign t[53204] = t[53203] ^ n[53204];
assign t[53205] = t[53204] ^ n[53205];
assign t[53206] = t[53205] ^ n[53206];
assign t[53207] = t[53206] ^ n[53207];
assign t[53208] = t[53207] ^ n[53208];
assign t[53209] = t[53208] ^ n[53209];
assign t[53210] = t[53209] ^ n[53210];
assign t[53211] = t[53210] ^ n[53211];
assign t[53212] = t[53211] ^ n[53212];
assign t[53213] = t[53212] ^ n[53213];
assign t[53214] = t[53213] ^ n[53214];
assign t[53215] = t[53214] ^ n[53215];
assign t[53216] = t[53215] ^ n[53216];
assign t[53217] = t[53216] ^ n[53217];
assign t[53218] = t[53217] ^ n[53218];
assign t[53219] = t[53218] ^ n[53219];
assign t[53220] = t[53219] ^ n[53220];
assign t[53221] = t[53220] ^ n[53221];
assign t[53222] = t[53221] ^ n[53222];
assign t[53223] = t[53222] ^ n[53223];
assign t[53224] = t[53223] ^ n[53224];
assign t[53225] = t[53224] ^ n[53225];
assign t[53226] = t[53225] ^ n[53226];
assign t[53227] = t[53226] ^ n[53227];
assign t[53228] = t[53227] ^ n[53228];
assign t[53229] = t[53228] ^ n[53229];
assign t[53230] = t[53229] ^ n[53230];
assign t[53231] = t[53230] ^ n[53231];
assign t[53232] = t[53231] ^ n[53232];
assign t[53233] = t[53232] ^ n[53233];
assign t[53234] = t[53233] ^ n[53234];
assign t[53235] = t[53234] ^ n[53235];
assign t[53236] = t[53235] ^ n[53236];
assign t[53237] = t[53236] ^ n[53237];
assign t[53238] = t[53237] ^ n[53238];
assign t[53239] = t[53238] ^ n[53239];
assign t[53240] = t[53239] ^ n[53240];
assign t[53241] = t[53240] ^ n[53241];
assign t[53242] = t[53241] ^ n[53242];
assign t[53243] = t[53242] ^ n[53243];
assign t[53244] = t[53243] ^ n[53244];
assign t[53245] = t[53244] ^ n[53245];
assign t[53246] = t[53245] ^ n[53246];
assign t[53247] = t[53246] ^ n[53247];
assign t[53248] = t[53247] ^ n[53248];
assign t[53249] = t[53248] ^ n[53249];
assign t[53250] = t[53249] ^ n[53250];
assign t[53251] = t[53250] ^ n[53251];
assign t[53252] = t[53251] ^ n[53252];
assign t[53253] = t[53252] ^ n[53253];
assign t[53254] = t[53253] ^ n[53254];
assign t[53255] = t[53254] ^ n[53255];
assign t[53256] = t[53255] ^ n[53256];
assign t[53257] = t[53256] ^ n[53257];
assign t[53258] = t[53257] ^ n[53258];
assign t[53259] = t[53258] ^ n[53259];
assign t[53260] = t[53259] ^ n[53260];
assign t[53261] = t[53260] ^ n[53261];
assign t[53262] = t[53261] ^ n[53262];
assign t[53263] = t[53262] ^ n[53263];
assign t[53264] = t[53263] ^ n[53264];
assign t[53265] = t[53264] ^ n[53265];
assign t[53266] = t[53265] ^ n[53266];
assign t[53267] = t[53266] ^ n[53267];
assign t[53268] = t[53267] ^ n[53268];
assign t[53269] = t[53268] ^ n[53269];
assign t[53270] = t[53269] ^ n[53270];
assign t[53271] = t[53270] ^ n[53271];
assign t[53272] = t[53271] ^ n[53272];
assign t[53273] = t[53272] ^ n[53273];
assign t[53274] = t[53273] ^ n[53274];
assign t[53275] = t[53274] ^ n[53275];
assign t[53276] = t[53275] ^ n[53276];
assign t[53277] = t[53276] ^ n[53277];
assign t[53278] = t[53277] ^ n[53278];
assign t[53279] = t[53278] ^ n[53279];
assign t[53280] = t[53279] ^ n[53280];
assign t[53281] = t[53280] ^ n[53281];
assign t[53282] = t[53281] ^ n[53282];
assign t[53283] = t[53282] ^ n[53283];
assign t[53284] = t[53283] ^ n[53284];
assign t[53285] = t[53284] ^ n[53285];
assign t[53286] = t[53285] ^ n[53286];
assign t[53287] = t[53286] ^ n[53287];
assign t[53288] = t[53287] ^ n[53288];
assign t[53289] = t[53288] ^ n[53289];
assign t[53290] = t[53289] ^ n[53290];
assign t[53291] = t[53290] ^ n[53291];
assign t[53292] = t[53291] ^ n[53292];
assign t[53293] = t[53292] ^ n[53293];
assign t[53294] = t[53293] ^ n[53294];
assign t[53295] = t[53294] ^ n[53295];
assign t[53296] = t[53295] ^ n[53296];
assign t[53297] = t[53296] ^ n[53297];
assign t[53298] = t[53297] ^ n[53298];
assign t[53299] = t[53298] ^ n[53299];
assign t[53300] = t[53299] ^ n[53300];
assign t[53301] = t[53300] ^ n[53301];
assign t[53302] = t[53301] ^ n[53302];
assign t[53303] = t[53302] ^ n[53303];
assign t[53304] = t[53303] ^ n[53304];
assign t[53305] = t[53304] ^ n[53305];
assign t[53306] = t[53305] ^ n[53306];
assign t[53307] = t[53306] ^ n[53307];
assign t[53308] = t[53307] ^ n[53308];
assign t[53309] = t[53308] ^ n[53309];
assign t[53310] = t[53309] ^ n[53310];
assign t[53311] = t[53310] ^ n[53311];
assign t[53312] = t[53311] ^ n[53312];
assign t[53313] = t[53312] ^ n[53313];
assign t[53314] = t[53313] ^ n[53314];
assign t[53315] = t[53314] ^ n[53315];
assign t[53316] = t[53315] ^ n[53316];
assign t[53317] = t[53316] ^ n[53317];
assign t[53318] = t[53317] ^ n[53318];
assign t[53319] = t[53318] ^ n[53319];
assign t[53320] = t[53319] ^ n[53320];
assign t[53321] = t[53320] ^ n[53321];
assign t[53322] = t[53321] ^ n[53322];
assign t[53323] = t[53322] ^ n[53323];
assign t[53324] = t[53323] ^ n[53324];
assign t[53325] = t[53324] ^ n[53325];
assign t[53326] = t[53325] ^ n[53326];
assign t[53327] = t[53326] ^ n[53327];
assign t[53328] = t[53327] ^ n[53328];
assign t[53329] = t[53328] ^ n[53329];
assign t[53330] = t[53329] ^ n[53330];
assign t[53331] = t[53330] ^ n[53331];
assign t[53332] = t[53331] ^ n[53332];
assign t[53333] = t[53332] ^ n[53333];
assign t[53334] = t[53333] ^ n[53334];
assign t[53335] = t[53334] ^ n[53335];
assign t[53336] = t[53335] ^ n[53336];
assign t[53337] = t[53336] ^ n[53337];
assign t[53338] = t[53337] ^ n[53338];
assign t[53339] = t[53338] ^ n[53339];
assign t[53340] = t[53339] ^ n[53340];
assign t[53341] = t[53340] ^ n[53341];
assign t[53342] = t[53341] ^ n[53342];
assign t[53343] = t[53342] ^ n[53343];
assign t[53344] = t[53343] ^ n[53344];
assign t[53345] = t[53344] ^ n[53345];
assign t[53346] = t[53345] ^ n[53346];
assign t[53347] = t[53346] ^ n[53347];
assign t[53348] = t[53347] ^ n[53348];
assign t[53349] = t[53348] ^ n[53349];
assign t[53350] = t[53349] ^ n[53350];
assign t[53351] = t[53350] ^ n[53351];
assign t[53352] = t[53351] ^ n[53352];
assign t[53353] = t[53352] ^ n[53353];
assign t[53354] = t[53353] ^ n[53354];
assign t[53355] = t[53354] ^ n[53355];
assign t[53356] = t[53355] ^ n[53356];
assign t[53357] = t[53356] ^ n[53357];
assign t[53358] = t[53357] ^ n[53358];
assign t[53359] = t[53358] ^ n[53359];
assign t[53360] = t[53359] ^ n[53360];
assign t[53361] = t[53360] ^ n[53361];
assign t[53362] = t[53361] ^ n[53362];
assign t[53363] = t[53362] ^ n[53363];
assign t[53364] = t[53363] ^ n[53364];
assign t[53365] = t[53364] ^ n[53365];
assign t[53366] = t[53365] ^ n[53366];
assign t[53367] = t[53366] ^ n[53367];
assign t[53368] = t[53367] ^ n[53368];
assign t[53369] = t[53368] ^ n[53369];
assign t[53370] = t[53369] ^ n[53370];
assign t[53371] = t[53370] ^ n[53371];
assign t[53372] = t[53371] ^ n[53372];
assign t[53373] = t[53372] ^ n[53373];
assign t[53374] = t[53373] ^ n[53374];
assign t[53375] = t[53374] ^ n[53375];
assign t[53376] = t[53375] ^ n[53376];
assign t[53377] = t[53376] ^ n[53377];
assign t[53378] = t[53377] ^ n[53378];
assign t[53379] = t[53378] ^ n[53379];
assign t[53380] = t[53379] ^ n[53380];
assign t[53381] = t[53380] ^ n[53381];
assign t[53382] = t[53381] ^ n[53382];
assign t[53383] = t[53382] ^ n[53383];
assign t[53384] = t[53383] ^ n[53384];
assign t[53385] = t[53384] ^ n[53385];
assign t[53386] = t[53385] ^ n[53386];
assign t[53387] = t[53386] ^ n[53387];
assign t[53388] = t[53387] ^ n[53388];
assign t[53389] = t[53388] ^ n[53389];
assign t[53390] = t[53389] ^ n[53390];
assign t[53391] = t[53390] ^ n[53391];
assign t[53392] = t[53391] ^ n[53392];
assign t[53393] = t[53392] ^ n[53393];
assign t[53394] = t[53393] ^ n[53394];
assign t[53395] = t[53394] ^ n[53395];
assign t[53396] = t[53395] ^ n[53396];
assign t[53397] = t[53396] ^ n[53397];
assign t[53398] = t[53397] ^ n[53398];
assign t[53399] = t[53398] ^ n[53399];
assign t[53400] = t[53399] ^ n[53400];
assign t[53401] = t[53400] ^ n[53401];
assign t[53402] = t[53401] ^ n[53402];
assign t[53403] = t[53402] ^ n[53403];
assign t[53404] = t[53403] ^ n[53404];
assign t[53405] = t[53404] ^ n[53405];
assign t[53406] = t[53405] ^ n[53406];
assign t[53407] = t[53406] ^ n[53407];
assign t[53408] = t[53407] ^ n[53408];
assign t[53409] = t[53408] ^ n[53409];
assign t[53410] = t[53409] ^ n[53410];
assign t[53411] = t[53410] ^ n[53411];
assign t[53412] = t[53411] ^ n[53412];
assign t[53413] = t[53412] ^ n[53413];
assign t[53414] = t[53413] ^ n[53414];
assign t[53415] = t[53414] ^ n[53415];
assign t[53416] = t[53415] ^ n[53416];
assign t[53417] = t[53416] ^ n[53417];
assign t[53418] = t[53417] ^ n[53418];
assign t[53419] = t[53418] ^ n[53419];
assign t[53420] = t[53419] ^ n[53420];
assign t[53421] = t[53420] ^ n[53421];
assign t[53422] = t[53421] ^ n[53422];
assign t[53423] = t[53422] ^ n[53423];
assign t[53424] = t[53423] ^ n[53424];
assign t[53425] = t[53424] ^ n[53425];
assign t[53426] = t[53425] ^ n[53426];
assign t[53427] = t[53426] ^ n[53427];
assign t[53428] = t[53427] ^ n[53428];
assign t[53429] = t[53428] ^ n[53429];
assign t[53430] = t[53429] ^ n[53430];
assign t[53431] = t[53430] ^ n[53431];
assign t[53432] = t[53431] ^ n[53432];
assign t[53433] = t[53432] ^ n[53433];
assign t[53434] = t[53433] ^ n[53434];
assign t[53435] = t[53434] ^ n[53435];
assign t[53436] = t[53435] ^ n[53436];
assign t[53437] = t[53436] ^ n[53437];
assign t[53438] = t[53437] ^ n[53438];
assign t[53439] = t[53438] ^ n[53439];
assign t[53440] = t[53439] ^ n[53440];
assign t[53441] = t[53440] ^ n[53441];
assign t[53442] = t[53441] ^ n[53442];
assign t[53443] = t[53442] ^ n[53443];
assign t[53444] = t[53443] ^ n[53444];
assign t[53445] = t[53444] ^ n[53445];
assign t[53446] = t[53445] ^ n[53446];
assign t[53447] = t[53446] ^ n[53447];
assign t[53448] = t[53447] ^ n[53448];
assign t[53449] = t[53448] ^ n[53449];
assign t[53450] = t[53449] ^ n[53450];
assign t[53451] = t[53450] ^ n[53451];
assign t[53452] = t[53451] ^ n[53452];
assign t[53453] = t[53452] ^ n[53453];
assign t[53454] = t[53453] ^ n[53454];
assign t[53455] = t[53454] ^ n[53455];
assign t[53456] = t[53455] ^ n[53456];
assign t[53457] = t[53456] ^ n[53457];
assign t[53458] = t[53457] ^ n[53458];
assign t[53459] = t[53458] ^ n[53459];
assign t[53460] = t[53459] ^ n[53460];
assign t[53461] = t[53460] ^ n[53461];
assign t[53462] = t[53461] ^ n[53462];
assign t[53463] = t[53462] ^ n[53463];
assign t[53464] = t[53463] ^ n[53464];
assign t[53465] = t[53464] ^ n[53465];
assign t[53466] = t[53465] ^ n[53466];
assign t[53467] = t[53466] ^ n[53467];
assign t[53468] = t[53467] ^ n[53468];
assign t[53469] = t[53468] ^ n[53469];
assign t[53470] = t[53469] ^ n[53470];
assign t[53471] = t[53470] ^ n[53471];
assign t[53472] = t[53471] ^ n[53472];
assign t[53473] = t[53472] ^ n[53473];
assign t[53474] = t[53473] ^ n[53474];
assign t[53475] = t[53474] ^ n[53475];
assign t[53476] = t[53475] ^ n[53476];
assign t[53477] = t[53476] ^ n[53477];
assign t[53478] = t[53477] ^ n[53478];
assign t[53479] = t[53478] ^ n[53479];
assign t[53480] = t[53479] ^ n[53480];
assign t[53481] = t[53480] ^ n[53481];
assign t[53482] = t[53481] ^ n[53482];
assign t[53483] = t[53482] ^ n[53483];
assign t[53484] = t[53483] ^ n[53484];
assign t[53485] = t[53484] ^ n[53485];
assign t[53486] = t[53485] ^ n[53486];
assign t[53487] = t[53486] ^ n[53487];
assign t[53488] = t[53487] ^ n[53488];
assign t[53489] = t[53488] ^ n[53489];
assign t[53490] = t[53489] ^ n[53490];
assign t[53491] = t[53490] ^ n[53491];
assign t[53492] = t[53491] ^ n[53492];
assign t[53493] = t[53492] ^ n[53493];
assign t[53494] = t[53493] ^ n[53494];
assign t[53495] = t[53494] ^ n[53495];
assign t[53496] = t[53495] ^ n[53496];
assign t[53497] = t[53496] ^ n[53497];
assign t[53498] = t[53497] ^ n[53498];
assign t[53499] = t[53498] ^ n[53499];
assign t[53500] = t[53499] ^ n[53500];
assign t[53501] = t[53500] ^ n[53501];
assign t[53502] = t[53501] ^ n[53502];
assign t[53503] = t[53502] ^ n[53503];
assign t[53504] = t[53503] ^ n[53504];
assign t[53505] = t[53504] ^ n[53505];
assign t[53506] = t[53505] ^ n[53506];
assign t[53507] = t[53506] ^ n[53507];
assign t[53508] = t[53507] ^ n[53508];
assign t[53509] = t[53508] ^ n[53509];
assign t[53510] = t[53509] ^ n[53510];
assign t[53511] = t[53510] ^ n[53511];
assign t[53512] = t[53511] ^ n[53512];
assign t[53513] = t[53512] ^ n[53513];
assign t[53514] = t[53513] ^ n[53514];
assign t[53515] = t[53514] ^ n[53515];
assign t[53516] = t[53515] ^ n[53516];
assign t[53517] = t[53516] ^ n[53517];
assign t[53518] = t[53517] ^ n[53518];
assign t[53519] = t[53518] ^ n[53519];
assign t[53520] = t[53519] ^ n[53520];
assign t[53521] = t[53520] ^ n[53521];
assign t[53522] = t[53521] ^ n[53522];
assign t[53523] = t[53522] ^ n[53523];
assign t[53524] = t[53523] ^ n[53524];
assign t[53525] = t[53524] ^ n[53525];
assign t[53526] = t[53525] ^ n[53526];
assign t[53527] = t[53526] ^ n[53527];
assign t[53528] = t[53527] ^ n[53528];
assign t[53529] = t[53528] ^ n[53529];
assign t[53530] = t[53529] ^ n[53530];
assign t[53531] = t[53530] ^ n[53531];
assign t[53532] = t[53531] ^ n[53532];
assign t[53533] = t[53532] ^ n[53533];
assign t[53534] = t[53533] ^ n[53534];
assign t[53535] = t[53534] ^ n[53535];
assign t[53536] = t[53535] ^ n[53536];
assign t[53537] = t[53536] ^ n[53537];
assign t[53538] = t[53537] ^ n[53538];
assign t[53539] = t[53538] ^ n[53539];
assign t[53540] = t[53539] ^ n[53540];
assign t[53541] = t[53540] ^ n[53541];
assign t[53542] = t[53541] ^ n[53542];
assign t[53543] = t[53542] ^ n[53543];
assign t[53544] = t[53543] ^ n[53544];
assign t[53545] = t[53544] ^ n[53545];
assign t[53546] = t[53545] ^ n[53546];
assign t[53547] = t[53546] ^ n[53547];
assign t[53548] = t[53547] ^ n[53548];
assign t[53549] = t[53548] ^ n[53549];
assign t[53550] = t[53549] ^ n[53550];
assign t[53551] = t[53550] ^ n[53551];
assign t[53552] = t[53551] ^ n[53552];
assign t[53553] = t[53552] ^ n[53553];
assign t[53554] = t[53553] ^ n[53554];
assign t[53555] = t[53554] ^ n[53555];
assign t[53556] = t[53555] ^ n[53556];
assign t[53557] = t[53556] ^ n[53557];
assign t[53558] = t[53557] ^ n[53558];
assign t[53559] = t[53558] ^ n[53559];
assign t[53560] = t[53559] ^ n[53560];
assign t[53561] = t[53560] ^ n[53561];
assign t[53562] = t[53561] ^ n[53562];
assign t[53563] = t[53562] ^ n[53563];
assign t[53564] = t[53563] ^ n[53564];
assign t[53565] = t[53564] ^ n[53565];
assign t[53566] = t[53565] ^ n[53566];
assign t[53567] = t[53566] ^ n[53567];
assign t[53568] = t[53567] ^ n[53568];
assign t[53569] = t[53568] ^ n[53569];
assign t[53570] = t[53569] ^ n[53570];
assign t[53571] = t[53570] ^ n[53571];
assign t[53572] = t[53571] ^ n[53572];
assign t[53573] = t[53572] ^ n[53573];
assign t[53574] = t[53573] ^ n[53574];
assign t[53575] = t[53574] ^ n[53575];
assign t[53576] = t[53575] ^ n[53576];
assign t[53577] = t[53576] ^ n[53577];
assign t[53578] = t[53577] ^ n[53578];
assign t[53579] = t[53578] ^ n[53579];
assign t[53580] = t[53579] ^ n[53580];
assign t[53581] = t[53580] ^ n[53581];
assign t[53582] = t[53581] ^ n[53582];
assign t[53583] = t[53582] ^ n[53583];
assign t[53584] = t[53583] ^ n[53584];
assign t[53585] = t[53584] ^ n[53585];
assign t[53586] = t[53585] ^ n[53586];
assign t[53587] = t[53586] ^ n[53587];
assign t[53588] = t[53587] ^ n[53588];
assign t[53589] = t[53588] ^ n[53589];
assign t[53590] = t[53589] ^ n[53590];
assign t[53591] = t[53590] ^ n[53591];
assign t[53592] = t[53591] ^ n[53592];
assign t[53593] = t[53592] ^ n[53593];
assign t[53594] = t[53593] ^ n[53594];
assign t[53595] = t[53594] ^ n[53595];
assign t[53596] = t[53595] ^ n[53596];
assign t[53597] = t[53596] ^ n[53597];
assign t[53598] = t[53597] ^ n[53598];
assign t[53599] = t[53598] ^ n[53599];
assign t[53600] = t[53599] ^ n[53600];
assign t[53601] = t[53600] ^ n[53601];
assign t[53602] = t[53601] ^ n[53602];
assign t[53603] = t[53602] ^ n[53603];
assign t[53604] = t[53603] ^ n[53604];
assign t[53605] = t[53604] ^ n[53605];
assign t[53606] = t[53605] ^ n[53606];
assign t[53607] = t[53606] ^ n[53607];
assign t[53608] = t[53607] ^ n[53608];
assign t[53609] = t[53608] ^ n[53609];
assign t[53610] = t[53609] ^ n[53610];
assign t[53611] = t[53610] ^ n[53611];
assign t[53612] = t[53611] ^ n[53612];
assign t[53613] = t[53612] ^ n[53613];
assign t[53614] = t[53613] ^ n[53614];
assign t[53615] = t[53614] ^ n[53615];
assign t[53616] = t[53615] ^ n[53616];
assign t[53617] = t[53616] ^ n[53617];
assign t[53618] = t[53617] ^ n[53618];
assign t[53619] = t[53618] ^ n[53619];
assign t[53620] = t[53619] ^ n[53620];
assign t[53621] = t[53620] ^ n[53621];
assign t[53622] = t[53621] ^ n[53622];
assign t[53623] = t[53622] ^ n[53623];
assign t[53624] = t[53623] ^ n[53624];
assign t[53625] = t[53624] ^ n[53625];
assign t[53626] = t[53625] ^ n[53626];
assign t[53627] = t[53626] ^ n[53627];
assign t[53628] = t[53627] ^ n[53628];
assign t[53629] = t[53628] ^ n[53629];
assign t[53630] = t[53629] ^ n[53630];
assign t[53631] = t[53630] ^ n[53631];
assign t[53632] = t[53631] ^ n[53632];
assign t[53633] = t[53632] ^ n[53633];
assign t[53634] = t[53633] ^ n[53634];
assign t[53635] = t[53634] ^ n[53635];
assign t[53636] = t[53635] ^ n[53636];
assign t[53637] = t[53636] ^ n[53637];
assign t[53638] = t[53637] ^ n[53638];
assign t[53639] = t[53638] ^ n[53639];
assign t[53640] = t[53639] ^ n[53640];
assign t[53641] = t[53640] ^ n[53641];
assign t[53642] = t[53641] ^ n[53642];
assign t[53643] = t[53642] ^ n[53643];
assign t[53644] = t[53643] ^ n[53644];
assign t[53645] = t[53644] ^ n[53645];
assign t[53646] = t[53645] ^ n[53646];
assign t[53647] = t[53646] ^ n[53647];
assign t[53648] = t[53647] ^ n[53648];
assign t[53649] = t[53648] ^ n[53649];
assign t[53650] = t[53649] ^ n[53650];
assign t[53651] = t[53650] ^ n[53651];
assign t[53652] = t[53651] ^ n[53652];
assign t[53653] = t[53652] ^ n[53653];
assign t[53654] = t[53653] ^ n[53654];
assign t[53655] = t[53654] ^ n[53655];
assign t[53656] = t[53655] ^ n[53656];
assign t[53657] = t[53656] ^ n[53657];
assign t[53658] = t[53657] ^ n[53658];
assign t[53659] = t[53658] ^ n[53659];
assign t[53660] = t[53659] ^ n[53660];
assign t[53661] = t[53660] ^ n[53661];
assign t[53662] = t[53661] ^ n[53662];
assign t[53663] = t[53662] ^ n[53663];
assign t[53664] = t[53663] ^ n[53664];
assign t[53665] = t[53664] ^ n[53665];
assign t[53666] = t[53665] ^ n[53666];
assign t[53667] = t[53666] ^ n[53667];
assign t[53668] = t[53667] ^ n[53668];
assign t[53669] = t[53668] ^ n[53669];
assign t[53670] = t[53669] ^ n[53670];
assign t[53671] = t[53670] ^ n[53671];
assign t[53672] = t[53671] ^ n[53672];
assign t[53673] = t[53672] ^ n[53673];
assign t[53674] = t[53673] ^ n[53674];
assign t[53675] = t[53674] ^ n[53675];
assign t[53676] = t[53675] ^ n[53676];
assign t[53677] = t[53676] ^ n[53677];
assign t[53678] = t[53677] ^ n[53678];
assign t[53679] = t[53678] ^ n[53679];
assign t[53680] = t[53679] ^ n[53680];
assign t[53681] = t[53680] ^ n[53681];
assign t[53682] = t[53681] ^ n[53682];
assign t[53683] = t[53682] ^ n[53683];
assign t[53684] = t[53683] ^ n[53684];
assign t[53685] = t[53684] ^ n[53685];
assign t[53686] = t[53685] ^ n[53686];
assign t[53687] = t[53686] ^ n[53687];
assign t[53688] = t[53687] ^ n[53688];
assign t[53689] = t[53688] ^ n[53689];
assign t[53690] = t[53689] ^ n[53690];
assign t[53691] = t[53690] ^ n[53691];
assign t[53692] = t[53691] ^ n[53692];
assign t[53693] = t[53692] ^ n[53693];
assign t[53694] = t[53693] ^ n[53694];
assign t[53695] = t[53694] ^ n[53695];
assign t[53696] = t[53695] ^ n[53696];
assign t[53697] = t[53696] ^ n[53697];
assign t[53698] = t[53697] ^ n[53698];
assign t[53699] = t[53698] ^ n[53699];
assign t[53700] = t[53699] ^ n[53700];
assign t[53701] = t[53700] ^ n[53701];
assign t[53702] = t[53701] ^ n[53702];
assign t[53703] = t[53702] ^ n[53703];
assign t[53704] = t[53703] ^ n[53704];
assign t[53705] = t[53704] ^ n[53705];
assign t[53706] = t[53705] ^ n[53706];
assign t[53707] = t[53706] ^ n[53707];
assign t[53708] = t[53707] ^ n[53708];
assign t[53709] = t[53708] ^ n[53709];
assign t[53710] = t[53709] ^ n[53710];
assign t[53711] = t[53710] ^ n[53711];
assign t[53712] = t[53711] ^ n[53712];
assign t[53713] = t[53712] ^ n[53713];
assign t[53714] = t[53713] ^ n[53714];
assign t[53715] = t[53714] ^ n[53715];
assign t[53716] = t[53715] ^ n[53716];
assign t[53717] = t[53716] ^ n[53717];
assign t[53718] = t[53717] ^ n[53718];
assign t[53719] = t[53718] ^ n[53719];
assign t[53720] = t[53719] ^ n[53720];
assign t[53721] = t[53720] ^ n[53721];
assign t[53722] = t[53721] ^ n[53722];
assign t[53723] = t[53722] ^ n[53723];
assign t[53724] = t[53723] ^ n[53724];
assign t[53725] = t[53724] ^ n[53725];
assign t[53726] = t[53725] ^ n[53726];
assign t[53727] = t[53726] ^ n[53727];
assign t[53728] = t[53727] ^ n[53728];
assign t[53729] = t[53728] ^ n[53729];
assign t[53730] = t[53729] ^ n[53730];
assign t[53731] = t[53730] ^ n[53731];
assign t[53732] = t[53731] ^ n[53732];
assign t[53733] = t[53732] ^ n[53733];
assign t[53734] = t[53733] ^ n[53734];
assign t[53735] = t[53734] ^ n[53735];
assign t[53736] = t[53735] ^ n[53736];
assign t[53737] = t[53736] ^ n[53737];
assign t[53738] = t[53737] ^ n[53738];
assign t[53739] = t[53738] ^ n[53739];
assign t[53740] = t[53739] ^ n[53740];
assign t[53741] = t[53740] ^ n[53741];
assign t[53742] = t[53741] ^ n[53742];
assign t[53743] = t[53742] ^ n[53743];
assign t[53744] = t[53743] ^ n[53744];
assign t[53745] = t[53744] ^ n[53745];
assign t[53746] = t[53745] ^ n[53746];
assign t[53747] = t[53746] ^ n[53747];
assign t[53748] = t[53747] ^ n[53748];
assign t[53749] = t[53748] ^ n[53749];
assign t[53750] = t[53749] ^ n[53750];
assign t[53751] = t[53750] ^ n[53751];
assign t[53752] = t[53751] ^ n[53752];
assign t[53753] = t[53752] ^ n[53753];
assign t[53754] = t[53753] ^ n[53754];
assign t[53755] = t[53754] ^ n[53755];
assign t[53756] = t[53755] ^ n[53756];
assign t[53757] = t[53756] ^ n[53757];
assign t[53758] = t[53757] ^ n[53758];
assign t[53759] = t[53758] ^ n[53759];
assign t[53760] = t[53759] ^ n[53760];
assign t[53761] = t[53760] ^ n[53761];
assign t[53762] = t[53761] ^ n[53762];
assign t[53763] = t[53762] ^ n[53763];
assign t[53764] = t[53763] ^ n[53764];
assign t[53765] = t[53764] ^ n[53765];
assign t[53766] = t[53765] ^ n[53766];
assign t[53767] = t[53766] ^ n[53767];
assign t[53768] = t[53767] ^ n[53768];
assign t[53769] = t[53768] ^ n[53769];
assign t[53770] = t[53769] ^ n[53770];
assign t[53771] = t[53770] ^ n[53771];
assign t[53772] = t[53771] ^ n[53772];
assign t[53773] = t[53772] ^ n[53773];
assign t[53774] = t[53773] ^ n[53774];
assign t[53775] = t[53774] ^ n[53775];
assign t[53776] = t[53775] ^ n[53776];
assign t[53777] = t[53776] ^ n[53777];
assign t[53778] = t[53777] ^ n[53778];
assign t[53779] = t[53778] ^ n[53779];
assign t[53780] = t[53779] ^ n[53780];
assign t[53781] = t[53780] ^ n[53781];
assign t[53782] = t[53781] ^ n[53782];
assign t[53783] = t[53782] ^ n[53783];
assign t[53784] = t[53783] ^ n[53784];
assign t[53785] = t[53784] ^ n[53785];
assign t[53786] = t[53785] ^ n[53786];
assign t[53787] = t[53786] ^ n[53787];
assign t[53788] = t[53787] ^ n[53788];
assign t[53789] = t[53788] ^ n[53789];
assign t[53790] = t[53789] ^ n[53790];
assign t[53791] = t[53790] ^ n[53791];
assign t[53792] = t[53791] ^ n[53792];
assign t[53793] = t[53792] ^ n[53793];
assign t[53794] = t[53793] ^ n[53794];
assign t[53795] = t[53794] ^ n[53795];
assign t[53796] = t[53795] ^ n[53796];
assign t[53797] = t[53796] ^ n[53797];
assign t[53798] = t[53797] ^ n[53798];
assign t[53799] = t[53798] ^ n[53799];
assign t[53800] = t[53799] ^ n[53800];
assign t[53801] = t[53800] ^ n[53801];
assign t[53802] = t[53801] ^ n[53802];
assign t[53803] = t[53802] ^ n[53803];
assign t[53804] = t[53803] ^ n[53804];
assign t[53805] = t[53804] ^ n[53805];
assign t[53806] = t[53805] ^ n[53806];
assign t[53807] = t[53806] ^ n[53807];
assign t[53808] = t[53807] ^ n[53808];
assign t[53809] = t[53808] ^ n[53809];
assign t[53810] = t[53809] ^ n[53810];
assign t[53811] = t[53810] ^ n[53811];
assign t[53812] = t[53811] ^ n[53812];
assign t[53813] = t[53812] ^ n[53813];
assign t[53814] = t[53813] ^ n[53814];
assign t[53815] = t[53814] ^ n[53815];
assign t[53816] = t[53815] ^ n[53816];
assign t[53817] = t[53816] ^ n[53817];
assign t[53818] = t[53817] ^ n[53818];
assign t[53819] = t[53818] ^ n[53819];
assign t[53820] = t[53819] ^ n[53820];
assign t[53821] = t[53820] ^ n[53821];
assign t[53822] = t[53821] ^ n[53822];
assign t[53823] = t[53822] ^ n[53823];
assign t[53824] = t[53823] ^ n[53824];
assign t[53825] = t[53824] ^ n[53825];
assign t[53826] = t[53825] ^ n[53826];
assign t[53827] = t[53826] ^ n[53827];
assign t[53828] = t[53827] ^ n[53828];
assign t[53829] = t[53828] ^ n[53829];
assign t[53830] = t[53829] ^ n[53830];
assign t[53831] = t[53830] ^ n[53831];
assign t[53832] = t[53831] ^ n[53832];
assign t[53833] = t[53832] ^ n[53833];
assign t[53834] = t[53833] ^ n[53834];
assign t[53835] = t[53834] ^ n[53835];
assign t[53836] = t[53835] ^ n[53836];
assign t[53837] = t[53836] ^ n[53837];
assign t[53838] = t[53837] ^ n[53838];
assign t[53839] = t[53838] ^ n[53839];
assign t[53840] = t[53839] ^ n[53840];
assign t[53841] = t[53840] ^ n[53841];
assign t[53842] = t[53841] ^ n[53842];
assign t[53843] = t[53842] ^ n[53843];
assign t[53844] = t[53843] ^ n[53844];
assign t[53845] = t[53844] ^ n[53845];
assign t[53846] = t[53845] ^ n[53846];
assign t[53847] = t[53846] ^ n[53847];
assign t[53848] = t[53847] ^ n[53848];
assign t[53849] = t[53848] ^ n[53849];
assign t[53850] = t[53849] ^ n[53850];
assign t[53851] = t[53850] ^ n[53851];
assign t[53852] = t[53851] ^ n[53852];
assign t[53853] = t[53852] ^ n[53853];
assign t[53854] = t[53853] ^ n[53854];
assign t[53855] = t[53854] ^ n[53855];
assign t[53856] = t[53855] ^ n[53856];
assign t[53857] = t[53856] ^ n[53857];
assign t[53858] = t[53857] ^ n[53858];
assign t[53859] = t[53858] ^ n[53859];
assign t[53860] = t[53859] ^ n[53860];
assign t[53861] = t[53860] ^ n[53861];
assign t[53862] = t[53861] ^ n[53862];
assign t[53863] = t[53862] ^ n[53863];
assign t[53864] = t[53863] ^ n[53864];
assign t[53865] = t[53864] ^ n[53865];
assign t[53866] = t[53865] ^ n[53866];
assign t[53867] = t[53866] ^ n[53867];
assign t[53868] = t[53867] ^ n[53868];
assign t[53869] = t[53868] ^ n[53869];
assign t[53870] = t[53869] ^ n[53870];
assign t[53871] = t[53870] ^ n[53871];
assign t[53872] = t[53871] ^ n[53872];
assign t[53873] = t[53872] ^ n[53873];
assign t[53874] = t[53873] ^ n[53874];
assign t[53875] = t[53874] ^ n[53875];
assign t[53876] = t[53875] ^ n[53876];
assign t[53877] = t[53876] ^ n[53877];
assign t[53878] = t[53877] ^ n[53878];
assign t[53879] = t[53878] ^ n[53879];
assign t[53880] = t[53879] ^ n[53880];
assign t[53881] = t[53880] ^ n[53881];
assign t[53882] = t[53881] ^ n[53882];
assign t[53883] = t[53882] ^ n[53883];
assign t[53884] = t[53883] ^ n[53884];
assign t[53885] = t[53884] ^ n[53885];
assign t[53886] = t[53885] ^ n[53886];
assign t[53887] = t[53886] ^ n[53887];
assign t[53888] = t[53887] ^ n[53888];
assign t[53889] = t[53888] ^ n[53889];
assign t[53890] = t[53889] ^ n[53890];
assign t[53891] = t[53890] ^ n[53891];
assign t[53892] = t[53891] ^ n[53892];
assign t[53893] = t[53892] ^ n[53893];
assign t[53894] = t[53893] ^ n[53894];
assign t[53895] = t[53894] ^ n[53895];
assign t[53896] = t[53895] ^ n[53896];
assign t[53897] = t[53896] ^ n[53897];
assign t[53898] = t[53897] ^ n[53898];
assign t[53899] = t[53898] ^ n[53899];
assign t[53900] = t[53899] ^ n[53900];
assign t[53901] = t[53900] ^ n[53901];
assign t[53902] = t[53901] ^ n[53902];
assign t[53903] = t[53902] ^ n[53903];
assign t[53904] = t[53903] ^ n[53904];
assign t[53905] = t[53904] ^ n[53905];
assign t[53906] = t[53905] ^ n[53906];
assign t[53907] = t[53906] ^ n[53907];
assign t[53908] = t[53907] ^ n[53908];
assign t[53909] = t[53908] ^ n[53909];
assign t[53910] = t[53909] ^ n[53910];
assign t[53911] = t[53910] ^ n[53911];
assign t[53912] = t[53911] ^ n[53912];
assign t[53913] = t[53912] ^ n[53913];
assign t[53914] = t[53913] ^ n[53914];
assign t[53915] = t[53914] ^ n[53915];
assign t[53916] = t[53915] ^ n[53916];
assign t[53917] = t[53916] ^ n[53917];
assign t[53918] = t[53917] ^ n[53918];
assign t[53919] = t[53918] ^ n[53919];
assign t[53920] = t[53919] ^ n[53920];
assign t[53921] = t[53920] ^ n[53921];
assign t[53922] = t[53921] ^ n[53922];
assign t[53923] = t[53922] ^ n[53923];
assign t[53924] = t[53923] ^ n[53924];
assign t[53925] = t[53924] ^ n[53925];
assign t[53926] = t[53925] ^ n[53926];
assign t[53927] = t[53926] ^ n[53927];
assign t[53928] = t[53927] ^ n[53928];
assign t[53929] = t[53928] ^ n[53929];
assign t[53930] = t[53929] ^ n[53930];
assign t[53931] = t[53930] ^ n[53931];
assign t[53932] = t[53931] ^ n[53932];
assign t[53933] = t[53932] ^ n[53933];
assign t[53934] = t[53933] ^ n[53934];
assign t[53935] = t[53934] ^ n[53935];
assign t[53936] = t[53935] ^ n[53936];
assign t[53937] = t[53936] ^ n[53937];
assign t[53938] = t[53937] ^ n[53938];
assign t[53939] = t[53938] ^ n[53939];
assign t[53940] = t[53939] ^ n[53940];
assign t[53941] = t[53940] ^ n[53941];
assign t[53942] = t[53941] ^ n[53942];
assign t[53943] = t[53942] ^ n[53943];
assign t[53944] = t[53943] ^ n[53944];
assign t[53945] = t[53944] ^ n[53945];
assign t[53946] = t[53945] ^ n[53946];
assign t[53947] = t[53946] ^ n[53947];
assign t[53948] = t[53947] ^ n[53948];
assign t[53949] = t[53948] ^ n[53949];
assign t[53950] = t[53949] ^ n[53950];
assign t[53951] = t[53950] ^ n[53951];
assign t[53952] = t[53951] ^ n[53952];
assign t[53953] = t[53952] ^ n[53953];
assign t[53954] = t[53953] ^ n[53954];
assign t[53955] = t[53954] ^ n[53955];
assign t[53956] = t[53955] ^ n[53956];
assign t[53957] = t[53956] ^ n[53957];
assign t[53958] = t[53957] ^ n[53958];
assign t[53959] = t[53958] ^ n[53959];
assign t[53960] = t[53959] ^ n[53960];
assign t[53961] = t[53960] ^ n[53961];
assign t[53962] = t[53961] ^ n[53962];
assign t[53963] = t[53962] ^ n[53963];
assign t[53964] = t[53963] ^ n[53964];
assign t[53965] = t[53964] ^ n[53965];
assign t[53966] = t[53965] ^ n[53966];
assign t[53967] = t[53966] ^ n[53967];
assign t[53968] = t[53967] ^ n[53968];
assign t[53969] = t[53968] ^ n[53969];
assign t[53970] = t[53969] ^ n[53970];
assign t[53971] = t[53970] ^ n[53971];
assign t[53972] = t[53971] ^ n[53972];
assign t[53973] = t[53972] ^ n[53973];
assign t[53974] = t[53973] ^ n[53974];
assign t[53975] = t[53974] ^ n[53975];
assign t[53976] = t[53975] ^ n[53976];
assign t[53977] = t[53976] ^ n[53977];
assign t[53978] = t[53977] ^ n[53978];
assign t[53979] = t[53978] ^ n[53979];
assign t[53980] = t[53979] ^ n[53980];
assign t[53981] = t[53980] ^ n[53981];
assign t[53982] = t[53981] ^ n[53982];
assign t[53983] = t[53982] ^ n[53983];
assign t[53984] = t[53983] ^ n[53984];
assign t[53985] = t[53984] ^ n[53985];
assign t[53986] = t[53985] ^ n[53986];
assign t[53987] = t[53986] ^ n[53987];
assign t[53988] = t[53987] ^ n[53988];
assign t[53989] = t[53988] ^ n[53989];
assign t[53990] = t[53989] ^ n[53990];
assign t[53991] = t[53990] ^ n[53991];
assign t[53992] = t[53991] ^ n[53992];
assign t[53993] = t[53992] ^ n[53993];
assign t[53994] = t[53993] ^ n[53994];
assign t[53995] = t[53994] ^ n[53995];
assign t[53996] = t[53995] ^ n[53996];
assign t[53997] = t[53996] ^ n[53997];
assign t[53998] = t[53997] ^ n[53998];
assign t[53999] = t[53998] ^ n[53999];
assign t[54000] = t[53999] ^ n[54000];
assign t[54001] = t[54000] ^ n[54001];
assign t[54002] = t[54001] ^ n[54002];
assign t[54003] = t[54002] ^ n[54003];
assign t[54004] = t[54003] ^ n[54004];
assign t[54005] = t[54004] ^ n[54005];
assign t[54006] = t[54005] ^ n[54006];
assign t[54007] = t[54006] ^ n[54007];
assign t[54008] = t[54007] ^ n[54008];
assign t[54009] = t[54008] ^ n[54009];
assign t[54010] = t[54009] ^ n[54010];
assign t[54011] = t[54010] ^ n[54011];
assign t[54012] = t[54011] ^ n[54012];
assign t[54013] = t[54012] ^ n[54013];
assign t[54014] = t[54013] ^ n[54014];
assign t[54015] = t[54014] ^ n[54015];
assign t[54016] = t[54015] ^ n[54016];
assign t[54017] = t[54016] ^ n[54017];
assign t[54018] = t[54017] ^ n[54018];
assign t[54019] = t[54018] ^ n[54019];
assign t[54020] = t[54019] ^ n[54020];
assign t[54021] = t[54020] ^ n[54021];
assign t[54022] = t[54021] ^ n[54022];
assign t[54023] = t[54022] ^ n[54023];
assign t[54024] = t[54023] ^ n[54024];
assign t[54025] = t[54024] ^ n[54025];
assign t[54026] = t[54025] ^ n[54026];
assign t[54027] = t[54026] ^ n[54027];
assign t[54028] = t[54027] ^ n[54028];
assign t[54029] = t[54028] ^ n[54029];
assign t[54030] = t[54029] ^ n[54030];
assign t[54031] = t[54030] ^ n[54031];
assign t[54032] = t[54031] ^ n[54032];
assign t[54033] = t[54032] ^ n[54033];
assign t[54034] = t[54033] ^ n[54034];
assign t[54035] = t[54034] ^ n[54035];
assign t[54036] = t[54035] ^ n[54036];
assign t[54037] = t[54036] ^ n[54037];
assign t[54038] = t[54037] ^ n[54038];
assign t[54039] = t[54038] ^ n[54039];
assign t[54040] = t[54039] ^ n[54040];
assign t[54041] = t[54040] ^ n[54041];
assign t[54042] = t[54041] ^ n[54042];
assign t[54043] = t[54042] ^ n[54043];
assign t[54044] = t[54043] ^ n[54044];
assign t[54045] = t[54044] ^ n[54045];
assign t[54046] = t[54045] ^ n[54046];
assign t[54047] = t[54046] ^ n[54047];
assign t[54048] = t[54047] ^ n[54048];
assign t[54049] = t[54048] ^ n[54049];
assign t[54050] = t[54049] ^ n[54050];
assign t[54051] = t[54050] ^ n[54051];
assign t[54052] = t[54051] ^ n[54052];
assign t[54053] = t[54052] ^ n[54053];
assign t[54054] = t[54053] ^ n[54054];
assign t[54055] = t[54054] ^ n[54055];
assign t[54056] = t[54055] ^ n[54056];
assign t[54057] = t[54056] ^ n[54057];
assign t[54058] = t[54057] ^ n[54058];
assign t[54059] = t[54058] ^ n[54059];
assign t[54060] = t[54059] ^ n[54060];
assign t[54061] = t[54060] ^ n[54061];
assign t[54062] = t[54061] ^ n[54062];
assign t[54063] = t[54062] ^ n[54063];
assign t[54064] = t[54063] ^ n[54064];
assign t[54065] = t[54064] ^ n[54065];
assign t[54066] = t[54065] ^ n[54066];
assign t[54067] = t[54066] ^ n[54067];
assign t[54068] = t[54067] ^ n[54068];
assign t[54069] = t[54068] ^ n[54069];
assign t[54070] = t[54069] ^ n[54070];
assign t[54071] = t[54070] ^ n[54071];
assign t[54072] = t[54071] ^ n[54072];
assign t[54073] = t[54072] ^ n[54073];
assign t[54074] = t[54073] ^ n[54074];
assign t[54075] = t[54074] ^ n[54075];
assign t[54076] = t[54075] ^ n[54076];
assign t[54077] = t[54076] ^ n[54077];
assign t[54078] = t[54077] ^ n[54078];
assign t[54079] = t[54078] ^ n[54079];
assign t[54080] = t[54079] ^ n[54080];
assign t[54081] = t[54080] ^ n[54081];
assign t[54082] = t[54081] ^ n[54082];
assign t[54083] = t[54082] ^ n[54083];
assign t[54084] = t[54083] ^ n[54084];
assign t[54085] = t[54084] ^ n[54085];
assign t[54086] = t[54085] ^ n[54086];
assign t[54087] = t[54086] ^ n[54087];
assign t[54088] = t[54087] ^ n[54088];
assign t[54089] = t[54088] ^ n[54089];
assign t[54090] = t[54089] ^ n[54090];
assign t[54091] = t[54090] ^ n[54091];
assign t[54092] = t[54091] ^ n[54092];
assign t[54093] = t[54092] ^ n[54093];
assign t[54094] = t[54093] ^ n[54094];
assign t[54095] = t[54094] ^ n[54095];
assign t[54096] = t[54095] ^ n[54096];
assign t[54097] = t[54096] ^ n[54097];
assign t[54098] = t[54097] ^ n[54098];
assign t[54099] = t[54098] ^ n[54099];
assign t[54100] = t[54099] ^ n[54100];
assign t[54101] = t[54100] ^ n[54101];
assign t[54102] = t[54101] ^ n[54102];
assign t[54103] = t[54102] ^ n[54103];
assign t[54104] = t[54103] ^ n[54104];
assign t[54105] = t[54104] ^ n[54105];
assign t[54106] = t[54105] ^ n[54106];
assign t[54107] = t[54106] ^ n[54107];
assign t[54108] = t[54107] ^ n[54108];
assign t[54109] = t[54108] ^ n[54109];
assign t[54110] = t[54109] ^ n[54110];
assign t[54111] = t[54110] ^ n[54111];
assign t[54112] = t[54111] ^ n[54112];
assign t[54113] = t[54112] ^ n[54113];
assign t[54114] = t[54113] ^ n[54114];
assign t[54115] = t[54114] ^ n[54115];
assign t[54116] = t[54115] ^ n[54116];
assign t[54117] = t[54116] ^ n[54117];
assign t[54118] = t[54117] ^ n[54118];
assign t[54119] = t[54118] ^ n[54119];
assign t[54120] = t[54119] ^ n[54120];
assign t[54121] = t[54120] ^ n[54121];
assign t[54122] = t[54121] ^ n[54122];
assign t[54123] = t[54122] ^ n[54123];
assign t[54124] = t[54123] ^ n[54124];
assign t[54125] = t[54124] ^ n[54125];
assign t[54126] = t[54125] ^ n[54126];
assign t[54127] = t[54126] ^ n[54127];
assign t[54128] = t[54127] ^ n[54128];
assign t[54129] = t[54128] ^ n[54129];
assign t[54130] = t[54129] ^ n[54130];
assign t[54131] = t[54130] ^ n[54131];
assign t[54132] = t[54131] ^ n[54132];
assign t[54133] = t[54132] ^ n[54133];
assign t[54134] = t[54133] ^ n[54134];
assign t[54135] = t[54134] ^ n[54135];
assign t[54136] = t[54135] ^ n[54136];
assign t[54137] = t[54136] ^ n[54137];
assign t[54138] = t[54137] ^ n[54138];
assign t[54139] = t[54138] ^ n[54139];
assign t[54140] = t[54139] ^ n[54140];
assign t[54141] = t[54140] ^ n[54141];
assign t[54142] = t[54141] ^ n[54142];
assign t[54143] = t[54142] ^ n[54143];
assign t[54144] = t[54143] ^ n[54144];
assign t[54145] = t[54144] ^ n[54145];
assign t[54146] = t[54145] ^ n[54146];
assign t[54147] = t[54146] ^ n[54147];
assign t[54148] = t[54147] ^ n[54148];
assign t[54149] = t[54148] ^ n[54149];
assign t[54150] = t[54149] ^ n[54150];
assign t[54151] = t[54150] ^ n[54151];
assign t[54152] = t[54151] ^ n[54152];
assign t[54153] = t[54152] ^ n[54153];
assign t[54154] = t[54153] ^ n[54154];
assign t[54155] = t[54154] ^ n[54155];
assign t[54156] = t[54155] ^ n[54156];
assign t[54157] = t[54156] ^ n[54157];
assign t[54158] = t[54157] ^ n[54158];
assign t[54159] = t[54158] ^ n[54159];
assign t[54160] = t[54159] ^ n[54160];
assign t[54161] = t[54160] ^ n[54161];
assign t[54162] = t[54161] ^ n[54162];
assign t[54163] = t[54162] ^ n[54163];
assign t[54164] = t[54163] ^ n[54164];
assign t[54165] = t[54164] ^ n[54165];
assign t[54166] = t[54165] ^ n[54166];
assign t[54167] = t[54166] ^ n[54167];
assign t[54168] = t[54167] ^ n[54168];
assign t[54169] = t[54168] ^ n[54169];
assign t[54170] = t[54169] ^ n[54170];
assign t[54171] = t[54170] ^ n[54171];
assign t[54172] = t[54171] ^ n[54172];
assign t[54173] = t[54172] ^ n[54173];
assign t[54174] = t[54173] ^ n[54174];
assign t[54175] = t[54174] ^ n[54175];
assign t[54176] = t[54175] ^ n[54176];
assign t[54177] = t[54176] ^ n[54177];
assign t[54178] = t[54177] ^ n[54178];
assign t[54179] = t[54178] ^ n[54179];
assign t[54180] = t[54179] ^ n[54180];
assign t[54181] = t[54180] ^ n[54181];
assign t[54182] = t[54181] ^ n[54182];
assign t[54183] = t[54182] ^ n[54183];
assign t[54184] = t[54183] ^ n[54184];
assign t[54185] = t[54184] ^ n[54185];
assign t[54186] = t[54185] ^ n[54186];
assign t[54187] = t[54186] ^ n[54187];
assign t[54188] = t[54187] ^ n[54188];
assign t[54189] = t[54188] ^ n[54189];
assign t[54190] = t[54189] ^ n[54190];
assign t[54191] = t[54190] ^ n[54191];
assign t[54192] = t[54191] ^ n[54192];
assign t[54193] = t[54192] ^ n[54193];
assign t[54194] = t[54193] ^ n[54194];
assign t[54195] = t[54194] ^ n[54195];
assign t[54196] = t[54195] ^ n[54196];
assign t[54197] = t[54196] ^ n[54197];
assign t[54198] = t[54197] ^ n[54198];
assign t[54199] = t[54198] ^ n[54199];
assign t[54200] = t[54199] ^ n[54200];
assign t[54201] = t[54200] ^ n[54201];
assign t[54202] = t[54201] ^ n[54202];
assign t[54203] = t[54202] ^ n[54203];
assign t[54204] = t[54203] ^ n[54204];
assign t[54205] = t[54204] ^ n[54205];
assign t[54206] = t[54205] ^ n[54206];
assign t[54207] = t[54206] ^ n[54207];
assign t[54208] = t[54207] ^ n[54208];
assign t[54209] = t[54208] ^ n[54209];
assign t[54210] = t[54209] ^ n[54210];
assign t[54211] = t[54210] ^ n[54211];
assign t[54212] = t[54211] ^ n[54212];
assign t[54213] = t[54212] ^ n[54213];
assign t[54214] = t[54213] ^ n[54214];
assign t[54215] = t[54214] ^ n[54215];
assign t[54216] = t[54215] ^ n[54216];
assign t[54217] = t[54216] ^ n[54217];
assign t[54218] = t[54217] ^ n[54218];
assign t[54219] = t[54218] ^ n[54219];
assign t[54220] = t[54219] ^ n[54220];
assign t[54221] = t[54220] ^ n[54221];
assign t[54222] = t[54221] ^ n[54222];
assign t[54223] = t[54222] ^ n[54223];
assign t[54224] = t[54223] ^ n[54224];
assign t[54225] = t[54224] ^ n[54225];
assign t[54226] = t[54225] ^ n[54226];
assign t[54227] = t[54226] ^ n[54227];
assign t[54228] = t[54227] ^ n[54228];
assign t[54229] = t[54228] ^ n[54229];
assign t[54230] = t[54229] ^ n[54230];
assign t[54231] = t[54230] ^ n[54231];
assign t[54232] = t[54231] ^ n[54232];
assign t[54233] = t[54232] ^ n[54233];
assign t[54234] = t[54233] ^ n[54234];
assign t[54235] = t[54234] ^ n[54235];
assign t[54236] = t[54235] ^ n[54236];
assign t[54237] = t[54236] ^ n[54237];
assign t[54238] = t[54237] ^ n[54238];
assign t[54239] = t[54238] ^ n[54239];
assign t[54240] = t[54239] ^ n[54240];
assign t[54241] = t[54240] ^ n[54241];
assign t[54242] = t[54241] ^ n[54242];
assign t[54243] = t[54242] ^ n[54243];
assign t[54244] = t[54243] ^ n[54244];
assign t[54245] = t[54244] ^ n[54245];
assign t[54246] = t[54245] ^ n[54246];
assign t[54247] = t[54246] ^ n[54247];
assign t[54248] = t[54247] ^ n[54248];
assign t[54249] = t[54248] ^ n[54249];
assign t[54250] = t[54249] ^ n[54250];
assign t[54251] = t[54250] ^ n[54251];
assign t[54252] = t[54251] ^ n[54252];
assign t[54253] = t[54252] ^ n[54253];
assign t[54254] = t[54253] ^ n[54254];
assign t[54255] = t[54254] ^ n[54255];
assign t[54256] = t[54255] ^ n[54256];
assign t[54257] = t[54256] ^ n[54257];
assign t[54258] = t[54257] ^ n[54258];
assign t[54259] = t[54258] ^ n[54259];
assign t[54260] = t[54259] ^ n[54260];
assign t[54261] = t[54260] ^ n[54261];
assign t[54262] = t[54261] ^ n[54262];
assign t[54263] = t[54262] ^ n[54263];
assign t[54264] = t[54263] ^ n[54264];
assign t[54265] = t[54264] ^ n[54265];
assign t[54266] = t[54265] ^ n[54266];
assign t[54267] = t[54266] ^ n[54267];
assign t[54268] = t[54267] ^ n[54268];
assign t[54269] = t[54268] ^ n[54269];
assign t[54270] = t[54269] ^ n[54270];
assign t[54271] = t[54270] ^ n[54271];
assign t[54272] = t[54271] ^ n[54272];
assign t[54273] = t[54272] ^ n[54273];
assign t[54274] = t[54273] ^ n[54274];
assign t[54275] = t[54274] ^ n[54275];
assign t[54276] = t[54275] ^ n[54276];
assign t[54277] = t[54276] ^ n[54277];
assign t[54278] = t[54277] ^ n[54278];
assign t[54279] = t[54278] ^ n[54279];
assign t[54280] = t[54279] ^ n[54280];
assign t[54281] = t[54280] ^ n[54281];
assign t[54282] = t[54281] ^ n[54282];
assign t[54283] = t[54282] ^ n[54283];
assign t[54284] = t[54283] ^ n[54284];
assign t[54285] = t[54284] ^ n[54285];
assign t[54286] = t[54285] ^ n[54286];
assign t[54287] = t[54286] ^ n[54287];
assign t[54288] = t[54287] ^ n[54288];
assign t[54289] = t[54288] ^ n[54289];
assign t[54290] = t[54289] ^ n[54290];
assign t[54291] = t[54290] ^ n[54291];
assign t[54292] = t[54291] ^ n[54292];
assign t[54293] = t[54292] ^ n[54293];
assign t[54294] = t[54293] ^ n[54294];
assign t[54295] = t[54294] ^ n[54295];
assign t[54296] = t[54295] ^ n[54296];
assign t[54297] = t[54296] ^ n[54297];
assign t[54298] = t[54297] ^ n[54298];
assign t[54299] = t[54298] ^ n[54299];
assign t[54300] = t[54299] ^ n[54300];
assign t[54301] = t[54300] ^ n[54301];
assign t[54302] = t[54301] ^ n[54302];
assign t[54303] = t[54302] ^ n[54303];
assign t[54304] = t[54303] ^ n[54304];
assign t[54305] = t[54304] ^ n[54305];
assign t[54306] = t[54305] ^ n[54306];
assign t[54307] = t[54306] ^ n[54307];
assign t[54308] = t[54307] ^ n[54308];
assign t[54309] = t[54308] ^ n[54309];
assign t[54310] = t[54309] ^ n[54310];
assign t[54311] = t[54310] ^ n[54311];
assign t[54312] = t[54311] ^ n[54312];
assign t[54313] = t[54312] ^ n[54313];
assign t[54314] = t[54313] ^ n[54314];
assign t[54315] = t[54314] ^ n[54315];
assign t[54316] = t[54315] ^ n[54316];
assign t[54317] = t[54316] ^ n[54317];
assign t[54318] = t[54317] ^ n[54318];
assign t[54319] = t[54318] ^ n[54319];
assign t[54320] = t[54319] ^ n[54320];
assign t[54321] = t[54320] ^ n[54321];
assign t[54322] = t[54321] ^ n[54322];
assign t[54323] = t[54322] ^ n[54323];
assign t[54324] = t[54323] ^ n[54324];
assign t[54325] = t[54324] ^ n[54325];
assign t[54326] = t[54325] ^ n[54326];
assign t[54327] = t[54326] ^ n[54327];
assign t[54328] = t[54327] ^ n[54328];
assign t[54329] = t[54328] ^ n[54329];
assign t[54330] = t[54329] ^ n[54330];
assign t[54331] = t[54330] ^ n[54331];
assign t[54332] = t[54331] ^ n[54332];
assign t[54333] = t[54332] ^ n[54333];
assign t[54334] = t[54333] ^ n[54334];
assign t[54335] = t[54334] ^ n[54335];
assign t[54336] = t[54335] ^ n[54336];
assign t[54337] = t[54336] ^ n[54337];
assign t[54338] = t[54337] ^ n[54338];
assign t[54339] = t[54338] ^ n[54339];
assign t[54340] = t[54339] ^ n[54340];
assign t[54341] = t[54340] ^ n[54341];
assign t[54342] = t[54341] ^ n[54342];
assign t[54343] = t[54342] ^ n[54343];
assign t[54344] = t[54343] ^ n[54344];
assign t[54345] = t[54344] ^ n[54345];
assign t[54346] = t[54345] ^ n[54346];
assign t[54347] = t[54346] ^ n[54347];
assign t[54348] = t[54347] ^ n[54348];
assign t[54349] = t[54348] ^ n[54349];
assign t[54350] = t[54349] ^ n[54350];
assign t[54351] = t[54350] ^ n[54351];
assign t[54352] = t[54351] ^ n[54352];
assign t[54353] = t[54352] ^ n[54353];
assign t[54354] = t[54353] ^ n[54354];
assign t[54355] = t[54354] ^ n[54355];
assign t[54356] = t[54355] ^ n[54356];
assign t[54357] = t[54356] ^ n[54357];
assign t[54358] = t[54357] ^ n[54358];
assign t[54359] = t[54358] ^ n[54359];
assign t[54360] = t[54359] ^ n[54360];
assign t[54361] = t[54360] ^ n[54361];
assign t[54362] = t[54361] ^ n[54362];
assign t[54363] = t[54362] ^ n[54363];
assign t[54364] = t[54363] ^ n[54364];
assign t[54365] = t[54364] ^ n[54365];
assign t[54366] = t[54365] ^ n[54366];
assign t[54367] = t[54366] ^ n[54367];
assign t[54368] = t[54367] ^ n[54368];
assign t[54369] = t[54368] ^ n[54369];
assign t[54370] = t[54369] ^ n[54370];
assign t[54371] = t[54370] ^ n[54371];
assign t[54372] = t[54371] ^ n[54372];
assign t[54373] = t[54372] ^ n[54373];
assign t[54374] = t[54373] ^ n[54374];
assign t[54375] = t[54374] ^ n[54375];
assign t[54376] = t[54375] ^ n[54376];
assign t[54377] = t[54376] ^ n[54377];
assign t[54378] = t[54377] ^ n[54378];
assign t[54379] = t[54378] ^ n[54379];
assign t[54380] = t[54379] ^ n[54380];
assign t[54381] = t[54380] ^ n[54381];
assign t[54382] = t[54381] ^ n[54382];
assign t[54383] = t[54382] ^ n[54383];
assign t[54384] = t[54383] ^ n[54384];
assign t[54385] = t[54384] ^ n[54385];
assign t[54386] = t[54385] ^ n[54386];
assign t[54387] = t[54386] ^ n[54387];
assign t[54388] = t[54387] ^ n[54388];
assign t[54389] = t[54388] ^ n[54389];
assign t[54390] = t[54389] ^ n[54390];
assign t[54391] = t[54390] ^ n[54391];
assign t[54392] = t[54391] ^ n[54392];
assign t[54393] = t[54392] ^ n[54393];
assign t[54394] = t[54393] ^ n[54394];
assign t[54395] = t[54394] ^ n[54395];
assign t[54396] = t[54395] ^ n[54396];
assign t[54397] = t[54396] ^ n[54397];
assign t[54398] = t[54397] ^ n[54398];
assign t[54399] = t[54398] ^ n[54399];
assign t[54400] = t[54399] ^ n[54400];
assign t[54401] = t[54400] ^ n[54401];
assign t[54402] = t[54401] ^ n[54402];
assign t[54403] = t[54402] ^ n[54403];
assign t[54404] = t[54403] ^ n[54404];
assign t[54405] = t[54404] ^ n[54405];
assign t[54406] = t[54405] ^ n[54406];
assign t[54407] = t[54406] ^ n[54407];
assign t[54408] = t[54407] ^ n[54408];
assign t[54409] = t[54408] ^ n[54409];
assign t[54410] = t[54409] ^ n[54410];
assign t[54411] = t[54410] ^ n[54411];
assign t[54412] = t[54411] ^ n[54412];
assign t[54413] = t[54412] ^ n[54413];
assign t[54414] = t[54413] ^ n[54414];
assign t[54415] = t[54414] ^ n[54415];
assign t[54416] = t[54415] ^ n[54416];
assign t[54417] = t[54416] ^ n[54417];
assign t[54418] = t[54417] ^ n[54418];
assign t[54419] = t[54418] ^ n[54419];
assign t[54420] = t[54419] ^ n[54420];
assign t[54421] = t[54420] ^ n[54421];
assign t[54422] = t[54421] ^ n[54422];
assign t[54423] = t[54422] ^ n[54423];
assign t[54424] = t[54423] ^ n[54424];
assign t[54425] = t[54424] ^ n[54425];
assign t[54426] = t[54425] ^ n[54426];
assign t[54427] = t[54426] ^ n[54427];
assign t[54428] = t[54427] ^ n[54428];
assign t[54429] = t[54428] ^ n[54429];
assign t[54430] = t[54429] ^ n[54430];
assign t[54431] = t[54430] ^ n[54431];
assign t[54432] = t[54431] ^ n[54432];
assign t[54433] = t[54432] ^ n[54433];
assign t[54434] = t[54433] ^ n[54434];
assign t[54435] = t[54434] ^ n[54435];
assign t[54436] = t[54435] ^ n[54436];
assign t[54437] = t[54436] ^ n[54437];
assign t[54438] = t[54437] ^ n[54438];
assign t[54439] = t[54438] ^ n[54439];
assign t[54440] = t[54439] ^ n[54440];
assign t[54441] = t[54440] ^ n[54441];
assign t[54442] = t[54441] ^ n[54442];
assign t[54443] = t[54442] ^ n[54443];
assign t[54444] = t[54443] ^ n[54444];
assign t[54445] = t[54444] ^ n[54445];
assign t[54446] = t[54445] ^ n[54446];
assign t[54447] = t[54446] ^ n[54447];
assign t[54448] = t[54447] ^ n[54448];
assign t[54449] = t[54448] ^ n[54449];
assign t[54450] = t[54449] ^ n[54450];
assign t[54451] = t[54450] ^ n[54451];
assign t[54452] = t[54451] ^ n[54452];
assign t[54453] = t[54452] ^ n[54453];
assign t[54454] = t[54453] ^ n[54454];
assign t[54455] = t[54454] ^ n[54455];
assign t[54456] = t[54455] ^ n[54456];
assign t[54457] = t[54456] ^ n[54457];
assign t[54458] = t[54457] ^ n[54458];
assign t[54459] = t[54458] ^ n[54459];
assign t[54460] = t[54459] ^ n[54460];
assign t[54461] = t[54460] ^ n[54461];
assign t[54462] = t[54461] ^ n[54462];
assign t[54463] = t[54462] ^ n[54463];
assign t[54464] = t[54463] ^ n[54464];
assign t[54465] = t[54464] ^ n[54465];
assign t[54466] = t[54465] ^ n[54466];
assign t[54467] = t[54466] ^ n[54467];
assign t[54468] = t[54467] ^ n[54468];
assign t[54469] = t[54468] ^ n[54469];
assign t[54470] = t[54469] ^ n[54470];
assign t[54471] = t[54470] ^ n[54471];
assign t[54472] = t[54471] ^ n[54472];
assign t[54473] = t[54472] ^ n[54473];
assign t[54474] = t[54473] ^ n[54474];
assign t[54475] = t[54474] ^ n[54475];
assign t[54476] = t[54475] ^ n[54476];
assign t[54477] = t[54476] ^ n[54477];
assign t[54478] = t[54477] ^ n[54478];
assign t[54479] = t[54478] ^ n[54479];
assign t[54480] = t[54479] ^ n[54480];
assign t[54481] = t[54480] ^ n[54481];
assign t[54482] = t[54481] ^ n[54482];
assign t[54483] = t[54482] ^ n[54483];
assign t[54484] = t[54483] ^ n[54484];
assign t[54485] = t[54484] ^ n[54485];
assign t[54486] = t[54485] ^ n[54486];
assign t[54487] = t[54486] ^ n[54487];
assign t[54488] = t[54487] ^ n[54488];
assign t[54489] = t[54488] ^ n[54489];
assign t[54490] = t[54489] ^ n[54490];
assign t[54491] = t[54490] ^ n[54491];
assign t[54492] = t[54491] ^ n[54492];
assign t[54493] = t[54492] ^ n[54493];
assign t[54494] = t[54493] ^ n[54494];
assign t[54495] = t[54494] ^ n[54495];
assign t[54496] = t[54495] ^ n[54496];
assign t[54497] = t[54496] ^ n[54497];
assign t[54498] = t[54497] ^ n[54498];
assign t[54499] = t[54498] ^ n[54499];
assign t[54500] = t[54499] ^ n[54500];
assign t[54501] = t[54500] ^ n[54501];
assign t[54502] = t[54501] ^ n[54502];
assign t[54503] = t[54502] ^ n[54503];
assign t[54504] = t[54503] ^ n[54504];
assign t[54505] = t[54504] ^ n[54505];
assign t[54506] = t[54505] ^ n[54506];
assign t[54507] = t[54506] ^ n[54507];
assign t[54508] = t[54507] ^ n[54508];
assign t[54509] = t[54508] ^ n[54509];
assign t[54510] = t[54509] ^ n[54510];
assign t[54511] = t[54510] ^ n[54511];
assign t[54512] = t[54511] ^ n[54512];
assign t[54513] = t[54512] ^ n[54513];
assign t[54514] = t[54513] ^ n[54514];
assign t[54515] = t[54514] ^ n[54515];
assign t[54516] = t[54515] ^ n[54516];
assign t[54517] = t[54516] ^ n[54517];
assign t[54518] = t[54517] ^ n[54518];
assign t[54519] = t[54518] ^ n[54519];
assign t[54520] = t[54519] ^ n[54520];
assign t[54521] = t[54520] ^ n[54521];
assign t[54522] = t[54521] ^ n[54522];
assign t[54523] = t[54522] ^ n[54523];
assign t[54524] = t[54523] ^ n[54524];
assign t[54525] = t[54524] ^ n[54525];
assign t[54526] = t[54525] ^ n[54526];
assign t[54527] = t[54526] ^ n[54527];
assign t[54528] = t[54527] ^ n[54528];
assign t[54529] = t[54528] ^ n[54529];
assign t[54530] = t[54529] ^ n[54530];
assign t[54531] = t[54530] ^ n[54531];
assign t[54532] = t[54531] ^ n[54532];
assign t[54533] = t[54532] ^ n[54533];
assign t[54534] = t[54533] ^ n[54534];
assign t[54535] = t[54534] ^ n[54535];
assign t[54536] = t[54535] ^ n[54536];
assign t[54537] = t[54536] ^ n[54537];
assign t[54538] = t[54537] ^ n[54538];
assign t[54539] = t[54538] ^ n[54539];
assign t[54540] = t[54539] ^ n[54540];
assign t[54541] = t[54540] ^ n[54541];
assign t[54542] = t[54541] ^ n[54542];
assign t[54543] = t[54542] ^ n[54543];
assign t[54544] = t[54543] ^ n[54544];
assign t[54545] = t[54544] ^ n[54545];
assign t[54546] = t[54545] ^ n[54546];
assign t[54547] = t[54546] ^ n[54547];
assign t[54548] = t[54547] ^ n[54548];
assign t[54549] = t[54548] ^ n[54549];
assign t[54550] = t[54549] ^ n[54550];
assign t[54551] = t[54550] ^ n[54551];
assign t[54552] = t[54551] ^ n[54552];
assign t[54553] = t[54552] ^ n[54553];
assign t[54554] = t[54553] ^ n[54554];
assign t[54555] = t[54554] ^ n[54555];
assign t[54556] = t[54555] ^ n[54556];
assign t[54557] = t[54556] ^ n[54557];
assign t[54558] = t[54557] ^ n[54558];
assign t[54559] = t[54558] ^ n[54559];
assign t[54560] = t[54559] ^ n[54560];
assign t[54561] = t[54560] ^ n[54561];
assign t[54562] = t[54561] ^ n[54562];
assign t[54563] = t[54562] ^ n[54563];
assign t[54564] = t[54563] ^ n[54564];
assign t[54565] = t[54564] ^ n[54565];
assign t[54566] = t[54565] ^ n[54566];
assign t[54567] = t[54566] ^ n[54567];
assign t[54568] = t[54567] ^ n[54568];
assign t[54569] = t[54568] ^ n[54569];
assign t[54570] = t[54569] ^ n[54570];
assign t[54571] = t[54570] ^ n[54571];
assign t[54572] = t[54571] ^ n[54572];
assign t[54573] = t[54572] ^ n[54573];
assign t[54574] = t[54573] ^ n[54574];
assign t[54575] = t[54574] ^ n[54575];
assign t[54576] = t[54575] ^ n[54576];
assign t[54577] = t[54576] ^ n[54577];
assign t[54578] = t[54577] ^ n[54578];
assign t[54579] = t[54578] ^ n[54579];
assign t[54580] = t[54579] ^ n[54580];
assign t[54581] = t[54580] ^ n[54581];
assign t[54582] = t[54581] ^ n[54582];
assign t[54583] = t[54582] ^ n[54583];
assign t[54584] = t[54583] ^ n[54584];
assign t[54585] = t[54584] ^ n[54585];
assign t[54586] = t[54585] ^ n[54586];
assign t[54587] = t[54586] ^ n[54587];
assign t[54588] = t[54587] ^ n[54588];
assign t[54589] = t[54588] ^ n[54589];
assign t[54590] = t[54589] ^ n[54590];
assign t[54591] = t[54590] ^ n[54591];
assign t[54592] = t[54591] ^ n[54592];
assign t[54593] = t[54592] ^ n[54593];
assign t[54594] = t[54593] ^ n[54594];
assign t[54595] = t[54594] ^ n[54595];
assign t[54596] = t[54595] ^ n[54596];
assign t[54597] = t[54596] ^ n[54597];
assign t[54598] = t[54597] ^ n[54598];
assign t[54599] = t[54598] ^ n[54599];
assign t[54600] = t[54599] ^ n[54600];
assign t[54601] = t[54600] ^ n[54601];
assign t[54602] = t[54601] ^ n[54602];
assign t[54603] = t[54602] ^ n[54603];
assign t[54604] = t[54603] ^ n[54604];
assign t[54605] = t[54604] ^ n[54605];
assign t[54606] = t[54605] ^ n[54606];
assign t[54607] = t[54606] ^ n[54607];
assign t[54608] = t[54607] ^ n[54608];
assign t[54609] = t[54608] ^ n[54609];
assign t[54610] = t[54609] ^ n[54610];
assign t[54611] = t[54610] ^ n[54611];
assign t[54612] = t[54611] ^ n[54612];
assign t[54613] = t[54612] ^ n[54613];
assign t[54614] = t[54613] ^ n[54614];
assign t[54615] = t[54614] ^ n[54615];
assign t[54616] = t[54615] ^ n[54616];
assign t[54617] = t[54616] ^ n[54617];
assign t[54618] = t[54617] ^ n[54618];
assign t[54619] = t[54618] ^ n[54619];
assign t[54620] = t[54619] ^ n[54620];
assign t[54621] = t[54620] ^ n[54621];
assign t[54622] = t[54621] ^ n[54622];
assign t[54623] = t[54622] ^ n[54623];
assign t[54624] = t[54623] ^ n[54624];
assign t[54625] = t[54624] ^ n[54625];
assign t[54626] = t[54625] ^ n[54626];
assign t[54627] = t[54626] ^ n[54627];
assign t[54628] = t[54627] ^ n[54628];
assign t[54629] = t[54628] ^ n[54629];
assign t[54630] = t[54629] ^ n[54630];
assign t[54631] = t[54630] ^ n[54631];
assign t[54632] = t[54631] ^ n[54632];
assign t[54633] = t[54632] ^ n[54633];
assign t[54634] = t[54633] ^ n[54634];
assign t[54635] = t[54634] ^ n[54635];
assign t[54636] = t[54635] ^ n[54636];
assign t[54637] = t[54636] ^ n[54637];
assign t[54638] = t[54637] ^ n[54638];
assign t[54639] = t[54638] ^ n[54639];
assign t[54640] = t[54639] ^ n[54640];
assign t[54641] = t[54640] ^ n[54641];
assign t[54642] = t[54641] ^ n[54642];
assign t[54643] = t[54642] ^ n[54643];
assign t[54644] = t[54643] ^ n[54644];
assign t[54645] = t[54644] ^ n[54645];
assign t[54646] = t[54645] ^ n[54646];
assign t[54647] = t[54646] ^ n[54647];
assign t[54648] = t[54647] ^ n[54648];
assign t[54649] = t[54648] ^ n[54649];
assign t[54650] = t[54649] ^ n[54650];
assign t[54651] = t[54650] ^ n[54651];
assign t[54652] = t[54651] ^ n[54652];
assign t[54653] = t[54652] ^ n[54653];
assign t[54654] = t[54653] ^ n[54654];
assign t[54655] = t[54654] ^ n[54655];
assign t[54656] = t[54655] ^ n[54656];
assign t[54657] = t[54656] ^ n[54657];
assign t[54658] = t[54657] ^ n[54658];
assign t[54659] = t[54658] ^ n[54659];
assign t[54660] = t[54659] ^ n[54660];
assign t[54661] = t[54660] ^ n[54661];
assign t[54662] = t[54661] ^ n[54662];
assign t[54663] = t[54662] ^ n[54663];
assign t[54664] = t[54663] ^ n[54664];
assign t[54665] = t[54664] ^ n[54665];
assign t[54666] = t[54665] ^ n[54666];
assign t[54667] = t[54666] ^ n[54667];
assign t[54668] = t[54667] ^ n[54668];
assign t[54669] = t[54668] ^ n[54669];
assign t[54670] = t[54669] ^ n[54670];
assign t[54671] = t[54670] ^ n[54671];
assign t[54672] = t[54671] ^ n[54672];
assign t[54673] = t[54672] ^ n[54673];
assign t[54674] = t[54673] ^ n[54674];
assign t[54675] = t[54674] ^ n[54675];
assign t[54676] = t[54675] ^ n[54676];
assign t[54677] = t[54676] ^ n[54677];
assign t[54678] = t[54677] ^ n[54678];
assign t[54679] = t[54678] ^ n[54679];
assign t[54680] = t[54679] ^ n[54680];
assign t[54681] = t[54680] ^ n[54681];
assign t[54682] = t[54681] ^ n[54682];
assign t[54683] = t[54682] ^ n[54683];
assign t[54684] = t[54683] ^ n[54684];
assign t[54685] = t[54684] ^ n[54685];
assign t[54686] = t[54685] ^ n[54686];
assign t[54687] = t[54686] ^ n[54687];
assign t[54688] = t[54687] ^ n[54688];
assign t[54689] = t[54688] ^ n[54689];
assign t[54690] = t[54689] ^ n[54690];
assign t[54691] = t[54690] ^ n[54691];
assign t[54692] = t[54691] ^ n[54692];
assign t[54693] = t[54692] ^ n[54693];
assign t[54694] = t[54693] ^ n[54694];
assign t[54695] = t[54694] ^ n[54695];
assign t[54696] = t[54695] ^ n[54696];
assign t[54697] = t[54696] ^ n[54697];
assign t[54698] = t[54697] ^ n[54698];
assign t[54699] = t[54698] ^ n[54699];
assign t[54700] = t[54699] ^ n[54700];
assign t[54701] = t[54700] ^ n[54701];
assign t[54702] = t[54701] ^ n[54702];
assign t[54703] = t[54702] ^ n[54703];
assign t[54704] = t[54703] ^ n[54704];
assign t[54705] = t[54704] ^ n[54705];
assign t[54706] = t[54705] ^ n[54706];
assign t[54707] = t[54706] ^ n[54707];
assign t[54708] = t[54707] ^ n[54708];
assign t[54709] = t[54708] ^ n[54709];
assign t[54710] = t[54709] ^ n[54710];
assign t[54711] = t[54710] ^ n[54711];
assign t[54712] = t[54711] ^ n[54712];
assign t[54713] = t[54712] ^ n[54713];
assign t[54714] = t[54713] ^ n[54714];
assign t[54715] = t[54714] ^ n[54715];
assign t[54716] = t[54715] ^ n[54716];
assign t[54717] = t[54716] ^ n[54717];
assign t[54718] = t[54717] ^ n[54718];
assign t[54719] = t[54718] ^ n[54719];
assign t[54720] = t[54719] ^ n[54720];
assign t[54721] = t[54720] ^ n[54721];
assign t[54722] = t[54721] ^ n[54722];
assign t[54723] = t[54722] ^ n[54723];
assign t[54724] = t[54723] ^ n[54724];
assign t[54725] = t[54724] ^ n[54725];
assign t[54726] = t[54725] ^ n[54726];
assign t[54727] = t[54726] ^ n[54727];
assign t[54728] = t[54727] ^ n[54728];
assign t[54729] = t[54728] ^ n[54729];
assign t[54730] = t[54729] ^ n[54730];
assign t[54731] = t[54730] ^ n[54731];
assign t[54732] = t[54731] ^ n[54732];
assign t[54733] = t[54732] ^ n[54733];
assign t[54734] = t[54733] ^ n[54734];
assign t[54735] = t[54734] ^ n[54735];
assign t[54736] = t[54735] ^ n[54736];
assign t[54737] = t[54736] ^ n[54737];
assign t[54738] = t[54737] ^ n[54738];
assign t[54739] = t[54738] ^ n[54739];
assign t[54740] = t[54739] ^ n[54740];
assign t[54741] = t[54740] ^ n[54741];
assign t[54742] = t[54741] ^ n[54742];
assign t[54743] = t[54742] ^ n[54743];
assign t[54744] = t[54743] ^ n[54744];
assign t[54745] = t[54744] ^ n[54745];
assign t[54746] = t[54745] ^ n[54746];
assign t[54747] = t[54746] ^ n[54747];
assign t[54748] = t[54747] ^ n[54748];
assign t[54749] = t[54748] ^ n[54749];
assign t[54750] = t[54749] ^ n[54750];
assign t[54751] = t[54750] ^ n[54751];
assign t[54752] = t[54751] ^ n[54752];
assign t[54753] = t[54752] ^ n[54753];
assign t[54754] = t[54753] ^ n[54754];
assign t[54755] = t[54754] ^ n[54755];
assign t[54756] = t[54755] ^ n[54756];
assign t[54757] = t[54756] ^ n[54757];
assign t[54758] = t[54757] ^ n[54758];
assign t[54759] = t[54758] ^ n[54759];
assign t[54760] = t[54759] ^ n[54760];
assign t[54761] = t[54760] ^ n[54761];
assign t[54762] = t[54761] ^ n[54762];
assign t[54763] = t[54762] ^ n[54763];
assign t[54764] = t[54763] ^ n[54764];
assign t[54765] = t[54764] ^ n[54765];
assign t[54766] = t[54765] ^ n[54766];
assign t[54767] = t[54766] ^ n[54767];
assign t[54768] = t[54767] ^ n[54768];
assign t[54769] = t[54768] ^ n[54769];
assign t[54770] = t[54769] ^ n[54770];
assign t[54771] = t[54770] ^ n[54771];
assign t[54772] = t[54771] ^ n[54772];
assign t[54773] = t[54772] ^ n[54773];
assign t[54774] = t[54773] ^ n[54774];
assign t[54775] = t[54774] ^ n[54775];
assign t[54776] = t[54775] ^ n[54776];
assign t[54777] = t[54776] ^ n[54777];
assign t[54778] = t[54777] ^ n[54778];
assign t[54779] = t[54778] ^ n[54779];
assign t[54780] = t[54779] ^ n[54780];
assign t[54781] = t[54780] ^ n[54781];
assign t[54782] = t[54781] ^ n[54782];
assign t[54783] = t[54782] ^ n[54783];
assign t[54784] = t[54783] ^ n[54784];
assign t[54785] = t[54784] ^ n[54785];
assign t[54786] = t[54785] ^ n[54786];
assign t[54787] = t[54786] ^ n[54787];
assign t[54788] = t[54787] ^ n[54788];
assign t[54789] = t[54788] ^ n[54789];
assign t[54790] = t[54789] ^ n[54790];
assign t[54791] = t[54790] ^ n[54791];
assign t[54792] = t[54791] ^ n[54792];
assign t[54793] = t[54792] ^ n[54793];
assign t[54794] = t[54793] ^ n[54794];
assign t[54795] = t[54794] ^ n[54795];
assign t[54796] = t[54795] ^ n[54796];
assign t[54797] = t[54796] ^ n[54797];
assign t[54798] = t[54797] ^ n[54798];
assign t[54799] = t[54798] ^ n[54799];
assign t[54800] = t[54799] ^ n[54800];
assign t[54801] = t[54800] ^ n[54801];
assign t[54802] = t[54801] ^ n[54802];
assign t[54803] = t[54802] ^ n[54803];
assign t[54804] = t[54803] ^ n[54804];
assign t[54805] = t[54804] ^ n[54805];
assign t[54806] = t[54805] ^ n[54806];
assign t[54807] = t[54806] ^ n[54807];
assign t[54808] = t[54807] ^ n[54808];
assign t[54809] = t[54808] ^ n[54809];
assign t[54810] = t[54809] ^ n[54810];
assign t[54811] = t[54810] ^ n[54811];
assign t[54812] = t[54811] ^ n[54812];
assign t[54813] = t[54812] ^ n[54813];
assign t[54814] = t[54813] ^ n[54814];
assign t[54815] = t[54814] ^ n[54815];
assign t[54816] = t[54815] ^ n[54816];
assign t[54817] = t[54816] ^ n[54817];
assign t[54818] = t[54817] ^ n[54818];
assign t[54819] = t[54818] ^ n[54819];
assign t[54820] = t[54819] ^ n[54820];
assign t[54821] = t[54820] ^ n[54821];
assign t[54822] = t[54821] ^ n[54822];
assign t[54823] = t[54822] ^ n[54823];
assign t[54824] = t[54823] ^ n[54824];
assign t[54825] = t[54824] ^ n[54825];
assign t[54826] = t[54825] ^ n[54826];
assign t[54827] = t[54826] ^ n[54827];
assign t[54828] = t[54827] ^ n[54828];
assign t[54829] = t[54828] ^ n[54829];
assign t[54830] = t[54829] ^ n[54830];
assign t[54831] = t[54830] ^ n[54831];
assign t[54832] = t[54831] ^ n[54832];
assign t[54833] = t[54832] ^ n[54833];
assign t[54834] = t[54833] ^ n[54834];
assign t[54835] = t[54834] ^ n[54835];
assign t[54836] = t[54835] ^ n[54836];
assign t[54837] = t[54836] ^ n[54837];
assign t[54838] = t[54837] ^ n[54838];
assign t[54839] = t[54838] ^ n[54839];
assign t[54840] = t[54839] ^ n[54840];
assign t[54841] = t[54840] ^ n[54841];
assign t[54842] = t[54841] ^ n[54842];
assign t[54843] = t[54842] ^ n[54843];
assign t[54844] = t[54843] ^ n[54844];
assign t[54845] = t[54844] ^ n[54845];
assign t[54846] = t[54845] ^ n[54846];
assign t[54847] = t[54846] ^ n[54847];
assign t[54848] = t[54847] ^ n[54848];
assign t[54849] = t[54848] ^ n[54849];
assign t[54850] = t[54849] ^ n[54850];
assign t[54851] = t[54850] ^ n[54851];
assign t[54852] = t[54851] ^ n[54852];
assign t[54853] = t[54852] ^ n[54853];
assign t[54854] = t[54853] ^ n[54854];
assign t[54855] = t[54854] ^ n[54855];
assign t[54856] = t[54855] ^ n[54856];
assign t[54857] = t[54856] ^ n[54857];
assign t[54858] = t[54857] ^ n[54858];
assign t[54859] = t[54858] ^ n[54859];
assign t[54860] = t[54859] ^ n[54860];
assign t[54861] = t[54860] ^ n[54861];
assign t[54862] = t[54861] ^ n[54862];
assign t[54863] = t[54862] ^ n[54863];
assign t[54864] = t[54863] ^ n[54864];
assign t[54865] = t[54864] ^ n[54865];
assign t[54866] = t[54865] ^ n[54866];
assign t[54867] = t[54866] ^ n[54867];
assign t[54868] = t[54867] ^ n[54868];
assign t[54869] = t[54868] ^ n[54869];
assign t[54870] = t[54869] ^ n[54870];
assign t[54871] = t[54870] ^ n[54871];
assign t[54872] = t[54871] ^ n[54872];
assign t[54873] = t[54872] ^ n[54873];
assign t[54874] = t[54873] ^ n[54874];
assign t[54875] = t[54874] ^ n[54875];
assign t[54876] = t[54875] ^ n[54876];
assign t[54877] = t[54876] ^ n[54877];
assign t[54878] = t[54877] ^ n[54878];
assign t[54879] = t[54878] ^ n[54879];
assign t[54880] = t[54879] ^ n[54880];
assign t[54881] = t[54880] ^ n[54881];
assign t[54882] = t[54881] ^ n[54882];
assign t[54883] = t[54882] ^ n[54883];
assign t[54884] = t[54883] ^ n[54884];
assign t[54885] = t[54884] ^ n[54885];
assign t[54886] = t[54885] ^ n[54886];
assign t[54887] = t[54886] ^ n[54887];
assign t[54888] = t[54887] ^ n[54888];
assign t[54889] = t[54888] ^ n[54889];
assign t[54890] = t[54889] ^ n[54890];
assign t[54891] = t[54890] ^ n[54891];
assign t[54892] = t[54891] ^ n[54892];
assign t[54893] = t[54892] ^ n[54893];
assign t[54894] = t[54893] ^ n[54894];
assign t[54895] = t[54894] ^ n[54895];
assign t[54896] = t[54895] ^ n[54896];
assign t[54897] = t[54896] ^ n[54897];
assign t[54898] = t[54897] ^ n[54898];
assign t[54899] = t[54898] ^ n[54899];
assign t[54900] = t[54899] ^ n[54900];
assign t[54901] = t[54900] ^ n[54901];
assign t[54902] = t[54901] ^ n[54902];
assign t[54903] = t[54902] ^ n[54903];
assign t[54904] = t[54903] ^ n[54904];
assign t[54905] = t[54904] ^ n[54905];
assign t[54906] = t[54905] ^ n[54906];
assign t[54907] = t[54906] ^ n[54907];
assign t[54908] = t[54907] ^ n[54908];
assign t[54909] = t[54908] ^ n[54909];
assign t[54910] = t[54909] ^ n[54910];
assign t[54911] = t[54910] ^ n[54911];
assign t[54912] = t[54911] ^ n[54912];
assign t[54913] = t[54912] ^ n[54913];
assign t[54914] = t[54913] ^ n[54914];
assign t[54915] = t[54914] ^ n[54915];
assign t[54916] = t[54915] ^ n[54916];
assign t[54917] = t[54916] ^ n[54917];
assign t[54918] = t[54917] ^ n[54918];
assign t[54919] = t[54918] ^ n[54919];
assign t[54920] = t[54919] ^ n[54920];
assign t[54921] = t[54920] ^ n[54921];
assign t[54922] = t[54921] ^ n[54922];
assign t[54923] = t[54922] ^ n[54923];
assign t[54924] = t[54923] ^ n[54924];
assign t[54925] = t[54924] ^ n[54925];
assign t[54926] = t[54925] ^ n[54926];
assign t[54927] = t[54926] ^ n[54927];
assign t[54928] = t[54927] ^ n[54928];
assign t[54929] = t[54928] ^ n[54929];
assign t[54930] = t[54929] ^ n[54930];
assign t[54931] = t[54930] ^ n[54931];
assign t[54932] = t[54931] ^ n[54932];
assign t[54933] = t[54932] ^ n[54933];
assign t[54934] = t[54933] ^ n[54934];
assign t[54935] = t[54934] ^ n[54935];
assign t[54936] = t[54935] ^ n[54936];
assign t[54937] = t[54936] ^ n[54937];
assign t[54938] = t[54937] ^ n[54938];
assign t[54939] = t[54938] ^ n[54939];
assign t[54940] = t[54939] ^ n[54940];
assign t[54941] = t[54940] ^ n[54941];
assign t[54942] = t[54941] ^ n[54942];
assign t[54943] = t[54942] ^ n[54943];
assign t[54944] = t[54943] ^ n[54944];
assign t[54945] = t[54944] ^ n[54945];
assign t[54946] = t[54945] ^ n[54946];
assign t[54947] = t[54946] ^ n[54947];
assign t[54948] = t[54947] ^ n[54948];
assign t[54949] = t[54948] ^ n[54949];
assign t[54950] = t[54949] ^ n[54950];
assign t[54951] = t[54950] ^ n[54951];
assign t[54952] = t[54951] ^ n[54952];
assign t[54953] = t[54952] ^ n[54953];
assign t[54954] = t[54953] ^ n[54954];
assign t[54955] = t[54954] ^ n[54955];
assign t[54956] = t[54955] ^ n[54956];
assign t[54957] = t[54956] ^ n[54957];
assign t[54958] = t[54957] ^ n[54958];
assign t[54959] = t[54958] ^ n[54959];
assign t[54960] = t[54959] ^ n[54960];
assign t[54961] = t[54960] ^ n[54961];
assign t[54962] = t[54961] ^ n[54962];
assign t[54963] = t[54962] ^ n[54963];
assign t[54964] = t[54963] ^ n[54964];
assign t[54965] = t[54964] ^ n[54965];
assign t[54966] = t[54965] ^ n[54966];
assign t[54967] = t[54966] ^ n[54967];
assign t[54968] = t[54967] ^ n[54968];
assign t[54969] = t[54968] ^ n[54969];
assign t[54970] = t[54969] ^ n[54970];
assign t[54971] = t[54970] ^ n[54971];
assign t[54972] = t[54971] ^ n[54972];
assign t[54973] = t[54972] ^ n[54973];
assign t[54974] = t[54973] ^ n[54974];
assign t[54975] = t[54974] ^ n[54975];
assign t[54976] = t[54975] ^ n[54976];
assign t[54977] = t[54976] ^ n[54977];
assign t[54978] = t[54977] ^ n[54978];
assign t[54979] = t[54978] ^ n[54979];
assign t[54980] = t[54979] ^ n[54980];
assign t[54981] = t[54980] ^ n[54981];
assign t[54982] = t[54981] ^ n[54982];
assign t[54983] = t[54982] ^ n[54983];
assign t[54984] = t[54983] ^ n[54984];
assign t[54985] = t[54984] ^ n[54985];
assign t[54986] = t[54985] ^ n[54986];
assign t[54987] = t[54986] ^ n[54987];
assign t[54988] = t[54987] ^ n[54988];
assign t[54989] = t[54988] ^ n[54989];
assign t[54990] = t[54989] ^ n[54990];
assign t[54991] = t[54990] ^ n[54991];
assign t[54992] = t[54991] ^ n[54992];
assign t[54993] = t[54992] ^ n[54993];
assign t[54994] = t[54993] ^ n[54994];
assign t[54995] = t[54994] ^ n[54995];
assign t[54996] = t[54995] ^ n[54996];
assign t[54997] = t[54996] ^ n[54997];
assign t[54998] = t[54997] ^ n[54998];
assign t[54999] = t[54998] ^ n[54999];
assign t[55000] = t[54999] ^ n[55000];
assign t[55001] = t[55000] ^ n[55001];
assign t[55002] = t[55001] ^ n[55002];
assign t[55003] = t[55002] ^ n[55003];
assign t[55004] = t[55003] ^ n[55004];
assign t[55005] = t[55004] ^ n[55005];
assign t[55006] = t[55005] ^ n[55006];
assign t[55007] = t[55006] ^ n[55007];
assign t[55008] = t[55007] ^ n[55008];
assign t[55009] = t[55008] ^ n[55009];
assign t[55010] = t[55009] ^ n[55010];
assign t[55011] = t[55010] ^ n[55011];
assign t[55012] = t[55011] ^ n[55012];
assign t[55013] = t[55012] ^ n[55013];
assign t[55014] = t[55013] ^ n[55014];
assign t[55015] = t[55014] ^ n[55015];
assign t[55016] = t[55015] ^ n[55016];
assign t[55017] = t[55016] ^ n[55017];
assign t[55018] = t[55017] ^ n[55018];
assign t[55019] = t[55018] ^ n[55019];
assign t[55020] = t[55019] ^ n[55020];
assign t[55021] = t[55020] ^ n[55021];
assign t[55022] = t[55021] ^ n[55022];
assign t[55023] = t[55022] ^ n[55023];
assign t[55024] = t[55023] ^ n[55024];
assign t[55025] = t[55024] ^ n[55025];
assign t[55026] = t[55025] ^ n[55026];
assign t[55027] = t[55026] ^ n[55027];
assign t[55028] = t[55027] ^ n[55028];
assign t[55029] = t[55028] ^ n[55029];
assign t[55030] = t[55029] ^ n[55030];
assign t[55031] = t[55030] ^ n[55031];
assign t[55032] = t[55031] ^ n[55032];
assign t[55033] = t[55032] ^ n[55033];
assign t[55034] = t[55033] ^ n[55034];
assign t[55035] = t[55034] ^ n[55035];
assign t[55036] = t[55035] ^ n[55036];
assign t[55037] = t[55036] ^ n[55037];
assign t[55038] = t[55037] ^ n[55038];
assign t[55039] = t[55038] ^ n[55039];
assign t[55040] = t[55039] ^ n[55040];
assign t[55041] = t[55040] ^ n[55041];
assign t[55042] = t[55041] ^ n[55042];
assign t[55043] = t[55042] ^ n[55043];
assign t[55044] = t[55043] ^ n[55044];
assign t[55045] = t[55044] ^ n[55045];
assign t[55046] = t[55045] ^ n[55046];
assign t[55047] = t[55046] ^ n[55047];
assign t[55048] = t[55047] ^ n[55048];
assign t[55049] = t[55048] ^ n[55049];
assign t[55050] = t[55049] ^ n[55050];
assign t[55051] = t[55050] ^ n[55051];
assign t[55052] = t[55051] ^ n[55052];
assign t[55053] = t[55052] ^ n[55053];
assign t[55054] = t[55053] ^ n[55054];
assign t[55055] = t[55054] ^ n[55055];
assign t[55056] = t[55055] ^ n[55056];
assign t[55057] = t[55056] ^ n[55057];
assign t[55058] = t[55057] ^ n[55058];
assign t[55059] = t[55058] ^ n[55059];
assign t[55060] = t[55059] ^ n[55060];
assign t[55061] = t[55060] ^ n[55061];
assign t[55062] = t[55061] ^ n[55062];
assign t[55063] = t[55062] ^ n[55063];
assign t[55064] = t[55063] ^ n[55064];
assign t[55065] = t[55064] ^ n[55065];
assign t[55066] = t[55065] ^ n[55066];
assign t[55067] = t[55066] ^ n[55067];
assign t[55068] = t[55067] ^ n[55068];
assign t[55069] = t[55068] ^ n[55069];
assign t[55070] = t[55069] ^ n[55070];
assign t[55071] = t[55070] ^ n[55071];
assign t[55072] = t[55071] ^ n[55072];
assign t[55073] = t[55072] ^ n[55073];
assign t[55074] = t[55073] ^ n[55074];
assign t[55075] = t[55074] ^ n[55075];
assign t[55076] = t[55075] ^ n[55076];
assign t[55077] = t[55076] ^ n[55077];
assign t[55078] = t[55077] ^ n[55078];
assign t[55079] = t[55078] ^ n[55079];
assign t[55080] = t[55079] ^ n[55080];
assign t[55081] = t[55080] ^ n[55081];
assign t[55082] = t[55081] ^ n[55082];
assign t[55083] = t[55082] ^ n[55083];
assign t[55084] = t[55083] ^ n[55084];
assign t[55085] = t[55084] ^ n[55085];
assign t[55086] = t[55085] ^ n[55086];
assign t[55087] = t[55086] ^ n[55087];
assign t[55088] = t[55087] ^ n[55088];
assign t[55089] = t[55088] ^ n[55089];
assign t[55090] = t[55089] ^ n[55090];
assign t[55091] = t[55090] ^ n[55091];
assign t[55092] = t[55091] ^ n[55092];
assign t[55093] = t[55092] ^ n[55093];
assign t[55094] = t[55093] ^ n[55094];
assign t[55095] = t[55094] ^ n[55095];
assign t[55096] = t[55095] ^ n[55096];
assign t[55097] = t[55096] ^ n[55097];
assign t[55098] = t[55097] ^ n[55098];
assign t[55099] = t[55098] ^ n[55099];
assign t[55100] = t[55099] ^ n[55100];
assign t[55101] = t[55100] ^ n[55101];
assign t[55102] = t[55101] ^ n[55102];
assign t[55103] = t[55102] ^ n[55103];
assign t[55104] = t[55103] ^ n[55104];
assign t[55105] = t[55104] ^ n[55105];
assign t[55106] = t[55105] ^ n[55106];
assign t[55107] = t[55106] ^ n[55107];
assign t[55108] = t[55107] ^ n[55108];
assign t[55109] = t[55108] ^ n[55109];
assign t[55110] = t[55109] ^ n[55110];
assign t[55111] = t[55110] ^ n[55111];
assign t[55112] = t[55111] ^ n[55112];
assign t[55113] = t[55112] ^ n[55113];
assign t[55114] = t[55113] ^ n[55114];
assign t[55115] = t[55114] ^ n[55115];
assign t[55116] = t[55115] ^ n[55116];
assign t[55117] = t[55116] ^ n[55117];
assign t[55118] = t[55117] ^ n[55118];
assign t[55119] = t[55118] ^ n[55119];
assign t[55120] = t[55119] ^ n[55120];
assign t[55121] = t[55120] ^ n[55121];
assign t[55122] = t[55121] ^ n[55122];
assign t[55123] = t[55122] ^ n[55123];
assign t[55124] = t[55123] ^ n[55124];
assign t[55125] = t[55124] ^ n[55125];
assign t[55126] = t[55125] ^ n[55126];
assign t[55127] = t[55126] ^ n[55127];
assign t[55128] = t[55127] ^ n[55128];
assign t[55129] = t[55128] ^ n[55129];
assign t[55130] = t[55129] ^ n[55130];
assign t[55131] = t[55130] ^ n[55131];
assign t[55132] = t[55131] ^ n[55132];
assign t[55133] = t[55132] ^ n[55133];
assign t[55134] = t[55133] ^ n[55134];
assign t[55135] = t[55134] ^ n[55135];
assign t[55136] = t[55135] ^ n[55136];
assign t[55137] = t[55136] ^ n[55137];
assign t[55138] = t[55137] ^ n[55138];
assign t[55139] = t[55138] ^ n[55139];
assign t[55140] = t[55139] ^ n[55140];
assign t[55141] = t[55140] ^ n[55141];
assign t[55142] = t[55141] ^ n[55142];
assign t[55143] = t[55142] ^ n[55143];
assign t[55144] = t[55143] ^ n[55144];
assign t[55145] = t[55144] ^ n[55145];
assign t[55146] = t[55145] ^ n[55146];
assign t[55147] = t[55146] ^ n[55147];
assign t[55148] = t[55147] ^ n[55148];
assign t[55149] = t[55148] ^ n[55149];
assign t[55150] = t[55149] ^ n[55150];
assign t[55151] = t[55150] ^ n[55151];
assign t[55152] = t[55151] ^ n[55152];
assign t[55153] = t[55152] ^ n[55153];
assign t[55154] = t[55153] ^ n[55154];
assign t[55155] = t[55154] ^ n[55155];
assign t[55156] = t[55155] ^ n[55156];
assign t[55157] = t[55156] ^ n[55157];
assign t[55158] = t[55157] ^ n[55158];
assign t[55159] = t[55158] ^ n[55159];
assign t[55160] = t[55159] ^ n[55160];
assign t[55161] = t[55160] ^ n[55161];
assign t[55162] = t[55161] ^ n[55162];
assign t[55163] = t[55162] ^ n[55163];
assign t[55164] = t[55163] ^ n[55164];
assign t[55165] = t[55164] ^ n[55165];
assign t[55166] = t[55165] ^ n[55166];
assign t[55167] = t[55166] ^ n[55167];
assign t[55168] = t[55167] ^ n[55168];
assign t[55169] = t[55168] ^ n[55169];
assign t[55170] = t[55169] ^ n[55170];
assign t[55171] = t[55170] ^ n[55171];
assign t[55172] = t[55171] ^ n[55172];
assign t[55173] = t[55172] ^ n[55173];
assign t[55174] = t[55173] ^ n[55174];
assign t[55175] = t[55174] ^ n[55175];
assign t[55176] = t[55175] ^ n[55176];
assign t[55177] = t[55176] ^ n[55177];
assign t[55178] = t[55177] ^ n[55178];
assign t[55179] = t[55178] ^ n[55179];
assign t[55180] = t[55179] ^ n[55180];
assign t[55181] = t[55180] ^ n[55181];
assign t[55182] = t[55181] ^ n[55182];
assign t[55183] = t[55182] ^ n[55183];
assign t[55184] = t[55183] ^ n[55184];
assign t[55185] = t[55184] ^ n[55185];
assign t[55186] = t[55185] ^ n[55186];
assign t[55187] = t[55186] ^ n[55187];
assign t[55188] = t[55187] ^ n[55188];
assign t[55189] = t[55188] ^ n[55189];
assign t[55190] = t[55189] ^ n[55190];
assign t[55191] = t[55190] ^ n[55191];
assign t[55192] = t[55191] ^ n[55192];
assign t[55193] = t[55192] ^ n[55193];
assign t[55194] = t[55193] ^ n[55194];
assign t[55195] = t[55194] ^ n[55195];
assign t[55196] = t[55195] ^ n[55196];
assign t[55197] = t[55196] ^ n[55197];
assign t[55198] = t[55197] ^ n[55198];
assign t[55199] = t[55198] ^ n[55199];
assign t[55200] = t[55199] ^ n[55200];
assign t[55201] = t[55200] ^ n[55201];
assign t[55202] = t[55201] ^ n[55202];
assign t[55203] = t[55202] ^ n[55203];
assign t[55204] = t[55203] ^ n[55204];
assign t[55205] = t[55204] ^ n[55205];
assign t[55206] = t[55205] ^ n[55206];
assign t[55207] = t[55206] ^ n[55207];
assign t[55208] = t[55207] ^ n[55208];
assign t[55209] = t[55208] ^ n[55209];
assign t[55210] = t[55209] ^ n[55210];
assign t[55211] = t[55210] ^ n[55211];
assign t[55212] = t[55211] ^ n[55212];
assign t[55213] = t[55212] ^ n[55213];
assign t[55214] = t[55213] ^ n[55214];
assign t[55215] = t[55214] ^ n[55215];
assign t[55216] = t[55215] ^ n[55216];
assign t[55217] = t[55216] ^ n[55217];
assign t[55218] = t[55217] ^ n[55218];
assign t[55219] = t[55218] ^ n[55219];
assign t[55220] = t[55219] ^ n[55220];
assign t[55221] = t[55220] ^ n[55221];
assign t[55222] = t[55221] ^ n[55222];
assign t[55223] = t[55222] ^ n[55223];
assign t[55224] = t[55223] ^ n[55224];
assign t[55225] = t[55224] ^ n[55225];
assign t[55226] = t[55225] ^ n[55226];
assign t[55227] = t[55226] ^ n[55227];
assign t[55228] = t[55227] ^ n[55228];
assign t[55229] = t[55228] ^ n[55229];
assign t[55230] = t[55229] ^ n[55230];
assign t[55231] = t[55230] ^ n[55231];
assign t[55232] = t[55231] ^ n[55232];
assign t[55233] = t[55232] ^ n[55233];
assign t[55234] = t[55233] ^ n[55234];
assign t[55235] = t[55234] ^ n[55235];
assign t[55236] = t[55235] ^ n[55236];
assign t[55237] = t[55236] ^ n[55237];
assign t[55238] = t[55237] ^ n[55238];
assign t[55239] = t[55238] ^ n[55239];
assign t[55240] = t[55239] ^ n[55240];
assign t[55241] = t[55240] ^ n[55241];
assign t[55242] = t[55241] ^ n[55242];
assign t[55243] = t[55242] ^ n[55243];
assign t[55244] = t[55243] ^ n[55244];
assign t[55245] = t[55244] ^ n[55245];
assign t[55246] = t[55245] ^ n[55246];
assign t[55247] = t[55246] ^ n[55247];
assign t[55248] = t[55247] ^ n[55248];
assign t[55249] = t[55248] ^ n[55249];
assign t[55250] = t[55249] ^ n[55250];
assign t[55251] = t[55250] ^ n[55251];
assign t[55252] = t[55251] ^ n[55252];
assign t[55253] = t[55252] ^ n[55253];
assign t[55254] = t[55253] ^ n[55254];
assign t[55255] = t[55254] ^ n[55255];
assign t[55256] = t[55255] ^ n[55256];
assign t[55257] = t[55256] ^ n[55257];
assign t[55258] = t[55257] ^ n[55258];
assign t[55259] = t[55258] ^ n[55259];
assign t[55260] = t[55259] ^ n[55260];
assign t[55261] = t[55260] ^ n[55261];
assign t[55262] = t[55261] ^ n[55262];
assign t[55263] = t[55262] ^ n[55263];
assign t[55264] = t[55263] ^ n[55264];
assign t[55265] = t[55264] ^ n[55265];
assign t[55266] = t[55265] ^ n[55266];
assign t[55267] = t[55266] ^ n[55267];
assign t[55268] = t[55267] ^ n[55268];
assign t[55269] = t[55268] ^ n[55269];
assign t[55270] = t[55269] ^ n[55270];
assign t[55271] = t[55270] ^ n[55271];
assign t[55272] = t[55271] ^ n[55272];
assign t[55273] = t[55272] ^ n[55273];
assign t[55274] = t[55273] ^ n[55274];
assign t[55275] = t[55274] ^ n[55275];
assign t[55276] = t[55275] ^ n[55276];
assign t[55277] = t[55276] ^ n[55277];
assign t[55278] = t[55277] ^ n[55278];
assign t[55279] = t[55278] ^ n[55279];
assign t[55280] = t[55279] ^ n[55280];
assign t[55281] = t[55280] ^ n[55281];
assign t[55282] = t[55281] ^ n[55282];
assign t[55283] = t[55282] ^ n[55283];
assign t[55284] = t[55283] ^ n[55284];
assign t[55285] = t[55284] ^ n[55285];
assign t[55286] = t[55285] ^ n[55286];
assign t[55287] = t[55286] ^ n[55287];
assign t[55288] = t[55287] ^ n[55288];
assign t[55289] = t[55288] ^ n[55289];
assign t[55290] = t[55289] ^ n[55290];
assign t[55291] = t[55290] ^ n[55291];
assign t[55292] = t[55291] ^ n[55292];
assign t[55293] = t[55292] ^ n[55293];
assign t[55294] = t[55293] ^ n[55294];
assign t[55295] = t[55294] ^ n[55295];
assign t[55296] = t[55295] ^ n[55296];
assign t[55297] = t[55296] ^ n[55297];
assign t[55298] = t[55297] ^ n[55298];
assign t[55299] = t[55298] ^ n[55299];
assign t[55300] = t[55299] ^ n[55300];
assign t[55301] = t[55300] ^ n[55301];
assign t[55302] = t[55301] ^ n[55302];
assign t[55303] = t[55302] ^ n[55303];
assign t[55304] = t[55303] ^ n[55304];
assign t[55305] = t[55304] ^ n[55305];
assign t[55306] = t[55305] ^ n[55306];
assign t[55307] = t[55306] ^ n[55307];
assign t[55308] = t[55307] ^ n[55308];
assign t[55309] = t[55308] ^ n[55309];
assign t[55310] = t[55309] ^ n[55310];
assign t[55311] = t[55310] ^ n[55311];
assign t[55312] = t[55311] ^ n[55312];
assign t[55313] = t[55312] ^ n[55313];
assign t[55314] = t[55313] ^ n[55314];
assign t[55315] = t[55314] ^ n[55315];
assign t[55316] = t[55315] ^ n[55316];
assign t[55317] = t[55316] ^ n[55317];
assign t[55318] = t[55317] ^ n[55318];
assign t[55319] = t[55318] ^ n[55319];
assign t[55320] = t[55319] ^ n[55320];
assign t[55321] = t[55320] ^ n[55321];
assign t[55322] = t[55321] ^ n[55322];
assign t[55323] = t[55322] ^ n[55323];
assign t[55324] = t[55323] ^ n[55324];
assign t[55325] = t[55324] ^ n[55325];
assign t[55326] = t[55325] ^ n[55326];
assign t[55327] = t[55326] ^ n[55327];
assign t[55328] = t[55327] ^ n[55328];
assign t[55329] = t[55328] ^ n[55329];
assign t[55330] = t[55329] ^ n[55330];
assign t[55331] = t[55330] ^ n[55331];
assign t[55332] = t[55331] ^ n[55332];
assign t[55333] = t[55332] ^ n[55333];
assign t[55334] = t[55333] ^ n[55334];
assign t[55335] = t[55334] ^ n[55335];
assign t[55336] = t[55335] ^ n[55336];
assign t[55337] = t[55336] ^ n[55337];
assign t[55338] = t[55337] ^ n[55338];
assign t[55339] = t[55338] ^ n[55339];
assign t[55340] = t[55339] ^ n[55340];
assign t[55341] = t[55340] ^ n[55341];
assign t[55342] = t[55341] ^ n[55342];
assign t[55343] = t[55342] ^ n[55343];
assign t[55344] = t[55343] ^ n[55344];
assign t[55345] = t[55344] ^ n[55345];
assign t[55346] = t[55345] ^ n[55346];
assign t[55347] = t[55346] ^ n[55347];
assign t[55348] = t[55347] ^ n[55348];
assign t[55349] = t[55348] ^ n[55349];
assign t[55350] = t[55349] ^ n[55350];
assign t[55351] = t[55350] ^ n[55351];
assign t[55352] = t[55351] ^ n[55352];
assign t[55353] = t[55352] ^ n[55353];
assign t[55354] = t[55353] ^ n[55354];
assign t[55355] = t[55354] ^ n[55355];
assign t[55356] = t[55355] ^ n[55356];
assign t[55357] = t[55356] ^ n[55357];
assign t[55358] = t[55357] ^ n[55358];
assign t[55359] = t[55358] ^ n[55359];
assign t[55360] = t[55359] ^ n[55360];
assign t[55361] = t[55360] ^ n[55361];
assign t[55362] = t[55361] ^ n[55362];
assign t[55363] = t[55362] ^ n[55363];
assign t[55364] = t[55363] ^ n[55364];
assign t[55365] = t[55364] ^ n[55365];
assign t[55366] = t[55365] ^ n[55366];
assign t[55367] = t[55366] ^ n[55367];
assign t[55368] = t[55367] ^ n[55368];
assign t[55369] = t[55368] ^ n[55369];
assign t[55370] = t[55369] ^ n[55370];
assign t[55371] = t[55370] ^ n[55371];
assign t[55372] = t[55371] ^ n[55372];
assign t[55373] = t[55372] ^ n[55373];
assign t[55374] = t[55373] ^ n[55374];
assign t[55375] = t[55374] ^ n[55375];
assign t[55376] = t[55375] ^ n[55376];
assign t[55377] = t[55376] ^ n[55377];
assign t[55378] = t[55377] ^ n[55378];
assign t[55379] = t[55378] ^ n[55379];
assign t[55380] = t[55379] ^ n[55380];
assign t[55381] = t[55380] ^ n[55381];
assign t[55382] = t[55381] ^ n[55382];
assign t[55383] = t[55382] ^ n[55383];
assign t[55384] = t[55383] ^ n[55384];
assign t[55385] = t[55384] ^ n[55385];
assign t[55386] = t[55385] ^ n[55386];
assign t[55387] = t[55386] ^ n[55387];
assign t[55388] = t[55387] ^ n[55388];
assign t[55389] = t[55388] ^ n[55389];
assign t[55390] = t[55389] ^ n[55390];
assign t[55391] = t[55390] ^ n[55391];
assign t[55392] = t[55391] ^ n[55392];
assign t[55393] = t[55392] ^ n[55393];
assign t[55394] = t[55393] ^ n[55394];
assign t[55395] = t[55394] ^ n[55395];
assign t[55396] = t[55395] ^ n[55396];
assign t[55397] = t[55396] ^ n[55397];
assign t[55398] = t[55397] ^ n[55398];
assign t[55399] = t[55398] ^ n[55399];
assign t[55400] = t[55399] ^ n[55400];
assign t[55401] = t[55400] ^ n[55401];
assign t[55402] = t[55401] ^ n[55402];
assign t[55403] = t[55402] ^ n[55403];
assign t[55404] = t[55403] ^ n[55404];
assign t[55405] = t[55404] ^ n[55405];
assign t[55406] = t[55405] ^ n[55406];
assign t[55407] = t[55406] ^ n[55407];
assign t[55408] = t[55407] ^ n[55408];
assign t[55409] = t[55408] ^ n[55409];
assign t[55410] = t[55409] ^ n[55410];
assign t[55411] = t[55410] ^ n[55411];
assign t[55412] = t[55411] ^ n[55412];
assign t[55413] = t[55412] ^ n[55413];
assign t[55414] = t[55413] ^ n[55414];
assign t[55415] = t[55414] ^ n[55415];
assign t[55416] = t[55415] ^ n[55416];
assign t[55417] = t[55416] ^ n[55417];
assign t[55418] = t[55417] ^ n[55418];
assign t[55419] = t[55418] ^ n[55419];
assign t[55420] = t[55419] ^ n[55420];
assign t[55421] = t[55420] ^ n[55421];
assign t[55422] = t[55421] ^ n[55422];
assign t[55423] = t[55422] ^ n[55423];
assign t[55424] = t[55423] ^ n[55424];
assign t[55425] = t[55424] ^ n[55425];
assign t[55426] = t[55425] ^ n[55426];
assign t[55427] = t[55426] ^ n[55427];
assign t[55428] = t[55427] ^ n[55428];
assign t[55429] = t[55428] ^ n[55429];
assign t[55430] = t[55429] ^ n[55430];
assign t[55431] = t[55430] ^ n[55431];
assign t[55432] = t[55431] ^ n[55432];
assign t[55433] = t[55432] ^ n[55433];
assign t[55434] = t[55433] ^ n[55434];
assign t[55435] = t[55434] ^ n[55435];
assign t[55436] = t[55435] ^ n[55436];
assign t[55437] = t[55436] ^ n[55437];
assign t[55438] = t[55437] ^ n[55438];
assign t[55439] = t[55438] ^ n[55439];
assign t[55440] = t[55439] ^ n[55440];
assign t[55441] = t[55440] ^ n[55441];
assign t[55442] = t[55441] ^ n[55442];
assign t[55443] = t[55442] ^ n[55443];
assign t[55444] = t[55443] ^ n[55444];
assign t[55445] = t[55444] ^ n[55445];
assign t[55446] = t[55445] ^ n[55446];
assign t[55447] = t[55446] ^ n[55447];
assign t[55448] = t[55447] ^ n[55448];
assign t[55449] = t[55448] ^ n[55449];
assign t[55450] = t[55449] ^ n[55450];
assign t[55451] = t[55450] ^ n[55451];
assign t[55452] = t[55451] ^ n[55452];
assign t[55453] = t[55452] ^ n[55453];
assign t[55454] = t[55453] ^ n[55454];
assign t[55455] = t[55454] ^ n[55455];
assign t[55456] = t[55455] ^ n[55456];
assign t[55457] = t[55456] ^ n[55457];
assign t[55458] = t[55457] ^ n[55458];
assign t[55459] = t[55458] ^ n[55459];
assign t[55460] = t[55459] ^ n[55460];
assign t[55461] = t[55460] ^ n[55461];
assign t[55462] = t[55461] ^ n[55462];
assign t[55463] = t[55462] ^ n[55463];
assign t[55464] = t[55463] ^ n[55464];
assign t[55465] = t[55464] ^ n[55465];
assign t[55466] = t[55465] ^ n[55466];
assign t[55467] = t[55466] ^ n[55467];
assign t[55468] = t[55467] ^ n[55468];
assign t[55469] = t[55468] ^ n[55469];
assign t[55470] = t[55469] ^ n[55470];
assign t[55471] = t[55470] ^ n[55471];
assign t[55472] = t[55471] ^ n[55472];
assign t[55473] = t[55472] ^ n[55473];
assign t[55474] = t[55473] ^ n[55474];
assign t[55475] = t[55474] ^ n[55475];
assign t[55476] = t[55475] ^ n[55476];
assign t[55477] = t[55476] ^ n[55477];
assign t[55478] = t[55477] ^ n[55478];
assign t[55479] = t[55478] ^ n[55479];
assign t[55480] = t[55479] ^ n[55480];
assign t[55481] = t[55480] ^ n[55481];
assign t[55482] = t[55481] ^ n[55482];
assign t[55483] = t[55482] ^ n[55483];
assign t[55484] = t[55483] ^ n[55484];
assign t[55485] = t[55484] ^ n[55485];
assign t[55486] = t[55485] ^ n[55486];
assign t[55487] = t[55486] ^ n[55487];
assign t[55488] = t[55487] ^ n[55488];
assign t[55489] = t[55488] ^ n[55489];
assign t[55490] = t[55489] ^ n[55490];
assign t[55491] = t[55490] ^ n[55491];
assign t[55492] = t[55491] ^ n[55492];
assign t[55493] = t[55492] ^ n[55493];
assign t[55494] = t[55493] ^ n[55494];
assign t[55495] = t[55494] ^ n[55495];
assign t[55496] = t[55495] ^ n[55496];
assign t[55497] = t[55496] ^ n[55497];
assign t[55498] = t[55497] ^ n[55498];
assign t[55499] = t[55498] ^ n[55499];
assign t[55500] = t[55499] ^ n[55500];
assign t[55501] = t[55500] ^ n[55501];
assign t[55502] = t[55501] ^ n[55502];
assign t[55503] = t[55502] ^ n[55503];
assign t[55504] = t[55503] ^ n[55504];
assign t[55505] = t[55504] ^ n[55505];
assign t[55506] = t[55505] ^ n[55506];
assign t[55507] = t[55506] ^ n[55507];
assign t[55508] = t[55507] ^ n[55508];
assign t[55509] = t[55508] ^ n[55509];
assign t[55510] = t[55509] ^ n[55510];
assign t[55511] = t[55510] ^ n[55511];
assign t[55512] = t[55511] ^ n[55512];
assign t[55513] = t[55512] ^ n[55513];
assign t[55514] = t[55513] ^ n[55514];
assign t[55515] = t[55514] ^ n[55515];
assign t[55516] = t[55515] ^ n[55516];
assign t[55517] = t[55516] ^ n[55517];
assign t[55518] = t[55517] ^ n[55518];
assign t[55519] = t[55518] ^ n[55519];
assign t[55520] = t[55519] ^ n[55520];
assign t[55521] = t[55520] ^ n[55521];
assign t[55522] = t[55521] ^ n[55522];
assign t[55523] = t[55522] ^ n[55523];
assign t[55524] = t[55523] ^ n[55524];
assign t[55525] = t[55524] ^ n[55525];
assign t[55526] = t[55525] ^ n[55526];
assign t[55527] = t[55526] ^ n[55527];
assign t[55528] = t[55527] ^ n[55528];
assign t[55529] = t[55528] ^ n[55529];
assign t[55530] = t[55529] ^ n[55530];
assign t[55531] = t[55530] ^ n[55531];
assign t[55532] = t[55531] ^ n[55532];
assign t[55533] = t[55532] ^ n[55533];
assign t[55534] = t[55533] ^ n[55534];
assign t[55535] = t[55534] ^ n[55535];
assign t[55536] = t[55535] ^ n[55536];
assign t[55537] = t[55536] ^ n[55537];
assign t[55538] = t[55537] ^ n[55538];
assign t[55539] = t[55538] ^ n[55539];
assign t[55540] = t[55539] ^ n[55540];
assign t[55541] = t[55540] ^ n[55541];
assign t[55542] = t[55541] ^ n[55542];
assign t[55543] = t[55542] ^ n[55543];
assign t[55544] = t[55543] ^ n[55544];
assign t[55545] = t[55544] ^ n[55545];
assign t[55546] = t[55545] ^ n[55546];
assign t[55547] = t[55546] ^ n[55547];
assign t[55548] = t[55547] ^ n[55548];
assign t[55549] = t[55548] ^ n[55549];
assign t[55550] = t[55549] ^ n[55550];
assign t[55551] = t[55550] ^ n[55551];
assign t[55552] = t[55551] ^ n[55552];
assign t[55553] = t[55552] ^ n[55553];
assign t[55554] = t[55553] ^ n[55554];
assign t[55555] = t[55554] ^ n[55555];
assign t[55556] = t[55555] ^ n[55556];
assign t[55557] = t[55556] ^ n[55557];
assign t[55558] = t[55557] ^ n[55558];
assign t[55559] = t[55558] ^ n[55559];
assign t[55560] = t[55559] ^ n[55560];
assign t[55561] = t[55560] ^ n[55561];
assign t[55562] = t[55561] ^ n[55562];
assign t[55563] = t[55562] ^ n[55563];
assign t[55564] = t[55563] ^ n[55564];
assign t[55565] = t[55564] ^ n[55565];
assign t[55566] = t[55565] ^ n[55566];
assign t[55567] = t[55566] ^ n[55567];
assign t[55568] = t[55567] ^ n[55568];
assign t[55569] = t[55568] ^ n[55569];
assign t[55570] = t[55569] ^ n[55570];
assign t[55571] = t[55570] ^ n[55571];
assign t[55572] = t[55571] ^ n[55572];
assign t[55573] = t[55572] ^ n[55573];
assign t[55574] = t[55573] ^ n[55574];
assign t[55575] = t[55574] ^ n[55575];
assign t[55576] = t[55575] ^ n[55576];
assign t[55577] = t[55576] ^ n[55577];
assign t[55578] = t[55577] ^ n[55578];
assign t[55579] = t[55578] ^ n[55579];
assign t[55580] = t[55579] ^ n[55580];
assign t[55581] = t[55580] ^ n[55581];
assign t[55582] = t[55581] ^ n[55582];
assign t[55583] = t[55582] ^ n[55583];
assign t[55584] = t[55583] ^ n[55584];
assign t[55585] = t[55584] ^ n[55585];
assign t[55586] = t[55585] ^ n[55586];
assign t[55587] = t[55586] ^ n[55587];
assign t[55588] = t[55587] ^ n[55588];
assign t[55589] = t[55588] ^ n[55589];
assign t[55590] = t[55589] ^ n[55590];
assign t[55591] = t[55590] ^ n[55591];
assign t[55592] = t[55591] ^ n[55592];
assign t[55593] = t[55592] ^ n[55593];
assign t[55594] = t[55593] ^ n[55594];
assign t[55595] = t[55594] ^ n[55595];
assign t[55596] = t[55595] ^ n[55596];
assign t[55597] = t[55596] ^ n[55597];
assign t[55598] = t[55597] ^ n[55598];
assign t[55599] = t[55598] ^ n[55599];
assign t[55600] = t[55599] ^ n[55600];
assign t[55601] = t[55600] ^ n[55601];
assign t[55602] = t[55601] ^ n[55602];
assign t[55603] = t[55602] ^ n[55603];
assign t[55604] = t[55603] ^ n[55604];
assign t[55605] = t[55604] ^ n[55605];
assign t[55606] = t[55605] ^ n[55606];
assign t[55607] = t[55606] ^ n[55607];
assign t[55608] = t[55607] ^ n[55608];
assign t[55609] = t[55608] ^ n[55609];
assign t[55610] = t[55609] ^ n[55610];
assign t[55611] = t[55610] ^ n[55611];
assign t[55612] = t[55611] ^ n[55612];
assign t[55613] = t[55612] ^ n[55613];
assign t[55614] = t[55613] ^ n[55614];
assign t[55615] = t[55614] ^ n[55615];
assign t[55616] = t[55615] ^ n[55616];
assign t[55617] = t[55616] ^ n[55617];
assign t[55618] = t[55617] ^ n[55618];
assign t[55619] = t[55618] ^ n[55619];
assign t[55620] = t[55619] ^ n[55620];
assign t[55621] = t[55620] ^ n[55621];
assign t[55622] = t[55621] ^ n[55622];
assign t[55623] = t[55622] ^ n[55623];
assign t[55624] = t[55623] ^ n[55624];
assign t[55625] = t[55624] ^ n[55625];
assign t[55626] = t[55625] ^ n[55626];
assign t[55627] = t[55626] ^ n[55627];
assign t[55628] = t[55627] ^ n[55628];
assign t[55629] = t[55628] ^ n[55629];
assign t[55630] = t[55629] ^ n[55630];
assign t[55631] = t[55630] ^ n[55631];
assign t[55632] = t[55631] ^ n[55632];
assign t[55633] = t[55632] ^ n[55633];
assign t[55634] = t[55633] ^ n[55634];
assign t[55635] = t[55634] ^ n[55635];
assign t[55636] = t[55635] ^ n[55636];
assign t[55637] = t[55636] ^ n[55637];
assign t[55638] = t[55637] ^ n[55638];
assign t[55639] = t[55638] ^ n[55639];
assign t[55640] = t[55639] ^ n[55640];
assign t[55641] = t[55640] ^ n[55641];
assign t[55642] = t[55641] ^ n[55642];
assign t[55643] = t[55642] ^ n[55643];
assign t[55644] = t[55643] ^ n[55644];
assign t[55645] = t[55644] ^ n[55645];
assign t[55646] = t[55645] ^ n[55646];
assign t[55647] = t[55646] ^ n[55647];
assign t[55648] = t[55647] ^ n[55648];
assign t[55649] = t[55648] ^ n[55649];
assign t[55650] = t[55649] ^ n[55650];
assign t[55651] = t[55650] ^ n[55651];
assign t[55652] = t[55651] ^ n[55652];
assign t[55653] = t[55652] ^ n[55653];
assign t[55654] = t[55653] ^ n[55654];
assign t[55655] = t[55654] ^ n[55655];
assign t[55656] = t[55655] ^ n[55656];
assign t[55657] = t[55656] ^ n[55657];
assign t[55658] = t[55657] ^ n[55658];
assign t[55659] = t[55658] ^ n[55659];
assign t[55660] = t[55659] ^ n[55660];
assign t[55661] = t[55660] ^ n[55661];
assign t[55662] = t[55661] ^ n[55662];
assign t[55663] = t[55662] ^ n[55663];
assign t[55664] = t[55663] ^ n[55664];
assign t[55665] = t[55664] ^ n[55665];
assign t[55666] = t[55665] ^ n[55666];
assign t[55667] = t[55666] ^ n[55667];
assign t[55668] = t[55667] ^ n[55668];
assign t[55669] = t[55668] ^ n[55669];
assign t[55670] = t[55669] ^ n[55670];
assign t[55671] = t[55670] ^ n[55671];
assign t[55672] = t[55671] ^ n[55672];
assign t[55673] = t[55672] ^ n[55673];
assign t[55674] = t[55673] ^ n[55674];
assign t[55675] = t[55674] ^ n[55675];
assign t[55676] = t[55675] ^ n[55676];
assign t[55677] = t[55676] ^ n[55677];
assign t[55678] = t[55677] ^ n[55678];
assign t[55679] = t[55678] ^ n[55679];
assign t[55680] = t[55679] ^ n[55680];
assign t[55681] = t[55680] ^ n[55681];
assign t[55682] = t[55681] ^ n[55682];
assign t[55683] = t[55682] ^ n[55683];
assign t[55684] = t[55683] ^ n[55684];
assign t[55685] = t[55684] ^ n[55685];
assign t[55686] = t[55685] ^ n[55686];
assign t[55687] = t[55686] ^ n[55687];
assign t[55688] = t[55687] ^ n[55688];
assign t[55689] = t[55688] ^ n[55689];
assign t[55690] = t[55689] ^ n[55690];
assign t[55691] = t[55690] ^ n[55691];
assign t[55692] = t[55691] ^ n[55692];
assign t[55693] = t[55692] ^ n[55693];
assign t[55694] = t[55693] ^ n[55694];
assign t[55695] = t[55694] ^ n[55695];
assign t[55696] = t[55695] ^ n[55696];
assign t[55697] = t[55696] ^ n[55697];
assign t[55698] = t[55697] ^ n[55698];
assign t[55699] = t[55698] ^ n[55699];
assign t[55700] = t[55699] ^ n[55700];
assign t[55701] = t[55700] ^ n[55701];
assign t[55702] = t[55701] ^ n[55702];
assign t[55703] = t[55702] ^ n[55703];
assign t[55704] = t[55703] ^ n[55704];
assign t[55705] = t[55704] ^ n[55705];
assign t[55706] = t[55705] ^ n[55706];
assign t[55707] = t[55706] ^ n[55707];
assign t[55708] = t[55707] ^ n[55708];
assign t[55709] = t[55708] ^ n[55709];
assign t[55710] = t[55709] ^ n[55710];
assign t[55711] = t[55710] ^ n[55711];
assign t[55712] = t[55711] ^ n[55712];
assign t[55713] = t[55712] ^ n[55713];
assign t[55714] = t[55713] ^ n[55714];
assign t[55715] = t[55714] ^ n[55715];
assign t[55716] = t[55715] ^ n[55716];
assign t[55717] = t[55716] ^ n[55717];
assign t[55718] = t[55717] ^ n[55718];
assign t[55719] = t[55718] ^ n[55719];
assign t[55720] = t[55719] ^ n[55720];
assign t[55721] = t[55720] ^ n[55721];
assign t[55722] = t[55721] ^ n[55722];
assign t[55723] = t[55722] ^ n[55723];
assign t[55724] = t[55723] ^ n[55724];
assign t[55725] = t[55724] ^ n[55725];
assign t[55726] = t[55725] ^ n[55726];
assign t[55727] = t[55726] ^ n[55727];
assign t[55728] = t[55727] ^ n[55728];
assign t[55729] = t[55728] ^ n[55729];
assign t[55730] = t[55729] ^ n[55730];
assign t[55731] = t[55730] ^ n[55731];
assign t[55732] = t[55731] ^ n[55732];
assign t[55733] = t[55732] ^ n[55733];
assign t[55734] = t[55733] ^ n[55734];
assign t[55735] = t[55734] ^ n[55735];
assign t[55736] = t[55735] ^ n[55736];
assign t[55737] = t[55736] ^ n[55737];
assign t[55738] = t[55737] ^ n[55738];
assign t[55739] = t[55738] ^ n[55739];
assign t[55740] = t[55739] ^ n[55740];
assign t[55741] = t[55740] ^ n[55741];
assign t[55742] = t[55741] ^ n[55742];
assign t[55743] = t[55742] ^ n[55743];
assign t[55744] = t[55743] ^ n[55744];
assign t[55745] = t[55744] ^ n[55745];
assign t[55746] = t[55745] ^ n[55746];
assign t[55747] = t[55746] ^ n[55747];
assign t[55748] = t[55747] ^ n[55748];
assign t[55749] = t[55748] ^ n[55749];
assign t[55750] = t[55749] ^ n[55750];
assign t[55751] = t[55750] ^ n[55751];
assign t[55752] = t[55751] ^ n[55752];
assign t[55753] = t[55752] ^ n[55753];
assign t[55754] = t[55753] ^ n[55754];
assign t[55755] = t[55754] ^ n[55755];
assign t[55756] = t[55755] ^ n[55756];
assign t[55757] = t[55756] ^ n[55757];
assign t[55758] = t[55757] ^ n[55758];
assign t[55759] = t[55758] ^ n[55759];
assign t[55760] = t[55759] ^ n[55760];
assign t[55761] = t[55760] ^ n[55761];
assign t[55762] = t[55761] ^ n[55762];
assign t[55763] = t[55762] ^ n[55763];
assign t[55764] = t[55763] ^ n[55764];
assign t[55765] = t[55764] ^ n[55765];
assign t[55766] = t[55765] ^ n[55766];
assign t[55767] = t[55766] ^ n[55767];
assign t[55768] = t[55767] ^ n[55768];
assign t[55769] = t[55768] ^ n[55769];
assign t[55770] = t[55769] ^ n[55770];
assign t[55771] = t[55770] ^ n[55771];
assign t[55772] = t[55771] ^ n[55772];
assign t[55773] = t[55772] ^ n[55773];
assign t[55774] = t[55773] ^ n[55774];
assign t[55775] = t[55774] ^ n[55775];
assign t[55776] = t[55775] ^ n[55776];
assign t[55777] = t[55776] ^ n[55777];
assign t[55778] = t[55777] ^ n[55778];
assign t[55779] = t[55778] ^ n[55779];
assign t[55780] = t[55779] ^ n[55780];
assign t[55781] = t[55780] ^ n[55781];
assign t[55782] = t[55781] ^ n[55782];
assign t[55783] = t[55782] ^ n[55783];
assign t[55784] = t[55783] ^ n[55784];
assign t[55785] = t[55784] ^ n[55785];
assign t[55786] = t[55785] ^ n[55786];
assign t[55787] = t[55786] ^ n[55787];
assign t[55788] = t[55787] ^ n[55788];
assign t[55789] = t[55788] ^ n[55789];
assign t[55790] = t[55789] ^ n[55790];
assign t[55791] = t[55790] ^ n[55791];
assign t[55792] = t[55791] ^ n[55792];
assign t[55793] = t[55792] ^ n[55793];
assign t[55794] = t[55793] ^ n[55794];
assign t[55795] = t[55794] ^ n[55795];
assign t[55796] = t[55795] ^ n[55796];
assign t[55797] = t[55796] ^ n[55797];
assign t[55798] = t[55797] ^ n[55798];
assign t[55799] = t[55798] ^ n[55799];
assign t[55800] = t[55799] ^ n[55800];
assign t[55801] = t[55800] ^ n[55801];
assign t[55802] = t[55801] ^ n[55802];
assign t[55803] = t[55802] ^ n[55803];
assign t[55804] = t[55803] ^ n[55804];
assign t[55805] = t[55804] ^ n[55805];
assign t[55806] = t[55805] ^ n[55806];
assign t[55807] = t[55806] ^ n[55807];
assign t[55808] = t[55807] ^ n[55808];
assign t[55809] = t[55808] ^ n[55809];
assign t[55810] = t[55809] ^ n[55810];
assign t[55811] = t[55810] ^ n[55811];
assign t[55812] = t[55811] ^ n[55812];
assign t[55813] = t[55812] ^ n[55813];
assign t[55814] = t[55813] ^ n[55814];
assign t[55815] = t[55814] ^ n[55815];
assign t[55816] = t[55815] ^ n[55816];
assign t[55817] = t[55816] ^ n[55817];
assign t[55818] = t[55817] ^ n[55818];
assign t[55819] = t[55818] ^ n[55819];
assign t[55820] = t[55819] ^ n[55820];
assign t[55821] = t[55820] ^ n[55821];
assign t[55822] = t[55821] ^ n[55822];
assign t[55823] = t[55822] ^ n[55823];
assign t[55824] = t[55823] ^ n[55824];
assign t[55825] = t[55824] ^ n[55825];
assign t[55826] = t[55825] ^ n[55826];
assign t[55827] = t[55826] ^ n[55827];
assign t[55828] = t[55827] ^ n[55828];
assign t[55829] = t[55828] ^ n[55829];
assign t[55830] = t[55829] ^ n[55830];
assign t[55831] = t[55830] ^ n[55831];
assign t[55832] = t[55831] ^ n[55832];
assign t[55833] = t[55832] ^ n[55833];
assign t[55834] = t[55833] ^ n[55834];
assign t[55835] = t[55834] ^ n[55835];
assign t[55836] = t[55835] ^ n[55836];
assign t[55837] = t[55836] ^ n[55837];
assign t[55838] = t[55837] ^ n[55838];
assign t[55839] = t[55838] ^ n[55839];
assign t[55840] = t[55839] ^ n[55840];
assign t[55841] = t[55840] ^ n[55841];
assign t[55842] = t[55841] ^ n[55842];
assign t[55843] = t[55842] ^ n[55843];
assign t[55844] = t[55843] ^ n[55844];
assign t[55845] = t[55844] ^ n[55845];
assign t[55846] = t[55845] ^ n[55846];
assign t[55847] = t[55846] ^ n[55847];
assign t[55848] = t[55847] ^ n[55848];
assign t[55849] = t[55848] ^ n[55849];
assign t[55850] = t[55849] ^ n[55850];
assign t[55851] = t[55850] ^ n[55851];
assign t[55852] = t[55851] ^ n[55852];
assign t[55853] = t[55852] ^ n[55853];
assign t[55854] = t[55853] ^ n[55854];
assign t[55855] = t[55854] ^ n[55855];
assign t[55856] = t[55855] ^ n[55856];
assign t[55857] = t[55856] ^ n[55857];
assign t[55858] = t[55857] ^ n[55858];
assign t[55859] = t[55858] ^ n[55859];
assign t[55860] = t[55859] ^ n[55860];
assign t[55861] = t[55860] ^ n[55861];
assign t[55862] = t[55861] ^ n[55862];
assign t[55863] = t[55862] ^ n[55863];
assign t[55864] = t[55863] ^ n[55864];
assign t[55865] = t[55864] ^ n[55865];
assign t[55866] = t[55865] ^ n[55866];
assign t[55867] = t[55866] ^ n[55867];
assign t[55868] = t[55867] ^ n[55868];
assign t[55869] = t[55868] ^ n[55869];
assign t[55870] = t[55869] ^ n[55870];
assign t[55871] = t[55870] ^ n[55871];
assign t[55872] = t[55871] ^ n[55872];
assign t[55873] = t[55872] ^ n[55873];
assign t[55874] = t[55873] ^ n[55874];
assign t[55875] = t[55874] ^ n[55875];
assign t[55876] = t[55875] ^ n[55876];
assign t[55877] = t[55876] ^ n[55877];
assign t[55878] = t[55877] ^ n[55878];
assign t[55879] = t[55878] ^ n[55879];
assign t[55880] = t[55879] ^ n[55880];
assign t[55881] = t[55880] ^ n[55881];
assign t[55882] = t[55881] ^ n[55882];
assign t[55883] = t[55882] ^ n[55883];
assign t[55884] = t[55883] ^ n[55884];
assign t[55885] = t[55884] ^ n[55885];
assign t[55886] = t[55885] ^ n[55886];
assign t[55887] = t[55886] ^ n[55887];
assign t[55888] = t[55887] ^ n[55888];
assign t[55889] = t[55888] ^ n[55889];
assign t[55890] = t[55889] ^ n[55890];
assign t[55891] = t[55890] ^ n[55891];
assign t[55892] = t[55891] ^ n[55892];
assign t[55893] = t[55892] ^ n[55893];
assign t[55894] = t[55893] ^ n[55894];
assign t[55895] = t[55894] ^ n[55895];
assign t[55896] = t[55895] ^ n[55896];
assign t[55897] = t[55896] ^ n[55897];
assign t[55898] = t[55897] ^ n[55898];
assign t[55899] = t[55898] ^ n[55899];
assign t[55900] = t[55899] ^ n[55900];
assign t[55901] = t[55900] ^ n[55901];
assign t[55902] = t[55901] ^ n[55902];
assign t[55903] = t[55902] ^ n[55903];
assign t[55904] = t[55903] ^ n[55904];
assign t[55905] = t[55904] ^ n[55905];
assign t[55906] = t[55905] ^ n[55906];
assign t[55907] = t[55906] ^ n[55907];
assign t[55908] = t[55907] ^ n[55908];
assign t[55909] = t[55908] ^ n[55909];
assign t[55910] = t[55909] ^ n[55910];
assign t[55911] = t[55910] ^ n[55911];
assign t[55912] = t[55911] ^ n[55912];
assign t[55913] = t[55912] ^ n[55913];
assign t[55914] = t[55913] ^ n[55914];
assign t[55915] = t[55914] ^ n[55915];
assign t[55916] = t[55915] ^ n[55916];
assign t[55917] = t[55916] ^ n[55917];
assign t[55918] = t[55917] ^ n[55918];
assign t[55919] = t[55918] ^ n[55919];
assign t[55920] = t[55919] ^ n[55920];
assign t[55921] = t[55920] ^ n[55921];
assign t[55922] = t[55921] ^ n[55922];
assign t[55923] = t[55922] ^ n[55923];
assign t[55924] = t[55923] ^ n[55924];
assign t[55925] = t[55924] ^ n[55925];
assign t[55926] = t[55925] ^ n[55926];
assign t[55927] = t[55926] ^ n[55927];
assign t[55928] = t[55927] ^ n[55928];
assign t[55929] = t[55928] ^ n[55929];
assign t[55930] = t[55929] ^ n[55930];
assign t[55931] = t[55930] ^ n[55931];
assign t[55932] = t[55931] ^ n[55932];
assign t[55933] = t[55932] ^ n[55933];
assign t[55934] = t[55933] ^ n[55934];
assign t[55935] = t[55934] ^ n[55935];
assign t[55936] = t[55935] ^ n[55936];
assign t[55937] = t[55936] ^ n[55937];
assign t[55938] = t[55937] ^ n[55938];
assign t[55939] = t[55938] ^ n[55939];
assign t[55940] = t[55939] ^ n[55940];
assign t[55941] = t[55940] ^ n[55941];
assign t[55942] = t[55941] ^ n[55942];
assign t[55943] = t[55942] ^ n[55943];
assign t[55944] = t[55943] ^ n[55944];
assign t[55945] = t[55944] ^ n[55945];
assign t[55946] = t[55945] ^ n[55946];
assign t[55947] = t[55946] ^ n[55947];
assign t[55948] = t[55947] ^ n[55948];
assign t[55949] = t[55948] ^ n[55949];
assign t[55950] = t[55949] ^ n[55950];
assign t[55951] = t[55950] ^ n[55951];
assign t[55952] = t[55951] ^ n[55952];
assign t[55953] = t[55952] ^ n[55953];
assign t[55954] = t[55953] ^ n[55954];
assign t[55955] = t[55954] ^ n[55955];
assign t[55956] = t[55955] ^ n[55956];
assign t[55957] = t[55956] ^ n[55957];
assign t[55958] = t[55957] ^ n[55958];
assign t[55959] = t[55958] ^ n[55959];
assign t[55960] = t[55959] ^ n[55960];
assign t[55961] = t[55960] ^ n[55961];
assign t[55962] = t[55961] ^ n[55962];
assign t[55963] = t[55962] ^ n[55963];
assign t[55964] = t[55963] ^ n[55964];
assign t[55965] = t[55964] ^ n[55965];
assign t[55966] = t[55965] ^ n[55966];
assign t[55967] = t[55966] ^ n[55967];
assign t[55968] = t[55967] ^ n[55968];
assign t[55969] = t[55968] ^ n[55969];
assign t[55970] = t[55969] ^ n[55970];
assign t[55971] = t[55970] ^ n[55971];
assign t[55972] = t[55971] ^ n[55972];
assign t[55973] = t[55972] ^ n[55973];
assign t[55974] = t[55973] ^ n[55974];
assign t[55975] = t[55974] ^ n[55975];
assign t[55976] = t[55975] ^ n[55976];
assign t[55977] = t[55976] ^ n[55977];
assign t[55978] = t[55977] ^ n[55978];
assign t[55979] = t[55978] ^ n[55979];
assign t[55980] = t[55979] ^ n[55980];
assign t[55981] = t[55980] ^ n[55981];
assign t[55982] = t[55981] ^ n[55982];
assign t[55983] = t[55982] ^ n[55983];
assign t[55984] = t[55983] ^ n[55984];
assign t[55985] = t[55984] ^ n[55985];
assign t[55986] = t[55985] ^ n[55986];
assign t[55987] = t[55986] ^ n[55987];
assign t[55988] = t[55987] ^ n[55988];
assign t[55989] = t[55988] ^ n[55989];
assign t[55990] = t[55989] ^ n[55990];
assign t[55991] = t[55990] ^ n[55991];
assign t[55992] = t[55991] ^ n[55992];
assign t[55993] = t[55992] ^ n[55993];
assign t[55994] = t[55993] ^ n[55994];
assign t[55995] = t[55994] ^ n[55995];
assign t[55996] = t[55995] ^ n[55996];
assign t[55997] = t[55996] ^ n[55997];
assign t[55998] = t[55997] ^ n[55998];
assign t[55999] = t[55998] ^ n[55999];
assign t[56000] = t[55999] ^ n[56000];
assign t[56001] = t[56000] ^ n[56001];
assign t[56002] = t[56001] ^ n[56002];
assign t[56003] = t[56002] ^ n[56003];
assign t[56004] = t[56003] ^ n[56004];
assign t[56005] = t[56004] ^ n[56005];
assign t[56006] = t[56005] ^ n[56006];
assign t[56007] = t[56006] ^ n[56007];
assign t[56008] = t[56007] ^ n[56008];
assign t[56009] = t[56008] ^ n[56009];
assign t[56010] = t[56009] ^ n[56010];
assign t[56011] = t[56010] ^ n[56011];
assign t[56012] = t[56011] ^ n[56012];
assign t[56013] = t[56012] ^ n[56013];
assign t[56014] = t[56013] ^ n[56014];
assign t[56015] = t[56014] ^ n[56015];
assign t[56016] = t[56015] ^ n[56016];
assign t[56017] = t[56016] ^ n[56017];
assign t[56018] = t[56017] ^ n[56018];
assign t[56019] = t[56018] ^ n[56019];
assign t[56020] = t[56019] ^ n[56020];
assign t[56021] = t[56020] ^ n[56021];
assign t[56022] = t[56021] ^ n[56022];
assign t[56023] = t[56022] ^ n[56023];
assign t[56024] = t[56023] ^ n[56024];
assign t[56025] = t[56024] ^ n[56025];
assign t[56026] = t[56025] ^ n[56026];
assign t[56027] = t[56026] ^ n[56027];
assign t[56028] = t[56027] ^ n[56028];
assign t[56029] = t[56028] ^ n[56029];
assign t[56030] = t[56029] ^ n[56030];
assign t[56031] = t[56030] ^ n[56031];
assign t[56032] = t[56031] ^ n[56032];
assign t[56033] = t[56032] ^ n[56033];
assign t[56034] = t[56033] ^ n[56034];
assign t[56035] = t[56034] ^ n[56035];
assign t[56036] = t[56035] ^ n[56036];
assign t[56037] = t[56036] ^ n[56037];
assign t[56038] = t[56037] ^ n[56038];
assign t[56039] = t[56038] ^ n[56039];
assign t[56040] = t[56039] ^ n[56040];
assign t[56041] = t[56040] ^ n[56041];
assign t[56042] = t[56041] ^ n[56042];
assign t[56043] = t[56042] ^ n[56043];
assign t[56044] = t[56043] ^ n[56044];
assign t[56045] = t[56044] ^ n[56045];
assign t[56046] = t[56045] ^ n[56046];
assign t[56047] = t[56046] ^ n[56047];
assign t[56048] = t[56047] ^ n[56048];
assign t[56049] = t[56048] ^ n[56049];
assign t[56050] = t[56049] ^ n[56050];
assign t[56051] = t[56050] ^ n[56051];
assign t[56052] = t[56051] ^ n[56052];
assign t[56053] = t[56052] ^ n[56053];
assign t[56054] = t[56053] ^ n[56054];
assign t[56055] = t[56054] ^ n[56055];
assign t[56056] = t[56055] ^ n[56056];
assign t[56057] = t[56056] ^ n[56057];
assign t[56058] = t[56057] ^ n[56058];
assign t[56059] = t[56058] ^ n[56059];
assign t[56060] = t[56059] ^ n[56060];
assign t[56061] = t[56060] ^ n[56061];
assign t[56062] = t[56061] ^ n[56062];
assign t[56063] = t[56062] ^ n[56063];
assign t[56064] = t[56063] ^ n[56064];
assign t[56065] = t[56064] ^ n[56065];
assign t[56066] = t[56065] ^ n[56066];
assign t[56067] = t[56066] ^ n[56067];
assign t[56068] = t[56067] ^ n[56068];
assign t[56069] = t[56068] ^ n[56069];
assign t[56070] = t[56069] ^ n[56070];
assign t[56071] = t[56070] ^ n[56071];
assign t[56072] = t[56071] ^ n[56072];
assign t[56073] = t[56072] ^ n[56073];
assign t[56074] = t[56073] ^ n[56074];
assign t[56075] = t[56074] ^ n[56075];
assign t[56076] = t[56075] ^ n[56076];
assign t[56077] = t[56076] ^ n[56077];
assign t[56078] = t[56077] ^ n[56078];
assign t[56079] = t[56078] ^ n[56079];
assign t[56080] = t[56079] ^ n[56080];
assign t[56081] = t[56080] ^ n[56081];
assign t[56082] = t[56081] ^ n[56082];
assign t[56083] = t[56082] ^ n[56083];
assign t[56084] = t[56083] ^ n[56084];
assign t[56085] = t[56084] ^ n[56085];
assign t[56086] = t[56085] ^ n[56086];
assign t[56087] = t[56086] ^ n[56087];
assign t[56088] = t[56087] ^ n[56088];
assign t[56089] = t[56088] ^ n[56089];
assign t[56090] = t[56089] ^ n[56090];
assign t[56091] = t[56090] ^ n[56091];
assign t[56092] = t[56091] ^ n[56092];
assign t[56093] = t[56092] ^ n[56093];
assign t[56094] = t[56093] ^ n[56094];
assign t[56095] = t[56094] ^ n[56095];
assign t[56096] = t[56095] ^ n[56096];
assign t[56097] = t[56096] ^ n[56097];
assign t[56098] = t[56097] ^ n[56098];
assign t[56099] = t[56098] ^ n[56099];
assign t[56100] = t[56099] ^ n[56100];
assign t[56101] = t[56100] ^ n[56101];
assign t[56102] = t[56101] ^ n[56102];
assign t[56103] = t[56102] ^ n[56103];
assign t[56104] = t[56103] ^ n[56104];
assign t[56105] = t[56104] ^ n[56105];
assign t[56106] = t[56105] ^ n[56106];
assign t[56107] = t[56106] ^ n[56107];
assign t[56108] = t[56107] ^ n[56108];
assign t[56109] = t[56108] ^ n[56109];
assign t[56110] = t[56109] ^ n[56110];
assign t[56111] = t[56110] ^ n[56111];
assign t[56112] = t[56111] ^ n[56112];
assign t[56113] = t[56112] ^ n[56113];
assign t[56114] = t[56113] ^ n[56114];
assign t[56115] = t[56114] ^ n[56115];
assign t[56116] = t[56115] ^ n[56116];
assign t[56117] = t[56116] ^ n[56117];
assign t[56118] = t[56117] ^ n[56118];
assign t[56119] = t[56118] ^ n[56119];
assign t[56120] = t[56119] ^ n[56120];
assign t[56121] = t[56120] ^ n[56121];
assign t[56122] = t[56121] ^ n[56122];
assign t[56123] = t[56122] ^ n[56123];
assign t[56124] = t[56123] ^ n[56124];
assign t[56125] = t[56124] ^ n[56125];
assign t[56126] = t[56125] ^ n[56126];
assign t[56127] = t[56126] ^ n[56127];
assign t[56128] = t[56127] ^ n[56128];
assign t[56129] = t[56128] ^ n[56129];
assign t[56130] = t[56129] ^ n[56130];
assign t[56131] = t[56130] ^ n[56131];
assign t[56132] = t[56131] ^ n[56132];
assign t[56133] = t[56132] ^ n[56133];
assign t[56134] = t[56133] ^ n[56134];
assign t[56135] = t[56134] ^ n[56135];
assign t[56136] = t[56135] ^ n[56136];
assign t[56137] = t[56136] ^ n[56137];
assign t[56138] = t[56137] ^ n[56138];
assign t[56139] = t[56138] ^ n[56139];
assign t[56140] = t[56139] ^ n[56140];
assign t[56141] = t[56140] ^ n[56141];
assign t[56142] = t[56141] ^ n[56142];
assign t[56143] = t[56142] ^ n[56143];
assign t[56144] = t[56143] ^ n[56144];
assign t[56145] = t[56144] ^ n[56145];
assign t[56146] = t[56145] ^ n[56146];
assign t[56147] = t[56146] ^ n[56147];
assign t[56148] = t[56147] ^ n[56148];
assign t[56149] = t[56148] ^ n[56149];
assign t[56150] = t[56149] ^ n[56150];
assign t[56151] = t[56150] ^ n[56151];
assign t[56152] = t[56151] ^ n[56152];
assign t[56153] = t[56152] ^ n[56153];
assign t[56154] = t[56153] ^ n[56154];
assign t[56155] = t[56154] ^ n[56155];
assign t[56156] = t[56155] ^ n[56156];
assign t[56157] = t[56156] ^ n[56157];
assign t[56158] = t[56157] ^ n[56158];
assign t[56159] = t[56158] ^ n[56159];
assign t[56160] = t[56159] ^ n[56160];
assign t[56161] = t[56160] ^ n[56161];
assign t[56162] = t[56161] ^ n[56162];
assign t[56163] = t[56162] ^ n[56163];
assign t[56164] = t[56163] ^ n[56164];
assign t[56165] = t[56164] ^ n[56165];
assign t[56166] = t[56165] ^ n[56166];
assign t[56167] = t[56166] ^ n[56167];
assign t[56168] = t[56167] ^ n[56168];
assign t[56169] = t[56168] ^ n[56169];
assign t[56170] = t[56169] ^ n[56170];
assign t[56171] = t[56170] ^ n[56171];
assign t[56172] = t[56171] ^ n[56172];
assign t[56173] = t[56172] ^ n[56173];
assign t[56174] = t[56173] ^ n[56174];
assign t[56175] = t[56174] ^ n[56175];
assign t[56176] = t[56175] ^ n[56176];
assign t[56177] = t[56176] ^ n[56177];
assign t[56178] = t[56177] ^ n[56178];
assign t[56179] = t[56178] ^ n[56179];
assign t[56180] = t[56179] ^ n[56180];
assign t[56181] = t[56180] ^ n[56181];
assign t[56182] = t[56181] ^ n[56182];
assign t[56183] = t[56182] ^ n[56183];
assign t[56184] = t[56183] ^ n[56184];
assign t[56185] = t[56184] ^ n[56185];
assign t[56186] = t[56185] ^ n[56186];
assign t[56187] = t[56186] ^ n[56187];
assign t[56188] = t[56187] ^ n[56188];
assign t[56189] = t[56188] ^ n[56189];
assign t[56190] = t[56189] ^ n[56190];
assign t[56191] = t[56190] ^ n[56191];
assign t[56192] = t[56191] ^ n[56192];
assign t[56193] = t[56192] ^ n[56193];
assign t[56194] = t[56193] ^ n[56194];
assign t[56195] = t[56194] ^ n[56195];
assign t[56196] = t[56195] ^ n[56196];
assign t[56197] = t[56196] ^ n[56197];
assign t[56198] = t[56197] ^ n[56198];
assign t[56199] = t[56198] ^ n[56199];
assign t[56200] = t[56199] ^ n[56200];
assign t[56201] = t[56200] ^ n[56201];
assign t[56202] = t[56201] ^ n[56202];
assign t[56203] = t[56202] ^ n[56203];
assign t[56204] = t[56203] ^ n[56204];
assign t[56205] = t[56204] ^ n[56205];
assign t[56206] = t[56205] ^ n[56206];
assign t[56207] = t[56206] ^ n[56207];
assign t[56208] = t[56207] ^ n[56208];
assign t[56209] = t[56208] ^ n[56209];
assign t[56210] = t[56209] ^ n[56210];
assign t[56211] = t[56210] ^ n[56211];
assign t[56212] = t[56211] ^ n[56212];
assign t[56213] = t[56212] ^ n[56213];
assign t[56214] = t[56213] ^ n[56214];
assign t[56215] = t[56214] ^ n[56215];
assign t[56216] = t[56215] ^ n[56216];
assign t[56217] = t[56216] ^ n[56217];
assign t[56218] = t[56217] ^ n[56218];
assign t[56219] = t[56218] ^ n[56219];
assign t[56220] = t[56219] ^ n[56220];
assign t[56221] = t[56220] ^ n[56221];
assign t[56222] = t[56221] ^ n[56222];
assign t[56223] = t[56222] ^ n[56223];
assign t[56224] = t[56223] ^ n[56224];
assign t[56225] = t[56224] ^ n[56225];
assign t[56226] = t[56225] ^ n[56226];
assign t[56227] = t[56226] ^ n[56227];
assign t[56228] = t[56227] ^ n[56228];
assign t[56229] = t[56228] ^ n[56229];
assign t[56230] = t[56229] ^ n[56230];
assign t[56231] = t[56230] ^ n[56231];
assign t[56232] = t[56231] ^ n[56232];
assign t[56233] = t[56232] ^ n[56233];
assign t[56234] = t[56233] ^ n[56234];
assign t[56235] = t[56234] ^ n[56235];
assign t[56236] = t[56235] ^ n[56236];
assign t[56237] = t[56236] ^ n[56237];
assign t[56238] = t[56237] ^ n[56238];
assign t[56239] = t[56238] ^ n[56239];
assign t[56240] = t[56239] ^ n[56240];
assign t[56241] = t[56240] ^ n[56241];
assign t[56242] = t[56241] ^ n[56242];
assign t[56243] = t[56242] ^ n[56243];
assign t[56244] = t[56243] ^ n[56244];
assign t[56245] = t[56244] ^ n[56245];
assign t[56246] = t[56245] ^ n[56246];
assign t[56247] = t[56246] ^ n[56247];
assign t[56248] = t[56247] ^ n[56248];
assign t[56249] = t[56248] ^ n[56249];
assign t[56250] = t[56249] ^ n[56250];
assign t[56251] = t[56250] ^ n[56251];
assign t[56252] = t[56251] ^ n[56252];
assign t[56253] = t[56252] ^ n[56253];
assign t[56254] = t[56253] ^ n[56254];
assign t[56255] = t[56254] ^ n[56255];
assign t[56256] = t[56255] ^ n[56256];
assign t[56257] = t[56256] ^ n[56257];
assign t[56258] = t[56257] ^ n[56258];
assign t[56259] = t[56258] ^ n[56259];
assign t[56260] = t[56259] ^ n[56260];
assign t[56261] = t[56260] ^ n[56261];
assign t[56262] = t[56261] ^ n[56262];
assign t[56263] = t[56262] ^ n[56263];
assign t[56264] = t[56263] ^ n[56264];
assign t[56265] = t[56264] ^ n[56265];
assign t[56266] = t[56265] ^ n[56266];
assign t[56267] = t[56266] ^ n[56267];
assign t[56268] = t[56267] ^ n[56268];
assign t[56269] = t[56268] ^ n[56269];
assign t[56270] = t[56269] ^ n[56270];
assign t[56271] = t[56270] ^ n[56271];
assign t[56272] = t[56271] ^ n[56272];
assign t[56273] = t[56272] ^ n[56273];
assign t[56274] = t[56273] ^ n[56274];
assign t[56275] = t[56274] ^ n[56275];
assign t[56276] = t[56275] ^ n[56276];
assign t[56277] = t[56276] ^ n[56277];
assign t[56278] = t[56277] ^ n[56278];
assign t[56279] = t[56278] ^ n[56279];
assign t[56280] = t[56279] ^ n[56280];
assign t[56281] = t[56280] ^ n[56281];
assign t[56282] = t[56281] ^ n[56282];
assign t[56283] = t[56282] ^ n[56283];
assign t[56284] = t[56283] ^ n[56284];
assign t[56285] = t[56284] ^ n[56285];
assign t[56286] = t[56285] ^ n[56286];
assign t[56287] = t[56286] ^ n[56287];
assign t[56288] = t[56287] ^ n[56288];
assign t[56289] = t[56288] ^ n[56289];
assign t[56290] = t[56289] ^ n[56290];
assign t[56291] = t[56290] ^ n[56291];
assign t[56292] = t[56291] ^ n[56292];
assign t[56293] = t[56292] ^ n[56293];
assign t[56294] = t[56293] ^ n[56294];
assign t[56295] = t[56294] ^ n[56295];
assign t[56296] = t[56295] ^ n[56296];
assign t[56297] = t[56296] ^ n[56297];
assign t[56298] = t[56297] ^ n[56298];
assign t[56299] = t[56298] ^ n[56299];
assign t[56300] = t[56299] ^ n[56300];
assign t[56301] = t[56300] ^ n[56301];
assign t[56302] = t[56301] ^ n[56302];
assign t[56303] = t[56302] ^ n[56303];
assign t[56304] = t[56303] ^ n[56304];
assign t[56305] = t[56304] ^ n[56305];
assign t[56306] = t[56305] ^ n[56306];
assign t[56307] = t[56306] ^ n[56307];
assign t[56308] = t[56307] ^ n[56308];
assign t[56309] = t[56308] ^ n[56309];
assign t[56310] = t[56309] ^ n[56310];
assign t[56311] = t[56310] ^ n[56311];
assign t[56312] = t[56311] ^ n[56312];
assign t[56313] = t[56312] ^ n[56313];
assign t[56314] = t[56313] ^ n[56314];
assign t[56315] = t[56314] ^ n[56315];
assign t[56316] = t[56315] ^ n[56316];
assign t[56317] = t[56316] ^ n[56317];
assign t[56318] = t[56317] ^ n[56318];
assign t[56319] = t[56318] ^ n[56319];
assign t[56320] = t[56319] ^ n[56320];
assign t[56321] = t[56320] ^ n[56321];
assign t[56322] = t[56321] ^ n[56322];
assign t[56323] = t[56322] ^ n[56323];
assign t[56324] = t[56323] ^ n[56324];
assign t[56325] = t[56324] ^ n[56325];
assign t[56326] = t[56325] ^ n[56326];
assign t[56327] = t[56326] ^ n[56327];
assign t[56328] = t[56327] ^ n[56328];
assign t[56329] = t[56328] ^ n[56329];
assign t[56330] = t[56329] ^ n[56330];
assign t[56331] = t[56330] ^ n[56331];
assign t[56332] = t[56331] ^ n[56332];
assign t[56333] = t[56332] ^ n[56333];
assign t[56334] = t[56333] ^ n[56334];
assign t[56335] = t[56334] ^ n[56335];
assign t[56336] = t[56335] ^ n[56336];
assign t[56337] = t[56336] ^ n[56337];
assign t[56338] = t[56337] ^ n[56338];
assign t[56339] = t[56338] ^ n[56339];
assign t[56340] = t[56339] ^ n[56340];
assign t[56341] = t[56340] ^ n[56341];
assign t[56342] = t[56341] ^ n[56342];
assign t[56343] = t[56342] ^ n[56343];
assign t[56344] = t[56343] ^ n[56344];
assign t[56345] = t[56344] ^ n[56345];
assign t[56346] = t[56345] ^ n[56346];
assign t[56347] = t[56346] ^ n[56347];
assign t[56348] = t[56347] ^ n[56348];
assign t[56349] = t[56348] ^ n[56349];
assign t[56350] = t[56349] ^ n[56350];
assign t[56351] = t[56350] ^ n[56351];
assign t[56352] = t[56351] ^ n[56352];
assign t[56353] = t[56352] ^ n[56353];
assign t[56354] = t[56353] ^ n[56354];
assign t[56355] = t[56354] ^ n[56355];
assign t[56356] = t[56355] ^ n[56356];
assign t[56357] = t[56356] ^ n[56357];
assign t[56358] = t[56357] ^ n[56358];
assign t[56359] = t[56358] ^ n[56359];
assign t[56360] = t[56359] ^ n[56360];
assign t[56361] = t[56360] ^ n[56361];
assign t[56362] = t[56361] ^ n[56362];
assign t[56363] = t[56362] ^ n[56363];
assign t[56364] = t[56363] ^ n[56364];
assign t[56365] = t[56364] ^ n[56365];
assign t[56366] = t[56365] ^ n[56366];
assign t[56367] = t[56366] ^ n[56367];
assign t[56368] = t[56367] ^ n[56368];
assign t[56369] = t[56368] ^ n[56369];
assign t[56370] = t[56369] ^ n[56370];
assign t[56371] = t[56370] ^ n[56371];
assign t[56372] = t[56371] ^ n[56372];
assign t[56373] = t[56372] ^ n[56373];
assign t[56374] = t[56373] ^ n[56374];
assign t[56375] = t[56374] ^ n[56375];
assign t[56376] = t[56375] ^ n[56376];
assign t[56377] = t[56376] ^ n[56377];
assign t[56378] = t[56377] ^ n[56378];
assign t[56379] = t[56378] ^ n[56379];
assign t[56380] = t[56379] ^ n[56380];
assign t[56381] = t[56380] ^ n[56381];
assign t[56382] = t[56381] ^ n[56382];
assign t[56383] = t[56382] ^ n[56383];
assign t[56384] = t[56383] ^ n[56384];
assign t[56385] = t[56384] ^ n[56385];
assign t[56386] = t[56385] ^ n[56386];
assign t[56387] = t[56386] ^ n[56387];
assign t[56388] = t[56387] ^ n[56388];
assign t[56389] = t[56388] ^ n[56389];
assign t[56390] = t[56389] ^ n[56390];
assign t[56391] = t[56390] ^ n[56391];
assign t[56392] = t[56391] ^ n[56392];
assign t[56393] = t[56392] ^ n[56393];
assign t[56394] = t[56393] ^ n[56394];
assign t[56395] = t[56394] ^ n[56395];
assign t[56396] = t[56395] ^ n[56396];
assign t[56397] = t[56396] ^ n[56397];
assign t[56398] = t[56397] ^ n[56398];
assign t[56399] = t[56398] ^ n[56399];
assign t[56400] = t[56399] ^ n[56400];
assign t[56401] = t[56400] ^ n[56401];
assign t[56402] = t[56401] ^ n[56402];
assign t[56403] = t[56402] ^ n[56403];
assign t[56404] = t[56403] ^ n[56404];
assign t[56405] = t[56404] ^ n[56405];
assign t[56406] = t[56405] ^ n[56406];
assign t[56407] = t[56406] ^ n[56407];
assign t[56408] = t[56407] ^ n[56408];
assign t[56409] = t[56408] ^ n[56409];
assign t[56410] = t[56409] ^ n[56410];
assign t[56411] = t[56410] ^ n[56411];
assign t[56412] = t[56411] ^ n[56412];
assign t[56413] = t[56412] ^ n[56413];
assign t[56414] = t[56413] ^ n[56414];
assign t[56415] = t[56414] ^ n[56415];
assign t[56416] = t[56415] ^ n[56416];
assign t[56417] = t[56416] ^ n[56417];
assign t[56418] = t[56417] ^ n[56418];
assign t[56419] = t[56418] ^ n[56419];
assign t[56420] = t[56419] ^ n[56420];
assign t[56421] = t[56420] ^ n[56421];
assign t[56422] = t[56421] ^ n[56422];
assign t[56423] = t[56422] ^ n[56423];
assign t[56424] = t[56423] ^ n[56424];
assign t[56425] = t[56424] ^ n[56425];
assign t[56426] = t[56425] ^ n[56426];
assign t[56427] = t[56426] ^ n[56427];
assign t[56428] = t[56427] ^ n[56428];
assign t[56429] = t[56428] ^ n[56429];
assign t[56430] = t[56429] ^ n[56430];
assign t[56431] = t[56430] ^ n[56431];
assign t[56432] = t[56431] ^ n[56432];
assign t[56433] = t[56432] ^ n[56433];
assign t[56434] = t[56433] ^ n[56434];
assign t[56435] = t[56434] ^ n[56435];
assign t[56436] = t[56435] ^ n[56436];
assign t[56437] = t[56436] ^ n[56437];
assign t[56438] = t[56437] ^ n[56438];
assign t[56439] = t[56438] ^ n[56439];
assign t[56440] = t[56439] ^ n[56440];
assign t[56441] = t[56440] ^ n[56441];
assign t[56442] = t[56441] ^ n[56442];
assign t[56443] = t[56442] ^ n[56443];
assign t[56444] = t[56443] ^ n[56444];
assign t[56445] = t[56444] ^ n[56445];
assign t[56446] = t[56445] ^ n[56446];
assign t[56447] = t[56446] ^ n[56447];
assign t[56448] = t[56447] ^ n[56448];
assign t[56449] = t[56448] ^ n[56449];
assign t[56450] = t[56449] ^ n[56450];
assign t[56451] = t[56450] ^ n[56451];
assign t[56452] = t[56451] ^ n[56452];
assign t[56453] = t[56452] ^ n[56453];
assign t[56454] = t[56453] ^ n[56454];
assign t[56455] = t[56454] ^ n[56455];
assign t[56456] = t[56455] ^ n[56456];
assign t[56457] = t[56456] ^ n[56457];
assign t[56458] = t[56457] ^ n[56458];
assign t[56459] = t[56458] ^ n[56459];
assign t[56460] = t[56459] ^ n[56460];
assign t[56461] = t[56460] ^ n[56461];
assign t[56462] = t[56461] ^ n[56462];
assign t[56463] = t[56462] ^ n[56463];
assign t[56464] = t[56463] ^ n[56464];
assign t[56465] = t[56464] ^ n[56465];
assign t[56466] = t[56465] ^ n[56466];
assign t[56467] = t[56466] ^ n[56467];
assign t[56468] = t[56467] ^ n[56468];
assign t[56469] = t[56468] ^ n[56469];
assign t[56470] = t[56469] ^ n[56470];
assign t[56471] = t[56470] ^ n[56471];
assign t[56472] = t[56471] ^ n[56472];
assign t[56473] = t[56472] ^ n[56473];
assign t[56474] = t[56473] ^ n[56474];
assign t[56475] = t[56474] ^ n[56475];
assign t[56476] = t[56475] ^ n[56476];
assign t[56477] = t[56476] ^ n[56477];
assign t[56478] = t[56477] ^ n[56478];
assign t[56479] = t[56478] ^ n[56479];
assign t[56480] = t[56479] ^ n[56480];
assign t[56481] = t[56480] ^ n[56481];
assign t[56482] = t[56481] ^ n[56482];
assign t[56483] = t[56482] ^ n[56483];
assign t[56484] = t[56483] ^ n[56484];
assign t[56485] = t[56484] ^ n[56485];
assign t[56486] = t[56485] ^ n[56486];
assign t[56487] = t[56486] ^ n[56487];
assign t[56488] = t[56487] ^ n[56488];
assign t[56489] = t[56488] ^ n[56489];
assign t[56490] = t[56489] ^ n[56490];
assign t[56491] = t[56490] ^ n[56491];
assign t[56492] = t[56491] ^ n[56492];
assign t[56493] = t[56492] ^ n[56493];
assign t[56494] = t[56493] ^ n[56494];
assign t[56495] = t[56494] ^ n[56495];
assign t[56496] = t[56495] ^ n[56496];
assign t[56497] = t[56496] ^ n[56497];
assign t[56498] = t[56497] ^ n[56498];
assign t[56499] = t[56498] ^ n[56499];
assign t[56500] = t[56499] ^ n[56500];
assign t[56501] = t[56500] ^ n[56501];
assign t[56502] = t[56501] ^ n[56502];
assign t[56503] = t[56502] ^ n[56503];
assign t[56504] = t[56503] ^ n[56504];
assign t[56505] = t[56504] ^ n[56505];
assign t[56506] = t[56505] ^ n[56506];
assign t[56507] = t[56506] ^ n[56507];
assign t[56508] = t[56507] ^ n[56508];
assign t[56509] = t[56508] ^ n[56509];
assign t[56510] = t[56509] ^ n[56510];
assign t[56511] = t[56510] ^ n[56511];
assign t[56512] = t[56511] ^ n[56512];
assign t[56513] = t[56512] ^ n[56513];
assign t[56514] = t[56513] ^ n[56514];
assign t[56515] = t[56514] ^ n[56515];
assign t[56516] = t[56515] ^ n[56516];
assign t[56517] = t[56516] ^ n[56517];
assign t[56518] = t[56517] ^ n[56518];
assign t[56519] = t[56518] ^ n[56519];
assign t[56520] = t[56519] ^ n[56520];
assign t[56521] = t[56520] ^ n[56521];
assign t[56522] = t[56521] ^ n[56522];
assign t[56523] = t[56522] ^ n[56523];
assign t[56524] = t[56523] ^ n[56524];
assign t[56525] = t[56524] ^ n[56525];
assign t[56526] = t[56525] ^ n[56526];
assign t[56527] = t[56526] ^ n[56527];
assign t[56528] = t[56527] ^ n[56528];
assign t[56529] = t[56528] ^ n[56529];
assign t[56530] = t[56529] ^ n[56530];
assign t[56531] = t[56530] ^ n[56531];
assign t[56532] = t[56531] ^ n[56532];
assign t[56533] = t[56532] ^ n[56533];
assign t[56534] = t[56533] ^ n[56534];
assign t[56535] = t[56534] ^ n[56535];
assign t[56536] = t[56535] ^ n[56536];
assign t[56537] = t[56536] ^ n[56537];
assign t[56538] = t[56537] ^ n[56538];
assign t[56539] = t[56538] ^ n[56539];
assign t[56540] = t[56539] ^ n[56540];
assign t[56541] = t[56540] ^ n[56541];
assign t[56542] = t[56541] ^ n[56542];
assign t[56543] = t[56542] ^ n[56543];
assign t[56544] = t[56543] ^ n[56544];
assign t[56545] = t[56544] ^ n[56545];
assign t[56546] = t[56545] ^ n[56546];
assign t[56547] = t[56546] ^ n[56547];
assign t[56548] = t[56547] ^ n[56548];
assign t[56549] = t[56548] ^ n[56549];
assign t[56550] = t[56549] ^ n[56550];
assign t[56551] = t[56550] ^ n[56551];
assign t[56552] = t[56551] ^ n[56552];
assign t[56553] = t[56552] ^ n[56553];
assign t[56554] = t[56553] ^ n[56554];
assign t[56555] = t[56554] ^ n[56555];
assign t[56556] = t[56555] ^ n[56556];
assign t[56557] = t[56556] ^ n[56557];
assign t[56558] = t[56557] ^ n[56558];
assign t[56559] = t[56558] ^ n[56559];
assign t[56560] = t[56559] ^ n[56560];
assign t[56561] = t[56560] ^ n[56561];
assign t[56562] = t[56561] ^ n[56562];
assign t[56563] = t[56562] ^ n[56563];
assign t[56564] = t[56563] ^ n[56564];
assign t[56565] = t[56564] ^ n[56565];
assign t[56566] = t[56565] ^ n[56566];
assign t[56567] = t[56566] ^ n[56567];
assign t[56568] = t[56567] ^ n[56568];
assign t[56569] = t[56568] ^ n[56569];
assign t[56570] = t[56569] ^ n[56570];
assign t[56571] = t[56570] ^ n[56571];
assign t[56572] = t[56571] ^ n[56572];
assign t[56573] = t[56572] ^ n[56573];
assign t[56574] = t[56573] ^ n[56574];
assign t[56575] = t[56574] ^ n[56575];
assign t[56576] = t[56575] ^ n[56576];
assign t[56577] = t[56576] ^ n[56577];
assign t[56578] = t[56577] ^ n[56578];
assign t[56579] = t[56578] ^ n[56579];
assign t[56580] = t[56579] ^ n[56580];
assign t[56581] = t[56580] ^ n[56581];
assign t[56582] = t[56581] ^ n[56582];
assign t[56583] = t[56582] ^ n[56583];
assign t[56584] = t[56583] ^ n[56584];
assign t[56585] = t[56584] ^ n[56585];
assign t[56586] = t[56585] ^ n[56586];
assign t[56587] = t[56586] ^ n[56587];
assign t[56588] = t[56587] ^ n[56588];
assign t[56589] = t[56588] ^ n[56589];
assign t[56590] = t[56589] ^ n[56590];
assign t[56591] = t[56590] ^ n[56591];
assign t[56592] = t[56591] ^ n[56592];
assign t[56593] = t[56592] ^ n[56593];
assign t[56594] = t[56593] ^ n[56594];
assign t[56595] = t[56594] ^ n[56595];
assign t[56596] = t[56595] ^ n[56596];
assign t[56597] = t[56596] ^ n[56597];
assign t[56598] = t[56597] ^ n[56598];
assign t[56599] = t[56598] ^ n[56599];
assign t[56600] = t[56599] ^ n[56600];
assign t[56601] = t[56600] ^ n[56601];
assign t[56602] = t[56601] ^ n[56602];
assign t[56603] = t[56602] ^ n[56603];
assign t[56604] = t[56603] ^ n[56604];
assign t[56605] = t[56604] ^ n[56605];
assign t[56606] = t[56605] ^ n[56606];
assign t[56607] = t[56606] ^ n[56607];
assign t[56608] = t[56607] ^ n[56608];
assign t[56609] = t[56608] ^ n[56609];
assign t[56610] = t[56609] ^ n[56610];
assign t[56611] = t[56610] ^ n[56611];
assign t[56612] = t[56611] ^ n[56612];
assign t[56613] = t[56612] ^ n[56613];
assign t[56614] = t[56613] ^ n[56614];
assign t[56615] = t[56614] ^ n[56615];
assign t[56616] = t[56615] ^ n[56616];
assign t[56617] = t[56616] ^ n[56617];
assign t[56618] = t[56617] ^ n[56618];
assign t[56619] = t[56618] ^ n[56619];
assign t[56620] = t[56619] ^ n[56620];
assign t[56621] = t[56620] ^ n[56621];
assign t[56622] = t[56621] ^ n[56622];
assign t[56623] = t[56622] ^ n[56623];
assign t[56624] = t[56623] ^ n[56624];
assign t[56625] = t[56624] ^ n[56625];
assign t[56626] = t[56625] ^ n[56626];
assign t[56627] = t[56626] ^ n[56627];
assign t[56628] = t[56627] ^ n[56628];
assign t[56629] = t[56628] ^ n[56629];
assign t[56630] = t[56629] ^ n[56630];
assign t[56631] = t[56630] ^ n[56631];
assign t[56632] = t[56631] ^ n[56632];
assign t[56633] = t[56632] ^ n[56633];
assign t[56634] = t[56633] ^ n[56634];
assign t[56635] = t[56634] ^ n[56635];
assign t[56636] = t[56635] ^ n[56636];
assign t[56637] = t[56636] ^ n[56637];
assign t[56638] = t[56637] ^ n[56638];
assign t[56639] = t[56638] ^ n[56639];
assign t[56640] = t[56639] ^ n[56640];
assign t[56641] = t[56640] ^ n[56641];
assign t[56642] = t[56641] ^ n[56642];
assign t[56643] = t[56642] ^ n[56643];
assign t[56644] = t[56643] ^ n[56644];
assign t[56645] = t[56644] ^ n[56645];
assign t[56646] = t[56645] ^ n[56646];
assign t[56647] = t[56646] ^ n[56647];
assign t[56648] = t[56647] ^ n[56648];
assign t[56649] = t[56648] ^ n[56649];
assign t[56650] = t[56649] ^ n[56650];
assign t[56651] = t[56650] ^ n[56651];
assign t[56652] = t[56651] ^ n[56652];
assign t[56653] = t[56652] ^ n[56653];
assign t[56654] = t[56653] ^ n[56654];
assign t[56655] = t[56654] ^ n[56655];
assign t[56656] = t[56655] ^ n[56656];
assign t[56657] = t[56656] ^ n[56657];
assign t[56658] = t[56657] ^ n[56658];
assign t[56659] = t[56658] ^ n[56659];
assign t[56660] = t[56659] ^ n[56660];
assign t[56661] = t[56660] ^ n[56661];
assign t[56662] = t[56661] ^ n[56662];
assign t[56663] = t[56662] ^ n[56663];
assign t[56664] = t[56663] ^ n[56664];
assign t[56665] = t[56664] ^ n[56665];
assign t[56666] = t[56665] ^ n[56666];
assign t[56667] = t[56666] ^ n[56667];
assign t[56668] = t[56667] ^ n[56668];
assign t[56669] = t[56668] ^ n[56669];
assign t[56670] = t[56669] ^ n[56670];
assign t[56671] = t[56670] ^ n[56671];
assign t[56672] = t[56671] ^ n[56672];
assign t[56673] = t[56672] ^ n[56673];
assign t[56674] = t[56673] ^ n[56674];
assign t[56675] = t[56674] ^ n[56675];
assign t[56676] = t[56675] ^ n[56676];
assign t[56677] = t[56676] ^ n[56677];
assign t[56678] = t[56677] ^ n[56678];
assign t[56679] = t[56678] ^ n[56679];
assign t[56680] = t[56679] ^ n[56680];
assign t[56681] = t[56680] ^ n[56681];
assign t[56682] = t[56681] ^ n[56682];
assign t[56683] = t[56682] ^ n[56683];
assign t[56684] = t[56683] ^ n[56684];
assign t[56685] = t[56684] ^ n[56685];
assign t[56686] = t[56685] ^ n[56686];
assign t[56687] = t[56686] ^ n[56687];
assign t[56688] = t[56687] ^ n[56688];
assign t[56689] = t[56688] ^ n[56689];
assign t[56690] = t[56689] ^ n[56690];
assign t[56691] = t[56690] ^ n[56691];
assign t[56692] = t[56691] ^ n[56692];
assign t[56693] = t[56692] ^ n[56693];
assign t[56694] = t[56693] ^ n[56694];
assign t[56695] = t[56694] ^ n[56695];
assign t[56696] = t[56695] ^ n[56696];
assign t[56697] = t[56696] ^ n[56697];
assign t[56698] = t[56697] ^ n[56698];
assign t[56699] = t[56698] ^ n[56699];
assign t[56700] = t[56699] ^ n[56700];
assign t[56701] = t[56700] ^ n[56701];
assign t[56702] = t[56701] ^ n[56702];
assign t[56703] = t[56702] ^ n[56703];
assign t[56704] = t[56703] ^ n[56704];
assign t[56705] = t[56704] ^ n[56705];
assign t[56706] = t[56705] ^ n[56706];
assign t[56707] = t[56706] ^ n[56707];
assign t[56708] = t[56707] ^ n[56708];
assign t[56709] = t[56708] ^ n[56709];
assign t[56710] = t[56709] ^ n[56710];
assign t[56711] = t[56710] ^ n[56711];
assign t[56712] = t[56711] ^ n[56712];
assign t[56713] = t[56712] ^ n[56713];
assign t[56714] = t[56713] ^ n[56714];
assign t[56715] = t[56714] ^ n[56715];
assign t[56716] = t[56715] ^ n[56716];
assign t[56717] = t[56716] ^ n[56717];
assign t[56718] = t[56717] ^ n[56718];
assign t[56719] = t[56718] ^ n[56719];
assign t[56720] = t[56719] ^ n[56720];
assign t[56721] = t[56720] ^ n[56721];
assign t[56722] = t[56721] ^ n[56722];
assign t[56723] = t[56722] ^ n[56723];
assign t[56724] = t[56723] ^ n[56724];
assign t[56725] = t[56724] ^ n[56725];
assign t[56726] = t[56725] ^ n[56726];
assign t[56727] = t[56726] ^ n[56727];
assign t[56728] = t[56727] ^ n[56728];
assign t[56729] = t[56728] ^ n[56729];
assign t[56730] = t[56729] ^ n[56730];
assign t[56731] = t[56730] ^ n[56731];
assign t[56732] = t[56731] ^ n[56732];
assign t[56733] = t[56732] ^ n[56733];
assign t[56734] = t[56733] ^ n[56734];
assign t[56735] = t[56734] ^ n[56735];
assign t[56736] = t[56735] ^ n[56736];
assign t[56737] = t[56736] ^ n[56737];
assign t[56738] = t[56737] ^ n[56738];
assign t[56739] = t[56738] ^ n[56739];
assign t[56740] = t[56739] ^ n[56740];
assign t[56741] = t[56740] ^ n[56741];
assign t[56742] = t[56741] ^ n[56742];
assign t[56743] = t[56742] ^ n[56743];
assign t[56744] = t[56743] ^ n[56744];
assign t[56745] = t[56744] ^ n[56745];
assign t[56746] = t[56745] ^ n[56746];
assign t[56747] = t[56746] ^ n[56747];
assign t[56748] = t[56747] ^ n[56748];
assign t[56749] = t[56748] ^ n[56749];
assign t[56750] = t[56749] ^ n[56750];
assign t[56751] = t[56750] ^ n[56751];
assign t[56752] = t[56751] ^ n[56752];
assign t[56753] = t[56752] ^ n[56753];
assign t[56754] = t[56753] ^ n[56754];
assign t[56755] = t[56754] ^ n[56755];
assign t[56756] = t[56755] ^ n[56756];
assign t[56757] = t[56756] ^ n[56757];
assign t[56758] = t[56757] ^ n[56758];
assign t[56759] = t[56758] ^ n[56759];
assign t[56760] = t[56759] ^ n[56760];
assign t[56761] = t[56760] ^ n[56761];
assign t[56762] = t[56761] ^ n[56762];
assign t[56763] = t[56762] ^ n[56763];
assign t[56764] = t[56763] ^ n[56764];
assign t[56765] = t[56764] ^ n[56765];
assign t[56766] = t[56765] ^ n[56766];
assign t[56767] = t[56766] ^ n[56767];
assign t[56768] = t[56767] ^ n[56768];
assign t[56769] = t[56768] ^ n[56769];
assign t[56770] = t[56769] ^ n[56770];
assign t[56771] = t[56770] ^ n[56771];
assign t[56772] = t[56771] ^ n[56772];
assign t[56773] = t[56772] ^ n[56773];
assign t[56774] = t[56773] ^ n[56774];
assign t[56775] = t[56774] ^ n[56775];
assign t[56776] = t[56775] ^ n[56776];
assign t[56777] = t[56776] ^ n[56777];
assign t[56778] = t[56777] ^ n[56778];
assign t[56779] = t[56778] ^ n[56779];
assign t[56780] = t[56779] ^ n[56780];
assign t[56781] = t[56780] ^ n[56781];
assign t[56782] = t[56781] ^ n[56782];
assign t[56783] = t[56782] ^ n[56783];
assign t[56784] = t[56783] ^ n[56784];
assign t[56785] = t[56784] ^ n[56785];
assign t[56786] = t[56785] ^ n[56786];
assign t[56787] = t[56786] ^ n[56787];
assign t[56788] = t[56787] ^ n[56788];
assign t[56789] = t[56788] ^ n[56789];
assign t[56790] = t[56789] ^ n[56790];
assign t[56791] = t[56790] ^ n[56791];
assign t[56792] = t[56791] ^ n[56792];
assign t[56793] = t[56792] ^ n[56793];
assign t[56794] = t[56793] ^ n[56794];
assign t[56795] = t[56794] ^ n[56795];
assign t[56796] = t[56795] ^ n[56796];
assign t[56797] = t[56796] ^ n[56797];
assign t[56798] = t[56797] ^ n[56798];
assign t[56799] = t[56798] ^ n[56799];
assign t[56800] = t[56799] ^ n[56800];
assign t[56801] = t[56800] ^ n[56801];
assign t[56802] = t[56801] ^ n[56802];
assign t[56803] = t[56802] ^ n[56803];
assign t[56804] = t[56803] ^ n[56804];
assign t[56805] = t[56804] ^ n[56805];
assign t[56806] = t[56805] ^ n[56806];
assign t[56807] = t[56806] ^ n[56807];
assign t[56808] = t[56807] ^ n[56808];
assign t[56809] = t[56808] ^ n[56809];
assign t[56810] = t[56809] ^ n[56810];
assign t[56811] = t[56810] ^ n[56811];
assign t[56812] = t[56811] ^ n[56812];
assign t[56813] = t[56812] ^ n[56813];
assign t[56814] = t[56813] ^ n[56814];
assign t[56815] = t[56814] ^ n[56815];
assign t[56816] = t[56815] ^ n[56816];
assign t[56817] = t[56816] ^ n[56817];
assign t[56818] = t[56817] ^ n[56818];
assign t[56819] = t[56818] ^ n[56819];
assign t[56820] = t[56819] ^ n[56820];
assign t[56821] = t[56820] ^ n[56821];
assign t[56822] = t[56821] ^ n[56822];
assign t[56823] = t[56822] ^ n[56823];
assign t[56824] = t[56823] ^ n[56824];
assign t[56825] = t[56824] ^ n[56825];
assign t[56826] = t[56825] ^ n[56826];
assign t[56827] = t[56826] ^ n[56827];
assign t[56828] = t[56827] ^ n[56828];
assign t[56829] = t[56828] ^ n[56829];
assign t[56830] = t[56829] ^ n[56830];
assign t[56831] = t[56830] ^ n[56831];
assign t[56832] = t[56831] ^ n[56832];
assign t[56833] = t[56832] ^ n[56833];
assign t[56834] = t[56833] ^ n[56834];
assign t[56835] = t[56834] ^ n[56835];
assign t[56836] = t[56835] ^ n[56836];
assign t[56837] = t[56836] ^ n[56837];
assign t[56838] = t[56837] ^ n[56838];
assign t[56839] = t[56838] ^ n[56839];
assign t[56840] = t[56839] ^ n[56840];
assign t[56841] = t[56840] ^ n[56841];
assign t[56842] = t[56841] ^ n[56842];
assign t[56843] = t[56842] ^ n[56843];
assign t[56844] = t[56843] ^ n[56844];
assign t[56845] = t[56844] ^ n[56845];
assign t[56846] = t[56845] ^ n[56846];
assign t[56847] = t[56846] ^ n[56847];
assign t[56848] = t[56847] ^ n[56848];
assign t[56849] = t[56848] ^ n[56849];
assign t[56850] = t[56849] ^ n[56850];
assign t[56851] = t[56850] ^ n[56851];
assign t[56852] = t[56851] ^ n[56852];
assign t[56853] = t[56852] ^ n[56853];
assign t[56854] = t[56853] ^ n[56854];
assign t[56855] = t[56854] ^ n[56855];
assign t[56856] = t[56855] ^ n[56856];
assign t[56857] = t[56856] ^ n[56857];
assign t[56858] = t[56857] ^ n[56858];
assign t[56859] = t[56858] ^ n[56859];
assign t[56860] = t[56859] ^ n[56860];
assign t[56861] = t[56860] ^ n[56861];
assign t[56862] = t[56861] ^ n[56862];
assign t[56863] = t[56862] ^ n[56863];
assign t[56864] = t[56863] ^ n[56864];
assign t[56865] = t[56864] ^ n[56865];
assign t[56866] = t[56865] ^ n[56866];
assign t[56867] = t[56866] ^ n[56867];
assign t[56868] = t[56867] ^ n[56868];
assign t[56869] = t[56868] ^ n[56869];
assign t[56870] = t[56869] ^ n[56870];
assign t[56871] = t[56870] ^ n[56871];
assign t[56872] = t[56871] ^ n[56872];
assign t[56873] = t[56872] ^ n[56873];
assign t[56874] = t[56873] ^ n[56874];
assign t[56875] = t[56874] ^ n[56875];
assign t[56876] = t[56875] ^ n[56876];
assign t[56877] = t[56876] ^ n[56877];
assign t[56878] = t[56877] ^ n[56878];
assign t[56879] = t[56878] ^ n[56879];
assign t[56880] = t[56879] ^ n[56880];
assign t[56881] = t[56880] ^ n[56881];
assign t[56882] = t[56881] ^ n[56882];
assign t[56883] = t[56882] ^ n[56883];
assign t[56884] = t[56883] ^ n[56884];
assign t[56885] = t[56884] ^ n[56885];
assign t[56886] = t[56885] ^ n[56886];
assign t[56887] = t[56886] ^ n[56887];
assign t[56888] = t[56887] ^ n[56888];
assign t[56889] = t[56888] ^ n[56889];
assign t[56890] = t[56889] ^ n[56890];
assign t[56891] = t[56890] ^ n[56891];
assign t[56892] = t[56891] ^ n[56892];
assign t[56893] = t[56892] ^ n[56893];
assign t[56894] = t[56893] ^ n[56894];
assign t[56895] = t[56894] ^ n[56895];
assign t[56896] = t[56895] ^ n[56896];
assign t[56897] = t[56896] ^ n[56897];
assign t[56898] = t[56897] ^ n[56898];
assign t[56899] = t[56898] ^ n[56899];
assign t[56900] = t[56899] ^ n[56900];
assign t[56901] = t[56900] ^ n[56901];
assign t[56902] = t[56901] ^ n[56902];
assign t[56903] = t[56902] ^ n[56903];
assign t[56904] = t[56903] ^ n[56904];
assign t[56905] = t[56904] ^ n[56905];
assign t[56906] = t[56905] ^ n[56906];
assign t[56907] = t[56906] ^ n[56907];
assign t[56908] = t[56907] ^ n[56908];
assign t[56909] = t[56908] ^ n[56909];
assign t[56910] = t[56909] ^ n[56910];
assign t[56911] = t[56910] ^ n[56911];
assign t[56912] = t[56911] ^ n[56912];
assign t[56913] = t[56912] ^ n[56913];
assign t[56914] = t[56913] ^ n[56914];
assign t[56915] = t[56914] ^ n[56915];
assign t[56916] = t[56915] ^ n[56916];
assign t[56917] = t[56916] ^ n[56917];
assign t[56918] = t[56917] ^ n[56918];
assign t[56919] = t[56918] ^ n[56919];
assign t[56920] = t[56919] ^ n[56920];
assign t[56921] = t[56920] ^ n[56921];
assign t[56922] = t[56921] ^ n[56922];
assign t[56923] = t[56922] ^ n[56923];
assign t[56924] = t[56923] ^ n[56924];
assign t[56925] = t[56924] ^ n[56925];
assign t[56926] = t[56925] ^ n[56926];
assign t[56927] = t[56926] ^ n[56927];
assign t[56928] = t[56927] ^ n[56928];
assign t[56929] = t[56928] ^ n[56929];
assign t[56930] = t[56929] ^ n[56930];
assign t[56931] = t[56930] ^ n[56931];
assign t[56932] = t[56931] ^ n[56932];
assign t[56933] = t[56932] ^ n[56933];
assign t[56934] = t[56933] ^ n[56934];
assign t[56935] = t[56934] ^ n[56935];
assign t[56936] = t[56935] ^ n[56936];
assign t[56937] = t[56936] ^ n[56937];
assign t[56938] = t[56937] ^ n[56938];
assign t[56939] = t[56938] ^ n[56939];
assign t[56940] = t[56939] ^ n[56940];
assign t[56941] = t[56940] ^ n[56941];
assign t[56942] = t[56941] ^ n[56942];
assign t[56943] = t[56942] ^ n[56943];
assign t[56944] = t[56943] ^ n[56944];
assign t[56945] = t[56944] ^ n[56945];
assign t[56946] = t[56945] ^ n[56946];
assign t[56947] = t[56946] ^ n[56947];
assign t[56948] = t[56947] ^ n[56948];
assign t[56949] = t[56948] ^ n[56949];
assign t[56950] = t[56949] ^ n[56950];
assign t[56951] = t[56950] ^ n[56951];
assign t[56952] = t[56951] ^ n[56952];
assign t[56953] = t[56952] ^ n[56953];
assign t[56954] = t[56953] ^ n[56954];
assign t[56955] = t[56954] ^ n[56955];
assign t[56956] = t[56955] ^ n[56956];
assign t[56957] = t[56956] ^ n[56957];
assign t[56958] = t[56957] ^ n[56958];
assign t[56959] = t[56958] ^ n[56959];
assign t[56960] = t[56959] ^ n[56960];
assign t[56961] = t[56960] ^ n[56961];
assign t[56962] = t[56961] ^ n[56962];
assign t[56963] = t[56962] ^ n[56963];
assign t[56964] = t[56963] ^ n[56964];
assign t[56965] = t[56964] ^ n[56965];
assign t[56966] = t[56965] ^ n[56966];
assign t[56967] = t[56966] ^ n[56967];
assign t[56968] = t[56967] ^ n[56968];
assign t[56969] = t[56968] ^ n[56969];
assign t[56970] = t[56969] ^ n[56970];
assign t[56971] = t[56970] ^ n[56971];
assign t[56972] = t[56971] ^ n[56972];
assign t[56973] = t[56972] ^ n[56973];
assign t[56974] = t[56973] ^ n[56974];
assign t[56975] = t[56974] ^ n[56975];
assign t[56976] = t[56975] ^ n[56976];
assign t[56977] = t[56976] ^ n[56977];
assign t[56978] = t[56977] ^ n[56978];
assign t[56979] = t[56978] ^ n[56979];
assign t[56980] = t[56979] ^ n[56980];
assign t[56981] = t[56980] ^ n[56981];
assign t[56982] = t[56981] ^ n[56982];
assign t[56983] = t[56982] ^ n[56983];
assign t[56984] = t[56983] ^ n[56984];
assign t[56985] = t[56984] ^ n[56985];
assign t[56986] = t[56985] ^ n[56986];
assign t[56987] = t[56986] ^ n[56987];
assign t[56988] = t[56987] ^ n[56988];
assign t[56989] = t[56988] ^ n[56989];
assign t[56990] = t[56989] ^ n[56990];
assign t[56991] = t[56990] ^ n[56991];
assign t[56992] = t[56991] ^ n[56992];
assign t[56993] = t[56992] ^ n[56993];
assign t[56994] = t[56993] ^ n[56994];
assign t[56995] = t[56994] ^ n[56995];
assign t[56996] = t[56995] ^ n[56996];
assign t[56997] = t[56996] ^ n[56997];
assign t[56998] = t[56997] ^ n[56998];
assign t[56999] = t[56998] ^ n[56999];
assign t[57000] = t[56999] ^ n[57000];
assign t[57001] = t[57000] ^ n[57001];
assign t[57002] = t[57001] ^ n[57002];
assign t[57003] = t[57002] ^ n[57003];
assign t[57004] = t[57003] ^ n[57004];
assign t[57005] = t[57004] ^ n[57005];
assign t[57006] = t[57005] ^ n[57006];
assign t[57007] = t[57006] ^ n[57007];
assign t[57008] = t[57007] ^ n[57008];
assign t[57009] = t[57008] ^ n[57009];
assign t[57010] = t[57009] ^ n[57010];
assign t[57011] = t[57010] ^ n[57011];
assign t[57012] = t[57011] ^ n[57012];
assign t[57013] = t[57012] ^ n[57013];
assign t[57014] = t[57013] ^ n[57014];
assign t[57015] = t[57014] ^ n[57015];
assign t[57016] = t[57015] ^ n[57016];
assign t[57017] = t[57016] ^ n[57017];
assign t[57018] = t[57017] ^ n[57018];
assign t[57019] = t[57018] ^ n[57019];
assign t[57020] = t[57019] ^ n[57020];
assign t[57021] = t[57020] ^ n[57021];
assign t[57022] = t[57021] ^ n[57022];
assign t[57023] = t[57022] ^ n[57023];
assign t[57024] = t[57023] ^ n[57024];
assign t[57025] = t[57024] ^ n[57025];
assign t[57026] = t[57025] ^ n[57026];
assign t[57027] = t[57026] ^ n[57027];
assign t[57028] = t[57027] ^ n[57028];
assign t[57029] = t[57028] ^ n[57029];
assign t[57030] = t[57029] ^ n[57030];
assign t[57031] = t[57030] ^ n[57031];
assign t[57032] = t[57031] ^ n[57032];
assign t[57033] = t[57032] ^ n[57033];
assign t[57034] = t[57033] ^ n[57034];
assign t[57035] = t[57034] ^ n[57035];
assign t[57036] = t[57035] ^ n[57036];
assign t[57037] = t[57036] ^ n[57037];
assign t[57038] = t[57037] ^ n[57038];
assign t[57039] = t[57038] ^ n[57039];
assign t[57040] = t[57039] ^ n[57040];
assign t[57041] = t[57040] ^ n[57041];
assign t[57042] = t[57041] ^ n[57042];
assign t[57043] = t[57042] ^ n[57043];
assign t[57044] = t[57043] ^ n[57044];
assign t[57045] = t[57044] ^ n[57045];
assign t[57046] = t[57045] ^ n[57046];
assign t[57047] = t[57046] ^ n[57047];
assign t[57048] = t[57047] ^ n[57048];
assign t[57049] = t[57048] ^ n[57049];
assign t[57050] = t[57049] ^ n[57050];
assign t[57051] = t[57050] ^ n[57051];
assign t[57052] = t[57051] ^ n[57052];
assign t[57053] = t[57052] ^ n[57053];
assign t[57054] = t[57053] ^ n[57054];
assign t[57055] = t[57054] ^ n[57055];
assign t[57056] = t[57055] ^ n[57056];
assign t[57057] = t[57056] ^ n[57057];
assign t[57058] = t[57057] ^ n[57058];
assign t[57059] = t[57058] ^ n[57059];
assign t[57060] = t[57059] ^ n[57060];
assign t[57061] = t[57060] ^ n[57061];
assign t[57062] = t[57061] ^ n[57062];
assign t[57063] = t[57062] ^ n[57063];
assign t[57064] = t[57063] ^ n[57064];
assign t[57065] = t[57064] ^ n[57065];
assign t[57066] = t[57065] ^ n[57066];
assign t[57067] = t[57066] ^ n[57067];
assign t[57068] = t[57067] ^ n[57068];
assign t[57069] = t[57068] ^ n[57069];
assign t[57070] = t[57069] ^ n[57070];
assign t[57071] = t[57070] ^ n[57071];
assign t[57072] = t[57071] ^ n[57072];
assign t[57073] = t[57072] ^ n[57073];
assign t[57074] = t[57073] ^ n[57074];
assign t[57075] = t[57074] ^ n[57075];
assign t[57076] = t[57075] ^ n[57076];
assign t[57077] = t[57076] ^ n[57077];
assign t[57078] = t[57077] ^ n[57078];
assign t[57079] = t[57078] ^ n[57079];
assign t[57080] = t[57079] ^ n[57080];
assign t[57081] = t[57080] ^ n[57081];
assign t[57082] = t[57081] ^ n[57082];
assign t[57083] = t[57082] ^ n[57083];
assign t[57084] = t[57083] ^ n[57084];
assign t[57085] = t[57084] ^ n[57085];
assign t[57086] = t[57085] ^ n[57086];
assign t[57087] = t[57086] ^ n[57087];
assign t[57088] = t[57087] ^ n[57088];
assign t[57089] = t[57088] ^ n[57089];
assign t[57090] = t[57089] ^ n[57090];
assign t[57091] = t[57090] ^ n[57091];
assign t[57092] = t[57091] ^ n[57092];
assign t[57093] = t[57092] ^ n[57093];
assign t[57094] = t[57093] ^ n[57094];
assign t[57095] = t[57094] ^ n[57095];
assign t[57096] = t[57095] ^ n[57096];
assign t[57097] = t[57096] ^ n[57097];
assign t[57098] = t[57097] ^ n[57098];
assign t[57099] = t[57098] ^ n[57099];
assign t[57100] = t[57099] ^ n[57100];
assign t[57101] = t[57100] ^ n[57101];
assign t[57102] = t[57101] ^ n[57102];
assign t[57103] = t[57102] ^ n[57103];
assign t[57104] = t[57103] ^ n[57104];
assign t[57105] = t[57104] ^ n[57105];
assign t[57106] = t[57105] ^ n[57106];
assign t[57107] = t[57106] ^ n[57107];
assign t[57108] = t[57107] ^ n[57108];
assign t[57109] = t[57108] ^ n[57109];
assign t[57110] = t[57109] ^ n[57110];
assign t[57111] = t[57110] ^ n[57111];
assign t[57112] = t[57111] ^ n[57112];
assign t[57113] = t[57112] ^ n[57113];
assign t[57114] = t[57113] ^ n[57114];
assign t[57115] = t[57114] ^ n[57115];
assign t[57116] = t[57115] ^ n[57116];
assign t[57117] = t[57116] ^ n[57117];
assign t[57118] = t[57117] ^ n[57118];
assign t[57119] = t[57118] ^ n[57119];
assign t[57120] = t[57119] ^ n[57120];
assign t[57121] = t[57120] ^ n[57121];
assign t[57122] = t[57121] ^ n[57122];
assign t[57123] = t[57122] ^ n[57123];
assign t[57124] = t[57123] ^ n[57124];
assign t[57125] = t[57124] ^ n[57125];
assign t[57126] = t[57125] ^ n[57126];
assign t[57127] = t[57126] ^ n[57127];
assign t[57128] = t[57127] ^ n[57128];
assign t[57129] = t[57128] ^ n[57129];
assign t[57130] = t[57129] ^ n[57130];
assign t[57131] = t[57130] ^ n[57131];
assign t[57132] = t[57131] ^ n[57132];
assign t[57133] = t[57132] ^ n[57133];
assign t[57134] = t[57133] ^ n[57134];
assign t[57135] = t[57134] ^ n[57135];
assign t[57136] = t[57135] ^ n[57136];
assign t[57137] = t[57136] ^ n[57137];
assign t[57138] = t[57137] ^ n[57138];
assign t[57139] = t[57138] ^ n[57139];
assign t[57140] = t[57139] ^ n[57140];
assign t[57141] = t[57140] ^ n[57141];
assign t[57142] = t[57141] ^ n[57142];
assign t[57143] = t[57142] ^ n[57143];
assign t[57144] = t[57143] ^ n[57144];
assign t[57145] = t[57144] ^ n[57145];
assign t[57146] = t[57145] ^ n[57146];
assign t[57147] = t[57146] ^ n[57147];
assign t[57148] = t[57147] ^ n[57148];
assign t[57149] = t[57148] ^ n[57149];
assign t[57150] = t[57149] ^ n[57150];
assign t[57151] = t[57150] ^ n[57151];
assign t[57152] = t[57151] ^ n[57152];
assign t[57153] = t[57152] ^ n[57153];
assign t[57154] = t[57153] ^ n[57154];
assign t[57155] = t[57154] ^ n[57155];
assign t[57156] = t[57155] ^ n[57156];
assign t[57157] = t[57156] ^ n[57157];
assign t[57158] = t[57157] ^ n[57158];
assign t[57159] = t[57158] ^ n[57159];
assign t[57160] = t[57159] ^ n[57160];
assign t[57161] = t[57160] ^ n[57161];
assign t[57162] = t[57161] ^ n[57162];
assign t[57163] = t[57162] ^ n[57163];
assign t[57164] = t[57163] ^ n[57164];
assign t[57165] = t[57164] ^ n[57165];
assign t[57166] = t[57165] ^ n[57166];
assign t[57167] = t[57166] ^ n[57167];
assign t[57168] = t[57167] ^ n[57168];
assign t[57169] = t[57168] ^ n[57169];
assign t[57170] = t[57169] ^ n[57170];
assign t[57171] = t[57170] ^ n[57171];
assign t[57172] = t[57171] ^ n[57172];
assign t[57173] = t[57172] ^ n[57173];
assign t[57174] = t[57173] ^ n[57174];
assign t[57175] = t[57174] ^ n[57175];
assign t[57176] = t[57175] ^ n[57176];
assign t[57177] = t[57176] ^ n[57177];
assign t[57178] = t[57177] ^ n[57178];
assign t[57179] = t[57178] ^ n[57179];
assign t[57180] = t[57179] ^ n[57180];
assign t[57181] = t[57180] ^ n[57181];
assign t[57182] = t[57181] ^ n[57182];
assign t[57183] = t[57182] ^ n[57183];
assign t[57184] = t[57183] ^ n[57184];
assign t[57185] = t[57184] ^ n[57185];
assign t[57186] = t[57185] ^ n[57186];
assign t[57187] = t[57186] ^ n[57187];
assign t[57188] = t[57187] ^ n[57188];
assign t[57189] = t[57188] ^ n[57189];
assign t[57190] = t[57189] ^ n[57190];
assign t[57191] = t[57190] ^ n[57191];
assign t[57192] = t[57191] ^ n[57192];
assign t[57193] = t[57192] ^ n[57193];
assign t[57194] = t[57193] ^ n[57194];
assign t[57195] = t[57194] ^ n[57195];
assign t[57196] = t[57195] ^ n[57196];
assign t[57197] = t[57196] ^ n[57197];
assign t[57198] = t[57197] ^ n[57198];
assign t[57199] = t[57198] ^ n[57199];
assign t[57200] = t[57199] ^ n[57200];
assign t[57201] = t[57200] ^ n[57201];
assign t[57202] = t[57201] ^ n[57202];
assign t[57203] = t[57202] ^ n[57203];
assign t[57204] = t[57203] ^ n[57204];
assign t[57205] = t[57204] ^ n[57205];
assign t[57206] = t[57205] ^ n[57206];
assign t[57207] = t[57206] ^ n[57207];
assign t[57208] = t[57207] ^ n[57208];
assign t[57209] = t[57208] ^ n[57209];
assign t[57210] = t[57209] ^ n[57210];
assign t[57211] = t[57210] ^ n[57211];
assign t[57212] = t[57211] ^ n[57212];
assign t[57213] = t[57212] ^ n[57213];
assign t[57214] = t[57213] ^ n[57214];
assign t[57215] = t[57214] ^ n[57215];
assign t[57216] = t[57215] ^ n[57216];
assign t[57217] = t[57216] ^ n[57217];
assign t[57218] = t[57217] ^ n[57218];
assign t[57219] = t[57218] ^ n[57219];
assign t[57220] = t[57219] ^ n[57220];
assign t[57221] = t[57220] ^ n[57221];
assign t[57222] = t[57221] ^ n[57222];
assign t[57223] = t[57222] ^ n[57223];
assign t[57224] = t[57223] ^ n[57224];
assign t[57225] = t[57224] ^ n[57225];
assign t[57226] = t[57225] ^ n[57226];
assign t[57227] = t[57226] ^ n[57227];
assign t[57228] = t[57227] ^ n[57228];
assign t[57229] = t[57228] ^ n[57229];
assign t[57230] = t[57229] ^ n[57230];
assign t[57231] = t[57230] ^ n[57231];
assign t[57232] = t[57231] ^ n[57232];
assign t[57233] = t[57232] ^ n[57233];
assign t[57234] = t[57233] ^ n[57234];
assign t[57235] = t[57234] ^ n[57235];
assign t[57236] = t[57235] ^ n[57236];
assign t[57237] = t[57236] ^ n[57237];
assign t[57238] = t[57237] ^ n[57238];
assign t[57239] = t[57238] ^ n[57239];
assign t[57240] = t[57239] ^ n[57240];
assign t[57241] = t[57240] ^ n[57241];
assign t[57242] = t[57241] ^ n[57242];
assign t[57243] = t[57242] ^ n[57243];
assign t[57244] = t[57243] ^ n[57244];
assign t[57245] = t[57244] ^ n[57245];
assign t[57246] = t[57245] ^ n[57246];
assign t[57247] = t[57246] ^ n[57247];
assign t[57248] = t[57247] ^ n[57248];
assign t[57249] = t[57248] ^ n[57249];
assign t[57250] = t[57249] ^ n[57250];
assign t[57251] = t[57250] ^ n[57251];
assign t[57252] = t[57251] ^ n[57252];
assign t[57253] = t[57252] ^ n[57253];
assign t[57254] = t[57253] ^ n[57254];
assign t[57255] = t[57254] ^ n[57255];
assign t[57256] = t[57255] ^ n[57256];
assign t[57257] = t[57256] ^ n[57257];
assign t[57258] = t[57257] ^ n[57258];
assign t[57259] = t[57258] ^ n[57259];
assign t[57260] = t[57259] ^ n[57260];
assign t[57261] = t[57260] ^ n[57261];
assign t[57262] = t[57261] ^ n[57262];
assign t[57263] = t[57262] ^ n[57263];
assign t[57264] = t[57263] ^ n[57264];
assign t[57265] = t[57264] ^ n[57265];
assign t[57266] = t[57265] ^ n[57266];
assign t[57267] = t[57266] ^ n[57267];
assign t[57268] = t[57267] ^ n[57268];
assign t[57269] = t[57268] ^ n[57269];
assign t[57270] = t[57269] ^ n[57270];
assign t[57271] = t[57270] ^ n[57271];
assign t[57272] = t[57271] ^ n[57272];
assign t[57273] = t[57272] ^ n[57273];
assign t[57274] = t[57273] ^ n[57274];
assign t[57275] = t[57274] ^ n[57275];
assign t[57276] = t[57275] ^ n[57276];
assign t[57277] = t[57276] ^ n[57277];
assign t[57278] = t[57277] ^ n[57278];
assign t[57279] = t[57278] ^ n[57279];
assign t[57280] = t[57279] ^ n[57280];
assign t[57281] = t[57280] ^ n[57281];
assign t[57282] = t[57281] ^ n[57282];
assign t[57283] = t[57282] ^ n[57283];
assign t[57284] = t[57283] ^ n[57284];
assign t[57285] = t[57284] ^ n[57285];
assign t[57286] = t[57285] ^ n[57286];
assign t[57287] = t[57286] ^ n[57287];
assign t[57288] = t[57287] ^ n[57288];
assign t[57289] = t[57288] ^ n[57289];
assign t[57290] = t[57289] ^ n[57290];
assign t[57291] = t[57290] ^ n[57291];
assign t[57292] = t[57291] ^ n[57292];
assign t[57293] = t[57292] ^ n[57293];
assign t[57294] = t[57293] ^ n[57294];
assign t[57295] = t[57294] ^ n[57295];
assign t[57296] = t[57295] ^ n[57296];
assign t[57297] = t[57296] ^ n[57297];
assign t[57298] = t[57297] ^ n[57298];
assign t[57299] = t[57298] ^ n[57299];
assign t[57300] = t[57299] ^ n[57300];
assign t[57301] = t[57300] ^ n[57301];
assign t[57302] = t[57301] ^ n[57302];
assign t[57303] = t[57302] ^ n[57303];
assign t[57304] = t[57303] ^ n[57304];
assign t[57305] = t[57304] ^ n[57305];
assign t[57306] = t[57305] ^ n[57306];
assign t[57307] = t[57306] ^ n[57307];
assign t[57308] = t[57307] ^ n[57308];
assign t[57309] = t[57308] ^ n[57309];
assign t[57310] = t[57309] ^ n[57310];
assign t[57311] = t[57310] ^ n[57311];
assign t[57312] = t[57311] ^ n[57312];
assign t[57313] = t[57312] ^ n[57313];
assign t[57314] = t[57313] ^ n[57314];
assign t[57315] = t[57314] ^ n[57315];
assign t[57316] = t[57315] ^ n[57316];
assign t[57317] = t[57316] ^ n[57317];
assign t[57318] = t[57317] ^ n[57318];
assign t[57319] = t[57318] ^ n[57319];
assign t[57320] = t[57319] ^ n[57320];
assign t[57321] = t[57320] ^ n[57321];
assign t[57322] = t[57321] ^ n[57322];
assign t[57323] = t[57322] ^ n[57323];
assign t[57324] = t[57323] ^ n[57324];
assign t[57325] = t[57324] ^ n[57325];
assign t[57326] = t[57325] ^ n[57326];
assign t[57327] = t[57326] ^ n[57327];
assign t[57328] = t[57327] ^ n[57328];
assign t[57329] = t[57328] ^ n[57329];
assign t[57330] = t[57329] ^ n[57330];
assign t[57331] = t[57330] ^ n[57331];
assign t[57332] = t[57331] ^ n[57332];
assign t[57333] = t[57332] ^ n[57333];
assign t[57334] = t[57333] ^ n[57334];
assign t[57335] = t[57334] ^ n[57335];
assign t[57336] = t[57335] ^ n[57336];
assign t[57337] = t[57336] ^ n[57337];
assign t[57338] = t[57337] ^ n[57338];
assign t[57339] = t[57338] ^ n[57339];
assign t[57340] = t[57339] ^ n[57340];
assign t[57341] = t[57340] ^ n[57341];
assign t[57342] = t[57341] ^ n[57342];
assign t[57343] = t[57342] ^ n[57343];
assign t[57344] = t[57343] ^ n[57344];
assign t[57345] = t[57344] ^ n[57345];
assign t[57346] = t[57345] ^ n[57346];
assign t[57347] = t[57346] ^ n[57347];
assign t[57348] = t[57347] ^ n[57348];
assign t[57349] = t[57348] ^ n[57349];
assign t[57350] = t[57349] ^ n[57350];
assign t[57351] = t[57350] ^ n[57351];
assign t[57352] = t[57351] ^ n[57352];
assign t[57353] = t[57352] ^ n[57353];
assign t[57354] = t[57353] ^ n[57354];
assign t[57355] = t[57354] ^ n[57355];
assign t[57356] = t[57355] ^ n[57356];
assign t[57357] = t[57356] ^ n[57357];
assign t[57358] = t[57357] ^ n[57358];
assign t[57359] = t[57358] ^ n[57359];
assign t[57360] = t[57359] ^ n[57360];
assign t[57361] = t[57360] ^ n[57361];
assign t[57362] = t[57361] ^ n[57362];
assign t[57363] = t[57362] ^ n[57363];
assign t[57364] = t[57363] ^ n[57364];
assign t[57365] = t[57364] ^ n[57365];
assign t[57366] = t[57365] ^ n[57366];
assign t[57367] = t[57366] ^ n[57367];
assign t[57368] = t[57367] ^ n[57368];
assign t[57369] = t[57368] ^ n[57369];
assign t[57370] = t[57369] ^ n[57370];
assign t[57371] = t[57370] ^ n[57371];
assign t[57372] = t[57371] ^ n[57372];
assign t[57373] = t[57372] ^ n[57373];
assign t[57374] = t[57373] ^ n[57374];
assign t[57375] = t[57374] ^ n[57375];
assign t[57376] = t[57375] ^ n[57376];
assign t[57377] = t[57376] ^ n[57377];
assign t[57378] = t[57377] ^ n[57378];
assign t[57379] = t[57378] ^ n[57379];
assign t[57380] = t[57379] ^ n[57380];
assign t[57381] = t[57380] ^ n[57381];
assign t[57382] = t[57381] ^ n[57382];
assign t[57383] = t[57382] ^ n[57383];
assign t[57384] = t[57383] ^ n[57384];
assign t[57385] = t[57384] ^ n[57385];
assign t[57386] = t[57385] ^ n[57386];
assign t[57387] = t[57386] ^ n[57387];
assign t[57388] = t[57387] ^ n[57388];
assign t[57389] = t[57388] ^ n[57389];
assign t[57390] = t[57389] ^ n[57390];
assign t[57391] = t[57390] ^ n[57391];
assign t[57392] = t[57391] ^ n[57392];
assign t[57393] = t[57392] ^ n[57393];
assign t[57394] = t[57393] ^ n[57394];
assign t[57395] = t[57394] ^ n[57395];
assign t[57396] = t[57395] ^ n[57396];
assign t[57397] = t[57396] ^ n[57397];
assign t[57398] = t[57397] ^ n[57398];
assign t[57399] = t[57398] ^ n[57399];
assign t[57400] = t[57399] ^ n[57400];
assign t[57401] = t[57400] ^ n[57401];
assign t[57402] = t[57401] ^ n[57402];
assign t[57403] = t[57402] ^ n[57403];
assign t[57404] = t[57403] ^ n[57404];
assign t[57405] = t[57404] ^ n[57405];
assign t[57406] = t[57405] ^ n[57406];
assign t[57407] = t[57406] ^ n[57407];
assign t[57408] = t[57407] ^ n[57408];
assign t[57409] = t[57408] ^ n[57409];
assign t[57410] = t[57409] ^ n[57410];
assign t[57411] = t[57410] ^ n[57411];
assign t[57412] = t[57411] ^ n[57412];
assign t[57413] = t[57412] ^ n[57413];
assign t[57414] = t[57413] ^ n[57414];
assign t[57415] = t[57414] ^ n[57415];
assign t[57416] = t[57415] ^ n[57416];
assign t[57417] = t[57416] ^ n[57417];
assign t[57418] = t[57417] ^ n[57418];
assign t[57419] = t[57418] ^ n[57419];
assign t[57420] = t[57419] ^ n[57420];
assign t[57421] = t[57420] ^ n[57421];
assign t[57422] = t[57421] ^ n[57422];
assign t[57423] = t[57422] ^ n[57423];
assign t[57424] = t[57423] ^ n[57424];
assign t[57425] = t[57424] ^ n[57425];
assign t[57426] = t[57425] ^ n[57426];
assign t[57427] = t[57426] ^ n[57427];
assign t[57428] = t[57427] ^ n[57428];
assign t[57429] = t[57428] ^ n[57429];
assign t[57430] = t[57429] ^ n[57430];
assign t[57431] = t[57430] ^ n[57431];
assign t[57432] = t[57431] ^ n[57432];
assign t[57433] = t[57432] ^ n[57433];
assign t[57434] = t[57433] ^ n[57434];
assign t[57435] = t[57434] ^ n[57435];
assign t[57436] = t[57435] ^ n[57436];
assign t[57437] = t[57436] ^ n[57437];
assign t[57438] = t[57437] ^ n[57438];
assign t[57439] = t[57438] ^ n[57439];
assign t[57440] = t[57439] ^ n[57440];
assign t[57441] = t[57440] ^ n[57441];
assign t[57442] = t[57441] ^ n[57442];
assign t[57443] = t[57442] ^ n[57443];
assign t[57444] = t[57443] ^ n[57444];
assign t[57445] = t[57444] ^ n[57445];
assign t[57446] = t[57445] ^ n[57446];
assign t[57447] = t[57446] ^ n[57447];
assign t[57448] = t[57447] ^ n[57448];
assign t[57449] = t[57448] ^ n[57449];
assign t[57450] = t[57449] ^ n[57450];
assign t[57451] = t[57450] ^ n[57451];
assign t[57452] = t[57451] ^ n[57452];
assign t[57453] = t[57452] ^ n[57453];
assign t[57454] = t[57453] ^ n[57454];
assign t[57455] = t[57454] ^ n[57455];
assign t[57456] = t[57455] ^ n[57456];
assign t[57457] = t[57456] ^ n[57457];
assign t[57458] = t[57457] ^ n[57458];
assign t[57459] = t[57458] ^ n[57459];
assign t[57460] = t[57459] ^ n[57460];
assign t[57461] = t[57460] ^ n[57461];
assign t[57462] = t[57461] ^ n[57462];
assign t[57463] = t[57462] ^ n[57463];
assign t[57464] = t[57463] ^ n[57464];
assign t[57465] = t[57464] ^ n[57465];
assign t[57466] = t[57465] ^ n[57466];
assign t[57467] = t[57466] ^ n[57467];
assign t[57468] = t[57467] ^ n[57468];
assign t[57469] = t[57468] ^ n[57469];
assign t[57470] = t[57469] ^ n[57470];
assign t[57471] = t[57470] ^ n[57471];
assign t[57472] = t[57471] ^ n[57472];
assign t[57473] = t[57472] ^ n[57473];
assign t[57474] = t[57473] ^ n[57474];
assign t[57475] = t[57474] ^ n[57475];
assign t[57476] = t[57475] ^ n[57476];
assign t[57477] = t[57476] ^ n[57477];
assign t[57478] = t[57477] ^ n[57478];
assign t[57479] = t[57478] ^ n[57479];
assign t[57480] = t[57479] ^ n[57480];
assign t[57481] = t[57480] ^ n[57481];
assign t[57482] = t[57481] ^ n[57482];
assign t[57483] = t[57482] ^ n[57483];
assign t[57484] = t[57483] ^ n[57484];
assign t[57485] = t[57484] ^ n[57485];
assign t[57486] = t[57485] ^ n[57486];
assign t[57487] = t[57486] ^ n[57487];
assign t[57488] = t[57487] ^ n[57488];
assign t[57489] = t[57488] ^ n[57489];
assign t[57490] = t[57489] ^ n[57490];
assign t[57491] = t[57490] ^ n[57491];
assign t[57492] = t[57491] ^ n[57492];
assign t[57493] = t[57492] ^ n[57493];
assign t[57494] = t[57493] ^ n[57494];
assign t[57495] = t[57494] ^ n[57495];
assign t[57496] = t[57495] ^ n[57496];
assign t[57497] = t[57496] ^ n[57497];
assign t[57498] = t[57497] ^ n[57498];
assign t[57499] = t[57498] ^ n[57499];
assign t[57500] = t[57499] ^ n[57500];
assign t[57501] = t[57500] ^ n[57501];
assign t[57502] = t[57501] ^ n[57502];
assign t[57503] = t[57502] ^ n[57503];
assign t[57504] = t[57503] ^ n[57504];
assign t[57505] = t[57504] ^ n[57505];
assign t[57506] = t[57505] ^ n[57506];
assign t[57507] = t[57506] ^ n[57507];
assign t[57508] = t[57507] ^ n[57508];
assign t[57509] = t[57508] ^ n[57509];
assign t[57510] = t[57509] ^ n[57510];
assign t[57511] = t[57510] ^ n[57511];
assign t[57512] = t[57511] ^ n[57512];
assign t[57513] = t[57512] ^ n[57513];
assign t[57514] = t[57513] ^ n[57514];
assign t[57515] = t[57514] ^ n[57515];
assign t[57516] = t[57515] ^ n[57516];
assign t[57517] = t[57516] ^ n[57517];
assign t[57518] = t[57517] ^ n[57518];
assign t[57519] = t[57518] ^ n[57519];
assign t[57520] = t[57519] ^ n[57520];
assign t[57521] = t[57520] ^ n[57521];
assign t[57522] = t[57521] ^ n[57522];
assign t[57523] = t[57522] ^ n[57523];
assign t[57524] = t[57523] ^ n[57524];
assign t[57525] = t[57524] ^ n[57525];
assign t[57526] = t[57525] ^ n[57526];
assign t[57527] = t[57526] ^ n[57527];
assign t[57528] = t[57527] ^ n[57528];
assign t[57529] = t[57528] ^ n[57529];
assign t[57530] = t[57529] ^ n[57530];
assign t[57531] = t[57530] ^ n[57531];
assign t[57532] = t[57531] ^ n[57532];
assign t[57533] = t[57532] ^ n[57533];
assign t[57534] = t[57533] ^ n[57534];
assign t[57535] = t[57534] ^ n[57535];
assign t[57536] = t[57535] ^ n[57536];
assign t[57537] = t[57536] ^ n[57537];
assign t[57538] = t[57537] ^ n[57538];
assign t[57539] = t[57538] ^ n[57539];
assign t[57540] = t[57539] ^ n[57540];
assign t[57541] = t[57540] ^ n[57541];
assign t[57542] = t[57541] ^ n[57542];
assign t[57543] = t[57542] ^ n[57543];
assign t[57544] = t[57543] ^ n[57544];
assign t[57545] = t[57544] ^ n[57545];
assign t[57546] = t[57545] ^ n[57546];
assign t[57547] = t[57546] ^ n[57547];
assign t[57548] = t[57547] ^ n[57548];
assign t[57549] = t[57548] ^ n[57549];
assign t[57550] = t[57549] ^ n[57550];
assign t[57551] = t[57550] ^ n[57551];
assign t[57552] = t[57551] ^ n[57552];
assign t[57553] = t[57552] ^ n[57553];
assign t[57554] = t[57553] ^ n[57554];
assign t[57555] = t[57554] ^ n[57555];
assign t[57556] = t[57555] ^ n[57556];
assign t[57557] = t[57556] ^ n[57557];
assign t[57558] = t[57557] ^ n[57558];
assign t[57559] = t[57558] ^ n[57559];
assign t[57560] = t[57559] ^ n[57560];
assign t[57561] = t[57560] ^ n[57561];
assign t[57562] = t[57561] ^ n[57562];
assign t[57563] = t[57562] ^ n[57563];
assign t[57564] = t[57563] ^ n[57564];
assign t[57565] = t[57564] ^ n[57565];
assign t[57566] = t[57565] ^ n[57566];
assign t[57567] = t[57566] ^ n[57567];
assign t[57568] = t[57567] ^ n[57568];
assign t[57569] = t[57568] ^ n[57569];
assign t[57570] = t[57569] ^ n[57570];
assign t[57571] = t[57570] ^ n[57571];
assign t[57572] = t[57571] ^ n[57572];
assign t[57573] = t[57572] ^ n[57573];
assign t[57574] = t[57573] ^ n[57574];
assign t[57575] = t[57574] ^ n[57575];
assign t[57576] = t[57575] ^ n[57576];
assign t[57577] = t[57576] ^ n[57577];
assign t[57578] = t[57577] ^ n[57578];
assign t[57579] = t[57578] ^ n[57579];
assign t[57580] = t[57579] ^ n[57580];
assign t[57581] = t[57580] ^ n[57581];
assign t[57582] = t[57581] ^ n[57582];
assign t[57583] = t[57582] ^ n[57583];
assign t[57584] = t[57583] ^ n[57584];
assign t[57585] = t[57584] ^ n[57585];
assign t[57586] = t[57585] ^ n[57586];
assign t[57587] = t[57586] ^ n[57587];
assign t[57588] = t[57587] ^ n[57588];
assign t[57589] = t[57588] ^ n[57589];
assign t[57590] = t[57589] ^ n[57590];
assign t[57591] = t[57590] ^ n[57591];
assign t[57592] = t[57591] ^ n[57592];
assign t[57593] = t[57592] ^ n[57593];
assign t[57594] = t[57593] ^ n[57594];
assign t[57595] = t[57594] ^ n[57595];
assign t[57596] = t[57595] ^ n[57596];
assign t[57597] = t[57596] ^ n[57597];
assign t[57598] = t[57597] ^ n[57598];
assign t[57599] = t[57598] ^ n[57599];
assign t[57600] = t[57599] ^ n[57600];
assign t[57601] = t[57600] ^ n[57601];
assign t[57602] = t[57601] ^ n[57602];
assign t[57603] = t[57602] ^ n[57603];
assign t[57604] = t[57603] ^ n[57604];
assign t[57605] = t[57604] ^ n[57605];
assign t[57606] = t[57605] ^ n[57606];
assign t[57607] = t[57606] ^ n[57607];
assign t[57608] = t[57607] ^ n[57608];
assign t[57609] = t[57608] ^ n[57609];
assign t[57610] = t[57609] ^ n[57610];
assign t[57611] = t[57610] ^ n[57611];
assign t[57612] = t[57611] ^ n[57612];
assign t[57613] = t[57612] ^ n[57613];
assign t[57614] = t[57613] ^ n[57614];
assign t[57615] = t[57614] ^ n[57615];
assign t[57616] = t[57615] ^ n[57616];
assign t[57617] = t[57616] ^ n[57617];
assign t[57618] = t[57617] ^ n[57618];
assign t[57619] = t[57618] ^ n[57619];
assign t[57620] = t[57619] ^ n[57620];
assign t[57621] = t[57620] ^ n[57621];
assign t[57622] = t[57621] ^ n[57622];
assign t[57623] = t[57622] ^ n[57623];
assign t[57624] = t[57623] ^ n[57624];
assign t[57625] = t[57624] ^ n[57625];
assign t[57626] = t[57625] ^ n[57626];
assign t[57627] = t[57626] ^ n[57627];
assign t[57628] = t[57627] ^ n[57628];
assign t[57629] = t[57628] ^ n[57629];
assign t[57630] = t[57629] ^ n[57630];
assign t[57631] = t[57630] ^ n[57631];
assign t[57632] = t[57631] ^ n[57632];
assign t[57633] = t[57632] ^ n[57633];
assign t[57634] = t[57633] ^ n[57634];
assign t[57635] = t[57634] ^ n[57635];
assign t[57636] = t[57635] ^ n[57636];
assign t[57637] = t[57636] ^ n[57637];
assign t[57638] = t[57637] ^ n[57638];
assign t[57639] = t[57638] ^ n[57639];
assign t[57640] = t[57639] ^ n[57640];
assign t[57641] = t[57640] ^ n[57641];
assign t[57642] = t[57641] ^ n[57642];
assign t[57643] = t[57642] ^ n[57643];
assign t[57644] = t[57643] ^ n[57644];
assign t[57645] = t[57644] ^ n[57645];
assign t[57646] = t[57645] ^ n[57646];
assign t[57647] = t[57646] ^ n[57647];
assign t[57648] = t[57647] ^ n[57648];
assign t[57649] = t[57648] ^ n[57649];
assign t[57650] = t[57649] ^ n[57650];
assign t[57651] = t[57650] ^ n[57651];
assign t[57652] = t[57651] ^ n[57652];
assign t[57653] = t[57652] ^ n[57653];
assign t[57654] = t[57653] ^ n[57654];
assign t[57655] = t[57654] ^ n[57655];
assign t[57656] = t[57655] ^ n[57656];
assign t[57657] = t[57656] ^ n[57657];
assign t[57658] = t[57657] ^ n[57658];
assign t[57659] = t[57658] ^ n[57659];
assign t[57660] = t[57659] ^ n[57660];
assign t[57661] = t[57660] ^ n[57661];
assign t[57662] = t[57661] ^ n[57662];
assign t[57663] = t[57662] ^ n[57663];
assign t[57664] = t[57663] ^ n[57664];
assign t[57665] = t[57664] ^ n[57665];
assign t[57666] = t[57665] ^ n[57666];
assign t[57667] = t[57666] ^ n[57667];
assign t[57668] = t[57667] ^ n[57668];
assign t[57669] = t[57668] ^ n[57669];
assign t[57670] = t[57669] ^ n[57670];
assign t[57671] = t[57670] ^ n[57671];
assign t[57672] = t[57671] ^ n[57672];
assign t[57673] = t[57672] ^ n[57673];
assign t[57674] = t[57673] ^ n[57674];
assign t[57675] = t[57674] ^ n[57675];
assign t[57676] = t[57675] ^ n[57676];
assign t[57677] = t[57676] ^ n[57677];
assign t[57678] = t[57677] ^ n[57678];
assign t[57679] = t[57678] ^ n[57679];
assign t[57680] = t[57679] ^ n[57680];
assign t[57681] = t[57680] ^ n[57681];
assign t[57682] = t[57681] ^ n[57682];
assign t[57683] = t[57682] ^ n[57683];
assign t[57684] = t[57683] ^ n[57684];
assign t[57685] = t[57684] ^ n[57685];
assign t[57686] = t[57685] ^ n[57686];
assign t[57687] = t[57686] ^ n[57687];
assign t[57688] = t[57687] ^ n[57688];
assign t[57689] = t[57688] ^ n[57689];
assign t[57690] = t[57689] ^ n[57690];
assign t[57691] = t[57690] ^ n[57691];
assign t[57692] = t[57691] ^ n[57692];
assign t[57693] = t[57692] ^ n[57693];
assign t[57694] = t[57693] ^ n[57694];
assign t[57695] = t[57694] ^ n[57695];
assign t[57696] = t[57695] ^ n[57696];
assign t[57697] = t[57696] ^ n[57697];
assign t[57698] = t[57697] ^ n[57698];
assign t[57699] = t[57698] ^ n[57699];
assign t[57700] = t[57699] ^ n[57700];
assign t[57701] = t[57700] ^ n[57701];
assign t[57702] = t[57701] ^ n[57702];
assign t[57703] = t[57702] ^ n[57703];
assign t[57704] = t[57703] ^ n[57704];
assign t[57705] = t[57704] ^ n[57705];
assign t[57706] = t[57705] ^ n[57706];
assign t[57707] = t[57706] ^ n[57707];
assign t[57708] = t[57707] ^ n[57708];
assign t[57709] = t[57708] ^ n[57709];
assign t[57710] = t[57709] ^ n[57710];
assign t[57711] = t[57710] ^ n[57711];
assign t[57712] = t[57711] ^ n[57712];
assign t[57713] = t[57712] ^ n[57713];
assign t[57714] = t[57713] ^ n[57714];
assign t[57715] = t[57714] ^ n[57715];
assign t[57716] = t[57715] ^ n[57716];
assign t[57717] = t[57716] ^ n[57717];
assign t[57718] = t[57717] ^ n[57718];
assign t[57719] = t[57718] ^ n[57719];
assign t[57720] = t[57719] ^ n[57720];
assign t[57721] = t[57720] ^ n[57721];
assign t[57722] = t[57721] ^ n[57722];
assign t[57723] = t[57722] ^ n[57723];
assign t[57724] = t[57723] ^ n[57724];
assign t[57725] = t[57724] ^ n[57725];
assign t[57726] = t[57725] ^ n[57726];
assign t[57727] = t[57726] ^ n[57727];
assign t[57728] = t[57727] ^ n[57728];
assign t[57729] = t[57728] ^ n[57729];
assign t[57730] = t[57729] ^ n[57730];
assign t[57731] = t[57730] ^ n[57731];
assign t[57732] = t[57731] ^ n[57732];
assign t[57733] = t[57732] ^ n[57733];
assign t[57734] = t[57733] ^ n[57734];
assign t[57735] = t[57734] ^ n[57735];
assign t[57736] = t[57735] ^ n[57736];
assign t[57737] = t[57736] ^ n[57737];
assign t[57738] = t[57737] ^ n[57738];
assign t[57739] = t[57738] ^ n[57739];
assign t[57740] = t[57739] ^ n[57740];
assign t[57741] = t[57740] ^ n[57741];
assign t[57742] = t[57741] ^ n[57742];
assign t[57743] = t[57742] ^ n[57743];
assign t[57744] = t[57743] ^ n[57744];
assign t[57745] = t[57744] ^ n[57745];
assign t[57746] = t[57745] ^ n[57746];
assign t[57747] = t[57746] ^ n[57747];
assign t[57748] = t[57747] ^ n[57748];
assign t[57749] = t[57748] ^ n[57749];
assign t[57750] = t[57749] ^ n[57750];
assign t[57751] = t[57750] ^ n[57751];
assign t[57752] = t[57751] ^ n[57752];
assign t[57753] = t[57752] ^ n[57753];
assign t[57754] = t[57753] ^ n[57754];
assign t[57755] = t[57754] ^ n[57755];
assign t[57756] = t[57755] ^ n[57756];
assign t[57757] = t[57756] ^ n[57757];
assign t[57758] = t[57757] ^ n[57758];
assign t[57759] = t[57758] ^ n[57759];
assign t[57760] = t[57759] ^ n[57760];
assign t[57761] = t[57760] ^ n[57761];
assign t[57762] = t[57761] ^ n[57762];
assign t[57763] = t[57762] ^ n[57763];
assign t[57764] = t[57763] ^ n[57764];
assign t[57765] = t[57764] ^ n[57765];
assign t[57766] = t[57765] ^ n[57766];
assign t[57767] = t[57766] ^ n[57767];
assign t[57768] = t[57767] ^ n[57768];
assign t[57769] = t[57768] ^ n[57769];
assign t[57770] = t[57769] ^ n[57770];
assign t[57771] = t[57770] ^ n[57771];
assign t[57772] = t[57771] ^ n[57772];
assign t[57773] = t[57772] ^ n[57773];
assign t[57774] = t[57773] ^ n[57774];
assign t[57775] = t[57774] ^ n[57775];
assign t[57776] = t[57775] ^ n[57776];
assign t[57777] = t[57776] ^ n[57777];
assign t[57778] = t[57777] ^ n[57778];
assign t[57779] = t[57778] ^ n[57779];
assign t[57780] = t[57779] ^ n[57780];
assign t[57781] = t[57780] ^ n[57781];
assign t[57782] = t[57781] ^ n[57782];
assign t[57783] = t[57782] ^ n[57783];
assign t[57784] = t[57783] ^ n[57784];
assign t[57785] = t[57784] ^ n[57785];
assign t[57786] = t[57785] ^ n[57786];
assign t[57787] = t[57786] ^ n[57787];
assign t[57788] = t[57787] ^ n[57788];
assign t[57789] = t[57788] ^ n[57789];
assign t[57790] = t[57789] ^ n[57790];
assign t[57791] = t[57790] ^ n[57791];
assign t[57792] = t[57791] ^ n[57792];
assign t[57793] = t[57792] ^ n[57793];
assign t[57794] = t[57793] ^ n[57794];
assign t[57795] = t[57794] ^ n[57795];
assign t[57796] = t[57795] ^ n[57796];
assign t[57797] = t[57796] ^ n[57797];
assign t[57798] = t[57797] ^ n[57798];
assign t[57799] = t[57798] ^ n[57799];
assign t[57800] = t[57799] ^ n[57800];
assign t[57801] = t[57800] ^ n[57801];
assign t[57802] = t[57801] ^ n[57802];
assign t[57803] = t[57802] ^ n[57803];
assign t[57804] = t[57803] ^ n[57804];
assign t[57805] = t[57804] ^ n[57805];
assign t[57806] = t[57805] ^ n[57806];
assign t[57807] = t[57806] ^ n[57807];
assign t[57808] = t[57807] ^ n[57808];
assign t[57809] = t[57808] ^ n[57809];
assign t[57810] = t[57809] ^ n[57810];
assign t[57811] = t[57810] ^ n[57811];
assign t[57812] = t[57811] ^ n[57812];
assign t[57813] = t[57812] ^ n[57813];
assign t[57814] = t[57813] ^ n[57814];
assign t[57815] = t[57814] ^ n[57815];
assign t[57816] = t[57815] ^ n[57816];
assign t[57817] = t[57816] ^ n[57817];
assign t[57818] = t[57817] ^ n[57818];
assign t[57819] = t[57818] ^ n[57819];
assign t[57820] = t[57819] ^ n[57820];
assign t[57821] = t[57820] ^ n[57821];
assign t[57822] = t[57821] ^ n[57822];
assign t[57823] = t[57822] ^ n[57823];
assign t[57824] = t[57823] ^ n[57824];
assign t[57825] = t[57824] ^ n[57825];
assign t[57826] = t[57825] ^ n[57826];
assign t[57827] = t[57826] ^ n[57827];
assign t[57828] = t[57827] ^ n[57828];
assign t[57829] = t[57828] ^ n[57829];
assign t[57830] = t[57829] ^ n[57830];
assign t[57831] = t[57830] ^ n[57831];
assign t[57832] = t[57831] ^ n[57832];
assign t[57833] = t[57832] ^ n[57833];
assign t[57834] = t[57833] ^ n[57834];
assign t[57835] = t[57834] ^ n[57835];
assign t[57836] = t[57835] ^ n[57836];
assign t[57837] = t[57836] ^ n[57837];
assign t[57838] = t[57837] ^ n[57838];
assign t[57839] = t[57838] ^ n[57839];
assign t[57840] = t[57839] ^ n[57840];
assign t[57841] = t[57840] ^ n[57841];
assign t[57842] = t[57841] ^ n[57842];
assign t[57843] = t[57842] ^ n[57843];
assign t[57844] = t[57843] ^ n[57844];
assign t[57845] = t[57844] ^ n[57845];
assign t[57846] = t[57845] ^ n[57846];
assign t[57847] = t[57846] ^ n[57847];
assign t[57848] = t[57847] ^ n[57848];
assign t[57849] = t[57848] ^ n[57849];
assign t[57850] = t[57849] ^ n[57850];
assign t[57851] = t[57850] ^ n[57851];
assign t[57852] = t[57851] ^ n[57852];
assign t[57853] = t[57852] ^ n[57853];
assign t[57854] = t[57853] ^ n[57854];
assign t[57855] = t[57854] ^ n[57855];
assign t[57856] = t[57855] ^ n[57856];
assign t[57857] = t[57856] ^ n[57857];
assign t[57858] = t[57857] ^ n[57858];
assign t[57859] = t[57858] ^ n[57859];
assign t[57860] = t[57859] ^ n[57860];
assign t[57861] = t[57860] ^ n[57861];
assign t[57862] = t[57861] ^ n[57862];
assign t[57863] = t[57862] ^ n[57863];
assign t[57864] = t[57863] ^ n[57864];
assign t[57865] = t[57864] ^ n[57865];
assign t[57866] = t[57865] ^ n[57866];
assign t[57867] = t[57866] ^ n[57867];
assign t[57868] = t[57867] ^ n[57868];
assign t[57869] = t[57868] ^ n[57869];
assign t[57870] = t[57869] ^ n[57870];
assign t[57871] = t[57870] ^ n[57871];
assign t[57872] = t[57871] ^ n[57872];
assign t[57873] = t[57872] ^ n[57873];
assign t[57874] = t[57873] ^ n[57874];
assign t[57875] = t[57874] ^ n[57875];
assign t[57876] = t[57875] ^ n[57876];
assign t[57877] = t[57876] ^ n[57877];
assign t[57878] = t[57877] ^ n[57878];
assign t[57879] = t[57878] ^ n[57879];
assign t[57880] = t[57879] ^ n[57880];
assign t[57881] = t[57880] ^ n[57881];
assign t[57882] = t[57881] ^ n[57882];
assign t[57883] = t[57882] ^ n[57883];
assign t[57884] = t[57883] ^ n[57884];
assign t[57885] = t[57884] ^ n[57885];
assign t[57886] = t[57885] ^ n[57886];
assign t[57887] = t[57886] ^ n[57887];
assign t[57888] = t[57887] ^ n[57888];
assign t[57889] = t[57888] ^ n[57889];
assign t[57890] = t[57889] ^ n[57890];
assign t[57891] = t[57890] ^ n[57891];
assign t[57892] = t[57891] ^ n[57892];
assign t[57893] = t[57892] ^ n[57893];
assign t[57894] = t[57893] ^ n[57894];
assign t[57895] = t[57894] ^ n[57895];
assign t[57896] = t[57895] ^ n[57896];
assign t[57897] = t[57896] ^ n[57897];
assign t[57898] = t[57897] ^ n[57898];
assign t[57899] = t[57898] ^ n[57899];
assign t[57900] = t[57899] ^ n[57900];
assign t[57901] = t[57900] ^ n[57901];
assign t[57902] = t[57901] ^ n[57902];
assign t[57903] = t[57902] ^ n[57903];
assign t[57904] = t[57903] ^ n[57904];
assign t[57905] = t[57904] ^ n[57905];
assign t[57906] = t[57905] ^ n[57906];
assign t[57907] = t[57906] ^ n[57907];
assign t[57908] = t[57907] ^ n[57908];
assign t[57909] = t[57908] ^ n[57909];
assign t[57910] = t[57909] ^ n[57910];
assign t[57911] = t[57910] ^ n[57911];
assign t[57912] = t[57911] ^ n[57912];
assign t[57913] = t[57912] ^ n[57913];
assign t[57914] = t[57913] ^ n[57914];
assign t[57915] = t[57914] ^ n[57915];
assign t[57916] = t[57915] ^ n[57916];
assign t[57917] = t[57916] ^ n[57917];
assign t[57918] = t[57917] ^ n[57918];
assign t[57919] = t[57918] ^ n[57919];
assign t[57920] = t[57919] ^ n[57920];
assign t[57921] = t[57920] ^ n[57921];
assign t[57922] = t[57921] ^ n[57922];
assign t[57923] = t[57922] ^ n[57923];
assign t[57924] = t[57923] ^ n[57924];
assign t[57925] = t[57924] ^ n[57925];
assign t[57926] = t[57925] ^ n[57926];
assign t[57927] = t[57926] ^ n[57927];
assign t[57928] = t[57927] ^ n[57928];
assign t[57929] = t[57928] ^ n[57929];
assign t[57930] = t[57929] ^ n[57930];
assign t[57931] = t[57930] ^ n[57931];
assign t[57932] = t[57931] ^ n[57932];
assign t[57933] = t[57932] ^ n[57933];
assign t[57934] = t[57933] ^ n[57934];
assign t[57935] = t[57934] ^ n[57935];
assign t[57936] = t[57935] ^ n[57936];
assign t[57937] = t[57936] ^ n[57937];
assign t[57938] = t[57937] ^ n[57938];
assign t[57939] = t[57938] ^ n[57939];
assign t[57940] = t[57939] ^ n[57940];
assign t[57941] = t[57940] ^ n[57941];
assign t[57942] = t[57941] ^ n[57942];
assign t[57943] = t[57942] ^ n[57943];
assign t[57944] = t[57943] ^ n[57944];
assign t[57945] = t[57944] ^ n[57945];
assign t[57946] = t[57945] ^ n[57946];
assign t[57947] = t[57946] ^ n[57947];
assign t[57948] = t[57947] ^ n[57948];
assign t[57949] = t[57948] ^ n[57949];
assign t[57950] = t[57949] ^ n[57950];
assign t[57951] = t[57950] ^ n[57951];
assign t[57952] = t[57951] ^ n[57952];
assign t[57953] = t[57952] ^ n[57953];
assign t[57954] = t[57953] ^ n[57954];
assign t[57955] = t[57954] ^ n[57955];
assign t[57956] = t[57955] ^ n[57956];
assign t[57957] = t[57956] ^ n[57957];
assign t[57958] = t[57957] ^ n[57958];
assign t[57959] = t[57958] ^ n[57959];
assign t[57960] = t[57959] ^ n[57960];
assign t[57961] = t[57960] ^ n[57961];
assign t[57962] = t[57961] ^ n[57962];
assign t[57963] = t[57962] ^ n[57963];
assign t[57964] = t[57963] ^ n[57964];
assign t[57965] = t[57964] ^ n[57965];
assign t[57966] = t[57965] ^ n[57966];
assign t[57967] = t[57966] ^ n[57967];
assign t[57968] = t[57967] ^ n[57968];
assign t[57969] = t[57968] ^ n[57969];
assign t[57970] = t[57969] ^ n[57970];
assign t[57971] = t[57970] ^ n[57971];
assign t[57972] = t[57971] ^ n[57972];
assign t[57973] = t[57972] ^ n[57973];
assign t[57974] = t[57973] ^ n[57974];
assign t[57975] = t[57974] ^ n[57975];
assign t[57976] = t[57975] ^ n[57976];
assign t[57977] = t[57976] ^ n[57977];
assign t[57978] = t[57977] ^ n[57978];
assign t[57979] = t[57978] ^ n[57979];
assign t[57980] = t[57979] ^ n[57980];
assign t[57981] = t[57980] ^ n[57981];
assign t[57982] = t[57981] ^ n[57982];
assign t[57983] = t[57982] ^ n[57983];
assign t[57984] = t[57983] ^ n[57984];
assign t[57985] = t[57984] ^ n[57985];
assign t[57986] = t[57985] ^ n[57986];
assign t[57987] = t[57986] ^ n[57987];
assign t[57988] = t[57987] ^ n[57988];
assign t[57989] = t[57988] ^ n[57989];
assign t[57990] = t[57989] ^ n[57990];
assign t[57991] = t[57990] ^ n[57991];
assign t[57992] = t[57991] ^ n[57992];
assign t[57993] = t[57992] ^ n[57993];
assign t[57994] = t[57993] ^ n[57994];
assign t[57995] = t[57994] ^ n[57995];
assign t[57996] = t[57995] ^ n[57996];
assign t[57997] = t[57996] ^ n[57997];
assign t[57998] = t[57997] ^ n[57998];
assign t[57999] = t[57998] ^ n[57999];
assign t[58000] = t[57999] ^ n[58000];
assign t[58001] = t[58000] ^ n[58001];
assign t[58002] = t[58001] ^ n[58002];
assign t[58003] = t[58002] ^ n[58003];
assign t[58004] = t[58003] ^ n[58004];
assign t[58005] = t[58004] ^ n[58005];
assign t[58006] = t[58005] ^ n[58006];
assign t[58007] = t[58006] ^ n[58007];
assign t[58008] = t[58007] ^ n[58008];
assign t[58009] = t[58008] ^ n[58009];
assign t[58010] = t[58009] ^ n[58010];
assign t[58011] = t[58010] ^ n[58011];
assign t[58012] = t[58011] ^ n[58012];
assign t[58013] = t[58012] ^ n[58013];
assign t[58014] = t[58013] ^ n[58014];
assign t[58015] = t[58014] ^ n[58015];
assign t[58016] = t[58015] ^ n[58016];
assign t[58017] = t[58016] ^ n[58017];
assign t[58018] = t[58017] ^ n[58018];
assign t[58019] = t[58018] ^ n[58019];
assign t[58020] = t[58019] ^ n[58020];
assign t[58021] = t[58020] ^ n[58021];
assign t[58022] = t[58021] ^ n[58022];
assign t[58023] = t[58022] ^ n[58023];
assign t[58024] = t[58023] ^ n[58024];
assign t[58025] = t[58024] ^ n[58025];
assign t[58026] = t[58025] ^ n[58026];
assign t[58027] = t[58026] ^ n[58027];
assign t[58028] = t[58027] ^ n[58028];
assign t[58029] = t[58028] ^ n[58029];
assign t[58030] = t[58029] ^ n[58030];
assign t[58031] = t[58030] ^ n[58031];
assign t[58032] = t[58031] ^ n[58032];
assign t[58033] = t[58032] ^ n[58033];
assign t[58034] = t[58033] ^ n[58034];
assign t[58035] = t[58034] ^ n[58035];
assign t[58036] = t[58035] ^ n[58036];
assign t[58037] = t[58036] ^ n[58037];
assign t[58038] = t[58037] ^ n[58038];
assign t[58039] = t[58038] ^ n[58039];
assign t[58040] = t[58039] ^ n[58040];
assign t[58041] = t[58040] ^ n[58041];
assign t[58042] = t[58041] ^ n[58042];
assign t[58043] = t[58042] ^ n[58043];
assign t[58044] = t[58043] ^ n[58044];
assign t[58045] = t[58044] ^ n[58045];
assign t[58046] = t[58045] ^ n[58046];
assign t[58047] = t[58046] ^ n[58047];
assign t[58048] = t[58047] ^ n[58048];
assign t[58049] = t[58048] ^ n[58049];
assign t[58050] = t[58049] ^ n[58050];
assign t[58051] = t[58050] ^ n[58051];
assign t[58052] = t[58051] ^ n[58052];
assign t[58053] = t[58052] ^ n[58053];
assign t[58054] = t[58053] ^ n[58054];
assign t[58055] = t[58054] ^ n[58055];
assign t[58056] = t[58055] ^ n[58056];
assign t[58057] = t[58056] ^ n[58057];
assign t[58058] = t[58057] ^ n[58058];
assign t[58059] = t[58058] ^ n[58059];
assign t[58060] = t[58059] ^ n[58060];
assign t[58061] = t[58060] ^ n[58061];
assign t[58062] = t[58061] ^ n[58062];
assign t[58063] = t[58062] ^ n[58063];
assign t[58064] = t[58063] ^ n[58064];
assign t[58065] = t[58064] ^ n[58065];
assign t[58066] = t[58065] ^ n[58066];
assign t[58067] = t[58066] ^ n[58067];
assign t[58068] = t[58067] ^ n[58068];
assign t[58069] = t[58068] ^ n[58069];
assign t[58070] = t[58069] ^ n[58070];
assign t[58071] = t[58070] ^ n[58071];
assign t[58072] = t[58071] ^ n[58072];
assign t[58073] = t[58072] ^ n[58073];
assign t[58074] = t[58073] ^ n[58074];
assign t[58075] = t[58074] ^ n[58075];
assign t[58076] = t[58075] ^ n[58076];
assign t[58077] = t[58076] ^ n[58077];
assign t[58078] = t[58077] ^ n[58078];
assign t[58079] = t[58078] ^ n[58079];
assign t[58080] = t[58079] ^ n[58080];
assign t[58081] = t[58080] ^ n[58081];
assign t[58082] = t[58081] ^ n[58082];
assign t[58083] = t[58082] ^ n[58083];
assign t[58084] = t[58083] ^ n[58084];
assign t[58085] = t[58084] ^ n[58085];
assign t[58086] = t[58085] ^ n[58086];
assign t[58087] = t[58086] ^ n[58087];
assign t[58088] = t[58087] ^ n[58088];
assign t[58089] = t[58088] ^ n[58089];
assign t[58090] = t[58089] ^ n[58090];
assign t[58091] = t[58090] ^ n[58091];
assign t[58092] = t[58091] ^ n[58092];
assign t[58093] = t[58092] ^ n[58093];
assign t[58094] = t[58093] ^ n[58094];
assign t[58095] = t[58094] ^ n[58095];
assign t[58096] = t[58095] ^ n[58096];
assign t[58097] = t[58096] ^ n[58097];
assign t[58098] = t[58097] ^ n[58098];
assign t[58099] = t[58098] ^ n[58099];
assign t[58100] = t[58099] ^ n[58100];
assign t[58101] = t[58100] ^ n[58101];
assign t[58102] = t[58101] ^ n[58102];
assign t[58103] = t[58102] ^ n[58103];
assign t[58104] = t[58103] ^ n[58104];
assign t[58105] = t[58104] ^ n[58105];
assign t[58106] = t[58105] ^ n[58106];
assign t[58107] = t[58106] ^ n[58107];
assign t[58108] = t[58107] ^ n[58108];
assign t[58109] = t[58108] ^ n[58109];
assign t[58110] = t[58109] ^ n[58110];
assign t[58111] = t[58110] ^ n[58111];
assign t[58112] = t[58111] ^ n[58112];
assign t[58113] = t[58112] ^ n[58113];
assign t[58114] = t[58113] ^ n[58114];
assign t[58115] = t[58114] ^ n[58115];
assign t[58116] = t[58115] ^ n[58116];
assign t[58117] = t[58116] ^ n[58117];
assign t[58118] = t[58117] ^ n[58118];
assign t[58119] = t[58118] ^ n[58119];
assign t[58120] = t[58119] ^ n[58120];
assign t[58121] = t[58120] ^ n[58121];
assign t[58122] = t[58121] ^ n[58122];
assign t[58123] = t[58122] ^ n[58123];
assign t[58124] = t[58123] ^ n[58124];
assign t[58125] = t[58124] ^ n[58125];
assign t[58126] = t[58125] ^ n[58126];
assign t[58127] = t[58126] ^ n[58127];
assign t[58128] = t[58127] ^ n[58128];
assign t[58129] = t[58128] ^ n[58129];
assign t[58130] = t[58129] ^ n[58130];
assign t[58131] = t[58130] ^ n[58131];
assign t[58132] = t[58131] ^ n[58132];
assign t[58133] = t[58132] ^ n[58133];
assign t[58134] = t[58133] ^ n[58134];
assign t[58135] = t[58134] ^ n[58135];
assign t[58136] = t[58135] ^ n[58136];
assign t[58137] = t[58136] ^ n[58137];
assign t[58138] = t[58137] ^ n[58138];
assign t[58139] = t[58138] ^ n[58139];
assign t[58140] = t[58139] ^ n[58140];
assign t[58141] = t[58140] ^ n[58141];
assign t[58142] = t[58141] ^ n[58142];
assign t[58143] = t[58142] ^ n[58143];
assign t[58144] = t[58143] ^ n[58144];
assign t[58145] = t[58144] ^ n[58145];
assign t[58146] = t[58145] ^ n[58146];
assign t[58147] = t[58146] ^ n[58147];
assign t[58148] = t[58147] ^ n[58148];
assign t[58149] = t[58148] ^ n[58149];
assign t[58150] = t[58149] ^ n[58150];
assign t[58151] = t[58150] ^ n[58151];
assign t[58152] = t[58151] ^ n[58152];
assign t[58153] = t[58152] ^ n[58153];
assign t[58154] = t[58153] ^ n[58154];
assign t[58155] = t[58154] ^ n[58155];
assign t[58156] = t[58155] ^ n[58156];
assign t[58157] = t[58156] ^ n[58157];
assign t[58158] = t[58157] ^ n[58158];
assign t[58159] = t[58158] ^ n[58159];
assign t[58160] = t[58159] ^ n[58160];
assign t[58161] = t[58160] ^ n[58161];
assign t[58162] = t[58161] ^ n[58162];
assign t[58163] = t[58162] ^ n[58163];
assign t[58164] = t[58163] ^ n[58164];
assign t[58165] = t[58164] ^ n[58165];
assign t[58166] = t[58165] ^ n[58166];
assign t[58167] = t[58166] ^ n[58167];
assign t[58168] = t[58167] ^ n[58168];
assign t[58169] = t[58168] ^ n[58169];
assign t[58170] = t[58169] ^ n[58170];
assign t[58171] = t[58170] ^ n[58171];
assign t[58172] = t[58171] ^ n[58172];
assign t[58173] = t[58172] ^ n[58173];
assign t[58174] = t[58173] ^ n[58174];
assign t[58175] = t[58174] ^ n[58175];
assign t[58176] = t[58175] ^ n[58176];
assign t[58177] = t[58176] ^ n[58177];
assign t[58178] = t[58177] ^ n[58178];
assign t[58179] = t[58178] ^ n[58179];
assign t[58180] = t[58179] ^ n[58180];
assign t[58181] = t[58180] ^ n[58181];
assign t[58182] = t[58181] ^ n[58182];
assign t[58183] = t[58182] ^ n[58183];
assign t[58184] = t[58183] ^ n[58184];
assign t[58185] = t[58184] ^ n[58185];
assign t[58186] = t[58185] ^ n[58186];
assign t[58187] = t[58186] ^ n[58187];
assign t[58188] = t[58187] ^ n[58188];
assign t[58189] = t[58188] ^ n[58189];
assign t[58190] = t[58189] ^ n[58190];
assign t[58191] = t[58190] ^ n[58191];
assign t[58192] = t[58191] ^ n[58192];
assign t[58193] = t[58192] ^ n[58193];
assign t[58194] = t[58193] ^ n[58194];
assign t[58195] = t[58194] ^ n[58195];
assign t[58196] = t[58195] ^ n[58196];
assign t[58197] = t[58196] ^ n[58197];
assign t[58198] = t[58197] ^ n[58198];
assign t[58199] = t[58198] ^ n[58199];
assign t[58200] = t[58199] ^ n[58200];
assign t[58201] = t[58200] ^ n[58201];
assign t[58202] = t[58201] ^ n[58202];
assign t[58203] = t[58202] ^ n[58203];
assign t[58204] = t[58203] ^ n[58204];
assign t[58205] = t[58204] ^ n[58205];
assign t[58206] = t[58205] ^ n[58206];
assign t[58207] = t[58206] ^ n[58207];
assign t[58208] = t[58207] ^ n[58208];
assign t[58209] = t[58208] ^ n[58209];
assign t[58210] = t[58209] ^ n[58210];
assign t[58211] = t[58210] ^ n[58211];
assign t[58212] = t[58211] ^ n[58212];
assign t[58213] = t[58212] ^ n[58213];
assign t[58214] = t[58213] ^ n[58214];
assign t[58215] = t[58214] ^ n[58215];
assign t[58216] = t[58215] ^ n[58216];
assign t[58217] = t[58216] ^ n[58217];
assign t[58218] = t[58217] ^ n[58218];
assign t[58219] = t[58218] ^ n[58219];
assign t[58220] = t[58219] ^ n[58220];
assign t[58221] = t[58220] ^ n[58221];
assign t[58222] = t[58221] ^ n[58222];
assign t[58223] = t[58222] ^ n[58223];
assign t[58224] = t[58223] ^ n[58224];
assign t[58225] = t[58224] ^ n[58225];
assign t[58226] = t[58225] ^ n[58226];
assign t[58227] = t[58226] ^ n[58227];
assign t[58228] = t[58227] ^ n[58228];
assign t[58229] = t[58228] ^ n[58229];
assign t[58230] = t[58229] ^ n[58230];
assign t[58231] = t[58230] ^ n[58231];
assign t[58232] = t[58231] ^ n[58232];
assign t[58233] = t[58232] ^ n[58233];
assign t[58234] = t[58233] ^ n[58234];
assign t[58235] = t[58234] ^ n[58235];
assign t[58236] = t[58235] ^ n[58236];
assign t[58237] = t[58236] ^ n[58237];
assign t[58238] = t[58237] ^ n[58238];
assign t[58239] = t[58238] ^ n[58239];
assign t[58240] = t[58239] ^ n[58240];
assign t[58241] = t[58240] ^ n[58241];
assign t[58242] = t[58241] ^ n[58242];
assign t[58243] = t[58242] ^ n[58243];
assign t[58244] = t[58243] ^ n[58244];
assign t[58245] = t[58244] ^ n[58245];
assign t[58246] = t[58245] ^ n[58246];
assign t[58247] = t[58246] ^ n[58247];
assign t[58248] = t[58247] ^ n[58248];
assign t[58249] = t[58248] ^ n[58249];
assign t[58250] = t[58249] ^ n[58250];
assign t[58251] = t[58250] ^ n[58251];
assign t[58252] = t[58251] ^ n[58252];
assign t[58253] = t[58252] ^ n[58253];
assign t[58254] = t[58253] ^ n[58254];
assign t[58255] = t[58254] ^ n[58255];
assign t[58256] = t[58255] ^ n[58256];
assign t[58257] = t[58256] ^ n[58257];
assign t[58258] = t[58257] ^ n[58258];
assign t[58259] = t[58258] ^ n[58259];
assign t[58260] = t[58259] ^ n[58260];
assign t[58261] = t[58260] ^ n[58261];
assign t[58262] = t[58261] ^ n[58262];
assign t[58263] = t[58262] ^ n[58263];
assign t[58264] = t[58263] ^ n[58264];
assign t[58265] = t[58264] ^ n[58265];
assign t[58266] = t[58265] ^ n[58266];
assign t[58267] = t[58266] ^ n[58267];
assign t[58268] = t[58267] ^ n[58268];
assign t[58269] = t[58268] ^ n[58269];
assign t[58270] = t[58269] ^ n[58270];
assign t[58271] = t[58270] ^ n[58271];
assign t[58272] = t[58271] ^ n[58272];
assign t[58273] = t[58272] ^ n[58273];
assign t[58274] = t[58273] ^ n[58274];
assign t[58275] = t[58274] ^ n[58275];
assign t[58276] = t[58275] ^ n[58276];
assign t[58277] = t[58276] ^ n[58277];
assign t[58278] = t[58277] ^ n[58278];
assign t[58279] = t[58278] ^ n[58279];
assign t[58280] = t[58279] ^ n[58280];
assign t[58281] = t[58280] ^ n[58281];
assign t[58282] = t[58281] ^ n[58282];
assign t[58283] = t[58282] ^ n[58283];
assign t[58284] = t[58283] ^ n[58284];
assign t[58285] = t[58284] ^ n[58285];
assign t[58286] = t[58285] ^ n[58286];
assign t[58287] = t[58286] ^ n[58287];
assign t[58288] = t[58287] ^ n[58288];
assign t[58289] = t[58288] ^ n[58289];
assign t[58290] = t[58289] ^ n[58290];
assign t[58291] = t[58290] ^ n[58291];
assign t[58292] = t[58291] ^ n[58292];
assign t[58293] = t[58292] ^ n[58293];
assign t[58294] = t[58293] ^ n[58294];
assign t[58295] = t[58294] ^ n[58295];
assign t[58296] = t[58295] ^ n[58296];
assign t[58297] = t[58296] ^ n[58297];
assign t[58298] = t[58297] ^ n[58298];
assign t[58299] = t[58298] ^ n[58299];
assign t[58300] = t[58299] ^ n[58300];
assign t[58301] = t[58300] ^ n[58301];
assign t[58302] = t[58301] ^ n[58302];
assign t[58303] = t[58302] ^ n[58303];
assign t[58304] = t[58303] ^ n[58304];
assign t[58305] = t[58304] ^ n[58305];
assign t[58306] = t[58305] ^ n[58306];
assign t[58307] = t[58306] ^ n[58307];
assign t[58308] = t[58307] ^ n[58308];
assign t[58309] = t[58308] ^ n[58309];
assign t[58310] = t[58309] ^ n[58310];
assign t[58311] = t[58310] ^ n[58311];
assign t[58312] = t[58311] ^ n[58312];
assign t[58313] = t[58312] ^ n[58313];
assign t[58314] = t[58313] ^ n[58314];
assign t[58315] = t[58314] ^ n[58315];
assign t[58316] = t[58315] ^ n[58316];
assign t[58317] = t[58316] ^ n[58317];
assign t[58318] = t[58317] ^ n[58318];
assign t[58319] = t[58318] ^ n[58319];
assign t[58320] = t[58319] ^ n[58320];
assign t[58321] = t[58320] ^ n[58321];
assign t[58322] = t[58321] ^ n[58322];
assign t[58323] = t[58322] ^ n[58323];
assign t[58324] = t[58323] ^ n[58324];
assign t[58325] = t[58324] ^ n[58325];
assign t[58326] = t[58325] ^ n[58326];
assign t[58327] = t[58326] ^ n[58327];
assign t[58328] = t[58327] ^ n[58328];
assign t[58329] = t[58328] ^ n[58329];
assign t[58330] = t[58329] ^ n[58330];
assign t[58331] = t[58330] ^ n[58331];
assign t[58332] = t[58331] ^ n[58332];
assign t[58333] = t[58332] ^ n[58333];
assign t[58334] = t[58333] ^ n[58334];
assign t[58335] = t[58334] ^ n[58335];
assign t[58336] = t[58335] ^ n[58336];
assign t[58337] = t[58336] ^ n[58337];
assign t[58338] = t[58337] ^ n[58338];
assign t[58339] = t[58338] ^ n[58339];
assign t[58340] = t[58339] ^ n[58340];
assign t[58341] = t[58340] ^ n[58341];
assign t[58342] = t[58341] ^ n[58342];
assign t[58343] = t[58342] ^ n[58343];
assign t[58344] = t[58343] ^ n[58344];
assign t[58345] = t[58344] ^ n[58345];
assign t[58346] = t[58345] ^ n[58346];
assign t[58347] = t[58346] ^ n[58347];
assign t[58348] = t[58347] ^ n[58348];
assign t[58349] = t[58348] ^ n[58349];
assign t[58350] = t[58349] ^ n[58350];
assign t[58351] = t[58350] ^ n[58351];
assign t[58352] = t[58351] ^ n[58352];
assign t[58353] = t[58352] ^ n[58353];
assign t[58354] = t[58353] ^ n[58354];
assign t[58355] = t[58354] ^ n[58355];
assign t[58356] = t[58355] ^ n[58356];
assign t[58357] = t[58356] ^ n[58357];
assign t[58358] = t[58357] ^ n[58358];
assign t[58359] = t[58358] ^ n[58359];
assign t[58360] = t[58359] ^ n[58360];
assign t[58361] = t[58360] ^ n[58361];
assign t[58362] = t[58361] ^ n[58362];
assign t[58363] = t[58362] ^ n[58363];
assign t[58364] = t[58363] ^ n[58364];
assign t[58365] = t[58364] ^ n[58365];
assign t[58366] = t[58365] ^ n[58366];
assign t[58367] = t[58366] ^ n[58367];
assign t[58368] = t[58367] ^ n[58368];
assign t[58369] = t[58368] ^ n[58369];
assign t[58370] = t[58369] ^ n[58370];
assign t[58371] = t[58370] ^ n[58371];
assign t[58372] = t[58371] ^ n[58372];
assign t[58373] = t[58372] ^ n[58373];
assign t[58374] = t[58373] ^ n[58374];
assign t[58375] = t[58374] ^ n[58375];
assign t[58376] = t[58375] ^ n[58376];
assign t[58377] = t[58376] ^ n[58377];
assign t[58378] = t[58377] ^ n[58378];
assign t[58379] = t[58378] ^ n[58379];
assign t[58380] = t[58379] ^ n[58380];
assign t[58381] = t[58380] ^ n[58381];
assign t[58382] = t[58381] ^ n[58382];
assign t[58383] = t[58382] ^ n[58383];
assign t[58384] = t[58383] ^ n[58384];
assign t[58385] = t[58384] ^ n[58385];
assign t[58386] = t[58385] ^ n[58386];
assign t[58387] = t[58386] ^ n[58387];
assign t[58388] = t[58387] ^ n[58388];
assign t[58389] = t[58388] ^ n[58389];
assign t[58390] = t[58389] ^ n[58390];
assign t[58391] = t[58390] ^ n[58391];
assign t[58392] = t[58391] ^ n[58392];
assign t[58393] = t[58392] ^ n[58393];
assign t[58394] = t[58393] ^ n[58394];
assign t[58395] = t[58394] ^ n[58395];
assign t[58396] = t[58395] ^ n[58396];
assign t[58397] = t[58396] ^ n[58397];
assign t[58398] = t[58397] ^ n[58398];
assign t[58399] = t[58398] ^ n[58399];
assign t[58400] = t[58399] ^ n[58400];
assign t[58401] = t[58400] ^ n[58401];
assign t[58402] = t[58401] ^ n[58402];
assign t[58403] = t[58402] ^ n[58403];
assign t[58404] = t[58403] ^ n[58404];
assign t[58405] = t[58404] ^ n[58405];
assign t[58406] = t[58405] ^ n[58406];
assign t[58407] = t[58406] ^ n[58407];
assign t[58408] = t[58407] ^ n[58408];
assign t[58409] = t[58408] ^ n[58409];
assign t[58410] = t[58409] ^ n[58410];
assign t[58411] = t[58410] ^ n[58411];
assign t[58412] = t[58411] ^ n[58412];
assign t[58413] = t[58412] ^ n[58413];
assign t[58414] = t[58413] ^ n[58414];
assign t[58415] = t[58414] ^ n[58415];
assign t[58416] = t[58415] ^ n[58416];
assign t[58417] = t[58416] ^ n[58417];
assign t[58418] = t[58417] ^ n[58418];
assign t[58419] = t[58418] ^ n[58419];
assign t[58420] = t[58419] ^ n[58420];
assign t[58421] = t[58420] ^ n[58421];
assign t[58422] = t[58421] ^ n[58422];
assign t[58423] = t[58422] ^ n[58423];
assign t[58424] = t[58423] ^ n[58424];
assign t[58425] = t[58424] ^ n[58425];
assign t[58426] = t[58425] ^ n[58426];
assign t[58427] = t[58426] ^ n[58427];
assign t[58428] = t[58427] ^ n[58428];
assign t[58429] = t[58428] ^ n[58429];
assign t[58430] = t[58429] ^ n[58430];
assign t[58431] = t[58430] ^ n[58431];
assign t[58432] = t[58431] ^ n[58432];
assign t[58433] = t[58432] ^ n[58433];
assign t[58434] = t[58433] ^ n[58434];
assign t[58435] = t[58434] ^ n[58435];
assign t[58436] = t[58435] ^ n[58436];
assign t[58437] = t[58436] ^ n[58437];
assign t[58438] = t[58437] ^ n[58438];
assign t[58439] = t[58438] ^ n[58439];
assign t[58440] = t[58439] ^ n[58440];
assign t[58441] = t[58440] ^ n[58441];
assign t[58442] = t[58441] ^ n[58442];
assign t[58443] = t[58442] ^ n[58443];
assign t[58444] = t[58443] ^ n[58444];
assign t[58445] = t[58444] ^ n[58445];
assign t[58446] = t[58445] ^ n[58446];
assign t[58447] = t[58446] ^ n[58447];
assign t[58448] = t[58447] ^ n[58448];
assign t[58449] = t[58448] ^ n[58449];
assign t[58450] = t[58449] ^ n[58450];
assign t[58451] = t[58450] ^ n[58451];
assign t[58452] = t[58451] ^ n[58452];
assign t[58453] = t[58452] ^ n[58453];
assign t[58454] = t[58453] ^ n[58454];
assign t[58455] = t[58454] ^ n[58455];
assign t[58456] = t[58455] ^ n[58456];
assign t[58457] = t[58456] ^ n[58457];
assign t[58458] = t[58457] ^ n[58458];
assign t[58459] = t[58458] ^ n[58459];
assign t[58460] = t[58459] ^ n[58460];
assign t[58461] = t[58460] ^ n[58461];
assign t[58462] = t[58461] ^ n[58462];
assign t[58463] = t[58462] ^ n[58463];
assign t[58464] = t[58463] ^ n[58464];
assign t[58465] = t[58464] ^ n[58465];
assign t[58466] = t[58465] ^ n[58466];
assign t[58467] = t[58466] ^ n[58467];
assign t[58468] = t[58467] ^ n[58468];
assign t[58469] = t[58468] ^ n[58469];
assign t[58470] = t[58469] ^ n[58470];
assign t[58471] = t[58470] ^ n[58471];
assign t[58472] = t[58471] ^ n[58472];
assign t[58473] = t[58472] ^ n[58473];
assign t[58474] = t[58473] ^ n[58474];
assign t[58475] = t[58474] ^ n[58475];
assign t[58476] = t[58475] ^ n[58476];
assign t[58477] = t[58476] ^ n[58477];
assign t[58478] = t[58477] ^ n[58478];
assign t[58479] = t[58478] ^ n[58479];
assign t[58480] = t[58479] ^ n[58480];
assign t[58481] = t[58480] ^ n[58481];
assign t[58482] = t[58481] ^ n[58482];
assign t[58483] = t[58482] ^ n[58483];
assign t[58484] = t[58483] ^ n[58484];
assign t[58485] = t[58484] ^ n[58485];
assign t[58486] = t[58485] ^ n[58486];
assign t[58487] = t[58486] ^ n[58487];
assign t[58488] = t[58487] ^ n[58488];
assign t[58489] = t[58488] ^ n[58489];
assign t[58490] = t[58489] ^ n[58490];
assign t[58491] = t[58490] ^ n[58491];
assign t[58492] = t[58491] ^ n[58492];
assign t[58493] = t[58492] ^ n[58493];
assign t[58494] = t[58493] ^ n[58494];
assign t[58495] = t[58494] ^ n[58495];
assign t[58496] = t[58495] ^ n[58496];
assign t[58497] = t[58496] ^ n[58497];
assign t[58498] = t[58497] ^ n[58498];
assign t[58499] = t[58498] ^ n[58499];
assign t[58500] = t[58499] ^ n[58500];
assign t[58501] = t[58500] ^ n[58501];
assign t[58502] = t[58501] ^ n[58502];
assign t[58503] = t[58502] ^ n[58503];
assign t[58504] = t[58503] ^ n[58504];
assign t[58505] = t[58504] ^ n[58505];
assign t[58506] = t[58505] ^ n[58506];
assign t[58507] = t[58506] ^ n[58507];
assign t[58508] = t[58507] ^ n[58508];
assign t[58509] = t[58508] ^ n[58509];
assign t[58510] = t[58509] ^ n[58510];
assign t[58511] = t[58510] ^ n[58511];
assign t[58512] = t[58511] ^ n[58512];
assign t[58513] = t[58512] ^ n[58513];
assign t[58514] = t[58513] ^ n[58514];
assign t[58515] = t[58514] ^ n[58515];
assign t[58516] = t[58515] ^ n[58516];
assign t[58517] = t[58516] ^ n[58517];
assign t[58518] = t[58517] ^ n[58518];
assign t[58519] = t[58518] ^ n[58519];
assign t[58520] = t[58519] ^ n[58520];
assign t[58521] = t[58520] ^ n[58521];
assign t[58522] = t[58521] ^ n[58522];
assign t[58523] = t[58522] ^ n[58523];
assign t[58524] = t[58523] ^ n[58524];
assign t[58525] = t[58524] ^ n[58525];
assign t[58526] = t[58525] ^ n[58526];
assign t[58527] = t[58526] ^ n[58527];
assign t[58528] = t[58527] ^ n[58528];
assign t[58529] = t[58528] ^ n[58529];
assign t[58530] = t[58529] ^ n[58530];
assign t[58531] = t[58530] ^ n[58531];
assign t[58532] = t[58531] ^ n[58532];
assign t[58533] = t[58532] ^ n[58533];
assign t[58534] = t[58533] ^ n[58534];
assign t[58535] = t[58534] ^ n[58535];
assign t[58536] = t[58535] ^ n[58536];
assign t[58537] = t[58536] ^ n[58537];
assign t[58538] = t[58537] ^ n[58538];
assign t[58539] = t[58538] ^ n[58539];
assign t[58540] = t[58539] ^ n[58540];
assign t[58541] = t[58540] ^ n[58541];
assign t[58542] = t[58541] ^ n[58542];
assign t[58543] = t[58542] ^ n[58543];
assign t[58544] = t[58543] ^ n[58544];
assign t[58545] = t[58544] ^ n[58545];
assign t[58546] = t[58545] ^ n[58546];
assign t[58547] = t[58546] ^ n[58547];
assign t[58548] = t[58547] ^ n[58548];
assign t[58549] = t[58548] ^ n[58549];
assign t[58550] = t[58549] ^ n[58550];
assign t[58551] = t[58550] ^ n[58551];
assign t[58552] = t[58551] ^ n[58552];
assign t[58553] = t[58552] ^ n[58553];
assign t[58554] = t[58553] ^ n[58554];
assign t[58555] = t[58554] ^ n[58555];
assign t[58556] = t[58555] ^ n[58556];
assign t[58557] = t[58556] ^ n[58557];
assign t[58558] = t[58557] ^ n[58558];
assign t[58559] = t[58558] ^ n[58559];
assign t[58560] = t[58559] ^ n[58560];
assign t[58561] = t[58560] ^ n[58561];
assign t[58562] = t[58561] ^ n[58562];
assign t[58563] = t[58562] ^ n[58563];
assign t[58564] = t[58563] ^ n[58564];
assign t[58565] = t[58564] ^ n[58565];
assign t[58566] = t[58565] ^ n[58566];
assign t[58567] = t[58566] ^ n[58567];
assign t[58568] = t[58567] ^ n[58568];
assign t[58569] = t[58568] ^ n[58569];
assign t[58570] = t[58569] ^ n[58570];
assign t[58571] = t[58570] ^ n[58571];
assign t[58572] = t[58571] ^ n[58572];
assign t[58573] = t[58572] ^ n[58573];
assign t[58574] = t[58573] ^ n[58574];
assign t[58575] = t[58574] ^ n[58575];
assign t[58576] = t[58575] ^ n[58576];
assign t[58577] = t[58576] ^ n[58577];
assign t[58578] = t[58577] ^ n[58578];
assign t[58579] = t[58578] ^ n[58579];
assign t[58580] = t[58579] ^ n[58580];
assign t[58581] = t[58580] ^ n[58581];
assign t[58582] = t[58581] ^ n[58582];
assign t[58583] = t[58582] ^ n[58583];
assign t[58584] = t[58583] ^ n[58584];
assign t[58585] = t[58584] ^ n[58585];
assign t[58586] = t[58585] ^ n[58586];
assign t[58587] = t[58586] ^ n[58587];
assign t[58588] = t[58587] ^ n[58588];
assign t[58589] = t[58588] ^ n[58589];
assign t[58590] = t[58589] ^ n[58590];
assign t[58591] = t[58590] ^ n[58591];
assign t[58592] = t[58591] ^ n[58592];
assign t[58593] = t[58592] ^ n[58593];
assign t[58594] = t[58593] ^ n[58594];
assign t[58595] = t[58594] ^ n[58595];
assign t[58596] = t[58595] ^ n[58596];
assign t[58597] = t[58596] ^ n[58597];
assign t[58598] = t[58597] ^ n[58598];
assign t[58599] = t[58598] ^ n[58599];
assign t[58600] = t[58599] ^ n[58600];
assign t[58601] = t[58600] ^ n[58601];
assign t[58602] = t[58601] ^ n[58602];
assign t[58603] = t[58602] ^ n[58603];
assign t[58604] = t[58603] ^ n[58604];
assign t[58605] = t[58604] ^ n[58605];
assign t[58606] = t[58605] ^ n[58606];
assign t[58607] = t[58606] ^ n[58607];
assign t[58608] = t[58607] ^ n[58608];
assign t[58609] = t[58608] ^ n[58609];
assign t[58610] = t[58609] ^ n[58610];
assign t[58611] = t[58610] ^ n[58611];
assign t[58612] = t[58611] ^ n[58612];
assign t[58613] = t[58612] ^ n[58613];
assign t[58614] = t[58613] ^ n[58614];
assign t[58615] = t[58614] ^ n[58615];
assign t[58616] = t[58615] ^ n[58616];
assign t[58617] = t[58616] ^ n[58617];
assign t[58618] = t[58617] ^ n[58618];
assign t[58619] = t[58618] ^ n[58619];
assign t[58620] = t[58619] ^ n[58620];
assign t[58621] = t[58620] ^ n[58621];
assign t[58622] = t[58621] ^ n[58622];
assign t[58623] = t[58622] ^ n[58623];
assign t[58624] = t[58623] ^ n[58624];
assign t[58625] = t[58624] ^ n[58625];
assign t[58626] = t[58625] ^ n[58626];
assign t[58627] = t[58626] ^ n[58627];
assign t[58628] = t[58627] ^ n[58628];
assign t[58629] = t[58628] ^ n[58629];
assign t[58630] = t[58629] ^ n[58630];
assign t[58631] = t[58630] ^ n[58631];
assign t[58632] = t[58631] ^ n[58632];
assign t[58633] = t[58632] ^ n[58633];
assign t[58634] = t[58633] ^ n[58634];
assign t[58635] = t[58634] ^ n[58635];
assign t[58636] = t[58635] ^ n[58636];
assign t[58637] = t[58636] ^ n[58637];
assign t[58638] = t[58637] ^ n[58638];
assign t[58639] = t[58638] ^ n[58639];
assign t[58640] = t[58639] ^ n[58640];
assign t[58641] = t[58640] ^ n[58641];
assign t[58642] = t[58641] ^ n[58642];
assign t[58643] = t[58642] ^ n[58643];
assign t[58644] = t[58643] ^ n[58644];
assign t[58645] = t[58644] ^ n[58645];
assign t[58646] = t[58645] ^ n[58646];
assign t[58647] = t[58646] ^ n[58647];
assign t[58648] = t[58647] ^ n[58648];
assign t[58649] = t[58648] ^ n[58649];
assign t[58650] = t[58649] ^ n[58650];
assign t[58651] = t[58650] ^ n[58651];
assign t[58652] = t[58651] ^ n[58652];
assign t[58653] = t[58652] ^ n[58653];
assign t[58654] = t[58653] ^ n[58654];
assign t[58655] = t[58654] ^ n[58655];
assign t[58656] = t[58655] ^ n[58656];
assign t[58657] = t[58656] ^ n[58657];
assign t[58658] = t[58657] ^ n[58658];
assign t[58659] = t[58658] ^ n[58659];
assign t[58660] = t[58659] ^ n[58660];
assign t[58661] = t[58660] ^ n[58661];
assign t[58662] = t[58661] ^ n[58662];
assign t[58663] = t[58662] ^ n[58663];
assign t[58664] = t[58663] ^ n[58664];
assign t[58665] = t[58664] ^ n[58665];
assign t[58666] = t[58665] ^ n[58666];
assign t[58667] = t[58666] ^ n[58667];
assign t[58668] = t[58667] ^ n[58668];
assign t[58669] = t[58668] ^ n[58669];
assign t[58670] = t[58669] ^ n[58670];
assign t[58671] = t[58670] ^ n[58671];
assign t[58672] = t[58671] ^ n[58672];
assign t[58673] = t[58672] ^ n[58673];
assign t[58674] = t[58673] ^ n[58674];
assign t[58675] = t[58674] ^ n[58675];
assign t[58676] = t[58675] ^ n[58676];
assign t[58677] = t[58676] ^ n[58677];
assign t[58678] = t[58677] ^ n[58678];
assign t[58679] = t[58678] ^ n[58679];
assign t[58680] = t[58679] ^ n[58680];
assign t[58681] = t[58680] ^ n[58681];
assign t[58682] = t[58681] ^ n[58682];
assign t[58683] = t[58682] ^ n[58683];
assign t[58684] = t[58683] ^ n[58684];
assign t[58685] = t[58684] ^ n[58685];
assign t[58686] = t[58685] ^ n[58686];
assign t[58687] = t[58686] ^ n[58687];
assign t[58688] = t[58687] ^ n[58688];
assign t[58689] = t[58688] ^ n[58689];
assign t[58690] = t[58689] ^ n[58690];
assign t[58691] = t[58690] ^ n[58691];
assign t[58692] = t[58691] ^ n[58692];
assign t[58693] = t[58692] ^ n[58693];
assign t[58694] = t[58693] ^ n[58694];
assign t[58695] = t[58694] ^ n[58695];
assign t[58696] = t[58695] ^ n[58696];
assign t[58697] = t[58696] ^ n[58697];
assign t[58698] = t[58697] ^ n[58698];
assign t[58699] = t[58698] ^ n[58699];
assign t[58700] = t[58699] ^ n[58700];
assign t[58701] = t[58700] ^ n[58701];
assign t[58702] = t[58701] ^ n[58702];
assign t[58703] = t[58702] ^ n[58703];
assign t[58704] = t[58703] ^ n[58704];
assign t[58705] = t[58704] ^ n[58705];
assign t[58706] = t[58705] ^ n[58706];
assign t[58707] = t[58706] ^ n[58707];
assign t[58708] = t[58707] ^ n[58708];
assign t[58709] = t[58708] ^ n[58709];
assign t[58710] = t[58709] ^ n[58710];
assign t[58711] = t[58710] ^ n[58711];
assign t[58712] = t[58711] ^ n[58712];
assign t[58713] = t[58712] ^ n[58713];
assign t[58714] = t[58713] ^ n[58714];
assign t[58715] = t[58714] ^ n[58715];
assign t[58716] = t[58715] ^ n[58716];
assign t[58717] = t[58716] ^ n[58717];
assign t[58718] = t[58717] ^ n[58718];
assign t[58719] = t[58718] ^ n[58719];
assign t[58720] = t[58719] ^ n[58720];
assign t[58721] = t[58720] ^ n[58721];
assign t[58722] = t[58721] ^ n[58722];
assign t[58723] = t[58722] ^ n[58723];
assign t[58724] = t[58723] ^ n[58724];
assign t[58725] = t[58724] ^ n[58725];
assign t[58726] = t[58725] ^ n[58726];
assign t[58727] = t[58726] ^ n[58727];
assign t[58728] = t[58727] ^ n[58728];
assign t[58729] = t[58728] ^ n[58729];
assign t[58730] = t[58729] ^ n[58730];
assign t[58731] = t[58730] ^ n[58731];
assign t[58732] = t[58731] ^ n[58732];
assign t[58733] = t[58732] ^ n[58733];
assign t[58734] = t[58733] ^ n[58734];
assign t[58735] = t[58734] ^ n[58735];
assign t[58736] = t[58735] ^ n[58736];
assign t[58737] = t[58736] ^ n[58737];
assign t[58738] = t[58737] ^ n[58738];
assign t[58739] = t[58738] ^ n[58739];
assign t[58740] = t[58739] ^ n[58740];
assign t[58741] = t[58740] ^ n[58741];
assign t[58742] = t[58741] ^ n[58742];
assign t[58743] = t[58742] ^ n[58743];
assign t[58744] = t[58743] ^ n[58744];
assign t[58745] = t[58744] ^ n[58745];
assign t[58746] = t[58745] ^ n[58746];
assign t[58747] = t[58746] ^ n[58747];
assign t[58748] = t[58747] ^ n[58748];
assign t[58749] = t[58748] ^ n[58749];
assign t[58750] = t[58749] ^ n[58750];
assign t[58751] = t[58750] ^ n[58751];
assign t[58752] = t[58751] ^ n[58752];
assign t[58753] = t[58752] ^ n[58753];
assign t[58754] = t[58753] ^ n[58754];
assign t[58755] = t[58754] ^ n[58755];
assign t[58756] = t[58755] ^ n[58756];
assign t[58757] = t[58756] ^ n[58757];
assign t[58758] = t[58757] ^ n[58758];
assign t[58759] = t[58758] ^ n[58759];
assign t[58760] = t[58759] ^ n[58760];
assign t[58761] = t[58760] ^ n[58761];
assign t[58762] = t[58761] ^ n[58762];
assign t[58763] = t[58762] ^ n[58763];
assign t[58764] = t[58763] ^ n[58764];
assign t[58765] = t[58764] ^ n[58765];
assign t[58766] = t[58765] ^ n[58766];
assign t[58767] = t[58766] ^ n[58767];
assign t[58768] = t[58767] ^ n[58768];
assign t[58769] = t[58768] ^ n[58769];
assign t[58770] = t[58769] ^ n[58770];
assign t[58771] = t[58770] ^ n[58771];
assign t[58772] = t[58771] ^ n[58772];
assign t[58773] = t[58772] ^ n[58773];
assign t[58774] = t[58773] ^ n[58774];
assign t[58775] = t[58774] ^ n[58775];
assign t[58776] = t[58775] ^ n[58776];
assign t[58777] = t[58776] ^ n[58777];
assign t[58778] = t[58777] ^ n[58778];
assign t[58779] = t[58778] ^ n[58779];
assign t[58780] = t[58779] ^ n[58780];
assign t[58781] = t[58780] ^ n[58781];
assign t[58782] = t[58781] ^ n[58782];
assign t[58783] = t[58782] ^ n[58783];
assign t[58784] = t[58783] ^ n[58784];
assign t[58785] = t[58784] ^ n[58785];
assign t[58786] = t[58785] ^ n[58786];
assign t[58787] = t[58786] ^ n[58787];
assign t[58788] = t[58787] ^ n[58788];
assign t[58789] = t[58788] ^ n[58789];
assign t[58790] = t[58789] ^ n[58790];
assign t[58791] = t[58790] ^ n[58791];
assign t[58792] = t[58791] ^ n[58792];
assign t[58793] = t[58792] ^ n[58793];
assign t[58794] = t[58793] ^ n[58794];
assign t[58795] = t[58794] ^ n[58795];
assign t[58796] = t[58795] ^ n[58796];
assign t[58797] = t[58796] ^ n[58797];
assign t[58798] = t[58797] ^ n[58798];
assign t[58799] = t[58798] ^ n[58799];
assign t[58800] = t[58799] ^ n[58800];
assign t[58801] = t[58800] ^ n[58801];
assign t[58802] = t[58801] ^ n[58802];
assign t[58803] = t[58802] ^ n[58803];
assign t[58804] = t[58803] ^ n[58804];
assign t[58805] = t[58804] ^ n[58805];
assign t[58806] = t[58805] ^ n[58806];
assign t[58807] = t[58806] ^ n[58807];
assign t[58808] = t[58807] ^ n[58808];
assign t[58809] = t[58808] ^ n[58809];
assign t[58810] = t[58809] ^ n[58810];
assign t[58811] = t[58810] ^ n[58811];
assign t[58812] = t[58811] ^ n[58812];
assign t[58813] = t[58812] ^ n[58813];
assign t[58814] = t[58813] ^ n[58814];
assign t[58815] = t[58814] ^ n[58815];
assign t[58816] = t[58815] ^ n[58816];
assign t[58817] = t[58816] ^ n[58817];
assign t[58818] = t[58817] ^ n[58818];
assign t[58819] = t[58818] ^ n[58819];
assign t[58820] = t[58819] ^ n[58820];
assign t[58821] = t[58820] ^ n[58821];
assign t[58822] = t[58821] ^ n[58822];
assign t[58823] = t[58822] ^ n[58823];
assign t[58824] = t[58823] ^ n[58824];
assign t[58825] = t[58824] ^ n[58825];
assign t[58826] = t[58825] ^ n[58826];
assign t[58827] = t[58826] ^ n[58827];
assign t[58828] = t[58827] ^ n[58828];
assign t[58829] = t[58828] ^ n[58829];
assign t[58830] = t[58829] ^ n[58830];
assign t[58831] = t[58830] ^ n[58831];
assign t[58832] = t[58831] ^ n[58832];
assign t[58833] = t[58832] ^ n[58833];
assign t[58834] = t[58833] ^ n[58834];
assign t[58835] = t[58834] ^ n[58835];
assign t[58836] = t[58835] ^ n[58836];
assign t[58837] = t[58836] ^ n[58837];
assign t[58838] = t[58837] ^ n[58838];
assign t[58839] = t[58838] ^ n[58839];
assign t[58840] = t[58839] ^ n[58840];
assign t[58841] = t[58840] ^ n[58841];
assign t[58842] = t[58841] ^ n[58842];
assign t[58843] = t[58842] ^ n[58843];
assign t[58844] = t[58843] ^ n[58844];
assign t[58845] = t[58844] ^ n[58845];
assign t[58846] = t[58845] ^ n[58846];
assign t[58847] = t[58846] ^ n[58847];
assign t[58848] = t[58847] ^ n[58848];
assign t[58849] = t[58848] ^ n[58849];
assign t[58850] = t[58849] ^ n[58850];
assign t[58851] = t[58850] ^ n[58851];
assign t[58852] = t[58851] ^ n[58852];
assign t[58853] = t[58852] ^ n[58853];
assign t[58854] = t[58853] ^ n[58854];
assign t[58855] = t[58854] ^ n[58855];
assign t[58856] = t[58855] ^ n[58856];
assign t[58857] = t[58856] ^ n[58857];
assign t[58858] = t[58857] ^ n[58858];
assign t[58859] = t[58858] ^ n[58859];
assign t[58860] = t[58859] ^ n[58860];
assign t[58861] = t[58860] ^ n[58861];
assign t[58862] = t[58861] ^ n[58862];
assign t[58863] = t[58862] ^ n[58863];
assign t[58864] = t[58863] ^ n[58864];
assign t[58865] = t[58864] ^ n[58865];
assign t[58866] = t[58865] ^ n[58866];
assign t[58867] = t[58866] ^ n[58867];
assign t[58868] = t[58867] ^ n[58868];
assign t[58869] = t[58868] ^ n[58869];
assign t[58870] = t[58869] ^ n[58870];
assign t[58871] = t[58870] ^ n[58871];
assign t[58872] = t[58871] ^ n[58872];
assign t[58873] = t[58872] ^ n[58873];
assign t[58874] = t[58873] ^ n[58874];
assign t[58875] = t[58874] ^ n[58875];
assign t[58876] = t[58875] ^ n[58876];
assign t[58877] = t[58876] ^ n[58877];
assign t[58878] = t[58877] ^ n[58878];
assign t[58879] = t[58878] ^ n[58879];
assign t[58880] = t[58879] ^ n[58880];
assign t[58881] = t[58880] ^ n[58881];
assign t[58882] = t[58881] ^ n[58882];
assign t[58883] = t[58882] ^ n[58883];
assign t[58884] = t[58883] ^ n[58884];
assign t[58885] = t[58884] ^ n[58885];
assign t[58886] = t[58885] ^ n[58886];
assign t[58887] = t[58886] ^ n[58887];
assign t[58888] = t[58887] ^ n[58888];
assign t[58889] = t[58888] ^ n[58889];
assign t[58890] = t[58889] ^ n[58890];
assign t[58891] = t[58890] ^ n[58891];
assign t[58892] = t[58891] ^ n[58892];
assign t[58893] = t[58892] ^ n[58893];
assign t[58894] = t[58893] ^ n[58894];
assign t[58895] = t[58894] ^ n[58895];
assign t[58896] = t[58895] ^ n[58896];
assign t[58897] = t[58896] ^ n[58897];
assign t[58898] = t[58897] ^ n[58898];
assign t[58899] = t[58898] ^ n[58899];
assign t[58900] = t[58899] ^ n[58900];
assign t[58901] = t[58900] ^ n[58901];
assign t[58902] = t[58901] ^ n[58902];
assign t[58903] = t[58902] ^ n[58903];
assign t[58904] = t[58903] ^ n[58904];
assign t[58905] = t[58904] ^ n[58905];
assign t[58906] = t[58905] ^ n[58906];
assign t[58907] = t[58906] ^ n[58907];
assign t[58908] = t[58907] ^ n[58908];
assign t[58909] = t[58908] ^ n[58909];
assign t[58910] = t[58909] ^ n[58910];
assign t[58911] = t[58910] ^ n[58911];
assign t[58912] = t[58911] ^ n[58912];
assign t[58913] = t[58912] ^ n[58913];
assign t[58914] = t[58913] ^ n[58914];
assign t[58915] = t[58914] ^ n[58915];
assign t[58916] = t[58915] ^ n[58916];
assign t[58917] = t[58916] ^ n[58917];
assign t[58918] = t[58917] ^ n[58918];
assign t[58919] = t[58918] ^ n[58919];
assign t[58920] = t[58919] ^ n[58920];
assign t[58921] = t[58920] ^ n[58921];
assign t[58922] = t[58921] ^ n[58922];
assign t[58923] = t[58922] ^ n[58923];
assign t[58924] = t[58923] ^ n[58924];
assign t[58925] = t[58924] ^ n[58925];
assign t[58926] = t[58925] ^ n[58926];
assign t[58927] = t[58926] ^ n[58927];
assign t[58928] = t[58927] ^ n[58928];
assign t[58929] = t[58928] ^ n[58929];
assign t[58930] = t[58929] ^ n[58930];
assign t[58931] = t[58930] ^ n[58931];
assign t[58932] = t[58931] ^ n[58932];
assign t[58933] = t[58932] ^ n[58933];
assign t[58934] = t[58933] ^ n[58934];
assign t[58935] = t[58934] ^ n[58935];
assign t[58936] = t[58935] ^ n[58936];
assign t[58937] = t[58936] ^ n[58937];
assign t[58938] = t[58937] ^ n[58938];
assign t[58939] = t[58938] ^ n[58939];
assign t[58940] = t[58939] ^ n[58940];
assign t[58941] = t[58940] ^ n[58941];
assign t[58942] = t[58941] ^ n[58942];
assign t[58943] = t[58942] ^ n[58943];
assign t[58944] = t[58943] ^ n[58944];
assign t[58945] = t[58944] ^ n[58945];
assign t[58946] = t[58945] ^ n[58946];
assign t[58947] = t[58946] ^ n[58947];
assign t[58948] = t[58947] ^ n[58948];
assign t[58949] = t[58948] ^ n[58949];
assign t[58950] = t[58949] ^ n[58950];
assign t[58951] = t[58950] ^ n[58951];
assign t[58952] = t[58951] ^ n[58952];
assign t[58953] = t[58952] ^ n[58953];
assign t[58954] = t[58953] ^ n[58954];
assign t[58955] = t[58954] ^ n[58955];
assign t[58956] = t[58955] ^ n[58956];
assign t[58957] = t[58956] ^ n[58957];
assign t[58958] = t[58957] ^ n[58958];
assign t[58959] = t[58958] ^ n[58959];
assign t[58960] = t[58959] ^ n[58960];
assign t[58961] = t[58960] ^ n[58961];
assign t[58962] = t[58961] ^ n[58962];
assign t[58963] = t[58962] ^ n[58963];
assign t[58964] = t[58963] ^ n[58964];
assign t[58965] = t[58964] ^ n[58965];
assign t[58966] = t[58965] ^ n[58966];
assign t[58967] = t[58966] ^ n[58967];
assign t[58968] = t[58967] ^ n[58968];
assign t[58969] = t[58968] ^ n[58969];
assign t[58970] = t[58969] ^ n[58970];
assign t[58971] = t[58970] ^ n[58971];
assign t[58972] = t[58971] ^ n[58972];
assign t[58973] = t[58972] ^ n[58973];
assign t[58974] = t[58973] ^ n[58974];
assign t[58975] = t[58974] ^ n[58975];
assign t[58976] = t[58975] ^ n[58976];
assign t[58977] = t[58976] ^ n[58977];
assign t[58978] = t[58977] ^ n[58978];
assign t[58979] = t[58978] ^ n[58979];
assign t[58980] = t[58979] ^ n[58980];
assign t[58981] = t[58980] ^ n[58981];
assign t[58982] = t[58981] ^ n[58982];
assign t[58983] = t[58982] ^ n[58983];
assign t[58984] = t[58983] ^ n[58984];
assign t[58985] = t[58984] ^ n[58985];
assign t[58986] = t[58985] ^ n[58986];
assign t[58987] = t[58986] ^ n[58987];
assign t[58988] = t[58987] ^ n[58988];
assign t[58989] = t[58988] ^ n[58989];
assign t[58990] = t[58989] ^ n[58990];
assign t[58991] = t[58990] ^ n[58991];
assign t[58992] = t[58991] ^ n[58992];
assign t[58993] = t[58992] ^ n[58993];
assign t[58994] = t[58993] ^ n[58994];
assign t[58995] = t[58994] ^ n[58995];
assign t[58996] = t[58995] ^ n[58996];
assign t[58997] = t[58996] ^ n[58997];
assign t[58998] = t[58997] ^ n[58998];
assign t[58999] = t[58998] ^ n[58999];
assign t[59000] = t[58999] ^ n[59000];
assign t[59001] = t[59000] ^ n[59001];
assign t[59002] = t[59001] ^ n[59002];
assign t[59003] = t[59002] ^ n[59003];
assign t[59004] = t[59003] ^ n[59004];
assign t[59005] = t[59004] ^ n[59005];
assign t[59006] = t[59005] ^ n[59006];
assign t[59007] = t[59006] ^ n[59007];
assign t[59008] = t[59007] ^ n[59008];
assign t[59009] = t[59008] ^ n[59009];
assign t[59010] = t[59009] ^ n[59010];
assign t[59011] = t[59010] ^ n[59011];
assign t[59012] = t[59011] ^ n[59012];
assign t[59013] = t[59012] ^ n[59013];
assign t[59014] = t[59013] ^ n[59014];
assign t[59015] = t[59014] ^ n[59015];
assign t[59016] = t[59015] ^ n[59016];
assign t[59017] = t[59016] ^ n[59017];
assign t[59018] = t[59017] ^ n[59018];
assign t[59019] = t[59018] ^ n[59019];
assign t[59020] = t[59019] ^ n[59020];
assign t[59021] = t[59020] ^ n[59021];
assign t[59022] = t[59021] ^ n[59022];
assign t[59023] = t[59022] ^ n[59023];
assign t[59024] = t[59023] ^ n[59024];
assign t[59025] = t[59024] ^ n[59025];
assign t[59026] = t[59025] ^ n[59026];
assign t[59027] = t[59026] ^ n[59027];
assign t[59028] = t[59027] ^ n[59028];
assign t[59029] = t[59028] ^ n[59029];
assign t[59030] = t[59029] ^ n[59030];
assign t[59031] = t[59030] ^ n[59031];
assign t[59032] = t[59031] ^ n[59032];
assign t[59033] = t[59032] ^ n[59033];
assign t[59034] = t[59033] ^ n[59034];
assign t[59035] = t[59034] ^ n[59035];
assign t[59036] = t[59035] ^ n[59036];
assign t[59037] = t[59036] ^ n[59037];
assign t[59038] = t[59037] ^ n[59038];
assign t[59039] = t[59038] ^ n[59039];
assign t[59040] = t[59039] ^ n[59040];
assign t[59041] = t[59040] ^ n[59041];
assign t[59042] = t[59041] ^ n[59042];
assign t[59043] = t[59042] ^ n[59043];
assign t[59044] = t[59043] ^ n[59044];
assign t[59045] = t[59044] ^ n[59045];
assign t[59046] = t[59045] ^ n[59046];
assign t[59047] = t[59046] ^ n[59047];
assign t[59048] = t[59047] ^ n[59048];
assign t[59049] = t[59048] ^ n[59049];
assign t[59050] = t[59049] ^ n[59050];
assign t[59051] = t[59050] ^ n[59051];
assign t[59052] = t[59051] ^ n[59052];
assign t[59053] = t[59052] ^ n[59053];
assign t[59054] = t[59053] ^ n[59054];
assign t[59055] = t[59054] ^ n[59055];
assign t[59056] = t[59055] ^ n[59056];
assign t[59057] = t[59056] ^ n[59057];
assign t[59058] = t[59057] ^ n[59058];
assign t[59059] = t[59058] ^ n[59059];
assign t[59060] = t[59059] ^ n[59060];
assign t[59061] = t[59060] ^ n[59061];
assign t[59062] = t[59061] ^ n[59062];
assign t[59063] = t[59062] ^ n[59063];
assign t[59064] = t[59063] ^ n[59064];
assign t[59065] = t[59064] ^ n[59065];
assign t[59066] = t[59065] ^ n[59066];
assign t[59067] = t[59066] ^ n[59067];
assign t[59068] = t[59067] ^ n[59068];
assign t[59069] = t[59068] ^ n[59069];
assign t[59070] = t[59069] ^ n[59070];
assign t[59071] = t[59070] ^ n[59071];
assign t[59072] = t[59071] ^ n[59072];
assign t[59073] = t[59072] ^ n[59073];
assign t[59074] = t[59073] ^ n[59074];
assign t[59075] = t[59074] ^ n[59075];
assign t[59076] = t[59075] ^ n[59076];
assign t[59077] = t[59076] ^ n[59077];
assign t[59078] = t[59077] ^ n[59078];
assign t[59079] = t[59078] ^ n[59079];
assign t[59080] = t[59079] ^ n[59080];
assign t[59081] = t[59080] ^ n[59081];
assign t[59082] = t[59081] ^ n[59082];
assign t[59083] = t[59082] ^ n[59083];
assign t[59084] = t[59083] ^ n[59084];
assign t[59085] = t[59084] ^ n[59085];
assign t[59086] = t[59085] ^ n[59086];
assign t[59087] = t[59086] ^ n[59087];
assign t[59088] = t[59087] ^ n[59088];
assign t[59089] = t[59088] ^ n[59089];
assign t[59090] = t[59089] ^ n[59090];
assign t[59091] = t[59090] ^ n[59091];
assign t[59092] = t[59091] ^ n[59092];
assign t[59093] = t[59092] ^ n[59093];
assign t[59094] = t[59093] ^ n[59094];
assign t[59095] = t[59094] ^ n[59095];
assign t[59096] = t[59095] ^ n[59096];
assign t[59097] = t[59096] ^ n[59097];
assign t[59098] = t[59097] ^ n[59098];
assign t[59099] = t[59098] ^ n[59099];
assign t[59100] = t[59099] ^ n[59100];
assign t[59101] = t[59100] ^ n[59101];
assign t[59102] = t[59101] ^ n[59102];
assign t[59103] = t[59102] ^ n[59103];
assign t[59104] = t[59103] ^ n[59104];
assign t[59105] = t[59104] ^ n[59105];
assign t[59106] = t[59105] ^ n[59106];
assign t[59107] = t[59106] ^ n[59107];
assign t[59108] = t[59107] ^ n[59108];
assign t[59109] = t[59108] ^ n[59109];
assign t[59110] = t[59109] ^ n[59110];
assign t[59111] = t[59110] ^ n[59111];
assign t[59112] = t[59111] ^ n[59112];
assign t[59113] = t[59112] ^ n[59113];
assign t[59114] = t[59113] ^ n[59114];
assign t[59115] = t[59114] ^ n[59115];
assign t[59116] = t[59115] ^ n[59116];
assign t[59117] = t[59116] ^ n[59117];
assign t[59118] = t[59117] ^ n[59118];
assign t[59119] = t[59118] ^ n[59119];
assign t[59120] = t[59119] ^ n[59120];
assign t[59121] = t[59120] ^ n[59121];
assign t[59122] = t[59121] ^ n[59122];
assign t[59123] = t[59122] ^ n[59123];
assign t[59124] = t[59123] ^ n[59124];
assign t[59125] = t[59124] ^ n[59125];
assign t[59126] = t[59125] ^ n[59126];
assign t[59127] = t[59126] ^ n[59127];
assign t[59128] = t[59127] ^ n[59128];
assign t[59129] = t[59128] ^ n[59129];
assign t[59130] = t[59129] ^ n[59130];
assign t[59131] = t[59130] ^ n[59131];
assign t[59132] = t[59131] ^ n[59132];
assign t[59133] = t[59132] ^ n[59133];
assign t[59134] = t[59133] ^ n[59134];
assign t[59135] = t[59134] ^ n[59135];
assign t[59136] = t[59135] ^ n[59136];
assign t[59137] = t[59136] ^ n[59137];
assign t[59138] = t[59137] ^ n[59138];
assign t[59139] = t[59138] ^ n[59139];
assign t[59140] = t[59139] ^ n[59140];
assign t[59141] = t[59140] ^ n[59141];
assign t[59142] = t[59141] ^ n[59142];
assign t[59143] = t[59142] ^ n[59143];
assign t[59144] = t[59143] ^ n[59144];
assign t[59145] = t[59144] ^ n[59145];
assign t[59146] = t[59145] ^ n[59146];
assign t[59147] = t[59146] ^ n[59147];
assign t[59148] = t[59147] ^ n[59148];
assign t[59149] = t[59148] ^ n[59149];
assign t[59150] = t[59149] ^ n[59150];
assign t[59151] = t[59150] ^ n[59151];
assign t[59152] = t[59151] ^ n[59152];
assign t[59153] = t[59152] ^ n[59153];
assign t[59154] = t[59153] ^ n[59154];
assign t[59155] = t[59154] ^ n[59155];
assign t[59156] = t[59155] ^ n[59156];
assign t[59157] = t[59156] ^ n[59157];
assign t[59158] = t[59157] ^ n[59158];
assign t[59159] = t[59158] ^ n[59159];
assign t[59160] = t[59159] ^ n[59160];
assign t[59161] = t[59160] ^ n[59161];
assign t[59162] = t[59161] ^ n[59162];
assign t[59163] = t[59162] ^ n[59163];
assign t[59164] = t[59163] ^ n[59164];
assign t[59165] = t[59164] ^ n[59165];
assign t[59166] = t[59165] ^ n[59166];
assign t[59167] = t[59166] ^ n[59167];
assign t[59168] = t[59167] ^ n[59168];
assign t[59169] = t[59168] ^ n[59169];
assign t[59170] = t[59169] ^ n[59170];
assign t[59171] = t[59170] ^ n[59171];
assign t[59172] = t[59171] ^ n[59172];
assign t[59173] = t[59172] ^ n[59173];
assign t[59174] = t[59173] ^ n[59174];
assign t[59175] = t[59174] ^ n[59175];
assign t[59176] = t[59175] ^ n[59176];
assign t[59177] = t[59176] ^ n[59177];
assign t[59178] = t[59177] ^ n[59178];
assign t[59179] = t[59178] ^ n[59179];
assign t[59180] = t[59179] ^ n[59180];
assign t[59181] = t[59180] ^ n[59181];
assign t[59182] = t[59181] ^ n[59182];
assign t[59183] = t[59182] ^ n[59183];
assign t[59184] = t[59183] ^ n[59184];
assign t[59185] = t[59184] ^ n[59185];
assign t[59186] = t[59185] ^ n[59186];
assign t[59187] = t[59186] ^ n[59187];
assign t[59188] = t[59187] ^ n[59188];
assign t[59189] = t[59188] ^ n[59189];
assign t[59190] = t[59189] ^ n[59190];
assign t[59191] = t[59190] ^ n[59191];
assign t[59192] = t[59191] ^ n[59192];
assign t[59193] = t[59192] ^ n[59193];
assign t[59194] = t[59193] ^ n[59194];
assign t[59195] = t[59194] ^ n[59195];
assign t[59196] = t[59195] ^ n[59196];
assign t[59197] = t[59196] ^ n[59197];
assign t[59198] = t[59197] ^ n[59198];
assign t[59199] = t[59198] ^ n[59199];
assign t[59200] = t[59199] ^ n[59200];
assign t[59201] = t[59200] ^ n[59201];
assign t[59202] = t[59201] ^ n[59202];
assign t[59203] = t[59202] ^ n[59203];
assign t[59204] = t[59203] ^ n[59204];
assign t[59205] = t[59204] ^ n[59205];
assign t[59206] = t[59205] ^ n[59206];
assign t[59207] = t[59206] ^ n[59207];
assign t[59208] = t[59207] ^ n[59208];
assign t[59209] = t[59208] ^ n[59209];
assign t[59210] = t[59209] ^ n[59210];
assign t[59211] = t[59210] ^ n[59211];
assign t[59212] = t[59211] ^ n[59212];
assign t[59213] = t[59212] ^ n[59213];
assign t[59214] = t[59213] ^ n[59214];
assign t[59215] = t[59214] ^ n[59215];
assign t[59216] = t[59215] ^ n[59216];
assign t[59217] = t[59216] ^ n[59217];
assign t[59218] = t[59217] ^ n[59218];
assign t[59219] = t[59218] ^ n[59219];
assign t[59220] = t[59219] ^ n[59220];
assign t[59221] = t[59220] ^ n[59221];
assign t[59222] = t[59221] ^ n[59222];
assign t[59223] = t[59222] ^ n[59223];
assign t[59224] = t[59223] ^ n[59224];
assign t[59225] = t[59224] ^ n[59225];
assign t[59226] = t[59225] ^ n[59226];
assign t[59227] = t[59226] ^ n[59227];
assign t[59228] = t[59227] ^ n[59228];
assign t[59229] = t[59228] ^ n[59229];
assign t[59230] = t[59229] ^ n[59230];
assign t[59231] = t[59230] ^ n[59231];
assign t[59232] = t[59231] ^ n[59232];
assign t[59233] = t[59232] ^ n[59233];
assign t[59234] = t[59233] ^ n[59234];
assign t[59235] = t[59234] ^ n[59235];
assign t[59236] = t[59235] ^ n[59236];
assign t[59237] = t[59236] ^ n[59237];
assign t[59238] = t[59237] ^ n[59238];
assign t[59239] = t[59238] ^ n[59239];
assign t[59240] = t[59239] ^ n[59240];
assign t[59241] = t[59240] ^ n[59241];
assign t[59242] = t[59241] ^ n[59242];
assign t[59243] = t[59242] ^ n[59243];
assign t[59244] = t[59243] ^ n[59244];
assign t[59245] = t[59244] ^ n[59245];
assign t[59246] = t[59245] ^ n[59246];
assign t[59247] = t[59246] ^ n[59247];
assign t[59248] = t[59247] ^ n[59248];
assign t[59249] = t[59248] ^ n[59249];
assign t[59250] = t[59249] ^ n[59250];
assign t[59251] = t[59250] ^ n[59251];
assign t[59252] = t[59251] ^ n[59252];
assign t[59253] = t[59252] ^ n[59253];
assign t[59254] = t[59253] ^ n[59254];
assign t[59255] = t[59254] ^ n[59255];
assign t[59256] = t[59255] ^ n[59256];
assign t[59257] = t[59256] ^ n[59257];
assign t[59258] = t[59257] ^ n[59258];
assign t[59259] = t[59258] ^ n[59259];
assign t[59260] = t[59259] ^ n[59260];
assign t[59261] = t[59260] ^ n[59261];
assign t[59262] = t[59261] ^ n[59262];
assign t[59263] = t[59262] ^ n[59263];
assign t[59264] = t[59263] ^ n[59264];
assign t[59265] = t[59264] ^ n[59265];
assign t[59266] = t[59265] ^ n[59266];
assign t[59267] = t[59266] ^ n[59267];
assign t[59268] = t[59267] ^ n[59268];
assign t[59269] = t[59268] ^ n[59269];
assign t[59270] = t[59269] ^ n[59270];
assign t[59271] = t[59270] ^ n[59271];
assign t[59272] = t[59271] ^ n[59272];
assign t[59273] = t[59272] ^ n[59273];
assign t[59274] = t[59273] ^ n[59274];
assign t[59275] = t[59274] ^ n[59275];
assign t[59276] = t[59275] ^ n[59276];
assign t[59277] = t[59276] ^ n[59277];
assign t[59278] = t[59277] ^ n[59278];
assign t[59279] = t[59278] ^ n[59279];
assign t[59280] = t[59279] ^ n[59280];
assign t[59281] = t[59280] ^ n[59281];
assign t[59282] = t[59281] ^ n[59282];
assign t[59283] = t[59282] ^ n[59283];
assign t[59284] = t[59283] ^ n[59284];
assign t[59285] = t[59284] ^ n[59285];
assign t[59286] = t[59285] ^ n[59286];
assign t[59287] = t[59286] ^ n[59287];
assign t[59288] = t[59287] ^ n[59288];
assign t[59289] = t[59288] ^ n[59289];
assign t[59290] = t[59289] ^ n[59290];
assign t[59291] = t[59290] ^ n[59291];
assign t[59292] = t[59291] ^ n[59292];
assign t[59293] = t[59292] ^ n[59293];
assign t[59294] = t[59293] ^ n[59294];
assign t[59295] = t[59294] ^ n[59295];
assign t[59296] = t[59295] ^ n[59296];
assign t[59297] = t[59296] ^ n[59297];
assign t[59298] = t[59297] ^ n[59298];
assign t[59299] = t[59298] ^ n[59299];
assign t[59300] = t[59299] ^ n[59300];
assign t[59301] = t[59300] ^ n[59301];
assign t[59302] = t[59301] ^ n[59302];
assign t[59303] = t[59302] ^ n[59303];
assign t[59304] = t[59303] ^ n[59304];
assign t[59305] = t[59304] ^ n[59305];
assign t[59306] = t[59305] ^ n[59306];
assign t[59307] = t[59306] ^ n[59307];
assign t[59308] = t[59307] ^ n[59308];
assign t[59309] = t[59308] ^ n[59309];
assign t[59310] = t[59309] ^ n[59310];
assign t[59311] = t[59310] ^ n[59311];
assign t[59312] = t[59311] ^ n[59312];
assign t[59313] = t[59312] ^ n[59313];
assign t[59314] = t[59313] ^ n[59314];
assign t[59315] = t[59314] ^ n[59315];
assign t[59316] = t[59315] ^ n[59316];
assign t[59317] = t[59316] ^ n[59317];
assign t[59318] = t[59317] ^ n[59318];
assign t[59319] = t[59318] ^ n[59319];
assign t[59320] = t[59319] ^ n[59320];
assign t[59321] = t[59320] ^ n[59321];
assign t[59322] = t[59321] ^ n[59322];
assign t[59323] = t[59322] ^ n[59323];
assign t[59324] = t[59323] ^ n[59324];
assign t[59325] = t[59324] ^ n[59325];
assign t[59326] = t[59325] ^ n[59326];
assign t[59327] = t[59326] ^ n[59327];
assign t[59328] = t[59327] ^ n[59328];
assign t[59329] = t[59328] ^ n[59329];
assign t[59330] = t[59329] ^ n[59330];
assign t[59331] = t[59330] ^ n[59331];
assign t[59332] = t[59331] ^ n[59332];
assign t[59333] = t[59332] ^ n[59333];
assign t[59334] = t[59333] ^ n[59334];
assign t[59335] = t[59334] ^ n[59335];
assign t[59336] = t[59335] ^ n[59336];
assign t[59337] = t[59336] ^ n[59337];
assign t[59338] = t[59337] ^ n[59338];
assign t[59339] = t[59338] ^ n[59339];
assign t[59340] = t[59339] ^ n[59340];
assign t[59341] = t[59340] ^ n[59341];
assign t[59342] = t[59341] ^ n[59342];
assign t[59343] = t[59342] ^ n[59343];
assign t[59344] = t[59343] ^ n[59344];
assign t[59345] = t[59344] ^ n[59345];
assign t[59346] = t[59345] ^ n[59346];
assign t[59347] = t[59346] ^ n[59347];
assign t[59348] = t[59347] ^ n[59348];
assign t[59349] = t[59348] ^ n[59349];
assign t[59350] = t[59349] ^ n[59350];
assign t[59351] = t[59350] ^ n[59351];
assign t[59352] = t[59351] ^ n[59352];
assign t[59353] = t[59352] ^ n[59353];
assign t[59354] = t[59353] ^ n[59354];
assign t[59355] = t[59354] ^ n[59355];
assign t[59356] = t[59355] ^ n[59356];
assign t[59357] = t[59356] ^ n[59357];
assign t[59358] = t[59357] ^ n[59358];
assign t[59359] = t[59358] ^ n[59359];
assign t[59360] = t[59359] ^ n[59360];
assign t[59361] = t[59360] ^ n[59361];
assign t[59362] = t[59361] ^ n[59362];
assign t[59363] = t[59362] ^ n[59363];
assign t[59364] = t[59363] ^ n[59364];
assign t[59365] = t[59364] ^ n[59365];
assign t[59366] = t[59365] ^ n[59366];
assign t[59367] = t[59366] ^ n[59367];
assign t[59368] = t[59367] ^ n[59368];
assign t[59369] = t[59368] ^ n[59369];
assign t[59370] = t[59369] ^ n[59370];
assign t[59371] = t[59370] ^ n[59371];
assign t[59372] = t[59371] ^ n[59372];
assign t[59373] = t[59372] ^ n[59373];
assign t[59374] = t[59373] ^ n[59374];
assign t[59375] = t[59374] ^ n[59375];
assign t[59376] = t[59375] ^ n[59376];
assign t[59377] = t[59376] ^ n[59377];
assign t[59378] = t[59377] ^ n[59378];
assign t[59379] = t[59378] ^ n[59379];
assign t[59380] = t[59379] ^ n[59380];
assign t[59381] = t[59380] ^ n[59381];
assign t[59382] = t[59381] ^ n[59382];
assign t[59383] = t[59382] ^ n[59383];
assign t[59384] = t[59383] ^ n[59384];
assign t[59385] = t[59384] ^ n[59385];
assign t[59386] = t[59385] ^ n[59386];
assign t[59387] = t[59386] ^ n[59387];
assign t[59388] = t[59387] ^ n[59388];
assign t[59389] = t[59388] ^ n[59389];
assign t[59390] = t[59389] ^ n[59390];
assign t[59391] = t[59390] ^ n[59391];
assign t[59392] = t[59391] ^ n[59392];
assign t[59393] = t[59392] ^ n[59393];
assign t[59394] = t[59393] ^ n[59394];
assign t[59395] = t[59394] ^ n[59395];
assign t[59396] = t[59395] ^ n[59396];
assign t[59397] = t[59396] ^ n[59397];
assign t[59398] = t[59397] ^ n[59398];
assign t[59399] = t[59398] ^ n[59399];
assign t[59400] = t[59399] ^ n[59400];
assign t[59401] = t[59400] ^ n[59401];
assign t[59402] = t[59401] ^ n[59402];
assign t[59403] = t[59402] ^ n[59403];
assign t[59404] = t[59403] ^ n[59404];
assign t[59405] = t[59404] ^ n[59405];
assign t[59406] = t[59405] ^ n[59406];
assign t[59407] = t[59406] ^ n[59407];
assign t[59408] = t[59407] ^ n[59408];
assign t[59409] = t[59408] ^ n[59409];
assign t[59410] = t[59409] ^ n[59410];
assign t[59411] = t[59410] ^ n[59411];
assign t[59412] = t[59411] ^ n[59412];
assign t[59413] = t[59412] ^ n[59413];
assign t[59414] = t[59413] ^ n[59414];
assign t[59415] = t[59414] ^ n[59415];
assign t[59416] = t[59415] ^ n[59416];
assign t[59417] = t[59416] ^ n[59417];
assign t[59418] = t[59417] ^ n[59418];
assign t[59419] = t[59418] ^ n[59419];
assign t[59420] = t[59419] ^ n[59420];
assign t[59421] = t[59420] ^ n[59421];
assign t[59422] = t[59421] ^ n[59422];
assign t[59423] = t[59422] ^ n[59423];
assign t[59424] = t[59423] ^ n[59424];
assign t[59425] = t[59424] ^ n[59425];
assign t[59426] = t[59425] ^ n[59426];
assign t[59427] = t[59426] ^ n[59427];
assign t[59428] = t[59427] ^ n[59428];
assign t[59429] = t[59428] ^ n[59429];
assign t[59430] = t[59429] ^ n[59430];
assign t[59431] = t[59430] ^ n[59431];
assign t[59432] = t[59431] ^ n[59432];
assign t[59433] = t[59432] ^ n[59433];
assign t[59434] = t[59433] ^ n[59434];
assign t[59435] = t[59434] ^ n[59435];
assign t[59436] = t[59435] ^ n[59436];
assign t[59437] = t[59436] ^ n[59437];
assign t[59438] = t[59437] ^ n[59438];
assign t[59439] = t[59438] ^ n[59439];
assign t[59440] = t[59439] ^ n[59440];
assign t[59441] = t[59440] ^ n[59441];
assign t[59442] = t[59441] ^ n[59442];
assign t[59443] = t[59442] ^ n[59443];
assign t[59444] = t[59443] ^ n[59444];
assign t[59445] = t[59444] ^ n[59445];
assign t[59446] = t[59445] ^ n[59446];
assign t[59447] = t[59446] ^ n[59447];
assign t[59448] = t[59447] ^ n[59448];
assign t[59449] = t[59448] ^ n[59449];
assign t[59450] = t[59449] ^ n[59450];
assign t[59451] = t[59450] ^ n[59451];
assign t[59452] = t[59451] ^ n[59452];
assign t[59453] = t[59452] ^ n[59453];
assign t[59454] = t[59453] ^ n[59454];
assign t[59455] = t[59454] ^ n[59455];
assign t[59456] = t[59455] ^ n[59456];
assign t[59457] = t[59456] ^ n[59457];
assign t[59458] = t[59457] ^ n[59458];
assign t[59459] = t[59458] ^ n[59459];
assign t[59460] = t[59459] ^ n[59460];
assign t[59461] = t[59460] ^ n[59461];
assign t[59462] = t[59461] ^ n[59462];
assign t[59463] = t[59462] ^ n[59463];
assign t[59464] = t[59463] ^ n[59464];
assign t[59465] = t[59464] ^ n[59465];
assign t[59466] = t[59465] ^ n[59466];
assign t[59467] = t[59466] ^ n[59467];
assign t[59468] = t[59467] ^ n[59468];
assign t[59469] = t[59468] ^ n[59469];
assign t[59470] = t[59469] ^ n[59470];
assign t[59471] = t[59470] ^ n[59471];
assign t[59472] = t[59471] ^ n[59472];
assign t[59473] = t[59472] ^ n[59473];
assign t[59474] = t[59473] ^ n[59474];
assign t[59475] = t[59474] ^ n[59475];
assign t[59476] = t[59475] ^ n[59476];
assign t[59477] = t[59476] ^ n[59477];
assign t[59478] = t[59477] ^ n[59478];
assign t[59479] = t[59478] ^ n[59479];
assign t[59480] = t[59479] ^ n[59480];
assign t[59481] = t[59480] ^ n[59481];
assign t[59482] = t[59481] ^ n[59482];
assign t[59483] = t[59482] ^ n[59483];
assign t[59484] = t[59483] ^ n[59484];
assign t[59485] = t[59484] ^ n[59485];
assign t[59486] = t[59485] ^ n[59486];
assign t[59487] = t[59486] ^ n[59487];
assign t[59488] = t[59487] ^ n[59488];
assign t[59489] = t[59488] ^ n[59489];
assign t[59490] = t[59489] ^ n[59490];
assign t[59491] = t[59490] ^ n[59491];
assign t[59492] = t[59491] ^ n[59492];
assign t[59493] = t[59492] ^ n[59493];
assign t[59494] = t[59493] ^ n[59494];
assign t[59495] = t[59494] ^ n[59495];
assign t[59496] = t[59495] ^ n[59496];
assign t[59497] = t[59496] ^ n[59497];
assign t[59498] = t[59497] ^ n[59498];
assign t[59499] = t[59498] ^ n[59499];
assign t[59500] = t[59499] ^ n[59500];
assign t[59501] = t[59500] ^ n[59501];
assign t[59502] = t[59501] ^ n[59502];
assign t[59503] = t[59502] ^ n[59503];
assign t[59504] = t[59503] ^ n[59504];
assign t[59505] = t[59504] ^ n[59505];
assign t[59506] = t[59505] ^ n[59506];
assign t[59507] = t[59506] ^ n[59507];
assign t[59508] = t[59507] ^ n[59508];
assign t[59509] = t[59508] ^ n[59509];
assign t[59510] = t[59509] ^ n[59510];
assign t[59511] = t[59510] ^ n[59511];
assign t[59512] = t[59511] ^ n[59512];
assign t[59513] = t[59512] ^ n[59513];
assign t[59514] = t[59513] ^ n[59514];
assign t[59515] = t[59514] ^ n[59515];
assign t[59516] = t[59515] ^ n[59516];
assign t[59517] = t[59516] ^ n[59517];
assign t[59518] = t[59517] ^ n[59518];
assign t[59519] = t[59518] ^ n[59519];
assign t[59520] = t[59519] ^ n[59520];
assign t[59521] = t[59520] ^ n[59521];
assign t[59522] = t[59521] ^ n[59522];
assign t[59523] = t[59522] ^ n[59523];
assign t[59524] = t[59523] ^ n[59524];
assign t[59525] = t[59524] ^ n[59525];
assign t[59526] = t[59525] ^ n[59526];
assign t[59527] = t[59526] ^ n[59527];
assign t[59528] = t[59527] ^ n[59528];
assign t[59529] = t[59528] ^ n[59529];
assign t[59530] = t[59529] ^ n[59530];
assign t[59531] = t[59530] ^ n[59531];
assign t[59532] = t[59531] ^ n[59532];
assign t[59533] = t[59532] ^ n[59533];
assign t[59534] = t[59533] ^ n[59534];
assign t[59535] = t[59534] ^ n[59535];
assign t[59536] = t[59535] ^ n[59536];
assign t[59537] = t[59536] ^ n[59537];
assign t[59538] = t[59537] ^ n[59538];
assign t[59539] = t[59538] ^ n[59539];
assign t[59540] = t[59539] ^ n[59540];
assign t[59541] = t[59540] ^ n[59541];
assign t[59542] = t[59541] ^ n[59542];
assign t[59543] = t[59542] ^ n[59543];
assign t[59544] = t[59543] ^ n[59544];
assign t[59545] = t[59544] ^ n[59545];
assign t[59546] = t[59545] ^ n[59546];
assign t[59547] = t[59546] ^ n[59547];
assign t[59548] = t[59547] ^ n[59548];
assign t[59549] = t[59548] ^ n[59549];
assign t[59550] = t[59549] ^ n[59550];
assign t[59551] = t[59550] ^ n[59551];
assign t[59552] = t[59551] ^ n[59552];
assign t[59553] = t[59552] ^ n[59553];
assign t[59554] = t[59553] ^ n[59554];
assign t[59555] = t[59554] ^ n[59555];
assign t[59556] = t[59555] ^ n[59556];
assign t[59557] = t[59556] ^ n[59557];
assign t[59558] = t[59557] ^ n[59558];
assign t[59559] = t[59558] ^ n[59559];
assign t[59560] = t[59559] ^ n[59560];
assign t[59561] = t[59560] ^ n[59561];
assign t[59562] = t[59561] ^ n[59562];
assign t[59563] = t[59562] ^ n[59563];
assign t[59564] = t[59563] ^ n[59564];
assign t[59565] = t[59564] ^ n[59565];
assign t[59566] = t[59565] ^ n[59566];
assign t[59567] = t[59566] ^ n[59567];
assign t[59568] = t[59567] ^ n[59568];
assign t[59569] = t[59568] ^ n[59569];
assign t[59570] = t[59569] ^ n[59570];
assign t[59571] = t[59570] ^ n[59571];
assign t[59572] = t[59571] ^ n[59572];
assign t[59573] = t[59572] ^ n[59573];
assign t[59574] = t[59573] ^ n[59574];
assign t[59575] = t[59574] ^ n[59575];
assign t[59576] = t[59575] ^ n[59576];
assign t[59577] = t[59576] ^ n[59577];
assign t[59578] = t[59577] ^ n[59578];
assign t[59579] = t[59578] ^ n[59579];
assign t[59580] = t[59579] ^ n[59580];
assign t[59581] = t[59580] ^ n[59581];
assign t[59582] = t[59581] ^ n[59582];
assign t[59583] = t[59582] ^ n[59583];
assign t[59584] = t[59583] ^ n[59584];
assign t[59585] = t[59584] ^ n[59585];
assign t[59586] = t[59585] ^ n[59586];
assign t[59587] = t[59586] ^ n[59587];
assign t[59588] = t[59587] ^ n[59588];
assign t[59589] = t[59588] ^ n[59589];
assign t[59590] = t[59589] ^ n[59590];
assign t[59591] = t[59590] ^ n[59591];
assign t[59592] = t[59591] ^ n[59592];
assign t[59593] = t[59592] ^ n[59593];
assign t[59594] = t[59593] ^ n[59594];
assign t[59595] = t[59594] ^ n[59595];
assign t[59596] = t[59595] ^ n[59596];
assign t[59597] = t[59596] ^ n[59597];
assign t[59598] = t[59597] ^ n[59598];
assign t[59599] = t[59598] ^ n[59599];
assign t[59600] = t[59599] ^ n[59600];
assign t[59601] = t[59600] ^ n[59601];
assign t[59602] = t[59601] ^ n[59602];
assign t[59603] = t[59602] ^ n[59603];
assign t[59604] = t[59603] ^ n[59604];
assign t[59605] = t[59604] ^ n[59605];
assign t[59606] = t[59605] ^ n[59606];
assign t[59607] = t[59606] ^ n[59607];
assign t[59608] = t[59607] ^ n[59608];
assign t[59609] = t[59608] ^ n[59609];
assign t[59610] = t[59609] ^ n[59610];
assign t[59611] = t[59610] ^ n[59611];
assign t[59612] = t[59611] ^ n[59612];
assign t[59613] = t[59612] ^ n[59613];
assign t[59614] = t[59613] ^ n[59614];
assign t[59615] = t[59614] ^ n[59615];
assign t[59616] = t[59615] ^ n[59616];
assign t[59617] = t[59616] ^ n[59617];
assign t[59618] = t[59617] ^ n[59618];
assign t[59619] = t[59618] ^ n[59619];
assign t[59620] = t[59619] ^ n[59620];
assign t[59621] = t[59620] ^ n[59621];
assign t[59622] = t[59621] ^ n[59622];
assign t[59623] = t[59622] ^ n[59623];
assign t[59624] = t[59623] ^ n[59624];
assign t[59625] = t[59624] ^ n[59625];
assign t[59626] = t[59625] ^ n[59626];
assign t[59627] = t[59626] ^ n[59627];
assign t[59628] = t[59627] ^ n[59628];
assign t[59629] = t[59628] ^ n[59629];
assign t[59630] = t[59629] ^ n[59630];
assign t[59631] = t[59630] ^ n[59631];
assign t[59632] = t[59631] ^ n[59632];
assign t[59633] = t[59632] ^ n[59633];
assign t[59634] = t[59633] ^ n[59634];
assign t[59635] = t[59634] ^ n[59635];
assign t[59636] = t[59635] ^ n[59636];
assign t[59637] = t[59636] ^ n[59637];
assign t[59638] = t[59637] ^ n[59638];
assign t[59639] = t[59638] ^ n[59639];
assign t[59640] = t[59639] ^ n[59640];
assign t[59641] = t[59640] ^ n[59641];
assign t[59642] = t[59641] ^ n[59642];
assign t[59643] = t[59642] ^ n[59643];
assign t[59644] = t[59643] ^ n[59644];
assign t[59645] = t[59644] ^ n[59645];
assign t[59646] = t[59645] ^ n[59646];
assign t[59647] = t[59646] ^ n[59647];
assign t[59648] = t[59647] ^ n[59648];
assign t[59649] = t[59648] ^ n[59649];
assign t[59650] = t[59649] ^ n[59650];
assign t[59651] = t[59650] ^ n[59651];
assign t[59652] = t[59651] ^ n[59652];
assign t[59653] = t[59652] ^ n[59653];
assign t[59654] = t[59653] ^ n[59654];
assign t[59655] = t[59654] ^ n[59655];
assign t[59656] = t[59655] ^ n[59656];
assign t[59657] = t[59656] ^ n[59657];
assign t[59658] = t[59657] ^ n[59658];
assign t[59659] = t[59658] ^ n[59659];
assign t[59660] = t[59659] ^ n[59660];
assign t[59661] = t[59660] ^ n[59661];
assign t[59662] = t[59661] ^ n[59662];
assign t[59663] = t[59662] ^ n[59663];
assign t[59664] = t[59663] ^ n[59664];
assign t[59665] = t[59664] ^ n[59665];
assign t[59666] = t[59665] ^ n[59666];
assign t[59667] = t[59666] ^ n[59667];
assign t[59668] = t[59667] ^ n[59668];
assign t[59669] = t[59668] ^ n[59669];
assign t[59670] = t[59669] ^ n[59670];
assign t[59671] = t[59670] ^ n[59671];
assign t[59672] = t[59671] ^ n[59672];
assign t[59673] = t[59672] ^ n[59673];
assign t[59674] = t[59673] ^ n[59674];
assign t[59675] = t[59674] ^ n[59675];
assign t[59676] = t[59675] ^ n[59676];
assign t[59677] = t[59676] ^ n[59677];
assign t[59678] = t[59677] ^ n[59678];
assign t[59679] = t[59678] ^ n[59679];
assign t[59680] = t[59679] ^ n[59680];
assign t[59681] = t[59680] ^ n[59681];
assign t[59682] = t[59681] ^ n[59682];
assign t[59683] = t[59682] ^ n[59683];
assign t[59684] = t[59683] ^ n[59684];
assign t[59685] = t[59684] ^ n[59685];
assign t[59686] = t[59685] ^ n[59686];
assign t[59687] = t[59686] ^ n[59687];
assign t[59688] = t[59687] ^ n[59688];
assign t[59689] = t[59688] ^ n[59689];
assign t[59690] = t[59689] ^ n[59690];
assign t[59691] = t[59690] ^ n[59691];
assign t[59692] = t[59691] ^ n[59692];
assign t[59693] = t[59692] ^ n[59693];
assign t[59694] = t[59693] ^ n[59694];
assign t[59695] = t[59694] ^ n[59695];
assign t[59696] = t[59695] ^ n[59696];
assign t[59697] = t[59696] ^ n[59697];
assign t[59698] = t[59697] ^ n[59698];
assign t[59699] = t[59698] ^ n[59699];
assign t[59700] = t[59699] ^ n[59700];
assign t[59701] = t[59700] ^ n[59701];
assign t[59702] = t[59701] ^ n[59702];
assign t[59703] = t[59702] ^ n[59703];
assign t[59704] = t[59703] ^ n[59704];
assign t[59705] = t[59704] ^ n[59705];
assign t[59706] = t[59705] ^ n[59706];
assign t[59707] = t[59706] ^ n[59707];
assign t[59708] = t[59707] ^ n[59708];
assign t[59709] = t[59708] ^ n[59709];
assign t[59710] = t[59709] ^ n[59710];
assign t[59711] = t[59710] ^ n[59711];
assign t[59712] = t[59711] ^ n[59712];
assign t[59713] = t[59712] ^ n[59713];
assign t[59714] = t[59713] ^ n[59714];
assign t[59715] = t[59714] ^ n[59715];
assign t[59716] = t[59715] ^ n[59716];
assign t[59717] = t[59716] ^ n[59717];
assign t[59718] = t[59717] ^ n[59718];
assign t[59719] = t[59718] ^ n[59719];
assign t[59720] = t[59719] ^ n[59720];
assign t[59721] = t[59720] ^ n[59721];
assign t[59722] = t[59721] ^ n[59722];
assign t[59723] = t[59722] ^ n[59723];
assign t[59724] = t[59723] ^ n[59724];
assign t[59725] = t[59724] ^ n[59725];
assign t[59726] = t[59725] ^ n[59726];
assign t[59727] = t[59726] ^ n[59727];
assign t[59728] = t[59727] ^ n[59728];
assign t[59729] = t[59728] ^ n[59729];
assign t[59730] = t[59729] ^ n[59730];
assign t[59731] = t[59730] ^ n[59731];
assign t[59732] = t[59731] ^ n[59732];
assign t[59733] = t[59732] ^ n[59733];
assign t[59734] = t[59733] ^ n[59734];
assign t[59735] = t[59734] ^ n[59735];
assign t[59736] = t[59735] ^ n[59736];
assign t[59737] = t[59736] ^ n[59737];
assign t[59738] = t[59737] ^ n[59738];
assign t[59739] = t[59738] ^ n[59739];
assign t[59740] = t[59739] ^ n[59740];
assign t[59741] = t[59740] ^ n[59741];
assign t[59742] = t[59741] ^ n[59742];
assign t[59743] = t[59742] ^ n[59743];
assign t[59744] = t[59743] ^ n[59744];
assign t[59745] = t[59744] ^ n[59745];
assign t[59746] = t[59745] ^ n[59746];
assign t[59747] = t[59746] ^ n[59747];
assign t[59748] = t[59747] ^ n[59748];
assign t[59749] = t[59748] ^ n[59749];
assign t[59750] = t[59749] ^ n[59750];
assign t[59751] = t[59750] ^ n[59751];
assign t[59752] = t[59751] ^ n[59752];
assign t[59753] = t[59752] ^ n[59753];
assign t[59754] = t[59753] ^ n[59754];
assign t[59755] = t[59754] ^ n[59755];
assign t[59756] = t[59755] ^ n[59756];
assign t[59757] = t[59756] ^ n[59757];
assign t[59758] = t[59757] ^ n[59758];
assign t[59759] = t[59758] ^ n[59759];
assign t[59760] = t[59759] ^ n[59760];
assign t[59761] = t[59760] ^ n[59761];
assign t[59762] = t[59761] ^ n[59762];
assign t[59763] = t[59762] ^ n[59763];
assign t[59764] = t[59763] ^ n[59764];
assign t[59765] = t[59764] ^ n[59765];
assign t[59766] = t[59765] ^ n[59766];
assign t[59767] = t[59766] ^ n[59767];
assign t[59768] = t[59767] ^ n[59768];
assign t[59769] = t[59768] ^ n[59769];
assign t[59770] = t[59769] ^ n[59770];
assign t[59771] = t[59770] ^ n[59771];
assign t[59772] = t[59771] ^ n[59772];
assign t[59773] = t[59772] ^ n[59773];
assign t[59774] = t[59773] ^ n[59774];
assign t[59775] = t[59774] ^ n[59775];
assign t[59776] = t[59775] ^ n[59776];
assign t[59777] = t[59776] ^ n[59777];
assign t[59778] = t[59777] ^ n[59778];
assign t[59779] = t[59778] ^ n[59779];
assign t[59780] = t[59779] ^ n[59780];
assign t[59781] = t[59780] ^ n[59781];
assign t[59782] = t[59781] ^ n[59782];
assign t[59783] = t[59782] ^ n[59783];
assign t[59784] = t[59783] ^ n[59784];
assign t[59785] = t[59784] ^ n[59785];
assign t[59786] = t[59785] ^ n[59786];
assign t[59787] = t[59786] ^ n[59787];
assign t[59788] = t[59787] ^ n[59788];
assign t[59789] = t[59788] ^ n[59789];
assign t[59790] = t[59789] ^ n[59790];
assign t[59791] = t[59790] ^ n[59791];
assign t[59792] = t[59791] ^ n[59792];
assign t[59793] = t[59792] ^ n[59793];
assign t[59794] = t[59793] ^ n[59794];
assign t[59795] = t[59794] ^ n[59795];
assign t[59796] = t[59795] ^ n[59796];
assign t[59797] = t[59796] ^ n[59797];
assign t[59798] = t[59797] ^ n[59798];
assign t[59799] = t[59798] ^ n[59799];
assign t[59800] = t[59799] ^ n[59800];
assign t[59801] = t[59800] ^ n[59801];
assign t[59802] = t[59801] ^ n[59802];
assign t[59803] = t[59802] ^ n[59803];
assign t[59804] = t[59803] ^ n[59804];
assign t[59805] = t[59804] ^ n[59805];
assign t[59806] = t[59805] ^ n[59806];
assign t[59807] = t[59806] ^ n[59807];
assign t[59808] = t[59807] ^ n[59808];
assign t[59809] = t[59808] ^ n[59809];
assign t[59810] = t[59809] ^ n[59810];
assign t[59811] = t[59810] ^ n[59811];
assign t[59812] = t[59811] ^ n[59812];
assign t[59813] = t[59812] ^ n[59813];
assign t[59814] = t[59813] ^ n[59814];
assign t[59815] = t[59814] ^ n[59815];
assign t[59816] = t[59815] ^ n[59816];
assign t[59817] = t[59816] ^ n[59817];
assign t[59818] = t[59817] ^ n[59818];
assign t[59819] = t[59818] ^ n[59819];
assign t[59820] = t[59819] ^ n[59820];
assign t[59821] = t[59820] ^ n[59821];
assign t[59822] = t[59821] ^ n[59822];
assign t[59823] = t[59822] ^ n[59823];
assign t[59824] = t[59823] ^ n[59824];
assign t[59825] = t[59824] ^ n[59825];
assign t[59826] = t[59825] ^ n[59826];
assign t[59827] = t[59826] ^ n[59827];
assign t[59828] = t[59827] ^ n[59828];
assign t[59829] = t[59828] ^ n[59829];
assign t[59830] = t[59829] ^ n[59830];
assign t[59831] = t[59830] ^ n[59831];
assign t[59832] = t[59831] ^ n[59832];
assign t[59833] = t[59832] ^ n[59833];
assign t[59834] = t[59833] ^ n[59834];
assign t[59835] = t[59834] ^ n[59835];
assign t[59836] = t[59835] ^ n[59836];
assign t[59837] = t[59836] ^ n[59837];
assign t[59838] = t[59837] ^ n[59838];
assign t[59839] = t[59838] ^ n[59839];
assign t[59840] = t[59839] ^ n[59840];
assign t[59841] = t[59840] ^ n[59841];
assign t[59842] = t[59841] ^ n[59842];
assign t[59843] = t[59842] ^ n[59843];
assign t[59844] = t[59843] ^ n[59844];
assign t[59845] = t[59844] ^ n[59845];
assign t[59846] = t[59845] ^ n[59846];
assign t[59847] = t[59846] ^ n[59847];
assign t[59848] = t[59847] ^ n[59848];
assign t[59849] = t[59848] ^ n[59849];
assign t[59850] = t[59849] ^ n[59850];
assign t[59851] = t[59850] ^ n[59851];
assign t[59852] = t[59851] ^ n[59852];
assign t[59853] = t[59852] ^ n[59853];
assign t[59854] = t[59853] ^ n[59854];
assign t[59855] = t[59854] ^ n[59855];
assign t[59856] = t[59855] ^ n[59856];
assign t[59857] = t[59856] ^ n[59857];
assign t[59858] = t[59857] ^ n[59858];
assign t[59859] = t[59858] ^ n[59859];
assign t[59860] = t[59859] ^ n[59860];
assign t[59861] = t[59860] ^ n[59861];
assign t[59862] = t[59861] ^ n[59862];
assign t[59863] = t[59862] ^ n[59863];
assign t[59864] = t[59863] ^ n[59864];
assign t[59865] = t[59864] ^ n[59865];
assign t[59866] = t[59865] ^ n[59866];
assign t[59867] = t[59866] ^ n[59867];
assign t[59868] = t[59867] ^ n[59868];
assign t[59869] = t[59868] ^ n[59869];
assign t[59870] = t[59869] ^ n[59870];
assign t[59871] = t[59870] ^ n[59871];
assign t[59872] = t[59871] ^ n[59872];
assign t[59873] = t[59872] ^ n[59873];
assign t[59874] = t[59873] ^ n[59874];
assign t[59875] = t[59874] ^ n[59875];
assign t[59876] = t[59875] ^ n[59876];
assign t[59877] = t[59876] ^ n[59877];
assign t[59878] = t[59877] ^ n[59878];
assign t[59879] = t[59878] ^ n[59879];
assign t[59880] = t[59879] ^ n[59880];
assign t[59881] = t[59880] ^ n[59881];
assign t[59882] = t[59881] ^ n[59882];
assign t[59883] = t[59882] ^ n[59883];
assign t[59884] = t[59883] ^ n[59884];
assign t[59885] = t[59884] ^ n[59885];
assign t[59886] = t[59885] ^ n[59886];
assign t[59887] = t[59886] ^ n[59887];
assign t[59888] = t[59887] ^ n[59888];
assign t[59889] = t[59888] ^ n[59889];
assign t[59890] = t[59889] ^ n[59890];
assign t[59891] = t[59890] ^ n[59891];
assign t[59892] = t[59891] ^ n[59892];
assign t[59893] = t[59892] ^ n[59893];
assign t[59894] = t[59893] ^ n[59894];
assign t[59895] = t[59894] ^ n[59895];
assign t[59896] = t[59895] ^ n[59896];
assign t[59897] = t[59896] ^ n[59897];
assign t[59898] = t[59897] ^ n[59898];
assign t[59899] = t[59898] ^ n[59899];
assign t[59900] = t[59899] ^ n[59900];
assign t[59901] = t[59900] ^ n[59901];
assign t[59902] = t[59901] ^ n[59902];
assign t[59903] = t[59902] ^ n[59903];
assign t[59904] = t[59903] ^ n[59904];
assign t[59905] = t[59904] ^ n[59905];
assign t[59906] = t[59905] ^ n[59906];
assign t[59907] = t[59906] ^ n[59907];
assign t[59908] = t[59907] ^ n[59908];
assign t[59909] = t[59908] ^ n[59909];
assign t[59910] = t[59909] ^ n[59910];
assign t[59911] = t[59910] ^ n[59911];
assign t[59912] = t[59911] ^ n[59912];
assign t[59913] = t[59912] ^ n[59913];
assign t[59914] = t[59913] ^ n[59914];
assign t[59915] = t[59914] ^ n[59915];
assign t[59916] = t[59915] ^ n[59916];
assign t[59917] = t[59916] ^ n[59917];
assign t[59918] = t[59917] ^ n[59918];
assign t[59919] = t[59918] ^ n[59919];
assign t[59920] = t[59919] ^ n[59920];
assign t[59921] = t[59920] ^ n[59921];
assign t[59922] = t[59921] ^ n[59922];
assign t[59923] = t[59922] ^ n[59923];
assign t[59924] = t[59923] ^ n[59924];
assign t[59925] = t[59924] ^ n[59925];
assign t[59926] = t[59925] ^ n[59926];
assign t[59927] = t[59926] ^ n[59927];
assign t[59928] = t[59927] ^ n[59928];
assign t[59929] = t[59928] ^ n[59929];
assign t[59930] = t[59929] ^ n[59930];
assign t[59931] = t[59930] ^ n[59931];
assign t[59932] = t[59931] ^ n[59932];
assign t[59933] = t[59932] ^ n[59933];
assign t[59934] = t[59933] ^ n[59934];
assign t[59935] = t[59934] ^ n[59935];
assign t[59936] = t[59935] ^ n[59936];
assign t[59937] = t[59936] ^ n[59937];
assign t[59938] = t[59937] ^ n[59938];
assign t[59939] = t[59938] ^ n[59939];
assign t[59940] = t[59939] ^ n[59940];
assign t[59941] = t[59940] ^ n[59941];
assign t[59942] = t[59941] ^ n[59942];
assign t[59943] = t[59942] ^ n[59943];
assign t[59944] = t[59943] ^ n[59944];
assign t[59945] = t[59944] ^ n[59945];
assign t[59946] = t[59945] ^ n[59946];
assign t[59947] = t[59946] ^ n[59947];
assign t[59948] = t[59947] ^ n[59948];
assign t[59949] = t[59948] ^ n[59949];
assign t[59950] = t[59949] ^ n[59950];
assign t[59951] = t[59950] ^ n[59951];
assign t[59952] = t[59951] ^ n[59952];
assign t[59953] = t[59952] ^ n[59953];
assign t[59954] = t[59953] ^ n[59954];
assign t[59955] = t[59954] ^ n[59955];
assign t[59956] = t[59955] ^ n[59956];
assign t[59957] = t[59956] ^ n[59957];
assign t[59958] = t[59957] ^ n[59958];
assign t[59959] = t[59958] ^ n[59959];
assign t[59960] = t[59959] ^ n[59960];
assign t[59961] = t[59960] ^ n[59961];
assign t[59962] = t[59961] ^ n[59962];
assign t[59963] = t[59962] ^ n[59963];
assign t[59964] = t[59963] ^ n[59964];
assign t[59965] = t[59964] ^ n[59965];
assign t[59966] = t[59965] ^ n[59966];
assign t[59967] = t[59966] ^ n[59967];
assign t[59968] = t[59967] ^ n[59968];
assign t[59969] = t[59968] ^ n[59969];
assign t[59970] = t[59969] ^ n[59970];
assign t[59971] = t[59970] ^ n[59971];
assign t[59972] = t[59971] ^ n[59972];
assign t[59973] = t[59972] ^ n[59973];
assign t[59974] = t[59973] ^ n[59974];
assign t[59975] = t[59974] ^ n[59975];
assign t[59976] = t[59975] ^ n[59976];
assign t[59977] = t[59976] ^ n[59977];
assign t[59978] = t[59977] ^ n[59978];
assign t[59979] = t[59978] ^ n[59979];
assign t[59980] = t[59979] ^ n[59980];
assign t[59981] = t[59980] ^ n[59981];
assign t[59982] = t[59981] ^ n[59982];
assign t[59983] = t[59982] ^ n[59983];
assign t[59984] = t[59983] ^ n[59984];
assign t[59985] = t[59984] ^ n[59985];
assign t[59986] = t[59985] ^ n[59986];
assign t[59987] = t[59986] ^ n[59987];
assign t[59988] = t[59987] ^ n[59988];
assign t[59989] = t[59988] ^ n[59989];
assign t[59990] = t[59989] ^ n[59990];
assign t[59991] = t[59990] ^ n[59991];
assign t[59992] = t[59991] ^ n[59992];
assign t[59993] = t[59992] ^ n[59993];
assign t[59994] = t[59993] ^ n[59994];
assign t[59995] = t[59994] ^ n[59995];
assign t[59996] = t[59995] ^ n[59996];
assign t[59997] = t[59996] ^ n[59997];
assign t[59998] = t[59997] ^ n[59998];
assign t[59999] = t[59998] ^ n[59999];
assign t[60000] = t[59999] ^ n[60000];
assign t[60001] = t[60000] ^ n[60001];
assign t[60002] = t[60001] ^ n[60002];
assign t[60003] = t[60002] ^ n[60003];
assign t[60004] = t[60003] ^ n[60004];
assign t[60005] = t[60004] ^ n[60005];
assign t[60006] = t[60005] ^ n[60006];
assign t[60007] = t[60006] ^ n[60007];
assign t[60008] = t[60007] ^ n[60008];
assign t[60009] = t[60008] ^ n[60009];
assign t[60010] = t[60009] ^ n[60010];
assign t[60011] = t[60010] ^ n[60011];
assign t[60012] = t[60011] ^ n[60012];
assign t[60013] = t[60012] ^ n[60013];
assign t[60014] = t[60013] ^ n[60014];
assign t[60015] = t[60014] ^ n[60015];
assign t[60016] = t[60015] ^ n[60016];
assign t[60017] = t[60016] ^ n[60017];
assign t[60018] = t[60017] ^ n[60018];
assign t[60019] = t[60018] ^ n[60019];
assign t[60020] = t[60019] ^ n[60020];
assign t[60021] = t[60020] ^ n[60021];
assign t[60022] = t[60021] ^ n[60022];
assign t[60023] = t[60022] ^ n[60023];
assign t[60024] = t[60023] ^ n[60024];
assign t[60025] = t[60024] ^ n[60025];
assign t[60026] = t[60025] ^ n[60026];
assign t[60027] = t[60026] ^ n[60027];
assign t[60028] = t[60027] ^ n[60028];
assign t[60029] = t[60028] ^ n[60029];
assign t[60030] = t[60029] ^ n[60030];
assign t[60031] = t[60030] ^ n[60031];
assign t[60032] = t[60031] ^ n[60032];
assign t[60033] = t[60032] ^ n[60033];
assign t[60034] = t[60033] ^ n[60034];
assign t[60035] = t[60034] ^ n[60035];
assign t[60036] = t[60035] ^ n[60036];
assign t[60037] = t[60036] ^ n[60037];
assign t[60038] = t[60037] ^ n[60038];
assign t[60039] = t[60038] ^ n[60039];
assign t[60040] = t[60039] ^ n[60040];
assign t[60041] = t[60040] ^ n[60041];
assign t[60042] = t[60041] ^ n[60042];
assign t[60043] = t[60042] ^ n[60043];
assign t[60044] = t[60043] ^ n[60044];
assign t[60045] = t[60044] ^ n[60045];
assign t[60046] = t[60045] ^ n[60046];
assign t[60047] = t[60046] ^ n[60047];
assign t[60048] = t[60047] ^ n[60048];
assign t[60049] = t[60048] ^ n[60049];
assign t[60050] = t[60049] ^ n[60050];
assign t[60051] = t[60050] ^ n[60051];
assign t[60052] = t[60051] ^ n[60052];
assign t[60053] = t[60052] ^ n[60053];
assign t[60054] = t[60053] ^ n[60054];
assign t[60055] = t[60054] ^ n[60055];
assign t[60056] = t[60055] ^ n[60056];
assign t[60057] = t[60056] ^ n[60057];
assign t[60058] = t[60057] ^ n[60058];
assign t[60059] = t[60058] ^ n[60059];
assign t[60060] = t[60059] ^ n[60060];
assign t[60061] = t[60060] ^ n[60061];
assign t[60062] = t[60061] ^ n[60062];
assign t[60063] = t[60062] ^ n[60063];
assign t[60064] = t[60063] ^ n[60064];
assign t[60065] = t[60064] ^ n[60065];
assign t[60066] = t[60065] ^ n[60066];
assign t[60067] = t[60066] ^ n[60067];
assign t[60068] = t[60067] ^ n[60068];
assign t[60069] = t[60068] ^ n[60069];
assign t[60070] = t[60069] ^ n[60070];
assign t[60071] = t[60070] ^ n[60071];
assign t[60072] = t[60071] ^ n[60072];
assign t[60073] = t[60072] ^ n[60073];
assign t[60074] = t[60073] ^ n[60074];
assign t[60075] = t[60074] ^ n[60075];
assign t[60076] = t[60075] ^ n[60076];
assign t[60077] = t[60076] ^ n[60077];
assign t[60078] = t[60077] ^ n[60078];
assign t[60079] = t[60078] ^ n[60079];
assign t[60080] = t[60079] ^ n[60080];
assign t[60081] = t[60080] ^ n[60081];
assign t[60082] = t[60081] ^ n[60082];
assign t[60083] = t[60082] ^ n[60083];
assign t[60084] = t[60083] ^ n[60084];
assign t[60085] = t[60084] ^ n[60085];
assign t[60086] = t[60085] ^ n[60086];
assign t[60087] = t[60086] ^ n[60087];
assign t[60088] = t[60087] ^ n[60088];
assign t[60089] = t[60088] ^ n[60089];
assign t[60090] = t[60089] ^ n[60090];
assign t[60091] = t[60090] ^ n[60091];
assign t[60092] = t[60091] ^ n[60092];
assign t[60093] = t[60092] ^ n[60093];
assign t[60094] = t[60093] ^ n[60094];
assign t[60095] = t[60094] ^ n[60095];
assign t[60096] = t[60095] ^ n[60096];
assign t[60097] = t[60096] ^ n[60097];
assign t[60098] = t[60097] ^ n[60098];
assign t[60099] = t[60098] ^ n[60099];
assign t[60100] = t[60099] ^ n[60100];
assign t[60101] = t[60100] ^ n[60101];
assign t[60102] = t[60101] ^ n[60102];
assign t[60103] = t[60102] ^ n[60103];
assign t[60104] = t[60103] ^ n[60104];
assign t[60105] = t[60104] ^ n[60105];
assign t[60106] = t[60105] ^ n[60106];
assign t[60107] = t[60106] ^ n[60107];
assign t[60108] = t[60107] ^ n[60108];
assign t[60109] = t[60108] ^ n[60109];
assign t[60110] = t[60109] ^ n[60110];
assign t[60111] = t[60110] ^ n[60111];
assign t[60112] = t[60111] ^ n[60112];
assign t[60113] = t[60112] ^ n[60113];
assign t[60114] = t[60113] ^ n[60114];
assign t[60115] = t[60114] ^ n[60115];
assign t[60116] = t[60115] ^ n[60116];
assign t[60117] = t[60116] ^ n[60117];
assign t[60118] = t[60117] ^ n[60118];
assign t[60119] = t[60118] ^ n[60119];
assign t[60120] = t[60119] ^ n[60120];
assign t[60121] = t[60120] ^ n[60121];
assign t[60122] = t[60121] ^ n[60122];
assign t[60123] = t[60122] ^ n[60123];
assign t[60124] = t[60123] ^ n[60124];
assign t[60125] = t[60124] ^ n[60125];
assign t[60126] = t[60125] ^ n[60126];
assign t[60127] = t[60126] ^ n[60127];
assign t[60128] = t[60127] ^ n[60128];
assign t[60129] = t[60128] ^ n[60129];
assign t[60130] = t[60129] ^ n[60130];
assign t[60131] = t[60130] ^ n[60131];
assign t[60132] = t[60131] ^ n[60132];
assign t[60133] = t[60132] ^ n[60133];
assign t[60134] = t[60133] ^ n[60134];
assign t[60135] = t[60134] ^ n[60135];
assign t[60136] = t[60135] ^ n[60136];
assign t[60137] = t[60136] ^ n[60137];
assign t[60138] = t[60137] ^ n[60138];
assign t[60139] = t[60138] ^ n[60139];
assign t[60140] = t[60139] ^ n[60140];
assign t[60141] = t[60140] ^ n[60141];
assign t[60142] = t[60141] ^ n[60142];
assign t[60143] = t[60142] ^ n[60143];
assign t[60144] = t[60143] ^ n[60144];
assign t[60145] = t[60144] ^ n[60145];
assign t[60146] = t[60145] ^ n[60146];
assign t[60147] = t[60146] ^ n[60147];
assign t[60148] = t[60147] ^ n[60148];
assign t[60149] = t[60148] ^ n[60149];
assign t[60150] = t[60149] ^ n[60150];
assign t[60151] = t[60150] ^ n[60151];
assign t[60152] = t[60151] ^ n[60152];
assign t[60153] = t[60152] ^ n[60153];
assign t[60154] = t[60153] ^ n[60154];
assign t[60155] = t[60154] ^ n[60155];
assign t[60156] = t[60155] ^ n[60156];
assign t[60157] = t[60156] ^ n[60157];
assign t[60158] = t[60157] ^ n[60158];
assign t[60159] = t[60158] ^ n[60159];
assign t[60160] = t[60159] ^ n[60160];
assign t[60161] = t[60160] ^ n[60161];
assign t[60162] = t[60161] ^ n[60162];
assign t[60163] = t[60162] ^ n[60163];
assign t[60164] = t[60163] ^ n[60164];
assign t[60165] = t[60164] ^ n[60165];
assign t[60166] = t[60165] ^ n[60166];
assign t[60167] = t[60166] ^ n[60167];
assign t[60168] = t[60167] ^ n[60168];
assign t[60169] = t[60168] ^ n[60169];
assign t[60170] = t[60169] ^ n[60170];
assign t[60171] = t[60170] ^ n[60171];
assign t[60172] = t[60171] ^ n[60172];
assign t[60173] = t[60172] ^ n[60173];
assign t[60174] = t[60173] ^ n[60174];
assign t[60175] = t[60174] ^ n[60175];
assign t[60176] = t[60175] ^ n[60176];
assign t[60177] = t[60176] ^ n[60177];
assign t[60178] = t[60177] ^ n[60178];
assign t[60179] = t[60178] ^ n[60179];
assign t[60180] = t[60179] ^ n[60180];
assign t[60181] = t[60180] ^ n[60181];
assign t[60182] = t[60181] ^ n[60182];
assign t[60183] = t[60182] ^ n[60183];
assign t[60184] = t[60183] ^ n[60184];
assign t[60185] = t[60184] ^ n[60185];
assign t[60186] = t[60185] ^ n[60186];
assign t[60187] = t[60186] ^ n[60187];
assign t[60188] = t[60187] ^ n[60188];
assign t[60189] = t[60188] ^ n[60189];
assign t[60190] = t[60189] ^ n[60190];
assign t[60191] = t[60190] ^ n[60191];
assign t[60192] = t[60191] ^ n[60192];
assign t[60193] = t[60192] ^ n[60193];
assign t[60194] = t[60193] ^ n[60194];
assign t[60195] = t[60194] ^ n[60195];
assign t[60196] = t[60195] ^ n[60196];
assign t[60197] = t[60196] ^ n[60197];
assign t[60198] = t[60197] ^ n[60198];
assign t[60199] = t[60198] ^ n[60199];
assign t[60200] = t[60199] ^ n[60200];
assign t[60201] = t[60200] ^ n[60201];
assign t[60202] = t[60201] ^ n[60202];
assign t[60203] = t[60202] ^ n[60203];
assign t[60204] = t[60203] ^ n[60204];
assign t[60205] = t[60204] ^ n[60205];
assign t[60206] = t[60205] ^ n[60206];
assign t[60207] = t[60206] ^ n[60207];
assign t[60208] = t[60207] ^ n[60208];
assign t[60209] = t[60208] ^ n[60209];
assign t[60210] = t[60209] ^ n[60210];
assign t[60211] = t[60210] ^ n[60211];
assign t[60212] = t[60211] ^ n[60212];
assign t[60213] = t[60212] ^ n[60213];
assign t[60214] = t[60213] ^ n[60214];
assign t[60215] = t[60214] ^ n[60215];
assign t[60216] = t[60215] ^ n[60216];
assign t[60217] = t[60216] ^ n[60217];
assign t[60218] = t[60217] ^ n[60218];
assign t[60219] = t[60218] ^ n[60219];
assign t[60220] = t[60219] ^ n[60220];
assign t[60221] = t[60220] ^ n[60221];
assign t[60222] = t[60221] ^ n[60222];
assign t[60223] = t[60222] ^ n[60223];
assign t[60224] = t[60223] ^ n[60224];
assign t[60225] = t[60224] ^ n[60225];
assign t[60226] = t[60225] ^ n[60226];
assign t[60227] = t[60226] ^ n[60227];
assign t[60228] = t[60227] ^ n[60228];
assign t[60229] = t[60228] ^ n[60229];
assign t[60230] = t[60229] ^ n[60230];
assign t[60231] = t[60230] ^ n[60231];
assign t[60232] = t[60231] ^ n[60232];
assign t[60233] = t[60232] ^ n[60233];
assign t[60234] = t[60233] ^ n[60234];
assign t[60235] = t[60234] ^ n[60235];
assign t[60236] = t[60235] ^ n[60236];
assign t[60237] = t[60236] ^ n[60237];
assign t[60238] = t[60237] ^ n[60238];
assign t[60239] = t[60238] ^ n[60239];
assign t[60240] = t[60239] ^ n[60240];
assign t[60241] = t[60240] ^ n[60241];
assign t[60242] = t[60241] ^ n[60242];
assign t[60243] = t[60242] ^ n[60243];
assign t[60244] = t[60243] ^ n[60244];
assign t[60245] = t[60244] ^ n[60245];
assign t[60246] = t[60245] ^ n[60246];
assign t[60247] = t[60246] ^ n[60247];
assign t[60248] = t[60247] ^ n[60248];
assign t[60249] = t[60248] ^ n[60249];
assign t[60250] = t[60249] ^ n[60250];
assign t[60251] = t[60250] ^ n[60251];
assign t[60252] = t[60251] ^ n[60252];
assign t[60253] = t[60252] ^ n[60253];
assign t[60254] = t[60253] ^ n[60254];
assign t[60255] = t[60254] ^ n[60255];
assign t[60256] = t[60255] ^ n[60256];
assign t[60257] = t[60256] ^ n[60257];
assign t[60258] = t[60257] ^ n[60258];
assign t[60259] = t[60258] ^ n[60259];
assign t[60260] = t[60259] ^ n[60260];
assign t[60261] = t[60260] ^ n[60261];
assign t[60262] = t[60261] ^ n[60262];
assign t[60263] = t[60262] ^ n[60263];
assign t[60264] = t[60263] ^ n[60264];
assign t[60265] = t[60264] ^ n[60265];
assign t[60266] = t[60265] ^ n[60266];
assign t[60267] = t[60266] ^ n[60267];
assign t[60268] = t[60267] ^ n[60268];
assign t[60269] = t[60268] ^ n[60269];
assign t[60270] = t[60269] ^ n[60270];
assign t[60271] = t[60270] ^ n[60271];
assign t[60272] = t[60271] ^ n[60272];
assign t[60273] = t[60272] ^ n[60273];
assign t[60274] = t[60273] ^ n[60274];
assign t[60275] = t[60274] ^ n[60275];
assign t[60276] = t[60275] ^ n[60276];
assign t[60277] = t[60276] ^ n[60277];
assign t[60278] = t[60277] ^ n[60278];
assign t[60279] = t[60278] ^ n[60279];
assign t[60280] = t[60279] ^ n[60280];
assign t[60281] = t[60280] ^ n[60281];
assign t[60282] = t[60281] ^ n[60282];
assign t[60283] = t[60282] ^ n[60283];
assign t[60284] = t[60283] ^ n[60284];
assign t[60285] = t[60284] ^ n[60285];
assign t[60286] = t[60285] ^ n[60286];
assign t[60287] = t[60286] ^ n[60287];
assign t[60288] = t[60287] ^ n[60288];
assign t[60289] = t[60288] ^ n[60289];
assign t[60290] = t[60289] ^ n[60290];
assign t[60291] = t[60290] ^ n[60291];
assign t[60292] = t[60291] ^ n[60292];
assign t[60293] = t[60292] ^ n[60293];
assign t[60294] = t[60293] ^ n[60294];
assign t[60295] = t[60294] ^ n[60295];
assign t[60296] = t[60295] ^ n[60296];
assign t[60297] = t[60296] ^ n[60297];
assign t[60298] = t[60297] ^ n[60298];
assign t[60299] = t[60298] ^ n[60299];
assign t[60300] = t[60299] ^ n[60300];
assign t[60301] = t[60300] ^ n[60301];
assign t[60302] = t[60301] ^ n[60302];
assign t[60303] = t[60302] ^ n[60303];
assign t[60304] = t[60303] ^ n[60304];
assign t[60305] = t[60304] ^ n[60305];
assign t[60306] = t[60305] ^ n[60306];
assign t[60307] = t[60306] ^ n[60307];
assign t[60308] = t[60307] ^ n[60308];
assign t[60309] = t[60308] ^ n[60309];
assign t[60310] = t[60309] ^ n[60310];
assign t[60311] = t[60310] ^ n[60311];
assign t[60312] = t[60311] ^ n[60312];
assign t[60313] = t[60312] ^ n[60313];
assign t[60314] = t[60313] ^ n[60314];
assign t[60315] = t[60314] ^ n[60315];
assign t[60316] = t[60315] ^ n[60316];
assign t[60317] = t[60316] ^ n[60317];
assign t[60318] = t[60317] ^ n[60318];
assign t[60319] = t[60318] ^ n[60319];
assign t[60320] = t[60319] ^ n[60320];
assign t[60321] = t[60320] ^ n[60321];
assign t[60322] = t[60321] ^ n[60322];
assign t[60323] = t[60322] ^ n[60323];
assign t[60324] = t[60323] ^ n[60324];
assign t[60325] = t[60324] ^ n[60325];
assign t[60326] = t[60325] ^ n[60326];
assign t[60327] = t[60326] ^ n[60327];
assign t[60328] = t[60327] ^ n[60328];
assign t[60329] = t[60328] ^ n[60329];
assign t[60330] = t[60329] ^ n[60330];
assign t[60331] = t[60330] ^ n[60331];
assign t[60332] = t[60331] ^ n[60332];
assign t[60333] = t[60332] ^ n[60333];
assign t[60334] = t[60333] ^ n[60334];
assign t[60335] = t[60334] ^ n[60335];
assign t[60336] = t[60335] ^ n[60336];
assign t[60337] = t[60336] ^ n[60337];
assign t[60338] = t[60337] ^ n[60338];
assign t[60339] = t[60338] ^ n[60339];
assign t[60340] = t[60339] ^ n[60340];
assign t[60341] = t[60340] ^ n[60341];
assign t[60342] = t[60341] ^ n[60342];
assign t[60343] = t[60342] ^ n[60343];
assign t[60344] = t[60343] ^ n[60344];
assign t[60345] = t[60344] ^ n[60345];
assign t[60346] = t[60345] ^ n[60346];
assign t[60347] = t[60346] ^ n[60347];
assign t[60348] = t[60347] ^ n[60348];
assign t[60349] = t[60348] ^ n[60349];
assign t[60350] = t[60349] ^ n[60350];
assign t[60351] = t[60350] ^ n[60351];
assign t[60352] = t[60351] ^ n[60352];
assign t[60353] = t[60352] ^ n[60353];
assign t[60354] = t[60353] ^ n[60354];
assign t[60355] = t[60354] ^ n[60355];
assign t[60356] = t[60355] ^ n[60356];
assign t[60357] = t[60356] ^ n[60357];
assign t[60358] = t[60357] ^ n[60358];
assign t[60359] = t[60358] ^ n[60359];
assign t[60360] = t[60359] ^ n[60360];
assign t[60361] = t[60360] ^ n[60361];
assign t[60362] = t[60361] ^ n[60362];
assign t[60363] = t[60362] ^ n[60363];
assign t[60364] = t[60363] ^ n[60364];
assign t[60365] = t[60364] ^ n[60365];
assign t[60366] = t[60365] ^ n[60366];
assign t[60367] = t[60366] ^ n[60367];
assign t[60368] = t[60367] ^ n[60368];
assign t[60369] = t[60368] ^ n[60369];
assign t[60370] = t[60369] ^ n[60370];
assign t[60371] = t[60370] ^ n[60371];
assign t[60372] = t[60371] ^ n[60372];
assign t[60373] = t[60372] ^ n[60373];
assign t[60374] = t[60373] ^ n[60374];
assign t[60375] = t[60374] ^ n[60375];
assign t[60376] = t[60375] ^ n[60376];
assign t[60377] = t[60376] ^ n[60377];
assign t[60378] = t[60377] ^ n[60378];
assign t[60379] = t[60378] ^ n[60379];
assign t[60380] = t[60379] ^ n[60380];
assign t[60381] = t[60380] ^ n[60381];
assign t[60382] = t[60381] ^ n[60382];
assign t[60383] = t[60382] ^ n[60383];
assign t[60384] = t[60383] ^ n[60384];
assign t[60385] = t[60384] ^ n[60385];
assign t[60386] = t[60385] ^ n[60386];
assign t[60387] = t[60386] ^ n[60387];
assign t[60388] = t[60387] ^ n[60388];
assign t[60389] = t[60388] ^ n[60389];
assign t[60390] = t[60389] ^ n[60390];
assign t[60391] = t[60390] ^ n[60391];
assign t[60392] = t[60391] ^ n[60392];
assign t[60393] = t[60392] ^ n[60393];
assign t[60394] = t[60393] ^ n[60394];
assign t[60395] = t[60394] ^ n[60395];
assign t[60396] = t[60395] ^ n[60396];
assign t[60397] = t[60396] ^ n[60397];
assign t[60398] = t[60397] ^ n[60398];
assign t[60399] = t[60398] ^ n[60399];
assign t[60400] = t[60399] ^ n[60400];
assign t[60401] = t[60400] ^ n[60401];
assign t[60402] = t[60401] ^ n[60402];
assign t[60403] = t[60402] ^ n[60403];
assign t[60404] = t[60403] ^ n[60404];
assign t[60405] = t[60404] ^ n[60405];
assign t[60406] = t[60405] ^ n[60406];
assign t[60407] = t[60406] ^ n[60407];
assign t[60408] = t[60407] ^ n[60408];
assign t[60409] = t[60408] ^ n[60409];
assign t[60410] = t[60409] ^ n[60410];
assign t[60411] = t[60410] ^ n[60411];
assign t[60412] = t[60411] ^ n[60412];
assign t[60413] = t[60412] ^ n[60413];
assign t[60414] = t[60413] ^ n[60414];
assign t[60415] = t[60414] ^ n[60415];
assign t[60416] = t[60415] ^ n[60416];
assign t[60417] = t[60416] ^ n[60417];
assign t[60418] = t[60417] ^ n[60418];
assign t[60419] = t[60418] ^ n[60419];
assign t[60420] = t[60419] ^ n[60420];
assign t[60421] = t[60420] ^ n[60421];
assign t[60422] = t[60421] ^ n[60422];
assign t[60423] = t[60422] ^ n[60423];
assign t[60424] = t[60423] ^ n[60424];
assign t[60425] = t[60424] ^ n[60425];
assign t[60426] = t[60425] ^ n[60426];
assign t[60427] = t[60426] ^ n[60427];
assign t[60428] = t[60427] ^ n[60428];
assign t[60429] = t[60428] ^ n[60429];
assign t[60430] = t[60429] ^ n[60430];
assign t[60431] = t[60430] ^ n[60431];
assign t[60432] = t[60431] ^ n[60432];
assign t[60433] = t[60432] ^ n[60433];
assign t[60434] = t[60433] ^ n[60434];
assign t[60435] = t[60434] ^ n[60435];
assign t[60436] = t[60435] ^ n[60436];
assign t[60437] = t[60436] ^ n[60437];
assign t[60438] = t[60437] ^ n[60438];
assign t[60439] = t[60438] ^ n[60439];
assign t[60440] = t[60439] ^ n[60440];
assign t[60441] = t[60440] ^ n[60441];
assign t[60442] = t[60441] ^ n[60442];
assign t[60443] = t[60442] ^ n[60443];
assign t[60444] = t[60443] ^ n[60444];
assign t[60445] = t[60444] ^ n[60445];
assign t[60446] = t[60445] ^ n[60446];
assign t[60447] = t[60446] ^ n[60447];
assign t[60448] = t[60447] ^ n[60448];
assign t[60449] = t[60448] ^ n[60449];
assign t[60450] = t[60449] ^ n[60450];
assign t[60451] = t[60450] ^ n[60451];
assign t[60452] = t[60451] ^ n[60452];
assign t[60453] = t[60452] ^ n[60453];
assign t[60454] = t[60453] ^ n[60454];
assign t[60455] = t[60454] ^ n[60455];
assign t[60456] = t[60455] ^ n[60456];
assign t[60457] = t[60456] ^ n[60457];
assign t[60458] = t[60457] ^ n[60458];
assign t[60459] = t[60458] ^ n[60459];
assign t[60460] = t[60459] ^ n[60460];
assign t[60461] = t[60460] ^ n[60461];
assign t[60462] = t[60461] ^ n[60462];
assign t[60463] = t[60462] ^ n[60463];
assign t[60464] = t[60463] ^ n[60464];
assign t[60465] = t[60464] ^ n[60465];
assign t[60466] = t[60465] ^ n[60466];
assign t[60467] = t[60466] ^ n[60467];
assign t[60468] = t[60467] ^ n[60468];
assign t[60469] = t[60468] ^ n[60469];
assign t[60470] = t[60469] ^ n[60470];
assign t[60471] = t[60470] ^ n[60471];
assign t[60472] = t[60471] ^ n[60472];
assign t[60473] = t[60472] ^ n[60473];
assign t[60474] = t[60473] ^ n[60474];
assign t[60475] = t[60474] ^ n[60475];
assign t[60476] = t[60475] ^ n[60476];
assign t[60477] = t[60476] ^ n[60477];
assign t[60478] = t[60477] ^ n[60478];
assign t[60479] = t[60478] ^ n[60479];
assign t[60480] = t[60479] ^ n[60480];
assign t[60481] = t[60480] ^ n[60481];
assign t[60482] = t[60481] ^ n[60482];
assign t[60483] = t[60482] ^ n[60483];
assign t[60484] = t[60483] ^ n[60484];
assign t[60485] = t[60484] ^ n[60485];
assign t[60486] = t[60485] ^ n[60486];
assign t[60487] = t[60486] ^ n[60487];
assign t[60488] = t[60487] ^ n[60488];
assign t[60489] = t[60488] ^ n[60489];
assign t[60490] = t[60489] ^ n[60490];
assign t[60491] = t[60490] ^ n[60491];
assign t[60492] = t[60491] ^ n[60492];
assign t[60493] = t[60492] ^ n[60493];
assign t[60494] = t[60493] ^ n[60494];
assign t[60495] = t[60494] ^ n[60495];
assign t[60496] = t[60495] ^ n[60496];
assign t[60497] = t[60496] ^ n[60497];
assign t[60498] = t[60497] ^ n[60498];
assign t[60499] = t[60498] ^ n[60499];
assign t[60500] = t[60499] ^ n[60500];
assign t[60501] = t[60500] ^ n[60501];
assign t[60502] = t[60501] ^ n[60502];
assign t[60503] = t[60502] ^ n[60503];
assign t[60504] = t[60503] ^ n[60504];
assign t[60505] = t[60504] ^ n[60505];
assign t[60506] = t[60505] ^ n[60506];
assign t[60507] = t[60506] ^ n[60507];
assign t[60508] = t[60507] ^ n[60508];
assign t[60509] = t[60508] ^ n[60509];
assign t[60510] = t[60509] ^ n[60510];
assign t[60511] = t[60510] ^ n[60511];
assign t[60512] = t[60511] ^ n[60512];
assign t[60513] = t[60512] ^ n[60513];
assign t[60514] = t[60513] ^ n[60514];
assign t[60515] = t[60514] ^ n[60515];
assign t[60516] = t[60515] ^ n[60516];
assign t[60517] = t[60516] ^ n[60517];
assign t[60518] = t[60517] ^ n[60518];
assign t[60519] = t[60518] ^ n[60519];
assign t[60520] = t[60519] ^ n[60520];
assign t[60521] = t[60520] ^ n[60521];
assign t[60522] = t[60521] ^ n[60522];
assign t[60523] = t[60522] ^ n[60523];
assign t[60524] = t[60523] ^ n[60524];
assign t[60525] = t[60524] ^ n[60525];
assign t[60526] = t[60525] ^ n[60526];
assign t[60527] = t[60526] ^ n[60527];
assign t[60528] = t[60527] ^ n[60528];
assign t[60529] = t[60528] ^ n[60529];
assign t[60530] = t[60529] ^ n[60530];
assign t[60531] = t[60530] ^ n[60531];
assign t[60532] = t[60531] ^ n[60532];
assign t[60533] = t[60532] ^ n[60533];
assign t[60534] = t[60533] ^ n[60534];
assign t[60535] = t[60534] ^ n[60535];
assign t[60536] = t[60535] ^ n[60536];
assign t[60537] = t[60536] ^ n[60537];
assign t[60538] = t[60537] ^ n[60538];
assign t[60539] = t[60538] ^ n[60539];
assign t[60540] = t[60539] ^ n[60540];
assign t[60541] = t[60540] ^ n[60541];
assign t[60542] = t[60541] ^ n[60542];
assign t[60543] = t[60542] ^ n[60543];
assign t[60544] = t[60543] ^ n[60544];
assign t[60545] = t[60544] ^ n[60545];
assign t[60546] = t[60545] ^ n[60546];
assign t[60547] = t[60546] ^ n[60547];
assign t[60548] = t[60547] ^ n[60548];
assign t[60549] = t[60548] ^ n[60549];
assign t[60550] = t[60549] ^ n[60550];
assign t[60551] = t[60550] ^ n[60551];
assign t[60552] = t[60551] ^ n[60552];
assign t[60553] = t[60552] ^ n[60553];
assign t[60554] = t[60553] ^ n[60554];
assign t[60555] = t[60554] ^ n[60555];
assign t[60556] = t[60555] ^ n[60556];
assign t[60557] = t[60556] ^ n[60557];
assign t[60558] = t[60557] ^ n[60558];
assign t[60559] = t[60558] ^ n[60559];
assign t[60560] = t[60559] ^ n[60560];
assign t[60561] = t[60560] ^ n[60561];
assign t[60562] = t[60561] ^ n[60562];
assign t[60563] = t[60562] ^ n[60563];
assign t[60564] = t[60563] ^ n[60564];
assign t[60565] = t[60564] ^ n[60565];
assign t[60566] = t[60565] ^ n[60566];
assign t[60567] = t[60566] ^ n[60567];
assign t[60568] = t[60567] ^ n[60568];
assign t[60569] = t[60568] ^ n[60569];
assign t[60570] = t[60569] ^ n[60570];
assign t[60571] = t[60570] ^ n[60571];
assign t[60572] = t[60571] ^ n[60572];
assign t[60573] = t[60572] ^ n[60573];
assign t[60574] = t[60573] ^ n[60574];
assign t[60575] = t[60574] ^ n[60575];
assign t[60576] = t[60575] ^ n[60576];
assign t[60577] = t[60576] ^ n[60577];
assign t[60578] = t[60577] ^ n[60578];
assign t[60579] = t[60578] ^ n[60579];
assign t[60580] = t[60579] ^ n[60580];
assign t[60581] = t[60580] ^ n[60581];
assign t[60582] = t[60581] ^ n[60582];
assign t[60583] = t[60582] ^ n[60583];
assign t[60584] = t[60583] ^ n[60584];
assign t[60585] = t[60584] ^ n[60585];
assign t[60586] = t[60585] ^ n[60586];
assign t[60587] = t[60586] ^ n[60587];
assign t[60588] = t[60587] ^ n[60588];
assign t[60589] = t[60588] ^ n[60589];
assign t[60590] = t[60589] ^ n[60590];
assign t[60591] = t[60590] ^ n[60591];
assign t[60592] = t[60591] ^ n[60592];
assign t[60593] = t[60592] ^ n[60593];
assign t[60594] = t[60593] ^ n[60594];
assign t[60595] = t[60594] ^ n[60595];
assign t[60596] = t[60595] ^ n[60596];
assign t[60597] = t[60596] ^ n[60597];
assign t[60598] = t[60597] ^ n[60598];
assign t[60599] = t[60598] ^ n[60599];
assign t[60600] = t[60599] ^ n[60600];
assign t[60601] = t[60600] ^ n[60601];
assign t[60602] = t[60601] ^ n[60602];
assign t[60603] = t[60602] ^ n[60603];
assign t[60604] = t[60603] ^ n[60604];
assign t[60605] = t[60604] ^ n[60605];
assign t[60606] = t[60605] ^ n[60606];
assign t[60607] = t[60606] ^ n[60607];
assign t[60608] = t[60607] ^ n[60608];
assign t[60609] = t[60608] ^ n[60609];
assign t[60610] = t[60609] ^ n[60610];
assign t[60611] = t[60610] ^ n[60611];
assign t[60612] = t[60611] ^ n[60612];
assign t[60613] = t[60612] ^ n[60613];
assign t[60614] = t[60613] ^ n[60614];
assign t[60615] = t[60614] ^ n[60615];
assign t[60616] = t[60615] ^ n[60616];
assign t[60617] = t[60616] ^ n[60617];
assign t[60618] = t[60617] ^ n[60618];
assign t[60619] = t[60618] ^ n[60619];
assign t[60620] = t[60619] ^ n[60620];
assign t[60621] = t[60620] ^ n[60621];
assign t[60622] = t[60621] ^ n[60622];
assign t[60623] = t[60622] ^ n[60623];
assign t[60624] = t[60623] ^ n[60624];
assign t[60625] = t[60624] ^ n[60625];
assign t[60626] = t[60625] ^ n[60626];
assign t[60627] = t[60626] ^ n[60627];
assign t[60628] = t[60627] ^ n[60628];
assign t[60629] = t[60628] ^ n[60629];
assign t[60630] = t[60629] ^ n[60630];
assign t[60631] = t[60630] ^ n[60631];
assign t[60632] = t[60631] ^ n[60632];
assign t[60633] = t[60632] ^ n[60633];
assign t[60634] = t[60633] ^ n[60634];
assign t[60635] = t[60634] ^ n[60635];
assign t[60636] = t[60635] ^ n[60636];
assign t[60637] = t[60636] ^ n[60637];
assign t[60638] = t[60637] ^ n[60638];
assign t[60639] = t[60638] ^ n[60639];
assign t[60640] = t[60639] ^ n[60640];
assign t[60641] = t[60640] ^ n[60641];
assign t[60642] = t[60641] ^ n[60642];
assign t[60643] = t[60642] ^ n[60643];
assign t[60644] = t[60643] ^ n[60644];
assign t[60645] = t[60644] ^ n[60645];
assign t[60646] = t[60645] ^ n[60646];
assign t[60647] = t[60646] ^ n[60647];
assign t[60648] = t[60647] ^ n[60648];
assign t[60649] = t[60648] ^ n[60649];
assign t[60650] = t[60649] ^ n[60650];
assign t[60651] = t[60650] ^ n[60651];
assign t[60652] = t[60651] ^ n[60652];
assign t[60653] = t[60652] ^ n[60653];
assign t[60654] = t[60653] ^ n[60654];
assign t[60655] = t[60654] ^ n[60655];
assign t[60656] = t[60655] ^ n[60656];
assign t[60657] = t[60656] ^ n[60657];
assign t[60658] = t[60657] ^ n[60658];
assign t[60659] = t[60658] ^ n[60659];
assign t[60660] = t[60659] ^ n[60660];
assign t[60661] = t[60660] ^ n[60661];
assign t[60662] = t[60661] ^ n[60662];
assign t[60663] = t[60662] ^ n[60663];
assign t[60664] = t[60663] ^ n[60664];
assign t[60665] = t[60664] ^ n[60665];
assign t[60666] = t[60665] ^ n[60666];
assign t[60667] = t[60666] ^ n[60667];
assign t[60668] = t[60667] ^ n[60668];
assign t[60669] = t[60668] ^ n[60669];
assign t[60670] = t[60669] ^ n[60670];
assign t[60671] = t[60670] ^ n[60671];
assign t[60672] = t[60671] ^ n[60672];
assign t[60673] = t[60672] ^ n[60673];
assign t[60674] = t[60673] ^ n[60674];
assign t[60675] = t[60674] ^ n[60675];
assign t[60676] = t[60675] ^ n[60676];
assign t[60677] = t[60676] ^ n[60677];
assign t[60678] = t[60677] ^ n[60678];
assign t[60679] = t[60678] ^ n[60679];
assign t[60680] = t[60679] ^ n[60680];
assign t[60681] = t[60680] ^ n[60681];
assign t[60682] = t[60681] ^ n[60682];
assign t[60683] = t[60682] ^ n[60683];
assign t[60684] = t[60683] ^ n[60684];
assign t[60685] = t[60684] ^ n[60685];
assign t[60686] = t[60685] ^ n[60686];
assign t[60687] = t[60686] ^ n[60687];
assign t[60688] = t[60687] ^ n[60688];
assign t[60689] = t[60688] ^ n[60689];
assign t[60690] = t[60689] ^ n[60690];
assign t[60691] = t[60690] ^ n[60691];
assign t[60692] = t[60691] ^ n[60692];
assign t[60693] = t[60692] ^ n[60693];
assign t[60694] = t[60693] ^ n[60694];
assign t[60695] = t[60694] ^ n[60695];
assign t[60696] = t[60695] ^ n[60696];
assign t[60697] = t[60696] ^ n[60697];
assign t[60698] = t[60697] ^ n[60698];
assign t[60699] = t[60698] ^ n[60699];
assign t[60700] = t[60699] ^ n[60700];
assign t[60701] = t[60700] ^ n[60701];
assign t[60702] = t[60701] ^ n[60702];
assign t[60703] = t[60702] ^ n[60703];
assign t[60704] = t[60703] ^ n[60704];
assign t[60705] = t[60704] ^ n[60705];
assign t[60706] = t[60705] ^ n[60706];
assign t[60707] = t[60706] ^ n[60707];
assign t[60708] = t[60707] ^ n[60708];
assign t[60709] = t[60708] ^ n[60709];
assign t[60710] = t[60709] ^ n[60710];
assign t[60711] = t[60710] ^ n[60711];
assign t[60712] = t[60711] ^ n[60712];
assign t[60713] = t[60712] ^ n[60713];
assign t[60714] = t[60713] ^ n[60714];
assign t[60715] = t[60714] ^ n[60715];
assign t[60716] = t[60715] ^ n[60716];
assign t[60717] = t[60716] ^ n[60717];
assign t[60718] = t[60717] ^ n[60718];
assign t[60719] = t[60718] ^ n[60719];
assign t[60720] = t[60719] ^ n[60720];
assign t[60721] = t[60720] ^ n[60721];
assign t[60722] = t[60721] ^ n[60722];
assign t[60723] = t[60722] ^ n[60723];
assign t[60724] = t[60723] ^ n[60724];
assign t[60725] = t[60724] ^ n[60725];
assign t[60726] = t[60725] ^ n[60726];
assign t[60727] = t[60726] ^ n[60727];
assign t[60728] = t[60727] ^ n[60728];
assign t[60729] = t[60728] ^ n[60729];
assign t[60730] = t[60729] ^ n[60730];
assign t[60731] = t[60730] ^ n[60731];
assign t[60732] = t[60731] ^ n[60732];
assign t[60733] = t[60732] ^ n[60733];
assign t[60734] = t[60733] ^ n[60734];
assign t[60735] = t[60734] ^ n[60735];
assign t[60736] = t[60735] ^ n[60736];
assign t[60737] = t[60736] ^ n[60737];
assign t[60738] = t[60737] ^ n[60738];
assign t[60739] = t[60738] ^ n[60739];
assign t[60740] = t[60739] ^ n[60740];
assign t[60741] = t[60740] ^ n[60741];
assign t[60742] = t[60741] ^ n[60742];
assign t[60743] = t[60742] ^ n[60743];
assign t[60744] = t[60743] ^ n[60744];
assign t[60745] = t[60744] ^ n[60745];
assign t[60746] = t[60745] ^ n[60746];
assign t[60747] = t[60746] ^ n[60747];
assign t[60748] = t[60747] ^ n[60748];
assign t[60749] = t[60748] ^ n[60749];
assign t[60750] = t[60749] ^ n[60750];
assign t[60751] = t[60750] ^ n[60751];
assign t[60752] = t[60751] ^ n[60752];
assign t[60753] = t[60752] ^ n[60753];
assign t[60754] = t[60753] ^ n[60754];
assign t[60755] = t[60754] ^ n[60755];
assign t[60756] = t[60755] ^ n[60756];
assign t[60757] = t[60756] ^ n[60757];
assign t[60758] = t[60757] ^ n[60758];
assign t[60759] = t[60758] ^ n[60759];
assign t[60760] = t[60759] ^ n[60760];
assign t[60761] = t[60760] ^ n[60761];
assign t[60762] = t[60761] ^ n[60762];
assign t[60763] = t[60762] ^ n[60763];
assign t[60764] = t[60763] ^ n[60764];
assign t[60765] = t[60764] ^ n[60765];
assign t[60766] = t[60765] ^ n[60766];
assign t[60767] = t[60766] ^ n[60767];
assign t[60768] = t[60767] ^ n[60768];
assign t[60769] = t[60768] ^ n[60769];
assign t[60770] = t[60769] ^ n[60770];
assign t[60771] = t[60770] ^ n[60771];
assign t[60772] = t[60771] ^ n[60772];
assign t[60773] = t[60772] ^ n[60773];
assign t[60774] = t[60773] ^ n[60774];
assign t[60775] = t[60774] ^ n[60775];
assign t[60776] = t[60775] ^ n[60776];
assign t[60777] = t[60776] ^ n[60777];
assign t[60778] = t[60777] ^ n[60778];
assign t[60779] = t[60778] ^ n[60779];
assign t[60780] = t[60779] ^ n[60780];
assign t[60781] = t[60780] ^ n[60781];
assign t[60782] = t[60781] ^ n[60782];
assign t[60783] = t[60782] ^ n[60783];
assign t[60784] = t[60783] ^ n[60784];
assign t[60785] = t[60784] ^ n[60785];
assign t[60786] = t[60785] ^ n[60786];
assign t[60787] = t[60786] ^ n[60787];
assign t[60788] = t[60787] ^ n[60788];
assign t[60789] = t[60788] ^ n[60789];
assign t[60790] = t[60789] ^ n[60790];
assign t[60791] = t[60790] ^ n[60791];
assign t[60792] = t[60791] ^ n[60792];
assign t[60793] = t[60792] ^ n[60793];
assign t[60794] = t[60793] ^ n[60794];
assign t[60795] = t[60794] ^ n[60795];
assign t[60796] = t[60795] ^ n[60796];
assign t[60797] = t[60796] ^ n[60797];
assign t[60798] = t[60797] ^ n[60798];
assign t[60799] = t[60798] ^ n[60799];
assign t[60800] = t[60799] ^ n[60800];
assign t[60801] = t[60800] ^ n[60801];
assign t[60802] = t[60801] ^ n[60802];
assign t[60803] = t[60802] ^ n[60803];
assign t[60804] = t[60803] ^ n[60804];
assign t[60805] = t[60804] ^ n[60805];
assign t[60806] = t[60805] ^ n[60806];
assign t[60807] = t[60806] ^ n[60807];
assign t[60808] = t[60807] ^ n[60808];
assign t[60809] = t[60808] ^ n[60809];
assign t[60810] = t[60809] ^ n[60810];
assign t[60811] = t[60810] ^ n[60811];
assign t[60812] = t[60811] ^ n[60812];
assign t[60813] = t[60812] ^ n[60813];
assign t[60814] = t[60813] ^ n[60814];
assign t[60815] = t[60814] ^ n[60815];
assign t[60816] = t[60815] ^ n[60816];
assign t[60817] = t[60816] ^ n[60817];
assign t[60818] = t[60817] ^ n[60818];
assign t[60819] = t[60818] ^ n[60819];
assign t[60820] = t[60819] ^ n[60820];
assign t[60821] = t[60820] ^ n[60821];
assign t[60822] = t[60821] ^ n[60822];
assign t[60823] = t[60822] ^ n[60823];
assign t[60824] = t[60823] ^ n[60824];
assign t[60825] = t[60824] ^ n[60825];
assign t[60826] = t[60825] ^ n[60826];
assign t[60827] = t[60826] ^ n[60827];
assign t[60828] = t[60827] ^ n[60828];
assign t[60829] = t[60828] ^ n[60829];
assign t[60830] = t[60829] ^ n[60830];
assign t[60831] = t[60830] ^ n[60831];
assign t[60832] = t[60831] ^ n[60832];
assign t[60833] = t[60832] ^ n[60833];
assign t[60834] = t[60833] ^ n[60834];
assign t[60835] = t[60834] ^ n[60835];
assign t[60836] = t[60835] ^ n[60836];
assign t[60837] = t[60836] ^ n[60837];
assign t[60838] = t[60837] ^ n[60838];
assign t[60839] = t[60838] ^ n[60839];
assign t[60840] = t[60839] ^ n[60840];
assign t[60841] = t[60840] ^ n[60841];
assign t[60842] = t[60841] ^ n[60842];
assign t[60843] = t[60842] ^ n[60843];
assign t[60844] = t[60843] ^ n[60844];
assign t[60845] = t[60844] ^ n[60845];
assign t[60846] = t[60845] ^ n[60846];
assign t[60847] = t[60846] ^ n[60847];
assign t[60848] = t[60847] ^ n[60848];
assign t[60849] = t[60848] ^ n[60849];
assign t[60850] = t[60849] ^ n[60850];
assign t[60851] = t[60850] ^ n[60851];
assign t[60852] = t[60851] ^ n[60852];
assign t[60853] = t[60852] ^ n[60853];
assign t[60854] = t[60853] ^ n[60854];
assign t[60855] = t[60854] ^ n[60855];
assign t[60856] = t[60855] ^ n[60856];
assign t[60857] = t[60856] ^ n[60857];
assign t[60858] = t[60857] ^ n[60858];
assign t[60859] = t[60858] ^ n[60859];
assign t[60860] = t[60859] ^ n[60860];
assign t[60861] = t[60860] ^ n[60861];
assign t[60862] = t[60861] ^ n[60862];
assign t[60863] = t[60862] ^ n[60863];
assign t[60864] = t[60863] ^ n[60864];
assign t[60865] = t[60864] ^ n[60865];
assign t[60866] = t[60865] ^ n[60866];
assign t[60867] = t[60866] ^ n[60867];
assign t[60868] = t[60867] ^ n[60868];
assign t[60869] = t[60868] ^ n[60869];
assign t[60870] = t[60869] ^ n[60870];
assign t[60871] = t[60870] ^ n[60871];
assign t[60872] = t[60871] ^ n[60872];
assign t[60873] = t[60872] ^ n[60873];
assign t[60874] = t[60873] ^ n[60874];
assign t[60875] = t[60874] ^ n[60875];
assign t[60876] = t[60875] ^ n[60876];
assign t[60877] = t[60876] ^ n[60877];
assign t[60878] = t[60877] ^ n[60878];
assign t[60879] = t[60878] ^ n[60879];
assign t[60880] = t[60879] ^ n[60880];
assign t[60881] = t[60880] ^ n[60881];
assign t[60882] = t[60881] ^ n[60882];
assign t[60883] = t[60882] ^ n[60883];
assign t[60884] = t[60883] ^ n[60884];
assign t[60885] = t[60884] ^ n[60885];
assign t[60886] = t[60885] ^ n[60886];
assign t[60887] = t[60886] ^ n[60887];
assign t[60888] = t[60887] ^ n[60888];
assign t[60889] = t[60888] ^ n[60889];
assign t[60890] = t[60889] ^ n[60890];
assign t[60891] = t[60890] ^ n[60891];
assign t[60892] = t[60891] ^ n[60892];
assign t[60893] = t[60892] ^ n[60893];
assign t[60894] = t[60893] ^ n[60894];
assign t[60895] = t[60894] ^ n[60895];
assign t[60896] = t[60895] ^ n[60896];
assign t[60897] = t[60896] ^ n[60897];
assign t[60898] = t[60897] ^ n[60898];
assign t[60899] = t[60898] ^ n[60899];
assign t[60900] = t[60899] ^ n[60900];
assign t[60901] = t[60900] ^ n[60901];
assign t[60902] = t[60901] ^ n[60902];
assign t[60903] = t[60902] ^ n[60903];
assign t[60904] = t[60903] ^ n[60904];
assign t[60905] = t[60904] ^ n[60905];
assign t[60906] = t[60905] ^ n[60906];
assign t[60907] = t[60906] ^ n[60907];
assign t[60908] = t[60907] ^ n[60908];
assign t[60909] = t[60908] ^ n[60909];
assign t[60910] = t[60909] ^ n[60910];
assign t[60911] = t[60910] ^ n[60911];
assign t[60912] = t[60911] ^ n[60912];
assign t[60913] = t[60912] ^ n[60913];
assign t[60914] = t[60913] ^ n[60914];
assign t[60915] = t[60914] ^ n[60915];
assign t[60916] = t[60915] ^ n[60916];
assign t[60917] = t[60916] ^ n[60917];
assign t[60918] = t[60917] ^ n[60918];
assign t[60919] = t[60918] ^ n[60919];
assign t[60920] = t[60919] ^ n[60920];
assign t[60921] = t[60920] ^ n[60921];
assign t[60922] = t[60921] ^ n[60922];
assign t[60923] = t[60922] ^ n[60923];
assign t[60924] = t[60923] ^ n[60924];
assign t[60925] = t[60924] ^ n[60925];
assign t[60926] = t[60925] ^ n[60926];
assign t[60927] = t[60926] ^ n[60927];
assign t[60928] = t[60927] ^ n[60928];
assign t[60929] = t[60928] ^ n[60929];
assign t[60930] = t[60929] ^ n[60930];
assign t[60931] = t[60930] ^ n[60931];
assign t[60932] = t[60931] ^ n[60932];
assign t[60933] = t[60932] ^ n[60933];
assign t[60934] = t[60933] ^ n[60934];
assign t[60935] = t[60934] ^ n[60935];
assign t[60936] = t[60935] ^ n[60936];
assign t[60937] = t[60936] ^ n[60937];
assign t[60938] = t[60937] ^ n[60938];
assign t[60939] = t[60938] ^ n[60939];
assign t[60940] = t[60939] ^ n[60940];
assign t[60941] = t[60940] ^ n[60941];
assign t[60942] = t[60941] ^ n[60942];
assign t[60943] = t[60942] ^ n[60943];
assign t[60944] = t[60943] ^ n[60944];
assign t[60945] = t[60944] ^ n[60945];
assign t[60946] = t[60945] ^ n[60946];
assign t[60947] = t[60946] ^ n[60947];
assign t[60948] = t[60947] ^ n[60948];
assign t[60949] = t[60948] ^ n[60949];
assign t[60950] = t[60949] ^ n[60950];
assign t[60951] = t[60950] ^ n[60951];
assign t[60952] = t[60951] ^ n[60952];
assign t[60953] = t[60952] ^ n[60953];
assign t[60954] = t[60953] ^ n[60954];
assign t[60955] = t[60954] ^ n[60955];
assign t[60956] = t[60955] ^ n[60956];
assign t[60957] = t[60956] ^ n[60957];
assign t[60958] = t[60957] ^ n[60958];
assign t[60959] = t[60958] ^ n[60959];
assign t[60960] = t[60959] ^ n[60960];
assign t[60961] = t[60960] ^ n[60961];
assign t[60962] = t[60961] ^ n[60962];
assign t[60963] = t[60962] ^ n[60963];
assign t[60964] = t[60963] ^ n[60964];
assign t[60965] = t[60964] ^ n[60965];
assign t[60966] = t[60965] ^ n[60966];
assign t[60967] = t[60966] ^ n[60967];
assign t[60968] = t[60967] ^ n[60968];
assign t[60969] = t[60968] ^ n[60969];
assign t[60970] = t[60969] ^ n[60970];
assign t[60971] = t[60970] ^ n[60971];
assign t[60972] = t[60971] ^ n[60972];
assign t[60973] = t[60972] ^ n[60973];
assign t[60974] = t[60973] ^ n[60974];
assign t[60975] = t[60974] ^ n[60975];
assign t[60976] = t[60975] ^ n[60976];
assign t[60977] = t[60976] ^ n[60977];
assign t[60978] = t[60977] ^ n[60978];
assign t[60979] = t[60978] ^ n[60979];
assign t[60980] = t[60979] ^ n[60980];
assign t[60981] = t[60980] ^ n[60981];
assign t[60982] = t[60981] ^ n[60982];
assign t[60983] = t[60982] ^ n[60983];
assign t[60984] = t[60983] ^ n[60984];
assign t[60985] = t[60984] ^ n[60985];
assign t[60986] = t[60985] ^ n[60986];
assign t[60987] = t[60986] ^ n[60987];
assign t[60988] = t[60987] ^ n[60988];
assign t[60989] = t[60988] ^ n[60989];
assign t[60990] = t[60989] ^ n[60990];
assign t[60991] = t[60990] ^ n[60991];
assign t[60992] = t[60991] ^ n[60992];
assign t[60993] = t[60992] ^ n[60993];
assign t[60994] = t[60993] ^ n[60994];
assign t[60995] = t[60994] ^ n[60995];
assign t[60996] = t[60995] ^ n[60996];
assign t[60997] = t[60996] ^ n[60997];
assign t[60998] = t[60997] ^ n[60998];
assign t[60999] = t[60998] ^ n[60999];
assign t[61000] = t[60999] ^ n[61000];
assign t[61001] = t[61000] ^ n[61001];
assign t[61002] = t[61001] ^ n[61002];
assign t[61003] = t[61002] ^ n[61003];
assign t[61004] = t[61003] ^ n[61004];
assign t[61005] = t[61004] ^ n[61005];
assign t[61006] = t[61005] ^ n[61006];
assign t[61007] = t[61006] ^ n[61007];
assign t[61008] = t[61007] ^ n[61008];
assign t[61009] = t[61008] ^ n[61009];
assign t[61010] = t[61009] ^ n[61010];
assign t[61011] = t[61010] ^ n[61011];
assign t[61012] = t[61011] ^ n[61012];
assign t[61013] = t[61012] ^ n[61013];
assign t[61014] = t[61013] ^ n[61014];
assign t[61015] = t[61014] ^ n[61015];
assign t[61016] = t[61015] ^ n[61016];
assign t[61017] = t[61016] ^ n[61017];
assign t[61018] = t[61017] ^ n[61018];
assign t[61019] = t[61018] ^ n[61019];
assign t[61020] = t[61019] ^ n[61020];
assign t[61021] = t[61020] ^ n[61021];
assign t[61022] = t[61021] ^ n[61022];
assign t[61023] = t[61022] ^ n[61023];
assign t[61024] = t[61023] ^ n[61024];
assign t[61025] = t[61024] ^ n[61025];
assign t[61026] = t[61025] ^ n[61026];
assign t[61027] = t[61026] ^ n[61027];
assign t[61028] = t[61027] ^ n[61028];
assign t[61029] = t[61028] ^ n[61029];
assign t[61030] = t[61029] ^ n[61030];
assign t[61031] = t[61030] ^ n[61031];
assign t[61032] = t[61031] ^ n[61032];
assign t[61033] = t[61032] ^ n[61033];
assign t[61034] = t[61033] ^ n[61034];
assign t[61035] = t[61034] ^ n[61035];
assign t[61036] = t[61035] ^ n[61036];
assign t[61037] = t[61036] ^ n[61037];
assign t[61038] = t[61037] ^ n[61038];
assign t[61039] = t[61038] ^ n[61039];
assign t[61040] = t[61039] ^ n[61040];
assign t[61041] = t[61040] ^ n[61041];
assign t[61042] = t[61041] ^ n[61042];
assign t[61043] = t[61042] ^ n[61043];
assign t[61044] = t[61043] ^ n[61044];
assign t[61045] = t[61044] ^ n[61045];
assign t[61046] = t[61045] ^ n[61046];
assign t[61047] = t[61046] ^ n[61047];
assign t[61048] = t[61047] ^ n[61048];
assign t[61049] = t[61048] ^ n[61049];
assign t[61050] = t[61049] ^ n[61050];
assign t[61051] = t[61050] ^ n[61051];
assign t[61052] = t[61051] ^ n[61052];
assign t[61053] = t[61052] ^ n[61053];
assign t[61054] = t[61053] ^ n[61054];
assign t[61055] = t[61054] ^ n[61055];
assign t[61056] = t[61055] ^ n[61056];
assign t[61057] = t[61056] ^ n[61057];
assign t[61058] = t[61057] ^ n[61058];
assign t[61059] = t[61058] ^ n[61059];
assign t[61060] = t[61059] ^ n[61060];
assign t[61061] = t[61060] ^ n[61061];
assign t[61062] = t[61061] ^ n[61062];
assign t[61063] = t[61062] ^ n[61063];
assign t[61064] = t[61063] ^ n[61064];
assign t[61065] = t[61064] ^ n[61065];
assign t[61066] = t[61065] ^ n[61066];
assign t[61067] = t[61066] ^ n[61067];
assign t[61068] = t[61067] ^ n[61068];
assign t[61069] = t[61068] ^ n[61069];
assign t[61070] = t[61069] ^ n[61070];
assign t[61071] = t[61070] ^ n[61071];
assign t[61072] = t[61071] ^ n[61072];
assign t[61073] = t[61072] ^ n[61073];
assign t[61074] = t[61073] ^ n[61074];
assign t[61075] = t[61074] ^ n[61075];
assign t[61076] = t[61075] ^ n[61076];
assign t[61077] = t[61076] ^ n[61077];
assign t[61078] = t[61077] ^ n[61078];
assign t[61079] = t[61078] ^ n[61079];
assign t[61080] = t[61079] ^ n[61080];
assign t[61081] = t[61080] ^ n[61081];
assign t[61082] = t[61081] ^ n[61082];
assign t[61083] = t[61082] ^ n[61083];
assign t[61084] = t[61083] ^ n[61084];
assign t[61085] = t[61084] ^ n[61085];
assign t[61086] = t[61085] ^ n[61086];
assign t[61087] = t[61086] ^ n[61087];
assign t[61088] = t[61087] ^ n[61088];
assign t[61089] = t[61088] ^ n[61089];
assign t[61090] = t[61089] ^ n[61090];
assign t[61091] = t[61090] ^ n[61091];
assign t[61092] = t[61091] ^ n[61092];
assign t[61093] = t[61092] ^ n[61093];
assign t[61094] = t[61093] ^ n[61094];
assign t[61095] = t[61094] ^ n[61095];
assign t[61096] = t[61095] ^ n[61096];
assign t[61097] = t[61096] ^ n[61097];
assign t[61098] = t[61097] ^ n[61098];
assign t[61099] = t[61098] ^ n[61099];
assign t[61100] = t[61099] ^ n[61100];
assign t[61101] = t[61100] ^ n[61101];
assign t[61102] = t[61101] ^ n[61102];
assign t[61103] = t[61102] ^ n[61103];
assign t[61104] = t[61103] ^ n[61104];
assign t[61105] = t[61104] ^ n[61105];
assign t[61106] = t[61105] ^ n[61106];
assign t[61107] = t[61106] ^ n[61107];
assign t[61108] = t[61107] ^ n[61108];
assign t[61109] = t[61108] ^ n[61109];
assign t[61110] = t[61109] ^ n[61110];
assign t[61111] = t[61110] ^ n[61111];
assign t[61112] = t[61111] ^ n[61112];
assign t[61113] = t[61112] ^ n[61113];
assign t[61114] = t[61113] ^ n[61114];
assign t[61115] = t[61114] ^ n[61115];
assign t[61116] = t[61115] ^ n[61116];
assign t[61117] = t[61116] ^ n[61117];
assign t[61118] = t[61117] ^ n[61118];
assign t[61119] = t[61118] ^ n[61119];
assign t[61120] = t[61119] ^ n[61120];
assign t[61121] = t[61120] ^ n[61121];
assign t[61122] = t[61121] ^ n[61122];
assign t[61123] = t[61122] ^ n[61123];
assign t[61124] = t[61123] ^ n[61124];
assign t[61125] = t[61124] ^ n[61125];
assign t[61126] = t[61125] ^ n[61126];
assign t[61127] = t[61126] ^ n[61127];
assign t[61128] = t[61127] ^ n[61128];
assign t[61129] = t[61128] ^ n[61129];
assign t[61130] = t[61129] ^ n[61130];
assign t[61131] = t[61130] ^ n[61131];
assign t[61132] = t[61131] ^ n[61132];
assign t[61133] = t[61132] ^ n[61133];
assign t[61134] = t[61133] ^ n[61134];
assign t[61135] = t[61134] ^ n[61135];
assign t[61136] = t[61135] ^ n[61136];
assign t[61137] = t[61136] ^ n[61137];
assign t[61138] = t[61137] ^ n[61138];
assign t[61139] = t[61138] ^ n[61139];
assign t[61140] = t[61139] ^ n[61140];
assign t[61141] = t[61140] ^ n[61141];
assign t[61142] = t[61141] ^ n[61142];
assign t[61143] = t[61142] ^ n[61143];
assign t[61144] = t[61143] ^ n[61144];
assign t[61145] = t[61144] ^ n[61145];
assign t[61146] = t[61145] ^ n[61146];
assign t[61147] = t[61146] ^ n[61147];
assign t[61148] = t[61147] ^ n[61148];
assign t[61149] = t[61148] ^ n[61149];
assign t[61150] = t[61149] ^ n[61150];
assign t[61151] = t[61150] ^ n[61151];
assign t[61152] = t[61151] ^ n[61152];
assign t[61153] = t[61152] ^ n[61153];
assign t[61154] = t[61153] ^ n[61154];
assign t[61155] = t[61154] ^ n[61155];
assign t[61156] = t[61155] ^ n[61156];
assign t[61157] = t[61156] ^ n[61157];
assign t[61158] = t[61157] ^ n[61158];
assign t[61159] = t[61158] ^ n[61159];
assign t[61160] = t[61159] ^ n[61160];
assign t[61161] = t[61160] ^ n[61161];
assign t[61162] = t[61161] ^ n[61162];
assign t[61163] = t[61162] ^ n[61163];
assign t[61164] = t[61163] ^ n[61164];
assign t[61165] = t[61164] ^ n[61165];
assign t[61166] = t[61165] ^ n[61166];
assign t[61167] = t[61166] ^ n[61167];
assign t[61168] = t[61167] ^ n[61168];
assign t[61169] = t[61168] ^ n[61169];
assign t[61170] = t[61169] ^ n[61170];
assign t[61171] = t[61170] ^ n[61171];
assign t[61172] = t[61171] ^ n[61172];
assign t[61173] = t[61172] ^ n[61173];
assign t[61174] = t[61173] ^ n[61174];
assign t[61175] = t[61174] ^ n[61175];
assign t[61176] = t[61175] ^ n[61176];
assign t[61177] = t[61176] ^ n[61177];
assign t[61178] = t[61177] ^ n[61178];
assign t[61179] = t[61178] ^ n[61179];
assign t[61180] = t[61179] ^ n[61180];
assign t[61181] = t[61180] ^ n[61181];
assign t[61182] = t[61181] ^ n[61182];
assign t[61183] = t[61182] ^ n[61183];
assign t[61184] = t[61183] ^ n[61184];
assign t[61185] = t[61184] ^ n[61185];
assign t[61186] = t[61185] ^ n[61186];
assign t[61187] = t[61186] ^ n[61187];
assign t[61188] = t[61187] ^ n[61188];
assign t[61189] = t[61188] ^ n[61189];
assign t[61190] = t[61189] ^ n[61190];
assign t[61191] = t[61190] ^ n[61191];
assign t[61192] = t[61191] ^ n[61192];
assign t[61193] = t[61192] ^ n[61193];
assign t[61194] = t[61193] ^ n[61194];
assign t[61195] = t[61194] ^ n[61195];
assign t[61196] = t[61195] ^ n[61196];
assign t[61197] = t[61196] ^ n[61197];
assign t[61198] = t[61197] ^ n[61198];
assign t[61199] = t[61198] ^ n[61199];
assign t[61200] = t[61199] ^ n[61200];
assign t[61201] = t[61200] ^ n[61201];
assign t[61202] = t[61201] ^ n[61202];
assign t[61203] = t[61202] ^ n[61203];
assign t[61204] = t[61203] ^ n[61204];
assign t[61205] = t[61204] ^ n[61205];
assign t[61206] = t[61205] ^ n[61206];
assign t[61207] = t[61206] ^ n[61207];
assign t[61208] = t[61207] ^ n[61208];
assign t[61209] = t[61208] ^ n[61209];
assign t[61210] = t[61209] ^ n[61210];
assign t[61211] = t[61210] ^ n[61211];
assign t[61212] = t[61211] ^ n[61212];
assign t[61213] = t[61212] ^ n[61213];
assign t[61214] = t[61213] ^ n[61214];
assign t[61215] = t[61214] ^ n[61215];
assign t[61216] = t[61215] ^ n[61216];
assign t[61217] = t[61216] ^ n[61217];
assign t[61218] = t[61217] ^ n[61218];
assign t[61219] = t[61218] ^ n[61219];
assign t[61220] = t[61219] ^ n[61220];
assign t[61221] = t[61220] ^ n[61221];
assign t[61222] = t[61221] ^ n[61222];
assign t[61223] = t[61222] ^ n[61223];
assign t[61224] = t[61223] ^ n[61224];
assign t[61225] = t[61224] ^ n[61225];
assign t[61226] = t[61225] ^ n[61226];
assign t[61227] = t[61226] ^ n[61227];
assign t[61228] = t[61227] ^ n[61228];
assign t[61229] = t[61228] ^ n[61229];
assign t[61230] = t[61229] ^ n[61230];
assign t[61231] = t[61230] ^ n[61231];
assign t[61232] = t[61231] ^ n[61232];
assign t[61233] = t[61232] ^ n[61233];
assign t[61234] = t[61233] ^ n[61234];
assign t[61235] = t[61234] ^ n[61235];
assign t[61236] = t[61235] ^ n[61236];
assign t[61237] = t[61236] ^ n[61237];
assign t[61238] = t[61237] ^ n[61238];
assign t[61239] = t[61238] ^ n[61239];
assign t[61240] = t[61239] ^ n[61240];
assign t[61241] = t[61240] ^ n[61241];
assign t[61242] = t[61241] ^ n[61242];
assign t[61243] = t[61242] ^ n[61243];
assign t[61244] = t[61243] ^ n[61244];
assign t[61245] = t[61244] ^ n[61245];
assign t[61246] = t[61245] ^ n[61246];
assign t[61247] = t[61246] ^ n[61247];
assign t[61248] = t[61247] ^ n[61248];
assign t[61249] = t[61248] ^ n[61249];
assign t[61250] = t[61249] ^ n[61250];
assign t[61251] = t[61250] ^ n[61251];
assign t[61252] = t[61251] ^ n[61252];
assign t[61253] = t[61252] ^ n[61253];
assign t[61254] = t[61253] ^ n[61254];
assign t[61255] = t[61254] ^ n[61255];
assign t[61256] = t[61255] ^ n[61256];
assign t[61257] = t[61256] ^ n[61257];
assign t[61258] = t[61257] ^ n[61258];
assign t[61259] = t[61258] ^ n[61259];
assign t[61260] = t[61259] ^ n[61260];
assign t[61261] = t[61260] ^ n[61261];
assign t[61262] = t[61261] ^ n[61262];
assign t[61263] = t[61262] ^ n[61263];
assign t[61264] = t[61263] ^ n[61264];
assign t[61265] = t[61264] ^ n[61265];
assign t[61266] = t[61265] ^ n[61266];
assign t[61267] = t[61266] ^ n[61267];
assign t[61268] = t[61267] ^ n[61268];
assign t[61269] = t[61268] ^ n[61269];
assign t[61270] = t[61269] ^ n[61270];
assign t[61271] = t[61270] ^ n[61271];
assign t[61272] = t[61271] ^ n[61272];
assign t[61273] = t[61272] ^ n[61273];
assign t[61274] = t[61273] ^ n[61274];
assign t[61275] = t[61274] ^ n[61275];
assign t[61276] = t[61275] ^ n[61276];
assign t[61277] = t[61276] ^ n[61277];
assign t[61278] = t[61277] ^ n[61278];
assign t[61279] = t[61278] ^ n[61279];
assign t[61280] = t[61279] ^ n[61280];
assign t[61281] = t[61280] ^ n[61281];
assign t[61282] = t[61281] ^ n[61282];
assign t[61283] = t[61282] ^ n[61283];
assign t[61284] = t[61283] ^ n[61284];
assign t[61285] = t[61284] ^ n[61285];
assign t[61286] = t[61285] ^ n[61286];
assign t[61287] = t[61286] ^ n[61287];
assign t[61288] = t[61287] ^ n[61288];
assign t[61289] = t[61288] ^ n[61289];
assign t[61290] = t[61289] ^ n[61290];
assign t[61291] = t[61290] ^ n[61291];
assign t[61292] = t[61291] ^ n[61292];
assign t[61293] = t[61292] ^ n[61293];
assign t[61294] = t[61293] ^ n[61294];
assign t[61295] = t[61294] ^ n[61295];
assign t[61296] = t[61295] ^ n[61296];
assign t[61297] = t[61296] ^ n[61297];
assign t[61298] = t[61297] ^ n[61298];
assign t[61299] = t[61298] ^ n[61299];
assign t[61300] = t[61299] ^ n[61300];
assign t[61301] = t[61300] ^ n[61301];
assign t[61302] = t[61301] ^ n[61302];
assign t[61303] = t[61302] ^ n[61303];
assign t[61304] = t[61303] ^ n[61304];
assign t[61305] = t[61304] ^ n[61305];
assign t[61306] = t[61305] ^ n[61306];
assign t[61307] = t[61306] ^ n[61307];
assign t[61308] = t[61307] ^ n[61308];
assign t[61309] = t[61308] ^ n[61309];
assign t[61310] = t[61309] ^ n[61310];
assign t[61311] = t[61310] ^ n[61311];
assign t[61312] = t[61311] ^ n[61312];
assign t[61313] = t[61312] ^ n[61313];
assign t[61314] = t[61313] ^ n[61314];
assign t[61315] = t[61314] ^ n[61315];
assign t[61316] = t[61315] ^ n[61316];
assign t[61317] = t[61316] ^ n[61317];
assign t[61318] = t[61317] ^ n[61318];
assign t[61319] = t[61318] ^ n[61319];
assign t[61320] = t[61319] ^ n[61320];
assign t[61321] = t[61320] ^ n[61321];
assign t[61322] = t[61321] ^ n[61322];
assign t[61323] = t[61322] ^ n[61323];
assign t[61324] = t[61323] ^ n[61324];
assign t[61325] = t[61324] ^ n[61325];
assign t[61326] = t[61325] ^ n[61326];
assign t[61327] = t[61326] ^ n[61327];
assign t[61328] = t[61327] ^ n[61328];
assign t[61329] = t[61328] ^ n[61329];
assign t[61330] = t[61329] ^ n[61330];
assign t[61331] = t[61330] ^ n[61331];
assign t[61332] = t[61331] ^ n[61332];
assign t[61333] = t[61332] ^ n[61333];
assign t[61334] = t[61333] ^ n[61334];
assign t[61335] = t[61334] ^ n[61335];
assign t[61336] = t[61335] ^ n[61336];
assign t[61337] = t[61336] ^ n[61337];
assign t[61338] = t[61337] ^ n[61338];
assign t[61339] = t[61338] ^ n[61339];
assign t[61340] = t[61339] ^ n[61340];
assign t[61341] = t[61340] ^ n[61341];
assign t[61342] = t[61341] ^ n[61342];
assign t[61343] = t[61342] ^ n[61343];
assign t[61344] = t[61343] ^ n[61344];
assign t[61345] = t[61344] ^ n[61345];
assign t[61346] = t[61345] ^ n[61346];
assign t[61347] = t[61346] ^ n[61347];
assign t[61348] = t[61347] ^ n[61348];
assign t[61349] = t[61348] ^ n[61349];
assign t[61350] = t[61349] ^ n[61350];
assign t[61351] = t[61350] ^ n[61351];
assign t[61352] = t[61351] ^ n[61352];
assign t[61353] = t[61352] ^ n[61353];
assign t[61354] = t[61353] ^ n[61354];
assign t[61355] = t[61354] ^ n[61355];
assign t[61356] = t[61355] ^ n[61356];
assign t[61357] = t[61356] ^ n[61357];
assign t[61358] = t[61357] ^ n[61358];
assign t[61359] = t[61358] ^ n[61359];
assign t[61360] = t[61359] ^ n[61360];
assign t[61361] = t[61360] ^ n[61361];
assign t[61362] = t[61361] ^ n[61362];
assign t[61363] = t[61362] ^ n[61363];
assign t[61364] = t[61363] ^ n[61364];
assign t[61365] = t[61364] ^ n[61365];
assign t[61366] = t[61365] ^ n[61366];
assign t[61367] = t[61366] ^ n[61367];
assign t[61368] = t[61367] ^ n[61368];
assign t[61369] = t[61368] ^ n[61369];
assign t[61370] = t[61369] ^ n[61370];
assign t[61371] = t[61370] ^ n[61371];
assign t[61372] = t[61371] ^ n[61372];
assign t[61373] = t[61372] ^ n[61373];
assign t[61374] = t[61373] ^ n[61374];
assign t[61375] = t[61374] ^ n[61375];
assign t[61376] = t[61375] ^ n[61376];
assign t[61377] = t[61376] ^ n[61377];
assign t[61378] = t[61377] ^ n[61378];
assign t[61379] = t[61378] ^ n[61379];
assign t[61380] = t[61379] ^ n[61380];
assign t[61381] = t[61380] ^ n[61381];
assign t[61382] = t[61381] ^ n[61382];
assign t[61383] = t[61382] ^ n[61383];
assign t[61384] = t[61383] ^ n[61384];
assign t[61385] = t[61384] ^ n[61385];
assign t[61386] = t[61385] ^ n[61386];
assign t[61387] = t[61386] ^ n[61387];
assign t[61388] = t[61387] ^ n[61388];
assign t[61389] = t[61388] ^ n[61389];
assign t[61390] = t[61389] ^ n[61390];
assign t[61391] = t[61390] ^ n[61391];
assign t[61392] = t[61391] ^ n[61392];
assign t[61393] = t[61392] ^ n[61393];
assign t[61394] = t[61393] ^ n[61394];
assign t[61395] = t[61394] ^ n[61395];
assign t[61396] = t[61395] ^ n[61396];
assign t[61397] = t[61396] ^ n[61397];
assign t[61398] = t[61397] ^ n[61398];
assign t[61399] = t[61398] ^ n[61399];
assign t[61400] = t[61399] ^ n[61400];
assign t[61401] = t[61400] ^ n[61401];
assign t[61402] = t[61401] ^ n[61402];
assign t[61403] = t[61402] ^ n[61403];
assign t[61404] = t[61403] ^ n[61404];
assign t[61405] = t[61404] ^ n[61405];
assign t[61406] = t[61405] ^ n[61406];
assign t[61407] = t[61406] ^ n[61407];
assign t[61408] = t[61407] ^ n[61408];
assign t[61409] = t[61408] ^ n[61409];
assign t[61410] = t[61409] ^ n[61410];
assign t[61411] = t[61410] ^ n[61411];
assign t[61412] = t[61411] ^ n[61412];
assign t[61413] = t[61412] ^ n[61413];
assign t[61414] = t[61413] ^ n[61414];
assign t[61415] = t[61414] ^ n[61415];
assign t[61416] = t[61415] ^ n[61416];
assign t[61417] = t[61416] ^ n[61417];
assign t[61418] = t[61417] ^ n[61418];
assign t[61419] = t[61418] ^ n[61419];
assign t[61420] = t[61419] ^ n[61420];
assign t[61421] = t[61420] ^ n[61421];
assign t[61422] = t[61421] ^ n[61422];
assign t[61423] = t[61422] ^ n[61423];
assign t[61424] = t[61423] ^ n[61424];
assign t[61425] = t[61424] ^ n[61425];
assign t[61426] = t[61425] ^ n[61426];
assign t[61427] = t[61426] ^ n[61427];
assign t[61428] = t[61427] ^ n[61428];
assign t[61429] = t[61428] ^ n[61429];
assign t[61430] = t[61429] ^ n[61430];
assign t[61431] = t[61430] ^ n[61431];
assign t[61432] = t[61431] ^ n[61432];
assign t[61433] = t[61432] ^ n[61433];
assign t[61434] = t[61433] ^ n[61434];
assign t[61435] = t[61434] ^ n[61435];
assign t[61436] = t[61435] ^ n[61436];
assign t[61437] = t[61436] ^ n[61437];
assign t[61438] = t[61437] ^ n[61438];
assign t[61439] = t[61438] ^ n[61439];
assign t[61440] = t[61439] ^ n[61440];
assign t[61441] = t[61440] ^ n[61441];
assign t[61442] = t[61441] ^ n[61442];
assign t[61443] = t[61442] ^ n[61443];
assign t[61444] = t[61443] ^ n[61444];
assign t[61445] = t[61444] ^ n[61445];
assign t[61446] = t[61445] ^ n[61446];
assign t[61447] = t[61446] ^ n[61447];
assign t[61448] = t[61447] ^ n[61448];
assign t[61449] = t[61448] ^ n[61449];
assign t[61450] = t[61449] ^ n[61450];
assign t[61451] = t[61450] ^ n[61451];
assign t[61452] = t[61451] ^ n[61452];
assign t[61453] = t[61452] ^ n[61453];
assign t[61454] = t[61453] ^ n[61454];
assign t[61455] = t[61454] ^ n[61455];
assign t[61456] = t[61455] ^ n[61456];
assign t[61457] = t[61456] ^ n[61457];
assign t[61458] = t[61457] ^ n[61458];
assign t[61459] = t[61458] ^ n[61459];
assign t[61460] = t[61459] ^ n[61460];
assign t[61461] = t[61460] ^ n[61461];
assign t[61462] = t[61461] ^ n[61462];
assign t[61463] = t[61462] ^ n[61463];
assign t[61464] = t[61463] ^ n[61464];
assign t[61465] = t[61464] ^ n[61465];
assign t[61466] = t[61465] ^ n[61466];
assign t[61467] = t[61466] ^ n[61467];
assign t[61468] = t[61467] ^ n[61468];
assign t[61469] = t[61468] ^ n[61469];
assign t[61470] = t[61469] ^ n[61470];
assign t[61471] = t[61470] ^ n[61471];
assign t[61472] = t[61471] ^ n[61472];
assign t[61473] = t[61472] ^ n[61473];
assign t[61474] = t[61473] ^ n[61474];
assign t[61475] = t[61474] ^ n[61475];
assign t[61476] = t[61475] ^ n[61476];
assign t[61477] = t[61476] ^ n[61477];
assign t[61478] = t[61477] ^ n[61478];
assign t[61479] = t[61478] ^ n[61479];
assign t[61480] = t[61479] ^ n[61480];
assign t[61481] = t[61480] ^ n[61481];
assign t[61482] = t[61481] ^ n[61482];
assign t[61483] = t[61482] ^ n[61483];
assign t[61484] = t[61483] ^ n[61484];
assign t[61485] = t[61484] ^ n[61485];
assign t[61486] = t[61485] ^ n[61486];
assign t[61487] = t[61486] ^ n[61487];
assign t[61488] = t[61487] ^ n[61488];
assign t[61489] = t[61488] ^ n[61489];
assign t[61490] = t[61489] ^ n[61490];
assign t[61491] = t[61490] ^ n[61491];
assign t[61492] = t[61491] ^ n[61492];
assign t[61493] = t[61492] ^ n[61493];
assign t[61494] = t[61493] ^ n[61494];
assign t[61495] = t[61494] ^ n[61495];
assign t[61496] = t[61495] ^ n[61496];
assign t[61497] = t[61496] ^ n[61497];
assign t[61498] = t[61497] ^ n[61498];
assign t[61499] = t[61498] ^ n[61499];
assign t[61500] = t[61499] ^ n[61500];
assign t[61501] = t[61500] ^ n[61501];
assign t[61502] = t[61501] ^ n[61502];
assign t[61503] = t[61502] ^ n[61503];
assign t[61504] = t[61503] ^ n[61504];
assign t[61505] = t[61504] ^ n[61505];
assign t[61506] = t[61505] ^ n[61506];
assign t[61507] = t[61506] ^ n[61507];
assign t[61508] = t[61507] ^ n[61508];
assign t[61509] = t[61508] ^ n[61509];
assign t[61510] = t[61509] ^ n[61510];
assign t[61511] = t[61510] ^ n[61511];
assign t[61512] = t[61511] ^ n[61512];
assign t[61513] = t[61512] ^ n[61513];
assign t[61514] = t[61513] ^ n[61514];
assign t[61515] = t[61514] ^ n[61515];
assign t[61516] = t[61515] ^ n[61516];
assign t[61517] = t[61516] ^ n[61517];
assign t[61518] = t[61517] ^ n[61518];
assign t[61519] = t[61518] ^ n[61519];
assign t[61520] = t[61519] ^ n[61520];
assign t[61521] = t[61520] ^ n[61521];
assign t[61522] = t[61521] ^ n[61522];
assign t[61523] = t[61522] ^ n[61523];
assign t[61524] = t[61523] ^ n[61524];
assign t[61525] = t[61524] ^ n[61525];
assign t[61526] = t[61525] ^ n[61526];
assign t[61527] = t[61526] ^ n[61527];
assign t[61528] = t[61527] ^ n[61528];
assign t[61529] = t[61528] ^ n[61529];
assign t[61530] = t[61529] ^ n[61530];
assign t[61531] = t[61530] ^ n[61531];
assign t[61532] = t[61531] ^ n[61532];
assign t[61533] = t[61532] ^ n[61533];
assign t[61534] = t[61533] ^ n[61534];
assign t[61535] = t[61534] ^ n[61535];
assign t[61536] = t[61535] ^ n[61536];
assign t[61537] = t[61536] ^ n[61537];
assign t[61538] = t[61537] ^ n[61538];
assign t[61539] = t[61538] ^ n[61539];
assign t[61540] = t[61539] ^ n[61540];
assign t[61541] = t[61540] ^ n[61541];
assign t[61542] = t[61541] ^ n[61542];
assign t[61543] = t[61542] ^ n[61543];
assign t[61544] = t[61543] ^ n[61544];
assign t[61545] = t[61544] ^ n[61545];
assign t[61546] = t[61545] ^ n[61546];
assign t[61547] = t[61546] ^ n[61547];
assign t[61548] = t[61547] ^ n[61548];
assign t[61549] = t[61548] ^ n[61549];
assign t[61550] = t[61549] ^ n[61550];
assign t[61551] = t[61550] ^ n[61551];
assign t[61552] = t[61551] ^ n[61552];
assign t[61553] = t[61552] ^ n[61553];
assign t[61554] = t[61553] ^ n[61554];
assign t[61555] = t[61554] ^ n[61555];
assign t[61556] = t[61555] ^ n[61556];
assign t[61557] = t[61556] ^ n[61557];
assign t[61558] = t[61557] ^ n[61558];
assign t[61559] = t[61558] ^ n[61559];
assign t[61560] = t[61559] ^ n[61560];
assign t[61561] = t[61560] ^ n[61561];
assign t[61562] = t[61561] ^ n[61562];
assign t[61563] = t[61562] ^ n[61563];
assign t[61564] = t[61563] ^ n[61564];
assign t[61565] = t[61564] ^ n[61565];
assign t[61566] = t[61565] ^ n[61566];
assign t[61567] = t[61566] ^ n[61567];
assign t[61568] = t[61567] ^ n[61568];
assign t[61569] = t[61568] ^ n[61569];
assign t[61570] = t[61569] ^ n[61570];
assign t[61571] = t[61570] ^ n[61571];
assign t[61572] = t[61571] ^ n[61572];
assign t[61573] = t[61572] ^ n[61573];
assign t[61574] = t[61573] ^ n[61574];
assign t[61575] = t[61574] ^ n[61575];
assign t[61576] = t[61575] ^ n[61576];
assign t[61577] = t[61576] ^ n[61577];
assign t[61578] = t[61577] ^ n[61578];
assign t[61579] = t[61578] ^ n[61579];
assign t[61580] = t[61579] ^ n[61580];
assign t[61581] = t[61580] ^ n[61581];
assign t[61582] = t[61581] ^ n[61582];
assign t[61583] = t[61582] ^ n[61583];
assign t[61584] = t[61583] ^ n[61584];
assign t[61585] = t[61584] ^ n[61585];
assign t[61586] = t[61585] ^ n[61586];
assign t[61587] = t[61586] ^ n[61587];
assign t[61588] = t[61587] ^ n[61588];
assign t[61589] = t[61588] ^ n[61589];
assign t[61590] = t[61589] ^ n[61590];
assign t[61591] = t[61590] ^ n[61591];
assign t[61592] = t[61591] ^ n[61592];
assign t[61593] = t[61592] ^ n[61593];
assign t[61594] = t[61593] ^ n[61594];
assign t[61595] = t[61594] ^ n[61595];
assign t[61596] = t[61595] ^ n[61596];
assign t[61597] = t[61596] ^ n[61597];
assign t[61598] = t[61597] ^ n[61598];
assign t[61599] = t[61598] ^ n[61599];
assign t[61600] = t[61599] ^ n[61600];
assign t[61601] = t[61600] ^ n[61601];
assign t[61602] = t[61601] ^ n[61602];
assign t[61603] = t[61602] ^ n[61603];
assign t[61604] = t[61603] ^ n[61604];
assign t[61605] = t[61604] ^ n[61605];
assign t[61606] = t[61605] ^ n[61606];
assign t[61607] = t[61606] ^ n[61607];
assign t[61608] = t[61607] ^ n[61608];
assign t[61609] = t[61608] ^ n[61609];
assign t[61610] = t[61609] ^ n[61610];
assign t[61611] = t[61610] ^ n[61611];
assign t[61612] = t[61611] ^ n[61612];
assign t[61613] = t[61612] ^ n[61613];
assign t[61614] = t[61613] ^ n[61614];
assign t[61615] = t[61614] ^ n[61615];
assign t[61616] = t[61615] ^ n[61616];
assign t[61617] = t[61616] ^ n[61617];
assign t[61618] = t[61617] ^ n[61618];
assign t[61619] = t[61618] ^ n[61619];
assign t[61620] = t[61619] ^ n[61620];
assign t[61621] = t[61620] ^ n[61621];
assign t[61622] = t[61621] ^ n[61622];
assign t[61623] = t[61622] ^ n[61623];
assign t[61624] = t[61623] ^ n[61624];
assign t[61625] = t[61624] ^ n[61625];
assign t[61626] = t[61625] ^ n[61626];
assign t[61627] = t[61626] ^ n[61627];
assign t[61628] = t[61627] ^ n[61628];
assign t[61629] = t[61628] ^ n[61629];
assign t[61630] = t[61629] ^ n[61630];
assign t[61631] = t[61630] ^ n[61631];
assign t[61632] = t[61631] ^ n[61632];
assign t[61633] = t[61632] ^ n[61633];
assign t[61634] = t[61633] ^ n[61634];
assign t[61635] = t[61634] ^ n[61635];
assign t[61636] = t[61635] ^ n[61636];
assign t[61637] = t[61636] ^ n[61637];
assign t[61638] = t[61637] ^ n[61638];
assign t[61639] = t[61638] ^ n[61639];
assign t[61640] = t[61639] ^ n[61640];
assign t[61641] = t[61640] ^ n[61641];
assign t[61642] = t[61641] ^ n[61642];
assign t[61643] = t[61642] ^ n[61643];
assign t[61644] = t[61643] ^ n[61644];
assign t[61645] = t[61644] ^ n[61645];
assign t[61646] = t[61645] ^ n[61646];
assign t[61647] = t[61646] ^ n[61647];
assign t[61648] = t[61647] ^ n[61648];
assign t[61649] = t[61648] ^ n[61649];
assign t[61650] = t[61649] ^ n[61650];
assign t[61651] = t[61650] ^ n[61651];
assign t[61652] = t[61651] ^ n[61652];
assign t[61653] = t[61652] ^ n[61653];
assign t[61654] = t[61653] ^ n[61654];
assign t[61655] = t[61654] ^ n[61655];
assign t[61656] = t[61655] ^ n[61656];
assign t[61657] = t[61656] ^ n[61657];
assign t[61658] = t[61657] ^ n[61658];
assign t[61659] = t[61658] ^ n[61659];
assign t[61660] = t[61659] ^ n[61660];
assign t[61661] = t[61660] ^ n[61661];
assign t[61662] = t[61661] ^ n[61662];
assign t[61663] = t[61662] ^ n[61663];
assign t[61664] = t[61663] ^ n[61664];
assign t[61665] = t[61664] ^ n[61665];
assign t[61666] = t[61665] ^ n[61666];
assign t[61667] = t[61666] ^ n[61667];
assign t[61668] = t[61667] ^ n[61668];
assign t[61669] = t[61668] ^ n[61669];
assign t[61670] = t[61669] ^ n[61670];
assign t[61671] = t[61670] ^ n[61671];
assign t[61672] = t[61671] ^ n[61672];
assign t[61673] = t[61672] ^ n[61673];
assign t[61674] = t[61673] ^ n[61674];
assign t[61675] = t[61674] ^ n[61675];
assign t[61676] = t[61675] ^ n[61676];
assign t[61677] = t[61676] ^ n[61677];
assign t[61678] = t[61677] ^ n[61678];
assign t[61679] = t[61678] ^ n[61679];
assign t[61680] = t[61679] ^ n[61680];
assign t[61681] = t[61680] ^ n[61681];
assign t[61682] = t[61681] ^ n[61682];
assign t[61683] = t[61682] ^ n[61683];
assign t[61684] = t[61683] ^ n[61684];
assign t[61685] = t[61684] ^ n[61685];
assign t[61686] = t[61685] ^ n[61686];
assign t[61687] = t[61686] ^ n[61687];
assign t[61688] = t[61687] ^ n[61688];
assign t[61689] = t[61688] ^ n[61689];
assign t[61690] = t[61689] ^ n[61690];
assign t[61691] = t[61690] ^ n[61691];
assign t[61692] = t[61691] ^ n[61692];
assign t[61693] = t[61692] ^ n[61693];
assign t[61694] = t[61693] ^ n[61694];
assign t[61695] = t[61694] ^ n[61695];
assign t[61696] = t[61695] ^ n[61696];
assign t[61697] = t[61696] ^ n[61697];
assign t[61698] = t[61697] ^ n[61698];
assign t[61699] = t[61698] ^ n[61699];
assign t[61700] = t[61699] ^ n[61700];
assign t[61701] = t[61700] ^ n[61701];
assign t[61702] = t[61701] ^ n[61702];
assign t[61703] = t[61702] ^ n[61703];
assign t[61704] = t[61703] ^ n[61704];
assign t[61705] = t[61704] ^ n[61705];
assign t[61706] = t[61705] ^ n[61706];
assign t[61707] = t[61706] ^ n[61707];
assign t[61708] = t[61707] ^ n[61708];
assign t[61709] = t[61708] ^ n[61709];
assign t[61710] = t[61709] ^ n[61710];
assign t[61711] = t[61710] ^ n[61711];
assign t[61712] = t[61711] ^ n[61712];
assign t[61713] = t[61712] ^ n[61713];
assign t[61714] = t[61713] ^ n[61714];
assign t[61715] = t[61714] ^ n[61715];
assign t[61716] = t[61715] ^ n[61716];
assign t[61717] = t[61716] ^ n[61717];
assign t[61718] = t[61717] ^ n[61718];
assign t[61719] = t[61718] ^ n[61719];
assign t[61720] = t[61719] ^ n[61720];
assign t[61721] = t[61720] ^ n[61721];
assign t[61722] = t[61721] ^ n[61722];
assign t[61723] = t[61722] ^ n[61723];
assign t[61724] = t[61723] ^ n[61724];
assign t[61725] = t[61724] ^ n[61725];
assign t[61726] = t[61725] ^ n[61726];
assign t[61727] = t[61726] ^ n[61727];
assign t[61728] = t[61727] ^ n[61728];
assign t[61729] = t[61728] ^ n[61729];
assign t[61730] = t[61729] ^ n[61730];
assign t[61731] = t[61730] ^ n[61731];
assign t[61732] = t[61731] ^ n[61732];
assign t[61733] = t[61732] ^ n[61733];
assign t[61734] = t[61733] ^ n[61734];
assign t[61735] = t[61734] ^ n[61735];
assign t[61736] = t[61735] ^ n[61736];
assign t[61737] = t[61736] ^ n[61737];
assign t[61738] = t[61737] ^ n[61738];
assign t[61739] = t[61738] ^ n[61739];
assign t[61740] = t[61739] ^ n[61740];
assign t[61741] = t[61740] ^ n[61741];
assign t[61742] = t[61741] ^ n[61742];
assign t[61743] = t[61742] ^ n[61743];
assign t[61744] = t[61743] ^ n[61744];
assign t[61745] = t[61744] ^ n[61745];
assign t[61746] = t[61745] ^ n[61746];
assign t[61747] = t[61746] ^ n[61747];
assign t[61748] = t[61747] ^ n[61748];
assign t[61749] = t[61748] ^ n[61749];
assign t[61750] = t[61749] ^ n[61750];
assign t[61751] = t[61750] ^ n[61751];
assign t[61752] = t[61751] ^ n[61752];
assign t[61753] = t[61752] ^ n[61753];
assign t[61754] = t[61753] ^ n[61754];
assign t[61755] = t[61754] ^ n[61755];
assign t[61756] = t[61755] ^ n[61756];
assign t[61757] = t[61756] ^ n[61757];
assign t[61758] = t[61757] ^ n[61758];
assign t[61759] = t[61758] ^ n[61759];
assign t[61760] = t[61759] ^ n[61760];
assign t[61761] = t[61760] ^ n[61761];
assign t[61762] = t[61761] ^ n[61762];
assign t[61763] = t[61762] ^ n[61763];
assign t[61764] = t[61763] ^ n[61764];
assign t[61765] = t[61764] ^ n[61765];
assign t[61766] = t[61765] ^ n[61766];
assign t[61767] = t[61766] ^ n[61767];
assign t[61768] = t[61767] ^ n[61768];
assign t[61769] = t[61768] ^ n[61769];
assign t[61770] = t[61769] ^ n[61770];
assign t[61771] = t[61770] ^ n[61771];
assign t[61772] = t[61771] ^ n[61772];
assign t[61773] = t[61772] ^ n[61773];
assign t[61774] = t[61773] ^ n[61774];
assign t[61775] = t[61774] ^ n[61775];
assign t[61776] = t[61775] ^ n[61776];
assign t[61777] = t[61776] ^ n[61777];
assign t[61778] = t[61777] ^ n[61778];
assign t[61779] = t[61778] ^ n[61779];
assign t[61780] = t[61779] ^ n[61780];
assign t[61781] = t[61780] ^ n[61781];
assign t[61782] = t[61781] ^ n[61782];
assign t[61783] = t[61782] ^ n[61783];
assign t[61784] = t[61783] ^ n[61784];
assign t[61785] = t[61784] ^ n[61785];
assign t[61786] = t[61785] ^ n[61786];
assign t[61787] = t[61786] ^ n[61787];
assign t[61788] = t[61787] ^ n[61788];
assign t[61789] = t[61788] ^ n[61789];
assign t[61790] = t[61789] ^ n[61790];
assign t[61791] = t[61790] ^ n[61791];
assign t[61792] = t[61791] ^ n[61792];
assign t[61793] = t[61792] ^ n[61793];
assign t[61794] = t[61793] ^ n[61794];
assign t[61795] = t[61794] ^ n[61795];
assign t[61796] = t[61795] ^ n[61796];
assign t[61797] = t[61796] ^ n[61797];
assign t[61798] = t[61797] ^ n[61798];
assign t[61799] = t[61798] ^ n[61799];
assign t[61800] = t[61799] ^ n[61800];
assign t[61801] = t[61800] ^ n[61801];
assign t[61802] = t[61801] ^ n[61802];
assign t[61803] = t[61802] ^ n[61803];
assign t[61804] = t[61803] ^ n[61804];
assign t[61805] = t[61804] ^ n[61805];
assign t[61806] = t[61805] ^ n[61806];
assign t[61807] = t[61806] ^ n[61807];
assign t[61808] = t[61807] ^ n[61808];
assign t[61809] = t[61808] ^ n[61809];
assign t[61810] = t[61809] ^ n[61810];
assign t[61811] = t[61810] ^ n[61811];
assign t[61812] = t[61811] ^ n[61812];
assign t[61813] = t[61812] ^ n[61813];
assign t[61814] = t[61813] ^ n[61814];
assign t[61815] = t[61814] ^ n[61815];
assign t[61816] = t[61815] ^ n[61816];
assign t[61817] = t[61816] ^ n[61817];
assign t[61818] = t[61817] ^ n[61818];
assign t[61819] = t[61818] ^ n[61819];
assign t[61820] = t[61819] ^ n[61820];
assign t[61821] = t[61820] ^ n[61821];
assign t[61822] = t[61821] ^ n[61822];
assign t[61823] = t[61822] ^ n[61823];
assign t[61824] = t[61823] ^ n[61824];
assign t[61825] = t[61824] ^ n[61825];
assign t[61826] = t[61825] ^ n[61826];
assign t[61827] = t[61826] ^ n[61827];
assign t[61828] = t[61827] ^ n[61828];
assign t[61829] = t[61828] ^ n[61829];
assign t[61830] = t[61829] ^ n[61830];
assign t[61831] = t[61830] ^ n[61831];
assign t[61832] = t[61831] ^ n[61832];
assign t[61833] = t[61832] ^ n[61833];
assign t[61834] = t[61833] ^ n[61834];
assign t[61835] = t[61834] ^ n[61835];
assign t[61836] = t[61835] ^ n[61836];
assign t[61837] = t[61836] ^ n[61837];
assign t[61838] = t[61837] ^ n[61838];
assign t[61839] = t[61838] ^ n[61839];
assign t[61840] = t[61839] ^ n[61840];
assign t[61841] = t[61840] ^ n[61841];
assign t[61842] = t[61841] ^ n[61842];
assign t[61843] = t[61842] ^ n[61843];
assign t[61844] = t[61843] ^ n[61844];
assign t[61845] = t[61844] ^ n[61845];
assign t[61846] = t[61845] ^ n[61846];
assign t[61847] = t[61846] ^ n[61847];
assign t[61848] = t[61847] ^ n[61848];
assign t[61849] = t[61848] ^ n[61849];
assign t[61850] = t[61849] ^ n[61850];
assign t[61851] = t[61850] ^ n[61851];
assign t[61852] = t[61851] ^ n[61852];
assign t[61853] = t[61852] ^ n[61853];
assign t[61854] = t[61853] ^ n[61854];
assign t[61855] = t[61854] ^ n[61855];
assign t[61856] = t[61855] ^ n[61856];
assign t[61857] = t[61856] ^ n[61857];
assign t[61858] = t[61857] ^ n[61858];
assign t[61859] = t[61858] ^ n[61859];
assign t[61860] = t[61859] ^ n[61860];
assign t[61861] = t[61860] ^ n[61861];
assign t[61862] = t[61861] ^ n[61862];
assign t[61863] = t[61862] ^ n[61863];
assign t[61864] = t[61863] ^ n[61864];
assign t[61865] = t[61864] ^ n[61865];
assign t[61866] = t[61865] ^ n[61866];
assign t[61867] = t[61866] ^ n[61867];
assign t[61868] = t[61867] ^ n[61868];
assign t[61869] = t[61868] ^ n[61869];
assign t[61870] = t[61869] ^ n[61870];
assign t[61871] = t[61870] ^ n[61871];
assign t[61872] = t[61871] ^ n[61872];
assign t[61873] = t[61872] ^ n[61873];
assign t[61874] = t[61873] ^ n[61874];
assign t[61875] = t[61874] ^ n[61875];
assign t[61876] = t[61875] ^ n[61876];
assign t[61877] = t[61876] ^ n[61877];
assign t[61878] = t[61877] ^ n[61878];
assign t[61879] = t[61878] ^ n[61879];
assign t[61880] = t[61879] ^ n[61880];
assign t[61881] = t[61880] ^ n[61881];
assign t[61882] = t[61881] ^ n[61882];
assign t[61883] = t[61882] ^ n[61883];
assign t[61884] = t[61883] ^ n[61884];
assign t[61885] = t[61884] ^ n[61885];
assign t[61886] = t[61885] ^ n[61886];
assign t[61887] = t[61886] ^ n[61887];
assign t[61888] = t[61887] ^ n[61888];
assign t[61889] = t[61888] ^ n[61889];
assign t[61890] = t[61889] ^ n[61890];
assign t[61891] = t[61890] ^ n[61891];
assign t[61892] = t[61891] ^ n[61892];
assign t[61893] = t[61892] ^ n[61893];
assign t[61894] = t[61893] ^ n[61894];
assign t[61895] = t[61894] ^ n[61895];
assign t[61896] = t[61895] ^ n[61896];
assign t[61897] = t[61896] ^ n[61897];
assign t[61898] = t[61897] ^ n[61898];
assign t[61899] = t[61898] ^ n[61899];
assign t[61900] = t[61899] ^ n[61900];
assign t[61901] = t[61900] ^ n[61901];
assign t[61902] = t[61901] ^ n[61902];
assign t[61903] = t[61902] ^ n[61903];
assign t[61904] = t[61903] ^ n[61904];
assign t[61905] = t[61904] ^ n[61905];
assign t[61906] = t[61905] ^ n[61906];
assign t[61907] = t[61906] ^ n[61907];
assign t[61908] = t[61907] ^ n[61908];
assign t[61909] = t[61908] ^ n[61909];
assign t[61910] = t[61909] ^ n[61910];
assign t[61911] = t[61910] ^ n[61911];
assign t[61912] = t[61911] ^ n[61912];
assign t[61913] = t[61912] ^ n[61913];
assign t[61914] = t[61913] ^ n[61914];
assign t[61915] = t[61914] ^ n[61915];
assign t[61916] = t[61915] ^ n[61916];
assign t[61917] = t[61916] ^ n[61917];
assign t[61918] = t[61917] ^ n[61918];
assign t[61919] = t[61918] ^ n[61919];
assign t[61920] = t[61919] ^ n[61920];
assign t[61921] = t[61920] ^ n[61921];
assign t[61922] = t[61921] ^ n[61922];
assign t[61923] = t[61922] ^ n[61923];
assign t[61924] = t[61923] ^ n[61924];
assign t[61925] = t[61924] ^ n[61925];
assign t[61926] = t[61925] ^ n[61926];
assign t[61927] = t[61926] ^ n[61927];
assign t[61928] = t[61927] ^ n[61928];
assign t[61929] = t[61928] ^ n[61929];
assign t[61930] = t[61929] ^ n[61930];
assign t[61931] = t[61930] ^ n[61931];
assign t[61932] = t[61931] ^ n[61932];
assign t[61933] = t[61932] ^ n[61933];
assign t[61934] = t[61933] ^ n[61934];
assign t[61935] = t[61934] ^ n[61935];
assign t[61936] = t[61935] ^ n[61936];
assign t[61937] = t[61936] ^ n[61937];
assign t[61938] = t[61937] ^ n[61938];
assign t[61939] = t[61938] ^ n[61939];
assign t[61940] = t[61939] ^ n[61940];
assign t[61941] = t[61940] ^ n[61941];
assign t[61942] = t[61941] ^ n[61942];
assign t[61943] = t[61942] ^ n[61943];
assign t[61944] = t[61943] ^ n[61944];
assign t[61945] = t[61944] ^ n[61945];
assign t[61946] = t[61945] ^ n[61946];
assign t[61947] = t[61946] ^ n[61947];
assign t[61948] = t[61947] ^ n[61948];
assign t[61949] = t[61948] ^ n[61949];
assign t[61950] = t[61949] ^ n[61950];
assign t[61951] = t[61950] ^ n[61951];
assign t[61952] = t[61951] ^ n[61952];
assign t[61953] = t[61952] ^ n[61953];
assign t[61954] = t[61953] ^ n[61954];
assign t[61955] = t[61954] ^ n[61955];
assign t[61956] = t[61955] ^ n[61956];
assign t[61957] = t[61956] ^ n[61957];
assign t[61958] = t[61957] ^ n[61958];
assign t[61959] = t[61958] ^ n[61959];
assign t[61960] = t[61959] ^ n[61960];
assign t[61961] = t[61960] ^ n[61961];
assign t[61962] = t[61961] ^ n[61962];
assign t[61963] = t[61962] ^ n[61963];
assign t[61964] = t[61963] ^ n[61964];
assign t[61965] = t[61964] ^ n[61965];
assign t[61966] = t[61965] ^ n[61966];
assign t[61967] = t[61966] ^ n[61967];
assign t[61968] = t[61967] ^ n[61968];
assign t[61969] = t[61968] ^ n[61969];
assign t[61970] = t[61969] ^ n[61970];
assign t[61971] = t[61970] ^ n[61971];
assign t[61972] = t[61971] ^ n[61972];
assign t[61973] = t[61972] ^ n[61973];
assign t[61974] = t[61973] ^ n[61974];
assign t[61975] = t[61974] ^ n[61975];
assign t[61976] = t[61975] ^ n[61976];
assign t[61977] = t[61976] ^ n[61977];
assign t[61978] = t[61977] ^ n[61978];
assign t[61979] = t[61978] ^ n[61979];
assign t[61980] = t[61979] ^ n[61980];
assign t[61981] = t[61980] ^ n[61981];
assign t[61982] = t[61981] ^ n[61982];
assign t[61983] = t[61982] ^ n[61983];
assign t[61984] = t[61983] ^ n[61984];
assign t[61985] = t[61984] ^ n[61985];
assign t[61986] = t[61985] ^ n[61986];
assign t[61987] = t[61986] ^ n[61987];
assign t[61988] = t[61987] ^ n[61988];
assign t[61989] = t[61988] ^ n[61989];
assign t[61990] = t[61989] ^ n[61990];
assign t[61991] = t[61990] ^ n[61991];
assign t[61992] = t[61991] ^ n[61992];
assign t[61993] = t[61992] ^ n[61993];
assign t[61994] = t[61993] ^ n[61994];
assign t[61995] = t[61994] ^ n[61995];
assign t[61996] = t[61995] ^ n[61996];
assign t[61997] = t[61996] ^ n[61997];
assign t[61998] = t[61997] ^ n[61998];
assign t[61999] = t[61998] ^ n[61999];
assign t[62000] = t[61999] ^ n[62000];
assign t[62001] = t[62000] ^ n[62001];
assign t[62002] = t[62001] ^ n[62002];
assign t[62003] = t[62002] ^ n[62003];
assign t[62004] = t[62003] ^ n[62004];
assign t[62005] = t[62004] ^ n[62005];
assign t[62006] = t[62005] ^ n[62006];
assign t[62007] = t[62006] ^ n[62007];
assign t[62008] = t[62007] ^ n[62008];
assign t[62009] = t[62008] ^ n[62009];
assign t[62010] = t[62009] ^ n[62010];
assign t[62011] = t[62010] ^ n[62011];
assign t[62012] = t[62011] ^ n[62012];
assign t[62013] = t[62012] ^ n[62013];
assign t[62014] = t[62013] ^ n[62014];
assign t[62015] = t[62014] ^ n[62015];
assign t[62016] = t[62015] ^ n[62016];
assign t[62017] = t[62016] ^ n[62017];
assign t[62018] = t[62017] ^ n[62018];
assign t[62019] = t[62018] ^ n[62019];
assign t[62020] = t[62019] ^ n[62020];
assign t[62021] = t[62020] ^ n[62021];
assign t[62022] = t[62021] ^ n[62022];
assign t[62023] = t[62022] ^ n[62023];
assign t[62024] = t[62023] ^ n[62024];
assign t[62025] = t[62024] ^ n[62025];
assign t[62026] = t[62025] ^ n[62026];
assign t[62027] = t[62026] ^ n[62027];
assign t[62028] = t[62027] ^ n[62028];
assign t[62029] = t[62028] ^ n[62029];
assign t[62030] = t[62029] ^ n[62030];
assign t[62031] = t[62030] ^ n[62031];
assign t[62032] = t[62031] ^ n[62032];
assign t[62033] = t[62032] ^ n[62033];
assign t[62034] = t[62033] ^ n[62034];
assign t[62035] = t[62034] ^ n[62035];
assign t[62036] = t[62035] ^ n[62036];
assign t[62037] = t[62036] ^ n[62037];
assign t[62038] = t[62037] ^ n[62038];
assign t[62039] = t[62038] ^ n[62039];
assign t[62040] = t[62039] ^ n[62040];
assign t[62041] = t[62040] ^ n[62041];
assign t[62042] = t[62041] ^ n[62042];
assign t[62043] = t[62042] ^ n[62043];
assign t[62044] = t[62043] ^ n[62044];
assign t[62045] = t[62044] ^ n[62045];
assign t[62046] = t[62045] ^ n[62046];
assign t[62047] = t[62046] ^ n[62047];
assign t[62048] = t[62047] ^ n[62048];
assign t[62049] = t[62048] ^ n[62049];
assign t[62050] = t[62049] ^ n[62050];
assign t[62051] = t[62050] ^ n[62051];
assign t[62052] = t[62051] ^ n[62052];
assign t[62053] = t[62052] ^ n[62053];
assign t[62054] = t[62053] ^ n[62054];
assign t[62055] = t[62054] ^ n[62055];
assign t[62056] = t[62055] ^ n[62056];
assign t[62057] = t[62056] ^ n[62057];
assign t[62058] = t[62057] ^ n[62058];
assign t[62059] = t[62058] ^ n[62059];
assign t[62060] = t[62059] ^ n[62060];
assign t[62061] = t[62060] ^ n[62061];
assign t[62062] = t[62061] ^ n[62062];
assign t[62063] = t[62062] ^ n[62063];
assign t[62064] = t[62063] ^ n[62064];
assign t[62065] = t[62064] ^ n[62065];
assign t[62066] = t[62065] ^ n[62066];
assign t[62067] = t[62066] ^ n[62067];
assign t[62068] = t[62067] ^ n[62068];
assign t[62069] = t[62068] ^ n[62069];
assign t[62070] = t[62069] ^ n[62070];
assign t[62071] = t[62070] ^ n[62071];
assign t[62072] = t[62071] ^ n[62072];
assign t[62073] = t[62072] ^ n[62073];
assign t[62074] = t[62073] ^ n[62074];
assign t[62075] = t[62074] ^ n[62075];
assign t[62076] = t[62075] ^ n[62076];
assign t[62077] = t[62076] ^ n[62077];
assign t[62078] = t[62077] ^ n[62078];
assign t[62079] = t[62078] ^ n[62079];
assign t[62080] = t[62079] ^ n[62080];
assign t[62081] = t[62080] ^ n[62081];
assign t[62082] = t[62081] ^ n[62082];
assign t[62083] = t[62082] ^ n[62083];
assign t[62084] = t[62083] ^ n[62084];
assign t[62085] = t[62084] ^ n[62085];
assign t[62086] = t[62085] ^ n[62086];
assign t[62087] = t[62086] ^ n[62087];
assign t[62088] = t[62087] ^ n[62088];
assign t[62089] = t[62088] ^ n[62089];
assign t[62090] = t[62089] ^ n[62090];
assign t[62091] = t[62090] ^ n[62091];
assign t[62092] = t[62091] ^ n[62092];
assign t[62093] = t[62092] ^ n[62093];
assign t[62094] = t[62093] ^ n[62094];
assign t[62095] = t[62094] ^ n[62095];
assign t[62096] = t[62095] ^ n[62096];
assign t[62097] = t[62096] ^ n[62097];
assign t[62098] = t[62097] ^ n[62098];
assign t[62099] = t[62098] ^ n[62099];
assign t[62100] = t[62099] ^ n[62100];
assign t[62101] = t[62100] ^ n[62101];
assign t[62102] = t[62101] ^ n[62102];
assign t[62103] = t[62102] ^ n[62103];
assign t[62104] = t[62103] ^ n[62104];
assign t[62105] = t[62104] ^ n[62105];
assign t[62106] = t[62105] ^ n[62106];
assign t[62107] = t[62106] ^ n[62107];
assign t[62108] = t[62107] ^ n[62108];
assign t[62109] = t[62108] ^ n[62109];
assign t[62110] = t[62109] ^ n[62110];
assign t[62111] = t[62110] ^ n[62111];
assign t[62112] = t[62111] ^ n[62112];
assign t[62113] = t[62112] ^ n[62113];
assign t[62114] = t[62113] ^ n[62114];
assign t[62115] = t[62114] ^ n[62115];
assign t[62116] = t[62115] ^ n[62116];
assign t[62117] = t[62116] ^ n[62117];
assign t[62118] = t[62117] ^ n[62118];
assign t[62119] = t[62118] ^ n[62119];
assign t[62120] = t[62119] ^ n[62120];
assign t[62121] = t[62120] ^ n[62121];
assign t[62122] = t[62121] ^ n[62122];
assign t[62123] = t[62122] ^ n[62123];
assign t[62124] = t[62123] ^ n[62124];
assign t[62125] = t[62124] ^ n[62125];
assign t[62126] = t[62125] ^ n[62126];
assign t[62127] = t[62126] ^ n[62127];
assign t[62128] = t[62127] ^ n[62128];
assign t[62129] = t[62128] ^ n[62129];
assign t[62130] = t[62129] ^ n[62130];
assign t[62131] = t[62130] ^ n[62131];
assign t[62132] = t[62131] ^ n[62132];
assign t[62133] = t[62132] ^ n[62133];
assign t[62134] = t[62133] ^ n[62134];
assign t[62135] = t[62134] ^ n[62135];
assign t[62136] = t[62135] ^ n[62136];
assign t[62137] = t[62136] ^ n[62137];
assign t[62138] = t[62137] ^ n[62138];
assign t[62139] = t[62138] ^ n[62139];
assign t[62140] = t[62139] ^ n[62140];
assign t[62141] = t[62140] ^ n[62141];
assign t[62142] = t[62141] ^ n[62142];
assign t[62143] = t[62142] ^ n[62143];
assign t[62144] = t[62143] ^ n[62144];
assign t[62145] = t[62144] ^ n[62145];
assign t[62146] = t[62145] ^ n[62146];
assign t[62147] = t[62146] ^ n[62147];
assign t[62148] = t[62147] ^ n[62148];
assign t[62149] = t[62148] ^ n[62149];
assign t[62150] = t[62149] ^ n[62150];
assign t[62151] = t[62150] ^ n[62151];
assign t[62152] = t[62151] ^ n[62152];
assign t[62153] = t[62152] ^ n[62153];
assign t[62154] = t[62153] ^ n[62154];
assign t[62155] = t[62154] ^ n[62155];
assign t[62156] = t[62155] ^ n[62156];
assign t[62157] = t[62156] ^ n[62157];
assign t[62158] = t[62157] ^ n[62158];
assign t[62159] = t[62158] ^ n[62159];
assign t[62160] = t[62159] ^ n[62160];
assign t[62161] = t[62160] ^ n[62161];
assign t[62162] = t[62161] ^ n[62162];
assign t[62163] = t[62162] ^ n[62163];
assign t[62164] = t[62163] ^ n[62164];
assign t[62165] = t[62164] ^ n[62165];
assign t[62166] = t[62165] ^ n[62166];
assign t[62167] = t[62166] ^ n[62167];
assign t[62168] = t[62167] ^ n[62168];
assign t[62169] = t[62168] ^ n[62169];
assign t[62170] = t[62169] ^ n[62170];
assign t[62171] = t[62170] ^ n[62171];
assign t[62172] = t[62171] ^ n[62172];
assign t[62173] = t[62172] ^ n[62173];
assign t[62174] = t[62173] ^ n[62174];
assign t[62175] = t[62174] ^ n[62175];
assign t[62176] = t[62175] ^ n[62176];
assign t[62177] = t[62176] ^ n[62177];
assign t[62178] = t[62177] ^ n[62178];
assign t[62179] = t[62178] ^ n[62179];
assign t[62180] = t[62179] ^ n[62180];
assign t[62181] = t[62180] ^ n[62181];
assign t[62182] = t[62181] ^ n[62182];
assign t[62183] = t[62182] ^ n[62183];
assign t[62184] = t[62183] ^ n[62184];
assign t[62185] = t[62184] ^ n[62185];
assign t[62186] = t[62185] ^ n[62186];
assign t[62187] = t[62186] ^ n[62187];
assign t[62188] = t[62187] ^ n[62188];
assign t[62189] = t[62188] ^ n[62189];
assign t[62190] = t[62189] ^ n[62190];
assign t[62191] = t[62190] ^ n[62191];
assign t[62192] = t[62191] ^ n[62192];
assign t[62193] = t[62192] ^ n[62193];
assign t[62194] = t[62193] ^ n[62194];
assign t[62195] = t[62194] ^ n[62195];
assign t[62196] = t[62195] ^ n[62196];
assign t[62197] = t[62196] ^ n[62197];
assign t[62198] = t[62197] ^ n[62198];
assign t[62199] = t[62198] ^ n[62199];
assign t[62200] = t[62199] ^ n[62200];
assign t[62201] = t[62200] ^ n[62201];
assign t[62202] = t[62201] ^ n[62202];
assign t[62203] = t[62202] ^ n[62203];
assign t[62204] = t[62203] ^ n[62204];
assign t[62205] = t[62204] ^ n[62205];
assign t[62206] = t[62205] ^ n[62206];
assign t[62207] = t[62206] ^ n[62207];
assign t[62208] = t[62207] ^ n[62208];
assign t[62209] = t[62208] ^ n[62209];
assign t[62210] = t[62209] ^ n[62210];
assign t[62211] = t[62210] ^ n[62211];
assign t[62212] = t[62211] ^ n[62212];
assign t[62213] = t[62212] ^ n[62213];
assign t[62214] = t[62213] ^ n[62214];
assign t[62215] = t[62214] ^ n[62215];
assign t[62216] = t[62215] ^ n[62216];
assign t[62217] = t[62216] ^ n[62217];
assign t[62218] = t[62217] ^ n[62218];
assign t[62219] = t[62218] ^ n[62219];
assign t[62220] = t[62219] ^ n[62220];
assign t[62221] = t[62220] ^ n[62221];
assign t[62222] = t[62221] ^ n[62222];
assign t[62223] = t[62222] ^ n[62223];
assign t[62224] = t[62223] ^ n[62224];
assign t[62225] = t[62224] ^ n[62225];
assign t[62226] = t[62225] ^ n[62226];
assign t[62227] = t[62226] ^ n[62227];
assign t[62228] = t[62227] ^ n[62228];
assign t[62229] = t[62228] ^ n[62229];
assign t[62230] = t[62229] ^ n[62230];
assign t[62231] = t[62230] ^ n[62231];
assign t[62232] = t[62231] ^ n[62232];
assign t[62233] = t[62232] ^ n[62233];
assign t[62234] = t[62233] ^ n[62234];
assign t[62235] = t[62234] ^ n[62235];
assign t[62236] = t[62235] ^ n[62236];
assign t[62237] = t[62236] ^ n[62237];
assign t[62238] = t[62237] ^ n[62238];
assign t[62239] = t[62238] ^ n[62239];
assign t[62240] = t[62239] ^ n[62240];
assign t[62241] = t[62240] ^ n[62241];
assign t[62242] = t[62241] ^ n[62242];
assign t[62243] = t[62242] ^ n[62243];
assign t[62244] = t[62243] ^ n[62244];
assign t[62245] = t[62244] ^ n[62245];
assign t[62246] = t[62245] ^ n[62246];
assign t[62247] = t[62246] ^ n[62247];
assign t[62248] = t[62247] ^ n[62248];
assign t[62249] = t[62248] ^ n[62249];
assign t[62250] = t[62249] ^ n[62250];
assign t[62251] = t[62250] ^ n[62251];
assign t[62252] = t[62251] ^ n[62252];
assign t[62253] = t[62252] ^ n[62253];
assign t[62254] = t[62253] ^ n[62254];
assign t[62255] = t[62254] ^ n[62255];
assign t[62256] = t[62255] ^ n[62256];
assign t[62257] = t[62256] ^ n[62257];
assign t[62258] = t[62257] ^ n[62258];
assign t[62259] = t[62258] ^ n[62259];
assign t[62260] = t[62259] ^ n[62260];
assign t[62261] = t[62260] ^ n[62261];
assign t[62262] = t[62261] ^ n[62262];
assign t[62263] = t[62262] ^ n[62263];
assign t[62264] = t[62263] ^ n[62264];
assign t[62265] = t[62264] ^ n[62265];
assign t[62266] = t[62265] ^ n[62266];
assign t[62267] = t[62266] ^ n[62267];
assign t[62268] = t[62267] ^ n[62268];
assign t[62269] = t[62268] ^ n[62269];
assign t[62270] = t[62269] ^ n[62270];
assign t[62271] = t[62270] ^ n[62271];
assign t[62272] = t[62271] ^ n[62272];
assign t[62273] = t[62272] ^ n[62273];
assign t[62274] = t[62273] ^ n[62274];
assign t[62275] = t[62274] ^ n[62275];
assign t[62276] = t[62275] ^ n[62276];
assign t[62277] = t[62276] ^ n[62277];
assign t[62278] = t[62277] ^ n[62278];
assign t[62279] = t[62278] ^ n[62279];
assign t[62280] = t[62279] ^ n[62280];
assign t[62281] = t[62280] ^ n[62281];
assign t[62282] = t[62281] ^ n[62282];
assign t[62283] = t[62282] ^ n[62283];
assign t[62284] = t[62283] ^ n[62284];
assign t[62285] = t[62284] ^ n[62285];
assign t[62286] = t[62285] ^ n[62286];
assign t[62287] = t[62286] ^ n[62287];
assign t[62288] = t[62287] ^ n[62288];
assign t[62289] = t[62288] ^ n[62289];
assign t[62290] = t[62289] ^ n[62290];
assign t[62291] = t[62290] ^ n[62291];
assign t[62292] = t[62291] ^ n[62292];
assign t[62293] = t[62292] ^ n[62293];
assign t[62294] = t[62293] ^ n[62294];
assign t[62295] = t[62294] ^ n[62295];
assign t[62296] = t[62295] ^ n[62296];
assign t[62297] = t[62296] ^ n[62297];
assign t[62298] = t[62297] ^ n[62298];
assign t[62299] = t[62298] ^ n[62299];
assign t[62300] = t[62299] ^ n[62300];
assign t[62301] = t[62300] ^ n[62301];
assign t[62302] = t[62301] ^ n[62302];
assign t[62303] = t[62302] ^ n[62303];
assign t[62304] = t[62303] ^ n[62304];
assign t[62305] = t[62304] ^ n[62305];
assign t[62306] = t[62305] ^ n[62306];
assign t[62307] = t[62306] ^ n[62307];
assign t[62308] = t[62307] ^ n[62308];
assign t[62309] = t[62308] ^ n[62309];
assign t[62310] = t[62309] ^ n[62310];
assign t[62311] = t[62310] ^ n[62311];
assign t[62312] = t[62311] ^ n[62312];
assign t[62313] = t[62312] ^ n[62313];
assign t[62314] = t[62313] ^ n[62314];
assign t[62315] = t[62314] ^ n[62315];
assign t[62316] = t[62315] ^ n[62316];
assign t[62317] = t[62316] ^ n[62317];
assign t[62318] = t[62317] ^ n[62318];
assign t[62319] = t[62318] ^ n[62319];
assign t[62320] = t[62319] ^ n[62320];
assign t[62321] = t[62320] ^ n[62321];
assign t[62322] = t[62321] ^ n[62322];
assign t[62323] = t[62322] ^ n[62323];
assign t[62324] = t[62323] ^ n[62324];
assign t[62325] = t[62324] ^ n[62325];
assign t[62326] = t[62325] ^ n[62326];
assign t[62327] = t[62326] ^ n[62327];
assign t[62328] = t[62327] ^ n[62328];
assign t[62329] = t[62328] ^ n[62329];
assign t[62330] = t[62329] ^ n[62330];
assign t[62331] = t[62330] ^ n[62331];
assign t[62332] = t[62331] ^ n[62332];
assign t[62333] = t[62332] ^ n[62333];
assign t[62334] = t[62333] ^ n[62334];
assign t[62335] = t[62334] ^ n[62335];
assign t[62336] = t[62335] ^ n[62336];
assign t[62337] = t[62336] ^ n[62337];
assign t[62338] = t[62337] ^ n[62338];
assign t[62339] = t[62338] ^ n[62339];
assign t[62340] = t[62339] ^ n[62340];
assign t[62341] = t[62340] ^ n[62341];
assign t[62342] = t[62341] ^ n[62342];
assign t[62343] = t[62342] ^ n[62343];
assign t[62344] = t[62343] ^ n[62344];
assign t[62345] = t[62344] ^ n[62345];
assign t[62346] = t[62345] ^ n[62346];
assign t[62347] = t[62346] ^ n[62347];
assign t[62348] = t[62347] ^ n[62348];
assign t[62349] = t[62348] ^ n[62349];
assign t[62350] = t[62349] ^ n[62350];
assign t[62351] = t[62350] ^ n[62351];
assign t[62352] = t[62351] ^ n[62352];
assign t[62353] = t[62352] ^ n[62353];
assign t[62354] = t[62353] ^ n[62354];
assign t[62355] = t[62354] ^ n[62355];
assign t[62356] = t[62355] ^ n[62356];
assign t[62357] = t[62356] ^ n[62357];
assign t[62358] = t[62357] ^ n[62358];
assign t[62359] = t[62358] ^ n[62359];
assign t[62360] = t[62359] ^ n[62360];
assign t[62361] = t[62360] ^ n[62361];
assign t[62362] = t[62361] ^ n[62362];
assign t[62363] = t[62362] ^ n[62363];
assign t[62364] = t[62363] ^ n[62364];
assign t[62365] = t[62364] ^ n[62365];
assign t[62366] = t[62365] ^ n[62366];
assign t[62367] = t[62366] ^ n[62367];
assign t[62368] = t[62367] ^ n[62368];
assign t[62369] = t[62368] ^ n[62369];
assign t[62370] = t[62369] ^ n[62370];
assign t[62371] = t[62370] ^ n[62371];
assign t[62372] = t[62371] ^ n[62372];
assign t[62373] = t[62372] ^ n[62373];
assign t[62374] = t[62373] ^ n[62374];
assign t[62375] = t[62374] ^ n[62375];
assign t[62376] = t[62375] ^ n[62376];
assign t[62377] = t[62376] ^ n[62377];
assign t[62378] = t[62377] ^ n[62378];
assign t[62379] = t[62378] ^ n[62379];
assign t[62380] = t[62379] ^ n[62380];
assign t[62381] = t[62380] ^ n[62381];
assign t[62382] = t[62381] ^ n[62382];
assign t[62383] = t[62382] ^ n[62383];
assign t[62384] = t[62383] ^ n[62384];
assign t[62385] = t[62384] ^ n[62385];
assign t[62386] = t[62385] ^ n[62386];
assign t[62387] = t[62386] ^ n[62387];
assign t[62388] = t[62387] ^ n[62388];
assign t[62389] = t[62388] ^ n[62389];
assign t[62390] = t[62389] ^ n[62390];
assign t[62391] = t[62390] ^ n[62391];
assign t[62392] = t[62391] ^ n[62392];
assign t[62393] = t[62392] ^ n[62393];
assign t[62394] = t[62393] ^ n[62394];
assign t[62395] = t[62394] ^ n[62395];
assign t[62396] = t[62395] ^ n[62396];
assign t[62397] = t[62396] ^ n[62397];
assign t[62398] = t[62397] ^ n[62398];
assign t[62399] = t[62398] ^ n[62399];
assign t[62400] = t[62399] ^ n[62400];
assign t[62401] = t[62400] ^ n[62401];
assign t[62402] = t[62401] ^ n[62402];
assign t[62403] = t[62402] ^ n[62403];
assign t[62404] = t[62403] ^ n[62404];
assign t[62405] = t[62404] ^ n[62405];
assign t[62406] = t[62405] ^ n[62406];
assign t[62407] = t[62406] ^ n[62407];
assign t[62408] = t[62407] ^ n[62408];
assign t[62409] = t[62408] ^ n[62409];
assign t[62410] = t[62409] ^ n[62410];
assign t[62411] = t[62410] ^ n[62411];
assign t[62412] = t[62411] ^ n[62412];
assign t[62413] = t[62412] ^ n[62413];
assign t[62414] = t[62413] ^ n[62414];
assign t[62415] = t[62414] ^ n[62415];
assign t[62416] = t[62415] ^ n[62416];
assign t[62417] = t[62416] ^ n[62417];
assign t[62418] = t[62417] ^ n[62418];
assign t[62419] = t[62418] ^ n[62419];
assign t[62420] = t[62419] ^ n[62420];
assign t[62421] = t[62420] ^ n[62421];
assign t[62422] = t[62421] ^ n[62422];
assign t[62423] = t[62422] ^ n[62423];
assign t[62424] = t[62423] ^ n[62424];
assign t[62425] = t[62424] ^ n[62425];
assign t[62426] = t[62425] ^ n[62426];
assign t[62427] = t[62426] ^ n[62427];
assign t[62428] = t[62427] ^ n[62428];
assign t[62429] = t[62428] ^ n[62429];
assign t[62430] = t[62429] ^ n[62430];
assign t[62431] = t[62430] ^ n[62431];
assign t[62432] = t[62431] ^ n[62432];
assign t[62433] = t[62432] ^ n[62433];
assign t[62434] = t[62433] ^ n[62434];
assign t[62435] = t[62434] ^ n[62435];
assign t[62436] = t[62435] ^ n[62436];
assign t[62437] = t[62436] ^ n[62437];
assign t[62438] = t[62437] ^ n[62438];
assign t[62439] = t[62438] ^ n[62439];
assign t[62440] = t[62439] ^ n[62440];
assign t[62441] = t[62440] ^ n[62441];
assign t[62442] = t[62441] ^ n[62442];
assign t[62443] = t[62442] ^ n[62443];
assign t[62444] = t[62443] ^ n[62444];
assign t[62445] = t[62444] ^ n[62445];
assign t[62446] = t[62445] ^ n[62446];
assign t[62447] = t[62446] ^ n[62447];
assign t[62448] = t[62447] ^ n[62448];
assign t[62449] = t[62448] ^ n[62449];
assign t[62450] = t[62449] ^ n[62450];
assign t[62451] = t[62450] ^ n[62451];
assign t[62452] = t[62451] ^ n[62452];
assign t[62453] = t[62452] ^ n[62453];
assign t[62454] = t[62453] ^ n[62454];
assign t[62455] = t[62454] ^ n[62455];
assign t[62456] = t[62455] ^ n[62456];
assign t[62457] = t[62456] ^ n[62457];
assign t[62458] = t[62457] ^ n[62458];
assign t[62459] = t[62458] ^ n[62459];
assign t[62460] = t[62459] ^ n[62460];
assign t[62461] = t[62460] ^ n[62461];
assign t[62462] = t[62461] ^ n[62462];
assign t[62463] = t[62462] ^ n[62463];
assign t[62464] = t[62463] ^ n[62464];
assign t[62465] = t[62464] ^ n[62465];
assign t[62466] = t[62465] ^ n[62466];
assign t[62467] = t[62466] ^ n[62467];
assign t[62468] = t[62467] ^ n[62468];
assign t[62469] = t[62468] ^ n[62469];
assign t[62470] = t[62469] ^ n[62470];
assign t[62471] = t[62470] ^ n[62471];
assign t[62472] = t[62471] ^ n[62472];
assign t[62473] = t[62472] ^ n[62473];
assign t[62474] = t[62473] ^ n[62474];
assign t[62475] = t[62474] ^ n[62475];
assign t[62476] = t[62475] ^ n[62476];
assign t[62477] = t[62476] ^ n[62477];
assign t[62478] = t[62477] ^ n[62478];
assign t[62479] = t[62478] ^ n[62479];
assign t[62480] = t[62479] ^ n[62480];
assign t[62481] = t[62480] ^ n[62481];
assign t[62482] = t[62481] ^ n[62482];
assign t[62483] = t[62482] ^ n[62483];
assign t[62484] = t[62483] ^ n[62484];
assign t[62485] = t[62484] ^ n[62485];
assign t[62486] = t[62485] ^ n[62486];
assign t[62487] = t[62486] ^ n[62487];
assign t[62488] = t[62487] ^ n[62488];
assign t[62489] = t[62488] ^ n[62489];
assign t[62490] = t[62489] ^ n[62490];
assign t[62491] = t[62490] ^ n[62491];
assign t[62492] = t[62491] ^ n[62492];
assign t[62493] = t[62492] ^ n[62493];
assign t[62494] = t[62493] ^ n[62494];
assign t[62495] = t[62494] ^ n[62495];
assign t[62496] = t[62495] ^ n[62496];
assign t[62497] = t[62496] ^ n[62497];
assign t[62498] = t[62497] ^ n[62498];
assign t[62499] = t[62498] ^ n[62499];
assign t[62500] = t[62499] ^ n[62500];
assign t[62501] = t[62500] ^ n[62501];
assign t[62502] = t[62501] ^ n[62502];
assign t[62503] = t[62502] ^ n[62503];
assign t[62504] = t[62503] ^ n[62504];
assign t[62505] = t[62504] ^ n[62505];
assign t[62506] = t[62505] ^ n[62506];
assign t[62507] = t[62506] ^ n[62507];
assign t[62508] = t[62507] ^ n[62508];
assign t[62509] = t[62508] ^ n[62509];
assign t[62510] = t[62509] ^ n[62510];
assign t[62511] = t[62510] ^ n[62511];
assign t[62512] = t[62511] ^ n[62512];
assign t[62513] = t[62512] ^ n[62513];
assign t[62514] = t[62513] ^ n[62514];
assign t[62515] = t[62514] ^ n[62515];
assign t[62516] = t[62515] ^ n[62516];
assign t[62517] = t[62516] ^ n[62517];
assign t[62518] = t[62517] ^ n[62518];
assign t[62519] = t[62518] ^ n[62519];
assign t[62520] = t[62519] ^ n[62520];
assign t[62521] = t[62520] ^ n[62521];
assign t[62522] = t[62521] ^ n[62522];
assign t[62523] = t[62522] ^ n[62523];
assign t[62524] = t[62523] ^ n[62524];
assign t[62525] = t[62524] ^ n[62525];
assign t[62526] = t[62525] ^ n[62526];
assign t[62527] = t[62526] ^ n[62527];
assign t[62528] = t[62527] ^ n[62528];
assign t[62529] = t[62528] ^ n[62529];
assign t[62530] = t[62529] ^ n[62530];
assign t[62531] = t[62530] ^ n[62531];
assign t[62532] = t[62531] ^ n[62532];
assign t[62533] = t[62532] ^ n[62533];
assign t[62534] = t[62533] ^ n[62534];
assign t[62535] = t[62534] ^ n[62535];
assign t[62536] = t[62535] ^ n[62536];
assign t[62537] = t[62536] ^ n[62537];
assign t[62538] = t[62537] ^ n[62538];
assign t[62539] = t[62538] ^ n[62539];
assign t[62540] = t[62539] ^ n[62540];
assign t[62541] = t[62540] ^ n[62541];
assign t[62542] = t[62541] ^ n[62542];
assign t[62543] = t[62542] ^ n[62543];
assign t[62544] = t[62543] ^ n[62544];
assign t[62545] = t[62544] ^ n[62545];
assign t[62546] = t[62545] ^ n[62546];
assign t[62547] = t[62546] ^ n[62547];
assign t[62548] = t[62547] ^ n[62548];
assign t[62549] = t[62548] ^ n[62549];
assign t[62550] = t[62549] ^ n[62550];
assign t[62551] = t[62550] ^ n[62551];
assign t[62552] = t[62551] ^ n[62552];
assign t[62553] = t[62552] ^ n[62553];
assign t[62554] = t[62553] ^ n[62554];
assign t[62555] = t[62554] ^ n[62555];
assign t[62556] = t[62555] ^ n[62556];
assign t[62557] = t[62556] ^ n[62557];
assign t[62558] = t[62557] ^ n[62558];
assign t[62559] = t[62558] ^ n[62559];
assign t[62560] = t[62559] ^ n[62560];
assign t[62561] = t[62560] ^ n[62561];
assign t[62562] = t[62561] ^ n[62562];
assign t[62563] = t[62562] ^ n[62563];
assign t[62564] = t[62563] ^ n[62564];
assign t[62565] = t[62564] ^ n[62565];
assign t[62566] = t[62565] ^ n[62566];
assign t[62567] = t[62566] ^ n[62567];
assign t[62568] = t[62567] ^ n[62568];
assign t[62569] = t[62568] ^ n[62569];
assign t[62570] = t[62569] ^ n[62570];
assign t[62571] = t[62570] ^ n[62571];
assign t[62572] = t[62571] ^ n[62572];
assign t[62573] = t[62572] ^ n[62573];
assign t[62574] = t[62573] ^ n[62574];
assign t[62575] = t[62574] ^ n[62575];
assign t[62576] = t[62575] ^ n[62576];
assign t[62577] = t[62576] ^ n[62577];
assign t[62578] = t[62577] ^ n[62578];
assign t[62579] = t[62578] ^ n[62579];
assign t[62580] = t[62579] ^ n[62580];
assign t[62581] = t[62580] ^ n[62581];
assign t[62582] = t[62581] ^ n[62582];
assign t[62583] = t[62582] ^ n[62583];
assign t[62584] = t[62583] ^ n[62584];
assign t[62585] = t[62584] ^ n[62585];
assign t[62586] = t[62585] ^ n[62586];
assign t[62587] = t[62586] ^ n[62587];
assign t[62588] = t[62587] ^ n[62588];
assign t[62589] = t[62588] ^ n[62589];
assign t[62590] = t[62589] ^ n[62590];
assign t[62591] = t[62590] ^ n[62591];
assign t[62592] = t[62591] ^ n[62592];
assign t[62593] = t[62592] ^ n[62593];
assign t[62594] = t[62593] ^ n[62594];
assign t[62595] = t[62594] ^ n[62595];
assign t[62596] = t[62595] ^ n[62596];
assign t[62597] = t[62596] ^ n[62597];
assign t[62598] = t[62597] ^ n[62598];
assign t[62599] = t[62598] ^ n[62599];
assign t[62600] = t[62599] ^ n[62600];
assign t[62601] = t[62600] ^ n[62601];
assign t[62602] = t[62601] ^ n[62602];
assign t[62603] = t[62602] ^ n[62603];
assign t[62604] = t[62603] ^ n[62604];
assign t[62605] = t[62604] ^ n[62605];
assign t[62606] = t[62605] ^ n[62606];
assign t[62607] = t[62606] ^ n[62607];
assign t[62608] = t[62607] ^ n[62608];
assign t[62609] = t[62608] ^ n[62609];
assign t[62610] = t[62609] ^ n[62610];
assign t[62611] = t[62610] ^ n[62611];
assign t[62612] = t[62611] ^ n[62612];
assign t[62613] = t[62612] ^ n[62613];
assign t[62614] = t[62613] ^ n[62614];
assign t[62615] = t[62614] ^ n[62615];
assign t[62616] = t[62615] ^ n[62616];
assign t[62617] = t[62616] ^ n[62617];
assign t[62618] = t[62617] ^ n[62618];
assign t[62619] = t[62618] ^ n[62619];
assign t[62620] = t[62619] ^ n[62620];
assign t[62621] = t[62620] ^ n[62621];
assign t[62622] = t[62621] ^ n[62622];
assign t[62623] = t[62622] ^ n[62623];
assign t[62624] = t[62623] ^ n[62624];
assign t[62625] = t[62624] ^ n[62625];
assign t[62626] = t[62625] ^ n[62626];
assign t[62627] = t[62626] ^ n[62627];
assign t[62628] = t[62627] ^ n[62628];
assign t[62629] = t[62628] ^ n[62629];
assign t[62630] = t[62629] ^ n[62630];
assign t[62631] = t[62630] ^ n[62631];
assign t[62632] = t[62631] ^ n[62632];
assign t[62633] = t[62632] ^ n[62633];
assign t[62634] = t[62633] ^ n[62634];
assign t[62635] = t[62634] ^ n[62635];
assign t[62636] = t[62635] ^ n[62636];
assign t[62637] = t[62636] ^ n[62637];
assign t[62638] = t[62637] ^ n[62638];
assign t[62639] = t[62638] ^ n[62639];
assign t[62640] = t[62639] ^ n[62640];
assign t[62641] = t[62640] ^ n[62641];
assign t[62642] = t[62641] ^ n[62642];
assign t[62643] = t[62642] ^ n[62643];
assign t[62644] = t[62643] ^ n[62644];
assign t[62645] = t[62644] ^ n[62645];
assign t[62646] = t[62645] ^ n[62646];
assign t[62647] = t[62646] ^ n[62647];
assign t[62648] = t[62647] ^ n[62648];
assign t[62649] = t[62648] ^ n[62649];
assign t[62650] = t[62649] ^ n[62650];
assign t[62651] = t[62650] ^ n[62651];
assign t[62652] = t[62651] ^ n[62652];
assign t[62653] = t[62652] ^ n[62653];
assign t[62654] = t[62653] ^ n[62654];
assign t[62655] = t[62654] ^ n[62655];
assign t[62656] = t[62655] ^ n[62656];
assign t[62657] = t[62656] ^ n[62657];
assign t[62658] = t[62657] ^ n[62658];
assign t[62659] = t[62658] ^ n[62659];
assign t[62660] = t[62659] ^ n[62660];
assign t[62661] = t[62660] ^ n[62661];
assign t[62662] = t[62661] ^ n[62662];
assign t[62663] = t[62662] ^ n[62663];
assign t[62664] = t[62663] ^ n[62664];
assign t[62665] = t[62664] ^ n[62665];
assign t[62666] = t[62665] ^ n[62666];
assign t[62667] = t[62666] ^ n[62667];
assign t[62668] = t[62667] ^ n[62668];
assign t[62669] = t[62668] ^ n[62669];
assign t[62670] = t[62669] ^ n[62670];
assign t[62671] = t[62670] ^ n[62671];
assign t[62672] = t[62671] ^ n[62672];
assign t[62673] = t[62672] ^ n[62673];
assign t[62674] = t[62673] ^ n[62674];
assign t[62675] = t[62674] ^ n[62675];
assign t[62676] = t[62675] ^ n[62676];
assign t[62677] = t[62676] ^ n[62677];
assign t[62678] = t[62677] ^ n[62678];
assign t[62679] = t[62678] ^ n[62679];
assign t[62680] = t[62679] ^ n[62680];
assign t[62681] = t[62680] ^ n[62681];
assign t[62682] = t[62681] ^ n[62682];
assign t[62683] = t[62682] ^ n[62683];
assign t[62684] = t[62683] ^ n[62684];
assign t[62685] = t[62684] ^ n[62685];
assign t[62686] = t[62685] ^ n[62686];
assign t[62687] = t[62686] ^ n[62687];
assign t[62688] = t[62687] ^ n[62688];
assign t[62689] = t[62688] ^ n[62689];
assign t[62690] = t[62689] ^ n[62690];
assign t[62691] = t[62690] ^ n[62691];
assign t[62692] = t[62691] ^ n[62692];
assign t[62693] = t[62692] ^ n[62693];
assign t[62694] = t[62693] ^ n[62694];
assign t[62695] = t[62694] ^ n[62695];
assign t[62696] = t[62695] ^ n[62696];
assign t[62697] = t[62696] ^ n[62697];
assign t[62698] = t[62697] ^ n[62698];
assign t[62699] = t[62698] ^ n[62699];
assign t[62700] = t[62699] ^ n[62700];
assign t[62701] = t[62700] ^ n[62701];
assign t[62702] = t[62701] ^ n[62702];
assign t[62703] = t[62702] ^ n[62703];
assign t[62704] = t[62703] ^ n[62704];
assign t[62705] = t[62704] ^ n[62705];
assign t[62706] = t[62705] ^ n[62706];
assign t[62707] = t[62706] ^ n[62707];
assign t[62708] = t[62707] ^ n[62708];
assign t[62709] = t[62708] ^ n[62709];
assign t[62710] = t[62709] ^ n[62710];
assign t[62711] = t[62710] ^ n[62711];
assign t[62712] = t[62711] ^ n[62712];
assign t[62713] = t[62712] ^ n[62713];
assign t[62714] = t[62713] ^ n[62714];
assign t[62715] = t[62714] ^ n[62715];
assign t[62716] = t[62715] ^ n[62716];
assign t[62717] = t[62716] ^ n[62717];
assign t[62718] = t[62717] ^ n[62718];
assign t[62719] = t[62718] ^ n[62719];
assign t[62720] = t[62719] ^ n[62720];
assign t[62721] = t[62720] ^ n[62721];
assign t[62722] = t[62721] ^ n[62722];
assign t[62723] = t[62722] ^ n[62723];
assign t[62724] = t[62723] ^ n[62724];
assign t[62725] = t[62724] ^ n[62725];
assign t[62726] = t[62725] ^ n[62726];
assign t[62727] = t[62726] ^ n[62727];
assign t[62728] = t[62727] ^ n[62728];
assign t[62729] = t[62728] ^ n[62729];
assign t[62730] = t[62729] ^ n[62730];
assign t[62731] = t[62730] ^ n[62731];
assign t[62732] = t[62731] ^ n[62732];
assign t[62733] = t[62732] ^ n[62733];
assign t[62734] = t[62733] ^ n[62734];
assign t[62735] = t[62734] ^ n[62735];
assign t[62736] = t[62735] ^ n[62736];
assign t[62737] = t[62736] ^ n[62737];
assign t[62738] = t[62737] ^ n[62738];
assign t[62739] = t[62738] ^ n[62739];
assign t[62740] = t[62739] ^ n[62740];
assign t[62741] = t[62740] ^ n[62741];
assign t[62742] = t[62741] ^ n[62742];
assign t[62743] = t[62742] ^ n[62743];
assign t[62744] = t[62743] ^ n[62744];
assign t[62745] = t[62744] ^ n[62745];
assign t[62746] = t[62745] ^ n[62746];
assign t[62747] = t[62746] ^ n[62747];
assign t[62748] = t[62747] ^ n[62748];
assign t[62749] = t[62748] ^ n[62749];
assign t[62750] = t[62749] ^ n[62750];
assign t[62751] = t[62750] ^ n[62751];
assign t[62752] = t[62751] ^ n[62752];
assign t[62753] = t[62752] ^ n[62753];
assign t[62754] = t[62753] ^ n[62754];
assign t[62755] = t[62754] ^ n[62755];
assign t[62756] = t[62755] ^ n[62756];
assign t[62757] = t[62756] ^ n[62757];
assign t[62758] = t[62757] ^ n[62758];
assign t[62759] = t[62758] ^ n[62759];
assign t[62760] = t[62759] ^ n[62760];
assign t[62761] = t[62760] ^ n[62761];
assign t[62762] = t[62761] ^ n[62762];
assign t[62763] = t[62762] ^ n[62763];
assign t[62764] = t[62763] ^ n[62764];
assign t[62765] = t[62764] ^ n[62765];
assign t[62766] = t[62765] ^ n[62766];
assign t[62767] = t[62766] ^ n[62767];
assign t[62768] = t[62767] ^ n[62768];
assign t[62769] = t[62768] ^ n[62769];
assign t[62770] = t[62769] ^ n[62770];
assign t[62771] = t[62770] ^ n[62771];
assign t[62772] = t[62771] ^ n[62772];
assign t[62773] = t[62772] ^ n[62773];
assign t[62774] = t[62773] ^ n[62774];
assign t[62775] = t[62774] ^ n[62775];
assign t[62776] = t[62775] ^ n[62776];
assign t[62777] = t[62776] ^ n[62777];
assign t[62778] = t[62777] ^ n[62778];
assign t[62779] = t[62778] ^ n[62779];
assign t[62780] = t[62779] ^ n[62780];
assign t[62781] = t[62780] ^ n[62781];
assign t[62782] = t[62781] ^ n[62782];
assign t[62783] = t[62782] ^ n[62783];
assign t[62784] = t[62783] ^ n[62784];
assign t[62785] = t[62784] ^ n[62785];
assign t[62786] = t[62785] ^ n[62786];
assign t[62787] = t[62786] ^ n[62787];
assign t[62788] = t[62787] ^ n[62788];
assign t[62789] = t[62788] ^ n[62789];
assign t[62790] = t[62789] ^ n[62790];
assign t[62791] = t[62790] ^ n[62791];
assign t[62792] = t[62791] ^ n[62792];
assign t[62793] = t[62792] ^ n[62793];
assign t[62794] = t[62793] ^ n[62794];
assign t[62795] = t[62794] ^ n[62795];
assign t[62796] = t[62795] ^ n[62796];
assign t[62797] = t[62796] ^ n[62797];
assign t[62798] = t[62797] ^ n[62798];
assign t[62799] = t[62798] ^ n[62799];
assign t[62800] = t[62799] ^ n[62800];
assign t[62801] = t[62800] ^ n[62801];
assign t[62802] = t[62801] ^ n[62802];
assign t[62803] = t[62802] ^ n[62803];
assign t[62804] = t[62803] ^ n[62804];
assign t[62805] = t[62804] ^ n[62805];
assign t[62806] = t[62805] ^ n[62806];
assign t[62807] = t[62806] ^ n[62807];
assign t[62808] = t[62807] ^ n[62808];
assign t[62809] = t[62808] ^ n[62809];
assign t[62810] = t[62809] ^ n[62810];
assign t[62811] = t[62810] ^ n[62811];
assign t[62812] = t[62811] ^ n[62812];
assign t[62813] = t[62812] ^ n[62813];
assign t[62814] = t[62813] ^ n[62814];
assign t[62815] = t[62814] ^ n[62815];
assign t[62816] = t[62815] ^ n[62816];
assign t[62817] = t[62816] ^ n[62817];
assign t[62818] = t[62817] ^ n[62818];
assign t[62819] = t[62818] ^ n[62819];
assign t[62820] = t[62819] ^ n[62820];
assign t[62821] = t[62820] ^ n[62821];
assign t[62822] = t[62821] ^ n[62822];
assign t[62823] = t[62822] ^ n[62823];
assign t[62824] = t[62823] ^ n[62824];
assign t[62825] = t[62824] ^ n[62825];
assign t[62826] = t[62825] ^ n[62826];
assign t[62827] = t[62826] ^ n[62827];
assign t[62828] = t[62827] ^ n[62828];
assign t[62829] = t[62828] ^ n[62829];
assign t[62830] = t[62829] ^ n[62830];
assign t[62831] = t[62830] ^ n[62831];
assign t[62832] = t[62831] ^ n[62832];
assign t[62833] = t[62832] ^ n[62833];
assign t[62834] = t[62833] ^ n[62834];
assign t[62835] = t[62834] ^ n[62835];
assign t[62836] = t[62835] ^ n[62836];
assign t[62837] = t[62836] ^ n[62837];
assign t[62838] = t[62837] ^ n[62838];
assign t[62839] = t[62838] ^ n[62839];
assign t[62840] = t[62839] ^ n[62840];
assign t[62841] = t[62840] ^ n[62841];
assign t[62842] = t[62841] ^ n[62842];
assign t[62843] = t[62842] ^ n[62843];
assign t[62844] = t[62843] ^ n[62844];
assign t[62845] = t[62844] ^ n[62845];
assign t[62846] = t[62845] ^ n[62846];
assign t[62847] = t[62846] ^ n[62847];
assign t[62848] = t[62847] ^ n[62848];
assign t[62849] = t[62848] ^ n[62849];
assign t[62850] = t[62849] ^ n[62850];
assign t[62851] = t[62850] ^ n[62851];
assign t[62852] = t[62851] ^ n[62852];
assign t[62853] = t[62852] ^ n[62853];
assign t[62854] = t[62853] ^ n[62854];
assign t[62855] = t[62854] ^ n[62855];
assign t[62856] = t[62855] ^ n[62856];
assign t[62857] = t[62856] ^ n[62857];
assign t[62858] = t[62857] ^ n[62858];
assign t[62859] = t[62858] ^ n[62859];
assign t[62860] = t[62859] ^ n[62860];
assign t[62861] = t[62860] ^ n[62861];
assign t[62862] = t[62861] ^ n[62862];
assign t[62863] = t[62862] ^ n[62863];
assign t[62864] = t[62863] ^ n[62864];
assign t[62865] = t[62864] ^ n[62865];
assign t[62866] = t[62865] ^ n[62866];
assign t[62867] = t[62866] ^ n[62867];
assign t[62868] = t[62867] ^ n[62868];
assign t[62869] = t[62868] ^ n[62869];
assign t[62870] = t[62869] ^ n[62870];
assign t[62871] = t[62870] ^ n[62871];
assign t[62872] = t[62871] ^ n[62872];
assign t[62873] = t[62872] ^ n[62873];
assign t[62874] = t[62873] ^ n[62874];
assign t[62875] = t[62874] ^ n[62875];
assign t[62876] = t[62875] ^ n[62876];
assign t[62877] = t[62876] ^ n[62877];
assign t[62878] = t[62877] ^ n[62878];
assign t[62879] = t[62878] ^ n[62879];
assign t[62880] = t[62879] ^ n[62880];
assign t[62881] = t[62880] ^ n[62881];
assign t[62882] = t[62881] ^ n[62882];
assign t[62883] = t[62882] ^ n[62883];
assign t[62884] = t[62883] ^ n[62884];
assign t[62885] = t[62884] ^ n[62885];
assign t[62886] = t[62885] ^ n[62886];
assign t[62887] = t[62886] ^ n[62887];
assign t[62888] = t[62887] ^ n[62888];
assign t[62889] = t[62888] ^ n[62889];
assign t[62890] = t[62889] ^ n[62890];
assign t[62891] = t[62890] ^ n[62891];
assign t[62892] = t[62891] ^ n[62892];
assign t[62893] = t[62892] ^ n[62893];
assign t[62894] = t[62893] ^ n[62894];
assign t[62895] = t[62894] ^ n[62895];
assign t[62896] = t[62895] ^ n[62896];
assign t[62897] = t[62896] ^ n[62897];
assign t[62898] = t[62897] ^ n[62898];
assign t[62899] = t[62898] ^ n[62899];
assign t[62900] = t[62899] ^ n[62900];
assign t[62901] = t[62900] ^ n[62901];
assign t[62902] = t[62901] ^ n[62902];
assign t[62903] = t[62902] ^ n[62903];
assign t[62904] = t[62903] ^ n[62904];
assign t[62905] = t[62904] ^ n[62905];
assign t[62906] = t[62905] ^ n[62906];
assign t[62907] = t[62906] ^ n[62907];
assign t[62908] = t[62907] ^ n[62908];
assign t[62909] = t[62908] ^ n[62909];
assign t[62910] = t[62909] ^ n[62910];
assign t[62911] = t[62910] ^ n[62911];
assign t[62912] = t[62911] ^ n[62912];
assign t[62913] = t[62912] ^ n[62913];
assign t[62914] = t[62913] ^ n[62914];
assign t[62915] = t[62914] ^ n[62915];
assign t[62916] = t[62915] ^ n[62916];
assign t[62917] = t[62916] ^ n[62917];
assign t[62918] = t[62917] ^ n[62918];
assign t[62919] = t[62918] ^ n[62919];
assign t[62920] = t[62919] ^ n[62920];
assign t[62921] = t[62920] ^ n[62921];
assign t[62922] = t[62921] ^ n[62922];
assign t[62923] = t[62922] ^ n[62923];
assign t[62924] = t[62923] ^ n[62924];
assign t[62925] = t[62924] ^ n[62925];
assign t[62926] = t[62925] ^ n[62926];
assign t[62927] = t[62926] ^ n[62927];
assign t[62928] = t[62927] ^ n[62928];
assign t[62929] = t[62928] ^ n[62929];
assign t[62930] = t[62929] ^ n[62930];
assign t[62931] = t[62930] ^ n[62931];
assign t[62932] = t[62931] ^ n[62932];
assign t[62933] = t[62932] ^ n[62933];
assign t[62934] = t[62933] ^ n[62934];
assign t[62935] = t[62934] ^ n[62935];
assign t[62936] = t[62935] ^ n[62936];
assign t[62937] = t[62936] ^ n[62937];
assign t[62938] = t[62937] ^ n[62938];
assign t[62939] = t[62938] ^ n[62939];
assign t[62940] = t[62939] ^ n[62940];
assign t[62941] = t[62940] ^ n[62941];
assign t[62942] = t[62941] ^ n[62942];
assign t[62943] = t[62942] ^ n[62943];
assign t[62944] = t[62943] ^ n[62944];
assign t[62945] = t[62944] ^ n[62945];
assign t[62946] = t[62945] ^ n[62946];
assign t[62947] = t[62946] ^ n[62947];
assign t[62948] = t[62947] ^ n[62948];
assign t[62949] = t[62948] ^ n[62949];
assign t[62950] = t[62949] ^ n[62950];
assign t[62951] = t[62950] ^ n[62951];
assign t[62952] = t[62951] ^ n[62952];
assign t[62953] = t[62952] ^ n[62953];
assign t[62954] = t[62953] ^ n[62954];
assign t[62955] = t[62954] ^ n[62955];
assign t[62956] = t[62955] ^ n[62956];
assign t[62957] = t[62956] ^ n[62957];
assign t[62958] = t[62957] ^ n[62958];
assign t[62959] = t[62958] ^ n[62959];
assign t[62960] = t[62959] ^ n[62960];
assign t[62961] = t[62960] ^ n[62961];
assign t[62962] = t[62961] ^ n[62962];
assign t[62963] = t[62962] ^ n[62963];
assign t[62964] = t[62963] ^ n[62964];
assign t[62965] = t[62964] ^ n[62965];
assign t[62966] = t[62965] ^ n[62966];
assign t[62967] = t[62966] ^ n[62967];
assign t[62968] = t[62967] ^ n[62968];
assign t[62969] = t[62968] ^ n[62969];
assign t[62970] = t[62969] ^ n[62970];
assign t[62971] = t[62970] ^ n[62971];
assign t[62972] = t[62971] ^ n[62972];
assign t[62973] = t[62972] ^ n[62973];
assign t[62974] = t[62973] ^ n[62974];
assign t[62975] = t[62974] ^ n[62975];
assign t[62976] = t[62975] ^ n[62976];
assign t[62977] = t[62976] ^ n[62977];
assign t[62978] = t[62977] ^ n[62978];
assign t[62979] = t[62978] ^ n[62979];
assign t[62980] = t[62979] ^ n[62980];
assign t[62981] = t[62980] ^ n[62981];
assign t[62982] = t[62981] ^ n[62982];
assign t[62983] = t[62982] ^ n[62983];
assign t[62984] = t[62983] ^ n[62984];
assign t[62985] = t[62984] ^ n[62985];
assign t[62986] = t[62985] ^ n[62986];
assign t[62987] = t[62986] ^ n[62987];
assign t[62988] = t[62987] ^ n[62988];
assign t[62989] = t[62988] ^ n[62989];
assign t[62990] = t[62989] ^ n[62990];
assign t[62991] = t[62990] ^ n[62991];
assign t[62992] = t[62991] ^ n[62992];
assign t[62993] = t[62992] ^ n[62993];
assign t[62994] = t[62993] ^ n[62994];
assign t[62995] = t[62994] ^ n[62995];
assign t[62996] = t[62995] ^ n[62996];
assign t[62997] = t[62996] ^ n[62997];
assign t[62998] = t[62997] ^ n[62998];
assign t[62999] = t[62998] ^ n[62999];
assign t[63000] = t[62999] ^ n[63000];
assign t[63001] = t[63000] ^ n[63001];
assign t[63002] = t[63001] ^ n[63002];
assign t[63003] = t[63002] ^ n[63003];
assign t[63004] = t[63003] ^ n[63004];
assign t[63005] = t[63004] ^ n[63005];
assign t[63006] = t[63005] ^ n[63006];
assign t[63007] = t[63006] ^ n[63007];
assign t[63008] = t[63007] ^ n[63008];
assign t[63009] = t[63008] ^ n[63009];
assign t[63010] = t[63009] ^ n[63010];
assign t[63011] = t[63010] ^ n[63011];
assign t[63012] = t[63011] ^ n[63012];
assign t[63013] = t[63012] ^ n[63013];
assign t[63014] = t[63013] ^ n[63014];
assign t[63015] = t[63014] ^ n[63015];
assign t[63016] = t[63015] ^ n[63016];
assign t[63017] = t[63016] ^ n[63017];
assign t[63018] = t[63017] ^ n[63018];
assign t[63019] = t[63018] ^ n[63019];
assign t[63020] = t[63019] ^ n[63020];
assign t[63021] = t[63020] ^ n[63021];
assign t[63022] = t[63021] ^ n[63022];
assign t[63023] = t[63022] ^ n[63023];
assign t[63024] = t[63023] ^ n[63024];
assign t[63025] = t[63024] ^ n[63025];
assign t[63026] = t[63025] ^ n[63026];
assign t[63027] = t[63026] ^ n[63027];
assign t[63028] = t[63027] ^ n[63028];
assign t[63029] = t[63028] ^ n[63029];
assign t[63030] = t[63029] ^ n[63030];
assign t[63031] = t[63030] ^ n[63031];
assign t[63032] = t[63031] ^ n[63032];
assign t[63033] = t[63032] ^ n[63033];
assign t[63034] = t[63033] ^ n[63034];
assign t[63035] = t[63034] ^ n[63035];
assign t[63036] = t[63035] ^ n[63036];
assign t[63037] = t[63036] ^ n[63037];
assign t[63038] = t[63037] ^ n[63038];
assign t[63039] = t[63038] ^ n[63039];
assign t[63040] = t[63039] ^ n[63040];
assign t[63041] = t[63040] ^ n[63041];
assign t[63042] = t[63041] ^ n[63042];
assign t[63043] = t[63042] ^ n[63043];
assign t[63044] = t[63043] ^ n[63044];
assign t[63045] = t[63044] ^ n[63045];
assign t[63046] = t[63045] ^ n[63046];
assign t[63047] = t[63046] ^ n[63047];
assign t[63048] = t[63047] ^ n[63048];
assign t[63049] = t[63048] ^ n[63049];
assign t[63050] = t[63049] ^ n[63050];
assign t[63051] = t[63050] ^ n[63051];
assign t[63052] = t[63051] ^ n[63052];
assign t[63053] = t[63052] ^ n[63053];
assign t[63054] = t[63053] ^ n[63054];
assign t[63055] = t[63054] ^ n[63055];
assign t[63056] = t[63055] ^ n[63056];
assign t[63057] = t[63056] ^ n[63057];
assign t[63058] = t[63057] ^ n[63058];
assign t[63059] = t[63058] ^ n[63059];
assign t[63060] = t[63059] ^ n[63060];
assign t[63061] = t[63060] ^ n[63061];
assign t[63062] = t[63061] ^ n[63062];
assign t[63063] = t[63062] ^ n[63063];
assign t[63064] = t[63063] ^ n[63064];
assign t[63065] = t[63064] ^ n[63065];
assign t[63066] = t[63065] ^ n[63066];
assign t[63067] = t[63066] ^ n[63067];
assign t[63068] = t[63067] ^ n[63068];
assign t[63069] = t[63068] ^ n[63069];
assign t[63070] = t[63069] ^ n[63070];
assign t[63071] = t[63070] ^ n[63071];
assign t[63072] = t[63071] ^ n[63072];
assign t[63073] = t[63072] ^ n[63073];
assign t[63074] = t[63073] ^ n[63074];
assign t[63075] = t[63074] ^ n[63075];
assign t[63076] = t[63075] ^ n[63076];
assign t[63077] = t[63076] ^ n[63077];
assign t[63078] = t[63077] ^ n[63078];
assign t[63079] = t[63078] ^ n[63079];
assign t[63080] = t[63079] ^ n[63080];
assign t[63081] = t[63080] ^ n[63081];
assign t[63082] = t[63081] ^ n[63082];
assign t[63083] = t[63082] ^ n[63083];
assign t[63084] = t[63083] ^ n[63084];
assign t[63085] = t[63084] ^ n[63085];
assign t[63086] = t[63085] ^ n[63086];
assign t[63087] = t[63086] ^ n[63087];
assign t[63088] = t[63087] ^ n[63088];
assign t[63089] = t[63088] ^ n[63089];
assign t[63090] = t[63089] ^ n[63090];
assign t[63091] = t[63090] ^ n[63091];
assign t[63092] = t[63091] ^ n[63092];
assign t[63093] = t[63092] ^ n[63093];
assign t[63094] = t[63093] ^ n[63094];
assign t[63095] = t[63094] ^ n[63095];
assign t[63096] = t[63095] ^ n[63096];
assign t[63097] = t[63096] ^ n[63097];
assign t[63098] = t[63097] ^ n[63098];
assign t[63099] = t[63098] ^ n[63099];
assign t[63100] = t[63099] ^ n[63100];
assign t[63101] = t[63100] ^ n[63101];
assign t[63102] = t[63101] ^ n[63102];
assign t[63103] = t[63102] ^ n[63103];
assign t[63104] = t[63103] ^ n[63104];
assign t[63105] = t[63104] ^ n[63105];
assign t[63106] = t[63105] ^ n[63106];
assign t[63107] = t[63106] ^ n[63107];
assign t[63108] = t[63107] ^ n[63108];
assign t[63109] = t[63108] ^ n[63109];
assign t[63110] = t[63109] ^ n[63110];
assign t[63111] = t[63110] ^ n[63111];
assign t[63112] = t[63111] ^ n[63112];
assign t[63113] = t[63112] ^ n[63113];
assign t[63114] = t[63113] ^ n[63114];
assign t[63115] = t[63114] ^ n[63115];
assign t[63116] = t[63115] ^ n[63116];
assign t[63117] = t[63116] ^ n[63117];
assign t[63118] = t[63117] ^ n[63118];
assign t[63119] = t[63118] ^ n[63119];
assign t[63120] = t[63119] ^ n[63120];
assign t[63121] = t[63120] ^ n[63121];
assign t[63122] = t[63121] ^ n[63122];
assign t[63123] = t[63122] ^ n[63123];
assign t[63124] = t[63123] ^ n[63124];
assign t[63125] = t[63124] ^ n[63125];
assign t[63126] = t[63125] ^ n[63126];
assign t[63127] = t[63126] ^ n[63127];
assign t[63128] = t[63127] ^ n[63128];
assign t[63129] = t[63128] ^ n[63129];
assign t[63130] = t[63129] ^ n[63130];
assign t[63131] = t[63130] ^ n[63131];
assign t[63132] = t[63131] ^ n[63132];
assign t[63133] = t[63132] ^ n[63133];
assign t[63134] = t[63133] ^ n[63134];
assign t[63135] = t[63134] ^ n[63135];
assign t[63136] = t[63135] ^ n[63136];
assign t[63137] = t[63136] ^ n[63137];
assign t[63138] = t[63137] ^ n[63138];
assign t[63139] = t[63138] ^ n[63139];
assign t[63140] = t[63139] ^ n[63140];
assign t[63141] = t[63140] ^ n[63141];
assign t[63142] = t[63141] ^ n[63142];
assign t[63143] = t[63142] ^ n[63143];
assign t[63144] = t[63143] ^ n[63144];
assign t[63145] = t[63144] ^ n[63145];
assign t[63146] = t[63145] ^ n[63146];
assign t[63147] = t[63146] ^ n[63147];
assign t[63148] = t[63147] ^ n[63148];
assign t[63149] = t[63148] ^ n[63149];
assign t[63150] = t[63149] ^ n[63150];
assign t[63151] = t[63150] ^ n[63151];
assign t[63152] = t[63151] ^ n[63152];
assign t[63153] = t[63152] ^ n[63153];
assign t[63154] = t[63153] ^ n[63154];
assign t[63155] = t[63154] ^ n[63155];
assign t[63156] = t[63155] ^ n[63156];
assign t[63157] = t[63156] ^ n[63157];
assign t[63158] = t[63157] ^ n[63158];
assign t[63159] = t[63158] ^ n[63159];
assign t[63160] = t[63159] ^ n[63160];
assign t[63161] = t[63160] ^ n[63161];
assign t[63162] = t[63161] ^ n[63162];
assign t[63163] = t[63162] ^ n[63163];
assign t[63164] = t[63163] ^ n[63164];
assign t[63165] = t[63164] ^ n[63165];
assign t[63166] = t[63165] ^ n[63166];
assign t[63167] = t[63166] ^ n[63167];
assign t[63168] = t[63167] ^ n[63168];
assign t[63169] = t[63168] ^ n[63169];
assign t[63170] = t[63169] ^ n[63170];
assign t[63171] = t[63170] ^ n[63171];
assign t[63172] = t[63171] ^ n[63172];
assign t[63173] = t[63172] ^ n[63173];
assign t[63174] = t[63173] ^ n[63174];
assign t[63175] = t[63174] ^ n[63175];
assign t[63176] = t[63175] ^ n[63176];
assign t[63177] = t[63176] ^ n[63177];
assign t[63178] = t[63177] ^ n[63178];
assign t[63179] = t[63178] ^ n[63179];
assign t[63180] = t[63179] ^ n[63180];
assign t[63181] = t[63180] ^ n[63181];
assign t[63182] = t[63181] ^ n[63182];
assign t[63183] = t[63182] ^ n[63183];
assign t[63184] = t[63183] ^ n[63184];
assign t[63185] = t[63184] ^ n[63185];
assign t[63186] = t[63185] ^ n[63186];
assign t[63187] = t[63186] ^ n[63187];
assign t[63188] = t[63187] ^ n[63188];
assign t[63189] = t[63188] ^ n[63189];
assign t[63190] = t[63189] ^ n[63190];
assign t[63191] = t[63190] ^ n[63191];
assign t[63192] = t[63191] ^ n[63192];
assign t[63193] = t[63192] ^ n[63193];
assign t[63194] = t[63193] ^ n[63194];
assign t[63195] = t[63194] ^ n[63195];
assign t[63196] = t[63195] ^ n[63196];
assign t[63197] = t[63196] ^ n[63197];
assign t[63198] = t[63197] ^ n[63198];
assign t[63199] = t[63198] ^ n[63199];
assign t[63200] = t[63199] ^ n[63200];
assign t[63201] = t[63200] ^ n[63201];
assign t[63202] = t[63201] ^ n[63202];
assign t[63203] = t[63202] ^ n[63203];
assign t[63204] = t[63203] ^ n[63204];
assign t[63205] = t[63204] ^ n[63205];
assign t[63206] = t[63205] ^ n[63206];
assign t[63207] = t[63206] ^ n[63207];
assign t[63208] = t[63207] ^ n[63208];
assign t[63209] = t[63208] ^ n[63209];
assign t[63210] = t[63209] ^ n[63210];
assign t[63211] = t[63210] ^ n[63211];
assign t[63212] = t[63211] ^ n[63212];
assign t[63213] = t[63212] ^ n[63213];
assign t[63214] = t[63213] ^ n[63214];
assign t[63215] = t[63214] ^ n[63215];
assign t[63216] = t[63215] ^ n[63216];
assign t[63217] = t[63216] ^ n[63217];
assign t[63218] = t[63217] ^ n[63218];
assign t[63219] = t[63218] ^ n[63219];
assign t[63220] = t[63219] ^ n[63220];
assign t[63221] = t[63220] ^ n[63221];
assign t[63222] = t[63221] ^ n[63222];
assign t[63223] = t[63222] ^ n[63223];
assign t[63224] = t[63223] ^ n[63224];
assign t[63225] = t[63224] ^ n[63225];
assign t[63226] = t[63225] ^ n[63226];
assign t[63227] = t[63226] ^ n[63227];
assign t[63228] = t[63227] ^ n[63228];
assign t[63229] = t[63228] ^ n[63229];
assign t[63230] = t[63229] ^ n[63230];
assign t[63231] = t[63230] ^ n[63231];
assign t[63232] = t[63231] ^ n[63232];
assign t[63233] = t[63232] ^ n[63233];
assign t[63234] = t[63233] ^ n[63234];
assign t[63235] = t[63234] ^ n[63235];
assign t[63236] = t[63235] ^ n[63236];
assign t[63237] = t[63236] ^ n[63237];
assign t[63238] = t[63237] ^ n[63238];
assign t[63239] = t[63238] ^ n[63239];
assign t[63240] = t[63239] ^ n[63240];
assign t[63241] = t[63240] ^ n[63241];
assign t[63242] = t[63241] ^ n[63242];
assign t[63243] = t[63242] ^ n[63243];
assign t[63244] = t[63243] ^ n[63244];
assign t[63245] = t[63244] ^ n[63245];
assign t[63246] = t[63245] ^ n[63246];
assign t[63247] = t[63246] ^ n[63247];
assign t[63248] = t[63247] ^ n[63248];
assign t[63249] = t[63248] ^ n[63249];
assign t[63250] = t[63249] ^ n[63250];
assign t[63251] = t[63250] ^ n[63251];
assign t[63252] = t[63251] ^ n[63252];
assign t[63253] = t[63252] ^ n[63253];
assign t[63254] = t[63253] ^ n[63254];
assign t[63255] = t[63254] ^ n[63255];
assign t[63256] = t[63255] ^ n[63256];
assign t[63257] = t[63256] ^ n[63257];
assign t[63258] = t[63257] ^ n[63258];
assign t[63259] = t[63258] ^ n[63259];
assign t[63260] = t[63259] ^ n[63260];
assign t[63261] = t[63260] ^ n[63261];
assign t[63262] = t[63261] ^ n[63262];
assign t[63263] = t[63262] ^ n[63263];
assign t[63264] = t[63263] ^ n[63264];
assign t[63265] = t[63264] ^ n[63265];
assign t[63266] = t[63265] ^ n[63266];
assign t[63267] = t[63266] ^ n[63267];
assign t[63268] = t[63267] ^ n[63268];
assign t[63269] = t[63268] ^ n[63269];
assign t[63270] = t[63269] ^ n[63270];
assign t[63271] = t[63270] ^ n[63271];
assign t[63272] = t[63271] ^ n[63272];
assign t[63273] = t[63272] ^ n[63273];
assign t[63274] = t[63273] ^ n[63274];
assign t[63275] = t[63274] ^ n[63275];
assign t[63276] = t[63275] ^ n[63276];
assign t[63277] = t[63276] ^ n[63277];
assign t[63278] = t[63277] ^ n[63278];
assign t[63279] = t[63278] ^ n[63279];
assign t[63280] = t[63279] ^ n[63280];
assign t[63281] = t[63280] ^ n[63281];
assign t[63282] = t[63281] ^ n[63282];
assign t[63283] = t[63282] ^ n[63283];
assign t[63284] = t[63283] ^ n[63284];
assign t[63285] = t[63284] ^ n[63285];
assign t[63286] = t[63285] ^ n[63286];
assign t[63287] = t[63286] ^ n[63287];
assign t[63288] = t[63287] ^ n[63288];
assign t[63289] = t[63288] ^ n[63289];
assign t[63290] = t[63289] ^ n[63290];
assign t[63291] = t[63290] ^ n[63291];
assign t[63292] = t[63291] ^ n[63292];
assign t[63293] = t[63292] ^ n[63293];
assign t[63294] = t[63293] ^ n[63294];
assign t[63295] = t[63294] ^ n[63295];
assign t[63296] = t[63295] ^ n[63296];
assign t[63297] = t[63296] ^ n[63297];
assign t[63298] = t[63297] ^ n[63298];
assign t[63299] = t[63298] ^ n[63299];
assign t[63300] = t[63299] ^ n[63300];
assign t[63301] = t[63300] ^ n[63301];
assign t[63302] = t[63301] ^ n[63302];
assign t[63303] = t[63302] ^ n[63303];
assign t[63304] = t[63303] ^ n[63304];
assign t[63305] = t[63304] ^ n[63305];
assign t[63306] = t[63305] ^ n[63306];
assign t[63307] = t[63306] ^ n[63307];
assign t[63308] = t[63307] ^ n[63308];
assign t[63309] = t[63308] ^ n[63309];
assign t[63310] = t[63309] ^ n[63310];
assign t[63311] = t[63310] ^ n[63311];
assign t[63312] = t[63311] ^ n[63312];
assign t[63313] = t[63312] ^ n[63313];
assign t[63314] = t[63313] ^ n[63314];
assign t[63315] = t[63314] ^ n[63315];
assign t[63316] = t[63315] ^ n[63316];
assign t[63317] = t[63316] ^ n[63317];
assign t[63318] = t[63317] ^ n[63318];
assign t[63319] = t[63318] ^ n[63319];
assign t[63320] = t[63319] ^ n[63320];
assign t[63321] = t[63320] ^ n[63321];
assign t[63322] = t[63321] ^ n[63322];
assign t[63323] = t[63322] ^ n[63323];
assign t[63324] = t[63323] ^ n[63324];
assign t[63325] = t[63324] ^ n[63325];
assign t[63326] = t[63325] ^ n[63326];
assign t[63327] = t[63326] ^ n[63327];
assign t[63328] = t[63327] ^ n[63328];
assign t[63329] = t[63328] ^ n[63329];
assign t[63330] = t[63329] ^ n[63330];
assign t[63331] = t[63330] ^ n[63331];
assign t[63332] = t[63331] ^ n[63332];
assign t[63333] = t[63332] ^ n[63333];
assign t[63334] = t[63333] ^ n[63334];
assign t[63335] = t[63334] ^ n[63335];
assign t[63336] = t[63335] ^ n[63336];
assign t[63337] = t[63336] ^ n[63337];
assign t[63338] = t[63337] ^ n[63338];
assign t[63339] = t[63338] ^ n[63339];
assign t[63340] = t[63339] ^ n[63340];
assign t[63341] = t[63340] ^ n[63341];
assign t[63342] = t[63341] ^ n[63342];
assign t[63343] = t[63342] ^ n[63343];
assign t[63344] = t[63343] ^ n[63344];
assign t[63345] = t[63344] ^ n[63345];
assign t[63346] = t[63345] ^ n[63346];
assign t[63347] = t[63346] ^ n[63347];
assign t[63348] = t[63347] ^ n[63348];
assign t[63349] = t[63348] ^ n[63349];
assign t[63350] = t[63349] ^ n[63350];
assign t[63351] = t[63350] ^ n[63351];
assign t[63352] = t[63351] ^ n[63352];
assign t[63353] = t[63352] ^ n[63353];
assign t[63354] = t[63353] ^ n[63354];
assign t[63355] = t[63354] ^ n[63355];
assign t[63356] = t[63355] ^ n[63356];
assign t[63357] = t[63356] ^ n[63357];
assign t[63358] = t[63357] ^ n[63358];
assign t[63359] = t[63358] ^ n[63359];
assign t[63360] = t[63359] ^ n[63360];
assign t[63361] = t[63360] ^ n[63361];
assign t[63362] = t[63361] ^ n[63362];
assign t[63363] = t[63362] ^ n[63363];
assign t[63364] = t[63363] ^ n[63364];
assign t[63365] = t[63364] ^ n[63365];
assign t[63366] = t[63365] ^ n[63366];
assign t[63367] = t[63366] ^ n[63367];
assign t[63368] = t[63367] ^ n[63368];
assign t[63369] = t[63368] ^ n[63369];
assign t[63370] = t[63369] ^ n[63370];
assign t[63371] = t[63370] ^ n[63371];
assign t[63372] = t[63371] ^ n[63372];
assign t[63373] = t[63372] ^ n[63373];
assign t[63374] = t[63373] ^ n[63374];
assign t[63375] = t[63374] ^ n[63375];
assign t[63376] = t[63375] ^ n[63376];
assign t[63377] = t[63376] ^ n[63377];
assign t[63378] = t[63377] ^ n[63378];
assign t[63379] = t[63378] ^ n[63379];
assign t[63380] = t[63379] ^ n[63380];
assign t[63381] = t[63380] ^ n[63381];
assign t[63382] = t[63381] ^ n[63382];
assign t[63383] = t[63382] ^ n[63383];
assign t[63384] = t[63383] ^ n[63384];
assign t[63385] = t[63384] ^ n[63385];
assign t[63386] = t[63385] ^ n[63386];
assign t[63387] = t[63386] ^ n[63387];
assign t[63388] = t[63387] ^ n[63388];
assign t[63389] = t[63388] ^ n[63389];
assign t[63390] = t[63389] ^ n[63390];
assign t[63391] = t[63390] ^ n[63391];
assign t[63392] = t[63391] ^ n[63392];
assign t[63393] = t[63392] ^ n[63393];
assign t[63394] = t[63393] ^ n[63394];
assign t[63395] = t[63394] ^ n[63395];
assign t[63396] = t[63395] ^ n[63396];
assign t[63397] = t[63396] ^ n[63397];
assign t[63398] = t[63397] ^ n[63398];
assign t[63399] = t[63398] ^ n[63399];
assign t[63400] = t[63399] ^ n[63400];
assign t[63401] = t[63400] ^ n[63401];
assign t[63402] = t[63401] ^ n[63402];
assign t[63403] = t[63402] ^ n[63403];
assign t[63404] = t[63403] ^ n[63404];
assign t[63405] = t[63404] ^ n[63405];
assign t[63406] = t[63405] ^ n[63406];
assign t[63407] = t[63406] ^ n[63407];
assign t[63408] = t[63407] ^ n[63408];
assign t[63409] = t[63408] ^ n[63409];
assign t[63410] = t[63409] ^ n[63410];
assign t[63411] = t[63410] ^ n[63411];
assign t[63412] = t[63411] ^ n[63412];
assign t[63413] = t[63412] ^ n[63413];
assign t[63414] = t[63413] ^ n[63414];
assign t[63415] = t[63414] ^ n[63415];
assign t[63416] = t[63415] ^ n[63416];
assign t[63417] = t[63416] ^ n[63417];
assign t[63418] = t[63417] ^ n[63418];
assign t[63419] = t[63418] ^ n[63419];
assign t[63420] = t[63419] ^ n[63420];
assign t[63421] = t[63420] ^ n[63421];
assign t[63422] = t[63421] ^ n[63422];
assign t[63423] = t[63422] ^ n[63423];
assign t[63424] = t[63423] ^ n[63424];
assign t[63425] = t[63424] ^ n[63425];
assign t[63426] = t[63425] ^ n[63426];
assign t[63427] = t[63426] ^ n[63427];
assign t[63428] = t[63427] ^ n[63428];
assign t[63429] = t[63428] ^ n[63429];
assign t[63430] = t[63429] ^ n[63430];
assign t[63431] = t[63430] ^ n[63431];
assign t[63432] = t[63431] ^ n[63432];
assign t[63433] = t[63432] ^ n[63433];
assign t[63434] = t[63433] ^ n[63434];
assign t[63435] = t[63434] ^ n[63435];
assign t[63436] = t[63435] ^ n[63436];
assign t[63437] = t[63436] ^ n[63437];
assign t[63438] = t[63437] ^ n[63438];
assign t[63439] = t[63438] ^ n[63439];
assign t[63440] = t[63439] ^ n[63440];
assign t[63441] = t[63440] ^ n[63441];
assign t[63442] = t[63441] ^ n[63442];
assign t[63443] = t[63442] ^ n[63443];
assign t[63444] = t[63443] ^ n[63444];
assign t[63445] = t[63444] ^ n[63445];
assign t[63446] = t[63445] ^ n[63446];
assign t[63447] = t[63446] ^ n[63447];
assign t[63448] = t[63447] ^ n[63448];
assign t[63449] = t[63448] ^ n[63449];
assign t[63450] = t[63449] ^ n[63450];
assign t[63451] = t[63450] ^ n[63451];
assign t[63452] = t[63451] ^ n[63452];
assign t[63453] = t[63452] ^ n[63453];
assign t[63454] = t[63453] ^ n[63454];
assign t[63455] = t[63454] ^ n[63455];
assign t[63456] = t[63455] ^ n[63456];
assign t[63457] = t[63456] ^ n[63457];
assign t[63458] = t[63457] ^ n[63458];
assign t[63459] = t[63458] ^ n[63459];
assign t[63460] = t[63459] ^ n[63460];
assign t[63461] = t[63460] ^ n[63461];
assign t[63462] = t[63461] ^ n[63462];
assign t[63463] = t[63462] ^ n[63463];
assign t[63464] = t[63463] ^ n[63464];
assign t[63465] = t[63464] ^ n[63465];
assign t[63466] = t[63465] ^ n[63466];
assign t[63467] = t[63466] ^ n[63467];
assign t[63468] = t[63467] ^ n[63468];
assign t[63469] = t[63468] ^ n[63469];
assign t[63470] = t[63469] ^ n[63470];
assign t[63471] = t[63470] ^ n[63471];
assign t[63472] = t[63471] ^ n[63472];
assign t[63473] = t[63472] ^ n[63473];
assign t[63474] = t[63473] ^ n[63474];
assign t[63475] = t[63474] ^ n[63475];
assign t[63476] = t[63475] ^ n[63476];
assign t[63477] = t[63476] ^ n[63477];
assign t[63478] = t[63477] ^ n[63478];
assign t[63479] = t[63478] ^ n[63479];
assign t[63480] = t[63479] ^ n[63480];
assign t[63481] = t[63480] ^ n[63481];
assign t[63482] = t[63481] ^ n[63482];
assign t[63483] = t[63482] ^ n[63483];
assign t[63484] = t[63483] ^ n[63484];
assign t[63485] = t[63484] ^ n[63485];
assign t[63486] = t[63485] ^ n[63486];
assign t[63487] = t[63486] ^ n[63487];
assign t[63488] = t[63487] ^ n[63488];
assign t[63489] = t[63488] ^ n[63489];
assign t[63490] = t[63489] ^ n[63490];
assign t[63491] = t[63490] ^ n[63491];
assign t[63492] = t[63491] ^ n[63492];
assign t[63493] = t[63492] ^ n[63493];
assign t[63494] = t[63493] ^ n[63494];
assign t[63495] = t[63494] ^ n[63495];
assign t[63496] = t[63495] ^ n[63496];
assign t[63497] = t[63496] ^ n[63497];
assign t[63498] = t[63497] ^ n[63498];
assign t[63499] = t[63498] ^ n[63499];
assign t[63500] = t[63499] ^ n[63500];
assign t[63501] = t[63500] ^ n[63501];
assign t[63502] = t[63501] ^ n[63502];
assign t[63503] = t[63502] ^ n[63503];
assign t[63504] = t[63503] ^ n[63504];
assign t[63505] = t[63504] ^ n[63505];
assign t[63506] = t[63505] ^ n[63506];
assign t[63507] = t[63506] ^ n[63507];
assign t[63508] = t[63507] ^ n[63508];
assign t[63509] = t[63508] ^ n[63509];
assign t[63510] = t[63509] ^ n[63510];
assign t[63511] = t[63510] ^ n[63511];
assign t[63512] = t[63511] ^ n[63512];
assign t[63513] = t[63512] ^ n[63513];
assign t[63514] = t[63513] ^ n[63514];
assign t[63515] = t[63514] ^ n[63515];
assign t[63516] = t[63515] ^ n[63516];
assign t[63517] = t[63516] ^ n[63517];
assign t[63518] = t[63517] ^ n[63518];
assign t[63519] = t[63518] ^ n[63519];
assign t[63520] = t[63519] ^ n[63520];
assign t[63521] = t[63520] ^ n[63521];
assign t[63522] = t[63521] ^ n[63522];
assign t[63523] = t[63522] ^ n[63523];
assign t[63524] = t[63523] ^ n[63524];
assign t[63525] = t[63524] ^ n[63525];
assign t[63526] = t[63525] ^ n[63526];
assign t[63527] = t[63526] ^ n[63527];
assign t[63528] = t[63527] ^ n[63528];
assign t[63529] = t[63528] ^ n[63529];
assign t[63530] = t[63529] ^ n[63530];
assign t[63531] = t[63530] ^ n[63531];
assign t[63532] = t[63531] ^ n[63532];
assign t[63533] = t[63532] ^ n[63533];
assign t[63534] = t[63533] ^ n[63534];
assign t[63535] = t[63534] ^ n[63535];
assign t[63536] = t[63535] ^ n[63536];
assign t[63537] = t[63536] ^ n[63537];
assign t[63538] = t[63537] ^ n[63538];
assign t[63539] = t[63538] ^ n[63539];
assign t[63540] = t[63539] ^ n[63540];
assign t[63541] = t[63540] ^ n[63541];
assign t[63542] = t[63541] ^ n[63542];
assign t[63543] = t[63542] ^ n[63543];
assign t[63544] = t[63543] ^ n[63544];
assign t[63545] = t[63544] ^ n[63545];
assign t[63546] = t[63545] ^ n[63546];
assign t[63547] = t[63546] ^ n[63547];
assign t[63548] = t[63547] ^ n[63548];
assign t[63549] = t[63548] ^ n[63549];
assign t[63550] = t[63549] ^ n[63550];
assign t[63551] = t[63550] ^ n[63551];
assign t[63552] = t[63551] ^ n[63552];
assign t[63553] = t[63552] ^ n[63553];
assign t[63554] = t[63553] ^ n[63554];
assign t[63555] = t[63554] ^ n[63555];
assign t[63556] = t[63555] ^ n[63556];
assign t[63557] = t[63556] ^ n[63557];
assign t[63558] = t[63557] ^ n[63558];
assign t[63559] = t[63558] ^ n[63559];
assign t[63560] = t[63559] ^ n[63560];
assign t[63561] = t[63560] ^ n[63561];
assign t[63562] = t[63561] ^ n[63562];
assign t[63563] = t[63562] ^ n[63563];
assign t[63564] = t[63563] ^ n[63564];
assign t[63565] = t[63564] ^ n[63565];
assign t[63566] = t[63565] ^ n[63566];
assign t[63567] = t[63566] ^ n[63567];
assign t[63568] = t[63567] ^ n[63568];
assign t[63569] = t[63568] ^ n[63569];
assign t[63570] = t[63569] ^ n[63570];
assign t[63571] = t[63570] ^ n[63571];
assign t[63572] = t[63571] ^ n[63572];
assign t[63573] = t[63572] ^ n[63573];
assign t[63574] = t[63573] ^ n[63574];
assign t[63575] = t[63574] ^ n[63575];
assign t[63576] = t[63575] ^ n[63576];
assign t[63577] = t[63576] ^ n[63577];
assign t[63578] = t[63577] ^ n[63578];
assign t[63579] = t[63578] ^ n[63579];
assign t[63580] = t[63579] ^ n[63580];
assign t[63581] = t[63580] ^ n[63581];
assign t[63582] = t[63581] ^ n[63582];
assign t[63583] = t[63582] ^ n[63583];
assign t[63584] = t[63583] ^ n[63584];
assign t[63585] = t[63584] ^ n[63585];
assign t[63586] = t[63585] ^ n[63586];
assign t[63587] = t[63586] ^ n[63587];
assign t[63588] = t[63587] ^ n[63588];
assign t[63589] = t[63588] ^ n[63589];
assign t[63590] = t[63589] ^ n[63590];
assign t[63591] = t[63590] ^ n[63591];
assign t[63592] = t[63591] ^ n[63592];
assign t[63593] = t[63592] ^ n[63593];
assign t[63594] = t[63593] ^ n[63594];
assign t[63595] = t[63594] ^ n[63595];
assign t[63596] = t[63595] ^ n[63596];
assign t[63597] = t[63596] ^ n[63597];
assign t[63598] = t[63597] ^ n[63598];
assign t[63599] = t[63598] ^ n[63599];
assign t[63600] = t[63599] ^ n[63600];
assign t[63601] = t[63600] ^ n[63601];
assign t[63602] = t[63601] ^ n[63602];
assign t[63603] = t[63602] ^ n[63603];
assign t[63604] = t[63603] ^ n[63604];
assign t[63605] = t[63604] ^ n[63605];
assign t[63606] = t[63605] ^ n[63606];
assign t[63607] = t[63606] ^ n[63607];
assign t[63608] = t[63607] ^ n[63608];
assign t[63609] = t[63608] ^ n[63609];
assign t[63610] = t[63609] ^ n[63610];
assign t[63611] = t[63610] ^ n[63611];
assign t[63612] = t[63611] ^ n[63612];
assign t[63613] = t[63612] ^ n[63613];
assign t[63614] = t[63613] ^ n[63614];
assign t[63615] = t[63614] ^ n[63615];
assign t[63616] = t[63615] ^ n[63616];
assign t[63617] = t[63616] ^ n[63617];
assign t[63618] = t[63617] ^ n[63618];
assign t[63619] = t[63618] ^ n[63619];
assign t[63620] = t[63619] ^ n[63620];
assign t[63621] = t[63620] ^ n[63621];
assign t[63622] = t[63621] ^ n[63622];
assign t[63623] = t[63622] ^ n[63623];
assign t[63624] = t[63623] ^ n[63624];
assign t[63625] = t[63624] ^ n[63625];
assign t[63626] = t[63625] ^ n[63626];
assign t[63627] = t[63626] ^ n[63627];
assign t[63628] = t[63627] ^ n[63628];
assign t[63629] = t[63628] ^ n[63629];
assign t[63630] = t[63629] ^ n[63630];
assign t[63631] = t[63630] ^ n[63631];
assign t[63632] = t[63631] ^ n[63632];
assign t[63633] = t[63632] ^ n[63633];
assign t[63634] = t[63633] ^ n[63634];
assign t[63635] = t[63634] ^ n[63635];
assign t[63636] = t[63635] ^ n[63636];
assign t[63637] = t[63636] ^ n[63637];
assign t[63638] = t[63637] ^ n[63638];
assign t[63639] = t[63638] ^ n[63639];
assign t[63640] = t[63639] ^ n[63640];
assign t[63641] = t[63640] ^ n[63641];
assign t[63642] = t[63641] ^ n[63642];
assign t[63643] = t[63642] ^ n[63643];
assign t[63644] = t[63643] ^ n[63644];
assign t[63645] = t[63644] ^ n[63645];
assign t[63646] = t[63645] ^ n[63646];
assign t[63647] = t[63646] ^ n[63647];
assign t[63648] = t[63647] ^ n[63648];
assign t[63649] = t[63648] ^ n[63649];
assign t[63650] = t[63649] ^ n[63650];
assign t[63651] = t[63650] ^ n[63651];
assign t[63652] = t[63651] ^ n[63652];
assign t[63653] = t[63652] ^ n[63653];
assign t[63654] = t[63653] ^ n[63654];
assign t[63655] = t[63654] ^ n[63655];
assign t[63656] = t[63655] ^ n[63656];
assign t[63657] = t[63656] ^ n[63657];
assign t[63658] = t[63657] ^ n[63658];
assign t[63659] = t[63658] ^ n[63659];
assign t[63660] = t[63659] ^ n[63660];
assign t[63661] = t[63660] ^ n[63661];
assign t[63662] = t[63661] ^ n[63662];
assign t[63663] = t[63662] ^ n[63663];
assign t[63664] = t[63663] ^ n[63664];
assign t[63665] = t[63664] ^ n[63665];
assign t[63666] = t[63665] ^ n[63666];
assign t[63667] = t[63666] ^ n[63667];
assign t[63668] = t[63667] ^ n[63668];
assign t[63669] = t[63668] ^ n[63669];
assign t[63670] = t[63669] ^ n[63670];
assign t[63671] = t[63670] ^ n[63671];
assign t[63672] = t[63671] ^ n[63672];
assign t[63673] = t[63672] ^ n[63673];
assign t[63674] = t[63673] ^ n[63674];
assign t[63675] = t[63674] ^ n[63675];
assign t[63676] = t[63675] ^ n[63676];
assign t[63677] = t[63676] ^ n[63677];
assign t[63678] = t[63677] ^ n[63678];
assign t[63679] = t[63678] ^ n[63679];
assign t[63680] = t[63679] ^ n[63680];
assign t[63681] = t[63680] ^ n[63681];
assign t[63682] = t[63681] ^ n[63682];
assign t[63683] = t[63682] ^ n[63683];
assign t[63684] = t[63683] ^ n[63684];
assign t[63685] = t[63684] ^ n[63685];
assign t[63686] = t[63685] ^ n[63686];
assign t[63687] = t[63686] ^ n[63687];
assign t[63688] = t[63687] ^ n[63688];
assign t[63689] = t[63688] ^ n[63689];
assign t[63690] = t[63689] ^ n[63690];
assign t[63691] = t[63690] ^ n[63691];
assign t[63692] = t[63691] ^ n[63692];
assign t[63693] = t[63692] ^ n[63693];
assign t[63694] = t[63693] ^ n[63694];
assign t[63695] = t[63694] ^ n[63695];
assign t[63696] = t[63695] ^ n[63696];
assign t[63697] = t[63696] ^ n[63697];
assign t[63698] = t[63697] ^ n[63698];
assign t[63699] = t[63698] ^ n[63699];
assign t[63700] = t[63699] ^ n[63700];
assign t[63701] = t[63700] ^ n[63701];
assign t[63702] = t[63701] ^ n[63702];
assign t[63703] = t[63702] ^ n[63703];
assign t[63704] = t[63703] ^ n[63704];
assign t[63705] = t[63704] ^ n[63705];
assign t[63706] = t[63705] ^ n[63706];
assign t[63707] = t[63706] ^ n[63707];
assign t[63708] = t[63707] ^ n[63708];
assign t[63709] = t[63708] ^ n[63709];
assign t[63710] = t[63709] ^ n[63710];
assign t[63711] = t[63710] ^ n[63711];
assign t[63712] = t[63711] ^ n[63712];
assign t[63713] = t[63712] ^ n[63713];
assign t[63714] = t[63713] ^ n[63714];
assign t[63715] = t[63714] ^ n[63715];
assign t[63716] = t[63715] ^ n[63716];
assign t[63717] = t[63716] ^ n[63717];
assign t[63718] = t[63717] ^ n[63718];
assign t[63719] = t[63718] ^ n[63719];
assign t[63720] = t[63719] ^ n[63720];
assign t[63721] = t[63720] ^ n[63721];
assign t[63722] = t[63721] ^ n[63722];
assign t[63723] = t[63722] ^ n[63723];
assign t[63724] = t[63723] ^ n[63724];
assign t[63725] = t[63724] ^ n[63725];
assign t[63726] = t[63725] ^ n[63726];
assign t[63727] = t[63726] ^ n[63727];
assign t[63728] = t[63727] ^ n[63728];
assign t[63729] = t[63728] ^ n[63729];
assign t[63730] = t[63729] ^ n[63730];
assign t[63731] = t[63730] ^ n[63731];
assign t[63732] = t[63731] ^ n[63732];
assign t[63733] = t[63732] ^ n[63733];
assign t[63734] = t[63733] ^ n[63734];
assign t[63735] = t[63734] ^ n[63735];
assign t[63736] = t[63735] ^ n[63736];
assign t[63737] = t[63736] ^ n[63737];
assign t[63738] = t[63737] ^ n[63738];
assign t[63739] = t[63738] ^ n[63739];
assign t[63740] = t[63739] ^ n[63740];
assign t[63741] = t[63740] ^ n[63741];
assign t[63742] = t[63741] ^ n[63742];
assign t[63743] = t[63742] ^ n[63743];
assign t[63744] = t[63743] ^ n[63744];
assign t[63745] = t[63744] ^ n[63745];
assign t[63746] = t[63745] ^ n[63746];
assign t[63747] = t[63746] ^ n[63747];
assign t[63748] = t[63747] ^ n[63748];
assign t[63749] = t[63748] ^ n[63749];
assign t[63750] = t[63749] ^ n[63750];
assign t[63751] = t[63750] ^ n[63751];
assign t[63752] = t[63751] ^ n[63752];
assign t[63753] = t[63752] ^ n[63753];
assign t[63754] = t[63753] ^ n[63754];
assign t[63755] = t[63754] ^ n[63755];
assign t[63756] = t[63755] ^ n[63756];
assign t[63757] = t[63756] ^ n[63757];
assign t[63758] = t[63757] ^ n[63758];
assign t[63759] = t[63758] ^ n[63759];
assign t[63760] = t[63759] ^ n[63760];
assign t[63761] = t[63760] ^ n[63761];
assign t[63762] = t[63761] ^ n[63762];
assign t[63763] = t[63762] ^ n[63763];
assign t[63764] = t[63763] ^ n[63764];
assign t[63765] = t[63764] ^ n[63765];
assign t[63766] = t[63765] ^ n[63766];
assign t[63767] = t[63766] ^ n[63767];
assign t[63768] = t[63767] ^ n[63768];
assign t[63769] = t[63768] ^ n[63769];
assign t[63770] = t[63769] ^ n[63770];
assign t[63771] = t[63770] ^ n[63771];
assign t[63772] = t[63771] ^ n[63772];
assign t[63773] = t[63772] ^ n[63773];
assign t[63774] = t[63773] ^ n[63774];
assign t[63775] = t[63774] ^ n[63775];
assign t[63776] = t[63775] ^ n[63776];
assign t[63777] = t[63776] ^ n[63777];
assign t[63778] = t[63777] ^ n[63778];
assign t[63779] = t[63778] ^ n[63779];
assign t[63780] = t[63779] ^ n[63780];
assign t[63781] = t[63780] ^ n[63781];
assign t[63782] = t[63781] ^ n[63782];
assign t[63783] = t[63782] ^ n[63783];
assign t[63784] = t[63783] ^ n[63784];
assign t[63785] = t[63784] ^ n[63785];
assign t[63786] = t[63785] ^ n[63786];
assign t[63787] = t[63786] ^ n[63787];
assign t[63788] = t[63787] ^ n[63788];
assign t[63789] = t[63788] ^ n[63789];
assign t[63790] = t[63789] ^ n[63790];
assign t[63791] = t[63790] ^ n[63791];
assign t[63792] = t[63791] ^ n[63792];
assign t[63793] = t[63792] ^ n[63793];
assign t[63794] = t[63793] ^ n[63794];
assign t[63795] = t[63794] ^ n[63795];
assign t[63796] = t[63795] ^ n[63796];
assign t[63797] = t[63796] ^ n[63797];
assign t[63798] = t[63797] ^ n[63798];
assign t[63799] = t[63798] ^ n[63799];
assign t[63800] = t[63799] ^ n[63800];
assign t[63801] = t[63800] ^ n[63801];
assign t[63802] = t[63801] ^ n[63802];
assign t[63803] = t[63802] ^ n[63803];
assign t[63804] = t[63803] ^ n[63804];
assign t[63805] = t[63804] ^ n[63805];
assign t[63806] = t[63805] ^ n[63806];
assign t[63807] = t[63806] ^ n[63807];
assign t[63808] = t[63807] ^ n[63808];
assign t[63809] = t[63808] ^ n[63809];
assign t[63810] = t[63809] ^ n[63810];
assign t[63811] = t[63810] ^ n[63811];
assign t[63812] = t[63811] ^ n[63812];
assign t[63813] = t[63812] ^ n[63813];
assign t[63814] = t[63813] ^ n[63814];
assign t[63815] = t[63814] ^ n[63815];
assign t[63816] = t[63815] ^ n[63816];
assign t[63817] = t[63816] ^ n[63817];
assign t[63818] = t[63817] ^ n[63818];
assign t[63819] = t[63818] ^ n[63819];
assign t[63820] = t[63819] ^ n[63820];
assign t[63821] = t[63820] ^ n[63821];
assign t[63822] = t[63821] ^ n[63822];
assign t[63823] = t[63822] ^ n[63823];
assign t[63824] = t[63823] ^ n[63824];
assign t[63825] = t[63824] ^ n[63825];
assign t[63826] = t[63825] ^ n[63826];
assign t[63827] = t[63826] ^ n[63827];
assign t[63828] = t[63827] ^ n[63828];
assign t[63829] = t[63828] ^ n[63829];
assign t[63830] = t[63829] ^ n[63830];
assign t[63831] = t[63830] ^ n[63831];
assign t[63832] = t[63831] ^ n[63832];
assign t[63833] = t[63832] ^ n[63833];
assign t[63834] = t[63833] ^ n[63834];
assign t[63835] = t[63834] ^ n[63835];
assign t[63836] = t[63835] ^ n[63836];
assign t[63837] = t[63836] ^ n[63837];
assign t[63838] = t[63837] ^ n[63838];
assign t[63839] = t[63838] ^ n[63839];
assign t[63840] = t[63839] ^ n[63840];
assign t[63841] = t[63840] ^ n[63841];
assign t[63842] = t[63841] ^ n[63842];
assign t[63843] = t[63842] ^ n[63843];
assign t[63844] = t[63843] ^ n[63844];
assign t[63845] = t[63844] ^ n[63845];
assign t[63846] = t[63845] ^ n[63846];
assign t[63847] = t[63846] ^ n[63847];
assign t[63848] = t[63847] ^ n[63848];
assign t[63849] = t[63848] ^ n[63849];
assign t[63850] = t[63849] ^ n[63850];
assign t[63851] = t[63850] ^ n[63851];
assign t[63852] = t[63851] ^ n[63852];
assign t[63853] = t[63852] ^ n[63853];
assign t[63854] = t[63853] ^ n[63854];
assign t[63855] = t[63854] ^ n[63855];
assign t[63856] = t[63855] ^ n[63856];
assign t[63857] = t[63856] ^ n[63857];
assign t[63858] = t[63857] ^ n[63858];
assign t[63859] = t[63858] ^ n[63859];
assign t[63860] = t[63859] ^ n[63860];
assign t[63861] = t[63860] ^ n[63861];
assign t[63862] = t[63861] ^ n[63862];
assign t[63863] = t[63862] ^ n[63863];
assign t[63864] = t[63863] ^ n[63864];
assign t[63865] = t[63864] ^ n[63865];
assign t[63866] = t[63865] ^ n[63866];
assign t[63867] = t[63866] ^ n[63867];
assign t[63868] = t[63867] ^ n[63868];
assign t[63869] = t[63868] ^ n[63869];
assign t[63870] = t[63869] ^ n[63870];
assign t[63871] = t[63870] ^ n[63871];
assign t[63872] = t[63871] ^ n[63872];
assign t[63873] = t[63872] ^ n[63873];
assign t[63874] = t[63873] ^ n[63874];
assign t[63875] = t[63874] ^ n[63875];
assign t[63876] = t[63875] ^ n[63876];
assign t[63877] = t[63876] ^ n[63877];
assign t[63878] = t[63877] ^ n[63878];
assign t[63879] = t[63878] ^ n[63879];
assign t[63880] = t[63879] ^ n[63880];
assign t[63881] = t[63880] ^ n[63881];
assign t[63882] = t[63881] ^ n[63882];
assign t[63883] = t[63882] ^ n[63883];
assign t[63884] = t[63883] ^ n[63884];
assign t[63885] = t[63884] ^ n[63885];
assign t[63886] = t[63885] ^ n[63886];
assign t[63887] = t[63886] ^ n[63887];
assign t[63888] = t[63887] ^ n[63888];
assign t[63889] = t[63888] ^ n[63889];
assign t[63890] = t[63889] ^ n[63890];
assign t[63891] = t[63890] ^ n[63891];
assign t[63892] = t[63891] ^ n[63892];
assign t[63893] = t[63892] ^ n[63893];
assign t[63894] = t[63893] ^ n[63894];
assign t[63895] = t[63894] ^ n[63895];
assign t[63896] = t[63895] ^ n[63896];
assign t[63897] = t[63896] ^ n[63897];
assign t[63898] = t[63897] ^ n[63898];
assign t[63899] = t[63898] ^ n[63899];
assign t[63900] = t[63899] ^ n[63900];
assign t[63901] = t[63900] ^ n[63901];
assign t[63902] = t[63901] ^ n[63902];
assign t[63903] = t[63902] ^ n[63903];
assign t[63904] = t[63903] ^ n[63904];
assign t[63905] = t[63904] ^ n[63905];
assign t[63906] = t[63905] ^ n[63906];
assign t[63907] = t[63906] ^ n[63907];
assign t[63908] = t[63907] ^ n[63908];
assign t[63909] = t[63908] ^ n[63909];
assign t[63910] = t[63909] ^ n[63910];
assign t[63911] = t[63910] ^ n[63911];
assign t[63912] = t[63911] ^ n[63912];
assign t[63913] = t[63912] ^ n[63913];
assign t[63914] = t[63913] ^ n[63914];
assign t[63915] = t[63914] ^ n[63915];
assign t[63916] = t[63915] ^ n[63916];
assign t[63917] = t[63916] ^ n[63917];
assign t[63918] = t[63917] ^ n[63918];
assign t[63919] = t[63918] ^ n[63919];
assign t[63920] = t[63919] ^ n[63920];
assign t[63921] = t[63920] ^ n[63921];
assign t[63922] = t[63921] ^ n[63922];
assign t[63923] = t[63922] ^ n[63923];
assign t[63924] = t[63923] ^ n[63924];
assign t[63925] = t[63924] ^ n[63925];
assign t[63926] = t[63925] ^ n[63926];
assign t[63927] = t[63926] ^ n[63927];
assign t[63928] = t[63927] ^ n[63928];
assign t[63929] = t[63928] ^ n[63929];
assign t[63930] = t[63929] ^ n[63930];
assign t[63931] = t[63930] ^ n[63931];
assign t[63932] = t[63931] ^ n[63932];
assign t[63933] = t[63932] ^ n[63933];
assign t[63934] = t[63933] ^ n[63934];
assign t[63935] = t[63934] ^ n[63935];
assign t[63936] = t[63935] ^ n[63936];
assign t[63937] = t[63936] ^ n[63937];
assign t[63938] = t[63937] ^ n[63938];
assign t[63939] = t[63938] ^ n[63939];
assign t[63940] = t[63939] ^ n[63940];
assign t[63941] = t[63940] ^ n[63941];
assign t[63942] = t[63941] ^ n[63942];
assign t[63943] = t[63942] ^ n[63943];
assign t[63944] = t[63943] ^ n[63944];
assign t[63945] = t[63944] ^ n[63945];
assign t[63946] = t[63945] ^ n[63946];
assign t[63947] = t[63946] ^ n[63947];
assign t[63948] = t[63947] ^ n[63948];
assign t[63949] = t[63948] ^ n[63949];
assign t[63950] = t[63949] ^ n[63950];
assign t[63951] = t[63950] ^ n[63951];
assign t[63952] = t[63951] ^ n[63952];
assign t[63953] = t[63952] ^ n[63953];
assign t[63954] = t[63953] ^ n[63954];
assign t[63955] = t[63954] ^ n[63955];
assign t[63956] = t[63955] ^ n[63956];
assign t[63957] = t[63956] ^ n[63957];
assign t[63958] = t[63957] ^ n[63958];
assign t[63959] = t[63958] ^ n[63959];
assign t[63960] = t[63959] ^ n[63960];
assign t[63961] = t[63960] ^ n[63961];
assign t[63962] = t[63961] ^ n[63962];
assign t[63963] = t[63962] ^ n[63963];
assign t[63964] = t[63963] ^ n[63964];
assign t[63965] = t[63964] ^ n[63965];
assign t[63966] = t[63965] ^ n[63966];
assign t[63967] = t[63966] ^ n[63967];
assign t[63968] = t[63967] ^ n[63968];
assign t[63969] = t[63968] ^ n[63969];
assign t[63970] = t[63969] ^ n[63970];
assign t[63971] = t[63970] ^ n[63971];
assign t[63972] = t[63971] ^ n[63972];
assign t[63973] = t[63972] ^ n[63973];
assign t[63974] = t[63973] ^ n[63974];
assign t[63975] = t[63974] ^ n[63975];
assign t[63976] = t[63975] ^ n[63976];
assign t[63977] = t[63976] ^ n[63977];
assign t[63978] = t[63977] ^ n[63978];
assign t[63979] = t[63978] ^ n[63979];
assign t[63980] = t[63979] ^ n[63980];
assign t[63981] = t[63980] ^ n[63981];
assign t[63982] = t[63981] ^ n[63982];
assign t[63983] = t[63982] ^ n[63983];
assign t[63984] = t[63983] ^ n[63984];
assign t[63985] = t[63984] ^ n[63985];
assign t[63986] = t[63985] ^ n[63986];
assign t[63987] = t[63986] ^ n[63987];
assign t[63988] = t[63987] ^ n[63988];
assign t[63989] = t[63988] ^ n[63989];
assign t[63990] = t[63989] ^ n[63990];
assign t[63991] = t[63990] ^ n[63991];
assign t[63992] = t[63991] ^ n[63992];
assign t[63993] = t[63992] ^ n[63993];
assign t[63994] = t[63993] ^ n[63994];
assign t[63995] = t[63994] ^ n[63995];
assign t[63996] = t[63995] ^ n[63996];
assign t[63997] = t[63996] ^ n[63997];
assign t[63998] = t[63997] ^ n[63998];
assign t[63999] = t[63998] ^ n[63999];
assign t[64000] = t[63999] ^ n[64000];
assign t[64001] = t[64000] ^ n[64001];
assign t[64002] = t[64001] ^ n[64002];
assign t[64003] = t[64002] ^ n[64003];
assign t[64004] = t[64003] ^ n[64004];
assign t[64005] = t[64004] ^ n[64005];
assign t[64006] = t[64005] ^ n[64006];
assign t[64007] = t[64006] ^ n[64007];
assign t[64008] = t[64007] ^ n[64008];
assign t[64009] = t[64008] ^ n[64009];
assign t[64010] = t[64009] ^ n[64010];
assign t[64011] = t[64010] ^ n[64011];
assign t[64012] = t[64011] ^ n[64012];
assign t[64013] = t[64012] ^ n[64013];
assign t[64014] = t[64013] ^ n[64014];
assign t[64015] = t[64014] ^ n[64015];
assign t[64016] = t[64015] ^ n[64016];
assign t[64017] = t[64016] ^ n[64017];
assign t[64018] = t[64017] ^ n[64018];
assign t[64019] = t[64018] ^ n[64019];
assign t[64020] = t[64019] ^ n[64020];
assign t[64021] = t[64020] ^ n[64021];
assign t[64022] = t[64021] ^ n[64022];
assign t[64023] = t[64022] ^ n[64023];
assign t[64024] = t[64023] ^ n[64024];
assign t[64025] = t[64024] ^ n[64025];
assign t[64026] = t[64025] ^ n[64026];
assign t[64027] = t[64026] ^ n[64027];
assign t[64028] = t[64027] ^ n[64028];
assign t[64029] = t[64028] ^ n[64029];
assign t[64030] = t[64029] ^ n[64030];
assign t[64031] = t[64030] ^ n[64031];
assign t[64032] = t[64031] ^ n[64032];
assign t[64033] = t[64032] ^ n[64033];
assign t[64034] = t[64033] ^ n[64034];
assign t[64035] = t[64034] ^ n[64035];
assign t[64036] = t[64035] ^ n[64036];
assign t[64037] = t[64036] ^ n[64037];
assign t[64038] = t[64037] ^ n[64038];
assign t[64039] = t[64038] ^ n[64039];
assign t[64040] = t[64039] ^ n[64040];
assign t[64041] = t[64040] ^ n[64041];
assign t[64042] = t[64041] ^ n[64042];
assign t[64043] = t[64042] ^ n[64043];
assign t[64044] = t[64043] ^ n[64044];
assign t[64045] = t[64044] ^ n[64045];
assign t[64046] = t[64045] ^ n[64046];
assign t[64047] = t[64046] ^ n[64047];
assign t[64048] = t[64047] ^ n[64048];
assign t[64049] = t[64048] ^ n[64049];
assign t[64050] = t[64049] ^ n[64050];
assign t[64051] = t[64050] ^ n[64051];
assign t[64052] = t[64051] ^ n[64052];
assign t[64053] = t[64052] ^ n[64053];
assign t[64054] = t[64053] ^ n[64054];
assign t[64055] = t[64054] ^ n[64055];
assign t[64056] = t[64055] ^ n[64056];
assign t[64057] = t[64056] ^ n[64057];
assign t[64058] = t[64057] ^ n[64058];
assign t[64059] = t[64058] ^ n[64059];
assign t[64060] = t[64059] ^ n[64060];
assign t[64061] = t[64060] ^ n[64061];
assign t[64062] = t[64061] ^ n[64062];
assign t[64063] = t[64062] ^ n[64063];
assign t[64064] = t[64063] ^ n[64064];
assign t[64065] = t[64064] ^ n[64065];
assign t[64066] = t[64065] ^ n[64066];
assign t[64067] = t[64066] ^ n[64067];
assign t[64068] = t[64067] ^ n[64068];
assign t[64069] = t[64068] ^ n[64069];
assign t[64070] = t[64069] ^ n[64070];
assign t[64071] = t[64070] ^ n[64071];
assign t[64072] = t[64071] ^ n[64072];
assign t[64073] = t[64072] ^ n[64073];
assign t[64074] = t[64073] ^ n[64074];
assign t[64075] = t[64074] ^ n[64075];
assign t[64076] = t[64075] ^ n[64076];
assign t[64077] = t[64076] ^ n[64077];
assign t[64078] = t[64077] ^ n[64078];
assign t[64079] = t[64078] ^ n[64079];
assign t[64080] = t[64079] ^ n[64080];
assign t[64081] = t[64080] ^ n[64081];
assign t[64082] = t[64081] ^ n[64082];
assign t[64083] = t[64082] ^ n[64083];
assign t[64084] = t[64083] ^ n[64084];
assign t[64085] = t[64084] ^ n[64085];
assign t[64086] = t[64085] ^ n[64086];
assign t[64087] = t[64086] ^ n[64087];
assign t[64088] = t[64087] ^ n[64088];
assign t[64089] = t[64088] ^ n[64089];
assign t[64090] = t[64089] ^ n[64090];
assign t[64091] = t[64090] ^ n[64091];
assign t[64092] = t[64091] ^ n[64092];
assign t[64093] = t[64092] ^ n[64093];
assign t[64094] = t[64093] ^ n[64094];
assign t[64095] = t[64094] ^ n[64095];
assign t[64096] = t[64095] ^ n[64096];
assign t[64097] = t[64096] ^ n[64097];
assign t[64098] = t[64097] ^ n[64098];
assign t[64099] = t[64098] ^ n[64099];
assign t[64100] = t[64099] ^ n[64100];
assign t[64101] = t[64100] ^ n[64101];
assign t[64102] = t[64101] ^ n[64102];
assign t[64103] = t[64102] ^ n[64103];
assign t[64104] = t[64103] ^ n[64104];
assign t[64105] = t[64104] ^ n[64105];
assign t[64106] = t[64105] ^ n[64106];
assign t[64107] = t[64106] ^ n[64107];
assign t[64108] = t[64107] ^ n[64108];
assign t[64109] = t[64108] ^ n[64109];
assign t[64110] = t[64109] ^ n[64110];
assign t[64111] = t[64110] ^ n[64111];
assign t[64112] = t[64111] ^ n[64112];
assign t[64113] = t[64112] ^ n[64113];
assign t[64114] = t[64113] ^ n[64114];
assign t[64115] = t[64114] ^ n[64115];
assign t[64116] = t[64115] ^ n[64116];
assign t[64117] = t[64116] ^ n[64117];
assign t[64118] = t[64117] ^ n[64118];
assign t[64119] = t[64118] ^ n[64119];
assign t[64120] = t[64119] ^ n[64120];
assign t[64121] = t[64120] ^ n[64121];
assign t[64122] = t[64121] ^ n[64122];
assign t[64123] = t[64122] ^ n[64123];
assign t[64124] = t[64123] ^ n[64124];
assign t[64125] = t[64124] ^ n[64125];
assign t[64126] = t[64125] ^ n[64126];
assign t[64127] = t[64126] ^ n[64127];
assign t[64128] = t[64127] ^ n[64128];
assign t[64129] = t[64128] ^ n[64129];
assign t[64130] = t[64129] ^ n[64130];
assign t[64131] = t[64130] ^ n[64131];
assign t[64132] = t[64131] ^ n[64132];
assign t[64133] = t[64132] ^ n[64133];
assign t[64134] = t[64133] ^ n[64134];
assign t[64135] = t[64134] ^ n[64135];
assign t[64136] = t[64135] ^ n[64136];
assign t[64137] = t[64136] ^ n[64137];
assign t[64138] = t[64137] ^ n[64138];
assign t[64139] = t[64138] ^ n[64139];
assign t[64140] = t[64139] ^ n[64140];
assign t[64141] = t[64140] ^ n[64141];
assign t[64142] = t[64141] ^ n[64142];
assign t[64143] = t[64142] ^ n[64143];
assign t[64144] = t[64143] ^ n[64144];
assign t[64145] = t[64144] ^ n[64145];
assign t[64146] = t[64145] ^ n[64146];
assign t[64147] = t[64146] ^ n[64147];
assign t[64148] = t[64147] ^ n[64148];
assign t[64149] = t[64148] ^ n[64149];
assign t[64150] = t[64149] ^ n[64150];
assign t[64151] = t[64150] ^ n[64151];
assign t[64152] = t[64151] ^ n[64152];
assign t[64153] = t[64152] ^ n[64153];
assign t[64154] = t[64153] ^ n[64154];
assign t[64155] = t[64154] ^ n[64155];
assign t[64156] = t[64155] ^ n[64156];
assign t[64157] = t[64156] ^ n[64157];
assign t[64158] = t[64157] ^ n[64158];
assign t[64159] = t[64158] ^ n[64159];
assign t[64160] = t[64159] ^ n[64160];
assign t[64161] = t[64160] ^ n[64161];
assign t[64162] = t[64161] ^ n[64162];
assign t[64163] = t[64162] ^ n[64163];
assign t[64164] = t[64163] ^ n[64164];
assign t[64165] = t[64164] ^ n[64165];
assign t[64166] = t[64165] ^ n[64166];
assign t[64167] = t[64166] ^ n[64167];
assign t[64168] = t[64167] ^ n[64168];
assign t[64169] = t[64168] ^ n[64169];
assign t[64170] = t[64169] ^ n[64170];
assign t[64171] = t[64170] ^ n[64171];
assign t[64172] = t[64171] ^ n[64172];
assign t[64173] = t[64172] ^ n[64173];
assign t[64174] = t[64173] ^ n[64174];
assign t[64175] = t[64174] ^ n[64175];
assign t[64176] = t[64175] ^ n[64176];
assign t[64177] = t[64176] ^ n[64177];
assign t[64178] = t[64177] ^ n[64178];
assign t[64179] = t[64178] ^ n[64179];
assign t[64180] = t[64179] ^ n[64180];
assign t[64181] = t[64180] ^ n[64181];
assign t[64182] = t[64181] ^ n[64182];
assign t[64183] = t[64182] ^ n[64183];
assign t[64184] = t[64183] ^ n[64184];
assign t[64185] = t[64184] ^ n[64185];
assign t[64186] = t[64185] ^ n[64186];
assign t[64187] = t[64186] ^ n[64187];
assign t[64188] = t[64187] ^ n[64188];
assign t[64189] = t[64188] ^ n[64189];
assign t[64190] = t[64189] ^ n[64190];
assign t[64191] = t[64190] ^ n[64191];
assign t[64192] = t[64191] ^ n[64192];
assign t[64193] = t[64192] ^ n[64193];
assign t[64194] = t[64193] ^ n[64194];
assign t[64195] = t[64194] ^ n[64195];
assign t[64196] = t[64195] ^ n[64196];
assign t[64197] = t[64196] ^ n[64197];
assign t[64198] = t[64197] ^ n[64198];
assign t[64199] = t[64198] ^ n[64199];
assign t[64200] = t[64199] ^ n[64200];
assign t[64201] = t[64200] ^ n[64201];
assign t[64202] = t[64201] ^ n[64202];
assign t[64203] = t[64202] ^ n[64203];
assign t[64204] = t[64203] ^ n[64204];
assign t[64205] = t[64204] ^ n[64205];
assign t[64206] = t[64205] ^ n[64206];
assign t[64207] = t[64206] ^ n[64207];
assign t[64208] = t[64207] ^ n[64208];
assign t[64209] = t[64208] ^ n[64209];
assign t[64210] = t[64209] ^ n[64210];
assign t[64211] = t[64210] ^ n[64211];
assign t[64212] = t[64211] ^ n[64212];
assign t[64213] = t[64212] ^ n[64213];
assign t[64214] = t[64213] ^ n[64214];
assign t[64215] = t[64214] ^ n[64215];
assign t[64216] = t[64215] ^ n[64216];
assign t[64217] = t[64216] ^ n[64217];
assign t[64218] = t[64217] ^ n[64218];
assign t[64219] = t[64218] ^ n[64219];
assign t[64220] = t[64219] ^ n[64220];
assign t[64221] = t[64220] ^ n[64221];
assign t[64222] = t[64221] ^ n[64222];
assign t[64223] = t[64222] ^ n[64223];
assign t[64224] = t[64223] ^ n[64224];
assign t[64225] = t[64224] ^ n[64225];
assign t[64226] = t[64225] ^ n[64226];
assign t[64227] = t[64226] ^ n[64227];
assign t[64228] = t[64227] ^ n[64228];
assign t[64229] = t[64228] ^ n[64229];
assign t[64230] = t[64229] ^ n[64230];
assign t[64231] = t[64230] ^ n[64231];
assign t[64232] = t[64231] ^ n[64232];
assign t[64233] = t[64232] ^ n[64233];
assign t[64234] = t[64233] ^ n[64234];
assign t[64235] = t[64234] ^ n[64235];
assign t[64236] = t[64235] ^ n[64236];
assign t[64237] = t[64236] ^ n[64237];
assign t[64238] = t[64237] ^ n[64238];
assign t[64239] = t[64238] ^ n[64239];
assign t[64240] = t[64239] ^ n[64240];
assign t[64241] = t[64240] ^ n[64241];
assign t[64242] = t[64241] ^ n[64242];
assign t[64243] = t[64242] ^ n[64243];
assign t[64244] = t[64243] ^ n[64244];
assign t[64245] = t[64244] ^ n[64245];
assign t[64246] = t[64245] ^ n[64246];
assign t[64247] = t[64246] ^ n[64247];
assign t[64248] = t[64247] ^ n[64248];
assign t[64249] = t[64248] ^ n[64249];
assign t[64250] = t[64249] ^ n[64250];
assign t[64251] = t[64250] ^ n[64251];
assign t[64252] = t[64251] ^ n[64252];
assign t[64253] = t[64252] ^ n[64253];
assign t[64254] = t[64253] ^ n[64254];
assign t[64255] = t[64254] ^ n[64255];
assign t[64256] = t[64255] ^ n[64256];
assign t[64257] = t[64256] ^ n[64257];
assign t[64258] = t[64257] ^ n[64258];
assign t[64259] = t[64258] ^ n[64259];
assign t[64260] = t[64259] ^ n[64260];
assign t[64261] = t[64260] ^ n[64261];
assign t[64262] = t[64261] ^ n[64262];
assign t[64263] = t[64262] ^ n[64263];
assign t[64264] = t[64263] ^ n[64264];
assign t[64265] = t[64264] ^ n[64265];
assign t[64266] = t[64265] ^ n[64266];
assign t[64267] = t[64266] ^ n[64267];
assign t[64268] = t[64267] ^ n[64268];
assign t[64269] = t[64268] ^ n[64269];
assign t[64270] = t[64269] ^ n[64270];
assign t[64271] = t[64270] ^ n[64271];
assign t[64272] = t[64271] ^ n[64272];
assign t[64273] = t[64272] ^ n[64273];
assign t[64274] = t[64273] ^ n[64274];
assign t[64275] = t[64274] ^ n[64275];
assign t[64276] = t[64275] ^ n[64276];
assign t[64277] = t[64276] ^ n[64277];
assign t[64278] = t[64277] ^ n[64278];
assign t[64279] = t[64278] ^ n[64279];
assign t[64280] = t[64279] ^ n[64280];
assign t[64281] = t[64280] ^ n[64281];
assign t[64282] = t[64281] ^ n[64282];
assign t[64283] = t[64282] ^ n[64283];
assign t[64284] = t[64283] ^ n[64284];
assign t[64285] = t[64284] ^ n[64285];
assign t[64286] = t[64285] ^ n[64286];
assign t[64287] = t[64286] ^ n[64287];
assign t[64288] = t[64287] ^ n[64288];
assign t[64289] = t[64288] ^ n[64289];
assign t[64290] = t[64289] ^ n[64290];
assign t[64291] = t[64290] ^ n[64291];
assign t[64292] = t[64291] ^ n[64292];
assign t[64293] = t[64292] ^ n[64293];
assign t[64294] = t[64293] ^ n[64294];
assign t[64295] = t[64294] ^ n[64295];
assign t[64296] = t[64295] ^ n[64296];
assign t[64297] = t[64296] ^ n[64297];
assign t[64298] = t[64297] ^ n[64298];
assign t[64299] = t[64298] ^ n[64299];
assign t[64300] = t[64299] ^ n[64300];
assign t[64301] = t[64300] ^ n[64301];
assign t[64302] = t[64301] ^ n[64302];
assign t[64303] = t[64302] ^ n[64303];
assign t[64304] = t[64303] ^ n[64304];
assign t[64305] = t[64304] ^ n[64305];
assign t[64306] = t[64305] ^ n[64306];
assign t[64307] = t[64306] ^ n[64307];
assign t[64308] = t[64307] ^ n[64308];
assign t[64309] = t[64308] ^ n[64309];
assign t[64310] = t[64309] ^ n[64310];
assign t[64311] = t[64310] ^ n[64311];
assign t[64312] = t[64311] ^ n[64312];
assign t[64313] = t[64312] ^ n[64313];
assign t[64314] = t[64313] ^ n[64314];
assign t[64315] = t[64314] ^ n[64315];
assign t[64316] = t[64315] ^ n[64316];
assign t[64317] = t[64316] ^ n[64317];
assign t[64318] = t[64317] ^ n[64318];
assign t[64319] = t[64318] ^ n[64319];
assign t[64320] = t[64319] ^ n[64320];
assign t[64321] = t[64320] ^ n[64321];
assign t[64322] = t[64321] ^ n[64322];
assign t[64323] = t[64322] ^ n[64323];
assign t[64324] = t[64323] ^ n[64324];
assign t[64325] = t[64324] ^ n[64325];
assign t[64326] = t[64325] ^ n[64326];
assign t[64327] = t[64326] ^ n[64327];
assign t[64328] = t[64327] ^ n[64328];
assign t[64329] = t[64328] ^ n[64329];
assign t[64330] = t[64329] ^ n[64330];
assign t[64331] = t[64330] ^ n[64331];
assign t[64332] = t[64331] ^ n[64332];
assign t[64333] = t[64332] ^ n[64333];
assign t[64334] = t[64333] ^ n[64334];
assign t[64335] = t[64334] ^ n[64335];
assign t[64336] = t[64335] ^ n[64336];
assign t[64337] = t[64336] ^ n[64337];
assign t[64338] = t[64337] ^ n[64338];
assign t[64339] = t[64338] ^ n[64339];
assign t[64340] = t[64339] ^ n[64340];
assign t[64341] = t[64340] ^ n[64341];
assign t[64342] = t[64341] ^ n[64342];
assign t[64343] = t[64342] ^ n[64343];
assign t[64344] = t[64343] ^ n[64344];
assign t[64345] = t[64344] ^ n[64345];
assign t[64346] = t[64345] ^ n[64346];
assign t[64347] = t[64346] ^ n[64347];
assign t[64348] = t[64347] ^ n[64348];
assign t[64349] = t[64348] ^ n[64349];
assign t[64350] = t[64349] ^ n[64350];
assign t[64351] = t[64350] ^ n[64351];
assign t[64352] = t[64351] ^ n[64352];
assign t[64353] = t[64352] ^ n[64353];
assign t[64354] = t[64353] ^ n[64354];
assign t[64355] = t[64354] ^ n[64355];
assign t[64356] = t[64355] ^ n[64356];
assign t[64357] = t[64356] ^ n[64357];
assign t[64358] = t[64357] ^ n[64358];
assign t[64359] = t[64358] ^ n[64359];
assign t[64360] = t[64359] ^ n[64360];
assign t[64361] = t[64360] ^ n[64361];
assign t[64362] = t[64361] ^ n[64362];
assign t[64363] = t[64362] ^ n[64363];
assign t[64364] = t[64363] ^ n[64364];
assign t[64365] = t[64364] ^ n[64365];
assign t[64366] = t[64365] ^ n[64366];
assign t[64367] = t[64366] ^ n[64367];
assign t[64368] = t[64367] ^ n[64368];
assign t[64369] = t[64368] ^ n[64369];
assign t[64370] = t[64369] ^ n[64370];
assign t[64371] = t[64370] ^ n[64371];
assign t[64372] = t[64371] ^ n[64372];
assign t[64373] = t[64372] ^ n[64373];
assign t[64374] = t[64373] ^ n[64374];
assign t[64375] = t[64374] ^ n[64375];
assign t[64376] = t[64375] ^ n[64376];
assign t[64377] = t[64376] ^ n[64377];
assign t[64378] = t[64377] ^ n[64378];
assign t[64379] = t[64378] ^ n[64379];
assign t[64380] = t[64379] ^ n[64380];
assign t[64381] = t[64380] ^ n[64381];
assign t[64382] = t[64381] ^ n[64382];
assign t[64383] = t[64382] ^ n[64383];
assign t[64384] = t[64383] ^ n[64384];
assign t[64385] = t[64384] ^ n[64385];
assign t[64386] = t[64385] ^ n[64386];
assign t[64387] = t[64386] ^ n[64387];
assign t[64388] = t[64387] ^ n[64388];
assign t[64389] = t[64388] ^ n[64389];
assign t[64390] = t[64389] ^ n[64390];
assign t[64391] = t[64390] ^ n[64391];
assign t[64392] = t[64391] ^ n[64392];
assign t[64393] = t[64392] ^ n[64393];
assign t[64394] = t[64393] ^ n[64394];
assign t[64395] = t[64394] ^ n[64395];
assign t[64396] = t[64395] ^ n[64396];
assign t[64397] = t[64396] ^ n[64397];
assign t[64398] = t[64397] ^ n[64398];
assign t[64399] = t[64398] ^ n[64399];
assign t[64400] = t[64399] ^ n[64400];
assign t[64401] = t[64400] ^ n[64401];
assign t[64402] = t[64401] ^ n[64402];
assign t[64403] = t[64402] ^ n[64403];
assign t[64404] = t[64403] ^ n[64404];
assign t[64405] = t[64404] ^ n[64405];
assign t[64406] = t[64405] ^ n[64406];
assign t[64407] = t[64406] ^ n[64407];
assign t[64408] = t[64407] ^ n[64408];
assign t[64409] = t[64408] ^ n[64409];
assign t[64410] = t[64409] ^ n[64410];
assign t[64411] = t[64410] ^ n[64411];
assign t[64412] = t[64411] ^ n[64412];
assign t[64413] = t[64412] ^ n[64413];
assign t[64414] = t[64413] ^ n[64414];
assign t[64415] = t[64414] ^ n[64415];
assign t[64416] = t[64415] ^ n[64416];
assign t[64417] = t[64416] ^ n[64417];
assign t[64418] = t[64417] ^ n[64418];
assign t[64419] = t[64418] ^ n[64419];
assign t[64420] = t[64419] ^ n[64420];
assign t[64421] = t[64420] ^ n[64421];
assign t[64422] = t[64421] ^ n[64422];
assign t[64423] = t[64422] ^ n[64423];
assign t[64424] = t[64423] ^ n[64424];
assign t[64425] = t[64424] ^ n[64425];
assign t[64426] = t[64425] ^ n[64426];
assign t[64427] = t[64426] ^ n[64427];
assign t[64428] = t[64427] ^ n[64428];
assign t[64429] = t[64428] ^ n[64429];
assign t[64430] = t[64429] ^ n[64430];
assign t[64431] = t[64430] ^ n[64431];
assign t[64432] = t[64431] ^ n[64432];
assign t[64433] = t[64432] ^ n[64433];
assign t[64434] = t[64433] ^ n[64434];
assign t[64435] = t[64434] ^ n[64435];
assign t[64436] = t[64435] ^ n[64436];
assign t[64437] = t[64436] ^ n[64437];
assign t[64438] = t[64437] ^ n[64438];
assign t[64439] = t[64438] ^ n[64439];
assign t[64440] = t[64439] ^ n[64440];
assign t[64441] = t[64440] ^ n[64441];
assign t[64442] = t[64441] ^ n[64442];
assign t[64443] = t[64442] ^ n[64443];
assign t[64444] = t[64443] ^ n[64444];
assign t[64445] = t[64444] ^ n[64445];
assign t[64446] = t[64445] ^ n[64446];
assign t[64447] = t[64446] ^ n[64447];
assign t[64448] = t[64447] ^ n[64448];
assign t[64449] = t[64448] ^ n[64449];
assign t[64450] = t[64449] ^ n[64450];
assign t[64451] = t[64450] ^ n[64451];
assign t[64452] = t[64451] ^ n[64452];
assign t[64453] = t[64452] ^ n[64453];
assign t[64454] = t[64453] ^ n[64454];
assign t[64455] = t[64454] ^ n[64455];
assign t[64456] = t[64455] ^ n[64456];
assign t[64457] = t[64456] ^ n[64457];
assign t[64458] = t[64457] ^ n[64458];
assign t[64459] = t[64458] ^ n[64459];
assign t[64460] = t[64459] ^ n[64460];
assign t[64461] = t[64460] ^ n[64461];
assign t[64462] = t[64461] ^ n[64462];
assign t[64463] = t[64462] ^ n[64463];
assign t[64464] = t[64463] ^ n[64464];
assign t[64465] = t[64464] ^ n[64465];
assign t[64466] = t[64465] ^ n[64466];
assign t[64467] = t[64466] ^ n[64467];
assign t[64468] = t[64467] ^ n[64468];
assign t[64469] = t[64468] ^ n[64469];
assign t[64470] = t[64469] ^ n[64470];
assign t[64471] = t[64470] ^ n[64471];
assign t[64472] = t[64471] ^ n[64472];
assign t[64473] = t[64472] ^ n[64473];
assign t[64474] = t[64473] ^ n[64474];
assign t[64475] = t[64474] ^ n[64475];
assign t[64476] = t[64475] ^ n[64476];
assign t[64477] = t[64476] ^ n[64477];
assign t[64478] = t[64477] ^ n[64478];
assign t[64479] = t[64478] ^ n[64479];
assign t[64480] = t[64479] ^ n[64480];
assign t[64481] = t[64480] ^ n[64481];
assign t[64482] = t[64481] ^ n[64482];
assign t[64483] = t[64482] ^ n[64483];
assign t[64484] = t[64483] ^ n[64484];
assign t[64485] = t[64484] ^ n[64485];
assign t[64486] = t[64485] ^ n[64486];
assign t[64487] = t[64486] ^ n[64487];
assign t[64488] = t[64487] ^ n[64488];
assign t[64489] = t[64488] ^ n[64489];
assign t[64490] = t[64489] ^ n[64490];
assign t[64491] = t[64490] ^ n[64491];
assign t[64492] = t[64491] ^ n[64492];
assign t[64493] = t[64492] ^ n[64493];
assign t[64494] = t[64493] ^ n[64494];
assign t[64495] = t[64494] ^ n[64495];
assign t[64496] = t[64495] ^ n[64496];
assign t[64497] = t[64496] ^ n[64497];
assign t[64498] = t[64497] ^ n[64498];
assign t[64499] = t[64498] ^ n[64499];
assign t[64500] = t[64499] ^ n[64500];
assign t[64501] = t[64500] ^ n[64501];
assign t[64502] = t[64501] ^ n[64502];
assign t[64503] = t[64502] ^ n[64503];
assign t[64504] = t[64503] ^ n[64504];
assign t[64505] = t[64504] ^ n[64505];
assign t[64506] = t[64505] ^ n[64506];
assign t[64507] = t[64506] ^ n[64507];
assign t[64508] = t[64507] ^ n[64508];
assign t[64509] = t[64508] ^ n[64509];
assign t[64510] = t[64509] ^ n[64510];
assign t[64511] = t[64510] ^ n[64511];
assign t[64512] = t[64511] ^ n[64512];
assign t[64513] = t[64512] ^ n[64513];
assign t[64514] = t[64513] ^ n[64514];
assign t[64515] = t[64514] ^ n[64515];
assign t[64516] = t[64515] ^ n[64516];
assign t[64517] = t[64516] ^ n[64517];
assign t[64518] = t[64517] ^ n[64518];
assign t[64519] = t[64518] ^ n[64519];
assign t[64520] = t[64519] ^ n[64520];
assign t[64521] = t[64520] ^ n[64521];
assign t[64522] = t[64521] ^ n[64522];
assign t[64523] = t[64522] ^ n[64523];
assign t[64524] = t[64523] ^ n[64524];
assign t[64525] = t[64524] ^ n[64525];
assign t[64526] = t[64525] ^ n[64526];
assign t[64527] = t[64526] ^ n[64527];
assign t[64528] = t[64527] ^ n[64528];
assign t[64529] = t[64528] ^ n[64529];
assign t[64530] = t[64529] ^ n[64530];
assign t[64531] = t[64530] ^ n[64531];
assign t[64532] = t[64531] ^ n[64532];
assign t[64533] = t[64532] ^ n[64533];
assign t[64534] = t[64533] ^ n[64534];
assign t[64535] = t[64534] ^ n[64535];
assign t[64536] = t[64535] ^ n[64536];
assign t[64537] = t[64536] ^ n[64537];
assign t[64538] = t[64537] ^ n[64538];
assign t[64539] = t[64538] ^ n[64539];
assign t[64540] = t[64539] ^ n[64540];
assign t[64541] = t[64540] ^ n[64541];
assign t[64542] = t[64541] ^ n[64542];
assign t[64543] = t[64542] ^ n[64543];
assign t[64544] = t[64543] ^ n[64544];
assign t[64545] = t[64544] ^ n[64545];
assign t[64546] = t[64545] ^ n[64546];
assign t[64547] = t[64546] ^ n[64547];
assign t[64548] = t[64547] ^ n[64548];
assign t[64549] = t[64548] ^ n[64549];
assign t[64550] = t[64549] ^ n[64550];
assign t[64551] = t[64550] ^ n[64551];
assign t[64552] = t[64551] ^ n[64552];
assign t[64553] = t[64552] ^ n[64553];
assign t[64554] = t[64553] ^ n[64554];
assign t[64555] = t[64554] ^ n[64555];
assign t[64556] = t[64555] ^ n[64556];
assign t[64557] = t[64556] ^ n[64557];
assign t[64558] = t[64557] ^ n[64558];
assign t[64559] = t[64558] ^ n[64559];
assign t[64560] = t[64559] ^ n[64560];
assign t[64561] = t[64560] ^ n[64561];
assign t[64562] = t[64561] ^ n[64562];
assign t[64563] = t[64562] ^ n[64563];
assign t[64564] = t[64563] ^ n[64564];
assign t[64565] = t[64564] ^ n[64565];
assign t[64566] = t[64565] ^ n[64566];
assign t[64567] = t[64566] ^ n[64567];
assign t[64568] = t[64567] ^ n[64568];
assign t[64569] = t[64568] ^ n[64569];
assign t[64570] = t[64569] ^ n[64570];
assign t[64571] = t[64570] ^ n[64571];
assign t[64572] = t[64571] ^ n[64572];
assign t[64573] = t[64572] ^ n[64573];
assign t[64574] = t[64573] ^ n[64574];
assign t[64575] = t[64574] ^ n[64575];
assign t[64576] = t[64575] ^ n[64576];
assign t[64577] = t[64576] ^ n[64577];
assign t[64578] = t[64577] ^ n[64578];
assign t[64579] = t[64578] ^ n[64579];
assign t[64580] = t[64579] ^ n[64580];
assign t[64581] = t[64580] ^ n[64581];
assign t[64582] = t[64581] ^ n[64582];
assign t[64583] = t[64582] ^ n[64583];
assign t[64584] = t[64583] ^ n[64584];
assign t[64585] = t[64584] ^ n[64585];
assign t[64586] = t[64585] ^ n[64586];
assign t[64587] = t[64586] ^ n[64587];
assign t[64588] = t[64587] ^ n[64588];
assign t[64589] = t[64588] ^ n[64589];
assign t[64590] = t[64589] ^ n[64590];
assign t[64591] = t[64590] ^ n[64591];
assign t[64592] = t[64591] ^ n[64592];
assign t[64593] = t[64592] ^ n[64593];
assign t[64594] = t[64593] ^ n[64594];
assign t[64595] = t[64594] ^ n[64595];
assign t[64596] = t[64595] ^ n[64596];
assign t[64597] = t[64596] ^ n[64597];
assign t[64598] = t[64597] ^ n[64598];
assign t[64599] = t[64598] ^ n[64599];
assign t[64600] = t[64599] ^ n[64600];
assign t[64601] = t[64600] ^ n[64601];
assign t[64602] = t[64601] ^ n[64602];
assign t[64603] = t[64602] ^ n[64603];
assign t[64604] = t[64603] ^ n[64604];
assign t[64605] = t[64604] ^ n[64605];
assign t[64606] = t[64605] ^ n[64606];
assign t[64607] = t[64606] ^ n[64607];
assign t[64608] = t[64607] ^ n[64608];
assign t[64609] = t[64608] ^ n[64609];
assign t[64610] = t[64609] ^ n[64610];
assign t[64611] = t[64610] ^ n[64611];
assign t[64612] = t[64611] ^ n[64612];
assign t[64613] = t[64612] ^ n[64613];
assign t[64614] = t[64613] ^ n[64614];
assign t[64615] = t[64614] ^ n[64615];
assign t[64616] = t[64615] ^ n[64616];
assign t[64617] = t[64616] ^ n[64617];
assign t[64618] = t[64617] ^ n[64618];
assign t[64619] = t[64618] ^ n[64619];
assign t[64620] = t[64619] ^ n[64620];
assign t[64621] = t[64620] ^ n[64621];
assign t[64622] = t[64621] ^ n[64622];
assign t[64623] = t[64622] ^ n[64623];
assign t[64624] = t[64623] ^ n[64624];
assign t[64625] = t[64624] ^ n[64625];
assign t[64626] = t[64625] ^ n[64626];
assign t[64627] = t[64626] ^ n[64627];
assign t[64628] = t[64627] ^ n[64628];
assign t[64629] = t[64628] ^ n[64629];
assign t[64630] = t[64629] ^ n[64630];
assign t[64631] = t[64630] ^ n[64631];
assign t[64632] = t[64631] ^ n[64632];
assign t[64633] = t[64632] ^ n[64633];
assign t[64634] = t[64633] ^ n[64634];
assign t[64635] = t[64634] ^ n[64635];
assign t[64636] = t[64635] ^ n[64636];
assign t[64637] = t[64636] ^ n[64637];
assign t[64638] = t[64637] ^ n[64638];
assign t[64639] = t[64638] ^ n[64639];
assign t[64640] = t[64639] ^ n[64640];
assign t[64641] = t[64640] ^ n[64641];
assign t[64642] = t[64641] ^ n[64642];
assign t[64643] = t[64642] ^ n[64643];
assign t[64644] = t[64643] ^ n[64644];
assign t[64645] = t[64644] ^ n[64645];
assign t[64646] = t[64645] ^ n[64646];
assign t[64647] = t[64646] ^ n[64647];
assign t[64648] = t[64647] ^ n[64648];
assign t[64649] = t[64648] ^ n[64649];
assign t[64650] = t[64649] ^ n[64650];
assign t[64651] = t[64650] ^ n[64651];
assign t[64652] = t[64651] ^ n[64652];
assign t[64653] = t[64652] ^ n[64653];
assign t[64654] = t[64653] ^ n[64654];
assign t[64655] = t[64654] ^ n[64655];
assign t[64656] = t[64655] ^ n[64656];
assign t[64657] = t[64656] ^ n[64657];
assign t[64658] = t[64657] ^ n[64658];
assign t[64659] = t[64658] ^ n[64659];
assign t[64660] = t[64659] ^ n[64660];
assign t[64661] = t[64660] ^ n[64661];
assign t[64662] = t[64661] ^ n[64662];
assign t[64663] = t[64662] ^ n[64663];
assign t[64664] = t[64663] ^ n[64664];
assign t[64665] = t[64664] ^ n[64665];
assign t[64666] = t[64665] ^ n[64666];
assign t[64667] = t[64666] ^ n[64667];
assign t[64668] = t[64667] ^ n[64668];
assign t[64669] = t[64668] ^ n[64669];
assign t[64670] = t[64669] ^ n[64670];
assign t[64671] = t[64670] ^ n[64671];
assign t[64672] = t[64671] ^ n[64672];
assign t[64673] = t[64672] ^ n[64673];
assign t[64674] = t[64673] ^ n[64674];
assign t[64675] = t[64674] ^ n[64675];
assign t[64676] = t[64675] ^ n[64676];
assign t[64677] = t[64676] ^ n[64677];
assign t[64678] = t[64677] ^ n[64678];
assign t[64679] = t[64678] ^ n[64679];
assign t[64680] = t[64679] ^ n[64680];
assign t[64681] = t[64680] ^ n[64681];
assign t[64682] = t[64681] ^ n[64682];
assign t[64683] = t[64682] ^ n[64683];
assign t[64684] = t[64683] ^ n[64684];
assign t[64685] = t[64684] ^ n[64685];
assign t[64686] = t[64685] ^ n[64686];
assign t[64687] = t[64686] ^ n[64687];
assign t[64688] = t[64687] ^ n[64688];
assign t[64689] = t[64688] ^ n[64689];
assign t[64690] = t[64689] ^ n[64690];
assign t[64691] = t[64690] ^ n[64691];
assign t[64692] = t[64691] ^ n[64692];
assign t[64693] = t[64692] ^ n[64693];
assign t[64694] = t[64693] ^ n[64694];
assign t[64695] = t[64694] ^ n[64695];
assign t[64696] = t[64695] ^ n[64696];
assign t[64697] = t[64696] ^ n[64697];
assign t[64698] = t[64697] ^ n[64698];
assign t[64699] = t[64698] ^ n[64699];
assign t[64700] = t[64699] ^ n[64700];
assign t[64701] = t[64700] ^ n[64701];
assign t[64702] = t[64701] ^ n[64702];
assign t[64703] = t[64702] ^ n[64703];
assign t[64704] = t[64703] ^ n[64704];
assign t[64705] = t[64704] ^ n[64705];
assign t[64706] = t[64705] ^ n[64706];
assign t[64707] = t[64706] ^ n[64707];
assign t[64708] = t[64707] ^ n[64708];
assign t[64709] = t[64708] ^ n[64709];
assign t[64710] = t[64709] ^ n[64710];
assign t[64711] = t[64710] ^ n[64711];
assign t[64712] = t[64711] ^ n[64712];
assign t[64713] = t[64712] ^ n[64713];
assign t[64714] = t[64713] ^ n[64714];
assign t[64715] = t[64714] ^ n[64715];
assign t[64716] = t[64715] ^ n[64716];
assign t[64717] = t[64716] ^ n[64717];
assign t[64718] = t[64717] ^ n[64718];
assign t[64719] = t[64718] ^ n[64719];
assign t[64720] = t[64719] ^ n[64720];
assign t[64721] = t[64720] ^ n[64721];
assign t[64722] = t[64721] ^ n[64722];
assign t[64723] = t[64722] ^ n[64723];
assign t[64724] = t[64723] ^ n[64724];
assign t[64725] = t[64724] ^ n[64725];
assign t[64726] = t[64725] ^ n[64726];
assign t[64727] = t[64726] ^ n[64727];
assign t[64728] = t[64727] ^ n[64728];
assign t[64729] = t[64728] ^ n[64729];
assign t[64730] = t[64729] ^ n[64730];
assign t[64731] = t[64730] ^ n[64731];
assign t[64732] = t[64731] ^ n[64732];
assign t[64733] = t[64732] ^ n[64733];
assign t[64734] = t[64733] ^ n[64734];
assign t[64735] = t[64734] ^ n[64735];
assign t[64736] = t[64735] ^ n[64736];
assign t[64737] = t[64736] ^ n[64737];
assign t[64738] = t[64737] ^ n[64738];
assign t[64739] = t[64738] ^ n[64739];
assign t[64740] = t[64739] ^ n[64740];
assign t[64741] = t[64740] ^ n[64741];
assign t[64742] = t[64741] ^ n[64742];
assign t[64743] = t[64742] ^ n[64743];
assign t[64744] = t[64743] ^ n[64744];
assign t[64745] = t[64744] ^ n[64745];
assign t[64746] = t[64745] ^ n[64746];
assign t[64747] = t[64746] ^ n[64747];
assign t[64748] = t[64747] ^ n[64748];
assign t[64749] = t[64748] ^ n[64749];
assign t[64750] = t[64749] ^ n[64750];
assign t[64751] = t[64750] ^ n[64751];
assign t[64752] = t[64751] ^ n[64752];
assign t[64753] = t[64752] ^ n[64753];
assign t[64754] = t[64753] ^ n[64754];
assign t[64755] = t[64754] ^ n[64755];
assign t[64756] = t[64755] ^ n[64756];
assign t[64757] = t[64756] ^ n[64757];
assign t[64758] = t[64757] ^ n[64758];
assign t[64759] = t[64758] ^ n[64759];
assign t[64760] = t[64759] ^ n[64760];
assign t[64761] = t[64760] ^ n[64761];
assign t[64762] = t[64761] ^ n[64762];
assign t[64763] = t[64762] ^ n[64763];
assign t[64764] = t[64763] ^ n[64764];
assign t[64765] = t[64764] ^ n[64765];
assign t[64766] = t[64765] ^ n[64766];
assign t[64767] = t[64766] ^ n[64767];
assign t[64768] = t[64767] ^ n[64768];
assign t[64769] = t[64768] ^ n[64769];
assign t[64770] = t[64769] ^ n[64770];
assign t[64771] = t[64770] ^ n[64771];
assign t[64772] = t[64771] ^ n[64772];
assign t[64773] = t[64772] ^ n[64773];
assign t[64774] = t[64773] ^ n[64774];
assign t[64775] = t[64774] ^ n[64775];
assign t[64776] = t[64775] ^ n[64776];
assign t[64777] = t[64776] ^ n[64777];
assign t[64778] = t[64777] ^ n[64778];
assign t[64779] = t[64778] ^ n[64779];
assign t[64780] = t[64779] ^ n[64780];
assign t[64781] = t[64780] ^ n[64781];
assign t[64782] = t[64781] ^ n[64782];
assign t[64783] = t[64782] ^ n[64783];
assign t[64784] = t[64783] ^ n[64784];
assign t[64785] = t[64784] ^ n[64785];
assign t[64786] = t[64785] ^ n[64786];
assign t[64787] = t[64786] ^ n[64787];
assign t[64788] = t[64787] ^ n[64788];
assign t[64789] = t[64788] ^ n[64789];
assign t[64790] = t[64789] ^ n[64790];
assign t[64791] = t[64790] ^ n[64791];
assign t[64792] = t[64791] ^ n[64792];
assign t[64793] = t[64792] ^ n[64793];
assign t[64794] = t[64793] ^ n[64794];
assign t[64795] = t[64794] ^ n[64795];
assign t[64796] = t[64795] ^ n[64796];
assign t[64797] = t[64796] ^ n[64797];
assign t[64798] = t[64797] ^ n[64798];
assign t[64799] = t[64798] ^ n[64799];
assign t[64800] = t[64799] ^ n[64800];
assign t[64801] = t[64800] ^ n[64801];
assign t[64802] = t[64801] ^ n[64802];
assign t[64803] = t[64802] ^ n[64803];
assign t[64804] = t[64803] ^ n[64804];
assign t[64805] = t[64804] ^ n[64805];
assign t[64806] = t[64805] ^ n[64806];
assign t[64807] = t[64806] ^ n[64807];
assign t[64808] = t[64807] ^ n[64808];
assign t[64809] = t[64808] ^ n[64809];
assign t[64810] = t[64809] ^ n[64810];
assign t[64811] = t[64810] ^ n[64811];
assign t[64812] = t[64811] ^ n[64812];
assign t[64813] = t[64812] ^ n[64813];
assign t[64814] = t[64813] ^ n[64814];
assign t[64815] = t[64814] ^ n[64815];
assign t[64816] = t[64815] ^ n[64816];
assign t[64817] = t[64816] ^ n[64817];
assign t[64818] = t[64817] ^ n[64818];
assign t[64819] = t[64818] ^ n[64819];
assign t[64820] = t[64819] ^ n[64820];
assign t[64821] = t[64820] ^ n[64821];
assign t[64822] = t[64821] ^ n[64822];
assign t[64823] = t[64822] ^ n[64823];
assign t[64824] = t[64823] ^ n[64824];
assign t[64825] = t[64824] ^ n[64825];
assign t[64826] = t[64825] ^ n[64826];
assign t[64827] = t[64826] ^ n[64827];
assign t[64828] = t[64827] ^ n[64828];
assign t[64829] = t[64828] ^ n[64829];
assign t[64830] = t[64829] ^ n[64830];
assign t[64831] = t[64830] ^ n[64831];
assign t[64832] = t[64831] ^ n[64832];
assign t[64833] = t[64832] ^ n[64833];
assign t[64834] = t[64833] ^ n[64834];
assign t[64835] = t[64834] ^ n[64835];
assign t[64836] = t[64835] ^ n[64836];
assign t[64837] = t[64836] ^ n[64837];
assign t[64838] = t[64837] ^ n[64838];
assign t[64839] = t[64838] ^ n[64839];
assign t[64840] = t[64839] ^ n[64840];
assign t[64841] = t[64840] ^ n[64841];
assign t[64842] = t[64841] ^ n[64842];
assign t[64843] = t[64842] ^ n[64843];
assign t[64844] = t[64843] ^ n[64844];
assign t[64845] = t[64844] ^ n[64845];
assign t[64846] = t[64845] ^ n[64846];
assign t[64847] = t[64846] ^ n[64847];
assign t[64848] = t[64847] ^ n[64848];
assign t[64849] = t[64848] ^ n[64849];
assign t[64850] = t[64849] ^ n[64850];
assign t[64851] = t[64850] ^ n[64851];
assign t[64852] = t[64851] ^ n[64852];
assign t[64853] = t[64852] ^ n[64853];
assign t[64854] = t[64853] ^ n[64854];
assign t[64855] = t[64854] ^ n[64855];
assign t[64856] = t[64855] ^ n[64856];
assign t[64857] = t[64856] ^ n[64857];
assign t[64858] = t[64857] ^ n[64858];
assign t[64859] = t[64858] ^ n[64859];
assign t[64860] = t[64859] ^ n[64860];
assign t[64861] = t[64860] ^ n[64861];
assign t[64862] = t[64861] ^ n[64862];
assign t[64863] = t[64862] ^ n[64863];
assign t[64864] = t[64863] ^ n[64864];
assign t[64865] = t[64864] ^ n[64865];
assign t[64866] = t[64865] ^ n[64866];
assign t[64867] = t[64866] ^ n[64867];
assign t[64868] = t[64867] ^ n[64868];
assign t[64869] = t[64868] ^ n[64869];
assign t[64870] = t[64869] ^ n[64870];
assign t[64871] = t[64870] ^ n[64871];
assign t[64872] = t[64871] ^ n[64872];
assign t[64873] = t[64872] ^ n[64873];
assign t[64874] = t[64873] ^ n[64874];
assign t[64875] = t[64874] ^ n[64875];
assign t[64876] = t[64875] ^ n[64876];
assign t[64877] = t[64876] ^ n[64877];
assign t[64878] = t[64877] ^ n[64878];
assign t[64879] = t[64878] ^ n[64879];
assign t[64880] = t[64879] ^ n[64880];
assign t[64881] = t[64880] ^ n[64881];
assign t[64882] = t[64881] ^ n[64882];
assign t[64883] = t[64882] ^ n[64883];
assign t[64884] = t[64883] ^ n[64884];
assign t[64885] = t[64884] ^ n[64885];
assign t[64886] = t[64885] ^ n[64886];
assign t[64887] = t[64886] ^ n[64887];
assign t[64888] = t[64887] ^ n[64888];
assign t[64889] = t[64888] ^ n[64889];
assign t[64890] = t[64889] ^ n[64890];
assign t[64891] = t[64890] ^ n[64891];
assign t[64892] = t[64891] ^ n[64892];
assign t[64893] = t[64892] ^ n[64893];
assign t[64894] = t[64893] ^ n[64894];
assign t[64895] = t[64894] ^ n[64895];
assign t[64896] = t[64895] ^ n[64896];
assign t[64897] = t[64896] ^ n[64897];
assign t[64898] = t[64897] ^ n[64898];
assign t[64899] = t[64898] ^ n[64899];
assign t[64900] = t[64899] ^ n[64900];
assign t[64901] = t[64900] ^ n[64901];
assign t[64902] = t[64901] ^ n[64902];
assign t[64903] = t[64902] ^ n[64903];
assign t[64904] = t[64903] ^ n[64904];
assign t[64905] = t[64904] ^ n[64905];
assign t[64906] = t[64905] ^ n[64906];
assign t[64907] = t[64906] ^ n[64907];
assign t[64908] = t[64907] ^ n[64908];
assign t[64909] = t[64908] ^ n[64909];
assign t[64910] = t[64909] ^ n[64910];
assign t[64911] = t[64910] ^ n[64911];
assign t[64912] = t[64911] ^ n[64912];
assign t[64913] = t[64912] ^ n[64913];
assign t[64914] = t[64913] ^ n[64914];
assign t[64915] = t[64914] ^ n[64915];
assign t[64916] = t[64915] ^ n[64916];
assign t[64917] = t[64916] ^ n[64917];
assign t[64918] = t[64917] ^ n[64918];
assign t[64919] = t[64918] ^ n[64919];
assign t[64920] = t[64919] ^ n[64920];
assign t[64921] = t[64920] ^ n[64921];
assign t[64922] = t[64921] ^ n[64922];
assign t[64923] = t[64922] ^ n[64923];
assign t[64924] = t[64923] ^ n[64924];
assign t[64925] = t[64924] ^ n[64925];
assign t[64926] = t[64925] ^ n[64926];
assign t[64927] = t[64926] ^ n[64927];
assign t[64928] = t[64927] ^ n[64928];
assign t[64929] = t[64928] ^ n[64929];
assign t[64930] = t[64929] ^ n[64930];
assign t[64931] = t[64930] ^ n[64931];
assign t[64932] = t[64931] ^ n[64932];
assign t[64933] = t[64932] ^ n[64933];
assign t[64934] = t[64933] ^ n[64934];
assign t[64935] = t[64934] ^ n[64935];
assign t[64936] = t[64935] ^ n[64936];
assign t[64937] = t[64936] ^ n[64937];
assign t[64938] = t[64937] ^ n[64938];
assign t[64939] = t[64938] ^ n[64939];
assign t[64940] = t[64939] ^ n[64940];
assign t[64941] = t[64940] ^ n[64941];
assign t[64942] = t[64941] ^ n[64942];
assign t[64943] = t[64942] ^ n[64943];
assign t[64944] = t[64943] ^ n[64944];
assign t[64945] = t[64944] ^ n[64945];
assign t[64946] = t[64945] ^ n[64946];
assign t[64947] = t[64946] ^ n[64947];
assign t[64948] = t[64947] ^ n[64948];
assign t[64949] = t[64948] ^ n[64949];
assign t[64950] = t[64949] ^ n[64950];
assign t[64951] = t[64950] ^ n[64951];
assign t[64952] = t[64951] ^ n[64952];
assign t[64953] = t[64952] ^ n[64953];
assign t[64954] = t[64953] ^ n[64954];
assign t[64955] = t[64954] ^ n[64955];
assign t[64956] = t[64955] ^ n[64956];
assign t[64957] = t[64956] ^ n[64957];
assign t[64958] = t[64957] ^ n[64958];
assign t[64959] = t[64958] ^ n[64959];
assign t[64960] = t[64959] ^ n[64960];
assign t[64961] = t[64960] ^ n[64961];
assign t[64962] = t[64961] ^ n[64962];
assign t[64963] = t[64962] ^ n[64963];
assign t[64964] = t[64963] ^ n[64964];
assign t[64965] = t[64964] ^ n[64965];
assign t[64966] = t[64965] ^ n[64966];
assign t[64967] = t[64966] ^ n[64967];
assign t[64968] = t[64967] ^ n[64968];
assign t[64969] = t[64968] ^ n[64969];
assign t[64970] = t[64969] ^ n[64970];
assign t[64971] = t[64970] ^ n[64971];
assign t[64972] = t[64971] ^ n[64972];
assign t[64973] = t[64972] ^ n[64973];
assign t[64974] = t[64973] ^ n[64974];
assign t[64975] = t[64974] ^ n[64975];
assign t[64976] = t[64975] ^ n[64976];
assign t[64977] = t[64976] ^ n[64977];
assign t[64978] = t[64977] ^ n[64978];
assign t[64979] = t[64978] ^ n[64979];
assign t[64980] = t[64979] ^ n[64980];
assign t[64981] = t[64980] ^ n[64981];
assign t[64982] = t[64981] ^ n[64982];
assign t[64983] = t[64982] ^ n[64983];
assign t[64984] = t[64983] ^ n[64984];
assign t[64985] = t[64984] ^ n[64985];
assign t[64986] = t[64985] ^ n[64986];
assign t[64987] = t[64986] ^ n[64987];
assign t[64988] = t[64987] ^ n[64988];
assign t[64989] = t[64988] ^ n[64989];
assign t[64990] = t[64989] ^ n[64990];
assign t[64991] = t[64990] ^ n[64991];
assign t[64992] = t[64991] ^ n[64992];
assign t[64993] = t[64992] ^ n[64993];
assign t[64994] = t[64993] ^ n[64994];
assign t[64995] = t[64994] ^ n[64995];
assign t[64996] = t[64995] ^ n[64996];
assign t[64997] = t[64996] ^ n[64997];
assign t[64998] = t[64997] ^ n[64998];
assign t[64999] = t[64998] ^ n[64999];
assign t[65000] = t[64999] ^ n[65000];
assign t[65001] = t[65000] ^ n[65001];
assign t[65002] = t[65001] ^ n[65002];
assign t[65003] = t[65002] ^ n[65003];
assign t[65004] = t[65003] ^ n[65004];
assign t[65005] = t[65004] ^ n[65005];
assign t[65006] = t[65005] ^ n[65006];
assign t[65007] = t[65006] ^ n[65007];
assign t[65008] = t[65007] ^ n[65008];
assign t[65009] = t[65008] ^ n[65009];
assign t[65010] = t[65009] ^ n[65010];
assign t[65011] = t[65010] ^ n[65011];
assign t[65012] = t[65011] ^ n[65012];
assign t[65013] = t[65012] ^ n[65013];
assign t[65014] = t[65013] ^ n[65014];
assign t[65015] = t[65014] ^ n[65015];
assign t[65016] = t[65015] ^ n[65016];
assign t[65017] = t[65016] ^ n[65017];
assign t[65018] = t[65017] ^ n[65018];
assign t[65019] = t[65018] ^ n[65019];
assign t[65020] = t[65019] ^ n[65020];
assign t[65021] = t[65020] ^ n[65021];
assign t[65022] = t[65021] ^ n[65022];
assign t[65023] = t[65022] ^ n[65023];
assign t[65024] = t[65023] ^ n[65024];
assign t[65025] = t[65024] ^ n[65025];
assign t[65026] = t[65025] ^ n[65026];
assign t[65027] = t[65026] ^ n[65027];
assign t[65028] = t[65027] ^ n[65028];
assign t[65029] = t[65028] ^ n[65029];
assign t[65030] = t[65029] ^ n[65030];
assign t[65031] = t[65030] ^ n[65031];
assign t[65032] = t[65031] ^ n[65032];
assign t[65033] = t[65032] ^ n[65033];
assign t[65034] = t[65033] ^ n[65034];
assign t[65035] = t[65034] ^ n[65035];
assign t[65036] = t[65035] ^ n[65036];
assign t[65037] = t[65036] ^ n[65037];
assign t[65038] = t[65037] ^ n[65038];
assign t[65039] = t[65038] ^ n[65039];
assign t[65040] = t[65039] ^ n[65040];
assign t[65041] = t[65040] ^ n[65041];
assign t[65042] = t[65041] ^ n[65042];
assign t[65043] = t[65042] ^ n[65043];
assign t[65044] = t[65043] ^ n[65044];
assign t[65045] = t[65044] ^ n[65045];
assign t[65046] = t[65045] ^ n[65046];
assign t[65047] = t[65046] ^ n[65047];
assign t[65048] = t[65047] ^ n[65048];
assign t[65049] = t[65048] ^ n[65049];
assign t[65050] = t[65049] ^ n[65050];
assign t[65051] = t[65050] ^ n[65051];
assign t[65052] = t[65051] ^ n[65052];
assign t[65053] = t[65052] ^ n[65053];
assign t[65054] = t[65053] ^ n[65054];
assign t[65055] = t[65054] ^ n[65055];
assign t[65056] = t[65055] ^ n[65056];
assign t[65057] = t[65056] ^ n[65057];
assign t[65058] = t[65057] ^ n[65058];
assign t[65059] = t[65058] ^ n[65059];
assign t[65060] = t[65059] ^ n[65060];
assign t[65061] = t[65060] ^ n[65061];
assign t[65062] = t[65061] ^ n[65062];
assign t[65063] = t[65062] ^ n[65063];
assign t[65064] = t[65063] ^ n[65064];
assign t[65065] = t[65064] ^ n[65065];
assign t[65066] = t[65065] ^ n[65066];
assign t[65067] = t[65066] ^ n[65067];
assign t[65068] = t[65067] ^ n[65068];
assign t[65069] = t[65068] ^ n[65069];
assign t[65070] = t[65069] ^ n[65070];
assign t[65071] = t[65070] ^ n[65071];
assign t[65072] = t[65071] ^ n[65072];
assign t[65073] = t[65072] ^ n[65073];
assign t[65074] = t[65073] ^ n[65074];
assign t[65075] = t[65074] ^ n[65075];
assign t[65076] = t[65075] ^ n[65076];
assign t[65077] = t[65076] ^ n[65077];
assign t[65078] = t[65077] ^ n[65078];
assign t[65079] = t[65078] ^ n[65079];
assign t[65080] = t[65079] ^ n[65080];
assign t[65081] = t[65080] ^ n[65081];
assign t[65082] = t[65081] ^ n[65082];
assign t[65083] = t[65082] ^ n[65083];
assign t[65084] = t[65083] ^ n[65084];
assign t[65085] = t[65084] ^ n[65085];
assign t[65086] = t[65085] ^ n[65086];
assign t[65087] = t[65086] ^ n[65087];
assign t[65088] = t[65087] ^ n[65088];
assign t[65089] = t[65088] ^ n[65089];
assign t[65090] = t[65089] ^ n[65090];
assign t[65091] = t[65090] ^ n[65091];
assign t[65092] = t[65091] ^ n[65092];
assign t[65093] = t[65092] ^ n[65093];
assign t[65094] = t[65093] ^ n[65094];
assign t[65095] = t[65094] ^ n[65095];
assign t[65096] = t[65095] ^ n[65096];
assign t[65097] = t[65096] ^ n[65097];
assign t[65098] = t[65097] ^ n[65098];
assign t[65099] = t[65098] ^ n[65099];
assign t[65100] = t[65099] ^ n[65100];
assign t[65101] = t[65100] ^ n[65101];
assign t[65102] = t[65101] ^ n[65102];
assign t[65103] = t[65102] ^ n[65103];
assign t[65104] = t[65103] ^ n[65104];
assign t[65105] = t[65104] ^ n[65105];
assign t[65106] = t[65105] ^ n[65106];
assign t[65107] = t[65106] ^ n[65107];
assign t[65108] = t[65107] ^ n[65108];
assign t[65109] = t[65108] ^ n[65109];
assign t[65110] = t[65109] ^ n[65110];
assign t[65111] = t[65110] ^ n[65111];
assign t[65112] = t[65111] ^ n[65112];
assign t[65113] = t[65112] ^ n[65113];
assign t[65114] = t[65113] ^ n[65114];
assign t[65115] = t[65114] ^ n[65115];
assign t[65116] = t[65115] ^ n[65116];
assign t[65117] = t[65116] ^ n[65117];
assign t[65118] = t[65117] ^ n[65118];
assign t[65119] = t[65118] ^ n[65119];
assign t[65120] = t[65119] ^ n[65120];
assign t[65121] = t[65120] ^ n[65121];
assign t[65122] = t[65121] ^ n[65122];
assign t[65123] = t[65122] ^ n[65123];
assign t[65124] = t[65123] ^ n[65124];
assign t[65125] = t[65124] ^ n[65125];
assign t[65126] = t[65125] ^ n[65126];
assign t[65127] = t[65126] ^ n[65127];
assign t[65128] = t[65127] ^ n[65128];
assign t[65129] = t[65128] ^ n[65129];
assign t[65130] = t[65129] ^ n[65130];
assign t[65131] = t[65130] ^ n[65131];
assign t[65132] = t[65131] ^ n[65132];
assign t[65133] = t[65132] ^ n[65133];
assign t[65134] = t[65133] ^ n[65134];
assign t[65135] = t[65134] ^ n[65135];
assign t[65136] = t[65135] ^ n[65136];
assign t[65137] = t[65136] ^ n[65137];
assign t[65138] = t[65137] ^ n[65138];
assign t[65139] = t[65138] ^ n[65139];
assign t[65140] = t[65139] ^ n[65140];
assign t[65141] = t[65140] ^ n[65141];
assign t[65142] = t[65141] ^ n[65142];
assign t[65143] = t[65142] ^ n[65143];
assign t[65144] = t[65143] ^ n[65144];
assign t[65145] = t[65144] ^ n[65145];
assign t[65146] = t[65145] ^ n[65146];
assign t[65147] = t[65146] ^ n[65147];
assign t[65148] = t[65147] ^ n[65148];
assign t[65149] = t[65148] ^ n[65149];
assign t[65150] = t[65149] ^ n[65150];
assign t[65151] = t[65150] ^ n[65151];
assign t[65152] = t[65151] ^ n[65152];
assign t[65153] = t[65152] ^ n[65153];
assign t[65154] = t[65153] ^ n[65154];
assign t[65155] = t[65154] ^ n[65155];
assign t[65156] = t[65155] ^ n[65156];
assign t[65157] = t[65156] ^ n[65157];
assign t[65158] = t[65157] ^ n[65158];
assign t[65159] = t[65158] ^ n[65159];
assign t[65160] = t[65159] ^ n[65160];
assign t[65161] = t[65160] ^ n[65161];
assign t[65162] = t[65161] ^ n[65162];
assign t[65163] = t[65162] ^ n[65163];
assign t[65164] = t[65163] ^ n[65164];
assign t[65165] = t[65164] ^ n[65165];
assign t[65166] = t[65165] ^ n[65166];
assign t[65167] = t[65166] ^ n[65167];
assign t[65168] = t[65167] ^ n[65168];
assign t[65169] = t[65168] ^ n[65169];
assign t[65170] = t[65169] ^ n[65170];
assign t[65171] = t[65170] ^ n[65171];
assign t[65172] = t[65171] ^ n[65172];
assign t[65173] = t[65172] ^ n[65173];
assign t[65174] = t[65173] ^ n[65174];
assign t[65175] = t[65174] ^ n[65175];
assign t[65176] = t[65175] ^ n[65176];
assign t[65177] = t[65176] ^ n[65177];
assign t[65178] = t[65177] ^ n[65178];
assign t[65179] = t[65178] ^ n[65179];
assign t[65180] = t[65179] ^ n[65180];
assign t[65181] = t[65180] ^ n[65181];
assign t[65182] = t[65181] ^ n[65182];
assign t[65183] = t[65182] ^ n[65183];
assign t[65184] = t[65183] ^ n[65184];
assign t[65185] = t[65184] ^ n[65185];
assign t[65186] = t[65185] ^ n[65186];
assign t[65187] = t[65186] ^ n[65187];
assign t[65188] = t[65187] ^ n[65188];
assign t[65189] = t[65188] ^ n[65189];
assign t[65190] = t[65189] ^ n[65190];
assign t[65191] = t[65190] ^ n[65191];
assign t[65192] = t[65191] ^ n[65192];
assign t[65193] = t[65192] ^ n[65193];
assign t[65194] = t[65193] ^ n[65194];
assign t[65195] = t[65194] ^ n[65195];
assign t[65196] = t[65195] ^ n[65196];
assign t[65197] = t[65196] ^ n[65197];
assign t[65198] = t[65197] ^ n[65198];
assign t[65199] = t[65198] ^ n[65199];
assign t[65200] = t[65199] ^ n[65200];
assign t[65201] = t[65200] ^ n[65201];
assign t[65202] = t[65201] ^ n[65202];
assign t[65203] = t[65202] ^ n[65203];
assign t[65204] = t[65203] ^ n[65204];
assign t[65205] = t[65204] ^ n[65205];
assign t[65206] = t[65205] ^ n[65206];
assign t[65207] = t[65206] ^ n[65207];
assign t[65208] = t[65207] ^ n[65208];
assign t[65209] = t[65208] ^ n[65209];
assign t[65210] = t[65209] ^ n[65210];
assign t[65211] = t[65210] ^ n[65211];
assign t[65212] = t[65211] ^ n[65212];
assign t[65213] = t[65212] ^ n[65213];
assign t[65214] = t[65213] ^ n[65214];
assign t[65215] = t[65214] ^ n[65215];
assign t[65216] = t[65215] ^ n[65216];
assign t[65217] = t[65216] ^ n[65217];
assign t[65218] = t[65217] ^ n[65218];
assign t[65219] = t[65218] ^ n[65219];
assign t[65220] = t[65219] ^ n[65220];
assign t[65221] = t[65220] ^ n[65221];
assign t[65222] = t[65221] ^ n[65222];
assign t[65223] = t[65222] ^ n[65223];
assign t[65224] = t[65223] ^ n[65224];
assign t[65225] = t[65224] ^ n[65225];
assign t[65226] = t[65225] ^ n[65226];
assign t[65227] = t[65226] ^ n[65227];
assign t[65228] = t[65227] ^ n[65228];
assign t[65229] = t[65228] ^ n[65229];
assign t[65230] = t[65229] ^ n[65230];
assign t[65231] = t[65230] ^ n[65231];
assign t[65232] = t[65231] ^ n[65232];
assign t[65233] = t[65232] ^ n[65233];
assign t[65234] = t[65233] ^ n[65234];
assign t[65235] = t[65234] ^ n[65235];
assign t[65236] = t[65235] ^ n[65236];
assign t[65237] = t[65236] ^ n[65237];
assign t[65238] = t[65237] ^ n[65238];
assign t[65239] = t[65238] ^ n[65239];
assign t[65240] = t[65239] ^ n[65240];
assign t[65241] = t[65240] ^ n[65241];
assign t[65242] = t[65241] ^ n[65242];
assign t[65243] = t[65242] ^ n[65243];
assign t[65244] = t[65243] ^ n[65244];
assign t[65245] = t[65244] ^ n[65245];
assign t[65246] = t[65245] ^ n[65246];
assign t[65247] = t[65246] ^ n[65247];
assign t[65248] = t[65247] ^ n[65248];
assign t[65249] = t[65248] ^ n[65249];
assign t[65250] = t[65249] ^ n[65250];
assign t[65251] = t[65250] ^ n[65251];
assign t[65252] = t[65251] ^ n[65252];
assign t[65253] = t[65252] ^ n[65253];
assign t[65254] = t[65253] ^ n[65254];
assign t[65255] = t[65254] ^ n[65255];
assign t[65256] = t[65255] ^ n[65256];
assign t[65257] = t[65256] ^ n[65257];
assign t[65258] = t[65257] ^ n[65258];
assign t[65259] = t[65258] ^ n[65259];
assign t[65260] = t[65259] ^ n[65260];
assign t[65261] = t[65260] ^ n[65261];
assign t[65262] = t[65261] ^ n[65262];
assign t[65263] = t[65262] ^ n[65263];
assign t[65264] = t[65263] ^ n[65264];
assign t[65265] = t[65264] ^ n[65265];
assign t[65266] = t[65265] ^ n[65266];
assign t[65267] = t[65266] ^ n[65267];
assign t[65268] = t[65267] ^ n[65268];
assign t[65269] = t[65268] ^ n[65269];
assign t[65270] = t[65269] ^ n[65270];
assign t[65271] = t[65270] ^ n[65271];
assign t[65272] = t[65271] ^ n[65272];
assign t[65273] = t[65272] ^ n[65273];
assign t[65274] = t[65273] ^ n[65274];
assign t[65275] = t[65274] ^ n[65275];
assign t[65276] = t[65275] ^ n[65276];
assign t[65277] = t[65276] ^ n[65277];
assign t[65278] = t[65277] ^ n[65278];
assign t[65279] = t[65278] ^ n[65279];
assign t[65280] = t[65279] ^ n[65280];
assign t[65281] = t[65280] ^ n[65281];
assign t[65282] = t[65281] ^ n[65282];
assign t[65283] = t[65282] ^ n[65283];
assign t[65284] = t[65283] ^ n[65284];
assign t[65285] = t[65284] ^ n[65285];
assign t[65286] = t[65285] ^ n[65286];
assign t[65287] = t[65286] ^ n[65287];
assign t[65288] = t[65287] ^ n[65288];
assign t[65289] = t[65288] ^ n[65289];
assign t[65290] = t[65289] ^ n[65290];
assign t[65291] = t[65290] ^ n[65291];
assign t[65292] = t[65291] ^ n[65292];
assign t[65293] = t[65292] ^ n[65293];
assign t[65294] = t[65293] ^ n[65294];
assign t[65295] = t[65294] ^ n[65295];
assign t[65296] = t[65295] ^ n[65296];
assign t[65297] = t[65296] ^ n[65297];
assign t[65298] = t[65297] ^ n[65298];
assign t[65299] = t[65298] ^ n[65299];
assign t[65300] = t[65299] ^ n[65300];
assign t[65301] = t[65300] ^ n[65301];
assign t[65302] = t[65301] ^ n[65302];
assign t[65303] = t[65302] ^ n[65303];
assign t[65304] = t[65303] ^ n[65304];
assign t[65305] = t[65304] ^ n[65305];
assign t[65306] = t[65305] ^ n[65306];
assign t[65307] = t[65306] ^ n[65307];
assign t[65308] = t[65307] ^ n[65308];
assign t[65309] = t[65308] ^ n[65309];
assign t[65310] = t[65309] ^ n[65310];
assign t[65311] = t[65310] ^ n[65311];
assign t[65312] = t[65311] ^ n[65312];
assign t[65313] = t[65312] ^ n[65313];
assign t[65314] = t[65313] ^ n[65314];
assign t[65315] = t[65314] ^ n[65315];
assign t[65316] = t[65315] ^ n[65316];
assign t[65317] = t[65316] ^ n[65317];
assign t[65318] = t[65317] ^ n[65318];
assign t[65319] = t[65318] ^ n[65319];
assign t[65320] = t[65319] ^ n[65320];
assign t[65321] = t[65320] ^ n[65321];
assign t[65322] = t[65321] ^ n[65322];
assign t[65323] = t[65322] ^ n[65323];
assign t[65324] = t[65323] ^ n[65324];
assign t[65325] = t[65324] ^ n[65325];
assign t[65326] = t[65325] ^ n[65326];
assign t[65327] = t[65326] ^ n[65327];
assign t[65328] = t[65327] ^ n[65328];
assign t[65329] = t[65328] ^ n[65329];
assign t[65330] = t[65329] ^ n[65330];
assign t[65331] = t[65330] ^ n[65331];
assign t[65332] = t[65331] ^ n[65332];
assign t[65333] = t[65332] ^ n[65333];
assign t[65334] = t[65333] ^ n[65334];
assign t[65335] = t[65334] ^ n[65335];
assign t[65336] = t[65335] ^ n[65336];
assign t[65337] = t[65336] ^ n[65337];
assign t[65338] = t[65337] ^ n[65338];
assign t[65339] = t[65338] ^ n[65339];
assign t[65340] = t[65339] ^ n[65340];
assign t[65341] = t[65340] ^ n[65341];
assign t[65342] = t[65341] ^ n[65342];
assign t[65343] = t[65342] ^ n[65343];
assign t[65344] = t[65343] ^ n[65344];
assign t[65345] = t[65344] ^ n[65345];
assign t[65346] = t[65345] ^ n[65346];
assign t[65347] = t[65346] ^ n[65347];
assign t[65348] = t[65347] ^ n[65348];
assign t[65349] = t[65348] ^ n[65349];
assign t[65350] = t[65349] ^ n[65350];
assign t[65351] = t[65350] ^ n[65351];
assign t[65352] = t[65351] ^ n[65352];
assign t[65353] = t[65352] ^ n[65353];
assign t[65354] = t[65353] ^ n[65354];
assign t[65355] = t[65354] ^ n[65355];
assign t[65356] = t[65355] ^ n[65356];
assign t[65357] = t[65356] ^ n[65357];
assign t[65358] = t[65357] ^ n[65358];
assign t[65359] = t[65358] ^ n[65359];
assign t[65360] = t[65359] ^ n[65360];
assign t[65361] = t[65360] ^ n[65361];
assign t[65362] = t[65361] ^ n[65362];
assign t[65363] = t[65362] ^ n[65363];
assign t[65364] = t[65363] ^ n[65364];
assign t[65365] = t[65364] ^ n[65365];
assign t[65366] = t[65365] ^ n[65366];
assign t[65367] = t[65366] ^ n[65367];
assign t[65368] = t[65367] ^ n[65368];
assign t[65369] = t[65368] ^ n[65369];
assign t[65370] = t[65369] ^ n[65370];
assign t[65371] = t[65370] ^ n[65371];
assign t[65372] = t[65371] ^ n[65372];
assign t[65373] = t[65372] ^ n[65373];
assign t[65374] = t[65373] ^ n[65374];
assign t[65375] = t[65374] ^ n[65375];
assign t[65376] = t[65375] ^ n[65376];
assign t[65377] = t[65376] ^ n[65377];
assign t[65378] = t[65377] ^ n[65378];
assign t[65379] = t[65378] ^ n[65379];
assign t[65380] = t[65379] ^ n[65380];
assign t[65381] = t[65380] ^ n[65381];
assign t[65382] = t[65381] ^ n[65382];
assign t[65383] = t[65382] ^ n[65383];
assign t[65384] = t[65383] ^ n[65384];
assign t[65385] = t[65384] ^ n[65385];
assign t[65386] = t[65385] ^ n[65386];
assign t[65387] = t[65386] ^ n[65387];
assign t[65388] = t[65387] ^ n[65388];
assign t[65389] = t[65388] ^ n[65389];
assign t[65390] = t[65389] ^ n[65390];
assign t[65391] = t[65390] ^ n[65391];
assign t[65392] = t[65391] ^ n[65392];
assign t[65393] = t[65392] ^ n[65393];
assign t[65394] = t[65393] ^ n[65394];
assign t[65395] = t[65394] ^ n[65395];
assign t[65396] = t[65395] ^ n[65396];
assign t[65397] = t[65396] ^ n[65397];
assign t[65398] = t[65397] ^ n[65398];
assign t[65399] = t[65398] ^ n[65399];
assign t[65400] = t[65399] ^ n[65400];
assign t[65401] = t[65400] ^ n[65401];
assign t[65402] = t[65401] ^ n[65402];
assign t[65403] = t[65402] ^ n[65403];
assign t[65404] = t[65403] ^ n[65404];
assign t[65405] = t[65404] ^ n[65405];
assign t[65406] = t[65405] ^ n[65406];
assign t[65407] = t[65406] ^ n[65407];
assign t[65408] = t[65407] ^ n[65408];
assign t[65409] = t[65408] ^ n[65409];
assign t[65410] = t[65409] ^ n[65410];
assign t[65411] = t[65410] ^ n[65411];
assign t[65412] = t[65411] ^ n[65412];
assign t[65413] = t[65412] ^ n[65413];
assign t[65414] = t[65413] ^ n[65414];
assign t[65415] = t[65414] ^ n[65415];
assign t[65416] = t[65415] ^ n[65416];
assign t[65417] = t[65416] ^ n[65417];
assign t[65418] = t[65417] ^ n[65418];
assign t[65419] = t[65418] ^ n[65419];
assign t[65420] = t[65419] ^ n[65420];
assign t[65421] = t[65420] ^ n[65421];
assign t[65422] = t[65421] ^ n[65422];
assign t[65423] = t[65422] ^ n[65423];
assign t[65424] = t[65423] ^ n[65424];
assign t[65425] = t[65424] ^ n[65425];
assign t[65426] = t[65425] ^ n[65426];
assign t[65427] = t[65426] ^ n[65427];
assign t[65428] = t[65427] ^ n[65428];
assign t[65429] = t[65428] ^ n[65429];
assign t[65430] = t[65429] ^ n[65430];
assign t[65431] = t[65430] ^ n[65431];
assign t[65432] = t[65431] ^ n[65432];
assign t[65433] = t[65432] ^ n[65433];
assign t[65434] = t[65433] ^ n[65434];
assign t[65435] = t[65434] ^ n[65435];
assign t[65436] = t[65435] ^ n[65436];
assign t[65437] = t[65436] ^ n[65437];
assign t[65438] = t[65437] ^ n[65438];
assign t[65439] = t[65438] ^ n[65439];
assign t[65440] = t[65439] ^ n[65440];
assign t[65441] = t[65440] ^ n[65441];
assign t[65442] = t[65441] ^ n[65442];
assign t[65443] = t[65442] ^ n[65443];
assign t[65444] = t[65443] ^ n[65444];
assign t[65445] = t[65444] ^ n[65445];
assign t[65446] = t[65445] ^ n[65446];
assign t[65447] = t[65446] ^ n[65447];
assign t[65448] = t[65447] ^ n[65448];
assign t[65449] = t[65448] ^ n[65449];
assign t[65450] = t[65449] ^ n[65450];
assign t[65451] = t[65450] ^ n[65451];
assign t[65452] = t[65451] ^ n[65452];
assign t[65453] = t[65452] ^ n[65453];
assign t[65454] = t[65453] ^ n[65454];
assign t[65455] = t[65454] ^ n[65455];
assign t[65456] = t[65455] ^ n[65456];
assign t[65457] = t[65456] ^ n[65457];
assign t[65458] = t[65457] ^ n[65458];
assign t[65459] = t[65458] ^ n[65459];
assign t[65460] = t[65459] ^ n[65460];
assign t[65461] = t[65460] ^ n[65461];
assign t[65462] = t[65461] ^ n[65462];
assign t[65463] = t[65462] ^ n[65463];
assign t[65464] = t[65463] ^ n[65464];
assign t[65465] = t[65464] ^ n[65465];
assign t[65466] = t[65465] ^ n[65466];
assign t[65467] = t[65466] ^ n[65467];
assign t[65468] = t[65467] ^ n[65468];
assign t[65469] = t[65468] ^ n[65469];
assign t[65470] = t[65469] ^ n[65470];
assign t[65471] = t[65470] ^ n[65471];
assign t[65472] = t[65471] ^ n[65472];
assign t[65473] = t[65472] ^ n[65473];
assign t[65474] = t[65473] ^ n[65474];
assign t[65475] = t[65474] ^ n[65475];
assign t[65476] = t[65475] ^ n[65476];
assign t[65477] = t[65476] ^ n[65477];
assign t[65478] = t[65477] ^ n[65478];
assign t[65479] = t[65478] ^ n[65479];
assign t[65480] = t[65479] ^ n[65480];
assign t[65481] = t[65480] ^ n[65481];
assign t[65482] = t[65481] ^ n[65482];
assign t[65483] = t[65482] ^ n[65483];
assign t[65484] = t[65483] ^ n[65484];
assign t[65485] = t[65484] ^ n[65485];
assign t[65486] = t[65485] ^ n[65486];
assign t[65487] = t[65486] ^ n[65487];
assign t[65488] = t[65487] ^ n[65488];
assign t[65489] = t[65488] ^ n[65489];
assign t[65490] = t[65489] ^ n[65490];
assign t[65491] = t[65490] ^ n[65491];
assign t[65492] = t[65491] ^ n[65492];
assign t[65493] = t[65492] ^ n[65493];
assign t[65494] = t[65493] ^ n[65494];
assign t[65495] = t[65494] ^ n[65495];
assign t[65496] = t[65495] ^ n[65496];
assign t[65497] = t[65496] ^ n[65497];
assign t[65498] = t[65497] ^ n[65498];
assign t[65499] = t[65498] ^ n[65499];
assign t[65500] = t[65499] ^ n[65500];
assign t[65501] = t[65500] ^ n[65501];
assign t[65502] = t[65501] ^ n[65502];
assign t[65503] = t[65502] ^ n[65503];
assign t[65504] = t[65503] ^ n[65504];
assign t[65505] = t[65504] ^ n[65505];
assign t[65506] = t[65505] ^ n[65506];
assign t[65507] = t[65506] ^ n[65507];
assign t[65508] = t[65507] ^ n[65508];
assign t[65509] = t[65508] ^ n[65509];
assign t[65510] = t[65509] ^ n[65510];
assign t[65511] = t[65510] ^ n[65511];
assign t[65512] = t[65511] ^ n[65512];
assign t[65513] = t[65512] ^ n[65513];
assign t[65514] = t[65513] ^ n[65514];
assign t[65515] = t[65514] ^ n[65515];
assign t[65516] = t[65515] ^ n[65516];
assign t[65517] = t[65516] ^ n[65517];
assign t[65518] = t[65517] ^ n[65518];

//asigning bit 15
assign s[15] = ( a[15] ^ b [15] ) ^ t[65518];

endmodule