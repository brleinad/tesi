module lut(index, lut_out);

input [7:0] index;
output [7:0] lut_out;

reg [7:0] lut_out;//[255:0]; //LUlut_out
always @(index)
begin
        case(index)
                0   : lut_out = 251; 
                1   : lut_out = 175; 
                2   : lut_out = 119; 
                3   : lut_out = 215; 
                4   : lut_out = 81; 
                5   : lut_out = 14; 
                6   : lut_out = 79; 
                7   : lut_out = 191; 
                8   : lut_out = 103; 
                9   : lut_out = 49; 
                10  : lut_out = 181; 
                11  : lut_out = 143; 
                12  : lut_out = 186; 
                13  : lut_out = 157; 
                14  : lut_out = 0;
                15  : lut_out = 232; 
                16  : lut_out = 31; 
                17  : lut_out = 32; 
                18  : lut_out = 55; 
                19  : lut_out = 60; 
                20  : lut_out = 152; 
                21  : lut_out = 58; 
                22  : lut_out = 17; 
                23  : lut_out = 237; 
                24  : lut_out = 174; 
                25  : lut_out = 70; 
                26  : lut_out = 160; 
                27  : lut_out = 144; 
                28  : lut_out = 220; 
                29  : lut_out = 90; 
                30  : lut_out = 57;
                31  : lut_out = 223; 
                32  : lut_out = 59;  
                33  : lut_out = 3; 
                34  : lut_out = 18; 
                35  : lut_out = 140; 
                36  : lut_out = 111; 
                37  : lut_out = 166; 
                38  : lut_out = 203; 
                39  : lut_out = 196; 
                40  : lut_out = 134; 
                41  : lut_out = 243; 
                42  : lut_out = 124; 
                43  : lut_out = 95; 
                44  : lut_out = 222; 
                45  : lut_out = 179;
                46  : lut_out = 197; 
                47  : lut_out = 65; 
                48  : lut_out = 180; 
                49  : lut_out = 48; 
                50  : lut_out = 36; 
                51  : lut_out = 15; 
                52  : lut_out = 107; 
                53  : lut_out = 46; 
                54  : lut_out = 233; 
                55  : lut_out = 130; 
                56  : lut_out = 165; 
                57  : lut_out = 30; 
                58  : lut_out = 123; 
                59  : lut_out = 161; 
                60  : lut_out = 209; 
                61  : lut_out = 23;
                62  : lut_out = 97; 
                63  : lut_out = 16; 
                64  : lut_out = 40; 
                65  : lut_out = 91; 
                66  : lut_out = 219; 
                67  : lut_out = 61; 
                68  : lut_out = 100; 
                69  : lut_out = 10; 
                70  : lut_out = 210; 
                71  : lut_out = 109; 
                72  : lut_out = 250; 
                73  : lut_out = 127; 
                74  : lut_out = 22; 
                75  : lut_out = 138; 
                76  : lut_out = 29; 
                77  : lut_out = 108;
                78  : lut_out = 244; 
                79  : lut_out = 67; 
                80  : lut_out = 207; 
                81  : lut_out = 9; 
                82  : lut_out = 178; 
                83  : lut_out = 204; 
                84  : lut_out = 74; 
                85  : lut_out = 98; 
                86  : lut_out = 126; 
                87  : lut_out = 249; 
                88  : lut_out = 167; 
                89  : lut_out = 116; 
                90  : lut_out = 34; 
                91  : lut_out = 77; 
                92  : lut_out = 193;
                93  : lut_out = 200; 
                94  : lut_out = 121; 
                95  : lut_out = 5; 
                96  : lut_out = 20; 
                97  : lut_out = 113; 
                98  : lut_out = 71; 
                99  : lut_out = 35; 
                100 : lut_out = 128; 
                101 : lut_out = 13; 
                102 : lut_out = 182; 
                103 : lut_out = 94; 
                104 : lut_out = 25; 
                105 : lut_out = 226; 
                106 : lut_out = 227; 
                107 : lut_out = 199; 
                108 : lut_out = 75;
                109 : lut_out = 27; 
                110 : lut_out = 41; 
                111 : lut_out = 245; 
                112 : lut_out = 230; 
                113 : lut_out = 224; 
                114 : lut_out = 43; 
                115 : lut_out = 225; 
                116 : lut_out = 177; 
                117 : lut_out = 26; 
                118 : lut_out = 155; 
                119 : lut_out = 150; 
                120 : lut_out = 212; 
                121 : lut_out = 142; 
                122 : lut_out = 218; 
                123 : lut_out = 115;
                124 : lut_out = 241; 
                125 : lut_out = 73; 
                126 : lut_out = 88; 
                127 : lut_out = 105; 
                128 : lut_out = 39; 
                129 : lut_out = 114; 
                130 : lut_out = 62; 
                131 : lut_out = 255; 
                132 : lut_out = 192; 
                133 : lut_out = 201; 
                134 : lut_out = 145; 
                135 : lut_out = 214; 
                136 : lut_out = 168; 
                137 : lut_out = 158; 
                138 : lut_out = 221;
                139 : lut_out = 148; 
                140 : lut_out = 154; 
                141 : lut_out = 122; 
                142 : lut_out = 12; 
                143 : lut_out = 84; 
                144 : lut_out = 82; 
                145 : lut_out = 163; 
                146 : lut_out = 44; 
                147 : lut_out = 139; 
                148 : lut_out = 228; 
                149 : lut_out = 236; 
                150 : lut_out = 205; 
                151 : lut_out = 242; 
                152 : lut_out = 217; 
                153 : lut_out = 11;
                154 : lut_out = 187; 
                155 : lut_out = 146; 
                156 : lut_out = 159; 
                157 : lut_out = 64; 
                158 : lut_out = 86; 
                159 : lut_out = 239; 
                160 : lut_out = 195; 
                161 : lut_out = 42; 
                162 : lut_out = 106; 
                163 : lut_out = 198; 
                164 : lut_out = 118; 
                165 : lut_out = 112; 
                166 : lut_out = 184; 
                167 : lut_out = 172; 
                168 : lut_out = 87;
                169 : lut_out = 2; 
                170 : lut_out = 173; 
                171 : lut_out = 117; 
                172 : lut_out = 176; 
                173 : lut_out = 229; 
                174 : lut_out = 247; 
                175 : lut_out = 253; 
                176 : lut_out = 137; 
                177 : lut_out = 185; 
                178 : lut_out = 99; 
                179 : lut_out = 164; 
                180 : lut_out = 102; 
                181 : lut_out = 147; 
                182 : lut_out = 45; 
                183 : lut_out = 66;
                184 : lut_out = 231; 
                185 : lut_out = 52; 
                186 : lut_out = 141; 
                187 : lut_out = 211; 
                188 : lut_out = 194; 
                189 : lut_out = 206; 
                190 : lut_out = 246; 
                191 : lut_out = 238; 
                192 : lut_out = 56; 
                193 : lut_out = 110; 
                194 : lut_out = 78; 
                195 : lut_out = 248; 
                196 : lut_out = 63; 
                197 : lut_out = 240; 
                198 : lut_out = 189;
                199 : lut_out = 93; 
                200 : lut_out = 92; 
                201 : lut_out = 51; 
                202 : lut_out = 53; 
                203 : lut_out = 183; 
                204 : lut_out = 19; 
                205 : lut_out = 171; 
                206 : lut_out = 72; 
                207 : lut_out = 50; 
                208 : lut_out = 33; 
                209 : lut_out = 104; 
                210 : lut_out = 101; 
                211 : lut_out = 69; 
                212 : lut_out = 8; 
                213 : lut_out = 252; 
                214 : lut_out = 83; 
                215 : lut_out = 120;
                216 : lut_out = 76; 
                217 : lut_out = 135; 
                218 : lut_out = 85; 
                219 : lut_out = 54; 
                220 : lut_out = 202; 
                221 : lut_out = 125; 
                222 : lut_out = 188; 
                223 : lut_out = 213; 
                224 : lut_out = 96; 
                225 : lut_out = 235; 
                226 : lut_out = 136; 
                227 : lut_out = 208; 
                228 : lut_out = 162; 
                229 : lut_out = 129; 
                230 : lut_out = 190;
                231 : lut_out = 132; 
                232 : lut_out = 156; 
                233 : lut_out = 38; 
                234 : lut_out = 47; 
                235 : lut_out = 1; 
                236 : lut_out = 7; 
                237 : lut_out = 254; 
                238 : lut_out = 24; 
                239 : lut_out = 4; 
                240 : lut_out = 216; 
                241 : lut_out = 131; 
                242 : lut_out = 89; 
                243 : lut_out = 21; 
                244 : lut_out = 28; 
                245 : lut_out = 133; 
                246 : lut_out = 37; 
                247 : lut_out = 153;
                248 : lut_out = 149; 
                249 : lut_out = 80; 
                250 : lut_out = 170; 
                251 : lut_out = 68; 
                252 : lut_out = 6; 
                253 : lut_out = 169; 
                254 : lut_out = 234; 
                255 : lut_out = 151;
                default: lut_out = 0;
    endcase
end

endmodule
