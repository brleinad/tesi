module adder4bit.out(a__0, a__1, a__2, a__3,b__0, b__1, b__2, b__3,s__0, s__1, s__2, s__3);
  input a__0, a__1, a__2, a__3;
  input b__0, b__1, b__2, b__3;
  output s__0, s__1, s__2, s__3;
  wire   n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign s__3 = n14 ^ n15;
  assign n15 = n16 | n17;
  assign n17 = a__2 & n18;
  assign n16 = b__2 & n19;
  assign n19 = a__2 | n18;
  assign n14 = b__3 ^ a__3;
  assign s__2 = n20 ^ n18;
  assign n18 = n21 | n22;
  assign n22 = b__1 & a__1;
  assign n21 = n23 & b__0;
  assign n23 = a__0 & n24;
  assign n24 = a__1 | b__1;
  assign n20 = b__2 ^ a__2;
  assign s__1 = n25 ^ n26;
  assign n26 = b__1 ^ a__1;
  assign n25 = b__0 & a__0;
  assign s__0 = b__0 ^ a__0;
