
module cla_adder ( a, b, s, cin, cout );
  input [63:0] a;
  input [63:0] b;
  output [63:0] s;
  input cin;
  output cout;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62;
  wire   [62:0] g;
  wire   [63:0] p;
  wire   [63:1] c;

  XOR2D0 C578 ( .A1(p[0]), .A2(cin), .Z(s[0]) );
  XOR2D0 C577 ( .A1(p[1]), .A2(c[1]), .Z(s[1]) );
  XOR2D0 C576 ( .A1(p[2]), .A2(c[2]), .Z(s[2]) );
  XOR2D0 C575 ( .A1(p[3]), .A2(c[3]), .Z(s[3]) );
  XOR2D0 C574 ( .A1(p[4]), .A2(c[4]), .Z(s[4]) );
  XOR2D0 C573 ( .A1(p[5]), .A2(c[5]), .Z(s[5]) );
  XOR2D0 C572 ( .A1(p[6]), .A2(c[6]), .Z(s[6]) );
  XOR2D0 C571 ( .A1(p[7]), .A2(c[7]), .Z(s[7]) );
  XOR2D0 C570 ( .A1(p[8]), .A2(c[8]), .Z(s[8]) );
  XOR2D0 C569 ( .A1(p[9]), .A2(c[9]), .Z(s[9]) );
  XOR2D0 C568 ( .A1(p[10]), .A2(c[10]), .Z(s[10]) );
  XOR2D0 C567 ( .A1(p[11]), .A2(c[11]), .Z(s[11]) );
  XOR2D0 C566 ( .A1(p[12]), .A2(c[12]), .Z(s[12]) );
  XOR2D0 C565 ( .A1(p[13]), .A2(c[13]), .Z(s[13]) );
  XOR2D0 C564 ( .A1(p[14]), .A2(c[14]), .Z(s[14]) );
  XOR2D0 C563 ( .A1(p[15]), .A2(c[15]), .Z(s[15]) );
  XOR2D0 C562 ( .A1(p[16]), .A2(c[16]), .Z(s[16]) );
  XOR2D0 C561 ( .A1(p[17]), .A2(c[17]), .Z(s[17]) );
  XOR2D0 C560 ( .A1(p[18]), .A2(c[18]), .Z(s[18]) );
  XOR2D0 C559 ( .A1(p[19]), .A2(c[19]), .Z(s[19]) );
  XOR2D0 C558 ( .A1(p[20]), .A2(c[20]), .Z(s[20]) );
  XOR2D0 C557 ( .A1(p[21]), .A2(c[21]), .Z(s[21]) );
  XOR2D0 C556 ( .A1(p[22]), .A2(c[22]), .Z(s[22]) );
  XOR2D0 C555 ( .A1(p[23]), .A2(c[23]), .Z(s[23]) );
  XOR2D0 C554 ( .A1(p[24]), .A2(c[24]), .Z(s[24]) );
  XOR2D0 C553 ( .A1(p[25]), .A2(c[25]), .Z(s[25]) );
  XOR2D0 C552 ( .A1(p[26]), .A2(c[26]), .Z(s[26]) );
  XOR2D0 C551 ( .A1(p[27]), .A2(c[27]), .Z(s[27]) );
  XOR2D0 C550 ( .A1(p[28]), .A2(c[28]), .Z(s[28]) );
  XOR2D0 C549 ( .A1(p[29]), .A2(c[29]), .Z(s[29]) );
  XOR2D0 C548 ( .A1(p[30]), .A2(c[30]), .Z(s[30]) );
  XOR2D0 C547 ( .A1(p[31]), .A2(c[31]), .Z(s[31]) );
  XOR2D0 C546 ( .A1(p[32]), .A2(c[32]), .Z(s[32]) );
  XOR2D0 C545 ( .A1(p[33]), .A2(c[33]), .Z(s[33]) );
  XOR2D0 C544 ( .A1(p[34]), .A2(c[34]), .Z(s[34]) );
  XOR2D0 C543 ( .A1(p[35]), .A2(c[35]), .Z(s[35]) );
  XOR2D0 C542 ( .A1(p[36]), .A2(c[36]), .Z(s[36]) );
  XOR2D0 C541 ( .A1(p[37]), .A2(c[37]), .Z(s[37]) );
  XOR2D0 C540 ( .A1(p[38]), .A2(c[38]), .Z(s[38]) );
  XOR2D0 C539 ( .A1(p[39]), .A2(c[39]), .Z(s[39]) );
  XOR2D0 C538 ( .A1(p[40]), .A2(c[40]), .Z(s[40]) );
  XOR2D0 C537 ( .A1(p[41]), .A2(c[41]), .Z(s[41]) );
  XOR2D0 C536 ( .A1(p[42]), .A2(c[42]), .Z(s[42]) );
  XOR2D0 C535 ( .A1(p[43]), .A2(c[43]), .Z(s[43]) );
  XOR2D0 C534 ( .A1(p[44]), .A2(c[44]), .Z(s[44]) );
  XOR2D0 C533 ( .A1(p[45]), .A2(c[45]), .Z(s[45]) );
  XOR2D0 C532 ( .A1(p[46]), .A2(c[46]), .Z(s[46]) );
  XOR2D0 C531 ( .A1(p[47]), .A2(c[47]), .Z(s[47]) );
  XOR2D0 C530 ( .A1(p[48]), .A2(c[48]), .Z(s[48]) );
  XOR2D0 C529 ( .A1(p[49]), .A2(c[49]), .Z(s[49]) );
  XOR2D0 C528 ( .A1(p[50]), .A2(c[50]), .Z(s[50]) );
  XOR2D0 C527 ( .A1(p[51]), .A2(c[51]), .Z(s[51]) );
  XOR2D0 C526 ( .A1(p[52]), .A2(c[52]), .Z(s[52]) );
  XOR2D0 C525 ( .A1(p[53]), .A2(c[53]), .Z(s[53]) );
  XOR2D0 C524 ( .A1(p[54]), .A2(c[54]), .Z(s[54]) );
  XOR2D0 C523 ( .A1(p[55]), .A2(c[55]), .Z(s[55]) );
  XOR2D0 C522 ( .A1(p[56]), .A2(c[56]), .Z(s[56]) );
  XOR2D0 C521 ( .A1(p[57]), .A2(c[57]), .Z(s[57]) );
  XOR2D0 C520 ( .A1(p[58]), .A2(c[58]), .Z(s[58]) );
  XOR2D0 C519 ( .A1(p[59]), .A2(c[59]), .Z(s[59]) );
  XOR2D0 C518 ( .A1(p[60]), .A2(c[60]), .Z(s[60]) );
  XOR2D0 C517 ( .A1(p[61]), .A2(c[61]), .Z(s[61]) );
  XOR2D0 C516 ( .A1(p[62]), .A2(c[62]), .Z(s[62]) );
  XOR2D0 C515 ( .A1(p[63]), .A2(c[63]), .Z(s[63]) );
  AN2D0 C514 ( .A1(p[62]), .A2(c[62]), .Z(N62) );
  OR2D0 C513 ( .A1(g[62]), .A2(N62), .Z(c[63]) );
  AN2D0 C512 ( .A1(p[61]), .A2(c[61]), .Z(N61) );
  OR2D0 C511 ( .A1(g[61]), .A2(N61), .Z(c[62]) );
  AN2D0 C510 ( .A1(p[60]), .A2(c[60]), .Z(N60) );
  OR2D0 C509 ( .A1(g[60]), .A2(N60), .Z(c[61]) );
  AN2D0 C508 ( .A1(p[59]), .A2(c[59]), .Z(N59) );
  OR2D0 C507 ( .A1(g[59]), .A2(N59), .Z(c[60]) );
  AN2D0 C506 ( .A1(p[58]), .A2(c[58]), .Z(N58) );
  OR2D0 C505 ( .A1(g[58]), .A2(N58), .Z(c[59]) );
  AN2D0 C504 ( .A1(p[57]), .A2(c[57]), .Z(N57) );
  OR2D0 C503 ( .A1(g[57]), .A2(N57), .Z(c[58]) );
  AN2D0 C502 ( .A1(p[56]), .A2(c[56]), .Z(N56) );
  OR2D0 C501 ( .A1(g[56]), .A2(N56), .Z(c[57]) );
  AN2D0 C500 ( .A1(p[55]), .A2(c[55]), .Z(N55) );
  OR2D0 C499 ( .A1(g[55]), .A2(N55), .Z(c[56]) );
  AN2D0 C498 ( .A1(p[54]), .A2(c[54]), .Z(N54) );
  OR2D0 C497 ( .A1(g[54]), .A2(N54), .Z(c[55]) );
  AN2D0 C496 ( .A1(p[53]), .A2(c[53]), .Z(N53) );
  OR2D0 C495 ( .A1(g[53]), .A2(N53), .Z(c[54]) );
  AN2D0 C494 ( .A1(p[52]), .A2(c[52]), .Z(N52) );
  OR2D0 C493 ( .A1(g[52]), .A2(N52), .Z(c[53]) );
  AN2D0 C492 ( .A1(p[51]), .A2(c[51]), .Z(N51) );
  OR2D0 C491 ( .A1(g[51]), .A2(N51), .Z(c[52]) );
  AN2D0 C490 ( .A1(p[50]), .A2(c[50]), .Z(N50) );
  OR2D0 C489 ( .A1(g[50]), .A2(N50), .Z(c[51]) );
  AN2D0 C488 ( .A1(p[49]), .A2(c[49]), .Z(N49) );
  OR2D0 C487 ( .A1(g[49]), .A2(N49), .Z(c[50]) );
  AN2D0 C486 ( .A1(p[48]), .A2(c[48]), .Z(N48) );
  OR2D0 C485 ( .A1(g[48]), .A2(N48), .Z(c[49]) );
  AN2D0 C484 ( .A1(p[47]), .A2(c[47]), .Z(N47) );
  OR2D0 C483 ( .A1(g[47]), .A2(N47), .Z(c[48]) );
  AN2D0 C482 ( .A1(p[46]), .A2(c[46]), .Z(N46) );
  OR2D0 C481 ( .A1(g[46]), .A2(N46), .Z(c[47]) );
  AN2D0 C480 ( .A1(p[45]), .A2(c[45]), .Z(N45) );
  OR2D0 C479 ( .A1(g[45]), .A2(N45), .Z(c[46]) );
  AN2D0 C478 ( .A1(p[44]), .A2(c[44]), .Z(N44) );
  OR2D0 C477 ( .A1(g[44]), .A2(N44), .Z(c[45]) );
  AN2D0 C476 ( .A1(p[43]), .A2(c[43]), .Z(N43) );
  OR2D0 C475 ( .A1(g[43]), .A2(N43), .Z(c[44]) );
  AN2D0 C474 ( .A1(p[42]), .A2(c[42]), .Z(N42) );
  OR2D0 C473 ( .A1(g[42]), .A2(N42), .Z(c[43]) );
  AN2D0 C472 ( .A1(p[41]), .A2(c[41]), .Z(N41) );
  OR2D0 C471 ( .A1(g[41]), .A2(N41), .Z(c[42]) );
  AN2D0 C470 ( .A1(p[40]), .A2(c[40]), .Z(N40) );
  OR2D0 C469 ( .A1(g[40]), .A2(N40), .Z(c[41]) );
  AN2D0 C468 ( .A1(p[39]), .A2(c[39]), .Z(N39) );
  OR2D0 C467 ( .A1(g[39]), .A2(N39), .Z(c[40]) );
  AN2D0 C466 ( .A1(p[38]), .A2(c[38]), .Z(N38) );
  OR2D0 C465 ( .A1(g[38]), .A2(N38), .Z(c[39]) );
  AN2D0 C464 ( .A1(p[37]), .A2(c[37]), .Z(N37) );
  OR2D0 C463 ( .A1(g[37]), .A2(N37), .Z(c[38]) );
  AN2D0 C462 ( .A1(p[36]), .A2(c[36]), .Z(N36) );
  OR2D0 C461 ( .A1(g[36]), .A2(N36), .Z(c[37]) );
  AN2D0 C460 ( .A1(p[35]), .A2(c[35]), .Z(N35) );
  OR2D0 C459 ( .A1(g[35]), .A2(N35), .Z(c[36]) );
  AN2D0 C458 ( .A1(p[34]), .A2(c[34]), .Z(N34) );
  OR2D0 C457 ( .A1(g[34]), .A2(N34), .Z(c[35]) );
  AN2D0 C456 ( .A1(p[33]), .A2(c[33]), .Z(N33) );
  OR2D0 C455 ( .A1(g[33]), .A2(N33), .Z(c[34]) );
  AN2D0 C454 ( .A1(p[32]), .A2(c[32]), .Z(N32) );
  OR2D0 C453 ( .A1(g[32]), .A2(N32), .Z(c[33]) );
  AN2D0 C452 ( .A1(p[31]), .A2(c[31]), .Z(N31) );
  OR2D0 C451 ( .A1(g[31]), .A2(N31), .Z(c[32]) );
  AN2D0 C450 ( .A1(p[30]), .A2(c[30]), .Z(N30) );
  OR2D0 C449 ( .A1(g[30]), .A2(N30), .Z(c[31]) );
  AN2D0 C448 ( .A1(p[29]), .A2(c[29]), .Z(N29) );
  OR2D0 C447 ( .A1(g[29]), .A2(N29), .Z(c[30]) );
  AN2D0 C446 ( .A1(p[28]), .A2(c[28]), .Z(N28) );
  OR2D0 C445 ( .A1(g[28]), .A2(N28), .Z(c[29]) );
  AN2D0 C444 ( .A1(p[27]), .A2(c[27]), .Z(N27) );
  OR2D0 C443 ( .A1(g[27]), .A2(N27), .Z(c[28]) );
  AN2D0 C442 ( .A1(p[26]), .A2(c[26]), .Z(N26) );
  OR2D0 C441 ( .A1(g[26]), .A2(N26), .Z(c[27]) );
  AN2D0 C440 ( .A1(p[25]), .A2(c[25]), .Z(N25) );
  OR2D0 C439 ( .A1(g[25]), .A2(N25), .Z(c[26]) );
  AN2D0 C438 ( .A1(p[24]), .A2(c[24]), .Z(N24) );
  OR2D0 C437 ( .A1(g[24]), .A2(N24), .Z(c[25]) );
  AN2D0 C436 ( .A1(p[23]), .A2(c[23]), .Z(N23) );
  OR2D0 C435 ( .A1(g[23]), .A2(N23), .Z(c[24]) );
  AN2D0 C434 ( .A1(p[22]), .A2(c[22]), .Z(N22) );
  OR2D0 C433 ( .A1(g[22]), .A2(N22), .Z(c[23]) );
  AN2D0 C432 ( .A1(p[21]), .A2(c[21]), .Z(N21) );
  OR2D0 C431 ( .A1(g[21]), .A2(N21), .Z(c[22]) );
  AN2D0 C430 ( .A1(p[20]), .A2(c[20]), .Z(N20) );
  OR2D0 C429 ( .A1(g[20]), .A2(N20), .Z(c[21]) );
  AN2D0 C428 ( .A1(p[19]), .A2(c[19]), .Z(N19) );
  OR2D0 C427 ( .A1(g[19]), .A2(N19), .Z(c[20]) );
  AN2D0 C426 ( .A1(p[18]), .A2(c[18]), .Z(N18) );
  OR2D0 C425 ( .A1(g[18]), .A2(N18), .Z(c[19]) );
  AN2D0 C424 ( .A1(p[17]), .A2(c[17]), .Z(N17) );
  OR2D0 C423 ( .A1(g[17]), .A2(N17), .Z(c[18]) );
  AN2D0 C422 ( .A1(p[16]), .A2(c[16]), .Z(N16) );
  OR2D0 C421 ( .A1(g[16]), .A2(N16), .Z(c[17]) );
  AN2D0 C420 ( .A1(p[15]), .A2(c[15]), .Z(N15) );
  OR2D0 C419 ( .A1(g[15]), .A2(N15), .Z(c[16]) );
  AN2D0 C418 ( .A1(p[14]), .A2(c[14]), .Z(N14) );
  OR2D0 C417 ( .A1(g[14]), .A2(N14), .Z(c[15]) );
  AN2D0 C416 ( .A1(p[13]), .A2(c[13]), .Z(N13) );
  OR2D0 C415 ( .A1(g[13]), .A2(N13), .Z(c[14]) );
  AN2D0 C414 ( .A1(p[12]), .A2(c[12]), .Z(N12) );
  OR2D0 C413 ( .A1(g[12]), .A2(N12), .Z(c[13]) );
  AN2D0 C412 ( .A1(p[11]), .A2(c[11]), .Z(N11) );
  OR2D0 C411 ( .A1(g[11]), .A2(N11), .Z(c[12]) );
  AN2D0 C410 ( .A1(p[10]), .A2(c[10]), .Z(N10) );
  OR2D0 C409 ( .A1(g[10]), .A2(N10), .Z(c[11]) );
  AN2D0 C408 ( .A1(p[9]), .A2(c[9]), .Z(N9) );
  OR2D0 C407 ( .A1(g[9]), .A2(N9), .Z(c[10]) );
  AN2D0 C406 ( .A1(p[8]), .A2(c[8]), .Z(N8) );
  OR2D0 C405 ( .A1(g[8]), .A2(N8), .Z(c[9]) );
  AN2D0 C404 ( .A1(p[7]), .A2(c[7]), .Z(N7) );
  OR2D0 C403 ( .A1(g[7]), .A2(N7), .Z(c[8]) );
  AN2D0 C402 ( .A1(p[6]), .A2(c[6]), .Z(N6) );
  OR2D0 C401 ( .A1(g[6]), .A2(N6), .Z(c[7]) );
  AN2D0 C400 ( .A1(p[5]), .A2(c[5]), .Z(N5) );
  OR2D0 C399 ( .A1(g[5]), .A2(N5), .Z(c[6]) );
  AN2D0 C398 ( .A1(p[4]), .A2(c[4]), .Z(N4) );
  OR2D0 C397 ( .A1(g[4]), .A2(N4), .Z(c[5]) );
  AN2D0 C396 ( .A1(p[3]), .A2(c[3]), .Z(N3) );
  OR2D0 C395 ( .A1(g[3]), .A2(N3), .Z(c[4]) );
  AN2D0 C394 ( .A1(p[2]), .A2(c[2]), .Z(N2) );
  OR2D0 C393 ( .A1(g[2]), .A2(N2), .Z(c[3]) );
  AN2D0 C392 ( .A1(p[1]), .A2(c[1]), .Z(N1) );
  OR2D0 C391 ( .A1(g[1]), .A2(N1), .Z(c[2]) );
  AN2D0 C390 ( .A1(p[0]), .A2(cin), .Z(N0) );
  OR2D0 C389 ( .A1(g[0]), .A2(N0), .Z(c[1]) );
  XOR2D0 C388 ( .A1(a[0]), .A2(b[0]), .Z(p[0]) );
  XOR2D0 C387 ( .A1(a[1]), .A2(b[1]), .Z(p[1]) );
  XOR2D0 C386 ( .A1(a[2]), .A2(b[2]), .Z(p[2]) );
  XOR2D0 C385 ( .A1(a[3]), .A2(b[3]), .Z(p[3]) );
  XOR2D0 C384 ( .A1(a[4]), .A2(b[4]), .Z(p[4]) );
  XOR2D0 C383 ( .A1(a[5]), .A2(b[5]), .Z(p[5]) );
  XOR2D0 C382 ( .A1(a[6]), .A2(b[6]), .Z(p[6]) );
  XOR2D0 C381 ( .A1(a[7]), .A2(b[7]), .Z(p[7]) );
  XOR2D0 C380 ( .A1(a[8]), .A2(b[8]), .Z(p[8]) );
  XOR2D0 C379 ( .A1(a[9]), .A2(b[9]), .Z(p[9]) );
  XOR2D0 C378 ( .A1(a[10]), .A2(b[10]), .Z(p[10]) );
  XOR2D0 C377 ( .A1(a[11]), .A2(b[11]), .Z(p[11]) );
  XOR2D0 C376 ( .A1(a[12]), .A2(b[12]), .Z(p[12]) );
  XOR2D0 C375 ( .A1(a[13]), .A2(b[13]), .Z(p[13]) );
  XOR2D0 C374 ( .A1(a[14]), .A2(b[14]), .Z(p[14]) );
  XOR2D0 C373 ( .A1(a[15]), .A2(b[15]), .Z(p[15]) );
  XOR2D0 C372 ( .A1(a[16]), .A2(b[16]), .Z(p[16]) );
  XOR2D0 C371 ( .A1(a[17]), .A2(b[17]), .Z(p[17]) );
  XOR2D0 C370 ( .A1(a[18]), .A2(b[18]), .Z(p[18]) );
  XOR2D0 C369 ( .A1(a[19]), .A2(b[19]), .Z(p[19]) );
  XOR2D0 C368 ( .A1(a[20]), .A2(b[20]), .Z(p[20]) );
  XOR2D0 C367 ( .A1(a[21]), .A2(b[21]), .Z(p[21]) );
  XOR2D0 C366 ( .A1(a[22]), .A2(b[22]), .Z(p[22]) );
  XOR2D0 C365 ( .A1(a[23]), .A2(b[23]), .Z(p[23]) );
  XOR2D0 C364 ( .A1(a[24]), .A2(b[24]), .Z(p[24]) );
  XOR2D0 C363 ( .A1(a[25]), .A2(b[25]), .Z(p[25]) );
  XOR2D0 C362 ( .A1(a[26]), .A2(b[26]), .Z(p[26]) );
  XOR2D0 C361 ( .A1(a[27]), .A2(b[27]), .Z(p[27]) );
  XOR2D0 C360 ( .A1(a[28]), .A2(b[28]), .Z(p[28]) );
  XOR2D0 C359 ( .A1(a[29]), .A2(b[29]), .Z(p[29]) );
  XOR2D0 C358 ( .A1(a[30]), .A2(b[30]), .Z(p[30]) );
  XOR2D0 C357 ( .A1(a[31]), .A2(b[31]), .Z(p[31]) );
  XOR2D0 C356 ( .A1(a[32]), .A2(b[32]), .Z(p[32]) );
  XOR2D0 C355 ( .A1(a[33]), .A2(b[33]), .Z(p[33]) );
  XOR2D0 C354 ( .A1(a[34]), .A2(b[34]), .Z(p[34]) );
  XOR2D0 C353 ( .A1(a[35]), .A2(b[35]), .Z(p[35]) );
  XOR2D0 C352 ( .A1(a[36]), .A2(b[36]), .Z(p[36]) );
  XOR2D0 C351 ( .A1(a[37]), .A2(b[37]), .Z(p[37]) );
  XOR2D0 C350 ( .A1(a[38]), .A2(b[38]), .Z(p[38]) );
  XOR2D0 C349 ( .A1(a[39]), .A2(b[39]), .Z(p[39]) );
  XOR2D0 C348 ( .A1(a[40]), .A2(b[40]), .Z(p[40]) );
  XOR2D0 C347 ( .A1(a[41]), .A2(b[41]), .Z(p[41]) );
  XOR2D0 C346 ( .A1(a[42]), .A2(b[42]), .Z(p[42]) );
  XOR2D0 C345 ( .A1(a[43]), .A2(b[43]), .Z(p[43]) );
  XOR2D0 C344 ( .A1(a[44]), .A2(b[44]), .Z(p[44]) );
  XOR2D0 C343 ( .A1(a[45]), .A2(b[45]), .Z(p[45]) );
  XOR2D0 C342 ( .A1(a[46]), .A2(b[46]), .Z(p[46]) );
  XOR2D0 C341 ( .A1(a[47]), .A2(b[47]), .Z(p[47]) );
  XOR2D0 C340 ( .A1(a[48]), .A2(b[48]), .Z(p[48]) );
  XOR2D0 C339 ( .A1(a[49]), .A2(b[49]), .Z(p[49]) );
  XOR2D0 C338 ( .A1(a[50]), .A2(b[50]), .Z(p[50]) );
  XOR2D0 C337 ( .A1(a[51]), .A2(b[51]), .Z(p[51]) );
  XOR2D0 C336 ( .A1(a[52]), .A2(b[52]), .Z(p[52]) );
  XOR2D0 C335 ( .A1(a[53]), .A2(b[53]), .Z(p[53]) );
  XOR2D0 C334 ( .A1(a[54]), .A2(b[54]), .Z(p[54]) );
  XOR2D0 C333 ( .A1(a[55]), .A2(b[55]), .Z(p[55]) );
  XOR2D0 C332 ( .A1(a[56]), .A2(b[56]), .Z(p[56]) );
  XOR2D0 C331 ( .A1(a[57]), .A2(b[57]), .Z(p[57]) );
  XOR2D0 C330 ( .A1(a[58]), .A2(b[58]), .Z(p[58]) );
  XOR2D0 C329 ( .A1(a[59]), .A2(b[59]), .Z(p[59]) );
  XOR2D0 C328 ( .A1(a[60]), .A2(b[60]), .Z(p[60]) );
  XOR2D0 C327 ( .A1(a[61]), .A2(b[61]), .Z(p[61]) );
  XOR2D0 C326 ( .A1(a[62]), .A2(b[62]), .Z(p[62]) );
  XOR2D0 C325 ( .A1(a[63]), .A2(b[63]), .Z(p[63]) );
  AN2D0 C324 ( .A1(a[0]), .A2(b[0]), .Z(g[0]) );
  AN2D0 C323 ( .A1(a[1]), .A2(b[1]), .Z(g[1]) );
  AN2D0 C322 ( .A1(a[2]), .A2(b[2]), .Z(g[2]) );
  AN2D0 C321 ( .A1(a[3]), .A2(b[3]), .Z(g[3]) );
  AN2D0 C320 ( .A1(a[4]), .A2(b[4]), .Z(g[4]) );
  AN2D0 C319 ( .A1(a[5]), .A2(b[5]), .Z(g[5]) );
  AN2D0 C318 ( .A1(a[6]), .A2(b[6]), .Z(g[6]) );
  AN2D0 C317 ( .A1(a[7]), .A2(b[7]), .Z(g[7]) );
  AN2D0 C316 ( .A1(a[8]), .A2(b[8]), .Z(g[8]) );
  AN2D0 C315 ( .A1(a[9]), .A2(b[9]), .Z(g[9]) );
  AN2D0 C314 ( .A1(a[10]), .A2(b[10]), .Z(g[10]) );
  AN2D0 C313 ( .A1(a[11]), .A2(b[11]), .Z(g[11]) );
  AN2D0 C312 ( .A1(a[12]), .A2(b[12]), .Z(g[12]) );
  AN2D0 C311 ( .A1(a[13]), .A2(b[13]), .Z(g[13]) );
  AN2D0 C310 ( .A1(a[14]), .A2(b[14]), .Z(g[14]) );
  AN2D0 C309 ( .A1(a[15]), .A2(b[15]), .Z(g[15]) );
  AN2D0 C308 ( .A1(a[16]), .A2(b[16]), .Z(g[16]) );
  AN2D0 C307 ( .A1(a[17]), .A2(b[17]), .Z(g[17]) );
  AN2D0 C306 ( .A1(a[18]), .A2(b[18]), .Z(g[18]) );
  AN2D0 C305 ( .A1(a[19]), .A2(b[19]), .Z(g[19]) );
  AN2D0 C304 ( .A1(a[20]), .A2(b[20]), .Z(g[20]) );
  AN2D0 C303 ( .A1(a[21]), .A2(b[21]), .Z(g[21]) );
  AN2D0 C302 ( .A1(a[22]), .A2(b[22]), .Z(g[22]) );
  AN2D0 C301 ( .A1(a[23]), .A2(b[23]), .Z(g[23]) );
  AN2D0 C300 ( .A1(a[24]), .A2(b[24]), .Z(g[24]) );
  AN2D0 C299 ( .A1(a[25]), .A2(b[25]), .Z(g[25]) );
  AN2D0 C298 ( .A1(a[26]), .A2(b[26]), .Z(g[26]) );
  AN2D0 C297 ( .A1(a[27]), .A2(b[27]), .Z(g[27]) );
  AN2D0 C296 ( .A1(a[28]), .A2(b[28]), .Z(g[28]) );
  AN2D0 C295 ( .A1(a[29]), .A2(b[29]), .Z(g[29]) );
  AN2D0 C294 ( .A1(a[30]), .A2(b[30]), .Z(g[30]) );
  AN2D0 C293 ( .A1(a[31]), .A2(b[31]), .Z(g[31]) );
  AN2D0 C292 ( .A1(a[32]), .A2(b[32]), .Z(g[32]) );
  AN2D0 C291 ( .A1(a[33]), .A2(b[33]), .Z(g[33]) );
  AN2D0 C290 ( .A1(a[34]), .A2(b[34]), .Z(g[34]) );
  AN2D0 C289 ( .A1(a[35]), .A2(b[35]), .Z(g[35]) );
  AN2D0 C288 ( .A1(a[36]), .A2(b[36]), .Z(g[36]) );
  AN2D0 C287 ( .A1(a[37]), .A2(b[37]), .Z(g[37]) );
  AN2D0 C286 ( .A1(a[38]), .A2(b[38]), .Z(g[38]) );
  AN2D0 C285 ( .A1(a[39]), .A2(b[39]), .Z(g[39]) );
  AN2D0 C284 ( .A1(a[40]), .A2(b[40]), .Z(g[40]) );
  AN2D0 C283 ( .A1(a[41]), .A2(b[41]), .Z(g[41]) );
  AN2D0 C282 ( .A1(a[42]), .A2(b[42]), .Z(g[42]) );
  AN2D0 C281 ( .A1(a[43]), .A2(b[43]), .Z(g[43]) );
  AN2D0 C280 ( .A1(a[44]), .A2(b[44]), .Z(g[44]) );
  AN2D0 C279 ( .A1(a[45]), .A2(b[45]), .Z(g[45]) );
  AN2D0 C278 ( .A1(a[46]), .A2(b[46]), .Z(g[46]) );
  AN2D0 C277 ( .A1(a[47]), .A2(b[47]), .Z(g[47]) );
  AN2D0 C276 ( .A1(a[48]), .A2(b[48]), .Z(g[48]) );
  AN2D0 C275 ( .A1(a[49]), .A2(b[49]), .Z(g[49]) );
  AN2D0 C274 ( .A1(a[50]), .A2(b[50]), .Z(g[50]) );
  AN2D0 C273 ( .A1(a[51]), .A2(b[51]), .Z(g[51]) );
  AN2D0 C272 ( .A1(a[52]), .A2(b[52]), .Z(g[52]) );
  AN2D0 C271 ( .A1(a[53]), .A2(b[53]), .Z(g[53]) );
  AN2D0 C270 ( .A1(a[54]), .A2(b[54]), .Z(g[54]) );
  AN2D0 C269 ( .A1(a[55]), .A2(b[55]), .Z(g[55]) );
  AN2D0 C268 ( .A1(a[56]), .A2(b[56]), .Z(g[56]) );
  AN2D0 C267 ( .A1(a[57]), .A2(b[57]), .Z(g[57]) );
  AN2D0 C266 ( .A1(a[58]), .A2(b[58]), .Z(g[58]) );
  AN2D0 C265 ( .A1(a[59]), .A2(b[59]), .Z(g[59]) );
  AN2D0 C264 ( .A1(a[60]), .A2(b[60]), .Z(g[60]) );
  AN2D0 C263 ( .A1(a[61]), .A2(b[61]), .Z(g[61]) );
  AN2D0 C262 ( .A1(a[62]), .A2(b[62]), .Z(g[62]) );
endmodule

