
module cla_adder ( a, b, s, cin, cout );
  input [15:0] a;
  input [15:0] b;
  output [15:0] s;
  input cin;
  output cout;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14;
  wire   [14:0] g;
  wire   [15:0] p;
  wire   [15:1] c;

  XOR2D0 C146 ( .A1(p[0]), .A2(cin), .Z(s[0]) );
  XOR2D0 C145 ( .A1(p[1]), .A2(c[1]), .Z(s[1]) );
  XOR2D0 C144 ( .A1(p[2]), .A2(c[2]), .Z(s[2]) );
  XOR2D0 C143 ( .A1(p[3]), .A2(c[3]), .Z(s[3]) );
  XOR2D0 C142 ( .A1(p[4]), .A2(c[4]), .Z(s[4]) );
  XOR2D0 C141 ( .A1(p[5]), .A2(c[5]), .Z(s[5]) );
  XOR2D0 C140 ( .A1(p[6]), .A2(c[6]), .Z(s[6]) );
  XOR2D0 C139 ( .A1(p[7]), .A2(c[7]), .Z(s[7]) );
  XOR2D0 C138 ( .A1(p[8]), .A2(c[8]), .Z(s[8]) );
  XOR2D0 C137 ( .A1(p[9]), .A2(c[9]), .Z(s[9]) );
  XOR2D0 C136 ( .A1(p[10]), .A2(c[10]), .Z(s[10]) );
  XOR2D0 C135 ( .A1(p[11]), .A2(c[11]), .Z(s[11]) );
  XOR2D0 C134 ( .A1(p[12]), .A2(c[12]), .Z(s[12]) );
  XOR2D0 C133 ( .A1(p[13]), .A2(c[13]), .Z(s[13]) );
  XOR2D0 C132 ( .A1(p[14]), .A2(c[14]), .Z(s[14]) );
  XOR2D0 C131 ( .A1(p[15]), .A2(c[15]), .Z(s[15]) );
  AN2D0 C130 ( .A1(p[14]), .A2(c[14]), .Z(N14) );
  OR2D0 C129 ( .A1(g[14]), .A2(N14), .Z(c[15]) );
  AN2D0 C128 ( .A1(p[13]), .A2(c[13]), .Z(N13) );
  OR2D0 C127 ( .A1(g[13]), .A2(N13), .Z(c[14]) );
  AN2D0 C126 ( .A1(p[12]), .A2(c[12]), .Z(N12) );
  OR2D0 C125 ( .A1(g[12]), .A2(N12), .Z(c[13]) );
  AN2D0 C124 ( .A1(p[11]), .A2(c[11]), .Z(N11) );
  OR2D0 C123 ( .A1(g[11]), .A2(N11), .Z(c[12]) );
  AN2D0 C122 ( .A1(p[10]), .A2(c[10]), .Z(N10) );
  OR2D0 C121 ( .A1(g[10]), .A2(N10), .Z(c[11]) );
  AN2D0 C120 ( .A1(p[9]), .A2(c[9]), .Z(N9) );
  OR2D0 C119 ( .A1(g[9]), .A2(N9), .Z(c[10]) );
  AN2D0 C118 ( .A1(p[8]), .A2(c[8]), .Z(N8) );
  OR2D0 C117 ( .A1(g[8]), .A2(N8), .Z(c[9]) );
  AN2D0 C116 ( .A1(p[7]), .A2(c[7]), .Z(N7) );
  OR2D0 C115 ( .A1(g[7]), .A2(N7), .Z(c[8]) );
  AN2D0 C114 ( .A1(p[6]), .A2(c[6]), .Z(N6) );
  OR2D0 C113 ( .A1(g[6]), .A2(N6), .Z(c[7]) );
  AN2D0 C112 ( .A1(p[5]), .A2(c[5]), .Z(N5) );
  OR2D0 C111 ( .A1(g[5]), .A2(N5), .Z(c[6]) );
  AN2D0 C110 ( .A1(p[4]), .A2(c[4]), .Z(N4) );
  OR2D0 C109 ( .A1(g[4]), .A2(N4), .Z(c[5]) );
  AN2D0 C108 ( .A1(p[3]), .A2(c[3]), .Z(N3) );
  OR2D0 C107 ( .A1(g[3]), .A2(N3), .Z(c[4]) );
  AN2D0 C106 ( .A1(p[2]), .A2(c[2]), .Z(N2) );
  OR2D0 C105 ( .A1(g[2]), .A2(N2), .Z(c[3]) );
  AN2D0 C104 ( .A1(p[1]), .A2(c[1]), .Z(N1) );
  OR2D0 C103 ( .A1(g[1]), .A2(N1), .Z(c[2]) );
  AN2D0 C102 ( .A1(p[0]), .A2(cin), .Z(N0) );
  OR2D0 C101 ( .A1(g[0]), .A2(N0), .Z(c[1]) );
  XOR2D0 C100 ( .A1(a[0]), .A2(b[0]), .Z(p[0]) );
  XOR2D0 C99 ( .A1(a[1]), .A2(b[1]), .Z(p[1]) );
  XOR2D0 C98 ( .A1(a[2]), .A2(b[2]), .Z(p[2]) );
  XOR2D0 C97 ( .A1(a[3]), .A2(b[3]), .Z(p[3]) );
  XOR2D0 C96 ( .A1(a[4]), .A2(b[4]), .Z(p[4]) );
  XOR2D0 C95 ( .A1(a[5]), .A2(b[5]), .Z(p[5]) );
  XOR2D0 C94 ( .A1(a[6]), .A2(b[6]), .Z(p[6]) );
  XOR2D0 C93 ( .A1(a[7]), .A2(b[7]), .Z(p[7]) );
  XOR2D0 C92 ( .A1(a[8]), .A2(b[8]), .Z(p[8]) );
  XOR2D0 C91 ( .A1(a[9]), .A2(b[9]), .Z(p[9]) );
  XOR2D0 C90 ( .A1(a[10]), .A2(b[10]), .Z(p[10]) );
  XOR2D0 C89 ( .A1(a[11]), .A2(b[11]), .Z(p[11]) );
  XOR2D0 C88 ( .A1(a[12]), .A2(b[12]), .Z(p[12]) );
  XOR2D0 C87 ( .A1(a[13]), .A2(b[13]), .Z(p[13]) );
  XOR2D0 C86 ( .A1(a[14]), .A2(b[14]), .Z(p[14]) );
  XOR2D0 C85 ( .A1(a[15]), .A2(b[15]), .Z(p[15]) );
  AN2D0 C84 ( .A1(a[0]), .A2(b[0]), .Z(g[0]) );
  AN2D0 C83 ( .A1(a[1]), .A2(b[1]), .Z(g[1]) );
  AN2D0 C82 ( .A1(a[2]), .A2(b[2]), .Z(g[2]) );
  AN2D0 C81 ( .A1(a[3]), .A2(b[3]), .Z(g[3]) );
  AN2D0 C80 ( .A1(a[4]), .A2(b[4]), .Z(g[4]) );
  AN2D0 C79 ( .A1(a[5]), .A2(b[5]), .Z(g[5]) );
  AN2D0 C78 ( .A1(a[6]), .A2(b[6]), .Z(g[6]) );
  AN2D0 C77 ( .A1(a[7]), .A2(b[7]), .Z(g[7]) );
  AN2D0 C76 ( .A1(a[8]), .A2(b[8]), .Z(g[8]) );
  AN2D0 C75 ( .A1(a[9]), .A2(b[9]), .Z(g[9]) );
  AN2D0 C74 ( .A1(a[10]), .A2(b[10]), .Z(g[10]) );
  AN2D0 C73 ( .A1(a[11]), .A2(b[11]), .Z(g[11]) );
  AN2D0 C72 ( .A1(a[12]), .A2(b[12]), .Z(g[12]) );
  AN2D0 C71 ( .A1(a[13]), .A2(b[13]), .Z(g[13]) );
  AN2D0 C70 ( .A1(a[14]), .A2(b[14]), .Z(g[14]) );
endmodule

