module gen_linear_part(a,b,n,s);

input  [7:0] a, b; //adder inputs
input [500:0] n; // non-linear outputs
output [7:0] s;

wire [500:0] t; // non-linear outputs
//asigning bit 0
assign s[0] = (a[0] ^ b[0]);
//asigning bit 1
assign t[0] = n[0];
assign t[1] = t[0] ^ n[1];
assign t[2] = t[1] ^ n[2];

assign s[1] = ( a[1] ^ b [1] ) ^ t[2];

//asigning bit 2
assign t[3] = n[3];
assign t[4] = t[3] ^ n[4];
assign t[5] = t[4] ^ n[5];
assign t[6] = t[5] ^ n[6];
assign t[7] = t[6] ^ n[7];
assign t[8] = t[7] ^ n[8];
assign t[9] = t[8] ^ n[9];

assign s[2] = ( a[2] ^ b [2] ) ^ t[9];

//asigning bit 3
assign t[10] = n[10];
assign t[11] = t[10] ^ n[11];
assign t[12] = t[11] ^ n[12];
assign t[13] = t[12] ^ n[13];
assign t[14] = t[13] ^ n[14];
assign t[15] = t[14] ^ n[15];
assign t[16] = t[15] ^ n[16];
assign t[17] = t[16] ^ n[17];
assign t[18] = t[17] ^ n[18];
assign t[19] = t[18] ^ n[19];
assign t[20] = t[19] ^ n[20];
assign t[21] = t[20] ^ n[21];
assign t[22] = t[21] ^ n[22];
assign t[23] = t[22] ^ n[23];
assign t[24] = t[23] ^ n[24];

assign s[3] = ( a[3] ^ b [3] ) ^ t[24];

//asigning bit 4
assign t[25] = n[25];
assign t[26] = t[25] ^ n[26];
assign t[27] = t[26] ^ n[27];
assign t[28] = t[27] ^ n[28];
assign t[29] = t[28] ^ n[29];
assign t[30] = t[29] ^ n[30];
assign t[31] = t[30] ^ n[31];
assign t[32] = t[31] ^ n[32];
assign t[33] = t[32] ^ n[33];
assign t[34] = t[33] ^ n[34];
assign t[35] = t[34] ^ n[35];
assign t[36] = t[35] ^ n[36];
assign t[37] = t[36] ^ n[37];
assign t[38] = t[37] ^ n[38];
assign t[39] = t[38] ^ n[39];
assign t[40] = t[39] ^ n[40];
assign t[41] = t[40] ^ n[41];
assign t[42] = t[41] ^ n[42];
assign t[43] = t[42] ^ n[43];
assign t[44] = t[43] ^ n[44];
assign t[45] = t[44] ^ n[45];
assign t[46] = t[45] ^ n[46];
assign t[47] = t[46] ^ n[47];
assign t[48] = t[47] ^ n[48];
assign t[49] = t[48] ^ n[49];
assign t[50] = t[49] ^ n[50];
assign t[51] = t[50] ^ n[51];
assign t[52] = t[51] ^ n[52];
assign t[53] = t[52] ^ n[53];
assign t[54] = t[53] ^ n[54];
assign t[55] = t[54] ^ n[55];

assign s[4] = ( a[4] ^ b [4] ) ^ t[55];

//asigning bit 5
assign t[56] = n[56];
assign t[57] = t[56] ^ n[57];
assign t[58] = t[57] ^ n[58];
assign t[59] = t[58] ^ n[59];
assign t[60] = t[59] ^ n[60];
assign t[61] = t[60] ^ n[61];
assign t[62] = t[61] ^ n[62];
assign t[63] = t[62] ^ n[63];
assign t[64] = t[63] ^ n[64];
assign t[65] = t[64] ^ n[65];
assign t[66] = t[65] ^ n[66];
assign t[67] = t[66] ^ n[67];
assign t[68] = t[67] ^ n[68];
assign t[69] = t[68] ^ n[69];
assign t[70] = t[69] ^ n[70];
assign t[71] = t[70] ^ n[71];
assign t[72] = t[71] ^ n[72];
assign t[73] = t[72] ^ n[73];
assign t[74] = t[73] ^ n[74];
assign t[75] = t[74] ^ n[75];
assign t[76] = t[75] ^ n[76];
assign t[77] = t[76] ^ n[77];
assign t[78] = t[77] ^ n[78];
assign t[79] = t[78] ^ n[79];
assign t[80] = t[79] ^ n[80];
assign t[81] = t[80] ^ n[81];
assign t[82] = t[81] ^ n[82];
assign t[83] = t[82] ^ n[83];
assign t[84] = t[83] ^ n[84];
assign t[85] = t[84] ^ n[85];
assign t[86] = t[85] ^ n[86];
assign t[87] = t[86] ^ n[87];
assign t[88] = t[87] ^ n[88];
assign t[89] = t[88] ^ n[89];
assign t[90] = t[89] ^ n[90];
assign t[91] = t[90] ^ n[91];
assign t[92] = t[91] ^ n[92];
assign t[93] = t[92] ^ n[93];
assign t[94] = t[93] ^ n[94];
assign t[95] = t[94] ^ n[95];
assign t[96] = t[95] ^ n[96];
assign t[97] = t[96] ^ n[97];
assign t[98] = t[97] ^ n[98];
assign t[99] = t[98] ^ n[99];
assign t[100] = t[99] ^ n[100];
assign t[101] = t[100] ^ n[101];
assign t[102] = t[101] ^ n[102];
assign t[103] = t[102] ^ n[103];
assign t[104] = t[103] ^ n[104];
assign t[105] = t[104] ^ n[105];
assign t[106] = t[105] ^ n[106];
assign t[107] = t[106] ^ n[107];
assign t[108] = t[107] ^ n[108];
assign t[109] = t[108] ^ n[109];
assign t[110] = t[109] ^ n[110];
assign t[111] = t[110] ^ n[111];
assign t[112] = t[111] ^ n[112];
assign t[113] = t[112] ^ n[113];
assign t[114] = t[113] ^ n[114];
assign t[115] = t[114] ^ n[115];
assign t[116] = t[115] ^ n[116];
assign t[117] = t[116] ^ n[117];
assign t[118] = t[117] ^ n[118];

assign s[5] = ( a[5] ^ b [5] ) ^ t[118];

//asigning bit 6
assign t[119] = n[119];
assign t[120] = t[119] ^ n[120];
assign t[121] = t[120] ^ n[121];
assign t[122] = t[121] ^ n[122];
assign t[123] = t[122] ^ n[123];
assign t[124] = t[123] ^ n[124];
assign t[125] = t[124] ^ n[125];
assign t[126] = t[125] ^ n[126];
assign t[127] = t[126] ^ n[127];
assign t[128] = t[127] ^ n[128];
assign t[129] = t[128] ^ n[129];
assign t[130] = t[129] ^ n[130];
assign t[131] = t[130] ^ n[131];
assign t[132] = t[131] ^ n[132];
assign t[133] = t[132] ^ n[133];
assign t[134] = t[133] ^ n[134];
assign t[135] = t[134] ^ n[135];
assign t[136] = t[135] ^ n[136];
assign t[137] = t[136] ^ n[137];
assign t[138] = t[137] ^ n[138];
assign t[139] = t[138] ^ n[139];
assign t[140] = t[139] ^ n[140];
assign t[141] = t[140] ^ n[141];
assign t[142] = t[141] ^ n[142];
assign t[143] = t[142] ^ n[143];
assign t[144] = t[143] ^ n[144];
assign t[145] = t[144] ^ n[145];
assign t[146] = t[145] ^ n[146];
assign t[147] = t[146] ^ n[147];
assign t[148] = t[147] ^ n[148];
assign t[149] = t[148] ^ n[149];
assign t[150] = t[149] ^ n[150];
assign t[151] = t[150] ^ n[151];
assign t[152] = t[151] ^ n[152];
assign t[153] = t[152] ^ n[153];
assign t[154] = t[153] ^ n[154];
assign t[155] = t[154] ^ n[155];
assign t[156] = t[155] ^ n[156];
assign t[157] = t[156] ^ n[157];
assign t[158] = t[157] ^ n[158];
assign t[159] = t[158] ^ n[159];
assign t[160] = t[159] ^ n[160];
assign t[161] = t[160] ^ n[161];
assign t[162] = t[161] ^ n[162];
assign t[163] = t[162] ^ n[163];
assign t[164] = t[163] ^ n[164];
assign t[165] = t[164] ^ n[165];
assign t[166] = t[165] ^ n[166];
assign t[167] = t[166] ^ n[167];
assign t[168] = t[167] ^ n[168];
assign t[169] = t[168] ^ n[169];
assign t[170] = t[169] ^ n[170];
assign t[171] = t[170] ^ n[171];
assign t[172] = t[171] ^ n[172];
assign t[173] = t[172] ^ n[173];
assign t[174] = t[173] ^ n[174];
assign t[175] = t[174] ^ n[175];
assign t[176] = t[175] ^ n[176];
assign t[177] = t[176] ^ n[177];
assign t[178] = t[177] ^ n[178];
assign t[179] = t[178] ^ n[179];
assign t[180] = t[179] ^ n[180];
assign t[181] = t[180] ^ n[181];
assign t[182] = t[181] ^ n[182];
assign t[183] = t[182] ^ n[183];
assign t[184] = t[183] ^ n[184];
assign t[185] = t[184] ^ n[185];
assign t[186] = t[185] ^ n[186];
assign t[187] = t[186] ^ n[187];
assign t[188] = t[187] ^ n[188];
assign t[189] = t[188] ^ n[189];
assign t[190] = t[189] ^ n[190];
assign t[191] = t[190] ^ n[191];
assign t[192] = t[191] ^ n[192];
assign t[193] = t[192] ^ n[193];
assign t[194] = t[193] ^ n[194];
assign t[195] = t[194] ^ n[195];
assign t[196] = t[195] ^ n[196];
assign t[197] = t[196] ^ n[197];
assign t[198] = t[197] ^ n[198];
assign t[199] = t[198] ^ n[199];
assign t[200] = t[199] ^ n[200];
assign t[201] = t[200] ^ n[201];
assign t[202] = t[201] ^ n[202];
assign t[203] = t[202] ^ n[203];
assign t[204] = t[203] ^ n[204];
assign t[205] = t[204] ^ n[205];
assign t[206] = t[205] ^ n[206];
assign t[207] = t[206] ^ n[207];
assign t[208] = t[207] ^ n[208];
assign t[209] = t[208] ^ n[209];
assign t[210] = t[209] ^ n[210];
assign t[211] = t[210] ^ n[211];
assign t[212] = t[211] ^ n[212];
assign t[213] = t[212] ^ n[213];
assign t[214] = t[213] ^ n[214];
assign t[215] = t[214] ^ n[215];
assign t[216] = t[215] ^ n[216];
assign t[217] = t[216] ^ n[217];
assign t[218] = t[217] ^ n[218];
assign t[219] = t[218] ^ n[219];
assign t[220] = t[219] ^ n[220];
assign t[221] = t[220] ^ n[221];
assign t[222] = t[221] ^ n[222];
assign t[223] = t[222] ^ n[223];
assign t[224] = t[223] ^ n[224];
assign t[225] = t[224] ^ n[225];
assign t[226] = t[225] ^ n[226];
assign t[227] = t[226] ^ n[227];
assign t[228] = t[227] ^ n[228];
assign t[229] = t[228] ^ n[229];
assign t[230] = t[229] ^ n[230];
assign t[231] = t[230] ^ n[231];
assign t[232] = t[231] ^ n[232];
assign t[233] = t[232] ^ n[233];
assign t[234] = t[233] ^ n[234];
assign t[235] = t[234] ^ n[235];
assign t[236] = t[235] ^ n[236];
assign t[237] = t[236] ^ n[237];
assign t[238] = t[237] ^ n[238];
assign t[239] = t[238] ^ n[239];
assign t[240] = t[239] ^ n[240];
assign t[241] = t[240] ^ n[241];
assign t[242] = t[241] ^ n[242];
assign t[243] = t[242] ^ n[243];
assign t[244] = t[243] ^ n[244];
assign t[245] = t[244] ^ n[245];

assign s[6] = ( a[6] ^ b [6] ) ^ t[245];

//asigning bit 7
assign t[246] = n[246];
assign t[247] = t[246] ^ n[247];
assign t[248] = t[247] ^ n[248];
assign t[249] = t[248] ^ n[249];
assign t[250] = t[249] ^ n[250];
assign t[251] = t[250] ^ n[251];
assign t[252] = t[251] ^ n[252];
assign t[253] = t[252] ^ n[253];
assign t[254] = t[253] ^ n[254];
assign t[255] = t[254] ^ n[255];
assign t[256] = t[255] ^ n[256];
assign t[257] = t[256] ^ n[257];
assign t[258] = t[257] ^ n[258];
assign t[259] = t[258] ^ n[259];
assign t[260] = t[259] ^ n[260];
assign t[261] = t[260] ^ n[261];
assign t[262] = t[261] ^ n[262];
assign t[263] = t[262] ^ n[263];
assign t[264] = t[263] ^ n[264];
assign t[265] = t[264] ^ n[265];
assign t[266] = t[265] ^ n[266];
assign t[267] = t[266] ^ n[267];
assign t[268] = t[267] ^ n[268];
assign t[269] = t[268] ^ n[269];
assign t[270] = t[269] ^ n[270];
assign t[271] = t[270] ^ n[271];
assign t[272] = t[271] ^ n[272];
assign t[273] = t[272] ^ n[273];
assign t[274] = t[273] ^ n[274];
assign t[275] = t[274] ^ n[275];
assign t[276] = t[275] ^ n[276];
assign t[277] = t[276] ^ n[277];
assign t[278] = t[277] ^ n[278];
assign t[279] = t[278] ^ n[279];
assign t[280] = t[279] ^ n[280];
assign t[281] = t[280] ^ n[281];
assign t[282] = t[281] ^ n[282];
assign t[283] = t[282] ^ n[283];
assign t[284] = t[283] ^ n[284];
assign t[285] = t[284] ^ n[285];
assign t[286] = t[285] ^ n[286];
assign t[287] = t[286] ^ n[287];
assign t[288] = t[287] ^ n[288];
assign t[289] = t[288] ^ n[289];
assign t[290] = t[289] ^ n[290];
assign t[291] = t[290] ^ n[291];
assign t[292] = t[291] ^ n[292];
assign t[293] = t[292] ^ n[293];
assign t[294] = t[293] ^ n[294];
assign t[295] = t[294] ^ n[295];
assign t[296] = t[295] ^ n[296];
assign t[297] = t[296] ^ n[297];
assign t[298] = t[297] ^ n[298];
assign t[299] = t[298] ^ n[299];
assign t[300] = t[299] ^ n[300];
assign t[301] = t[300] ^ n[301];
assign t[302] = t[301] ^ n[302];
assign t[303] = t[302] ^ n[303];
assign t[304] = t[303] ^ n[304];
assign t[305] = t[304] ^ n[305];
assign t[306] = t[305] ^ n[306];
assign t[307] = t[306] ^ n[307];
assign t[308] = t[307] ^ n[308];
assign t[309] = t[308] ^ n[309];
assign t[310] = t[309] ^ n[310];
assign t[311] = t[310] ^ n[311];
assign t[312] = t[311] ^ n[312];
assign t[313] = t[312] ^ n[313];
assign t[314] = t[313] ^ n[314];
assign t[315] = t[314] ^ n[315];
assign t[316] = t[315] ^ n[316];
assign t[317] = t[316] ^ n[317];
assign t[318] = t[317] ^ n[318];
assign t[319] = t[318] ^ n[319];
assign t[320] = t[319] ^ n[320];
assign t[321] = t[320] ^ n[321];
assign t[322] = t[321] ^ n[322];
assign t[323] = t[322] ^ n[323];
assign t[324] = t[323] ^ n[324];
assign t[325] = t[324] ^ n[325];
assign t[326] = t[325] ^ n[326];
assign t[327] = t[326] ^ n[327];
assign t[328] = t[327] ^ n[328];
assign t[329] = t[328] ^ n[329];
assign t[330] = t[329] ^ n[330];
assign t[331] = t[330] ^ n[331];
assign t[332] = t[331] ^ n[332];
assign t[333] = t[332] ^ n[333];
assign t[334] = t[333] ^ n[334];
assign t[335] = t[334] ^ n[335];
assign t[336] = t[335] ^ n[336];
assign t[337] = t[336] ^ n[337];
assign t[338] = t[337] ^ n[338];
assign t[339] = t[338] ^ n[339];
assign t[340] = t[339] ^ n[340];
assign t[341] = t[340] ^ n[341];
assign t[342] = t[341] ^ n[342];
assign t[343] = t[342] ^ n[343];
assign t[344] = t[343] ^ n[344];
assign t[345] = t[344] ^ n[345];
assign t[346] = t[345] ^ n[346];
assign t[347] = t[346] ^ n[347];
assign t[348] = t[347] ^ n[348];
assign t[349] = t[348] ^ n[349];
assign t[350] = t[349] ^ n[350];
assign t[351] = t[350] ^ n[351];
assign t[352] = t[351] ^ n[352];
assign t[353] = t[352] ^ n[353];
assign t[354] = t[353] ^ n[354];
assign t[355] = t[354] ^ n[355];
assign t[356] = t[355] ^ n[356];
assign t[357] = t[356] ^ n[357];
assign t[358] = t[357] ^ n[358];
assign t[359] = t[358] ^ n[359];
assign t[360] = t[359] ^ n[360];
assign t[361] = t[360] ^ n[361];
assign t[362] = t[361] ^ n[362];
assign t[363] = t[362] ^ n[363];
assign t[364] = t[363] ^ n[364];
assign t[365] = t[364] ^ n[365];
assign t[366] = t[365] ^ n[366];
assign t[367] = t[366] ^ n[367];
assign t[368] = t[367] ^ n[368];
assign t[369] = t[368] ^ n[369];
assign t[370] = t[369] ^ n[370];
assign t[371] = t[370] ^ n[371];
assign t[372] = t[371] ^ n[372];
assign t[373] = t[372] ^ n[373];
assign t[374] = t[373] ^ n[374];
assign t[375] = t[374] ^ n[375];
assign t[376] = t[375] ^ n[376];
assign t[377] = t[376] ^ n[377];
assign t[378] = t[377] ^ n[378];
assign t[379] = t[378] ^ n[379];
assign t[380] = t[379] ^ n[380];
assign t[381] = t[380] ^ n[381];
assign t[382] = t[381] ^ n[382];
assign t[383] = t[382] ^ n[383];
assign t[384] = t[383] ^ n[384];
assign t[385] = t[384] ^ n[385];
assign t[386] = t[385] ^ n[386];
assign t[387] = t[386] ^ n[387];
assign t[388] = t[387] ^ n[388];
assign t[389] = t[388] ^ n[389];
assign t[390] = t[389] ^ n[390];
assign t[391] = t[390] ^ n[391];
assign t[392] = t[391] ^ n[392];
assign t[393] = t[392] ^ n[393];
assign t[394] = t[393] ^ n[394];
assign t[395] = t[394] ^ n[395];
assign t[396] = t[395] ^ n[396];
assign t[397] = t[396] ^ n[397];
assign t[398] = t[397] ^ n[398];
assign t[399] = t[398] ^ n[399];
assign t[400] = t[399] ^ n[400];
assign t[401] = t[400] ^ n[401];
assign t[402] = t[401] ^ n[402];
assign t[403] = t[402] ^ n[403];
assign t[404] = t[403] ^ n[404];
assign t[405] = t[404] ^ n[405];
assign t[406] = t[405] ^ n[406];
assign t[407] = t[406] ^ n[407];
assign t[408] = t[407] ^ n[408];
assign t[409] = t[408] ^ n[409];
assign t[410] = t[409] ^ n[410];
assign t[411] = t[410] ^ n[411];
assign t[412] = t[411] ^ n[412];
assign t[413] = t[412] ^ n[413];
assign t[414] = t[413] ^ n[414];
assign t[415] = t[414] ^ n[415];
assign t[416] = t[415] ^ n[416];
assign t[417] = t[416] ^ n[417];
assign t[418] = t[417] ^ n[418];
assign t[419] = t[418] ^ n[419];
assign t[420] = t[419] ^ n[420];
assign t[421] = t[420] ^ n[421];
assign t[422] = t[421] ^ n[422];
assign t[423] = t[422] ^ n[423];
assign t[424] = t[423] ^ n[424];
assign t[425] = t[424] ^ n[425];
assign t[426] = t[425] ^ n[426];
assign t[427] = t[426] ^ n[427];
assign t[428] = t[427] ^ n[428];
assign t[429] = t[428] ^ n[429];
assign t[430] = t[429] ^ n[430];
assign t[431] = t[430] ^ n[431];
assign t[432] = t[431] ^ n[432];
assign t[433] = t[432] ^ n[433];
assign t[434] = t[433] ^ n[434];
assign t[435] = t[434] ^ n[435];
assign t[436] = t[435] ^ n[436];
assign t[437] = t[436] ^ n[437];
assign t[438] = t[437] ^ n[438];
assign t[439] = t[438] ^ n[439];
assign t[440] = t[439] ^ n[440];
assign t[441] = t[440] ^ n[441];
assign t[442] = t[441] ^ n[442];
assign t[443] = t[442] ^ n[443];
assign t[444] = t[443] ^ n[444];
assign t[445] = t[444] ^ n[445];
assign t[446] = t[445] ^ n[446];
assign t[447] = t[446] ^ n[447];
assign t[448] = t[447] ^ n[448];
assign t[449] = t[448] ^ n[449];
assign t[450] = t[449] ^ n[450];
assign t[451] = t[450] ^ n[451];
assign t[452] = t[451] ^ n[452];
assign t[453] = t[452] ^ n[453];
assign t[454] = t[453] ^ n[454];
assign t[455] = t[454] ^ n[455];
assign t[456] = t[455] ^ n[456];
assign t[457] = t[456] ^ n[457];
assign t[458] = t[457] ^ n[458];
assign t[459] = t[458] ^ n[459];
assign t[460] = t[459] ^ n[460];
assign t[461] = t[460] ^ n[461];
assign t[462] = t[461] ^ n[462];
assign t[463] = t[462] ^ n[463];
assign t[464] = t[463] ^ n[464];
assign t[465] = t[464] ^ n[465];
assign t[466] = t[465] ^ n[466];
assign t[467] = t[466] ^ n[467];
assign t[468] = t[467] ^ n[468];
assign t[469] = t[468] ^ n[469];
assign t[470] = t[469] ^ n[470];
assign t[471] = t[470] ^ n[471];
assign t[472] = t[471] ^ n[472];
assign t[473] = t[472] ^ n[473];
assign t[474] = t[473] ^ n[474];
assign t[475] = t[474] ^ n[475];
assign t[476] = t[475] ^ n[476];
assign t[477] = t[476] ^ n[477];
assign t[478] = t[477] ^ n[478];
assign t[479] = t[478] ^ n[479];
assign t[480] = t[479] ^ n[480];
assign t[481] = t[480] ^ n[481];
assign t[482] = t[481] ^ n[482];
assign t[483] = t[482] ^ n[483];
assign t[484] = t[483] ^ n[484];
assign t[485] = t[484] ^ n[485];
assign t[486] = t[485] ^ n[486];
assign t[487] = t[486] ^ n[487];
assign t[488] = t[487] ^ n[488];
assign t[489] = t[488] ^ n[489];
assign t[490] = t[489] ^ n[490];
assign t[491] = t[490] ^ n[491];
assign t[492] = t[491] ^ n[492];
assign t[493] = t[492] ^ n[493];
assign t[494] = t[493] ^ n[494];
assign t[495] = t[494] ^ n[495];
assign t[496] = t[495] ^ n[496];
assign t[497] = t[496] ^ n[497];
assign t[498] = t[497] ^ n[498];
assign t[499] = t[498] ^ n[499];
assign t[500] = t[499] ^ n[500];

assign s[7] = ( a[7] ^ b [7] ) ^ t[500];

endmodule