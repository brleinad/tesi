module adder7bit_P();

input [13:0]  c;
output [13:0] s;

s[0] = c[1] ^ c[4] ^ c[]

endmodule
