
module gen_linear_part ( a, b, n, s );
  input [6:0] a;
  input [6:0] b;
  input [245:0] n;
  output [6:0] s;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246;

  XOR2D0 U1 ( .A1(n1), .A2(n2), .Z(s[6]) );
  XOR2D0 U2 ( .A1(n[243]), .A2(n[242]), .Z(n2) );
  XOR2D0 U3 ( .A1(n3), .A2(n4), .Z(n1) );
  XOR2D0 U4 ( .A1(n5), .A2(n6), .Z(n4) );
  XOR2D0 U5 ( .A1(a[6]), .A2(n7), .Z(n6) );
  XOR2D0 U6 ( .A1(n8), .A2(n9), .Z(n7) );
  XOR2D0 U7 ( .A1(n10), .A2(n11), .Z(n9) );
  XOR2D0 U8 ( .A1(n[232]), .A2(n12), .Z(n11) );
  XOR2D0 U9 ( .A1(n13), .A2(n14), .Z(n12) );
  XOR2D0 U10 ( .A1(n15), .A2(n16), .Z(n14) );
  XOR2D0 U11 ( .A1(n[225]), .A2(n17), .Z(n16) );
  XOR2D0 U12 ( .A1(n18), .A2(n19), .Z(n17) );
  XOR2D0 U13 ( .A1(n20), .A2(n21), .Z(n19) );
  XOR2D0 U14 ( .A1(n[218]), .A2(n22), .Z(n21) );
  XOR2D0 U15 ( .A1(n23), .A2(n24), .Z(n22) );
  XOR2D0 U16 ( .A1(n25), .A2(n26), .Z(n24) );
  XOR2D0 U17 ( .A1(n[211]), .A2(n27), .Z(n26) );
  XOR2D0 U18 ( .A1(n28), .A2(n29), .Z(n27) );
  XOR2D0 U19 ( .A1(n30), .A2(n31), .Z(n29) );
  XOR2D0 U20 ( .A1(n[204]), .A2(n32), .Z(n31) );
  XOR2D0 U21 ( .A1(n33), .A2(n34), .Z(n32) );
  XOR2D0 U22 ( .A1(n35), .A2(n36), .Z(n34) );
  XOR2D0 U23 ( .A1(n[197]), .A2(n37), .Z(n36) );
  XOR2D0 U24 ( .A1(n38), .A2(n39), .Z(n37) );
  XOR2D0 U25 ( .A1(n40), .A2(n41), .Z(n39) );
  XOR2D0 U26 ( .A1(n[190]), .A2(n42), .Z(n41) );
  XOR2D0 U27 ( .A1(n43), .A2(n44), .Z(n42) );
  XOR2D0 U28 ( .A1(n45), .A2(n46), .Z(n44) );
  XOR2D0 U29 ( .A1(n[183]), .A2(n47), .Z(n46) );
  XOR2D0 U30 ( .A1(n48), .A2(n49), .Z(n47) );
  XOR2D0 U31 ( .A1(n50), .A2(n51), .Z(n49) );
  XOR2D0 U32 ( .A1(n[176]), .A2(n52), .Z(n51) );
  XOR2D0 U33 ( .A1(n53), .A2(n54), .Z(n52) );
  XOR2D0 U34 ( .A1(n55), .A2(n56), .Z(n54) );
  XOR2D0 U35 ( .A1(n[169]), .A2(n57), .Z(n56) );
  XOR2D0 U36 ( .A1(n58), .A2(n59), .Z(n57) );
  XOR2D0 U37 ( .A1(n60), .A2(n61), .Z(n59) );
  XOR2D0 U38 ( .A1(n[162]), .A2(n62), .Z(n61) );
  XOR2D0 U39 ( .A1(n63), .A2(n64), .Z(n62) );
  XOR2D0 U40 ( .A1(n65), .A2(n66), .Z(n64) );
  XOR2D0 U41 ( .A1(n[155]), .A2(n67), .Z(n66) );
  XOR2D0 U42 ( .A1(n68), .A2(n69), .Z(n67) );
  XOR2D0 U43 ( .A1(n70), .A2(n71), .Z(n69) );
  XOR2D0 U44 ( .A1(n[148]), .A2(n72), .Z(n71) );
  XOR2D0 U45 ( .A1(n73), .A2(n74), .Z(n72) );
  XOR2D0 U46 ( .A1(n75), .A2(n76), .Z(n74) );
  XOR2D0 U47 ( .A1(n[141]), .A2(n77), .Z(n76) );
  XOR2D0 U48 ( .A1(n78), .A2(n79), .Z(n77) );
  XOR2D0 U49 ( .A1(n80), .A2(n81), .Z(n79) );
  XOR2D0 U50 ( .A1(n[134]), .A2(n82), .Z(n81) );
  XOR2D0 U51 ( .A1(n83), .A2(n84), .Z(n82) );
  XOR2D0 U52 ( .A1(n85), .A2(n86), .Z(n84) );
  XOR2D0 U53 ( .A1(n[127]), .A2(n87), .Z(n86) );
  XOR2D0 U54 ( .A1(n88), .A2(n89), .Z(n87) );
  XOR2D0 U55 ( .A1(n90), .A2(n91), .Z(n89) );
  XOR2D0 U56 ( .A1(n[120]), .A2(n[119]), .Z(n91) );
  XOR2D0 U57 ( .A1(n[122]), .A2(n[121]), .Z(n90) );
  XOR2D0 U58 ( .A1(n92), .A2(n93), .Z(n88) );
  XOR2D0 U59 ( .A1(n[124]), .A2(n[123]), .Z(n93) );
  XOR2D0 U60 ( .A1(n[126]), .A2(n[125]), .Z(n92) );
  XOR2D0 U61 ( .A1(n[129]), .A2(n[128]), .Z(n85) );
  XOR2D0 U62 ( .A1(n94), .A2(n95), .Z(n83) );
  XOR2D0 U63 ( .A1(n[131]), .A2(n[130]), .Z(n95) );
  XOR2D0 U64 ( .A1(n[133]), .A2(n[132]), .Z(n94) );
  XOR2D0 U65 ( .A1(n[136]), .A2(n[135]), .Z(n80) );
  XOR2D0 U66 ( .A1(n96), .A2(n97), .Z(n78) );
  XOR2D0 U67 ( .A1(n[138]), .A2(n[137]), .Z(n97) );
  XOR2D0 U68 ( .A1(n[140]), .A2(n[139]), .Z(n96) );
  XOR2D0 U69 ( .A1(n[143]), .A2(n[142]), .Z(n75) );
  XOR2D0 U70 ( .A1(n98), .A2(n99), .Z(n73) );
  XOR2D0 U71 ( .A1(n[145]), .A2(n[144]), .Z(n99) );
  XOR2D0 U72 ( .A1(n[147]), .A2(n[146]), .Z(n98) );
  XOR2D0 U73 ( .A1(n[150]), .A2(n[149]), .Z(n70) );
  XOR2D0 U74 ( .A1(n100), .A2(n101), .Z(n68) );
  XOR2D0 U75 ( .A1(n[152]), .A2(n[151]), .Z(n101) );
  XOR2D0 U76 ( .A1(n[154]), .A2(n[153]), .Z(n100) );
  XOR2D0 U77 ( .A1(n[157]), .A2(n[156]), .Z(n65) );
  XOR2D0 U78 ( .A1(n102), .A2(n103), .Z(n63) );
  XOR2D0 U79 ( .A1(n[159]), .A2(n[158]), .Z(n103) );
  XOR2D0 U80 ( .A1(n[161]), .A2(n[160]), .Z(n102) );
  XOR2D0 U81 ( .A1(n[164]), .A2(n[163]), .Z(n60) );
  XOR2D0 U82 ( .A1(n104), .A2(n105), .Z(n58) );
  XOR2D0 U83 ( .A1(n[166]), .A2(n[165]), .Z(n105) );
  XOR2D0 U84 ( .A1(n[168]), .A2(n[167]), .Z(n104) );
  XOR2D0 U85 ( .A1(n[171]), .A2(n[170]), .Z(n55) );
  XOR2D0 U86 ( .A1(n106), .A2(n107), .Z(n53) );
  XOR2D0 U87 ( .A1(n[173]), .A2(n[172]), .Z(n107) );
  XOR2D0 U88 ( .A1(n[175]), .A2(n[174]), .Z(n106) );
  XOR2D0 U89 ( .A1(n[178]), .A2(n[177]), .Z(n50) );
  XOR2D0 U90 ( .A1(n108), .A2(n109), .Z(n48) );
  XOR2D0 U91 ( .A1(n[180]), .A2(n[179]), .Z(n109) );
  XOR2D0 U92 ( .A1(n[182]), .A2(n[181]), .Z(n108) );
  XOR2D0 U93 ( .A1(n[185]), .A2(n[184]), .Z(n45) );
  XOR2D0 U94 ( .A1(n110), .A2(n111), .Z(n43) );
  XOR2D0 U95 ( .A1(n[187]), .A2(n[186]), .Z(n111) );
  XOR2D0 U96 ( .A1(n[189]), .A2(n[188]), .Z(n110) );
  XOR2D0 U97 ( .A1(n[192]), .A2(n[191]), .Z(n40) );
  XOR2D0 U98 ( .A1(n112), .A2(n113), .Z(n38) );
  XOR2D0 U99 ( .A1(n[194]), .A2(n[193]), .Z(n113) );
  XOR2D0 U100 ( .A1(n[196]), .A2(n[195]), .Z(n112) );
  XOR2D0 U101 ( .A1(n[199]), .A2(n[198]), .Z(n35) );
  XOR2D0 U102 ( .A1(n114), .A2(n115), .Z(n33) );
  XOR2D0 U103 ( .A1(n[201]), .A2(n[200]), .Z(n115) );
  XOR2D0 U104 ( .A1(n[203]), .A2(n[202]), .Z(n114) );
  XOR2D0 U105 ( .A1(n[206]), .A2(n[205]), .Z(n30) );
  XOR2D0 U106 ( .A1(n116), .A2(n117), .Z(n28) );
  XOR2D0 U107 ( .A1(n[208]), .A2(n[207]), .Z(n117) );
  XOR2D0 U108 ( .A1(n[210]), .A2(n[209]), .Z(n116) );
  XOR2D0 U109 ( .A1(n[213]), .A2(n[212]), .Z(n25) );
  XOR2D0 U110 ( .A1(n118), .A2(n119), .Z(n23) );
  XOR2D0 U111 ( .A1(n[215]), .A2(n[214]), .Z(n119) );
  XOR2D0 U112 ( .A1(n[217]), .A2(n[216]), .Z(n118) );
  XOR2D0 U113 ( .A1(n[220]), .A2(n[219]), .Z(n20) );
  XOR2D0 U114 ( .A1(n120), .A2(n121), .Z(n18) );
  XOR2D0 U115 ( .A1(n[222]), .A2(n[221]), .Z(n121) );
  XOR2D0 U116 ( .A1(n[224]), .A2(n[223]), .Z(n120) );
  XOR2D0 U117 ( .A1(n[227]), .A2(n[226]), .Z(n15) );
  XOR2D0 U118 ( .A1(n122), .A2(n123), .Z(n13) );
  XOR2D0 U119 ( .A1(n[229]), .A2(n[228]), .Z(n123) );
  XOR2D0 U120 ( .A1(n[231]), .A2(n[230]), .Z(n122) );
  XOR2D0 U121 ( .A1(n[234]), .A2(n[233]), .Z(n10) );
  XOR2D0 U122 ( .A1(n124), .A2(n125), .Z(n8) );
  XOR2D0 U123 ( .A1(n[236]), .A2(n[235]), .Z(n125) );
  XOR2D0 U124 ( .A1(n[238]), .A2(n[237]), .Z(n124) );
  XOR2D0 U125 ( .A1(n[239]), .A2(b[6]), .Z(n5) );
  XOR2D0 U126 ( .A1(n126), .A2(n127), .Z(n3) );
  XOR2D0 U127 ( .A1(n[241]), .A2(n[240]), .Z(n127) );
  XOR2D0 U128 ( .A1(n[245]), .A2(n[244]), .Z(n126) );
  XOR2D0 U129 ( .A1(n128), .A2(n129), .Z(s[5]) );
  XOR2D0 U130 ( .A1(n[115]), .A2(n130), .Z(n129) );
  XOR2D0 U131 ( .A1(n131), .A2(n132), .Z(n130) );
  XOR2D0 U132 ( .A1(a[5]), .A2(n133), .Z(n132) );
  XOR2D0 U133 ( .A1(n134), .A2(n135), .Z(n133) );
  XOR2D0 U134 ( .A1(n136), .A2(n137), .Z(n135) );
  XOR2D0 U135 ( .A1(n[106]), .A2(n138), .Z(n137) );
  XOR2D0 U136 ( .A1(n139), .A2(n140), .Z(n138) );
  XOR2D0 U137 ( .A1(n141), .A2(n142), .Z(n140) );
  XOR2D0 U138 ( .A1(n[100]), .A2(n143), .Z(n142) );
  XOR2D0 U139 ( .A1(n144), .A2(n145), .Z(n143) );
  XOR2D0 U140 ( .A1(n146), .A2(n147), .Z(n145) );
  XOR2D0 U141 ( .A1(n[92]), .A2(n148), .Z(n147) );
  XOR2D0 U142 ( .A1(n149), .A2(n150), .Z(n148) );
  XOR2D0 U143 ( .A1(n151), .A2(n152), .Z(n150) );
  XOR2D0 U144 ( .A1(n[85]), .A2(n153), .Z(n152) );
  XOR2D0 U145 ( .A1(n154), .A2(n155), .Z(n153) );
  XOR2D0 U146 ( .A1(n156), .A2(n157), .Z(n155) );
  XOR2D0 U147 ( .A1(n[78]), .A2(n158), .Z(n157) );
  XOR2D0 U148 ( .A1(n159), .A2(n160), .Z(n158) );
  XOR2D0 U149 ( .A1(n161), .A2(n162), .Z(n160) );
  XOR2D0 U150 ( .A1(n[71]), .A2(n163), .Z(n162) );
  XOR2D0 U151 ( .A1(n164), .A2(n165), .Z(n163) );
  XOR2D0 U152 ( .A1(n166), .A2(n167), .Z(n165) );
  XOR2D0 U153 ( .A1(n[64]), .A2(n168), .Z(n167) );
  XOR2D0 U154 ( .A1(n169), .A2(n170), .Z(n168) );
  XOR2D0 U155 ( .A1(n171), .A2(n172), .Z(n170) );
  XOR2D0 U156 ( .A1(n[57]), .A2(n[56]), .Z(n172) );
  XOR2D0 U157 ( .A1(n[59]), .A2(n[58]), .Z(n171) );
  XOR2D0 U158 ( .A1(n173), .A2(n174), .Z(n169) );
  XOR2D0 U159 ( .A1(n[61]), .A2(n[60]), .Z(n174) );
  XOR2D0 U160 ( .A1(n[63]), .A2(n[62]), .Z(n173) );
  XOR2D0 U161 ( .A1(n[66]), .A2(n[65]), .Z(n166) );
  XOR2D0 U162 ( .A1(n175), .A2(n176), .Z(n164) );
  XOR2D0 U163 ( .A1(n[68]), .A2(n[67]), .Z(n176) );
  XOR2D0 U164 ( .A1(n[70]), .A2(n[69]), .Z(n175) );
  XOR2D0 U165 ( .A1(n[73]), .A2(n[72]), .Z(n161) );
  XOR2D0 U166 ( .A1(n177), .A2(n178), .Z(n159) );
  XOR2D0 U167 ( .A1(n[75]), .A2(n[74]), .Z(n178) );
  XOR2D0 U168 ( .A1(n[77]), .A2(n[76]), .Z(n177) );
  XOR2D0 U169 ( .A1(n[80]), .A2(n[79]), .Z(n156) );
  XOR2D0 U170 ( .A1(n179), .A2(n180), .Z(n154) );
  XOR2D0 U171 ( .A1(n[82]), .A2(n[81]), .Z(n180) );
  XOR2D0 U172 ( .A1(n[84]), .A2(n[83]), .Z(n179) );
  XOR2D0 U173 ( .A1(n[87]), .A2(n[86]), .Z(n151) );
  XOR2D0 U174 ( .A1(n181), .A2(n182), .Z(n149) );
  XOR2D0 U175 ( .A1(n[89]), .A2(n[88]), .Z(n182) );
  XOR2D0 U176 ( .A1(n[91]), .A2(n[90]), .Z(n181) );
  XOR2D0 U177 ( .A1(n[94]), .A2(n[93]), .Z(n146) );
  XOR2D0 U178 ( .A1(n183), .A2(n184), .Z(n144) );
  XOR2D0 U179 ( .A1(n[96]), .A2(n[95]), .Z(n184) );
  XOR2D0 U180 ( .A1(n[98]), .A2(n[97]), .Z(n183) );
  XOR2D0 U181 ( .A1(n[102]), .A2(n[101]), .Z(n141) );
  XOR2D0 U182 ( .A1(n185), .A2(n186), .Z(n139) );
  XOR2D0 U183 ( .A1(n[104]), .A2(n[103]), .Z(n186) );
  XOR2D0 U184 ( .A1(n[99]), .A2(n[105]), .Z(n185) );
  XOR2D0 U185 ( .A1(n[108]), .A2(n[107]), .Z(n136) );
  XOR2D0 U186 ( .A1(n187), .A2(n188), .Z(n134) );
  XOR2D0 U187 ( .A1(n[110]), .A2(n[109]), .Z(n188) );
  XOR2D0 U188 ( .A1(n[112]), .A2(n[111]), .Z(n187) );
  XOR2D0 U189 ( .A1(b[5]), .A2(n189), .Z(n131) );
  XOR2D0 U190 ( .A1(n[114]), .A2(n[113]), .Z(n189) );
  XOR2D0 U191 ( .A1(n[116]), .A2(n190), .Z(n128) );
  XOR2D0 U192 ( .A1(n[118]), .A2(n[117]), .Z(n190) );
  XOR2D0 U193 ( .A1(n191), .A2(n192), .Z(s[4]) );
  XOR2D0 U194 ( .A1(a[4]), .A2(n193), .Z(n192) );
  XOR2D0 U195 ( .A1(n194), .A2(n195), .Z(n193) );
  XOR2D0 U196 ( .A1(n196), .A2(n197), .Z(n195) );
  XOR2D0 U197 ( .A1(n[47]), .A2(n198), .Z(n197) );
  XOR2D0 U198 ( .A1(n199), .A2(n200), .Z(n198) );
  XOR2D0 U199 ( .A1(n201), .A2(n202), .Z(n200) );
  XOR2D0 U200 ( .A1(n[40]), .A2(n203), .Z(n202) );
  XOR2D0 U201 ( .A1(n204), .A2(n205), .Z(n203) );
  XOR2D0 U202 ( .A1(n206), .A2(n207), .Z(n205) );
  XOR2D0 U203 ( .A1(n[33]), .A2(n208), .Z(n207) );
  XOR2D0 U204 ( .A1(n209), .A2(n210), .Z(n208) );
  XOR2D0 U205 ( .A1(n211), .A2(n212), .Z(n210) );
  XOR2D0 U206 ( .A1(n[26]), .A2(n[25]), .Z(n212) );
  XOR2D0 U207 ( .A1(n[28]), .A2(n[27]), .Z(n211) );
  XOR2D0 U208 ( .A1(n213), .A2(n214), .Z(n209) );
  XOR2D0 U209 ( .A1(n[30]), .A2(n[29]), .Z(n214) );
  XOR2D0 U210 ( .A1(n[32]), .A2(n[31]), .Z(n213) );
  XOR2D0 U211 ( .A1(n[35]), .A2(n[34]), .Z(n206) );
  XOR2D0 U212 ( .A1(n215), .A2(n216), .Z(n204) );
  XOR2D0 U213 ( .A1(n[37]), .A2(n[36]), .Z(n216) );
  XOR2D0 U214 ( .A1(n[39]), .A2(n[38]), .Z(n215) );
  XOR2D0 U215 ( .A1(n[42]), .A2(n[41]), .Z(n201) );
  XOR2D0 U216 ( .A1(n217), .A2(n218), .Z(n199) );
  XOR2D0 U217 ( .A1(n[44]), .A2(n[43]), .Z(n218) );
  XOR2D0 U218 ( .A1(n[46]), .A2(n[45]), .Z(n217) );
  XOR2D0 U219 ( .A1(n[49]), .A2(n[48]), .Z(n196) );
  XOR2D0 U220 ( .A1(n219), .A2(n220), .Z(n194) );
  XOR2D0 U221 ( .A1(n[51]), .A2(n[50]), .Z(n220) );
  XOR2D0 U222 ( .A1(n[53]), .A2(n[52]), .Z(n219) );
  XOR2D0 U223 ( .A1(b[4]), .A2(n221), .Z(n191) );
  XOR2D0 U224 ( .A1(n[55]), .A2(n[54]), .Z(n221) );
  XOR2D0 U225 ( .A1(n222), .A2(n223), .Z(s[3]) );
  XOR2D0 U226 ( .A1(n[22]), .A2(n[21]), .Z(n223) );
  XOR2D0 U227 ( .A1(n224), .A2(n225), .Z(n222) );
  XOR2D0 U228 ( .A1(n226), .A2(n227), .Z(n225) );
  XOR2D0 U229 ( .A1(a[3]), .A2(n228), .Z(n227) );
  XOR2D0 U230 ( .A1(n229), .A2(n230), .Z(n228) );
  XOR2D0 U231 ( .A1(n231), .A2(n232), .Z(n230) );
  XOR2D0 U232 ( .A1(n[11]), .A2(n[10]), .Z(n232) );
  XOR2D0 U233 ( .A1(n[13]), .A2(n[12]), .Z(n231) );
  XOR2D0 U234 ( .A1(n233), .A2(n234), .Z(n229) );
  XOR2D0 U235 ( .A1(n[15]), .A2(n[14]), .Z(n234) );
  XOR2D0 U236 ( .A1(n[17]), .A2(n[16]), .Z(n233) );
  XOR2D0 U237 ( .A1(n[18]), .A2(b[3]), .Z(n226) );
  XOR2D0 U238 ( .A1(n235), .A2(n236), .Z(n224) );
  XOR2D0 U239 ( .A1(n[20]), .A2(n[19]), .Z(n236) );
  XOR2D0 U240 ( .A1(n[24]), .A2(n[23]), .Z(n235) );
  XOR2D0 U241 ( .A1(n[6]), .A2(n237), .Z(s[2]) );
  XOR2D0 U242 ( .A1(n238), .A2(n239), .Z(n237) );
  XOR2D0 U243 ( .A1(n240), .A2(n241), .Z(n239) );
  XOR2D0 U244 ( .A1(b[2]), .A2(a[2]), .Z(n241) );
  XOR2D0 U245 ( .A1(n[4]), .A2(n[3]), .Z(n240) );
  XOR2D0 U246 ( .A1(n242), .A2(n243), .Z(n238) );
  XOR2D0 U247 ( .A1(n[7]), .A2(n[5]), .Z(n243) );
  XOR2D0 U248 ( .A1(n[9]), .A2(n[8]), .Z(n242) );
  XOR2D0 U249 ( .A1(n244), .A2(n245), .Z(s[1]) );
  XOR2D0 U250 ( .A1(b[1]), .A2(a[1]), .Z(n245) );
  XOR2D0 U251 ( .A1(n[0]), .A2(n246), .Z(n244) );
  XOR2D0 U252 ( .A1(n[2]), .A2(n[1]), .Z(n246) );
  XOR2D0 U253 ( .A1(b[0]), .A2(a[0]), .Z(s[0]) );
endmodule


module gen_nonlinear_part ( a, b, n );
  input [6:0] a;
  input [6:0] b;
  output [245:0] n;
  wire   n_243, n_240, n_239, n_236, n_233, n_232, n_231, n_228, n_225, n_224,
         n_221, n_218, n_217, n_216, n_215, n_212, n_209, n_208, n_205, n_202,
         n_201, n_200, n_197, n_194, n_193, n_190, n_187, n_186, n_185, n_184,
         n_183, n_180, n_177, n_176, n_173, n_170, n_169, n_168, n_165, n_162,
         n_161, n_158, n_155, n_154, n_153, n_152, n_149, n_146, n_145, n_142,
         n_139, n_138, n_137, n_134, n_131, n_130, n_127, n_53, n_50, n_49,
         n_46, n_43, n_42, n_41, n_38, n_35, n_34, n_31, n_28, n_27, n_26,
         n_25, n_22, n_19, n_18, n_15, n_12, n_11, n_10, n_7, n_4, n_3, n_0,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285;
  assign n[243] = n_243;
  assign n[240] = n_240;
  assign n[239] = n_239;
  assign n[236] = n_236;
  assign n[233] = n_233;
  assign n[232] = n_232;
  assign n[231] = n_231;
  assign n[228] = n_228;
  assign n[225] = n_225;
  assign n[224] = n_224;
  assign n[221] = n_221;
  assign n[218] = n_218;
  assign n[217] = n_217;
  assign n[216] = n_216;
  assign n[215] = n_215;
  assign n[212] = n_212;
  assign n[209] = n_209;
  assign n[208] = n_208;
  assign n[205] = n_205;
  assign n[202] = n_202;
  assign n[201] = n_201;
  assign n[200] = n_200;
  assign n[197] = n_197;
  assign n[194] = n_194;
  assign n[193] = n_193;
  assign n[190] = n_190;
  assign n[187] = n_187;
  assign n[186] = n_186;
  assign n[185] = n_185;
  assign n[184] = n_184;
  assign n[183] = n_183;
  assign n[180] = n_180;
  assign n[177] = n_177;
  assign n[176] = n_176;
  assign n[173] = n_173;
  assign n[170] = n_170;
  assign n[169] = n_169;
  assign n[168] = n_168;
  assign n[165] = n_165;
  assign n[162] = n_162;
  assign n[161] = n_161;
  assign n[158] = n_158;
  assign n[155] = n_155;
  assign n[154] = n_154;
  assign n[153] = n_153;
  assign n[152] = n_152;
  assign n[149] = n_149;
  assign n[146] = n_146;
  assign n[145] = n_145;
  assign n[142] = n_142;
  assign n[139] = n_139;
  assign n[138] = n_138;
  assign n[137] = n_137;
  assign n[134] = n_134;
  assign n[131] = n_131;
  assign n[130] = n_130;
  assign n[127] = n_127;
  assign n[53] = n_53;
  assign n[50] = n_50;
  assign n[49] = n_49;
  assign n[46] = n_46;
  assign n[43] = n_43;
  assign n[42] = n_42;
  assign n[41] = n_41;
  assign n[38] = n_38;
  assign n[35] = n_35;
  assign n[34] = n_34;
  assign n[31] = n_31;
  assign n[28] = n_28;
  assign n[27] = n_27;
  assign n[26] = n_26;
  assign n[25] = n_25;
  assign n[22] = n_22;
  assign n[19] = n_19;
  assign n[18] = n_18;
  assign n[15] = n_15;
  assign n[12] = n_12;
  assign n[11] = n_11;
  assign n[10] = n_10;
  assign n[7] = n_7;
  assign n[4] = n_4;
  assign n[3] = n_3;
  assign n[0] = n_0;

  INVD1 U2 ( .I(1'b1), .ZN(n[1]) );
  INVD1 U4 ( .I(1'b1), .ZN(n[2]) );
  INVD1 U6 ( .I(1'b1), .ZN(n[5]) );
  INVD1 U8 ( .I(1'b1), .ZN(n[6]) );
  INVD1 U10 ( .I(1'b1), .ZN(n[8]) );
  INVD1 U12 ( .I(1'b1), .ZN(n[9]) );
  INVD1 U14 ( .I(1'b1), .ZN(n[13]) );
  INVD1 U16 ( .I(1'b1), .ZN(n[14]) );
  INVD1 U18 ( .I(1'b1), .ZN(n[16]) );
  INVD1 U20 ( .I(1'b1), .ZN(n[17]) );
  INVD1 U22 ( .I(1'b1), .ZN(n[20]) );
  INVD1 U24 ( .I(1'b1), .ZN(n[21]) );
  INVD1 U26 ( .I(1'b1), .ZN(n[23]) );
  INVD1 U28 ( .I(1'b1), .ZN(n[24]) );
  INVD1 U30 ( .I(1'b1), .ZN(n[29]) );
  INVD1 U32 ( .I(1'b1), .ZN(n[30]) );
  INVD1 U34 ( .I(1'b1), .ZN(n[32]) );
  INVD1 U36 ( .I(1'b1), .ZN(n[33]) );
  INVD1 U38 ( .I(1'b1), .ZN(n[36]) );
  INVD1 U40 ( .I(1'b1), .ZN(n[37]) );
  INVD1 U42 ( .I(1'b1), .ZN(n[39]) );
  INVD1 U44 ( .I(1'b1), .ZN(n[40]) );
  INVD1 U46 ( .I(1'b1), .ZN(n[44]) );
  INVD1 U48 ( .I(1'b1), .ZN(n[45]) );
  INVD1 U50 ( .I(1'b1), .ZN(n[47]) );
  INVD1 U52 ( .I(1'b1), .ZN(n[48]) );
  INVD1 U54 ( .I(1'b1), .ZN(n[51]) );
  INVD1 U56 ( .I(1'b1), .ZN(n[52]) );
  INVD1 U58 ( .I(1'b1), .ZN(n[54]) );
  INVD1 U60 ( .I(1'b1), .ZN(n[55]) );
  INVD1 U62 ( .I(1'b1), .ZN(n[61]) );
  INVD1 U64 ( .I(1'b1), .ZN(n[62]) );
  INVD1 U66 ( .I(1'b1), .ZN(n[64]) );
  INVD1 U68 ( .I(1'b1), .ZN(n[65]) );
  INVD1 U70 ( .I(1'b1), .ZN(n[68]) );
  INVD1 U72 ( .I(1'b1), .ZN(n[69]) );
  INVD1 U74 ( .I(1'b1), .ZN(n[71]) );
  INVD1 U76 ( .I(1'b1), .ZN(n[72]) );
  INVD1 U78 ( .I(1'b1), .ZN(n[76]) );
  INVD1 U80 ( .I(1'b1), .ZN(n[77]) );
  INVD1 U82 ( .I(1'b1), .ZN(n[79]) );
  INVD1 U84 ( .I(1'b1), .ZN(n[80]) );
  INVD1 U86 ( .I(1'b1), .ZN(n[83]) );
  INVD1 U88 ( .I(1'b1), .ZN(n[84]) );
  INVD1 U90 ( .I(1'b1), .ZN(n[86]) );
  INVD1 U92 ( .I(1'b1), .ZN(n[87]) );
  INVD1 U94 ( .I(1'b1), .ZN(n[92]) );
  INVD1 U96 ( .I(1'b1), .ZN(n[93]) );
  INVD1 U98 ( .I(1'b1), .ZN(n[95]) );
  INVD1 U100 ( .I(1'b1), .ZN(n[96]) );
  INVD1 U102 ( .I(1'b1), .ZN(n[99]) );
  INVD1 U104 ( .I(1'b1), .ZN(n[100]) );
  INVD1 U106 ( .I(1'b1), .ZN(n[102]) );
  INVD1 U108 ( .I(1'b1), .ZN(n[103]) );
  INVD1 U110 ( .I(1'b1), .ZN(n[107]) );
  INVD1 U112 ( .I(1'b1), .ZN(n[108]) );
  INVD1 U114 ( .I(1'b1), .ZN(n[110]) );
  INVD1 U116 ( .I(1'b1), .ZN(n[111]) );
  INVD1 U118 ( .I(1'b1), .ZN(n[114]) );
  INVD1 U120 ( .I(1'b1), .ZN(n[115]) );
  INVD1 U122 ( .I(1'b1), .ZN(n[117]) );
  INVD1 U124 ( .I(1'b1), .ZN(n[118]) );
  INVD1 U126 ( .I(1'b1), .ZN(n[125]) );
  INVD1 U128 ( .I(1'b1), .ZN(n[126]) );
  INVD1 U130 ( .I(1'b1), .ZN(n[128]) );
  INVD1 U132 ( .I(1'b1), .ZN(n[129]) );
  INVD1 U134 ( .I(1'b1), .ZN(n[132]) );
  INVD1 U136 ( .I(1'b1), .ZN(n[133]) );
  INVD1 U138 ( .I(1'b1), .ZN(n[135]) );
  INVD1 U140 ( .I(1'b1), .ZN(n[136]) );
  INVD1 U142 ( .I(1'b1), .ZN(n[140]) );
  INVD1 U144 ( .I(1'b1), .ZN(n[141]) );
  INVD1 U146 ( .I(1'b1), .ZN(n[143]) );
  INVD1 U148 ( .I(1'b1), .ZN(n[144]) );
  INVD1 U150 ( .I(1'b1), .ZN(n[147]) );
  INVD1 U152 ( .I(1'b1), .ZN(n[148]) );
  INVD1 U154 ( .I(1'b1), .ZN(n[150]) );
  INVD1 U156 ( .I(1'b1), .ZN(n[151]) );
  INVD1 U158 ( .I(1'b1), .ZN(n[156]) );
  INVD1 U160 ( .I(1'b1), .ZN(n[157]) );
  INVD1 U162 ( .I(1'b1), .ZN(n[159]) );
  INVD1 U164 ( .I(1'b1), .ZN(n[160]) );
  INVD1 U166 ( .I(1'b1), .ZN(n[163]) );
  INVD1 U168 ( .I(1'b1), .ZN(n[164]) );
  INVD1 U170 ( .I(1'b1), .ZN(n[166]) );
  INVD1 U172 ( .I(1'b1), .ZN(n[167]) );
  INVD1 U174 ( .I(1'b1), .ZN(n[171]) );
  INVD1 U176 ( .I(1'b1), .ZN(n[172]) );
  INVD1 U178 ( .I(1'b1), .ZN(n[174]) );
  INVD1 U180 ( .I(1'b1), .ZN(n[175]) );
  INVD1 U182 ( .I(1'b1), .ZN(n[178]) );
  INVD1 U184 ( .I(1'b1), .ZN(n[179]) );
  INVD1 U186 ( .I(1'b1), .ZN(n[181]) );
  INVD1 U188 ( .I(1'b1), .ZN(n[182]) );
  INVD1 U190 ( .I(1'b1), .ZN(n[188]) );
  INVD1 U192 ( .I(1'b1), .ZN(n[189]) );
  INVD1 U194 ( .I(1'b1), .ZN(n[191]) );
  INVD1 U196 ( .I(1'b1), .ZN(n[192]) );
  INVD1 U198 ( .I(1'b1), .ZN(n[195]) );
  INVD1 U200 ( .I(1'b1), .ZN(n[196]) );
  INVD1 U202 ( .I(1'b1), .ZN(n[198]) );
  INVD1 U204 ( .I(1'b1), .ZN(n[199]) );
  INVD1 U206 ( .I(1'b1), .ZN(n[203]) );
  INVD1 U208 ( .I(1'b1), .ZN(n[204]) );
  INVD1 U210 ( .I(1'b1), .ZN(n[206]) );
  INVD1 U212 ( .I(1'b1), .ZN(n[207]) );
  INVD1 U214 ( .I(1'b1), .ZN(n[210]) );
  INVD1 U216 ( .I(1'b1), .ZN(n[211]) );
  INVD1 U218 ( .I(1'b1), .ZN(n[213]) );
  INVD1 U220 ( .I(1'b1), .ZN(n[214]) );
  INVD1 U222 ( .I(1'b1), .ZN(n[219]) );
  INVD1 U224 ( .I(1'b1), .ZN(n[220]) );
  INVD1 U226 ( .I(1'b1), .ZN(n[222]) );
  INVD1 U228 ( .I(1'b1), .ZN(n[223]) );
  INVD1 U230 ( .I(1'b1), .ZN(n[226]) );
  INVD1 U232 ( .I(1'b1), .ZN(n[227]) );
  INVD1 U234 ( .I(1'b1), .ZN(n[229]) );
  INVD1 U236 ( .I(1'b1), .ZN(n[230]) );
  INVD1 U238 ( .I(1'b1), .ZN(n[234]) );
  INVD1 U240 ( .I(1'b1), .ZN(n[235]) );
  INVD1 U242 ( .I(1'b1), .ZN(n[237]) );
  INVD1 U244 ( .I(1'b1), .ZN(n[238]) );
  INVD1 U246 ( .I(1'b1), .ZN(n[241]) );
  INVD1 U248 ( .I(1'b1), .ZN(n[242]) );
  INVD1 U250 ( .I(1'b1), .ZN(n[244]) );
  INVD1 U252 ( .I(1'b1), .ZN(n[245]) );
  NR2D0 U254 ( .A1(n253), .A2(n254), .ZN(n_243) );
  NR2D0 U255 ( .A1(n254), .A2(n255), .ZN(n_240) );
  NR2D0 U256 ( .A1(n254), .A2(n256), .ZN(n_239) );
  NR2D0 U257 ( .A1(n254), .A2(n257), .ZN(n_236) );
  NR2D0 U258 ( .A1(n254), .A2(n258), .ZN(n_233) );
  NR2D0 U259 ( .A1(n254), .A2(n259), .ZN(n_232) );
  NR2D0 U260 ( .A1(n254), .A2(n260), .ZN(n_231) );
  NR2D0 U261 ( .A1(n254), .A2(n261), .ZN(n_228) );
  NR2D0 U262 ( .A1(n254), .A2(n262), .ZN(n_225) );
  NR2D0 U263 ( .A1(n254), .A2(n263), .ZN(n_224) );
  NR2D0 U264 ( .A1(n254), .A2(n264), .ZN(n_221) );
  NR2D0 U265 ( .A1(n254), .A2(n265), .ZN(n_218) );
  NR2D0 U266 ( .A1(n254), .A2(n266), .ZN(n_217) );
  NR2D0 U267 ( .A1(n254), .A2(n267), .ZN(n_216) );
  NR2D0 U268 ( .A1(n254), .A2(n268), .ZN(n_215) );
  NR2D0 U269 ( .A1(n254), .A2(n269), .ZN(n_212) );
  NR2D0 U270 ( .A1(n254), .A2(n270), .ZN(n_209) );
  NR2D0 U271 ( .A1(n254), .A2(n271), .ZN(n_208) );
  NR2D0 U272 ( .A1(n254), .A2(n272), .ZN(n_205) );
  NR2D0 U273 ( .A1(n254), .A2(n273), .ZN(n_202) );
  NR2D0 U274 ( .A1(n254), .A2(n274), .ZN(n_201) );
  NR2D0 U275 ( .A1(n254), .A2(n275), .ZN(n_200) );
  NR2D0 U276 ( .A1(n254), .A2(n276), .ZN(n_197) );
  NR2D0 U277 ( .A1(n254), .A2(n277), .ZN(n_194) );
  NR2D0 U278 ( .A1(n254), .A2(n278), .ZN(n_193) );
  NR2D0 U279 ( .A1(n254), .A2(n279), .ZN(n_190) );
  NR2D0 U280 ( .A1(n254), .A2(n280), .ZN(n_187) );
  NR2D0 U281 ( .A1(n254), .A2(n281), .ZN(n_186) );
  NR2D0 U282 ( .A1(n254), .A2(n282), .ZN(n_185) );
  NR2D0 U283 ( .A1(n254), .A2(n283), .ZN(n_184) );
  NR2D0 U284 ( .A1(n254), .A2(n284), .ZN(n_183) );
  NR2D0 U285 ( .A1(n253), .A2(n285), .ZN(n_180) );
  NR2D0 U286 ( .A1(n255), .A2(n285), .ZN(n_177) );
  NR2D0 U287 ( .A1(n256), .A2(n285), .ZN(n_176) );
  NR2D0 U288 ( .A1(n257), .A2(n285), .ZN(n_173) );
  NR2D0 U289 ( .A1(n258), .A2(n285), .ZN(n_170) );
  NR2D0 U290 ( .A1(n259), .A2(n285), .ZN(n_169) );
  NR2D0 U291 ( .A1(n260), .A2(n285), .ZN(n_168) );
  NR2D0 U292 ( .A1(n261), .A2(n285), .ZN(n_165) );
  NR2D0 U293 ( .A1(n262), .A2(n285), .ZN(n_162) );
  NR2D0 U294 ( .A1(n263), .A2(n285), .ZN(n_161) );
  NR2D0 U295 ( .A1(n264), .A2(n285), .ZN(n_158) );
  NR2D0 U296 ( .A1(n265), .A2(n285), .ZN(n_155) );
  NR2D0 U297 ( .A1(n266), .A2(n285), .ZN(n_154) );
  NR2D0 U298 ( .A1(n267), .A2(n285), .ZN(n_153) );
  NR2D0 U299 ( .A1(n268), .A2(n285), .ZN(n_152) );
  NR2D0 U300 ( .A1(n269), .A2(n285), .ZN(n_149) );
  NR2D0 U301 ( .A1(n270), .A2(n285), .ZN(n_146) );
  NR2D0 U302 ( .A1(n271), .A2(n285), .ZN(n_145) );
  NR2D0 U303 ( .A1(n272), .A2(n285), .ZN(n_142) );
  NR2D0 U304 ( .A1(n273), .A2(n285), .ZN(n_139) );
  NR2D0 U305 ( .A1(n274), .A2(n285), .ZN(n_138) );
  NR2D0 U306 ( .A1(n275), .A2(n285), .ZN(n_137) );
  NR2D0 U307 ( .A1(n276), .A2(n285), .ZN(n_134) );
  NR2D0 U308 ( .A1(n277), .A2(n285), .ZN(n_131) );
  NR2D0 U309 ( .A1(n278), .A2(n285), .ZN(n_130) );
  NR2D0 U310 ( .A1(n279), .A2(n285), .ZN(n_127) );
  INVD0 U311 ( .I(n262), .ZN(n[98]) );
  ND2D0 U312 ( .A1(n_35), .A2(b[4]), .ZN(n262) );
  INVD0 U313 ( .I(n263), .ZN(n[97]) );
  ND2D0 U314 ( .A1(n_34), .A2(b[4]), .ZN(n263) );
  INVD0 U315 ( .I(n264), .ZN(n[94]) );
  ND2D0 U316 ( .A1(n_31), .A2(b[4]), .ZN(n264) );
  INVD0 U317 ( .I(n265), .ZN(n[91]) );
  ND2D0 U318 ( .A1(n_28), .A2(b[4]), .ZN(n265) );
  INVD0 U319 ( .I(n266), .ZN(n[90]) );
  ND2D0 U320 ( .A1(n_27), .A2(b[4]), .ZN(n266) );
  INVD0 U321 ( .I(n267), .ZN(n[89]) );
  ND2D0 U322 ( .A1(n_26), .A2(b[4]), .ZN(n267) );
  INVD0 U323 ( .I(n268), .ZN(n[88]) );
  ND2D0 U324 ( .A1(n_25), .A2(b[4]), .ZN(n268) );
  INVD0 U325 ( .I(n269), .ZN(n[85]) );
  ND2D0 U326 ( .A1(a[4]), .A2(n_53), .ZN(n269) );
  INVD0 U327 ( .I(n270), .ZN(n[82]) );
  ND2D0 U328 ( .A1(a[4]), .A2(n_50), .ZN(n270) );
  INVD0 U329 ( .I(n271), .ZN(n[81]) );
  ND2D0 U330 ( .A1(a[4]), .A2(n_49), .ZN(n271) );
  INVD0 U331 ( .I(n272), .ZN(n[78]) );
  ND2D0 U332 ( .A1(a[4]), .A2(n_46), .ZN(n272) );
  INVD0 U333 ( .I(n273), .ZN(n[75]) );
  ND2D0 U334 ( .A1(a[4]), .A2(n_43), .ZN(n273) );
  INVD0 U335 ( .I(n274), .ZN(n[74]) );
  ND2D0 U336 ( .A1(a[4]), .A2(n_42), .ZN(n274) );
  INVD0 U337 ( .I(n275), .ZN(n[73]) );
  ND2D0 U338 ( .A1(a[4]), .A2(n_41), .ZN(n275) );
  INVD0 U339 ( .I(n276), .ZN(n[70]) );
  ND2D0 U340 ( .A1(a[4]), .A2(n_38), .ZN(n276) );
  INVD0 U341 ( .I(n277), .ZN(n[67]) );
  ND2D0 U342 ( .A1(a[4]), .A2(n_35), .ZN(n277) );
  AN2D0 U343 ( .A1(a[3]), .A2(n_19), .Z(n_35) );
  INVD0 U344 ( .I(n278), .ZN(n[66]) );
  ND2D0 U345 ( .A1(a[4]), .A2(n_34), .ZN(n278) );
  AN2D0 U346 ( .A1(a[3]), .A2(n_18), .Z(n_34) );
  INVD0 U347 ( .I(n279), .ZN(n[63]) );
  ND2D0 U348 ( .A1(a[4]), .A2(n_31), .ZN(n279) );
  AN2D0 U349 ( .A1(a[3]), .A2(n_15), .Z(n_31) );
  INVD0 U350 ( .I(n280), .ZN(n[60]) );
  INVD0 U351 ( .I(n281), .ZN(n[59]) );
  INVD0 U352 ( .I(n282), .ZN(n[58]) );
  INVD0 U353 ( .I(n283), .ZN(n[57]) );
  INVD0 U354 ( .I(n284), .ZN(n[56]) );
  NR2D0 U355 ( .A1(n280), .A2(n285), .ZN(n[124]) );
  ND2D0 U356 ( .A1(a[4]), .A2(n_28), .ZN(n280) );
  AN2D0 U357 ( .A1(a[3]), .A2(n_12), .Z(n_28) );
  NR2D0 U358 ( .A1(n281), .A2(n285), .ZN(n[123]) );
  ND2D0 U359 ( .A1(a[4]), .A2(n_27), .ZN(n281) );
  AN2D0 U360 ( .A1(a[3]), .A2(n_11), .Z(n_27) );
  NR2D0 U361 ( .A1(n282), .A2(n285), .ZN(n[122]) );
  ND2D0 U362 ( .A1(a[4]), .A2(n_26), .ZN(n282) );
  AN2D0 U363 ( .A1(a[3]), .A2(n_10), .Z(n_26) );
  NR2D0 U364 ( .A1(n283), .A2(n285), .ZN(n[121]) );
  ND2D0 U365 ( .A1(a[4]), .A2(n_25), .ZN(n283) );
  AN2D0 U366 ( .A1(a[3]), .A2(b[3]), .Z(n_25) );
  NR2D0 U367 ( .A1(n284), .A2(n285), .ZN(n[120]) );
  ND2D0 U368 ( .A1(a[4]), .A2(b[4]), .ZN(n284) );
  NR2D0 U369 ( .A1(n254), .A2(n285), .ZN(n[119]) );
  INVD0 U370 ( .I(a[5]), .ZN(n285) );
  INVD0 U371 ( .I(b[5]), .ZN(n254) );
  INVD0 U372 ( .I(n253), .ZN(n[116]) );
  ND2D0 U373 ( .A1(b[4]), .A2(n_53), .ZN(n253) );
  AN2D0 U374 ( .A1(b[3]), .A2(n_22), .Z(n_53) );
  INVD0 U375 ( .I(n255), .ZN(n[113]) );
  ND2D0 U376 ( .A1(n_50), .A2(b[4]), .ZN(n255) );
  AN2D0 U377 ( .A1(n_19), .A2(b[3]), .Z(n_50) );
  AN2D0 U378 ( .A1(n_4), .A2(b[2]), .Z(n_19) );
  INVD0 U379 ( .I(n256), .ZN(n[112]) );
  ND2D0 U380 ( .A1(n_49), .A2(b[4]), .ZN(n256) );
  AN2D0 U381 ( .A1(n_18), .A2(b[3]), .Z(n_49) );
  AN2D0 U382 ( .A1(n_3), .A2(b[2]), .Z(n_18) );
  INVD0 U383 ( .I(n257), .ZN(n[109]) );
  ND2D0 U384 ( .A1(n_46), .A2(b[4]), .ZN(n257) );
  AN2D0 U385 ( .A1(n_15), .A2(b[3]), .Z(n_46) );
  AN2D0 U386 ( .A1(a[2]), .A2(n_7), .Z(n_15) );
  INVD0 U387 ( .I(n258), .ZN(n[106]) );
  ND2D0 U388 ( .A1(n_43), .A2(b[4]), .ZN(n258) );
  AN2D0 U389 ( .A1(n_12), .A2(b[3]), .Z(n_43) );
  AN2D0 U390 ( .A1(a[2]), .A2(n_4), .Z(n_12) );
  AN2D0 U391 ( .A1(a[1]), .A2(n_0), .Z(n_4) );
  INVD0 U392 ( .I(n259), .ZN(n[105]) );
  ND2D0 U393 ( .A1(n_42), .A2(b[4]), .ZN(n259) );
  AN2D0 U394 ( .A1(n_11), .A2(b[3]), .Z(n_42) );
  AN2D0 U395 ( .A1(a[2]), .A2(n_3), .Z(n_11) );
  AN2D0 U396 ( .A1(a[1]), .A2(b[1]), .Z(n_3) );
  INVD0 U397 ( .I(n260), .ZN(n[104]) );
  ND2D0 U398 ( .A1(n_41), .A2(b[4]), .ZN(n260) );
  AN2D0 U399 ( .A1(n_10), .A2(b[3]), .Z(n_41) );
  AN2D0 U400 ( .A1(a[2]), .A2(b[2]), .Z(n_10) );
  INVD0 U401 ( .I(n261), .ZN(n[101]) );
  ND2D0 U402 ( .A1(n_38), .A2(b[4]), .ZN(n261) );
  AN2D0 U403 ( .A1(a[3]), .A2(n_22), .Z(n_38) );
  AN2D0 U404 ( .A1(b[2]), .A2(n_7), .Z(n_22) );
  AN2D0 U405 ( .A1(b[1]), .A2(n_0), .Z(n_7) );
  AN2D0 U406 ( .A1(b[0]), .A2(a[0]), .Z(n_0) );
endmodule


module gen_cla_decomposed ( a, b, s );
  input [6:0] a;
  input [6:0] b;
  output [6:0] s;

  wire   [245:0] n;

  gen_nonlinear_part NLIN ( .a(a), .b(b), .n(n) );
  gen_linear_part LIN ( .a(a), .b(b), .n({1'b0, 1'b0, n[243], 1'b0, 1'b0, 
        n[240:239], 1'b0, 1'b0, n[236], 1'b0, 1'b0, n[233:231], 1'b0, 1'b0, 
        n[228], 1'b0, 1'b0, n[225:224], 1'b0, 1'b0, n[221], 1'b0, 1'b0, 
        n[218:215], 1'b0, 1'b0, n[212], 1'b0, 1'b0, n[209:208], 1'b0, 1'b0, 
        n[205], 1'b0, 1'b0, n[202:200], 1'b0, 1'b0, n[197], 1'b0, 1'b0, 
        n[194:193], 1'b0, 1'b0, n[190], 1'b0, 1'b0, n[187:183], 1'b0, 1'b0, 
        n[180], 1'b0, 1'b0, n[177:176], 1'b0, 1'b0, n[173], 1'b0, 1'b0, 
        n[170:168], 1'b0, 1'b0, n[165], 1'b0, 1'b0, n[162:161], 1'b0, 1'b0, 
        n[158], 1'b0, 1'b0, n[155:152], 1'b0, 1'b0, n[149], 1'b0, 1'b0, 
        n[146:145], 1'b0, 1'b0, n[142], 1'b0, 1'b0, n[139:137], 1'b0, 1'b0, 
        n[134], 1'b0, 1'b0, n[131:130], 1'b0, 1'b0, n[127], 1'b0, 1'b0, 
        n[124:119], 1'b0, 1'b0, n[116], 1'b0, 1'b0, n[113:112], 1'b0, 1'b0, 
        n[109], 1'b0, 1'b0, n[106:104], 1'b0, 1'b0, n[101], 1'b0, 1'b0, 
        n[98:97], 1'b0, 1'b0, n[94], 1'b0, 1'b0, n[91:88], 1'b0, 1'b0, n[85], 
        1'b0, 1'b0, n[82:81], 1'b0, 1'b0, n[78], 1'b0, 1'b0, n[75:73], 1'b0, 
        1'b0, n[70], 1'b0, 1'b0, n[67:66], 1'b0, 1'b0, n[63], 1'b0, 1'b0, 
        n[60:56], 1'b0, 1'b0, n[53], 1'b0, 1'b0, n[50:49], 1'b0, 1'b0, n[46], 
        1'b0, 1'b0, n[43:41], 1'b0, 1'b0, n[38], 1'b0, 1'b0, n[35:34], 1'b0, 
        1'b0, n[31], 1'b0, 1'b0, n[28:25], 1'b0, 1'b0, n[22], 1'b0, 1'b0, 
        n[19:18], 1'b0, 1'b0, n[15], 1'b0, 1'b0, n[12:10], 1'b0, 1'b0, n[7], 
        1'b0, 1'b0, n[4:3], 1'b0, 1'b0, n[0]}), .s(s) );
endmodule

