
module gen_linear_part ( a, b, n, s );
  input [10:0] a;
  input [10:0] b;
  input [4081:0] n;
  output [10:0] s;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455;

  XOR4D0 U1 ( .A1(b[9]), .A2(a[9]), .A3(n1), .A4(n2), .Z(s[9]) );
  XOR4D0 U2 ( .A1(n[2028]), .A2(n3), .A3(n[2030]), .A4(n[2029]), .Z(n2) );
  XOR4D0 U3 ( .A1(n[2023]), .A2(n[2022]), .A3(n4), .A4(n5), .Z(n3) );
  XOR3D0 U4 ( .A1(n6), .A2(n7), .A3(n[2021]), .Z(n5) );
  XOR4D0 U5 ( .A1(n[2014]), .A2(n8), .A3(n[2016]), .A4(n[2015]), .Z(n7) );
  XOR4D0 U6 ( .A1(n[2009]), .A2(n[2008]), .A3(n9), .A4(n10), .Z(n8) );
  XOR3D0 U7 ( .A1(n11), .A2(n12), .A3(n[2007]), .Z(n10) );
  XOR4D0 U8 ( .A1(n[2000]), .A2(n13), .A3(n[2002]), .A4(n[2001]), .Z(n12) );
  XOR4D0 U9 ( .A1(n[1995]), .A2(n[1994]), .A3(n14), .A4(n15), .Z(n13) );
  XOR3D0 U10 ( .A1(n16), .A2(n17), .A3(n[1993]), .Z(n15) );
  XOR4D0 U11 ( .A1(n[1986]), .A2(n18), .A3(n[1988]), .A4(n[1987]), .Z(n17) );
  XOR4D0 U12 ( .A1(n[1981]), .A2(n[1980]), .A3(n19), .A4(n20), .Z(n18) );
  XOR3D0 U13 ( .A1(n21), .A2(n22), .A3(n[1979]), .Z(n20) );
  XOR4D0 U14 ( .A1(n[1972]), .A2(n23), .A3(n[1974]), .A4(n[1973]), .Z(n22) );
  XOR4D0 U15 ( .A1(n[1967]), .A2(n[1966]), .A3(n24), .A4(n25), .Z(n23) );
  XOR3D0 U16 ( .A1(n26), .A2(n27), .A3(n[1965]), .Z(n25) );
  XOR4D0 U17 ( .A1(n[1958]), .A2(n28), .A3(n[1960]), .A4(n[1959]), .Z(n27) );
  XOR4D0 U18 ( .A1(n[1953]), .A2(n[1952]), .A3(n29), .A4(n30), .Z(n28) );
  XOR3D0 U19 ( .A1(n31), .A2(n32), .A3(n[1951]), .Z(n30) );
  XOR4D0 U20 ( .A1(n[1944]), .A2(n33), .A3(n[1946]), .A4(n[1945]), .Z(n32) );
  XOR4D0 U21 ( .A1(n[1939]), .A2(n[1938]), .A3(n34), .A4(n35), .Z(n33) );
  XOR3D0 U22 ( .A1(n36), .A2(n37), .A3(n[1937]), .Z(n35) );
  XOR4D0 U23 ( .A1(n[1930]), .A2(n38), .A3(n[1932]), .A4(n[1931]), .Z(n37) );
  XOR4D0 U24 ( .A1(n[1925]), .A2(n[1924]), .A3(n39), .A4(n40), .Z(n38) );
  XOR3D0 U25 ( .A1(n41), .A2(n42), .A3(n[1923]), .Z(n40) );
  XOR4D0 U26 ( .A1(n[1916]), .A2(n43), .A3(n[1918]), .A4(n[1917]), .Z(n42) );
  XOR4D0 U27 ( .A1(n[1911]), .A2(n[1910]), .A3(n44), .A4(n45), .Z(n43) );
  XOR3D0 U28 ( .A1(n46), .A2(n47), .A3(n[1909]), .Z(n45) );
  XOR4D0 U29 ( .A1(n[1902]), .A2(n48), .A3(n[1904]), .A4(n[1903]), .Z(n47) );
  XOR4D0 U30 ( .A1(n[1897]), .A2(n[1896]), .A3(n49), .A4(n50), .Z(n48) );
  XOR3D0 U31 ( .A1(n51), .A2(n52), .A3(n[1895]), .Z(n50) );
  XOR4D0 U32 ( .A1(n[1888]), .A2(n53), .A3(n[1890]), .A4(n[1889]), .Z(n52) );
  XOR4D0 U33 ( .A1(n[1883]), .A2(n[1882]), .A3(n54), .A4(n55), .Z(n53) );
  XOR3D0 U34 ( .A1(n56), .A2(n57), .A3(n[1881]), .Z(n55) );
  XOR4D0 U35 ( .A1(n[1874]), .A2(n58), .A3(n[1876]), .A4(n[1875]), .Z(n57) );
  XOR4D0 U36 ( .A1(n[1869]), .A2(n[1868]), .A3(n59), .A4(n60), .Z(n58) );
  XOR3D0 U37 ( .A1(n61), .A2(n62), .A3(n[1867]), .Z(n60) );
  XOR4D0 U38 ( .A1(n[1860]), .A2(n63), .A3(n[1862]), .A4(n[1861]), .Z(n62) );
  XOR4D0 U39 ( .A1(n[1855]), .A2(n[1854]), .A3(n64), .A4(n65), .Z(n63) );
  XOR3D0 U40 ( .A1(n66), .A2(n67), .A3(n[1853]), .Z(n65) );
  XOR4D0 U41 ( .A1(n[1846]), .A2(n68), .A3(n[1848]), .A4(n[1847]), .Z(n67) );
  XOR4D0 U42 ( .A1(n[1841]), .A2(n[1840]), .A3(n69), .A4(n70), .Z(n68) );
  XOR3D0 U43 ( .A1(n71), .A2(n72), .A3(n[1839]), .Z(n70) );
  XOR4D0 U44 ( .A1(n[1832]), .A2(n73), .A3(n[1834]), .A4(n[1833]), .Z(n72) );
  XOR4D0 U45 ( .A1(n[1827]), .A2(n[1826]), .A3(n74), .A4(n75), .Z(n73) );
  XOR3D0 U46 ( .A1(n76), .A2(n77), .A3(n[1825]), .Z(n75) );
  XOR4D0 U47 ( .A1(n[1818]), .A2(n78), .A3(n[1820]), .A4(n[1819]), .Z(n77) );
  XOR4D0 U48 ( .A1(n[1813]), .A2(n[1812]), .A3(n79), .A4(n80), .Z(n78) );
  XOR3D0 U49 ( .A1(n81), .A2(n82), .A3(n[1811]), .Z(n80) );
  XOR4D0 U50 ( .A1(n[1804]), .A2(n83), .A3(n[1806]), .A4(n[1805]), .Z(n82) );
  XOR4D0 U51 ( .A1(n[1799]), .A2(n[1798]), .A3(n84), .A4(n85), .Z(n83) );
  XOR3D0 U52 ( .A1(n86), .A2(n87), .A3(n[1797]), .Z(n85) );
  XOR4D0 U53 ( .A1(n[1790]), .A2(n88), .A3(n[1792]), .A4(n[1791]), .Z(n87) );
  XOR4D0 U54 ( .A1(n[1785]), .A2(n[1784]), .A3(n89), .A4(n90), .Z(n88) );
  XOR3D0 U55 ( .A1(n91), .A2(n92), .A3(n[1783]), .Z(n90) );
  XOR4D0 U56 ( .A1(n[1776]), .A2(n93), .A3(n[1778]), .A4(n[1777]), .Z(n92) );
  XOR4D0 U57 ( .A1(n[1771]), .A2(n[1770]), .A3(n94), .A4(n95), .Z(n93) );
  XOR3D0 U58 ( .A1(n96), .A2(n97), .A3(n[1769]), .Z(n95) );
  XOR4D0 U59 ( .A1(n[1762]), .A2(n98), .A3(n[1764]), .A4(n[1763]), .Z(n97) );
  XOR4D0 U60 ( .A1(n[1757]), .A2(n[1756]), .A3(n99), .A4(n100), .Z(n98) );
  XOR3D0 U61 ( .A1(n101), .A2(n102), .A3(n[1755]), .Z(n100) );
  XOR4D0 U62 ( .A1(n[1748]), .A2(n103), .A3(n[1750]), .A4(n[1749]), .Z(n102)
         );
  XOR4D0 U63 ( .A1(n[1743]), .A2(n[1742]), .A3(n104), .A4(n105), .Z(n103) );
  XOR3D0 U64 ( .A1(n106), .A2(n107), .A3(n[1741]), .Z(n105) );
  XOR4D0 U65 ( .A1(n[1734]), .A2(n108), .A3(n[1736]), .A4(n[1735]), .Z(n107)
         );
  XOR4D0 U66 ( .A1(n[1729]), .A2(n[1728]), .A3(n109), .A4(n110), .Z(n108) );
  XOR3D0 U67 ( .A1(n111), .A2(n112), .A3(n[1727]), .Z(n110) );
  XOR4D0 U68 ( .A1(n[1720]), .A2(n113), .A3(n[1722]), .A4(n[1721]), .Z(n112)
         );
  XOR4D0 U69 ( .A1(n[1715]), .A2(n[1714]), .A3(n114), .A4(n115), .Z(n113) );
  XOR3D0 U70 ( .A1(n116), .A2(n117), .A3(n[1713]), .Z(n115) );
  XOR4D0 U71 ( .A1(n[1706]), .A2(n118), .A3(n[1708]), .A4(n[1707]), .Z(n117)
         );
  XOR4D0 U72 ( .A1(n[1701]), .A2(n[1700]), .A3(n119), .A4(n120), .Z(n118) );
  XOR3D0 U73 ( .A1(n121), .A2(n122), .A3(n[1699]), .Z(n120) );
  XOR4D0 U74 ( .A1(n[1692]), .A2(n123), .A3(n[1694]), .A4(n[1693]), .Z(n122)
         );
  XOR4D0 U75 ( .A1(n[1687]), .A2(n[1686]), .A3(n124), .A4(n125), .Z(n123) );
  XOR3D0 U76 ( .A1(n126), .A2(n127), .A3(n[1685]), .Z(n125) );
  XOR4D0 U77 ( .A1(n[1678]), .A2(n128), .A3(n[1680]), .A4(n[1679]), .Z(n127)
         );
  XOR4D0 U78 ( .A1(n[1673]), .A2(n[1672]), .A3(n129), .A4(n130), .Z(n128) );
  XOR3D0 U79 ( .A1(n131), .A2(n132), .A3(n[1671]), .Z(n130) );
  XOR4D0 U80 ( .A1(n[1664]), .A2(n133), .A3(n[1666]), .A4(n[1665]), .Z(n132)
         );
  XOR4D0 U81 ( .A1(n[1659]), .A2(n[1658]), .A3(n134), .A4(n135), .Z(n133) );
  XOR3D0 U82 ( .A1(n136), .A2(n137), .A3(n[1657]), .Z(n135) );
  XOR4D0 U83 ( .A1(n[1650]), .A2(n138), .A3(n[1652]), .A4(n[1651]), .Z(n137)
         );
  XOR4D0 U84 ( .A1(n[1645]), .A2(n[1644]), .A3(n139), .A4(n140), .Z(n138) );
  XOR3D0 U85 ( .A1(n141), .A2(n142), .A3(n[1643]), .Z(n140) );
  XOR4D0 U86 ( .A1(n[1636]), .A2(n143), .A3(n[1638]), .A4(n[1637]), .Z(n142)
         );
  XOR4D0 U87 ( .A1(n[1631]), .A2(n[1630]), .A3(n144), .A4(n145), .Z(n143) );
  XOR3D0 U88 ( .A1(n146), .A2(n147), .A3(n[1629]), .Z(n145) );
  XOR4D0 U89 ( .A1(n[1622]), .A2(n148), .A3(n[1624]), .A4(n[1623]), .Z(n147)
         );
  XOR4D0 U90 ( .A1(n[1617]), .A2(n[1616]), .A3(n149), .A4(n150), .Z(n148) );
  XOR3D0 U91 ( .A1(n151), .A2(n152), .A3(n[1615]), .Z(n150) );
  XOR4D0 U92 ( .A1(n[1608]), .A2(n153), .A3(n[1610]), .A4(n[1609]), .Z(n152)
         );
  XOR4D0 U93 ( .A1(n[1603]), .A2(n[1602]), .A3(n154), .A4(n155), .Z(n153) );
  XOR3D0 U94 ( .A1(n156), .A2(n157), .A3(n[1601]), .Z(n155) );
  XOR4D0 U95 ( .A1(n[1594]), .A2(n158), .A3(n[1596]), .A4(n[1595]), .Z(n157)
         );
  XOR4D0 U96 ( .A1(n[1589]), .A2(n[1588]), .A3(n159), .A4(n160), .Z(n158) );
  XOR3D0 U97 ( .A1(n161), .A2(n162), .A3(n[1587]), .Z(n160) );
  XOR4D0 U98 ( .A1(n[1580]), .A2(n163), .A3(n[1582]), .A4(n[1581]), .Z(n162)
         );
  XOR4D0 U99 ( .A1(n[1575]), .A2(n[1574]), .A3(n164), .A4(n165), .Z(n163) );
  XOR3D0 U100 ( .A1(n166), .A2(n167), .A3(n[1573]), .Z(n165) );
  XOR4D0 U101 ( .A1(n[1566]), .A2(n168), .A3(n[1568]), .A4(n[1567]), .Z(n167)
         );
  XOR4D0 U102 ( .A1(n[1561]), .A2(n[1560]), .A3(n169), .A4(n170), .Z(n168) );
  XOR3D0 U103 ( .A1(n171), .A2(n172), .A3(n[1559]), .Z(n170) );
  XOR4D0 U104 ( .A1(n[1552]), .A2(n173), .A3(n[1554]), .A4(n[1553]), .Z(n172)
         );
  XOR4D0 U105 ( .A1(n[1547]), .A2(n[1546]), .A3(n174), .A4(n175), .Z(n173) );
  XOR3D0 U106 ( .A1(n176), .A2(n177), .A3(n[1545]), .Z(n175) );
  XOR4D0 U107 ( .A1(n[1538]), .A2(n178), .A3(n[1540]), .A4(n[1539]), .Z(n177)
         );
  XOR4D0 U108 ( .A1(n[1533]), .A2(n[1532]), .A3(n179), .A4(n180), .Z(n178) );
  XOR3D0 U109 ( .A1(n181), .A2(n182), .A3(n[1531]), .Z(n180) );
  XOR4D0 U110 ( .A1(n[1524]), .A2(n183), .A3(n[1526]), .A4(n[1525]), .Z(n182)
         );
  XOR4D0 U111 ( .A1(n[1519]), .A2(n[1518]), .A3(n184), .A4(n185), .Z(n183) );
  XOR3D0 U112 ( .A1(n186), .A2(n187), .A3(n[1517]), .Z(n185) );
  XOR4D0 U113 ( .A1(n[1510]), .A2(n188), .A3(n[1512]), .A4(n[1511]), .Z(n187)
         );
  XOR4D0 U114 ( .A1(n[1505]), .A2(n[1504]), .A3(n189), .A4(n190), .Z(n188) );
  XOR3D0 U115 ( .A1(n191), .A2(n192), .A3(n[1503]), .Z(n190) );
  XOR4D0 U116 ( .A1(n[1496]), .A2(n193), .A3(n[1498]), .A4(n[1497]), .Z(n192)
         );
  XOR4D0 U117 ( .A1(n[1491]), .A2(n[1490]), .A3(n194), .A4(n195), .Z(n193) );
  XOR3D0 U118 ( .A1(n196), .A2(n197), .A3(n[1489]), .Z(n195) );
  XOR4D0 U119 ( .A1(n[1482]), .A2(n198), .A3(n[1484]), .A4(n[1483]), .Z(n197)
         );
  XOR4D0 U120 ( .A1(n[1477]), .A2(n[1476]), .A3(n199), .A4(n200), .Z(n198) );
  XOR3D0 U121 ( .A1(n201), .A2(n202), .A3(n[1475]), .Z(n200) );
  XOR4D0 U122 ( .A1(n[1468]), .A2(n203), .A3(n[1470]), .A4(n[1469]), .Z(n202)
         );
  XOR4D0 U123 ( .A1(n[1463]), .A2(n[1462]), .A3(n204), .A4(n205), .Z(n203) );
  XOR3D0 U124 ( .A1(n206), .A2(n207), .A3(n[1461]), .Z(n205) );
  XOR4D0 U125 ( .A1(n[1454]), .A2(n208), .A3(n[1456]), .A4(n[1455]), .Z(n207)
         );
  XOR4D0 U126 ( .A1(n[1449]), .A2(n[1448]), .A3(n209), .A4(n210), .Z(n208) );
  XOR3D0 U127 ( .A1(n211), .A2(n212), .A3(n[1447]), .Z(n210) );
  XOR4D0 U128 ( .A1(n[1440]), .A2(n213), .A3(n[1442]), .A4(n[1441]), .Z(n212)
         );
  XOR4D0 U129 ( .A1(n[1435]), .A2(n[1434]), .A3(n214), .A4(n215), .Z(n213) );
  XOR3D0 U130 ( .A1(n216), .A2(n217), .A3(n[1433]), .Z(n215) );
  XOR4D0 U131 ( .A1(n[1426]), .A2(n218), .A3(n[1428]), .A4(n[1427]), .Z(n217)
         );
  XOR4D0 U132 ( .A1(n[1421]), .A2(n[1420]), .A3(n219), .A4(n220), .Z(n218) );
  XOR3D0 U133 ( .A1(n221), .A2(n222), .A3(n[1419]), .Z(n220) );
  XOR4D0 U134 ( .A1(n[1412]), .A2(n223), .A3(n[1414]), .A4(n[1413]), .Z(n222)
         );
  XOR4D0 U135 ( .A1(n[1407]), .A2(n[1406]), .A3(n224), .A4(n225), .Z(n223) );
  XOR3D0 U136 ( .A1(n226), .A2(n227), .A3(n[1405]), .Z(n225) );
  XOR4D0 U137 ( .A1(n[1398]), .A2(n228), .A3(n[1400]), .A4(n[1399]), .Z(n227)
         );
  XOR4D0 U138 ( .A1(n[1393]), .A2(n[1392]), .A3(n229), .A4(n230), .Z(n228) );
  XOR3D0 U139 ( .A1(n231), .A2(n232), .A3(n[1391]), .Z(n230) );
  XOR4D0 U140 ( .A1(n[1384]), .A2(n233), .A3(n[1386]), .A4(n[1385]), .Z(n232)
         );
  XOR4D0 U141 ( .A1(n[1379]), .A2(n[1378]), .A3(n234), .A4(n235), .Z(n233) );
  XOR3D0 U142 ( .A1(n236), .A2(n237), .A3(n[1377]), .Z(n235) );
  XOR4D0 U143 ( .A1(n[1370]), .A2(n238), .A3(n[1372]), .A4(n[1371]), .Z(n237)
         );
  XOR4D0 U144 ( .A1(n[1365]), .A2(n[1364]), .A3(n239), .A4(n240), .Z(n238) );
  XOR3D0 U145 ( .A1(n241), .A2(n242), .A3(n[1363]), .Z(n240) );
  XOR4D0 U146 ( .A1(n[1356]), .A2(n243), .A3(n[1358]), .A4(n[1357]), .Z(n242)
         );
  XOR4D0 U147 ( .A1(n[1351]), .A2(n[1350]), .A3(n244), .A4(n245), .Z(n243) );
  XOR3D0 U148 ( .A1(n246), .A2(n247), .A3(n[1349]), .Z(n245) );
  XOR4D0 U149 ( .A1(n[1342]), .A2(n248), .A3(n[1344]), .A4(n[1343]), .Z(n247)
         );
  XOR4D0 U150 ( .A1(n[1337]), .A2(n[1336]), .A3(n249), .A4(n250), .Z(n248) );
  XOR3D0 U151 ( .A1(n251), .A2(n252), .A3(n[1335]), .Z(n250) );
  XOR4D0 U152 ( .A1(n[1328]), .A2(n253), .A3(n[1330]), .A4(n[1329]), .Z(n252)
         );
  XOR4D0 U153 ( .A1(n[1323]), .A2(n[1322]), .A3(n254), .A4(n255), .Z(n253) );
  XOR3D0 U154 ( .A1(n256), .A2(n257), .A3(n[1321]), .Z(n255) );
  XOR4D0 U155 ( .A1(n[1314]), .A2(n258), .A3(n[1316]), .A4(n[1315]), .Z(n257)
         );
  XOR4D0 U156 ( .A1(n[1309]), .A2(n[1308]), .A3(n259), .A4(n260), .Z(n258) );
  XOR3D0 U157 ( .A1(n261), .A2(n262), .A3(n[1307]), .Z(n260) );
  XOR4D0 U158 ( .A1(n[1300]), .A2(n263), .A3(n[1302]), .A4(n[1301]), .Z(n262)
         );
  XOR4D0 U159 ( .A1(n[1295]), .A2(n[1294]), .A3(n264), .A4(n265), .Z(n263) );
  XOR3D0 U160 ( .A1(n266), .A2(n267), .A3(n[1293]), .Z(n265) );
  XOR4D0 U161 ( .A1(n[1286]), .A2(n268), .A3(n[1288]), .A4(n[1287]), .Z(n267)
         );
  XOR4D0 U162 ( .A1(n[1281]), .A2(n[1280]), .A3(n269), .A4(n270), .Z(n268) );
  XOR3D0 U163 ( .A1(n271), .A2(n272), .A3(n[1279]), .Z(n270) );
  XOR4D0 U164 ( .A1(n[1272]), .A2(n273), .A3(n[1274]), .A4(n[1273]), .Z(n272)
         );
  XOR4D0 U165 ( .A1(n[1267]), .A2(n[1266]), .A3(n274), .A4(n275), .Z(n273) );
  XOR3D0 U166 ( .A1(n276), .A2(n277), .A3(n[1265]), .Z(n275) );
  XOR4D0 U167 ( .A1(n[1258]), .A2(n278), .A3(n[1260]), .A4(n[1259]), .Z(n277)
         );
  XOR4D0 U168 ( .A1(n[1253]), .A2(n[1252]), .A3(n279), .A4(n280), .Z(n278) );
  XOR3D0 U169 ( .A1(n281), .A2(n282), .A3(n[1251]), .Z(n280) );
  XOR4D0 U170 ( .A1(n[1244]), .A2(n283), .A3(n[1246]), .A4(n[1245]), .Z(n282)
         );
  XOR4D0 U171 ( .A1(n[1239]), .A2(n[1238]), .A3(n284), .A4(n285), .Z(n283) );
  XOR3D0 U172 ( .A1(n286), .A2(n287), .A3(n[1237]), .Z(n285) );
  XOR4D0 U173 ( .A1(n[1230]), .A2(n288), .A3(n[1232]), .A4(n[1231]), .Z(n287)
         );
  XOR4D0 U174 ( .A1(n[1225]), .A2(n[1224]), .A3(n289), .A4(n290), .Z(n288) );
  XOR3D0 U175 ( .A1(n291), .A2(n292), .A3(n[1223]), .Z(n290) );
  XOR4D0 U176 ( .A1(n[1216]), .A2(n293), .A3(n[1218]), .A4(n[1217]), .Z(n292)
         );
  XOR4D0 U177 ( .A1(n[1211]), .A2(n[1210]), .A3(n294), .A4(n295), .Z(n293) );
  XOR3D0 U178 ( .A1(n296), .A2(n297), .A3(n[1209]), .Z(n295) );
  XOR4D0 U179 ( .A1(n[1202]), .A2(n298), .A3(n[1204]), .A4(n[1203]), .Z(n297)
         );
  XOR4D0 U180 ( .A1(n[1197]), .A2(n[1196]), .A3(n299), .A4(n300), .Z(n298) );
  XOR3D0 U181 ( .A1(n301), .A2(n302), .A3(n[1195]), .Z(n300) );
  XOR4D0 U182 ( .A1(n[1188]), .A2(n303), .A3(n[1190]), .A4(n[1189]), .Z(n302)
         );
  XOR4D0 U183 ( .A1(n[1183]), .A2(n[1182]), .A3(n304), .A4(n305), .Z(n303) );
  XOR3D0 U184 ( .A1(n306), .A2(n307), .A3(n[1181]), .Z(n305) );
  XOR4D0 U185 ( .A1(n[1174]), .A2(n308), .A3(n[1176]), .A4(n[1175]), .Z(n307)
         );
  XOR4D0 U186 ( .A1(n[1169]), .A2(n[1168]), .A3(n309), .A4(n310), .Z(n308) );
  XOR3D0 U187 ( .A1(n311), .A2(n312), .A3(n[1167]), .Z(n310) );
  XOR4D0 U188 ( .A1(n[1160]), .A2(n313), .A3(n[1162]), .A4(n[1161]), .Z(n312)
         );
  XOR4D0 U189 ( .A1(n[1155]), .A2(n[1154]), .A3(n314), .A4(n315), .Z(n313) );
  XOR3D0 U190 ( .A1(n316), .A2(n317), .A3(n[1153]), .Z(n315) );
  XOR4D0 U191 ( .A1(n[1146]), .A2(n318), .A3(n[1148]), .A4(n[1147]), .Z(n317)
         );
  XOR4D0 U192 ( .A1(n[1141]), .A2(n[1140]), .A3(n319), .A4(n320), .Z(n318) );
  XOR3D0 U193 ( .A1(n321), .A2(n322), .A3(n[1139]), .Z(n320) );
  XOR4D0 U194 ( .A1(n[1132]), .A2(n323), .A3(n[1134]), .A4(n[1133]), .Z(n322)
         );
  XOR4D0 U195 ( .A1(n[1127]), .A2(n[1126]), .A3(n324), .A4(n325), .Z(n323) );
  XOR3D0 U196 ( .A1(n326), .A2(n327), .A3(n[1125]), .Z(n325) );
  XOR4D0 U197 ( .A1(n[1118]), .A2(n328), .A3(n[1120]), .A4(n[1119]), .Z(n327)
         );
  XOR4D0 U198 ( .A1(n[1113]), .A2(n[1112]), .A3(n329), .A4(n330), .Z(n328) );
  XOR3D0 U199 ( .A1(n331), .A2(n332), .A3(n[1111]), .Z(n330) );
  XOR4D0 U200 ( .A1(n[1104]), .A2(n333), .A3(n[1106]), .A4(n[1105]), .Z(n332)
         );
  XOR4D0 U201 ( .A1(n[1099]), .A2(n[1098]), .A3(n334), .A4(n335), .Z(n333) );
  XOR3D0 U202 ( .A1(n336), .A2(n337), .A3(n[1097]), .Z(n335) );
  XOR4D0 U203 ( .A1(n[1090]), .A2(n338), .A3(n[1092]), .A4(n[1091]), .Z(n337)
         );
  XOR4D0 U204 ( .A1(n[1085]), .A2(n[1084]), .A3(n339), .A4(n340), .Z(n338) );
  XOR3D0 U205 ( .A1(n341), .A2(n342), .A3(n[1083]), .Z(n340) );
  XOR4D0 U206 ( .A1(n[1076]), .A2(n343), .A3(n[1078]), .A4(n[1077]), .Z(n342)
         );
  XOR4D0 U207 ( .A1(n[1071]), .A2(n[1070]), .A3(n344), .A4(n345), .Z(n343) );
  XOR3D0 U208 ( .A1(n346), .A2(n347), .A3(n[1069]), .Z(n345) );
  XOR4D0 U209 ( .A1(n[1062]), .A2(n348), .A3(n[1064]), .A4(n[1063]), .Z(n347)
         );
  XOR4D0 U210 ( .A1(n[1057]), .A2(n[1056]), .A3(n349), .A4(n350), .Z(n348) );
  XOR3D0 U211 ( .A1(n351), .A2(n352), .A3(n[1055]), .Z(n350) );
  XOR4D0 U212 ( .A1(n[1048]), .A2(n353), .A3(n[1050]), .A4(n[1049]), .Z(n352)
         );
  XOR4D0 U213 ( .A1(n[1043]), .A2(n[1042]), .A3(n354), .A4(n355), .Z(n353) );
  XOR3D0 U214 ( .A1(n356), .A2(n357), .A3(n[1041]), .Z(n355) );
  XOR4D0 U215 ( .A1(n[1034]), .A2(n358), .A3(n[1036]), .A4(n[1035]), .Z(n357)
         );
  XOR4D0 U216 ( .A1(n[1029]), .A2(n[1028]), .A3(n359), .A4(n360), .Z(n358) );
  XOR3D0 U217 ( .A1(n361), .A2(n362), .A3(n[1027]), .Z(n360) );
  XOR3D0 U218 ( .A1(n[1022]), .A2(n[1021]), .A3(n363), .Z(n362) );
  XOR3D0 U219 ( .A1(n364), .A2(n365), .A3(n[1020]), .Z(n363) );
  XOR4D0 U220 ( .A1(n[1013]), .A2(n[1012]), .A3(n[1015]), .A4(n[1014]), .Z(
        n365) );
  XOR4D0 U221 ( .A1(n[1017]), .A2(n[1016]), .A3(n[1019]), .A4(n[1018]), .Z(
        n364) );
  XOR4D0 U222 ( .A1(n[1024]), .A2(n[1023]), .A3(n[1026]), .A4(n[1025]), .Z(
        n361) );
  XOR4D0 U223 ( .A1(n[1031]), .A2(n[1030]), .A3(n[1033]), .A4(n[1032]), .Z(
        n359) );
  XOR4D0 U224 ( .A1(n[1038]), .A2(n[1037]), .A3(n[1040]), .A4(n[1039]), .Z(
        n356) );
  XOR4D0 U225 ( .A1(n[1045]), .A2(n[1044]), .A3(n[1047]), .A4(n[1046]), .Z(
        n354) );
  XOR4D0 U226 ( .A1(n[1052]), .A2(n[1051]), .A3(n[1054]), .A4(n[1053]), .Z(
        n351) );
  XOR4D0 U227 ( .A1(n[1059]), .A2(n[1058]), .A3(n[1061]), .A4(n[1060]), .Z(
        n349) );
  XOR4D0 U228 ( .A1(n[1066]), .A2(n[1065]), .A3(n[1068]), .A4(n[1067]), .Z(
        n346) );
  XOR4D0 U229 ( .A1(n[1073]), .A2(n[1072]), .A3(n[1075]), .A4(n[1074]), .Z(
        n344) );
  XOR4D0 U230 ( .A1(n[1080]), .A2(n[1079]), .A3(n[1082]), .A4(n[1081]), .Z(
        n341) );
  XOR4D0 U231 ( .A1(n[1087]), .A2(n[1086]), .A3(n[1089]), .A4(n[1088]), .Z(
        n339) );
  XOR4D0 U232 ( .A1(n[1094]), .A2(n[1093]), .A3(n[1096]), .A4(n[1095]), .Z(
        n336) );
  XOR4D0 U233 ( .A1(n[1101]), .A2(n[1100]), .A3(n[1103]), .A4(n[1102]), .Z(
        n334) );
  XOR4D0 U234 ( .A1(n[1108]), .A2(n[1107]), .A3(n[1110]), .A4(n[1109]), .Z(
        n331) );
  XOR4D0 U235 ( .A1(n[1115]), .A2(n[1114]), .A3(n[1117]), .A4(n[1116]), .Z(
        n329) );
  XOR4D0 U236 ( .A1(n[1122]), .A2(n[1121]), .A3(n[1124]), .A4(n[1123]), .Z(
        n326) );
  XOR4D0 U237 ( .A1(n[1129]), .A2(n[1128]), .A3(n[1131]), .A4(n[1130]), .Z(
        n324) );
  XOR4D0 U238 ( .A1(n[1136]), .A2(n[1135]), .A3(n[1138]), .A4(n[1137]), .Z(
        n321) );
  XOR4D0 U239 ( .A1(n[1143]), .A2(n[1142]), .A3(n[1145]), .A4(n[1144]), .Z(
        n319) );
  XOR4D0 U240 ( .A1(n[1150]), .A2(n[1149]), .A3(n[1152]), .A4(n[1151]), .Z(
        n316) );
  XOR4D0 U241 ( .A1(n[1157]), .A2(n[1156]), .A3(n[1159]), .A4(n[1158]), .Z(
        n314) );
  XOR4D0 U242 ( .A1(n[1164]), .A2(n[1163]), .A3(n[1166]), .A4(n[1165]), .Z(
        n311) );
  XOR4D0 U243 ( .A1(n[1171]), .A2(n[1170]), .A3(n[1173]), .A4(n[1172]), .Z(
        n309) );
  XOR4D0 U244 ( .A1(n[1178]), .A2(n[1177]), .A3(n[1180]), .A4(n[1179]), .Z(
        n306) );
  XOR4D0 U245 ( .A1(n[1185]), .A2(n[1184]), .A3(n[1187]), .A4(n[1186]), .Z(
        n304) );
  XOR4D0 U246 ( .A1(n[1192]), .A2(n[1191]), .A3(n[1194]), .A4(n[1193]), .Z(
        n301) );
  XOR4D0 U247 ( .A1(n[1199]), .A2(n[1198]), .A3(n[1201]), .A4(n[1200]), .Z(
        n299) );
  XOR4D0 U248 ( .A1(n[1206]), .A2(n[1205]), .A3(n[1208]), .A4(n[1207]), .Z(
        n296) );
  XOR4D0 U249 ( .A1(n[1213]), .A2(n[1212]), .A3(n[1215]), .A4(n[1214]), .Z(
        n294) );
  XOR4D0 U250 ( .A1(n[1220]), .A2(n[1219]), .A3(n[1222]), .A4(n[1221]), .Z(
        n291) );
  XOR4D0 U251 ( .A1(n[1227]), .A2(n[1226]), .A3(n[1229]), .A4(n[1228]), .Z(
        n289) );
  XOR4D0 U252 ( .A1(n[1234]), .A2(n[1233]), .A3(n[1236]), .A4(n[1235]), .Z(
        n286) );
  XOR4D0 U253 ( .A1(n[1241]), .A2(n[1240]), .A3(n[1243]), .A4(n[1242]), .Z(
        n284) );
  XOR4D0 U254 ( .A1(n[1248]), .A2(n[1247]), .A3(n[1250]), .A4(n[1249]), .Z(
        n281) );
  XOR4D0 U255 ( .A1(n[1255]), .A2(n[1254]), .A3(n[1257]), .A4(n[1256]), .Z(
        n279) );
  XOR4D0 U256 ( .A1(n[1262]), .A2(n[1261]), .A3(n[1264]), .A4(n[1263]), .Z(
        n276) );
  XOR4D0 U257 ( .A1(n[1269]), .A2(n[1268]), .A3(n[1271]), .A4(n[1270]), .Z(
        n274) );
  XOR4D0 U258 ( .A1(n[1276]), .A2(n[1275]), .A3(n[1278]), .A4(n[1277]), .Z(
        n271) );
  XOR4D0 U259 ( .A1(n[1283]), .A2(n[1282]), .A3(n[1285]), .A4(n[1284]), .Z(
        n269) );
  XOR4D0 U260 ( .A1(n[1290]), .A2(n[1289]), .A3(n[1292]), .A4(n[1291]), .Z(
        n266) );
  XOR4D0 U261 ( .A1(n[1297]), .A2(n[1296]), .A3(n[1299]), .A4(n[1298]), .Z(
        n264) );
  XOR4D0 U262 ( .A1(n[1304]), .A2(n[1303]), .A3(n[1306]), .A4(n[1305]), .Z(
        n261) );
  XOR4D0 U263 ( .A1(n[1311]), .A2(n[1310]), .A3(n[1313]), .A4(n[1312]), .Z(
        n259) );
  XOR4D0 U264 ( .A1(n[1318]), .A2(n[1317]), .A3(n[1320]), .A4(n[1319]), .Z(
        n256) );
  XOR4D0 U265 ( .A1(n[1325]), .A2(n[1324]), .A3(n[1327]), .A4(n[1326]), .Z(
        n254) );
  XOR4D0 U266 ( .A1(n[1332]), .A2(n[1331]), .A3(n[1334]), .A4(n[1333]), .Z(
        n251) );
  XOR4D0 U267 ( .A1(n[1339]), .A2(n[1338]), .A3(n[1341]), .A4(n[1340]), .Z(
        n249) );
  XOR4D0 U268 ( .A1(n[1346]), .A2(n[1345]), .A3(n[1348]), .A4(n[1347]), .Z(
        n246) );
  XOR4D0 U269 ( .A1(n[1353]), .A2(n[1352]), .A3(n[1355]), .A4(n[1354]), .Z(
        n244) );
  XOR4D0 U270 ( .A1(n[1360]), .A2(n[1359]), .A3(n[1362]), .A4(n[1361]), .Z(
        n241) );
  XOR4D0 U271 ( .A1(n[1367]), .A2(n[1366]), .A3(n[1369]), .A4(n[1368]), .Z(
        n239) );
  XOR4D0 U272 ( .A1(n[1374]), .A2(n[1373]), .A3(n[1376]), .A4(n[1375]), .Z(
        n236) );
  XOR4D0 U273 ( .A1(n[1381]), .A2(n[1380]), .A3(n[1383]), .A4(n[1382]), .Z(
        n234) );
  XOR4D0 U274 ( .A1(n[1388]), .A2(n[1387]), .A3(n[1390]), .A4(n[1389]), .Z(
        n231) );
  XOR4D0 U275 ( .A1(n[1395]), .A2(n[1394]), .A3(n[1397]), .A4(n[1396]), .Z(
        n229) );
  XOR4D0 U276 ( .A1(n[1402]), .A2(n[1401]), .A3(n[1404]), .A4(n[1403]), .Z(
        n226) );
  XOR4D0 U277 ( .A1(n[1409]), .A2(n[1408]), .A3(n[1411]), .A4(n[1410]), .Z(
        n224) );
  XOR4D0 U278 ( .A1(n[1416]), .A2(n[1415]), .A3(n[1418]), .A4(n[1417]), .Z(
        n221) );
  XOR4D0 U279 ( .A1(n[1423]), .A2(n[1422]), .A3(n[1425]), .A4(n[1424]), .Z(
        n219) );
  XOR4D0 U280 ( .A1(n[1430]), .A2(n[1429]), .A3(n[1432]), .A4(n[1431]), .Z(
        n216) );
  XOR4D0 U281 ( .A1(n[1437]), .A2(n[1436]), .A3(n[1439]), .A4(n[1438]), .Z(
        n214) );
  XOR4D0 U282 ( .A1(n[1444]), .A2(n[1443]), .A3(n[1446]), .A4(n[1445]), .Z(
        n211) );
  XOR4D0 U283 ( .A1(n[1451]), .A2(n[1450]), .A3(n[1453]), .A4(n[1452]), .Z(
        n209) );
  XOR4D0 U284 ( .A1(n[1458]), .A2(n[1457]), .A3(n[1460]), .A4(n[1459]), .Z(
        n206) );
  XOR4D0 U285 ( .A1(n[1465]), .A2(n[1464]), .A3(n[1467]), .A4(n[1466]), .Z(
        n204) );
  XOR4D0 U286 ( .A1(n[1472]), .A2(n[1471]), .A3(n[1474]), .A4(n[1473]), .Z(
        n201) );
  XOR4D0 U287 ( .A1(n[1479]), .A2(n[1478]), .A3(n[1481]), .A4(n[1480]), .Z(
        n199) );
  XOR4D0 U288 ( .A1(n[1486]), .A2(n[1485]), .A3(n[1488]), .A4(n[1487]), .Z(
        n196) );
  XOR4D0 U289 ( .A1(n[1493]), .A2(n[1492]), .A3(n[1495]), .A4(n[1494]), .Z(
        n194) );
  XOR4D0 U290 ( .A1(n[1500]), .A2(n[1499]), .A3(n[1502]), .A4(n[1501]), .Z(
        n191) );
  XOR4D0 U291 ( .A1(n[1507]), .A2(n[1506]), .A3(n[1509]), .A4(n[1508]), .Z(
        n189) );
  XOR4D0 U292 ( .A1(n[1514]), .A2(n[1513]), .A3(n[1516]), .A4(n[1515]), .Z(
        n186) );
  XOR4D0 U293 ( .A1(n[1521]), .A2(n[1520]), .A3(n[1523]), .A4(n[1522]), .Z(
        n184) );
  XOR4D0 U294 ( .A1(n[1528]), .A2(n[1527]), .A3(n[1530]), .A4(n[1529]), .Z(
        n181) );
  XOR4D0 U295 ( .A1(n[1535]), .A2(n[1534]), .A3(n[1537]), .A4(n[1536]), .Z(
        n179) );
  XOR4D0 U296 ( .A1(n[1542]), .A2(n[1541]), .A3(n[1544]), .A4(n[1543]), .Z(
        n176) );
  XOR4D0 U297 ( .A1(n[1549]), .A2(n[1548]), .A3(n[1551]), .A4(n[1550]), .Z(
        n174) );
  XOR4D0 U298 ( .A1(n[1556]), .A2(n[1555]), .A3(n[1558]), .A4(n[1557]), .Z(
        n171) );
  XOR4D0 U299 ( .A1(n[1563]), .A2(n[1562]), .A3(n[1565]), .A4(n[1564]), .Z(
        n169) );
  XOR4D0 U300 ( .A1(n[1570]), .A2(n[1569]), .A3(n[1572]), .A4(n[1571]), .Z(
        n166) );
  XOR4D0 U301 ( .A1(n[1577]), .A2(n[1576]), .A3(n[1579]), .A4(n[1578]), .Z(
        n164) );
  XOR4D0 U302 ( .A1(n[1584]), .A2(n[1583]), .A3(n[1586]), .A4(n[1585]), .Z(
        n161) );
  XOR4D0 U303 ( .A1(n[1591]), .A2(n[1590]), .A3(n[1593]), .A4(n[1592]), .Z(
        n159) );
  XOR4D0 U304 ( .A1(n[1598]), .A2(n[1597]), .A3(n[1600]), .A4(n[1599]), .Z(
        n156) );
  XOR4D0 U305 ( .A1(n[1605]), .A2(n[1604]), .A3(n[1607]), .A4(n[1606]), .Z(
        n154) );
  XOR4D0 U306 ( .A1(n[1612]), .A2(n[1611]), .A3(n[1614]), .A4(n[1613]), .Z(
        n151) );
  XOR4D0 U307 ( .A1(n[1619]), .A2(n[1618]), .A3(n[1621]), .A4(n[1620]), .Z(
        n149) );
  XOR4D0 U308 ( .A1(n[1626]), .A2(n[1625]), .A3(n[1628]), .A4(n[1627]), .Z(
        n146) );
  XOR4D0 U309 ( .A1(n[1633]), .A2(n[1632]), .A3(n[1635]), .A4(n[1634]), .Z(
        n144) );
  XOR4D0 U310 ( .A1(n[1640]), .A2(n[1639]), .A3(n[1642]), .A4(n[1641]), .Z(
        n141) );
  XOR4D0 U311 ( .A1(n[1647]), .A2(n[1646]), .A3(n[1649]), .A4(n[1648]), .Z(
        n139) );
  XOR4D0 U312 ( .A1(n[1654]), .A2(n[1653]), .A3(n[1656]), .A4(n[1655]), .Z(
        n136) );
  XOR4D0 U313 ( .A1(n[1661]), .A2(n[1660]), .A3(n[1663]), .A4(n[1662]), .Z(
        n134) );
  XOR4D0 U314 ( .A1(n[1668]), .A2(n[1667]), .A3(n[1670]), .A4(n[1669]), .Z(
        n131) );
  XOR4D0 U315 ( .A1(n[1675]), .A2(n[1674]), .A3(n[1677]), .A4(n[1676]), .Z(
        n129) );
  XOR4D0 U316 ( .A1(n[1682]), .A2(n[1681]), .A3(n[1684]), .A4(n[1683]), .Z(
        n126) );
  XOR4D0 U317 ( .A1(n[1689]), .A2(n[1688]), .A3(n[1691]), .A4(n[1690]), .Z(
        n124) );
  XOR4D0 U318 ( .A1(n[1696]), .A2(n[1695]), .A3(n[1698]), .A4(n[1697]), .Z(
        n121) );
  XOR4D0 U319 ( .A1(n[1703]), .A2(n[1702]), .A3(n[1705]), .A4(n[1704]), .Z(
        n119) );
  XOR4D0 U320 ( .A1(n[1710]), .A2(n[1709]), .A3(n[1712]), .A4(n[1711]), .Z(
        n116) );
  XOR4D0 U321 ( .A1(n[1717]), .A2(n[1716]), .A3(n[1719]), .A4(n[1718]), .Z(
        n114) );
  XOR4D0 U322 ( .A1(n[1724]), .A2(n[1723]), .A3(n[1726]), .A4(n[1725]), .Z(
        n111) );
  XOR4D0 U323 ( .A1(n[1731]), .A2(n[1730]), .A3(n[1733]), .A4(n[1732]), .Z(
        n109) );
  XOR4D0 U324 ( .A1(n[1738]), .A2(n[1737]), .A3(n[1740]), .A4(n[1739]), .Z(
        n106) );
  XOR4D0 U325 ( .A1(n[1745]), .A2(n[1744]), .A3(n[1747]), .A4(n[1746]), .Z(
        n104) );
  XOR4D0 U326 ( .A1(n[1752]), .A2(n[1751]), .A3(n[1754]), .A4(n[1753]), .Z(
        n101) );
  XOR4D0 U327 ( .A1(n[1759]), .A2(n[1758]), .A3(n[1761]), .A4(n[1760]), .Z(n99) );
  XOR4D0 U328 ( .A1(n[1766]), .A2(n[1765]), .A3(n[1768]), .A4(n[1767]), .Z(n96) );
  XOR4D0 U329 ( .A1(n[1773]), .A2(n[1772]), .A3(n[1775]), .A4(n[1774]), .Z(n94) );
  XOR4D0 U330 ( .A1(n[1780]), .A2(n[1779]), .A3(n[1782]), .A4(n[1781]), .Z(n91) );
  XOR4D0 U331 ( .A1(n[1787]), .A2(n[1786]), .A3(n[1789]), .A4(n[1788]), .Z(n89) );
  XOR4D0 U332 ( .A1(n[1794]), .A2(n[1793]), .A3(n[1796]), .A4(n[1795]), .Z(n86) );
  XOR4D0 U333 ( .A1(n[1801]), .A2(n[1800]), .A3(n[1803]), .A4(n[1802]), .Z(n84) );
  XOR4D0 U334 ( .A1(n[1808]), .A2(n[1807]), .A3(n[1810]), .A4(n[1809]), .Z(n81) );
  XOR4D0 U335 ( .A1(n[1815]), .A2(n[1814]), .A3(n[1817]), .A4(n[1816]), .Z(n79) );
  XOR4D0 U336 ( .A1(n[1822]), .A2(n[1821]), .A3(n[1824]), .A4(n[1823]), .Z(n76) );
  XOR4D0 U337 ( .A1(n[1829]), .A2(n[1828]), .A3(n[1831]), .A4(n[1830]), .Z(n74) );
  XOR4D0 U338 ( .A1(n[1836]), .A2(n[1835]), .A3(n[1838]), .A4(n[1837]), .Z(n71) );
  XOR4D0 U339 ( .A1(n[1843]), .A2(n[1842]), .A3(n[1845]), .A4(n[1844]), .Z(n69) );
  XOR4D0 U340 ( .A1(n[1850]), .A2(n[1849]), .A3(n[1852]), .A4(n[1851]), .Z(n66) );
  XOR4D0 U341 ( .A1(n[1857]), .A2(n[1856]), .A3(n[1859]), .A4(n[1858]), .Z(n64) );
  XOR4D0 U342 ( .A1(n[1864]), .A2(n[1863]), .A3(n[1866]), .A4(n[1865]), .Z(n61) );
  XOR4D0 U343 ( .A1(n[1871]), .A2(n[1870]), .A3(n[1873]), .A4(n[1872]), .Z(n59) );
  XOR4D0 U344 ( .A1(n[1878]), .A2(n[1877]), .A3(n[1880]), .A4(n[1879]), .Z(n56) );
  XOR4D0 U345 ( .A1(n[1885]), .A2(n[1884]), .A3(n[1887]), .A4(n[1886]), .Z(n54) );
  XOR4D0 U346 ( .A1(n[1892]), .A2(n[1891]), .A3(n[1894]), .A4(n[1893]), .Z(n51) );
  XOR4D0 U347 ( .A1(n[1899]), .A2(n[1898]), .A3(n[1901]), .A4(n[1900]), .Z(n49) );
  XOR4D0 U348 ( .A1(n[1906]), .A2(n[1905]), .A3(n[1908]), .A4(n[1907]), .Z(n46) );
  XOR4D0 U349 ( .A1(n[1913]), .A2(n[1912]), .A3(n[1915]), .A4(n[1914]), .Z(n44) );
  XOR4D0 U350 ( .A1(n[1920]), .A2(n[1919]), .A3(n[1922]), .A4(n[1921]), .Z(n41) );
  XOR4D0 U351 ( .A1(n[1927]), .A2(n[1926]), .A3(n[1929]), .A4(n[1928]), .Z(n39) );
  XOR4D0 U352 ( .A1(n[1934]), .A2(n[1933]), .A3(n[1936]), .A4(n[1935]), .Z(n36) );
  XOR4D0 U353 ( .A1(n[1941]), .A2(n[1940]), .A3(n[1943]), .A4(n[1942]), .Z(n34) );
  XOR4D0 U354 ( .A1(n[1948]), .A2(n[1947]), .A3(n[1950]), .A4(n[1949]), .Z(n31) );
  XOR4D0 U355 ( .A1(n[1955]), .A2(n[1954]), .A3(n[1957]), .A4(n[1956]), .Z(n29) );
  XOR4D0 U356 ( .A1(n[1962]), .A2(n[1961]), .A3(n[1964]), .A4(n[1963]), .Z(n26) );
  XOR4D0 U357 ( .A1(n[1969]), .A2(n[1968]), .A3(n[1971]), .A4(n[1970]), .Z(n24) );
  XOR4D0 U358 ( .A1(n[1976]), .A2(n[1975]), .A3(n[1978]), .A4(n[1977]), .Z(n21) );
  XOR4D0 U359 ( .A1(n[1983]), .A2(n[1982]), .A3(n[1985]), .A4(n[1984]), .Z(n19) );
  XOR4D0 U360 ( .A1(n[1990]), .A2(n[1989]), .A3(n[1992]), .A4(n[1991]), .Z(n16) );
  XOR4D0 U361 ( .A1(n[1997]), .A2(n[1996]), .A3(n[1999]), .A4(n[1998]), .Z(n14) );
  XOR4D0 U362 ( .A1(n[2004]), .A2(n[2003]), .A3(n[2006]), .A4(n[2005]), .Z(n11) );
  XOR4D0 U363 ( .A1(n[2011]), .A2(n[2010]), .A3(n[2013]), .A4(n[2012]), .Z(n9)
         );
  XOR4D0 U364 ( .A1(n[2018]), .A2(n[2017]), .A3(n[2020]), .A4(n[2019]), .Z(n6)
         );
  XOR4D0 U365 ( .A1(n[2025]), .A2(n[2024]), .A3(n[2027]), .A4(n[2026]), .Z(n4)
         );
  XOR4D0 U366 ( .A1(n[2032]), .A2(n[2031]), .A3(n[2034]), .A4(n[2033]), .Z(n1)
         );
  XOR3D0 U367 ( .A1(n366), .A2(n367), .A3(n[1011]), .Z(s[8]) );
  XOR4D0 U368 ( .A1(a[8]), .A2(n368), .A3(n[1006]), .A4(b[8]), .Z(n367) );
  XOR4D0 U369 ( .A1(n[1002]), .A2(n[1001]), .A3(n369), .A4(n370), .Z(n368) );
  XOR3D0 U370 ( .A1(n371), .A2(n372), .A3(n[1000]), .Z(n370) );
  XOR4D0 U371 ( .A1(n[992]), .A2(n373), .A3(n[994]), .A4(n[993]), .Z(n372) );
  XOR4D0 U372 ( .A1(n[987]), .A2(n[986]), .A3(n374), .A4(n375), .Z(n373) );
  XOR3D0 U373 ( .A1(n376), .A2(n377), .A3(n[985]), .Z(n375) );
  XOR4D0 U374 ( .A1(n[978]), .A2(n378), .A3(n[980]), .A4(n[979]), .Z(n377) );
  XOR4D0 U375 ( .A1(n[973]), .A2(n[972]), .A3(n379), .A4(n380), .Z(n378) );
  XOR3D0 U376 ( .A1(n381), .A2(n382), .A3(n[971]), .Z(n380) );
  XOR4D0 U377 ( .A1(n[964]), .A2(n383), .A3(n[966]), .A4(n[965]), .Z(n382) );
  XOR4D0 U378 ( .A1(n[959]), .A2(n[958]), .A3(n384), .A4(n385), .Z(n383) );
  XOR3D0 U379 ( .A1(n386), .A2(n387), .A3(n[957]), .Z(n385) );
  XOR4D0 U380 ( .A1(n[950]), .A2(n388), .A3(n[952]), .A4(n[951]), .Z(n387) );
  XOR4D0 U381 ( .A1(n[945]), .A2(n[944]), .A3(n389), .A4(n390), .Z(n388) );
  XOR3D0 U382 ( .A1(n391), .A2(n392), .A3(n[943]), .Z(n390) );
  XOR4D0 U383 ( .A1(n[936]), .A2(n393), .A3(n[938]), .A4(n[937]), .Z(n392) );
  XOR4D0 U384 ( .A1(n[931]), .A2(n[930]), .A3(n394), .A4(n395), .Z(n393) );
  XOR3D0 U385 ( .A1(n396), .A2(n397), .A3(n[929]), .Z(n395) );
  XOR4D0 U386 ( .A1(n[922]), .A2(n398), .A3(n[924]), .A4(n[923]), .Z(n397) );
  XOR4D0 U387 ( .A1(n[917]), .A2(n[916]), .A3(n399), .A4(n400), .Z(n398) );
  XOR3D0 U388 ( .A1(n401), .A2(n402), .A3(n[915]), .Z(n400) );
  XOR4D0 U389 ( .A1(n[908]), .A2(n403), .A3(n[910]), .A4(n[909]), .Z(n402) );
  XOR4D0 U390 ( .A1(n[903]), .A2(n[902]), .A3(n404), .A4(n405), .Z(n403) );
  XOR3D0 U391 ( .A1(n406), .A2(n407), .A3(n[901]), .Z(n405) );
  XOR4D0 U392 ( .A1(n[894]), .A2(n408), .A3(n[896]), .A4(n[895]), .Z(n407) );
  XOR4D0 U393 ( .A1(n[889]), .A2(n[888]), .A3(n409), .A4(n410), .Z(n408) );
  XOR3D0 U394 ( .A1(n411), .A2(n412), .A3(n[887]), .Z(n410) );
  XOR4D0 U395 ( .A1(n[880]), .A2(n413), .A3(n[882]), .A4(n[881]), .Z(n412) );
  XOR4D0 U396 ( .A1(n[875]), .A2(n[874]), .A3(n414), .A4(n415), .Z(n413) );
  XOR3D0 U397 ( .A1(n416), .A2(n417), .A3(n[873]), .Z(n415) );
  XOR4D0 U398 ( .A1(n[866]), .A2(n418), .A3(n[868]), .A4(n[867]), .Z(n417) );
  XOR4D0 U399 ( .A1(n[861]), .A2(n[860]), .A3(n419), .A4(n420), .Z(n418) );
  XOR3D0 U400 ( .A1(n421), .A2(n422), .A3(n[859]), .Z(n420) );
  XOR4D0 U401 ( .A1(n[852]), .A2(n423), .A3(n[854]), .A4(n[853]), .Z(n422) );
  XOR4D0 U402 ( .A1(n[847]), .A2(n[846]), .A3(n424), .A4(n425), .Z(n423) );
  XOR3D0 U403 ( .A1(n426), .A2(n427), .A3(n[845]), .Z(n425) );
  XOR4D0 U404 ( .A1(n[838]), .A2(n428), .A3(n[840]), .A4(n[839]), .Z(n427) );
  XOR4D0 U405 ( .A1(n[833]), .A2(n[832]), .A3(n429), .A4(n430), .Z(n428) );
  XOR3D0 U406 ( .A1(n431), .A2(n432), .A3(n[831]), .Z(n430) );
  XOR4D0 U407 ( .A1(n[824]), .A2(n433), .A3(n[826]), .A4(n[825]), .Z(n432) );
  XOR4D0 U408 ( .A1(n[819]), .A2(n[818]), .A3(n434), .A4(n435), .Z(n433) );
  XOR3D0 U409 ( .A1(n436), .A2(n437), .A3(n[817]), .Z(n435) );
  XOR4D0 U410 ( .A1(n[810]), .A2(n438), .A3(n[812]), .A4(n[811]), .Z(n437) );
  XOR4D0 U411 ( .A1(n[805]), .A2(n[804]), .A3(n439), .A4(n440), .Z(n438) );
  XOR3D0 U412 ( .A1(n441), .A2(n442), .A3(n[803]), .Z(n440) );
  XOR4D0 U413 ( .A1(n[796]), .A2(n443), .A3(n[798]), .A4(n[797]), .Z(n442) );
  XOR4D0 U414 ( .A1(n[791]), .A2(n[790]), .A3(n444), .A4(n445), .Z(n443) );
  XOR3D0 U415 ( .A1(n446), .A2(n447), .A3(n[789]), .Z(n445) );
  XOR4D0 U416 ( .A1(n[782]), .A2(n448), .A3(n[784]), .A4(n[783]), .Z(n447) );
  XOR4D0 U417 ( .A1(n[777]), .A2(n[776]), .A3(n449), .A4(n450), .Z(n448) );
  XOR3D0 U418 ( .A1(n451), .A2(n452), .A3(n[775]), .Z(n450) );
  XOR4D0 U419 ( .A1(n[768]), .A2(n453), .A3(n[770]), .A4(n[769]), .Z(n452) );
  XOR4D0 U420 ( .A1(n[763]), .A2(n[762]), .A3(n454), .A4(n455), .Z(n453) );
  XOR3D0 U421 ( .A1(n456), .A2(n457), .A3(n[761]), .Z(n455) );
  XOR4D0 U422 ( .A1(n[754]), .A2(n458), .A3(n[756]), .A4(n[755]), .Z(n457) );
  XOR4D0 U423 ( .A1(n[749]), .A2(n[748]), .A3(n459), .A4(n460), .Z(n458) );
  XOR3D0 U424 ( .A1(n461), .A2(n462), .A3(n[747]), .Z(n460) );
  XOR4D0 U425 ( .A1(n[740]), .A2(n463), .A3(n[742]), .A4(n[741]), .Z(n462) );
  XOR4D0 U426 ( .A1(n[735]), .A2(n[734]), .A3(n464), .A4(n465), .Z(n463) );
  XOR3D0 U427 ( .A1(n466), .A2(n467), .A3(n[733]), .Z(n465) );
  XOR4D0 U428 ( .A1(n[726]), .A2(n468), .A3(n[728]), .A4(n[727]), .Z(n467) );
  XOR4D0 U429 ( .A1(n[721]), .A2(n[720]), .A3(n469), .A4(n470), .Z(n468) );
  XOR3D0 U430 ( .A1(n471), .A2(n472), .A3(n[719]), .Z(n470) );
  XOR4D0 U431 ( .A1(n[712]), .A2(n473), .A3(n[714]), .A4(n[713]), .Z(n472) );
  XOR4D0 U432 ( .A1(n[707]), .A2(n[706]), .A3(n474), .A4(n475), .Z(n473) );
  XOR3D0 U433 ( .A1(n476), .A2(n477), .A3(n[705]), .Z(n475) );
  XOR4D0 U434 ( .A1(n[698]), .A2(n478), .A3(n[700]), .A4(n[699]), .Z(n477) );
  XOR4D0 U435 ( .A1(n[693]), .A2(n[692]), .A3(n479), .A4(n480), .Z(n478) );
  XOR3D0 U436 ( .A1(n481), .A2(n482), .A3(n[691]), .Z(n480) );
  XOR4D0 U437 ( .A1(n[684]), .A2(n483), .A3(n[686]), .A4(n[685]), .Z(n482) );
  XOR4D0 U438 ( .A1(n[679]), .A2(n[678]), .A3(n484), .A4(n485), .Z(n483) );
  XOR3D0 U439 ( .A1(n486), .A2(n487), .A3(n[677]), .Z(n485) );
  XOR4D0 U440 ( .A1(n[670]), .A2(n488), .A3(n[672]), .A4(n[671]), .Z(n487) );
  XOR4D0 U441 ( .A1(n[665]), .A2(n[664]), .A3(n489), .A4(n490), .Z(n488) );
  XOR3D0 U442 ( .A1(n491), .A2(n492), .A3(n[663]), .Z(n490) );
  XOR4D0 U443 ( .A1(n[656]), .A2(n493), .A3(n[658]), .A4(n[657]), .Z(n492) );
  XOR4D0 U444 ( .A1(n[651]), .A2(n[650]), .A3(n494), .A4(n495), .Z(n493) );
  XOR3D0 U445 ( .A1(n496), .A2(n497), .A3(n[649]), .Z(n495) );
  XOR4D0 U446 ( .A1(n[642]), .A2(n498), .A3(n[644]), .A4(n[643]), .Z(n497) );
  XOR4D0 U447 ( .A1(n[637]), .A2(n[636]), .A3(n499), .A4(n500), .Z(n498) );
  XOR3D0 U448 ( .A1(n501), .A2(n502), .A3(n[635]), .Z(n500) );
  XOR4D0 U449 ( .A1(n[628]), .A2(n503), .A3(n[630]), .A4(n[629]), .Z(n502) );
  XOR4D0 U450 ( .A1(n[623]), .A2(n[622]), .A3(n504), .A4(n505), .Z(n503) );
  XOR3D0 U451 ( .A1(n506), .A2(n507), .A3(n[621]), .Z(n505) );
  XOR4D0 U452 ( .A1(n[614]), .A2(n508), .A3(n[616]), .A4(n[615]), .Z(n507) );
  XOR4D0 U453 ( .A1(n[609]), .A2(n[608]), .A3(n509), .A4(n510), .Z(n508) );
  XOR3D0 U454 ( .A1(n511), .A2(n512), .A3(n[607]), .Z(n510) );
  XOR4D0 U455 ( .A1(n[600]), .A2(n513), .A3(n[602]), .A4(n[601]), .Z(n512) );
  XOR4D0 U456 ( .A1(n[595]), .A2(n[594]), .A3(n514), .A4(n515), .Z(n513) );
  XOR3D0 U457 ( .A1(n516), .A2(n517), .A3(n[593]), .Z(n515) );
  XOR4D0 U458 ( .A1(n[586]), .A2(n518), .A3(n[588]), .A4(n[587]), .Z(n517) );
  XOR4D0 U459 ( .A1(n[581]), .A2(n[580]), .A3(n519), .A4(n520), .Z(n518) );
  XOR3D0 U460 ( .A1(n521), .A2(n522), .A3(n[579]), .Z(n520) );
  XOR4D0 U461 ( .A1(n[572]), .A2(n523), .A3(n[574]), .A4(n[573]), .Z(n522) );
  XOR4D0 U462 ( .A1(n[567]), .A2(n[566]), .A3(n524), .A4(n525), .Z(n523) );
  XOR3D0 U463 ( .A1(n526), .A2(n527), .A3(n[565]), .Z(n525) );
  XOR4D0 U464 ( .A1(n[558]), .A2(n528), .A3(n[560]), .A4(n[559]), .Z(n527) );
  XOR4D0 U465 ( .A1(n[553]), .A2(n[552]), .A3(n529), .A4(n530), .Z(n528) );
  XOR3D0 U466 ( .A1(n531), .A2(n532), .A3(n[551]), .Z(n530) );
  XOR4D0 U467 ( .A1(n[544]), .A2(n533), .A3(n[546]), .A4(n[545]), .Z(n532) );
  XOR4D0 U468 ( .A1(n[539]), .A2(n[538]), .A3(n534), .A4(n535), .Z(n533) );
  XOR3D0 U469 ( .A1(n536), .A2(n537), .A3(n[537]), .Z(n535) );
  XOR4D0 U470 ( .A1(n[530]), .A2(n538), .A3(n[532]), .A4(n[531]), .Z(n537) );
  XOR4D0 U471 ( .A1(n[525]), .A2(n[524]), .A3(n539), .A4(n540), .Z(n538) );
  XOR3D0 U472 ( .A1(n541), .A2(n542), .A3(n[523]), .Z(n540) );
  XOR4D0 U473 ( .A1(n[516]), .A2(n543), .A3(n[518]), .A4(n[517]), .Z(n542) );
  XOR4D0 U474 ( .A1(n[511]), .A2(n[510]), .A3(n544), .A4(n545), .Z(n543) );
  XOR3D0 U475 ( .A1(n546), .A2(n547), .A3(n[509]), .Z(n545) );
  XOR4D0 U476 ( .A1(n[502]), .A2(n[501]), .A3(n[504]), .A4(n[503]), .Z(n547)
         );
  XOR4D0 U477 ( .A1(n[506]), .A2(n[505]), .A3(n[508]), .A4(n[507]), .Z(n546)
         );
  XOR4D0 U478 ( .A1(n[513]), .A2(n[512]), .A3(n[515]), .A4(n[514]), .Z(n544)
         );
  XOR4D0 U479 ( .A1(n[520]), .A2(n[519]), .A3(n[522]), .A4(n[521]), .Z(n541)
         );
  XOR4D0 U480 ( .A1(n[527]), .A2(n[526]), .A3(n[529]), .A4(n[528]), .Z(n539)
         );
  XOR4D0 U481 ( .A1(n[534]), .A2(n[533]), .A3(n[536]), .A4(n[535]), .Z(n536)
         );
  XOR4D0 U482 ( .A1(n[541]), .A2(n[540]), .A3(n[543]), .A4(n[542]), .Z(n534)
         );
  XOR4D0 U483 ( .A1(n[548]), .A2(n[547]), .A3(n[550]), .A4(n[549]), .Z(n531)
         );
  XOR4D0 U484 ( .A1(n[555]), .A2(n[554]), .A3(n[557]), .A4(n[556]), .Z(n529)
         );
  XOR4D0 U485 ( .A1(n[562]), .A2(n[561]), .A3(n[564]), .A4(n[563]), .Z(n526)
         );
  XOR4D0 U486 ( .A1(n[569]), .A2(n[568]), .A3(n[571]), .A4(n[570]), .Z(n524)
         );
  XOR4D0 U487 ( .A1(n[576]), .A2(n[575]), .A3(n[578]), .A4(n[577]), .Z(n521)
         );
  XOR4D0 U488 ( .A1(n[583]), .A2(n[582]), .A3(n[585]), .A4(n[584]), .Z(n519)
         );
  XOR4D0 U489 ( .A1(n[590]), .A2(n[589]), .A3(n[592]), .A4(n[591]), .Z(n516)
         );
  XOR4D0 U490 ( .A1(n[597]), .A2(n[596]), .A3(n[599]), .A4(n[598]), .Z(n514)
         );
  XOR4D0 U491 ( .A1(n[604]), .A2(n[603]), .A3(n[606]), .A4(n[605]), .Z(n511)
         );
  XOR4D0 U492 ( .A1(n[611]), .A2(n[610]), .A3(n[613]), .A4(n[612]), .Z(n509)
         );
  XOR4D0 U493 ( .A1(n[618]), .A2(n[617]), .A3(n[620]), .A4(n[619]), .Z(n506)
         );
  XOR4D0 U494 ( .A1(n[625]), .A2(n[624]), .A3(n[627]), .A4(n[626]), .Z(n504)
         );
  XOR4D0 U495 ( .A1(n[632]), .A2(n[631]), .A3(n[634]), .A4(n[633]), .Z(n501)
         );
  XOR4D0 U496 ( .A1(n[639]), .A2(n[638]), .A3(n[641]), .A4(n[640]), .Z(n499)
         );
  XOR4D0 U497 ( .A1(n[646]), .A2(n[645]), .A3(n[648]), .A4(n[647]), .Z(n496)
         );
  XOR4D0 U498 ( .A1(n[653]), .A2(n[652]), .A3(n[655]), .A4(n[654]), .Z(n494)
         );
  XOR4D0 U499 ( .A1(n[660]), .A2(n[659]), .A3(n[662]), .A4(n[661]), .Z(n491)
         );
  XOR4D0 U500 ( .A1(n[667]), .A2(n[666]), .A3(n[669]), .A4(n[668]), .Z(n489)
         );
  XOR4D0 U501 ( .A1(n[674]), .A2(n[673]), .A3(n[676]), .A4(n[675]), .Z(n486)
         );
  XOR4D0 U502 ( .A1(n[681]), .A2(n[680]), .A3(n[683]), .A4(n[682]), .Z(n484)
         );
  XOR4D0 U503 ( .A1(n[688]), .A2(n[687]), .A3(n[690]), .A4(n[689]), .Z(n481)
         );
  XOR4D0 U504 ( .A1(n[695]), .A2(n[694]), .A3(n[697]), .A4(n[696]), .Z(n479)
         );
  XOR4D0 U505 ( .A1(n[702]), .A2(n[701]), .A3(n[704]), .A4(n[703]), .Z(n476)
         );
  XOR4D0 U506 ( .A1(n[709]), .A2(n[708]), .A3(n[711]), .A4(n[710]), .Z(n474)
         );
  XOR4D0 U507 ( .A1(n[716]), .A2(n[715]), .A3(n[718]), .A4(n[717]), .Z(n471)
         );
  XOR4D0 U508 ( .A1(n[723]), .A2(n[722]), .A3(n[725]), .A4(n[724]), .Z(n469)
         );
  XOR4D0 U509 ( .A1(n[730]), .A2(n[729]), .A3(n[732]), .A4(n[731]), .Z(n466)
         );
  XOR4D0 U510 ( .A1(n[737]), .A2(n[736]), .A3(n[739]), .A4(n[738]), .Z(n464)
         );
  XOR4D0 U511 ( .A1(n[744]), .A2(n[743]), .A3(n[746]), .A4(n[745]), .Z(n461)
         );
  XOR4D0 U512 ( .A1(n[751]), .A2(n[750]), .A3(n[753]), .A4(n[752]), .Z(n459)
         );
  XOR4D0 U513 ( .A1(n[758]), .A2(n[757]), .A3(n[760]), .A4(n[759]), .Z(n456)
         );
  XOR4D0 U514 ( .A1(n[765]), .A2(n[764]), .A3(n[767]), .A4(n[766]), .Z(n454)
         );
  XOR4D0 U515 ( .A1(n[772]), .A2(n[771]), .A3(n[774]), .A4(n[773]), .Z(n451)
         );
  XOR4D0 U516 ( .A1(n[779]), .A2(n[778]), .A3(n[781]), .A4(n[780]), .Z(n449)
         );
  XOR4D0 U517 ( .A1(n[786]), .A2(n[785]), .A3(n[788]), .A4(n[787]), .Z(n446)
         );
  XOR4D0 U518 ( .A1(n[793]), .A2(n[792]), .A3(n[795]), .A4(n[794]), .Z(n444)
         );
  XOR4D0 U519 ( .A1(n[800]), .A2(n[799]), .A3(n[802]), .A4(n[801]), .Z(n441)
         );
  XOR4D0 U520 ( .A1(n[807]), .A2(n[806]), .A3(n[809]), .A4(n[808]), .Z(n439)
         );
  XOR4D0 U521 ( .A1(n[814]), .A2(n[813]), .A3(n[816]), .A4(n[815]), .Z(n436)
         );
  XOR4D0 U522 ( .A1(n[821]), .A2(n[820]), .A3(n[823]), .A4(n[822]), .Z(n434)
         );
  XOR4D0 U523 ( .A1(n[828]), .A2(n[827]), .A3(n[830]), .A4(n[829]), .Z(n431)
         );
  XOR4D0 U524 ( .A1(n[835]), .A2(n[834]), .A3(n[837]), .A4(n[836]), .Z(n429)
         );
  XOR4D0 U525 ( .A1(n[842]), .A2(n[841]), .A3(n[844]), .A4(n[843]), .Z(n426)
         );
  XOR4D0 U526 ( .A1(n[849]), .A2(n[848]), .A3(n[851]), .A4(n[850]), .Z(n424)
         );
  XOR4D0 U527 ( .A1(n[856]), .A2(n[855]), .A3(n[858]), .A4(n[857]), .Z(n421)
         );
  XOR4D0 U528 ( .A1(n[863]), .A2(n[862]), .A3(n[865]), .A4(n[864]), .Z(n419)
         );
  XOR4D0 U529 ( .A1(n[870]), .A2(n[869]), .A3(n[872]), .A4(n[871]), .Z(n416)
         );
  XOR4D0 U530 ( .A1(n[877]), .A2(n[876]), .A3(n[879]), .A4(n[878]), .Z(n414)
         );
  XOR4D0 U531 ( .A1(n[884]), .A2(n[883]), .A3(n[886]), .A4(n[885]), .Z(n411)
         );
  XOR4D0 U532 ( .A1(n[891]), .A2(n[890]), .A3(n[893]), .A4(n[892]), .Z(n409)
         );
  XOR4D0 U533 ( .A1(n[898]), .A2(n[897]), .A3(n[900]), .A4(n[899]), .Z(n406)
         );
  XOR4D0 U534 ( .A1(n[905]), .A2(n[904]), .A3(n[907]), .A4(n[906]), .Z(n404)
         );
  XOR4D0 U535 ( .A1(n[912]), .A2(n[911]), .A3(n[914]), .A4(n[913]), .Z(n401)
         );
  XOR4D0 U536 ( .A1(n[919]), .A2(n[918]), .A3(n[921]), .A4(n[920]), .Z(n399)
         );
  XOR4D0 U537 ( .A1(n[926]), .A2(n[925]), .A3(n[928]), .A4(n[927]), .Z(n396)
         );
  XOR4D0 U538 ( .A1(n[933]), .A2(n[932]), .A3(n[935]), .A4(n[934]), .Z(n394)
         );
  XOR4D0 U539 ( .A1(n[940]), .A2(n[939]), .A3(n[942]), .A4(n[941]), .Z(n391)
         );
  XOR4D0 U540 ( .A1(n[947]), .A2(n[946]), .A3(n[949]), .A4(n[948]), .Z(n389)
         );
  XOR4D0 U541 ( .A1(n[954]), .A2(n[953]), .A3(n[956]), .A4(n[955]), .Z(n386)
         );
  XOR4D0 U542 ( .A1(n[961]), .A2(n[960]), .A3(n[963]), .A4(n[962]), .Z(n384)
         );
  XOR4D0 U543 ( .A1(n[968]), .A2(n[967]), .A3(n[970]), .A4(n[969]), .Z(n381)
         );
  XOR4D0 U544 ( .A1(n[975]), .A2(n[974]), .A3(n[977]), .A4(n[976]), .Z(n379)
         );
  XOR4D0 U545 ( .A1(n[982]), .A2(n[981]), .A3(n[984]), .A4(n[983]), .Z(n376)
         );
  XOR4D0 U546 ( .A1(n[989]), .A2(n[988]), .A3(n[991]), .A4(n[990]), .Z(n374)
         );
  XOR4D0 U547 ( .A1(n[996]), .A2(n[995]), .A3(n[998]), .A4(n[997]), .Z(n371)
         );
  XOR4D0 U548 ( .A1(n[1004]), .A2(n[1003]), .A3(n[999]), .A4(n[1005]), .Z(n369) );
  XOR4D0 U549 ( .A1(n[1008]), .A2(n[1007]), .A3(n[1010]), .A4(n[1009]), .Z(
        n366) );
  XOR4D0 U550 ( .A1(n548), .A2(n549), .A3(n550), .A4(n[495]), .Z(s[7]) );
  XOR3D0 U551 ( .A1(n[498]), .A2(n[497]), .A3(n[496]), .Z(n550) );
  XOR4D0 U552 ( .A1(a[7]), .A2(n551), .A3(n[492]), .A4(b[7]), .Z(n549) );
  XOR4D0 U553 ( .A1(n[487]), .A2(n[486]), .A3(n552), .A4(n553), .Z(n551) );
  XOR3D0 U554 ( .A1(n554), .A2(n555), .A3(n[485]), .Z(n553) );
  XOR4D0 U555 ( .A1(n[478]), .A2(n556), .A3(n[480]), .A4(n[479]), .Z(n555) );
  XOR4D0 U556 ( .A1(n[473]), .A2(n[472]), .A3(n557), .A4(n558), .Z(n556) );
  XOR3D0 U557 ( .A1(n559), .A2(n560), .A3(n[471]), .Z(n558) );
  XOR4D0 U558 ( .A1(n[464]), .A2(n561), .A3(n[466]), .A4(n[465]), .Z(n560) );
  XOR4D0 U559 ( .A1(n[459]), .A2(n[458]), .A3(n562), .A4(n563), .Z(n561) );
  XOR3D0 U560 ( .A1(n564), .A2(n565), .A3(n[457]), .Z(n563) );
  XOR4D0 U561 ( .A1(n[450]), .A2(n566), .A3(n[452]), .A4(n[451]), .Z(n565) );
  XOR4D0 U562 ( .A1(n[445]), .A2(n[444]), .A3(n567), .A4(n568), .Z(n566) );
  XOR3D0 U563 ( .A1(n569), .A2(n570), .A3(n[443]), .Z(n568) );
  XOR4D0 U564 ( .A1(n[436]), .A2(n571), .A3(n[438]), .A4(n[437]), .Z(n570) );
  XOR4D0 U565 ( .A1(n[431]), .A2(n[430]), .A3(n572), .A4(n573), .Z(n571) );
  XOR3D0 U566 ( .A1(n574), .A2(n575), .A3(n[429]), .Z(n573) );
  XOR4D0 U567 ( .A1(n[422]), .A2(n576), .A3(n[424]), .A4(n[423]), .Z(n575) );
  XOR4D0 U568 ( .A1(n[417]), .A2(n[416]), .A3(n577), .A4(n578), .Z(n576) );
  XOR3D0 U569 ( .A1(n579), .A2(n580), .A3(n[415]), .Z(n578) );
  XOR4D0 U570 ( .A1(n[408]), .A2(n581), .A3(n[410]), .A4(n[409]), .Z(n580) );
  XOR4D0 U571 ( .A1(n[403]), .A2(n[402]), .A3(n582), .A4(n583), .Z(n581) );
  XOR3D0 U572 ( .A1(n584), .A2(n585), .A3(n[401]), .Z(n583) );
  XOR4D0 U573 ( .A1(n[394]), .A2(n586), .A3(n[396]), .A4(n[395]), .Z(n585) );
  XOR4D0 U574 ( .A1(n[389]), .A2(n[388]), .A3(n587), .A4(n588), .Z(n586) );
  XOR3D0 U575 ( .A1(n589), .A2(n590), .A3(n[387]), .Z(n588) );
  XOR4D0 U576 ( .A1(n[380]), .A2(n591), .A3(n[382]), .A4(n[381]), .Z(n590) );
  XOR4D0 U577 ( .A1(n[375]), .A2(n[374]), .A3(n592), .A4(n593), .Z(n591) );
  XOR3D0 U578 ( .A1(n594), .A2(n595), .A3(n[373]), .Z(n593) );
  XOR4D0 U579 ( .A1(n[366]), .A2(n596), .A3(n[368]), .A4(n[367]), .Z(n595) );
  XOR4D0 U580 ( .A1(n[361]), .A2(n[360]), .A3(n597), .A4(n598), .Z(n596) );
  XOR3D0 U581 ( .A1(n599), .A2(n600), .A3(n[359]), .Z(n598) );
  XOR4D0 U582 ( .A1(n[352]), .A2(n601), .A3(n[354]), .A4(n[353]), .Z(n600) );
  XOR4D0 U583 ( .A1(n[347]), .A2(n[346]), .A3(n602), .A4(n603), .Z(n601) );
  XOR3D0 U584 ( .A1(n604), .A2(n605), .A3(n[345]), .Z(n603) );
  XOR4D0 U585 ( .A1(n[338]), .A2(n606), .A3(n[340]), .A4(n[339]), .Z(n605) );
  XOR4D0 U586 ( .A1(n[333]), .A2(n[332]), .A3(n607), .A4(n608), .Z(n606) );
  XOR3D0 U587 ( .A1(n609), .A2(n610), .A3(n[331]), .Z(n608) );
  XOR4D0 U588 ( .A1(n[324]), .A2(n611), .A3(n[326]), .A4(n[325]), .Z(n610) );
  XOR4D0 U589 ( .A1(n[319]), .A2(n[318]), .A3(n612), .A4(n613), .Z(n611) );
  XOR3D0 U590 ( .A1(n614), .A2(n615), .A3(n[317]), .Z(n613) );
  XOR4D0 U591 ( .A1(n[310]), .A2(n616), .A3(n[312]), .A4(n[311]), .Z(n615) );
  XOR4D0 U592 ( .A1(n[305]), .A2(n[304]), .A3(n617), .A4(n618), .Z(n616) );
  XOR3D0 U593 ( .A1(n619), .A2(n620), .A3(n[303]), .Z(n618) );
  XOR4D0 U594 ( .A1(n[296]), .A2(n621), .A3(n[298]), .A4(n[297]), .Z(n620) );
  XOR4D0 U595 ( .A1(n[291]), .A2(n[290]), .A3(n622), .A4(n623), .Z(n621) );
  XOR3D0 U596 ( .A1(n624), .A2(n625), .A3(n[289]), .Z(n623) );
  XOR4D0 U597 ( .A1(n[282]), .A2(n626), .A3(n[284]), .A4(n[283]), .Z(n625) );
  XOR4D0 U598 ( .A1(n[277]), .A2(n[276]), .A3(n627), .A4(n628), .Z(n626) );
  XOR3D0 U599 ( .A1(n629), .A2(n630), .A3(n[275]), .Z(n628) );
  XOR4D0 U600 ( .A1(n[268]), .A2(n631), .A3(n[270]), .A4(n[269]), .Z(n630) );
  XOR4D0 U601 ( .A1(n[263]), .A2(n[262]), .A3(n632), .A4(n633), .Z(n631) );
  XOR3D0 U602 ( .A1(n634), .A2(n635), .A3(n[261]), .Z(n633) );
  XOR3D0 U603 ( .A1(n[256]), .A2(n[255]), .A3(n636), .Z(n635) );
  XOR3D0 U604 ( .A1(n637), .A2(n638), .A3(n[254]), .Z(n636) );
  XOR4D0 U605 ( .A1(n[247]), .A2(n[246]), .A3(n[249]), .A4(n[248]), .Z(n638)
         );
  XOR4D0 U606 ( .A1(n[251]), .A2(n[250]), .A3(n[253]), .A4(n[252]), .Z(n637)
         );
  XOR4D0 U607 ( .A1(n[258]), .A2(n[257]), .A3(n[260]), .A4(n[259]), .Z(n634)
         );
  XOR4D0 U608 ( .A1(n[265]), .A2(n[264]), .A3(n[267]), .A4(n[266]), .Z(n632)
         );
  XOR4D0 U609 ( .A1(n[272]), .A2(n[271]), .A3(n[274]), .A4(n[273]), .Z(n629)
         );
  XOR4D0 U610 ( .A1(n[279]), .A2(n[278]), .A3(n[281]), .A4(n[280]), .Z(n627)
         );
  XOR4D0 U611 ( .A1(n[286]), .A2(n[285]), .A3(n[288]), .A4(n[287]), .Z(n624)
         );
  XOR4D0 U612 ( .A1(n[293]), .A2(n[292]), .A3(n[295]), .A4(n[294]), .Z(n622)
         );
  XOR4D0 U613 ( .A1(n[300]), .A2(n[299]), .A3(n[302]), .A4(n[301]), .Z(n619)
         );
  XOR4D0 U614 ( .A1(n[307]), .A2(n[306]), .A3(n[309]), .A4(n[308]), .Z(n617)
         );
  XOR4D0 U615 ( .A1(n[314]), .A2(n[313]), .A3(n[316]), .A4(n[315]), .Z(n614)
         );
  XOR4D0 U616 ( .A1(n[321]), .A2(n[320]), .A3(n[323]), .A4(n[322]), .Z(n612)
         );
  XOR4D0 U617 ( .A1(n[328]), .A2(n[327]), .A3(n[330]), .A4(n[329]), .Z(n609)
         );
  XOR4D0 U618 ( .A1(n[335]), .A2(n[334]), .A3(n[337]), .A4(n[336]), .Z(n607)
         );
  XOR4D0 U619 ( .A1(n[342]), .A2(n[341]), .A3(n[344]), .A4(n[343]), .Z(n604)
         );
  XOR4D0 U620 ( .A1(n[349]), .A2(n[348]), .A3(n[351]), .A4(n[350]), .Z(n602)
         );
  XOR4D0 U621 ( .A1(n[356]), .A2(n[355]), .A3(n[358]), .A4(n[357]), .Z(n599)
         );
  XOR4D0 U622 ( .A1(n[363]), .A2(n[362]), .A3(n[365]), .A4(n[364]), .Z(n597)
         );
  XOR4D0 U623 ( .A1(n[370]), .A2(n[369]), .A3(n[372]), .A4(n[371]), .Z(n594)
         );
  XOR4D0 U624 ( .A1(n[377]), .A2(n[376]), .A3(n[379]), .A4(n[378]), .Z(n592)
         );
  XOR4D0 U625 ( .A1(n[384]), .A2(n[383]), .A3(n[386]), .A4(n[385]), .Z(n589)
         );
  XOR4D0 U626 ( .A1(n[391]), .A2(n[390]), .A3(n[393]), .A4(n[392]), .Z(n587)
         );
  XOR4D0 U627 ( .A1(n[398]), .A2(n[397]), .A3(n[400]), .A4(n[399]), .Z(n584)
         );
  XOR4D0 U628 ( .A1(n[405]), .A2(n[404]), .A3(n[407]), .A4(n[406]), .Z(n582)
         );
  XOR4D0 U629 ( .A1(n[412]), .A2(n[411]), .A3(n[414]), .A4(n[413]), .Z(n579)
         );
  XOR4D0 U630 ( .A1(n[419]), .A2(n[418]), .A3(n[421]), .A4(n[420]), .Z(n577)
         );
  XOR4D0 U631 ( .A1(n[426]), .A2(n[425]), .A3(n[428]), .A4(n[427]), .Z(n574)
         );
  XOR4D0 U632 ( .A1(n[433]), .A2(n[432]), .A3(n[435]), .A4(n[434]), .Z(n572)
         );
  XOR4D0 U633 ( .A1(n[440]), .A2(n[439]), .A3(n[442]), .A4(n[441]), .Z(n569)
         );
  XOR4D0 U634 ( .A1(n[447]), .A2(n[446]), .A3(n[449]), .A4(n[448]), .Z(n567)
         );
  XOR4D0 U635 ( .A1(n[454]), .A2(n[453]), .A3(n[456]), .A4(n[455]), .Z(n564)
         );
  XOR4D0 U636 ( .A1(n[461]), .A2(n[460]), .A3(n[463]), .A4(n[462]), .Z(n562)
         );
  XOR4D0 U637 ( .A1(n[468]), .A2(n[467]), .A3(n[470]), .A4(n[469]), .Z(n559)
         );
  XOR4D0 U638 ( .A1(n[475]), .A2(n[474]), .A3(n[477]), .A4(n[476]), .Z(n557)
         );
  XOR4D0 U639 ( .A1(n[482]), .A2(n[481]), .A3(n[484]), .A4(n[483]), .Z(n554)
         );
  XOR4D0 U640 ( .A1(n[489]), .A2(n[488]), .A3(n[491]), .A4(n[490]), .Z(n552)
         );
  XOR4D0 U641 ( .A1(n[494]), .A2(n[493]), .A3(n[500]), .A4(n[499]), .Z(n548)
         );
  XOR4D0 U642 ( .A1(b[6]), .A2(a[6]), .A3(n639), .A4(n640), .Z(s[6]) );
  XOR4D0 U643 ( .A1(n[239]), .A2(n641), .A3(n[241]), .A4(n[240]), .Z(n640) );
  XOR4D0 U644 ( .A1(n[234]), .A2(n[233]), .A3(n642), .A4(n643), .Z(n641) );
  XOR3D0 U645 ( .A1(n644), .A2(n645), .A3(n[232]), .Z(n643) );
  XOR4D0 U646 ( .A1(n[225]), .A2(n646), .A3(n[227]), .A4(n[226]), .Z(n645) );
  XOR4D0 U647 ( .A1(n[220]), .A2(n[219]), .A3(n647), .A4(n648), .Z(n646) );
  XOR3D0 U648 ( .A1(n649), .A2(n650), .A3(n[218]), .Z(n648) );
  XOR4D0 U649 ( .A1(n[211]), .A2(n651), .A3(n[213]), .A4(n[212]), .Z(n650) );
  XOR4D0 U650 ( .A1(n[206]), .A2(n[205]), .A3(n652), .A4(n653), .Z(n651) );
  XOR3D0 U651 ( .A1(n654), .A2(n655), .A3(n[204]), .Z(n653) );
  XOR4D0 U652 ( .A1(n[197]), .A2(n656), .A3(n[199]), .A4(n[198]), .Z(n655) );
  XOR4D0 U653 ( .A1(n[192]), .A2(n[191]), .A3(n657), .A4(n658), .Z(n656) );
  XOR3D0 U654 ( .A1(n659), .A2(n660), .A3(n[190]), .Z(n658) );
  XOR4D0 U655 ( .A1(n[183]), .A2(n661), .A3(n[185]), .A4(n[184]), .Z(n660) );
  XOR4D0 U656 ( .A1(n[178]), .A2(n[177]), .A3(n662), .A4(n663), .Z(n661) );
  XOR3D0 U657 ( .A1(n664), .A2(n665), .A3(n[176]), .Z(n663) );
  XOR4D0 U658 ( .A1(n[169]), .A2(n666), .A3(n[171]), .A4(n[170]), .Z(n665) );
  XOR4D0 U659 ( .A1(n[164]), .A2(n[163]), .A3(n667), .A4(n668), .Z(n666) );
  XOR3D0 U660 ( .A1(n669), .A2(n670), .A3(n[162]), .Z(n668) );
  XOR4D0 U661 ( .A1(n[155]), .A2(n671), .A3(n[157]), .A4(n[156]), .Z(n670) );
  XOR4D0 U662 ( .A1(n[150]), .A2(n[149]), .A3(n672), .A4(n673), .Z(n671) );
  XOR3D0 U663 ( .A1(n674), .A2(n675), .A3(n[148]), .Z(n673) );
  XOR4D0 U664 ( .A1(n[141]), .A2(n676), .A3(n[143]), .A4(n[142]), .Z(n675) );
  XOR4D0 U665 ( .A1(n[136]), .A2(n[135]), .A3(n677), .A4(n678), .Z(n676) );
  XOR3D0 U666 ( .A1(n679), .A2(n680), .A3(n[134]), .Z(n678) );
  XOR3D0 U667 ( .A1(n[129]), .A2(n[128]), .A3(n681), .Z(n680) );
  XOR3D0 U668 ( .A1(n682), .A2(n683), .A3(n[127]), .Z(n681) );
  XOR4D0 U669 ( .A1(n[120]), .A2(n[119]), .A3(n[122]), .A4(n[121]), .Z(n683)
         );
  XOR4D0 U670 ( .A1(n[124]), .A2(n[123]), .A3(n[126]), .A4(n[125]), .Z(n682)
         );
  XOR4D0 U671 ( .A1(n[131]), .A2(n[130]), .A3(n[133]), .A4(n[132]), .Z(n679)
         );
  XOR4D0 U672 ( .A1(n[138]), .A2(n[137]), .A3(n[140]), .A4(n[139]), .Z(n677)
         );
  XOR4D0 U673 ( .A1(n[145]), .A2(n[144]), .A3(n[147]), .A4(n[146]), .Z(n674)
         );
  XOR4D0 U674 ( .A1(n[152]), .A2(n[151]), .A3(n[154]), .A4(n[153]), .Z(n672)
         );
  XOR4D0 U675 ( .A1(n[159]), .A2(n[158]), .A3(n[161]), .A4(n[160]), .Z(n669)
         );
  XOR4D0 U676 ( .A1(n[166]), .A2(n[165]), .A3(n[168]), .A4(n[167]), .Z(n667)
         );
  XOR4D0 U677 ( .A1(n[173]), .A2(n[172]), .A3(n[175]), .A4(n[174]), .Z(n664)
         );
  XOR4D0 U678 ( .A1(n[180]), .A2(n[179]), .A3(n[182]), .A4(n[181]), .Z(n662)
         );
  XOR4D0 U679 ( .A1(n[187]), .A2(n[186]), .A3(n[189]), .A4(n[188]), .Z(n659)
         );
  XOR4D0 U680 ( .A1(n[194]), .A2(n[193]), .A3(n[196]), .A4(n[195]), .Z(n657)
         );
  XOR4D0 U681 ( .A1(n[201]), .A2(n[200]), .A3(n[203]), .A4(n[202]), .Z(n654)
         );
  XOR4D0 U682 ( .A1(n[208]), .A2(n[207]), .A3(n[210]), .A4(n[209]), .Z(n652)
         );
  XOR4D0 U683 ( .A1(n[215]), .A2(n[214]), .A3(n[217]), .A4(n[216]), .Z(n649)
         );
  XOR4D0 U684 ( .A1(n[222]), .A2(n[221]), .A3(n[224]), .A4(n[223]), .Z(n647)
         );
  XOR4D0 U685 ( .A1(n[229]), .A2(n[228]), .A3(n[231]), .A4(n[230]), .Z(n644)
         );
  XOR4D0 U686 ( .A1(n[236]), .A2(n[235]), .A3(n[238]), .A4(n[237]), .Z(n642)
         );
  XOR4D0 U687 ( .A1(n[243]), .A2(n[242]), .A3(n[245]), .A4(n[244]), .Z(n639)
         );
  XOR3D0 U688 ( .A1(n684), .A2(n685), .A3(n[118]), .Z(s[5]) );
  XOR4D0 U689 ( .A1(a[5]), .A2(n686), .A3(n[113]), .A4(b[5]), .Z(n685) );
  XOR4D0 U690 ( .A1(n[108]), .A2(n[107]), .A3(n687), .A4(n688), .Z(n686) );
  XOR3D0 U691 ( .A1(n689), .A2(n690), .A3(n[106]), .Z(n688) );
  XOR4D0 U692 ( .A1(n[100]), .A2(n691), .A3(n[102]), .A4(n[101]), .Z(n690) );
  XOR4D0 U693 ( .A1(n[94]), .A2(n[93]), .A3(n692), .A4(n693), .Z(n691) );
  XOR3D0 U694 ( .A1(n694), .A2(n695), .A3(n[92]), .Z(n693) );
  XOR4D0 U695 ( .A1(n[85]), .A2(n696), .A3(n[87]), .A4(n[86]), .Z(n695) );
  XOR4D0 U696 ( .A1(n[80]), .A2(n[79]), .A3(n697), .A4(n698), .Z(n696) );
  XOR3D0 U697 ( .A1(n699), .A2(n700), .A3(n[78]), .Z(n698) );
  XOR4D0 U698 ( .A1(n[71]), .A2(n701), .A3(n[73]), .A4(n[72]), .Z(n700) );
  XOR4D0 U699 ( .A1(n[66]), .A2(n[65]), .A3(n702), .A4(n703), .Z(n701) );
  XOR3D0 U700 ( .A1(n704), .A2(n705), .A3(n[64]), .Z(n703) );
  XOR4D0 U701 ( .A1(n[57]), .A2(n[56]), .A3(n[59]), .A4(n[58]), .Z(n705) );
  XOR4D0 U702 ( .A1(n[61]), .A2(n[60]), .A3(n[63]), .A4(n[62]), .Z(n704) );
  XOR4D0 U703 ( .A1(n[68]), .A2(n[67]), .A3(n[70]), .A4(n[69]), .Z(n702) );
  XOR4D0 U704 ( .A1(n[75]), .A2(n[74]), .A3(n[77]), .A4(n[76]), .Z(n699) );
  XOR4D0 U705 ( .A1(n[82]), .A2(n[81]), .A3(n[84]), .A4(n[83]), .Z(n697) );
  XOR4D0 U706 ( .A1(n[89]), .A2(n[88]), .A3(n[91]), .A4(n[90]), .Z(n694) );
  XOR4D0 U707 ( .A1(n[96]), .A2(n[95]), .A3(n[98]), .A4(n[97]), .Z(n692) );
  XOR4D0 U708 ( .A1(n[104]), .A2(n[103]), .A3(n[99]), .A4(n[105]), .Z(n689) );
  XOR4D0 U709 ( .A1(n[110]), .A2(n[109]), .A3(n[112]), .A4(n[111]), .Z(n687)
         );
  XOR4D0 U710 ( .A1(n[115]), .A2(n[114]), .A3(n[117]), .A4(n[116]), .Z(n684)
         );
  XOR4D0 U711 ( .A1(n706), .A2(n707), .A3(n708), .A4(n[50]), .Z(s[4]) );
  XOR3D0 U712 ( .A1(n[53]), .A2(n[52]), .A3(n[51]), .Z(n708) );
  XOR4D0 U713 ( .A1(a[4]), .A2(n709), .A3(n[47]), .A4(b[4]), .Z(n707) );
  XOR4D0 U714 ( .A1(n[42]), .A2(n[41]), .A3(n710), .A4(n711), .Z(n709) );
  XOR3D0 U715 ( .A1(n712), .A2(n713), .A3(n[40]), .Z(n711) );
  XOR3D0 U716 ( .A1(n[35]), .A2(n[34]), .A3(n714), .Z(n713) );
  XOR3D0 U717 ( .A1(n715), .A2(n716), .A3(n[33]), .Z(n714) );
  XOR4D0 U718 ( .A1(n[26]), .A2(n[25]), .A3(n[28]), .A4(n[27]), .Z(n716) );
  XOR4D0 U719 ( .A1(n[30]), .A2(n[29]), .A3(n[32]), .A4(n[31]), .Z(n715) );
  XOR4D0 U720 ( .A1(n[37]), .A2(n[36]), .A3(n[39]), .A4(n[38]), .Z(n712) );
  XOR4D0 U721 ( .A1(n[44]), .A2(n[43]), .A3(n[46]), .A4(n[45]), .Z(n710) );
  XOR4D0 U722 ( .A1(n[49]), .A2(n[48]), .A3(n[55]), .A4(n[54]), .Z(n706) );
  XOR4D0 U723 ( .A1(b[3]), .A2(a[3]), .A3(n717), .A4(n718), .Z(s[3]) );
  XOR3D0 U724 ( .A1(n[20]), .A2(n[19]), .A3(n719), .Z(n718) );
  XOR3D0 U725 ( .A1(n720), .A2(n721), .A3(n[18]), .Z(n719) );
  XOR4D0 U726 ( .A1(n[11]), .A2(n[10]), .A3(n[13]), .A4(n[12]), .Z(n721) );
  XOR4D0 U727 ( .A1(n[15]), .A2(n[14]), .A3(n[17]), .A4(n[16]), .Z(n720) );
  XOR4D0 U728 ( .A1(n[22]), .A2(n[21]), .A3(n[24]), .A4(n[23]), .Z(n717) );
  XOR3D0 U729 ( .A1(n722), .A2(n723), .A3(n[9]), .Z(s[2]) );
  XOR4D0 U730 ( .A1(b[2]), .A2(a[2]), .A3(n[4]), .A4(n[3]), .Z(n723) );
  XOR4D0 U731 ( .A1(n[6]), .A2(n[5]), .A3(n[8]), .A4(n[7]), .Z(n722) );
  XOR3D0 U732 ( .A1(b[1]), .A2(a[1]), .A3(n724), .Z(s[1]) );
  XOR3D0 U733 ( .A1(n[2]), .A2(n[1]), .A3(n[0]), .Z(n724) );
  XOR4D0 U734 ( .A1(n725), .A2(n726), .A3(n727), .A4(n[4076]), .Z(s[10]) );
  XOR3D0 U735 ( .A1(n[4079]), .A2(n[4078]), .A3(n[4077]), .Z(n727) );
  XOR4D0 U736 ( .A1(a[10]), .A2(n728), .A3(n[4073]), .A4(b[10]), .Z(n726) );
  XOR4D0 U737 ( .A1(n[4068]), .A2(n[4067]), .A3(n729), .A4(n730), .Z(n728) );
  XOR3D0 U738 ( .A1(n731), .A2(n732), .A3(n[4066]), .Z(n730) );
  XOR4D0 U739 ( .A1(n[4059]), .A2(n733), .A3(n[4061]), .A4(n[4060]), .Z(n732)
         );
  XOR4D0 U740 ( .A1(n[4054]), .A2(n[4053]), .A3(n734), .A4(n735), .Z(n733) );
  XOR3D0 U741 ( .A1(n736), .A2(n737), .A3(n[4052]), .Z(n735) );
  XOR4D0 U742 ( .A1(n[4045]), .A2(n738), .A3(n[4047]), .A4(n[4046]), .Z(n737)
         );
  XOR4D0 U743 ( .A1(n[4040]), .A2(n[4039]), .A3(n739), .A4(n740), .Z(n738) );
  XOR3D0 U744 ( .A1(n741), .A2(n742), .A3(n[4038]), .Z(n740) );
  XOR4D0 U745 ( .A1(n[4031]), .A2(n743), .A3(n[4033]), .A4(n[4032]), .Z(n742)
         );
  XOR4D0 U746 ( .A1(n[4026]), .A2(n[4025]), .A3(n744), .A4(n745), .Z(n743) );
  XOR3D0 U747 ( .A1(n746), .A2(n747), .A3(n[4024]), .Z(n745) );
  XOR4D0 U748 ( .A1(n[4017]), .A2(n748), .A3(n[4019]), .A4(n[4018]), .Z(n747)
         );
  XOR4D0 U749 ( .A1(n[4012]), .A2(n[4011]), .A3(n749), .A4(n750), .Z(n748) );
  XOR3D0 U750 ( .A1(n751), .A2(n752), .A3(n[4010]), .Z(n750) );
  XOR4D0 U751 ( .A1(n[4003]), .A2(n753), .A3(n[4005]), .A4(n[4004]), .Z(n752)
         );
  XOR4D0 U752 ( .A1(n[3998]), .A2(n[3997]), .A3(n754), .A4(n755), .Z(n753) );
  XOR3D0 U753 ( .A1(n756), .A2(n757), .A3(n[3996]), .Z(n755) );
  XOR4D0 U754 ( .A1(n[3989]), .A2(n758), .A3(n[3991]), .A4(n[3990]), .Z(n757)
         );
  XOR4D0 U755 ( .A1(n[3984]), .A2(n[3983]), .A3(n759), .A4(n760), .Z(n758) );
  XOR3D0 U756 ( .A1(n761), .A2(n762), .A3(n[3982]), .Z(n760) );
  XOR4D0 U757 ( .A1(n[3975]), .A2(n763), .A3(n[3977]), .A4(n[3976]), .Z(n762)
         );
  XOR4D0 U758 ( .A1(n[3970]), .A2(n[3969]), .A3(n764), .A4(n765), .Z(n763) );
  XOR3D0 U759 ( .A1(n766), .A2(n767), .A3(n[3968]), .Z(n765) );
  XOR4D0 U760 ( .A1(n[3961]), .A2(n768), .A3(n[3963]), .A4(n[3962]), .Z(n767)
         );
  XOR4D0 U761 ( .A1(n[3956]), .A2(n[3955]), .A3(n769), .A4(n770), .Z(n768) );
  XOR3D0 U762 ( .A1(n771), .A2(n772), .A3(n[3954]), .Z(n770) );
  XOR4D0 U763 ( .A1(n[3947]), .A2(n773), .A3(n[3949]), .A4(n[3948]), .Z(n772)
         );
  XOR4D0 U764 ( .A1(n[3942]), .A2(n[3941]), .A3(n774), .A4(n775), .Z(n773) );
  XOR3D0 U765 ( .A1(n776), .A2(n777), .A3(n[3940]), .Z(n775) );
  XOR4D0 U766 ( .A1(n[3933]), .A2(n778), .A3(n[3935]), .A4(n[3934]), .Z(n777)
         );
  XOR4D0 U767 ( .A1(n[3928]), .A2(n[3927]), .A3(n779), .A4(n780), .Z(n778) );
  XOR3D0 U768 ( .A1(n781), .A2(n782), .A3(n[3926]), .Z(n780) );
  XOR4D0 U769 ( .A1(n[3919]), .A2(n783), .A3(n[3921]), .A4(n[3920]), .Z(n782)
         );
  XOR4D0 U770 ( .A1(n[3914]), .A2(n[3913]), .A3(n784), .A4(n785), .Z(n783) );
  XOR3D0 U771 ( .A1(n786), .A2(n787), .A3(n[3912]), .Z(n785) );
  XOR4D0 U772 ( .A1(n[3905]), .A2(n788), .A3(n[3907]), .A4(n[3906]), .Z(n787)
         );
  XOR4D0 U773 ( .A1(n[3900]), .A2(n[3899]), .A3(n789), .A4(n790), .Z(n788) );
  XOR3D0 U774 ( .A1(n791), .A2(n792), .A3(n[3898]), .Z(n790) );
  XOR4D0 U775 ( .A1(n[3891]), .A2(n793), .A3(n[3893]), .A4(n[3892]), .Z(n792)
         );
  XOR4D0 U776 ( .A1(n[3886]), .A2(n[3885]), .A3(n794), .A4(n795), .Z(n793) );
  XOR3D0 U777 ( .A1(n796), .A2(n797), .A3(n[3884]), .Z(n795) );
  XOR4D0 U778 ( .A1(n[3877]), .A2(n798), .A3(n[3879]), .A4(n[3878]), .Z(n797)
         );
  XOR4D0 U779 ( .A1(n[3872]), .A2(n[3871]), .A3(n799), .A4(n800), .Z(n798) );
  XOR3D0 U780 ( .A1(n801), .A2(n802), .A3(n[3870]), .Z(n800) );
  XOR4D0 U781 ( .A1(n[3863]), .A2(n803), .A3(n[3865]), .A4(n[3864]), .Z(n802)
         );
  XOR4D0 U782 ( .A1(n[3858]), .A2(n[3857]), .A3(n804), .A4(n805), .Z(n803) );
  XOR3D0 U783 ( .A1(n806), .A2(n807), .A3(n[3856]), .Z(n805) );
  XOR4D0 U784 ( .A1(n[3849]), .A2(n808), .A3(n[3851]), .A4(n[3850]), .Z(n807)
         );
  XOR4D0 U785 ( .A1(n[3844]), .A2(n[3843]), .A3(n809), .A4(n810), .Z(n808) );
  XOR3D0 U786 ( .A1(n811), .A2(n812), .A3(n[3842]), .Z(n810) );
  XOR4D0 U787 ( .A1(n[3835]), .A2(n813), .A3(n[3837]), .A4(n[3836]), .Z(n812)
         );
  XOR4D0 U788 ( .A1(n[3830]), .A2(n[3829]), .A3(n814), .A4(n815), .Z(n813) );
  XOR3D0 U789 ( .A1(n816), .A2(n817), .A3(n[3828]), .Z(n815) );
  XOR4D0 U790 ( .A1(n[3821]), .A2(n818), .A3(n[3823]), .A4(n[3822]), .Z(n817)
         );
  XOR4D0 U791 ( .A1(n[3816]), .A2(n[3815]), .A3(n819), .A4(n820), .Z(n818) );
  XOR3D0 U792 ( .A1(n821), .A2(n822), .A3(n[3814]), .Z(n820) );
  XOR4D0 U793 ( .A1(n[3807]), .A2(n823), .A3(n[3809]), .A4(n[3808]), .Z(n822)
         );
  XOR4D0 U794 ( .A1(n[3802]), .A2(n[3801]), .A3(n824), .A4(n825), .Z(n823) );
  XOR3D0 U795 ( .A1(n826), .A2(n827), .A3(n[3800]), .Z(n825) );
  XOR4D0 U796 ( .A1(n[3793]), .A2(n828), .A3(n[3795]), .A4(n[3794]), .Z(n827)
         );
  XOR4D0 U797 ( .A1(n[3788]), .A2(n[3787]), .A3(n829), .A4(n830), .Z(n828) );
  XOR3D0 U798 ( .A1(n831), .A2(n832), .A3(n[3786]), .Z(n830) );
  XOR4D0 U799 ( .A1(n[3779]), .A2(n833), .A3(n[3781]), .A4(n[3780]), .Z(n832)
         );
  XOR4D0 U800 ( .A1(n[3774]), .A2(n[3773]), .A3(n834), .A4(n835), .Z(n833) );
  XOR3D0 U801 ( .A1(n836), .A2(n837), .A3(n[3772]), .Z(n835) );
  XOR4D0 U802 ( .A1(n[3765]), .A2(n838), .A3(n[3767]), .A4(n[3766]), .Z(n837)
         );
  XOR4D0 U803 ( .A1(n[3760]), .A2(n[3759]), .A3(n839), .A4(n840), .Z(n838) );
  XOR3D0 U804 ( .A1(n841), .A2(n842), .A3(n[3758]), .Z(n840) );
  XOR4D0 U805 ( .A1(n[3751]), .A2(n843), .A3(n[3753]), .A4(n[3752]), .Z(n842)
         );
  XOR4D0 U806 ( .A1(n[3746]), .A2(n[3745]), .A3(n844), .A4(n845), .Z(n843) );
  XOR3D0 U807 ( .A1(n846), .A2(n847), .A3(n[3744]), .Z(n845) );
  XOR4D0 U808 ( .A1(n[3737]), .A2(n848), .A3(n[3739]), .A4(n[3738]), .Z(n847)
         );
  XOR4D0 U809 ( .A1(n[3732]), .A2(n[3731]), .A3(n849), .A4(n850), .Z(n848) );
  XOR3D0 U810 ( .A1(n851), .A2(n852), .A3(n[3730]), .Z(n850) );
  XOR4D0 U811 ( .A1(n[3723]), .A2(n853), .A3(n[3725]), .A4(n[3724]), .Z(n852)
         );
  XOR4D0 U812 ( .A1(n[3718]), .A2(n[3717]), .A3(n854), .A4(n855), .Z(n853) );
  XOR3D0 U813 ( .A1(n856), .A2(n857), .A3(n[3716]), .Z(n855) );
  XOR4D0 U814 ( .A1(n[3709]), .A2(n858), .A3(n[3711]), .A4(n[3710]), .Z(n857)
         );
  XOR4D0 U815 ( .A1(n[3704]), .A2(n[3703]), .A3(n859), .A4(n860), .Z(n858) );
  XOR3D0 U816 ( .A1(n861), .A2(n862), .A3(n[3702]), .Z(n860) );
  XOR4D0 U817 ( .A1(n[3695]), .A2(n863), .A3(n[3697]), .A4(n[3696]), .Z(n862)
         );
  XOR4D0 U818 ( .A1(n[3690]), .A2(n[3689]), .A3(n864), .A4(n865), .Z(n863) );
  XOR3D0 U819 ( .A1(n866), .A2(n867), .A3(n[3688]), .Z(n865) );
  XOR4D0 U820 ( .A1(n[3681]), .A2(n868), .A3(n[3683]), .A4(n[3682]), .Z(n867)
         );
  XOR4D0 U821 ( .A1(n[3676]), .A2(n[3675]), .A3(n869), .A4(n870), .Z(n868) );
  XOR3D0 U822 ( .A1(n871), .A2(n872), .A3(n[3674]), .Z(n870) );
  XOR4D0 U823 ( .A1(n[3667]), .A2(n873), .A3(n[3669]), .A4(n[3668]), .Z(n872)
         );
  XOR4D0 U824 ( .A1(n[3662]), .A2(n[3661]), .A3(n874), .A4(n875), .Z(n873) );
  XOR3D0 U825 ( .A1(n876), .A2(n877), .A3(n[3660]), .Z(n875) );
  XOR4D0 U826 ( .A1(n[3653]), .A2(n878), .A3(n[3655]), .A4(n[3654]), .Z(n877)
         );
  XOR4D0 U827 ( .A1(n[3648]), .A2(n[3647]), .A3(n879), .A4(n880), .Z(n878) );
  XOR3D0 U828 ( .A1(n881), .A2(n882), .A3(n[3646]), .Z(n880) );
  XOR4D0 U829 ( .A1(n[3639]), .A2(n883), .A3(n[3641]), .A4(n[3640]), .Z(n882)
         );
  XOR4D0 U830 ( .A1(n[3634]), .A2(n[3633]), .A3(n884), .A4(n885), .Z(n883) );
  XOR3D0 U831 ( .A1(n886), .A2(n887), .A3(n[3632]), .Z(n885) );
  XOR4D0 U832 ( .A1(n[3625]), .A2(n888), .A3(n[3627]), .A4(n[3626]), .Z(n887)
         );
  XOR4D0 U833 ( .A1(n[3620]), .A2(n[3619]), .A3(n889), .A4(n890), .Z(n888) );
  XOR3D0 U834 ( .A1(n891), .A2(n892), .A3(n[3618]), .Z(n890) );
  XOR4D0 U835 ( .A1(n[3611]), .A2(n893), .A3(n[3613]), .A4(n[3612]), .Z(n892)
         );
  XOR4D0 U836 ( .A1(n[3606]), .A2(n[3605]), .A3(n894), .A4(n895), .Z(n893) );
  XOR3D0 U837 ( .A1(n896), .A2(n897), .A3(n[3604]), .Z(n895) );
  XOR4D0 U838 ( .A1(n[3597]), .A2(n898), .A3(n[3599]), .A4(n[3598]), .Z(n897)
         );
  XOR4D0 U839 ( .A1(n[3592]), .A2(n[3591]), .A3(n899), .A4(n900), .Z(n898) );
  XOR3D0 U840 ( .A1(n901), .A2(n902), .A3(n[3590]), .Z(n900) );
  XOR4D0 U841 ( .A1(n[3583]), .A2(n903), .A3(n[3585]), .A4(n[3584]), .Z(n902)
         );
  XOR4D0 U842 ( .A1(n[3578]), .A2(n[3577]), .A3(n904), .A4(n905), .Z(n903) );
  XOR3D0 U843 ( .A1(n906), .A2(n907), .A3(n[3576]), .Z(n905) );
  XOR4D0 U844 ( .A1(n[3569]), .A2(n908), .A3(n[3571]), .A4(n[3570]), .Z(n907)
         );
  XOR4D0 U845 ( .A1(n[3564]), .A2(n[3563]), .A3(n909), .A4(n910), .Z(n908) );
  XOR3D0 U846 ( .A1(n911), .A2(n912), .A3(n[3562]), .Z(n910) );
  XOR4D0 U847 ( .A1(n[3555]), .A2(n913), .A3(n[3557]), .A4(n[3556]), .Z(n912)
         );
  XOR4D0 U848 ( .A1(n[3550]), .A2(n[3549]), .A3(n914), .A4(n915), .Z(n913) );
  XOR3D0 U849 ( .A1(n916), .A2(n917), .A3(n[3548]), .Z(n915) );
  XOR4D0 U850 ( .A1(n[3541]), .A2(n918), .A3(n[3543]), .A4(n[3542]), .Z(n917)
         );
  XOR4D0 U851 ( .A1(n[3536]), .A2(n[3535]), .A3(n919), .A4(n920), .Z(n918) );
  XOR3D0 U852 ( .A1(n921), .A2(n922), .A3(n[3534]), .Z(n920) );
  XOR4D0 U853 ( .A1(n[3527]), .A2(n923), .A3(n[3529]), .A4(n[3528]), .Z(n922)
         );
  XOR4D0 U854 ( .A1(n[3522]), .A2(n[3521]), .A3(n924), .A4(n925), .Z(n923) );
  XOR3D0 U855 ( .A1(n926), .A2(n927), .A3(n[3520]), .Z(n925) );
  XOR4D0 U856 ( .A1(n[3513]), .A2(n928), .A3(n[3515]), .A4(n[3514]), .Z(n927)
         );
  XOR4D0 U857 ( .A1(n[3508]), .A2(n[3507]), .A3(n929), .A4(n930), .Z(n928) );
  XOR3D0 U858 ( .A1(n931), .A2(n932), .A3(n[3506]), .Z(n930) );
  XOR4D0 U859 ( .A1(n[3499]), .A2(n933), .A3(n[3501]), .A4(n[3500]), .Z(n932)
         );
  XOR4D0 U860 ( .A1(n[3494]), .A2(n[3493]), .A3(n934), .A4(n935), .Z(n933) );
  XOR3D0 U861 ( .A1(n936), .A2(n937), .A3(n[3492]), .Z(n935) );
  XOR4D0 U862 ( .A1(n[3485]), .A2(n938), .A3(n[3487]), .A4(n[3486]), .Z(n937)
         );
  XOR4D0 U863 ( .A1(n[3480]), .A2(n[3479]), .A3(n939), .A4(n940), .Z(n938) );
  XOR3D0 U864 ( .A1(n941), .A2(n942), .A3(n[3478]), .Z(n940) );
  XOR4D0 U865 ( .A1(n[3471]), .A2(n943), .A3(n[3473]), .A4(n[3472]), .Z(n942)
         );
  XOR4D0 U866 ( .A1(n[3466]), .A2(n[3465]), .A3(n944), .A4(n945), .Z(n943) );
  XOR3D0 U867 ( .A1(n946), .A2(n947), .A3(n[3464]), .Z(n945) );
  XOR4D0 U868 ( .A1(n[3457]), .A2(n948), .A3(n[3459]), .A4(n[3458]), .Z(n947)
         );
  XOR4D0 U869 ( .A1(n[3452]), .A2(n[3451]), .A3(n949), .A4(n950), .Z(n948) );
  XOR3D0 U870 ( .A1(n951), .A2(n952), .A3(n[3450]), .Z(n950) );
  XOR4D0 U871 ( .A1(n[3443]), .A2(n953), .A3(n[3445]), .A4(n[3444]), .Z(n952)
         );
  XOR4D0 U872 ( .A1(n[3438]), .A2(n[3437]), .A3(n954), .A4(n955), .Z(n953) );
  XOR3D0 U873 ( .A1(n956), .A2(n957), .A3(n[3436]), .Z(n955) );
  XOR4D0 U874 ( .A1(n[3429]), .A2(n958), .A3(n[3431]), .A4(n[3430]), .Z(n957)
         );
  XOR4D0 U875 ( .A1(n[3424]), .A2(n[3423]), .A3(n959), .A4(n960), .Z(n958) );
  XOR3D0 U876 ( .A1(n961), .A2(n962), .A3(n[3422]), .Z(n960) );
  XOR4D0 U877 ( .A1(n[3415]), .A2(n963), .A3(n[3417]), .A4(n[3416]), .Z(n962)
         );
  XOR4D0 U878 ( .A1(n[3410]), .A2(n[3409]), .A3(n964), .A4(n965), .Z(n963) );
  XOR3D0 U879 ( .A1(n966), .A2(n967), .A3(n[3408]), .Z(n965) );
  XOR4D0 U880 ( .A1(n[3401]), .A2(n968), .A3(n[3403]), .A4(n[3402]), .Z(n967)
         );
  XOR4D0 U881 ( .A1(n[3396]), .A2(n[3395]), .A3(n969), .A4(n970), .Z(n968) );
  XOR3D0 U882 ( .A1(n971), .A2(n972), .A3(n[3394]), .Z(n970) );
  XOR4D0 U883 ( .A1(n[3387]), .A2(n973), .A3(n[3389]), .A4(n[3388]), .Z(n972)
         );
  XOR4D0 U884 ( .A1(n[3382]), .A2(n[3381]), .A3(n974), .A4(n975), .Z(n973) );
  XOR3D0 U885 ( .A1(n976), .A2(n977), .A3(n[3380]), .Z(n975) );
  XOR4D0 U886 ( .A1(n[3373]), .A2(n978), .A3(n[3375]), .A4(n[3374]), .Z(n977)
         );
  XOR4D0 U887 ( .A1(n[3368]), .A2(n[3367]), .A3(n979), .A4(n980), .Z(n978) );
  XOR3D0 U888 ( .A1(n981), .A2(n982), .A3(n[3366]), .Z(n980) );
  XOR4D0 U889 ( .A1(n[3359]), .A2(n983), .A3(n[3361]), .A4(n[3360]), .Z(n982)
         );
  XOR4D0 U890 ( .A1(n[3354]), .A2(n[3353]), .A3(n984), .A4(n985), .Z(n983) );
  XOR3D0 U891 ( .A1(n986), .A2(n987), .A3(n[3352]), .Z(n985) );
  XOR4D0 U892 ( .A1(n[3345]), .A2(n988), .A3(n[3347]), .A4(n[3346]), .Z(n987)
         );
  XOR4D0 U893 ( .A1(n[3340]), .A2(n[3339]), .A3(n989), .A4(n990), .Z(n988) );
  XOR3D0 U894 ( .A1(n991), .A2(n992), .A3(n[3338]), .Z(n990) );
  XOR4D0 U895 ( .A1(n[3331]), .A2(n993), .A3(n[3333]), .A4(n[3332]), .Z(n992)
         );
  XOR4D0 U896 ( .A1(n[3326]), .A2(n[3325]), .A3(n994), .A4(n995), .Z(n993) );
  XOR3D0 U897 ( .A1(n996), .A2(n997), .A3(n[3324]), .Z(n995) );
  XOR4D0 U898 ( .A1(n[3317]), .A2(n998), .A3(n[3319]), .A4(n[3318]), .Z(n997)
         );
  XOR4D0 U899 ( .A1(n[3312]), .A2(n[3311]), .A3(n999), .A4(n1000), .Z(n998) );
  XOR3D0 U900 ( .A1(n1001), .A2(n1002), .A3(n[3310]), .Z(n1000) );
  XOR4D0 U901 ( .A1(n[3303]), .A2(n1003), .A3(n[3305]), .A4(n[3304]), .Z(n1002) );
  XOR4D0 U902 ( .A1(n[3298]), .A2(n[3297]), .A3(n1004), .A4(n1005), .Z(n1003)
         );
  XOR3D0 U903 ( .A1(n1006), .A2(n1007), .A3(n[3296]), .Z(n1005) );
  XOR4D0 U904 ( .A1(n[3289]), .A2(n1008), .A3(n[3291]), .A4(n[3290]), .Z(n1007) );
  XOR4D0 U905 ( .A1(n[3284]), .A2(n[3283]), .A3(n1009), .A4(n1010), .Z(n1008)
         );
  XOR3D0 U906 ( .A1(n1011), .A2(n1012), .A3(n[3282]), .Z(n1010) );
  XOR4D0 U907 ( .A1(n[3275]), .A2(n1013), .A3(n[3277]), .A4(n[3276]), .Z(n1012) );
  XOR4D0 U908 ( .A1(n[3270]), .A2(n[3269]), .A3(n1014), .A4(n1015), .Z(n1013)
         );
  XOR3D0 U909 ( .A1(n1016), .A2(n1017), .A3(n[3268]), .Z(n1015) );
  XOR4D0 U910 ( .A1(n[3261]), .A2(n1018), .A3(n[3263]), .A4(n[3262]), .Z(n1017) );
  XOR4D0 U911 ( .A1(n[3256]), .A2(n[3255]), .A3(n1019), .A4(n1020), .Z(n1018)
         );
  XOR3D0 U912 ( .A1(n1021), .A2(n1022), .A3(n[3254]), .Z(n1020) );
  XOR4D0 U913 ( .A1(n[3247]), .A2(n1023), .A3(n[3249]), .A4(n[3248]), .Z(n1022) );
  XOR4D0 U914 ( .A1(n[3242]), .A2(n[3241]), .A3(n1024), .A4(n1025), .Z(n1023)
         );
  XOR3D0 U915 ( .A1(n1026), .A2(n1027), .A3(n[3240]), .Z(n1025) );
  XOR4D0 U916 ( .A1(n[3233]), .A2(n1028), .A3(n[3235]), .A4(n[3234]), .Z(n1027) );
  XOR4D0 U917 ( .A1(n[3228]), .A2(n[3227]), .A3(n1029), .A4(n1030), .Z(n1028)
         );
  XOR3D0 U918 ( .A1(n1031), .A2(n1032), .A3(n[3226]), .Z(n1030) );
  XOR4D0 U919 ( .A1(n[3219]), .A2(n1033), .A3(n[3221]), .A4(n[3220]), .Z(n1032) );
  XOR4D0 U920 ( .A1(n[3214]), .A2(n[3213]), .A3(n1034), .A4(n1035), .Z(n1033)
         );
  XOR3D0 U921 ( .A1(n1036), .A2(n1037), .A3(n[3212]), .Z(n1035) );
  XOR4D0 U922 ( .A1(n[3205]), .A2(n1038), .A3(n[3207]), .A4(n[3206]), .Z(n1037) );
  XOR4D0 U923 ( .A1(n[3200]), .A2(n[3199]), .A3(n1039), .A4(n1040), .Z(n1038)
         );
  XOR3D0 U924 ( .A1(n1041), .A2(n1042), .A3(n[3198]), .Z(n1040) );
  XOR4D0 U925 ( .A1(n[3191]), .A2(n1043), .A3(n[3193]), .A4(n[3192]), .Z(n1042) );
  XOR4D0 U926 ( .A1(n[3186]), .A2(n[3185]), .A3(n1044), .A4(n1045), .Z(n1043)
         );
  XOR3D0 U927 ( .A1(n1046), .A2(n1047), .A3(n[3184]), .Z(n1045) );
  XOR4D0 U928 ( .A1(n[3177]), .A2(n1048), .A3(n[3179]), .A4(n[3178]), .Z(n1047) );
  XOR4D0 U929 ( .A1(n[3172]), .A2(n[3171]), .A3(n1049), .A4(n1050), .Z(n1048)
         );
  XOR3D0 U930 ( .A1(n1051), .A2(n1052), .A3(n[3170]), .Z(n1050) );
  XOR4D0 U931 ( .A1(n[3163]), .A2(n1053), .A3(n[3165]), .A4(n[3164]), .Z(n1052) );
  XOR4D0 U932 ( .A1(n[3158]), .A2(n[3157]), .A3(n1054), .A4(n1055), .Z(n1053)
         );
  XOR3D0 U933 ( .A1(n1056), .A2(n1057), .A3(n[3156]), .Z(n1055) );
  XOR4D0 U934 ( .A1(n[3149]), .A2(n1058), .A3(n[3151]), .A4(n[3150]), .Z(n1057) );
  XOR4D0 U935 ( .A1(n[3144]), .A2(n[3143]), .A3(n1059), .A4(n1060), .Z(n1058)
         );
  XOR3D0 U936 ( .A1(n1061), .A2(n1062), .A3(n[3142]), .Z(n1060) );
  XOR4D0 U937 ( .A1(n[3135]), .A2(n1063), .A3(n[3137]), .A4(n[3136]), .Z(n1062) );
  XOR4D0 U938 ( .A1(n[3130]), .A2(n[3129]), .A3(n1064), .A4(n1065), .Z(n1063)
         );
  XOR3D0 U939 ( .A1(n1066), .A2(n1067), .A3(n[3128]), .Z(n1065) );
  XOR4D0 U940 ( .A1(n[3121]), .A2(n1068), .A3(n[3123]), .A4(n[3122]), .Z(n1067) );
  XOR4D0 U941 ( .A1(n[3116]), .A2(n[3115]), .A3(n1069), .A4(n1070), .Z(n1068)
         );
  XOR3D0 U942 ( .A1(n1071), .A2(n1072), .A3(n[3114]), .Z(n1070) );
  XOR4D0 U943 ( .A1(n[3107]), .A2(n1073), .A3(n[3109]), .A4(n[3108]), .Z(n1072) );
  XOR4D0 U944 ( .A1(n[3102]), .A2(n[3101]), .A3(n1074), .A4(n1075), .Z(n1073)
         );
  XOR3D0 U945 ( .A1(n1076), .A2(n1077), .A3(n[3100]), .Z(n1075) );
  XOR4D0 U946 ( .A1(n[3093]), .A2(n1078), .A3(n[3095]), .A4(n[3094]), .Z(n1077) );
  XOR4D0 U947 ( .A1(n[3088]), .A2(n[3087]), .A3(n1079), .A4(n1080), .Z(n1078)
         );
  XOR3D0 U948 ( .A1(n1081), .A2(n1082), .A3(n[3086]), .Z(n1080) );
  XOR4D0 U949 ( .A1(n[3079]), .A2(n1083), .A3(n[3081]), .A4(n[3080]), .Z(n1082) );
  XOR4D0 U950 ( .A1(n[3074]), .A2(n[3073]), .A3(n1084), .A4(n1085), .Z(n1083)
         );
  XOR3D0 U951 ( .A1(n1086), .A2(n1087), .A3(n[3072]), .Z(n1085) );
  XOR4D0 U952 ( .A1(n[3065]), .A2(n1088), .A3(n[3067]), .A4(n[3066]), .Z(n1087) );
  XOR4D0 U953 ( .A1(n[3060]), .A2(n[3059]), .A3(n1089), .A4(n1090), .Z(n1088)
         );
  XOR3D0 U954 ( .A1(n1091), .A2(n1092), .A3(n[3058]), .Z(n1090) );
  XOR4D0 U955 ( .A1(n[3051]), .A2(n1093), .A3(n[3053]), .A4(n[3052]), .Z(n1092) );
  XOR4D0 U956 ( .A1(n[3046]), .A2(n[3045]), .A3(n1094), .A4(n1095), .Z(n1093)
         );
  XOR3D0 U957 ( .A1(n1096), .A2(n1097), .A3(n[3044]), .Z(n1095) );
  XOR4D0 U958 ( .A1(n[3037]), .A2(n1098), .A3(n[3039]), .A4(n[3038]), .Z(n1097) );
  XOR4D0 U959 ( .A1(n[3032]), .A2(n[3031]), .A3(n1099), .A4(n1100), .Z(n1098)
         );
  XOR3D0 U960 ( .A1(n1101), .A2(n1102), .A3(n[3030]), .Z(n1100) );
  XOR4D0 U961 ( .A1(n[3023]), .A2(n1103), .A3(n[3025]), .A4(n[3024]), .Z(n1102) );
  XOR4D0 U962 ( .A1(n[3018]), .A2(n[3017]), .A3(n1104), .A4(n1105), .Z(n1103)
         );
  XOR3D0 U963 ( .A1(n1106), .A2(n1107), .A3(n[3016]), .Z(n1105) );
  XOR4D0 U964 ( .A1(n[3009]), .A2(n1108), .A3(n[3011]), .A4(n[3010]), .Z(n1107) );
  XOR4D0 U965 ( .A1(n[3004]), .A2(n[3003]), .A3(n1109), .A4(n1110), .Z(n1108)
         );
  XOR3D0 U966 ( .A1(n1111), .A2(n1112), .A3(n[3002]), .Z(n1110) );
  XOR4D0 U967 ( .A1(n[2995]), .A2(n1113), .A3(n[2997]), .A4(n[2996]), .Z(n1112) );
  XOR4D0 U968 ( .A1(n[2990]), .A2(n[2989]), .A3(n1114), .A4(n1115), .Z(n1113)
         );
  XOR3D0 U969 ( .A1(n1116), .A2(n1117), .A3(n[2988]), .Z(n1115) );
  XOR4D0 U970 ( .A1(n[2981]), .A2(n1118), .A3(n[2983]), .A4(n[2982]), .Z(n1117) );
  XOR4D0 U971 ( .A1(n[2976]), .A2(n[2975]), .A3(n1119), .A4(n1120), .Z(n1118)
         );
  XOR3D0 U972 ( .A1(n1121), .A2(n1122), .A3(n[2974]), .Z(n1120) );
  XOR4D0 U973 ( .A1(n[2967]), .A2(n1123), .A3(n[2969]), .A4(n[2968]), .Z(n1122) );
  XOR4D0 U974 ( .A1(n[2962]), .A2(n[2961]), .A3(n1124), .A4(n1125), .Z(n1123)
         );
  XOR3D0 U975 ( .A1(n1126), .A2(n1127), .A3(n[2960]), .Z(n1125) );
  XOR4D0 U976 ( .A1(n[2953]), .A2(n1128), .A3(n[2955]), .A4(n[2954]), .Z(n1127) );
  XOR4D0 U977 ( .A1(n[2948]), .A2(n[2947]), .A3(n1129), .A4(n1130), .Z(n1128)
         );
  XOR3D0 U978 ( .A1(n1131), .A2(n1132), .A3(n[2946]), .Z(n1130) );
  XOR4D0 U979 ( .A1(n[2939]), .A2(n1133), .A3(n[2941]), .A4(n[2940]), .Z(n1132) );
  XOR4D0 U980 ( .A1(n[2934]), .A2(n[2933]), .A3(n1134), .A4(n1135), .Z(n1133)
         );
  XOR3D0 U981 ( .A1(n1136), .A2(n1137), .A3(n[2932]), .Z(n1135) );
  XOR4D0 U982 ( .A1(n[2925]), .A2(n1138), .A3(n[2927]), .A4(n[2926]), .Z(n1137) );
  XOR4D0 U983 ( .A1(n[2920]), .A2(n[2919]), .A3(n1139), .A4(n1140), .Z(n1138)
         );
  XOR3D0 U984 ( .A1(n1141), .A2(n1142), .A3(n[2918]), .Z(n1140) );
  XOR4D0 U985 ( .A1(n[2911]), .A2(n1143), .A3(n[2913]), .A4(n[2912]), .Z(n1142) );
  XOR4D0 U986 ( .A1(n[2906]), .A2(n[2905]), .A3(n1144), .A4(n1145), .Z(n1143)
         );
  XOR3D0 U987 ( .A1(n1146), .A2(n1147), .A3(n[2904]), .Z(n1145) );
  XOR4D0 U988 ( .A1(n[2897]), .A2(n1148), .A3(n[2899]), .A4(n[2898]), .Z(n1147) );
  XOR4D0 U989 ( .A1(n[2892]), .A2(n[2891]), .A3(n1149), .A4(n1150), .Z(n1148)
         );
  XOR3D0 U990 ( .A1(n1151), .A2(n1152), .A3(n[2890]), .Z(n1150) );
  XOR4D0 U991 ( .A1(n[2883]), .A2(n1153), .A3(n[2885]), .A4(n[2884]), .Z(n1152) );
  XOR4D0 U992 ( .A1(n[2878]), .A2(n[2877]), .A3(n1154), .A4(n1155), .Z(n1153)
         );
  XOR3D0 U993 ( .A1(n1156), .A2(n1157), .A3(n[2876]), .Z(n1155) );
  XOR4D0 U994 ( .A1(n[2869]), .A2(n1158), .A3(n[2871]), .A4(n[2870]), .Z(n1157) );
  XOR4D0 U995 ( .A1(n[2864]), .A2(n[2863]), .A3(n1159), .A4(n1160), .Z(n1158)
         );
  XOR3D0 U996 ( .A1(n1161), .A2(n1162), .A3(n[2862]), .Z(n1160) );
  XOR4D0 U997 ( .A1(n[2855]), .A2(n1163), .A3(n[2857]), .A4(n[2856]), .Z(n1162) );
  XOR4D0 U998 ( .A1(n[2850]), .A2(n[2849]), .A3(n1164), .A4(n1165), .Z(n1163)
         );
  XOR3D0 U999 ( .A1(n1166), .A2(n1167), .A3(n[2848]), .Z(n1165) );
  XOR4D0 U1000 ( .A1(n[2841]), .A2(n1168), .A3(n[2843]), .A4(n[2842]), .Z(
        n1167) );
  XOR4D0 U1001 ( .A1(n[2836]), .A2(n[2835]), .A3(n1169), .A4(n1170), .Z(n1168)
         );
  XOR3D0 U1002 ( .A1(n1171), .A2(n1172), .A3(n[2834]), .Z(n1170) );
  XOR4D0 U1003 ( .A1(n[2827]), .A2(n1173), .A3(n[2829]), .A4(n[2828]), .Z(
        n1172) );
  XOR4D0 U1004 ( .A1(n[2822]), .A2(n[2821]), .A3(n1174), .A4(n1175), .Z(n1173)
         );
  XOR3D0 U1005 ( .A1(n1176), .A2(n1177), .A3(n[2820]), .Z(n1175) );
  XOR4D0 U1006 ( .A1(n[2813]), .A2(n1178), .A3(n[2815]), .A4(n[2814]), .Z(
        n1177) );
  XOR4D0 U1007 ( .A1(n[2808]), .A2(n[2807]), .A3(n1179), .A4(n1180), .Z(n1178)
         );
  XOR3D0 U1008 ( .A1(n1181), .A2(n1182), .A3(n[2806]), .Z(n1180) );
  XOR4D0 U1009 ( .A1(n[2799]), .A2(n1183), .A3(n[2801]), .A4(n[2800]), .Z(
        n1182) );
  XOR4D0 U1010 ( .A1(n[2794]), .A2(n[2793]), .A3(n1184), .A4(n1185), .Z(n1183)
         );
  XOR3D0 U1011 ( .A1(n1186), .A2(n1187), .A3(n[2792]), .Z(n1185) );
  XOR4D0 U1012 ( .A1(n[2785]), .A2(n1188), .A3(n[2787]), .A4(n[2786]), .Z(
        n1187) );
  XOR4D0 U1013 ( .A1(n[2780]), .A2(n[2779]), .A3(n1189), .A4(n1190), .Z(n1188)
         );
  XOR3D0 U1014 ( .A1(n1191), .A2(n1192), .A3(n[2778]), .Z(n1190) );
  XOR4D0 U1015 ( .A1(n[2771]), .A2(n1193), .A3(n[2773]), .A4(n[2772]), .Z(
        n1192) );
  XOR4D0 U1016 ( .A1(n[2766]), .A2(n[2765]), .A3(n1194), .A4(n1195), .Z(n1193)
         );
  XOR3D0 U1017 ( .A1(n1196), .A2(n1197), .A3(n[2764]), .Z(n1195) );
  XOR4D0 U1018 ( .A1(n[2757]), .A2(n1198), .A3(n[2759]), .A4(n[2758]), .Z(
        n1197) );
  XOR4D0 U1019 ( .A1(n[2752]), .A2(n[2751]), .A3(n1199), .A4(n1200), .Z(n1198)
         );
  XOR3D0 U1020 ( .A1(n1201), .A2(n1202), .A3(n[2750]), .Z(n1200) );
  XOR4D0 U1021 ( .A1(n[2743]), .A2(n1203), .A3(n[2745]), .A4(n[2744]), .Z(
        n1202) );
  XOR4D0 U1022 ( .A1(n[2738]), .A2(n[2737]), .A3(n1204), .A4(n1205), .Z(n1203)
         );
  XOR3D0 U1023 ( .A1(n1206), .A2(n1207), .A3(n[2736]), .Z(n1205) );
  XOR4D0 U1024 ( .A1(n[2729]), .A2(n1208), .A3(n[2731]), .A4(n[2730]), .Z(
        n1207) );
  XOR4D0 U1025 ( .A1(n[2724]), .A2(n[2723]), .A3(n1209), .A4(n1210), .Z(n1208)
         );
  XOR3D0 U1026 ( .A1(n1211), .A2(n1212), .A3(n[2722]), .Z(n1210) );
  XOR4D0 U1027 ( .A1(n[2715]), .A2(n1213), .A3(n[2717]), .A4(n[2716]), .Z(
        n1212) );
  XOR4D0 U1028 ( .A1(n[2710]), .A2(n[2709]), .A3(n1214), .A4(n1215), .Z(n1213)
         );
  XOR3D0 U1029 ( .A1(n1216), .A2(n1217), .A3(n[2708]), .Z(n1215) );
  XOR4D0 U1030 ( .A1(n[2701]), .A2(n1218), .A3(n[2703]), .A4(n[2702]), .Z(
        n1217) );
  XOR4D0 U1031 ( .A1(n[2696]), .A2(n[2695]), .A3(n1219), .A4(n1220), .Z(n1218)
         );
  XOR3D0 U1032 ( .A1(n1221), .A2(n1222), .A3(n[2694]), .Z(n1220) );
  XOR4D0 U1033 ( .A1(n[2687]), .A2(n1223), .A3(n[2689]), .A4(n[2688]), .Z(
        n1222) );
  XOR4D0 U1034 ( .A1(n[2682]), .A2(n[2681]), .A3(n1224), .A4(n1225), .Z(n1223)
         );
  XOR3D0 U1035 ( .A1(n1226), .A2(n1227), .A3(n[2680]), .Z(n1225) );
  XOR4D0 U1036 ( .A1(n[2673]), .A2(n1228), .A3(n[2675]), .A4(n[2674]), .Z(
        n1227) );
  XOR4D0 U1037 ( .A1(n[2668]), .A2(n[2667]), .A3(n1229), .A4(n1230), .Z(n1228)
         );
  XOR3D0 U1038 ( .A1(n1231), .A2(n1232), .A3(n[2666]), .Z(n1230) );
  XOR4D0 U1039 ( .A1(n[2659]), .A2(n1233), .A3(n[2661]), .A4(n[2660]), .Z(
        n1232) );
  XOR4D0 U1040 ( .A1(n[2654]), .A2(n[2653]), .A3(n1234), .A4(n1235), .Z(n1233)
         );
  XOR3D0 U1041 ( .A1(n1236), .A2(n1237), .A3(n[2652]), .Z(n1235) );
  XOR4D0 U1042 ( .A1(n[2645]), .A2(n1238), .A3(n[2647]), .A4(n[2646]), .Z(
        n1237) );
  XOR4D0 U1043 ( .A1(n[2640]), .A2(n[2639]), .A3(n1239), .A4(n1240), .Z(n1238)
         );
  XOR3D0 U1044 ( .A1(n1241), .A2(n1242), .A3(n[2638]), .Z(n1240) );
  XOR4D0 U1045 ( .A1(n[2631]), .A2(n1243), .A3(n[2633]), .A4(n[2632]), .Z(
        n1242) );
  XOR4D0 U1046 ( .A1(n[2626]), .A2(n[2625]), .A3(n1244), .A4(n1245), .Z(n1243)
         );
  XOR3D0 U1047 ( .A1(n1246), .A2(n1247), .A3(n[2624]), .Z(n1245) );
  XOR4D0 U1048 ( .A1(n[2617]), .A2(n1248), .A3(n[2619]), .A4(n[2618]), .Z(
        n1247) );
  XOR4D0 U1049 ( .A1(n[2612]), .A2(n[2611]), .A3(n1249), .A4(n1250), .Z(n1248)
         );
  XOR3D0 U1050 ( .A1(n1251), .A2(n1252), .A3(n[2610]), .Z(n1250) );
  XOR4D0 U1051 ( .A1(n[2603]), .A2(n1253), .A3(n[2605]), .A4(n[2604]), .Z(
        n1252) );
  XOR4D0 U1052 ( .A1(n[2598]), .A2(n[2597]), .A3(n1254), .A4(n1255), .Z(n1253)
         );
  XOR3D0 U1053 ( .A1(n1256), .A2(n1257), .A3(n[2596]), .Z(n1255) );
  XOR4D0 U1054 ( .A1(n[2589]), .A2(n1258), .A3(n[2591]), .A4(n[2590]), .Z(
        n1257) );
  XOR4D0 U1055 ( .A1(n[2584]), .A2(n[2583]), .A3(n1259), .A4(n1260), .Z(n1258)
         );
  XOR3D0 U1056 ( .A1(n1261), .A2(n1262), .A3(n[2582]), .Z(n1260) );
  XOR4D0 U1057 ( .A1(n[2575]), .A2(n1263), .A3(n[2577]), .A4(n[2576]), .Z(
        n1262) );
  XOR4D0 U1058 ( .A1(n[2570]), .A2(n[2569]), .A3(n1264), .A4(n1265), .Z(n1263)
         );
  XOR3D0 U1059 ( .A1(n1266), .A2(n1267), .A3(n[2568]), .Z(n1265) );
  XOR4D0 U1060 ( .A1(n[2561]), .A2(n1268), .A3(n[2563]), .A4(n[2562]), .Z(
        n1267) );
  XOR4D0 U1061 ( .A1(n[2556]), .A2(n[2555]), .A3(n1269), .A4(n1270), .Z(n1268)
         );
  XOR3D0 U1062 ( .A1(n1271), .A2(n1272), .A3(n[2554]), .Z(n1270) );
  XOR4D0 U1063 ( .A1(n[2547]), .A2(n1273), .A3(n[2549]), .A4(n[2548]), .Z(
        n1272) );
  XOR4D0 U1064 ( .A1(n[2542]), .A2(n[2541]), .A3(n1274), .A4(n1275), .Z(n1273)
         );
  XOR3D0 U1065 ( .A1(n1276), .A2(n1277), .A3(n[2540]), .Z(n1275) );
  XOR4D0 U1066 ( .A1(n[2533]), .A2(n1278), .A3(n[2535]), .A4(n[2534]), .Z(
        n1277) );
  XOR4D0 U1067 ( .A1(n[2528]), .A2(n[2527]), .A3(n1279), .A4(n1280), .Z(n1278)
         );
  XOR3D0 U1068 ( .A1(n1281), .A2(n1282), .A3(n[2526]), .Z(n1280) );
  XOR4D0 U1069 ( .A1(n[2519]), .A2(n1283), .A3(n[2521]), .A4(n[2520]), .Z(
        n1282) );
  XOR4D0 U1070 ( .A1(n[2514]), .A2(n[2513]), .A3(n1284), .A4(n1285), .Z(n1283)
         );
  XOR3D0 U1071 ( .A1(n1286), .A2(n1287), .A3(n[2512]), .Z(n1285) );
  XOR4D0 U1072 ( .A1(n[2505]), .A2(n1288), .A3(n[2507]), .A4(n[2506]), .Z(
        n1287) );
  XOR4D0 U1073 ( .A1(n[2500]), .A2(n[2499]), .A3(n1289), .A4(n1290), .Z(n1288)
         );
  XOR3D0 U1074 ( .A1(n1291), .A2(n1292), .A3(n[2498]), .Z(n1290) );
  XOR4D0 U1075 ( .A1(n[2491]), .A2(n1293), .A3(n[2493]), .A4(n[2492]), .Z(
        n1292) );
  XOR4D0 U1076 ( .A1(n[2486]), .A2(n[2485]), .A3(n1294), .A4(n1295), .Z(n1293)
         );
  XOR3D0 U1077 ( .A1(n1296), .A2(n1297), .A3(n[2484]), .Z(n1295) );
  XOR4D0 U1078 ( .A1(n[2477]), .A2(n1298), .A3(n[2479]), .A4(n[2478]), .Z(
        n1297) );
  XOR4D0 U1079 ( .A1(n[2472]), .A2(n[2471]), .A3(n1299), .A4(n1300), .Z(n1298)
         );
  XOR3D0 U1080 ( .A1(n1301), .A2(n1302), .A3(n[2470]), .Z(n1300) );
  XOR4D0 U1081 ( .A1(n[2463]), .A2(n1303), .A3(n[2465]), .A4(n[2464]), .Z(
        n1302) );
  XOR4D0 U1082 ( .A1(n[2458]), .A2(n[2457]), .A3(n1304), .A4(n1305), .Z(n1303)
         );
  XOR3D0 U1083 ( .A1(n1306), .A2(n1307), .A3(n[2456]), .Z(n1305) );
  XOR4D0 U1084 ( .A1(n[2449]), .A2(n1308), .A3(n[2451]), .A4(n[2450]), .Z(
        n1307) );
  XOR4D0 U1085 ( .A1(n[2444]), .A2(n[2443]), .A3(n1309), .A4(n1310), .Z(n1308)
         );
  XOR3D0 U1086 ( .A1(n1311), .A2(n1312), .A3(n[2442]), .Z(n1310) );
  XOR4D0 U1087 ( .A1(n[2435]), .A2(n1313), .A3(n[2437]), .A4(n[2436]), .Z(
        n1312) );
  XOR4D0 U1088 ( .A1(n[2430]), .A2(n[2429]), .A3(n1314), .A4(n1315), .Z(n1313)
         );
  XOR3D0 U1089 ( .A1(n1316), .A2(n1317), .A3(n[2428]), .Z(n1315) );
  XOR4D0 U1090 ( .A1(n[2421]), .A2(n1318), .A3(n[2423]), .A4(n[2422]), .Z(
        n1317) );
  XOR4D0 U1091 ( .A1(n[2416]), .A2(n[2415]), .A3(n1319), .A4(n1320), .Z(n1318)
         );
  XOR3D0 U1092 ( .A1(n1321), .A2(n1322), .A3(n[2414]), .Z(n1320) );
  XOR4D0 U1093 ( .A1(n[2407]), .A2(n1323), .A3(n[2409]), .A4(n[2408]), .Z(
        n1322) );
  XOR4D0 U1094 ( .A1(n[2402]), .A2(n[2401]), .A3(n1324), .A4(n1325), .Z(n1323)
         );
  XOR3D0 U1095 ( .A1(n1326), .A2(n1327), .A3(n[2400]), .Z(n1325) );
  XOR4D0 U1096 ( .A1(n[2393]), .A2(n1328), .A3(n[2395]), .A4(n[2394]), .Z(
        n1327) );
  XOR4D0 U1097 ( .A1(n[2388]), .A2(n[2387]), .A3(n1329), .A4(n1330), .Z(n1328)
         );
  XOR3D0 U1098 ( .A1(n1331), .A2(n1332), .A3(n[2386]), .Z(n1330) );
  XOR4D0 U1099 ( .A1(n[2379]), .A2(n1333), .A3(n[2381]), .A4(n[2380]), .Z(
        n1332) );
  XOR4D0 U1100 ( .A1(n[2374]), .A2(n[2373]), .A3(n1334), .A4(n1335), .Z(n1333)
         );
  XOR3D0 U1101 ( .A1(n1336), .A2(n1337), .A3(n[2372]), .Z(n1335) );
  XOR4D0 U1102 ( .A1(n[2365]), .A2(n1338), .A3(n[2367]), .A4(n[2366]), .Z(
        n1337) );
  XOR4D0 U1103 ( .A1(n[2360]), .A2(n[2359]), .A3(n1339), .A4(n1340), .Z(n1338)
         );
  XOR3D0 U1104 ( .A1(n1341), .A2(n1342), .A3(n[2358]), .Z(n1340) );
  XOR4D0 U1105 ( .A1(n[2351]), .A2(n1343), .A3(n[2353]), .A4(n[2352]), .Z(
        n1342) );
  XOR4D0 U1106 ( .A1(n[2346]), .A2(n[2345]), .A3(n1344), .A4(n1345), .Z(n1343)
         );
  XOR3D0 U1107 ( .A1(n1346), .A2(n1347), .A3(n[2344]), .Z(n1345) );
  XOR4D0 U1108 ( .A1(n[2337]), .A2(n1348), .A3(n[2339]), .A4(n[2338]), .Z(
        n1347) );
  XOR4D0 U1109 ( .A1(n[2332]), .A2(n[2331]), .A3(n1349), .A4(n1350), .Z(n1348)
         );
  XOR3D0 U1110 ( .A1(n1351), .A2(n1352), .A3(n[2330]), .Z(n1350) );
  XOR4D0 U1111 ( .A1(n[2323]), .A2(n1353), .A3(n[2325]), .A4(n[2324]), .Z(
        n1352) );
  XOR4D0 U1112 ( .A1(n[2318]), .A2(n[2317]), .A3(n1354), .A4(n1355), .Z(n1353)
         );
  XOR3D0 U1113 ( .A1(n1356), .A2(n1357), .A3(n[2316]), .Z(n1355) );
  XOR4D0 U1114 ( .A1(n[2309]), .A2(n1358), .A3(n[2311]), .A4(n[2310]), .Z(
        n1357) );
  XOR4D0 U1115 ( .A1(n[2304]), .A2(n[2303]), .A3(n1359), .A4(n1360), .Z(n1358)
         );
  XOR3D0 U1116 ( .A1(n1361), .A2(n1362), .A3(n[2302]), .Z(n1360) );
  XOR4D0 U1117 ( .A1(n[2295]), .A2(n1363), .A3(n[2297]), .A4(n[2296]), .Z(
        n1362) );
  XOR4D0 U1118 ( .A1(n[2290]), .A2(n[2289]), .A3(n1364), .A4(n1365), .Z(n1363)
         );
  XOR3D0 U1119 ( .A1(n1366), .A2(n1367), .A3(n[2288]), .Z(n1365) );
  XOR4D0 U1120 ( .A1(n[2281]), .A2(n1368), .A3(n[2283]), .A4(n[2282]), .Z(
        n1367) );
  XOR4D0 U1121 ( .A1(n[2276]), .A2(n[2275]), .A3(n1369), .A4(n1370), .Z(n1368)
         );
  XOR3D0 U1122 ( .A1(n1371), .A2(n1372), .A3(n[2274]), .Z(n1370) );
  XOR4D0 U1123 ( .A1(n[2267]), .A2(n1373), .A3(n[2269]), .A4(n[2268]), .Z(
        n1372) );
  XOR4D0 U1124 ( .A1(n[2262]), .A2(n[2261]), .A3(n1374), .A4(n1375), .Z(n1373)
         );
  XOR3D0 U1125 ( .A1(n1376), .A2(n1377), .A3(n[2260]), .Z(n1375) );
  XOR4D0 U1126 ( .A1(n[2253]), .A2(n1378), .A3(n[2255]), .A4(n[2254]), .Z(
        n1377) );
  XOR4D0 U1127 ( .A1(n[2248]), .A2(n[2247]), .A3(n1379), .A4(n1380), .Z(n1378)
         );
  XOR3D0 U1128 ( .A1(n1381), .A2(n1382), .A3(n[2246]), .Z(n1380) );
  XOR4D0 U1129 ( .A1(n[2239]), .A2(n1383), .A3(n[2241]), .A4(n[2240]), .Z(
        n1382) );
  XOR4D0 U1130 ( .A1(n[2234]), .A2(n[2233]), .A3(n1384), .A4(n1385), .Z(n1383)
         );
  XOR3D0 U1131 ( .A1(n1386), .A2(n1387), .A3(n[2232]), .Z(n1385) );
  XOR4D0 U1132 ( .A1(n[2225]), .A2(n1388), .A3(n[2227]), .A4(n[2226]), .Z(
        n1387) );
  XOR4D0 U1133 ( .A1(n[2220]), .A2(n[2219]), .A3(n1389), .A4(n1390), .Z(n1388)
         );
  XOR3D0 U1134 ( .A1(n1391), .A2(n1392), .A3(n[2218]), .Z(n1390) );
  XOR4D0 U1135 ( .A1(n[2211]), .A2(n1393), .A3(n[2213]), .A4(n[2212]), .Z(
        n1392) );
  XOR4D0 U1136 ( .A1(n[2206]), .A2(n[2205]), .A3(n1394), .A4(n1395), .Z(n1393)
         );
  XOR3D0 U1137 ( .A1(n1396), .A2(n1397), .A3(n[2204]), .Z(n1395) );
  XOR4D0 U1138 ( .A1(n[2197]), .A2(n1398), .A3(n[2199]), .A4(n[2198]), .Z(
        n1397) );
  XOR4D0 U1139 ( .A1(n[2192]), .A2(n[2191]), .A3(n1399), .A4(n1400), .Z(n1398)
         );
  XOR3D0 U1140 ( .A1(n1401), .A2(n1402), .A3(n[2190]), .Z(n1400) );
  XOR4D0 U1141 ( .A1(n[2183]), .A2(n1403), .A3(n[2185]), .A4(n[2184]), .Z(
        n1402) );
  XOR4D0 U1142 ( .A1(n[2178]), .A2(n[2177]), .A3(n1404), .A4(n1405), .Z(n1403)
         );
  XOR3D0 U1143 ( .A1(n1406), .A2(n1407), .A3(n[2176]), .Z(n1405) );
  XOR4D0 U1144 ( .A1(n[2169]), .A2(n1408), .A3(n[2171]), .A4(n[2170]), .Z(
        n1407) );
  XOR4D0 U1145 ( .A1(n[2164]), .A2(n[2163]), .A3(n1409), .A4(n1410), .Z(n1408)
         );
  XOR3D0 U1146 ( .A1(n1411), .A2(n1412), .A3(n[2162]), .Z(n1410) );
  XOR4D0 U1147 ( .A1(n[2155]), .A2(n1413), .A3(n[2157]), .A4(n[2156]), .Z(
        n1412) );
  XOR4D0 U1148 ( .A1(n[2150]), .A2(n[2149]), .A3(n1414), .A4(n1415), .Z(n1413)
         );
  XOR3D0 U1149 ( .A1(n1416), .A2(n1417), .A3(n[2148]), .Z(n1415) );
  XOR4D0 U1150 ( .A1(n[2141]), .A2(n1418), .A3(n[2143]), .A4(n[2142]), .Z(
        n1417) );
  XOR4D0 U1151 ( .A1(n[2136]), .A2(n[2135]), .A3(n1419), .A4(n1420), .Z(n1418)
         );
  XOR3D0 U1152 ( .A1(n1421), .A2(n1422), .A3(n[2134]), .Z(n1420) );
  XOR4D0 U1153 ( .A1(n[2127]), .A2(n1423), .A3(n[2129]), .A4(n[2128]), .Z(
        n1422) );
  XOR4D0 U1154 ( .A1(n[2122]), .A2(n[2121]), .A3(n1424), .A4(n1425), .Z(n1423)
         );
  XOR3D0 U1155 ( .A1(n1426), .A2(n1427), .A3(n[2120]), .Z(n1425) );
  XOR4D0 U1156 ( .A1(n[2113]), .A2(n1428), .A3(n[2115]), .A4(n[2114]), .Z(
        n1427) );
  XOR4D0 U1157 ( .A1(n[2108]), .A2(n[2107]), .A3(n1429), .A4(n1430), .Z(n1428)
         );
  XOR3D0 U1158 ( .A1(n1431), .A2(n1432), .A3(n[2106]), .Z(n1430) );
  XOR4D0 U1159 ( .A1(n[2099]), .A2(n1433), .A3(n[2101]), .A4(n[2100]), .Z(
        n1432) );
  XOR4D0 U1160 ( .A1(n[2094]), .A2(n[2093]), .A3(n1434), .A4(n1435), .Z(n1433)
         );
  XOR3D0 U1161 ( .A1(n1436), .A2(n1437), .A3(n[2092]), .Z(n1435) );
  XOR4D0 U1162 ( .A1(n[2085]), .A2(n1438), .A3(n[2087]), .A4(n[2086]), .Z(
        n1437) );
  XOR4D0 U1163 ( .A1(n[2080]), .A2(n[2079]), .A3(n1439), .A4(n1440), .Z(n1438)
         );
  XOR3D0 U1164 ( .A1(n1441), .A2(n1442), .A3(n[2078]), .Z(n1440) );
  XOR4D0 U1165 ( .A1(n[2071]), .A2(n1443), .A3(n[2073]), .A4(n[2072]), .Z(
        n1442) );
  XOR4D0 U1166 ( .A1(n[2066]), .A2(n[2065]), .A3(n1444), .A4(n1445), .Z(n1443)
         );
  XOR3D0 U1167 ( .A1(n1446), .A2(n1447), .A3(n[2064]), .Z(n1445) );
  XOR4D0 U1168 ( .A1(n[2057]), .A2(n1448), .A3(n[2059]), .A4(n[2058]), .Z(
        n1447) );
  XOR4D0 U1169 ( .A1(n[2052]), .A2(n[2051]), .A3(n1449), .A4(n1450), .Z(n1448)
         );
  XOR3D0 U1170 ( .A1(n1451), .A2(n1452), .A3(n[2050]), .Z(n1450) );
  XOR3D0 U1171 ( .A1(n[2045]), .A2(n[2044]), .A3(n1453), .Z(n1452) );
  XOR3D0 U1172 ( .A1(n1454), .A2(n1455), .A3(n[2043]), .Z(n1453) );
  XOR4D0 U1173 ( .A1(n[2036]), .A2(n[2035]), .A3(n[2038]), .A4(n[2037]), .Z(
        n1455) );
  XOR4D0 U1174 ( .A1(n[2040]), .A2(n[2039]), .A3(n[2042]), .A4(n[2041]), .Z(
        n1454) );
  XOR4D0 U1175 ( .A1(n[2047]), .A2(n[2046]), .A3(n[2049]), .A4(n[2048]), .Z(
        n1451) );
  XOR4D0 U1176 ( .A1(n[2054]), .A2(n[2053]), .A3(n[2056]), .A4(n[2055]), .Z(
        n1449) );
  XOR4D0 U1177 ( .A1(n[2061]), .A2(n[2060]), .A3(n[2063]), .A4(n[2062]), .Z(
        n1446) );
  XOR4D0 U1178 ( .A1(n[2068]), .A2(n[2067]), .A3(n[2070]), .A4(n[2069]), .Z(
        n1444) );
  XOR4D0 U1179 ( .A1(n[2075]), .A2(n[2074]), .A3(n[2077]), .A4(n[2076]), .Z(
        n1441) );
  XOR4D0 U1180 ( .A1(n[2082]), .A2(n[2081]), .A3(n[2084]), .A4(n[2083]), .Z(
        n1439) );
  XOR4D0 U1181 ( .A1(n[2089]), .A2(n[2088]), .A3(n[2091]), .A4(n[2090]), .Z(
        n1436) );
  XOR4D0 U1182 ( .A1(n[2096]), .A2(n[2095]), .A3(n[2098]), .A4(n[2097]), .Z(
        n1434) );
  XOR4D0 U1183 ( .A1(n[2103]), .A2(n[2102]), .A3(n[2105]), .A4(n[2104]), .Z(
        n1431) );
  XOR4D0 U1184 ( .A1(n[2110]), .A2(n[2109]), .A3(n[2112]), .A4(n[2111]), .Z(
        n1429) );
  XOR4D0 U1185 ( .A1(n[2117]), .A2(n[2116]), .A3(n[2119]), .A4(n[2118]), .Z(
        n1426) );
  XOR4D0 U1186 ( .A1(n[2124]), .A2(n[2123]), .A3(n[2126]), .A4(n[2125]), .Z(
        n1424) );
  XOR4D0 U1187 ( .A1(n[2131]), .A2(n[2130]), .A3(n[2133]), .A4(n[2132]), .Z(
        n1421) );
  XOR4D0 U1188 ( .A1(n[2138]), .A2(n[2137]), .A3(n[2140]), .A4(n[2139]), .Z(
        n1419) );
  XOR4D0 U1189 ( .A1(n[2145]), .A2(n[2144]), .A3(n[2147]), .A4(n[2146]), .Z(
        n1416) );
  XOR4D0 U1190 ( .A1(n[2152]), .A2(n[2151]), .A3(n[2154]), .A4(n[2153]), .Z(
        n1414) );
  XOR4D0 U1191 ( .A1(n[2159]), .A2(n[2158]), .A3(n[2161]), .A4(n[2160]), .Z(
        n1411) );
  XOR4D0 U1192 ( .A1(n[2166]), .A2(n[2165]), .A3(n[2168]), .A4(n[2167]), .Z(
        n1409) );
  XOR4D0 U1193 ( .A1(n[2173]), .A2(n[2172]), .A3(n[2175]), .A4(n[2174]), .Z(
        n1406) );
  XOR4D0 U1194 ( .A1(n[2180]), .A2(n[2179]), .A3(n[2182]), .A4(n[2181]), .Z(
        n1404) );
  XOR4D0 U1195 ( .A1(n[2187]), .A2(n[2186]), .A3(n[2189]), .A4(n[2188]), .Z(
        n1401) );
  XOR4D0 U1196 ( .A1(n[2194]), .A2(n[2193]), .A3(n[2196]), .A4(n[2195]), .Z(
        n1399) );
  XOR4D0 U1197 ( .A1(n[2201]), .A2(n[2200]), .A3(n[2203]), .A4(n[2202]), .Z(
        n1396) );
  XOR4D0 U1198 ( .A1(n[2208]), .A2(n[2207]), .A3(n[2210]), .A4(n[2209]), .Z(
        n1394) );
  XOR4D0 U1199 ( .A1(n[2215]), .A2(n[2214]), .A3(n[2217]), .A4(n[2216]), .Z(
        n1391) );
  XOR4D0 U1200 ( .A1(n[2222]), .A2(n[2221]), .A3(n[2224]), .A4(n[2223]), .Z(
        n1389) );
  XOR4D0 U1201 ( .A1(n[2229]), .A2(n[2228]), .A3(n[2231]), .A4(n[2230]), .Z(
        n1386) );
  XOR4D0 U1202 ( .A1(n[2236]), .A2(n[2235]), .A3(n[2238]), .A4(n[2237]), .Z(
        n1384) );
  XOR4D0 U1203 ( .A1(n[2243]), .A2(n[2242]), .A3(n[2245]), .A4(n[2244]), .Z(
        n1381) );
  XOR4D0 U1204 ( .A1(n[2250]), .A2(n[2249]), .A3(n[2252]), .A4(n[2251]), .Z(
        n1379) );
  XOR4D0 U1205 ( .A1(n[2257]), .A2(n[2256]), .A3(n[2259]), .A4(n[2258]), .Z(
        n1376) );
  XOR4D0 U1206 ( .A1(n[2264]), .A2(n[2263]), .A3(n[2266]), .A4(n[2265]), .Z(
        n1374) );
  XOR4D0 U1207 ( .A1(n[2271]), .A2(n[2270]), .A3(n[2273]), .A4(n[2272]), .Z(
        n1371) );
  XOR4D0 U1208 ( .A1(n[2278]), .A2(n[2277]), .A3(n[2280]), .A4(n[2279]), .Z(
        n1369) );
  XOR4D0 U1209 ( .A1(n[2285]), .A2(n[2284]), .A3(n[2287]), .A4(n[2286]), .Z(
        n1366) );
  XOR4D0 U1210 ( .A1(n[2292]), .A2(n[2291]), .A3(n[2294]), .A4(n[2293]), .Z(
        n1364) );
  XOR4D0 U1211 ( .A1(n[2299]), .A2(n[2298]), .A3(n[2301]), .A4(n[2300]), .Z(
        n1361) );
  XOR4D0 U1212 ( .A1(n[2306]), .A2(n[2305]), .A3(n[2308]), .A4(n[2307]), .Z(
        n1359) );
  XOR4D0 U1213 ( .A1(n[2313]), .A2(n[2312]), .A3(n[2315]), .A4(n[2314]), .Z(
        n1356) );
  XOR4D0 U1214 ( .A1(n[2320]), .A2(n[2319]), .A3(n[2322]), .A4(n[2321]), .Z(
        n1354) );
  XOR4D0 U1215 ( .A1(n[2327]), .A2(n[2326]), .A3(n[2329]), .A4(n[2328]), .Z(
        n1351) );
  XOR4D0 U1216 ( .A1(n[2334]), .A2(n[2333]), .A3(n[2336]), .A4(n[2335]), .Z(
        n1349) );
  XOR4D0 U1217 ( .A1(n[2341]), .A2(n[2340]), .A3(n[2343]), .A4(n[2342]), .Z(
        n1346) );
  XOR4D0 U1218 ( .A1(n[2348]), .A2(n[2347]), .A3(n[2350]), .A4(n[2349]), .Z(
        n1344) );
  XOR4D0 U1219 ( .A1(n[2355]), .A2(n[2354]), .A3(n[2357]), .A4(n[2356]), .Z(
        n1341) );
  XOR4D0 U1220 ( .A1(n[2362]), .A2(n[2361]), .A3(n[2364]), .A4(n[2363]), .Z(
        n1339) );
  XOR4D0 U1221 ( .A1(n[2369]), .A2(n[2368]), .A3(n[2371]), .A4(n[2370]), .Z(
        n1336) );
  XOR4D0 U1222 ( .A1(n[2376]), .A2(n[2375]), .A3(n[2378]), .A4(n[2377]), .Z(
        n1334) );
  XOR4D0 U1223 ( .A1(n[2383]), .A2(n[2382]), .A3(n[2385]), .A4(n[2384]), .Z(
        n1331) );
  XOR4D0 U1224 ( .A1(n[2390]), .A2(n[2389]), .A3(n[2392]), .A4(n[2391]), .Z(
        n1329) );
  XOR4D0 U1225 ( .A1(n[2397]), .A2(n[2396]), .A3(n[2399]), .A4(n[2398]), .Z(
        n1326) );
  XOR4D0 U1226 ( .A1(n[2404]), .A2(n[2403]), .A3(n[2406]), .A4(n[2405]), .Z(
        n1324) );
  XOR4D0 U1227 ( .A1(n[2411]), .A2(n[2410]), .A3(n[2413]), .A4(n[2412]), .Z(
        n1321) );
  XOR4D0 U1228 ( .A1(n[2418]), .A2(n[2417]), .A3(n[2420]), .A4(n[2419]), .Z(
        n1319) );
  XOR4D0 U1229 ( .A1(n[2425]), .A2(n[2424]), .A3(n[2427]), .A4(n[2426]), .Z(
        n1316) );
  XOR4D0 U1230 ( .A1(n[2432]), .A2(n[2431]), .A3(n[2434]), .A4(n[2433]), .Z(
        n1314) );
  XOR4D0 U1231 ( .A1(n[2439]), .A2(n[2438]), .A3(n[2441]), .A4(n[2440]), .Z(
        n1311) );
  XOR4D0 U1232 ( .A1(n[2446]), .A2(n[2445]), .A3(n[2448]), .A4(n[2447]), .Z(
        n1309) );
  XOR4D0 U1233 ( .A1(n[2453]), .A2(n[2452]), .A3(n[2455]), .A4(n[2454]), .Z(
        n1306) );
  XOR4D0 U1234 ( .A1(n[2460]), .A2(n[2459]), .A3(n[2462]), .A4(n[2461]), .Z(
        n1304) );
  XOR4D0 U1235 ( .A1(n[2467]), .A2(n[2466]), .A3(n[2469]), .A4(n[2468]), .Z(
        n1301) );
  XOR4D0 U1236 ( .A1(n[2474]), .A2(n[2473]), .A3(n[2476]), .A4(n[2475]), .Z(
        n1299) );
  XOR4D0 U1237 ( .A1(n[2481]), .A2(n[2480]), .A3(n[2483]), .A4(n[2482]), .Z(
        n1296) );
  XOR4D0 U1238 ( .A1(n[2488]), .A2(n[2487]), .A3(n[2490]), .A4(n[2489]), .Z(
        n1294) );
  XOR4D0 U1239 ( .A1(n[2495]), .A2(n[2494]), .A3(n[2497]), .A4(n[2496]), .Z(
        n1291) );
  XOR4D0 U1240 ( .A1(n[2502]), .A2(n[2501]), .A3(n[2504]), .A4(n[2503]), .Z(
        n1289) );
  XOR4D0 U1241 ( .A1(n[2509]), .A2(n[2508]), .A3(n[2511]), .A4(n[2510]), .Z(
        n1286) );
  XOR4D0 U1242 ( .A1(n[2516]), .A2(n[2515]), .A3(n[2518]), .A4(n[2517]), .Z(
        n1284) );
  XOR4D0 U1243 ( .A1(n[2523]), .A2(n[2522]), .A3(n[2525]), .A4(n[2524]), .Z(
        n1281) );
  XOR4D0 U1244 ( .A1(n[2530]), .A2(n[2529]), .A3(n[2532]), .A4(n[2531]), .Z(
        n1279) );
  XOR4D0 U1245 ( .A1(n[2537]), .A2(n[2536]), .A3(n[2539]), .A4(n[2538]), .Z(
        n1276) );
  XOR4D0 U1246 ( .A1(n[2544]), .A2(n[2543]), .A3(n[2546]), .A4(n[2545]), .Z(
        n1274) );
  XOR4D0 U1247 ( .A1(n[2551]), .A2(n[2550]), .A3(n[2553]), .A4(n[2552]), .Z(
        n1271) );
  XOR4D0 U1248 ( .A1(n[2558]), .A2(n[2557]), .A3(n[2560]), .A4(n[2559]), .Z(
        n1269) );
  XOR4D0 U1249 ( .A1(n[2565]), .A2(n[2564]), .A3(n[2567]), .A4(n[2566]), .Z(
        n1266) );
  XOR4D0 U1250 ( .A1(n[2572]), .A2(n[2571]), .A3(n[2574]), .A4(n[2573]), .Z(
        n1264) );
  XOR4D0 U1251 ( .A1(n[2579]), .A2(n[2578]), .A3(n[2581]), .A4(n[2580]), .Z(
        n1261) );
  XOR4D0 U1252 ( .A1(n[2586]), .A2(n[2585]), .A3(n[2588]), .A4(n[2587]), .Z(
        n1259) );
  XOR4D0 U1253 ( .A1(n[2593]), .A2(n[2592]), .A3(n[2595]), .A4(n[2594]), .Z(
        n1256) );
  XOR4D0 U1254 ( .A1(n[2600]), .A2(n[2599]), .A3(n[2602]), .A4(n[2601]), .Z(
        n1254) );
  XOR4D0 U1255 ( .A1(n[2607]), .A2(n[2606]), .A3(n[2609]), .A4(n[2608]), .Z(
        n1251) );
  XOR4D0 U1256 ( .A1(n[2614]), .A2(n[2613]), .A3(n[2616]), .A4(n[2615]), .Z(
        n1249) );
  XOR4D0 U1257 ( .A1(n[2621]), .A2(n[2620]), .A3(n[2623]), .A4(n[2622]), .Z(
        n1246) );
  XOR4D0 U1258 ( .A1(n[2628]), .A2(n[2627]), .A3(n[2630]), .A4(n[2629]), .Z(
        n1244) );
  XOR4D0 U1259 ( .A1(n[2635]), .A2(n[2634]), .A3(n[2637]), .A4(n[2636]), .Z(
        n1241) );
  XOR4D0 U1260 ( .A1(n[2642]), .A2(n[2641]), .A3(n[2644]), .A4(n[2643]), .Z(
        n1239) );
  XOR4D0 U1261 ( .A1(n[2649]), .A2(n[2648]), .A3(n[2651]), .A4(n[2650]), .Z(
        n1236) );
  XOR4D0 U1262 ( .A1(n[2656]), .A2(n[2655]), .A3(n[2658]), .A4(n[2657]), .Z(
        n1234) );
  XOR4D0 U1263 ( .A1(n[2663]), .A2(n[2662]), .A3(n[2665]), .A4(n[2664]), .Z(
        n1231) );
  XOR4D0 U1264 ( .A1(n[2670]), .A2(n[2669]), .A3(n[2672]), .A4(n[2671]), .Z(
        n1229) );
  XOR4D0 U1265 ( .A1(n[2677]), .A2(n[2676]), .A3(n[2679]), .A4(n[2678]), .Z(
        n1226) );
  XOR4D0 U1266 ( .A1(n[2684]), .A2(n[2683]), .A3(n[2686]), .A4(n[2685]), .Z(
        n1224) );
  XOR4D0 U1267 ( .A1(n[2691]), .A2(n[2690]), .A3(n[2693]), .A4(n[2692]), .Z(
        n1221) );
  XOR4D0 U1268 ( .A1(n[2698]), .A2(n[2697]), .A3(n[2700]), .A4(n[2699]), .Z(
        n1219) );
  XOR4D0 U1269 ( .A1(n[2705]), .A2(n[2704]), .A3(n[2707]), .A4(n[2706]), .Z(
        n1216) );
  XOR4D0 U1270 ( .A1(n[2712]), .A2(n[2711]), .A3(n[2714]), .A4(n[2713]), .Z(
        n1214) );
  XOR4D0 U1271 ( .A1(n[2719]), .A2(n[2718]), .A3(n[2721]), .A4(n[2720]), .Z(
        n1211) );
  XOR4D0 U1272 ( .A1(n[2726]), .A2(n[2725]), .A3(n[2728]), .A4(n[2727]), .Z(
        n1209) );
  XOR4D0 U1273 ( .A1(n[2733]), .A2(n[2732]), .A3(n[2735]), .A4(n[2734]), .Z(
        n1206) );
  XOR4D0 U1274 ( .A1(n[2740]), .A2(n[2739]), .A3(n[2742]), .A4(n[2741]), .Z(
        n1204) );
  XOR4D0 U1275 ( .A1(n[2747]), .A2(n[2746]), .A3(n[2749]), .A4(n[2748]), .Z(
        n1201) );
  XOR4D0 U1276 ( .A1(n[2754]), .A2(n[2753]), .A3(n[2756]), .A4(n[2755]), .Z(
        n1199) );
  XOR4D0 U1277 ( .A1(n[2761]), .A2(n[2760]), .A3(n[2763]), .A4(n[2762]), .Z(
        n1196) );
  XOR4D0 U1278 ( .A1(n[2768]), .A2(n[2767]), .A3(n[2770]), .A4(n[2769]), .Z(
        n1194) );
  XOR4D0 U1279 ( .A1(n[2775]), .A2(n[2774]), .A3(n[2777]), .A4(n[2776]), .Z(
        n1191) );
  XOR4D0 U1280 ( .A1(n[2782]), .A2(n[2781]), .A3(n[2784]), .A4(n[2783]), .Z(
        n1189) );
  XOR4D0 U1281 ( .A1(n[2789]), .A2(n[2788]), .A3(n[2791]), .A4(n[2790]), .Z(
        n1186) );
  XOR4D0 U1282 ( .A1(n[2796]), .A2(n[2795]), .A3(n[2798]), .A4(n[2797]), .Z(
        n1184) );
  XOR4D0 U1283 ( .A1(n[2803]), .A2(n[2802]), .A3(n[2805]), .A4(n[2804]), .Z(
        n1181) );
  XOR4D0 U1284 ( .A1(n[2810]), .A2(n[2809]), .A3(n[2812]), .A4(n[2811]), .Z(
        n1179) );
  XOR4D0 U1285 ( .A1(n[2817]), .A2(n[2816]), .A3(n[2819]), .A4(n[2818]), .Z(
        n1176) );
  XOR4D0 U1286 ( .A1(n[2824]), .A2(n[2823]), .A3(n[2826]), .A4(n[2825]), .Z(
        n1174) );
  XOR4D0 U1287 ( .A1(n[2831]), .A2(n[2830]), .A3(n[2833]), .A4(n[2832]), .Z(
        n1171) );
  XOR4D0 U1288 ( .A1(n[2838]), .A2(n[2837]), .A3(n[2840]), .A4(n[2839]), .Z(
        n1169) );
  XOR4D0 U1289 ( .A1(n[2845]), .A2(n[2844]), .A3(n[2847]), .A4(n[2846]), .Z(
        n1166) );
  XOR4D0 U1290 ( .A1(n[2852]), .A2(n[2851]), .A3(n[2854]), .A4(n[2853]), .Z(
        n1164) );
  XOR4D0 U1291 ( .A1(n[2859]), .A2(n[2858]), .A3(n[2861]), .A4(n[2860]), .Z(
        n1161) );
  XOR4D0 U1292 ( .A1(n[2866]), .A2(n[2865]), .A3(n[2868]), .A4(n[2867]), .Z(
        n1159) );
  XOR4D0 U1293 ( .A1(n[2873]), .A2(n[2872]), .A3(n[2875]), .A4(n[2874]), .Z(
        n1156) );
  XOR4D0 U1294 ( .A1(n[2880]), .A2(n[2879]), .A3(n[2882]), .A4(n[2881]), .Z(
        n1154) );
  XOR4D0 U1295 ( .A1(n[2887]), .A2(n[2886]), .A3(n[2889]), .A4(n[2888]), .Z(
        n1151) );
  XOR4D0 U1296 ( .A1(n[2894]), .A2(n[2893]), .A3(n[2896]), .A4(n[2895]), .Z(
        n1149) );
  XOR4D0 U1297 ( .A1(n[2901]), .A2(n[2900]), .A3(n[2903]), .A4(n[2902]), .Z(
        n1146) );
  XOR4D0 U1298 ( .A1(n[2908]), .A2(n[2907]), .A3(n[2910]), .A4(n[2909]), .Z(
        n1144) );
  XOR4D0 U1299 ( .A1(n[2915]), .A2(n[2914]), .A3(n[2917]), .A4(n[2916]), .Z(
        n1141) );
  XOR4D0 U1300 ( .A1(n[2922]), .A2(n[2921]), .A3(n[2924]), .A4(n[2923]), .Z(
        n1139) );
  XOR4D0 U1301 ( .A1(n[2929]), .A2(n[2928]), .A3(n[2931]), .A4(n[2930]), .Z(
        n1136) );
  XOR4D0 U1302 ( .A1(n[2936]), .A2(n[2935]), .A3(n[2938]), .A4(n[2937]), .Z(
        n1134) );
  XOR4D0 U1303 ( .A1(n[2943]), .A2(n[2942]), .A3(n[2945]), .A4(n[2944]), .Z(
        n1131) );
  XOR4D0 U1304 ( .A1(n[2950]), .A2(n[2949]), .A3(n[2952]), .A4(n[2951]), .Z(
        n1129) );
  XOR4D0 U1305 ( .A1(n[2957]), .A2(n[2956]), .A3(n[2959]), .A4(n[2958]), .Z(
        n1126) );
  XOR4D0 U1306 ( .A1(n[2964]), .A2(n[2963]), .A3(n[2966]), .A4(n[2965]), .Z(
        n1124) );
  XOR4D0 U1307 ( .A1(n[2971]), .A2(n[2970]), .A3(n[2973]), .A4(n[2972]), .Z(
        n1121) );
  XOR4D0 U1308 ( .A1(n[2978]), .A2(n[2977]), .A3(n[2980]), .A4(n[2979]), .Z(
        n1119) );
  XOR4D0 U1309 ( .A1(n[2985]), .A2(n[2984]), .A3(n[2987]), .A4(n[2986]), .Z(
        n1116) );
  XOR4D0 U1310 ( .A1(n[2992]), .A2(n[2991]), .A3(n[2994]), .A4(n[2993]), .Z(
        n1114) );
  XOR4D0 U1311 ( .A1(n[2999]), .A2(n[2998]), .A3(n[3001]), .A4(n[3000]), .Z(
        n1111) );
  XOR4D0 U1312 ( .A1(n[3006]), .A2(n[3005]), .A3(n[3008]), .A4(n[3007]), .Z(
        n1109) );
  XOR4D0 U1313 ( .A1(n[3013]), .A2(n[3012]), .A3(n[3015]), .A4(n[3014]), .Z(
        n1106) );
  XOR4D0 U1314 ( .A1(n[3020]), .A2(n[3019]), .A3(n[3022]), .A4(n[3021]), .Z(
        n1104) );
  XOR4D0 U1315 ( .A1(n[3027]), .A2(n[3026]), .A3(n[3029]), .A4(n[3028]), .Z(
        n1101) );
  XOR4D0 U1316 ( .A1(n[3034]), .A2(n[3033]), .A3(n[3036]), .A4(n[3035]), .Z(
        n1099) );
  XOR4D0 U1317 ( .A1(n[3041]), .A2(n[3040]), .A3(n[3043]), .A4(n[3042]), .Z(
        n1096) );
  XOR4D0 U1318 ( .A1(n[3048]), .A2(n[3047]), .A3(n[3050]), .A4(n[3049]), .Z(
        n1094) );
  XOR4D0 U1319 ( .A1(n[3055]), .A2(n[3054]), .A3(n[3057]), .A4(n[3056]), .Z(
        n1091) );
  XOR4D0 U1320 ( .A1(n[3062]), .A2(n[3061]), .A3(n[3064]), .A4(n[3063]), .Z(
        n1089) );
  XOR4D0 U1321 ( .A1(n[3069]), .A2(n[3068]), .A3(n[3071]), .A4(n[3070]), .Z(
        n1086) );
  XOR4D0 U1322 ( .A1(n[3076]), .A2(n[3075]), .A3(n[3078]), .A4(n[3077]), .Z(
        n1084) );
  XOR4D0 U1323 ( .A1(n[3083]), .A2(n[3082]), .A3(n[3085]), .A4(n[3084]), .Z(
        n1081) );
  XOR4D0 U1324 ( .A1(n[3090]), .A2(n[3089]), .A3(n[3092]), .A4(n[3091]), .Z(
        n1079) );
  XOR4D0 U1325 ( .A1(n[3097]), .A2(n[3096]), .A3(n[3099]), .A4(n[3098]), .Z(
        n1076) );
  XOR4D0 U1326 ( .A1(n[3104]), .A2(n[3103]), .A3(n[3106]), .A4(n[3105]), .Z(
        n1074) );
  XOR4D0 U1327 ( .A1(n[3111]), .A2(n[3110]), .A3(n[3113]), .A4(n[3112]), .Z(
        n1071) );
  XOR4D0 U1328 ( .A1(n[3118]), .A2(n[3117]), .A3(n[3120]), .A4(n[3119]), .Z(
        n1069) );
  XOR4D0 U1329 ( .A1(n[3125]), .A2(n[3124]), .A3(n[3127]), .A4(n[3126]), .Z(
        n1066) );
  XOR4D0 U1330 ( .A1(n[3132]), .A2(n[3131]), .A3(n[3134]), .A4(n[3133]), .Z(
        n1064) );
  XOR4D0 U1331 ( .A1(n[3139]), .A2(n[3138]), .A3(n[3141]), .A4(n[3140]), .Z(
        n1061) );
  XOR4D0 U1332 ( .A1(n[3146]), .A2(n[3145]), .A3(n[3148]), .A4(n[3147]), .Z(
        n1059) );
  XOR4D0 U1333 ( .A1(n[3153]), .A2(n[3152]), .A3(n[3155]), .A4(n[3154]), .Z(
        n1056) );
  XOR4D0 U1334 ( .A1(n[3160]), .A2(n[3159]), .A3(n[3162]), .A4(n[3161]), .Z(
        n1054) );
  XOR4D0 U1335 ( .A1(n[3167]), .A2(n[3166]), .A3(n[3169]), .A4(n[3168]), .Z(
        n1051) );
  XOR4D0 U1336 ( .A1(n[3174]), .A2(n[3173]), .A3(n[3176]), .A4(n[3175]), .Z(
        n1049) );
  XOR4D0 U1337 ( .A1(n[3181]), .A2(n[3180]), .A3(n[3183]), .A4(n[3182]), .Z(
        n1046) );
  XOR4D0 U1338 ( .A1(n[3188]), .A2(n[3187]), .A3(n[3190]), .A4(n[3189]), .Z(
        n1044) );
  XOR4D0 U1339 ( .A1(n[3195]), .A2(n[3194]), .A3(n[3197]), .A4(n[3196]), .Z(
        n1041) );
  XOR4D0 U1340 ( .A1(n[3202]), .A2(n[3201]), .A3(n[3204]), .A4(n[3203]), .Z(
        n1039) );
  XOR4D0 U1341 ( .A1(n[3209]), .A2(n[3208]), .A3(n[3211]), .A4(n[3210]), .Z(
        n1036) );
  XOR4D0 U1342 ( .A1(n[3216]), .A2(n[3215]), .A3(n[3218]), .A4(n[3217]), .Z(
        n1034) );
  XOR4D0 U1343 ( .A1(n[3223]), .A2(n[3222]), .A3(n[3225]), .A4(n[3224]), .Z(
        n1031) );
  XOR4D0 U1344 ( .A1(n[3230]), .A2(n[3229]), .A3(n[3232]), .A4(n[3231]), .Z(
        n1029) );
  XOR4D0 U1345 ( .A1(n[3237]), .A2(n[3236]), .A3(n[3239]), .A4(n[3238]), .Z(
        n1026) );
  XOR4D0 U1346 ( .A1(n[3244]), .A2(n[3243]), .A3(n[3246]), .A4(n[3245]), .Z(
        n1024) );
  XOR4D0 U1347 ( .A1(n[3251]), .A2(n[3250]), .A3(n[3253]), .A4(n[3252]), .Z(
        n1021) );
  XOR4D0 U1348 ( .A1(n[3258]), .A2(n[3257]), .A3(n[3260]), .A4(n[3259]), .Z(
        n1019) );
  XOR4D0 U1349 ( .A1(n[3265]), .A2(n[3264]), .A3(n[3267]), .A4(n[3266]), .Z(
        n1016) );
  XOR4D0 U1350 ( .A1(n[3272]), .A2(n[3271]), .A3(n[3274]), .A4(n[3273]), .Z(
        n1014) );
  XOR4D0 U1351 ( .A1(n[3279]), .A2(n[3278]), .A3(n[3281]), .A4(n[3280]), .Z(
        n1011) );
  XOR4D0 U1352 ( .A1(n[3286]), .A2(n[3285]), .A3(n[3288]), .A4(n[3287]), .Z(
        n1009) );
  XOR4D0 U1353 ( .A1(n[3293]), .A2(n[3292]), .A3(n[3295]), .A4(n[3294]), .Z(
        n1006) );
  XOR4D0 U1354 ( .A1(n[3300]), .A2(n[3299]), .A3(n[3302]), .A4(n[3301]), .Z(
        n1004) );
  XOR4D0 U1355 ( .A1(n[3307]), .A2(n[3306]), .A3(n[3309]), .A4(n[3308]), .Z(
        n1001) );
  XOR4D0 U1356 ( .A1(n[3314]), .A2(n[3313]), .A3(n[3316]), .A4(n[3315]), .Z(
        n999) );
  XOR4D0 U1357 ( .A1(n[3321]), .A2(n[3320]), .A3(n[3323]), .A4(n[3322]), .Z(
        n996) );
  XOR4D0 U1358 ( .A1(n[3328]), .A2(n[3327]), .A3(n[3330]), .A4(n[3329]), .Z(
        n994) );
  XOR4D0 U1359 ( .A1(n[3335]), .A2(n[3334]), .A3(n[3337]), .A4(n[3336]), .Z(
        n991) );
  XOR4D0 U1360 ( .A1(n[3342]), .A2(n[3341]), .A3(n[3344]), .A4(n[3343]), .Z(
        n989) );
  XOR4D0 U1361 ( .A1(n[3349]), .A2(n[3348]), .A3(n[3351]), .A4(n[3350]), .Z(
        n986) );
  XOR4D0 U1362 ( .A1(n[3356]), .A2(n[3355]), .A3(n[3358]), .A4(n[3357]), .Z(
        n984) );
  XOR4D0 U1363 ( .A1(n[3363]), .A2(n[3362]), .A3(n[3365]), .A4(n[3364]), .Z(
        n981) );
  XOR4D0 U1364 ( .A1(n[3370]), .A2(n[3369]), .A3(n[3372]), .A4(n[3371]), .Z(
        n979) );
  XOR4D0 U1365 ( .A1(n[3377]), .A2(n[3376]), .A3(n[3379]), .A4(n[3378]), .Z(
        n976) );
  XOR4D0 U1366 ( .A1(n[3384]), .A2(n[3383]), .A3(n[3386]), .A4(n[3385]), .Z(
        n974) );
  XOR4D0 U1367 ( .A1(n[3391]), .A2(n[3390]), .A3(n[3393]), .A4(n[3392]), .Z(
        n971) );
  XOR4D0 U1368 ( .A1(n[3398]), .A2(n[3397]), .A3(n[3400]), .A4(n[3399]), .Z(
        n969) );
  XOR4D0 U1369 ( .A1(n[3405]), .A2(n[3404]), .A3(n[3407]), .A4(n[3406]), .Z(
        n966) );
  XOR4D0 U1370 ( .A1(n[3412]), .A2(n[3411]), .A3(n[3414]), .A4(n[3413]), .Z(
        n964) );
  XOR4D0 U1371 ( .A1(n[3419]), .A2(n[3418]), .A3(n[3421]), .A4(n[3420]), .Z(
        n961) );
  XOR4D0 U1372 ( .A1(n[3426]), .A2(n[3425]), .A3(n[3428]), .A4(n[3427]), .Z(
        n959) );
  XOR4D0 U1373 ( .A1(n[3433]), .A2(n[3432]), .A3(n[3435]), .A4(n[3434]), .Z(
        n956) );
  XOR4D0 U1374 ( .A1(n[3440]), .A2(n[3439]), .A3(n[3442]), .A4(n[3441]), .Z(
        n954) );
  XOR4D0 U1375 ( .A1(n[3447]), .A2(n[3446]), .A3(n[3449]), .A4(n[3448]), .Z(
        n951) );
  XOR4D0 U1376 ( .A1(n[3454]), .A2(n[3453]), .A3(n[3456]), .A4(n[3455]), .Z(
        n949) );
  XOR4D0 U1377 ( .A1(n[3461]), .A2(n[3460]), .A3(n[3463]), .A4(n[3462]), .Z(
        n946) );
  XOR4D0 U1378 ( .A1(n[3468]), .A2(n[3467]), .A3(n[3470]), .A4(n[3469]), .Z(
        n944) );
  XOR4D0 U1379 ( .A1(n[3475]), .A2(n[3474]), .A3(n[3477]), .A4(n[3476]), .Z(
        n941) );
  XOR4D0 U1380 ( .A1(n[3482]), .A2(n[3481]), .A3(n[3484]), .A4(n[3483]), .Z(
        n939) );
  XOR4D0 U1381 ( .A1(n[3489]), .A2(n[3488]), .A3(n[3491]), .A4(n[3490]), .Z(
        n936) );
  XOR4D0 U1382 ( .A1(n[3496]), .A2(n[3495]), .A3(n[3498]), .A4(n[3497]), .Z(
        n934) );
  XOR4D0 U1383 ( .A1(n[3503]), .A2(n[3502]), .A3(n[3505]), .A4(n[3504]), .Z(
        n931) );
  XOR4D0 U1384 ( .A1(n[3510]), .A2(n[3509]), .A3(n[3512]), .A4(n[3511]), .Z(
        n929) );
  XOR4D0 U1385 ( .A1(n[3517]), .A2(n[3516]), .A3(n[3519]), .A4(n[3518]), .Z(
        n926) );
  XOR4D0 U1386 ( .A1(n[3524]), .A2(n[3523]), .A3(n[3526]), .A4(n[3525]), .Z(
        n924) );
  XOR4D0 U1387 ( .A1(n[3531]), .A2(n[3530]), .A3(n[3533]), .A4(n[3532]), .Z(
        n921) );
  XOR4D0 U1388 ( .A1(n[3538]), .A2(n[3537]), .A3(n[3540]), .A4(n[3539]), .Z(
        n919) );
  XOR4D0 U1389 ( .A1(n[3545]), .A2(n[3544]), .A3(n[3547]), .A4(n[3546]), .Z(
        n916) );
  XOR4D0 U1390 ( .A1(n[3552]), .A2(n[3551]), .A3(n[3554]), .A4(n[3553]), .Z(
        n914) );
  XOR4D0 U1391 ( .A1(n[3559]), .A2(n[3558]), .A3(n[3561]), .A4(n[3560]), .Z(
        n911) );
  XOR4D0 U1392 ( .A1(n[3566]), .A2(n[3565]), .A3(n[3568]), .A4(n[3567]), .Z(
        n909) );
  XOR4D0 U1393 ( .A1(n[3573]), .A2(n[3572]), .A3(n[3575]), .A4(n[3574]), .Z(
        n906) );
  XOR4D0 U1394 ( .A1(n[3580]), .A2(n[3579]), .A3(n[3582]), .A4(n[3581]), .Z(
        n904) );
  XOR4D0 U1395 ( .A1(n[3587]), .A2(n[3586]), .A3(n[3589]), .A4(n[3588]), .Z(
        n901) );
  XOR4D0 U1396 ( .A1(n[3594]), .A2(n[3593]), .A3(n[3596]), .A4(n[3595]), .Z(
        n899) );
  XOR4D0 U1397 ( .A1(n[3601]), .A2(n[3600]), .A3(n[3603]), .A4(n[3602]), .Z(
        n896) );
  XOR4D0 U1398 ( .A1(n[3608]), .A2(n[3607]), .A3(n[3610]), .A4(n[3609]), .Z(
        n894) );
  XOR4D0 U1399 ( .A1(n[3615]), .A2(n[3614]), .A3(n[3617]), .A4(n[3616]), .Z(
        n891) );
  XOR4D0 U1400 ( .A1(n[3622]), .A2(n[3621]), .A3(n[3624]), .A4(n[3623]), .Z(
        n889) );
  XOR4D0 U1401 ( .A1(n[3629]), .A2(n[3628]), .A3(n[3631]), .A4(n[3630]), .Z(
        n886) );
  XOR4D0 U1402 ( .A1(n[3636]), .A2(n[3635]), .A3(n[3638]), .A4(n[3637]), .Z(
        n884) );
  XOR4D0 U1403 ( .A1(n[3643]), .A2(n[3642]), .A3(n[3645]), .A4(n[3644]), .Z(
        n881) );
  XOR4D0 U1404 ( .A1(n[3650]), .A2(n[3649]), .A3(n[3652]), .A4(n[3651]), .Z(
        n879) );
  XOR4D0 U1405 ( .A1(n[3657]), .A2(n[3656]), .A3(n[3659]), .A4(n[3658]), .Z(
        n876) );
  XOR4D0 U1406 ( .A1(n[3664]), .A2(n[3663]), .A3(n[3666]), .A4(n[3665]), .Z(
        n874) );
  XOR4D0 U1407 ( .A1(n[3671]), .A2(n[3670]), .A3(n[3673]), .A4(n[3672]), .Z(
        n871) );
  XOR4D0 U1408 ( .A1(n[3678]), .A2(n[3677]), .A3(n[3680]), .A4(n[3679]), .Z(
        n869) );
  XOR4D0 U1409 ( .A1(n[3685]), .A2(n[3684]), .A3(n[3687]), .A4(n[3686]), .Z(
        n866) );
  XOR4D0 U1410 ( .A1(n[3692]), .A2(n[3691]), .A3(n[3694]), .A4(n[3693]), .Z(
        n864) );
  XOR4D0 U1411 ( .A1(n[3699]), .A2(n[3698]), .A3(n[3701]), .A4(n[3700]), .Z(
        n861) );
  XOR4D0 U1412 ( .A1(n[3706]), .A2(n[3705]), .A3(n[3708]), .A4(n[3707]), .Z(
        n859) );
  XOR4D0 U1413 ( .A1(n[3713]), .A2(n[3712]), .A3(n[3715]), .A4(n[3714]), .Z(
        n856) );
  XOR4D0 U1414 ( .A1(n[3720]), .A2(n[3719]), .A3(n[3722]), .A4(n[3721]), .Z(
        n854) );
  XOR4D0 U1415 ( .A1(n[3727]), .A2(n[3726]), .A3(n[3729]), .A4(n[3728]), .Z(
        n851) );
  XOR4D0 U1416 ( .A1(n[3734]), .A2(n[3733]), .A3(n[3736]), .A4(n[3735]), .Z(
        n849) );
  XOR4D0 U1417 ( .A1(n[3741]), .A2(n[3740]), .A3(n[3743]), .A4(n[3742]), .Z(
        n846) );
  XOR4D0 U1418 ( .A1(n[3748]), .A2(n[3747]), .A3(n[3750]), .A4(n[3749]), .Z(
        n844) );
  XOR4D0 U1419 ( .A1(n[3755]), .A2(n[3754]), .A3(n[3757]), .A4(n[3756]), .Z(
        n841) );
  XOR4D0 U1420 ( .A1(n[3762]), .A2(n[3761]), .A3(n[3764]), .A4(n[3763]), .Z(
        n839) );
  XOR4D0 U1421 ( .A1(n[3769]), .A2(n[3768]), .A3(n[3771]), .A4(n[3770]), .Z(
        n836) );
  XOR4D0 U1422 ( .A1(n[3776]), .A2(n[3775]), .A3(n[3778]), .A4(n[3777]), .Z(
        n834) );
  XOR4D0 U1423 ( .A1(n[3783]), .A2(n[3782]), .A3(n[3785]), .A4(n[3784]), .Z(
        n831) );
  XOR4D0 U1424 ( .A1(n[3790]), .A2(n[3789]), .A3(n[3792]), .A4(n[3791]), .Z(
        n829) );
  XOR4D0 U1425 ( .A1(n[3797]), .A2(n[3796]), .A3(n[3799]), .A4(n[3798]), .Z(
        n826) );
  XOR4D0 U1426 ( .A1(n[3804]), .A2(n[3803]), .A3(n[3806]), .A4(n[3805]), .Z(
        n824) );
  XOR4D0 U1427 ( .A1(n[3811]), .A2(n[3810]), .A3(n[3813]), .A4(n[3812]), .Z(
        n821) );
  XOR4D0 U1428 ( .A1(n[3818]), .A2(n[3817]), .A3(n[3820]), .A4(n[3819]), .Z(
        n819) );
  XOR4D0 U1429 ( .A1(n[3825]), .A2(n[3824]), .A3(n[3827]), .A4(n[3826]), .Z(
        n816) );
  XOR4D0 U1430 ( .A1(n[3832]), .A2(n[3831]), .A3(n[3834]), .A4(n[3833]), .Z(
        n814) );
  XOR4D0 U1431 ( .A1(n[3839]), .A2(n[3838]), .A3(n[3841]), .A4(n[3840]), .Z(
        n811) );
  XOR4D0 U1432 ( .A1(n[3846]), .A2(n[3845]), .A3(n[3848]), .A4(n[3847]), .Z(
        n809) );
  XOR4D0 U1433 ( .A1(n[3853]), .A2(n[3852]), .A3(n[3855]), .A4(n[3854]), .Z(
        n806) );
  XOR4D0 U1434 ( .A1(n[3860]), .A2(n[3859]), .A3(n[3862]), .A4(n[3861]), .Z(
        n804) );
  XOR4D0 U1435 ( .A1(n[3867]), .A2(n[3866]), .A3(n[3869]), .A4(n[3868]), .Z(
        n801) );
  XOR4D0 U1436 ( .A1(n[3874]), .A2(n[3873]), .A3(n[3876]), .A4(n[3875]), .Z(
        n799) );
  XOR4D0 U1437 ( .A1(n[3881]), .A2(n[3880]), .A3(n[3883]), .A4(n[3882]), .Z(
        n796) );
  XOR4D0 U1438 ( .A1(n[3888]), .A2(n[3887]), .A3(n[3890]), .A4(n[3889]), .Z(
        n794) );
  XOR4D0 U1439 ( .A1(n[3895]), .A2(n[3894]), .A3(n[3897]), .A4(n[3896]), .Z(
        n791) );
  XOR4D0 U1440 ( .A1(n[3902]), .A2(n[3901]), .A3(n[3904]), .A4(n[3903]), .Z(
        n789) );
  XOR4D0 U1441 ( .A1(n[3909]), .A2(n[3908]), .A3(n[3911]), .A4(n[3910]), .Z(
        n786) );
  XOR4D0 U1442 ( .A1(n[3916]), .A2(n[3915]), .A3(n[3918]), .A4(n[3917]), .Z(
        n784) );
  XOR4D0 U1443 ( .A1(n[3923]), .A2(n[3922]), .A3(n[3925]), .A4(n[3924]), .Z(
        n781) );
  XOR4D0 U1444 ( .A1(n[3930]), .A2(n[3929]), .A3(n[3932]), .A4(n[3931]), .Z(
        n779) );
  XOR4D0 U1445 ( .A1(n[3937]), .A2(n[3936]), .A3(n[3939]), .A4(n[3938]), .Z(
        n776) );
  XOR4D0 U1446 ( .A1(n[3944]), .A2(n[3943]), .A3(n[3946]), .A4(n[3945]), .Z(
        n774) );
  XOR4D0 U1447 ( .A1(n[3951]), .A2(n[3950]), .A3(n[3953]), .A4(n[3952]), .Z(
        n771) );
  XOR4D0 U1448 ( .A1(n[3958]), .A2(n[3957]), .A3(n[3960]), .A4(n[3959]), .Z(
        n769) );
  XOR4D0 U1449 ( .A1(n[3965]), .A2(n[3964]), .A3(n[3967]), .A4(n[3966]), .Z(
        n766) );
  XOR4D0 U1450 ( .A1(n[3972]), .A2(n[3971]), .A3(n[3974]), .A4(n[3973]), .Z(
        n764) );
  XOR4D0 U1451 ( .A1(n[3979]), .A2(n[3978]), .A3(n[3981]), .A4(n[3980]), .Z(
        n761) );
  XOR4D0 U1452 ( .A1(n[3986]), .A2(n[3985]), .A3(n[3988]), .A4(n[3987]), .Z(
        n759) );
  XOR4D0 U1453 ( .A1(n[3993]), .A2(n[3992]), .A3(n[3995]), .A4(n[3994]), .Z(
        n756) );
  XOR4D0 U1454 ( .A1(n[4000]), .A2(n[3999]), .A3(n[4002]), .A4(n[4001]), .Z(
        n754) );
  XOR4D0 U1455 ( .A1(n[4007]), .A2(n[4006]), .A3(n[4009]), .A4(n[4008]), .Z(
        n751) );
  XOR4D0 U1456 ( .A1(n[4014]), .A2(n[4013]), .A3(n[4016]), .A4(n[4015]), .Z(
        n749) );
  XOR4D0 U1457 ( .A1(n[4021]), .A2(n[4020]), .A3(n[4023]), .A4(n[4022]), .Z(
        n746) );
  XOR4D0 U1458 ( .A1(n[4028]), .A2(n[4027]), .A3(n[4030]), .A4(n[4029]), .Z(
        n744) );
  XOR4D0 U1459 ( .A1(n[4035]), .A2(n[4034]), .A3(n[4037]), .A4(n[4036]), .Z(
        n741) );
  XOR4D0 U1460 ( .A1(n[4042]), .A2(n[4041]), .A3(n[4044]), .A4(n[4043]), .Z(
        n739) );
  XOR4D0 U1461 ( .A1(n[4049]), .A2(n[4048]), .A3(n[4051]), .A4(n[4050]), .Z(
        n736) );
  XOR4D0 U1462 ( .A1(n[4056]), .A2(n[4055]), .A3(n[4058]), .A4(n[4057]), .Z(
        n734) );
  XOR4D0 U1463 ( .A1(n[4063]), .A2(n[4062]), .A3(n[4065]), .A4(n[4064]), .Z(
        n731) );
  XOR4D0 U1464 ( .A1(n[4070]), .A2(n[4069]), .A3(n[4072]), .A4(n[4071]), .Z(
        n729) );
  XOR4D0 U1465 ( .A1(n[4075]), .A2(n[4074]), .A3(n[4081]), .A4(n[4080]), .Z(
        n725) );
  XOR2D0 U1466 ( .A1(b[0]), .A2(a[0]), .Z(s[0]) );
endmodule


module gen_nonlinear_part ( a, b, n );
  input [10:0] a;
  input [10:0] b;
  output [4081:0] n;


  INVD0 U2 ( .I(1'b1), .ZN(n[1]) );
  INVD0 U4 ( .I(1'b1), .ZN(n[2]) );
  INVD0 U6 ( .I(1'b1), .ZN(n[5]) );
  INVD0 U8 ( .I(1'b1), .ZN(n[6]) );
  INVD0 U10 ( .I(1'b1), .ZN(n[8]) );
  INVD0 U12 ( .I(1'b1), .ZN(n[9]) );
  INVD0 U14 ( .I(1'b1), .ZN(n[13]) );
  INVD0 U16 ( .I(1'b1), .ZN(n[14]) );
  INVD0 U18 ( .I(1'b1), .ZN(n[16]) );
  INVD0 U20 ( .I(1'b1), .ZN(n[17]) );
  INVD0 U22 ( .I(1'b1), .ZN(n[20]) );
  INVD0 U24 ( .I(1'b1), .ZN(n[21]) );
  INVD0 U26 ( .I(1'b1), .ZN(n[23]) );
  INVD0 U28 ( .I(1'b1), .ZN(n[24]) );
  INVD0 U30 ( .I(1'b1), .ZN(n[29]) );
  INVD0 U32 ( .I(1'b1), .ZN(n[30]) );
  INVD0 U34 ( .I(1'b1), .ZN(n[32]) );
  INVD0 U36 ( .I(1'b1), .ZN(n[33]) );
  INVD0 U38 ( .I(1'b1), .ZN(n[36]) );
  INVD0 U40 ( .I(1'b1), .ZN(n[37]) );
  INVD0 U42 ( .I(1'b1), .ZN(n[39]) );
  INVD0 U44 ( .I(1'b1), .ZN(n[40]) );
  INVD0 U46 ( .I(1'b1), .ZN(n[44]) );
  INVD0 U48 ( .I(1'b1), .ZN(n[45]) );
  INVD0 U50 ( .I(1'b1), .ZN(n[47]) );
  INVD0 U52 ( .I(1'b1), .ZN(n[48]) );
  INVD0 U54 ( .I(1'b1), .ZN(n[51]) );
  INVD0 U56 ( .I(1'b1), .ZN(n[52]) );
  INVD0 U58 ( .I(1'b1), .ZN(n[54]) );
  INVD0 U60 ( .I(1'b1), .ZN(n[55]) );
  INVD0 U62 ( .I(1'b1), .ZN(n[61]) );
  INVD0 U64 ( .I(1'b1), .ZN(n[62]) );
  INVD0 U66 ( .I(1'b1), .ZN(n[64]) );
  INVD0 U68 ( .I(1'b1), .ZN(n[65]) );
  INVD0 U70 ( .I(1'b1), .ZN(n[68]) );
  INVD0 U72 ( .I(1'b1), .ZN(n[69]) );
  INVD0 U74 ( .I(1'b1), .ZN(n[71]) );
  INVD0 U76 ( .I(1'b1), .ZN(n[72]) );
  INVD0 U78 ( .I(1'b1), .ZN(n[76]) );
  INVD0 U80 ( .I(1'b1), .ZN(n[77]) );
  INVD0 U82 ( .I(1'b1), .ZN(n[79]) );
  INVD0 U84 ( .I(1'b1), .ZN(n[80]) );
  INVD0 U86 ( .I(1'b1), .ZN(n[83]) );
  INVD0 U88 ( .I(1'b1), .ZN(n[84]) );
  INVD0 U90 ( .I(1'b1), .ZN(n[86]) );
  INVD0 U92 ( .I(1'b1), .ZN(n[87]) );
  INVD0 U94 ( .I(1'b1), .ZN(n[92]) );
  INVD0 U96 ( .I(1'b1), .ZN(n[93]) );
  INVD0 U98 ( .I(1'b1), .ZN(n[95]) );
  INVD0 U100 ( .I(1'b1), .ZN(n[96]) );
  INVD0 U102 ( .I(1'b1), .ZN(n[99]) );
  INVD0 U104 ( .I(1'b1), .ZN(n[100]) );
  INVD0 U106 ( .I(1'b1), .ZN(n[102]) );
  INVD0 U108 ( .I(1'b1), .ZN(n[103]) );
  INVD0 U110 ( .I(1'b1), .ZN(n[107]) );
  INVD0 U112 ( .I(1'b1), .ZN(n[108]) );
  INVD0 U114 ( .I(1'b1), .ZN(n[110]) );
  INVD0 U116 ( .I(1'b1), .ZN(n[111]) );
  INVD0 U118 ( .I(1'b1), .ZN(n[114]) );
  INVD0 U120 ( .I(1'b1), .ZN(n[115]) );
  INVD0 U122 ( .I(1'b1), .ZN(n[117]) );
  INVD0 U124 ( .I(1'b1), .ZN(n[118]) );
  INVD0 U126 ( .I(1'b1), .ZN(n[125]) );
  INVD0 U128 ( .I(1'b1), .ZN(n[126]) );
  INVD0 U130 ( .I(1'b1), .ZN(n[128]) );
  INVD0 U132 ( .I(1'b1), .ZN(n[129]) );
  INVD0 U134 ( .I(1'b1), .ZN(n[132]) );
  INVD0 U136 ( .I(1'b1), .ZN(n[133]) );
  INVD0 U138 ( .I(1'b1), .ZN(n[135]) );
  INVD0 U140 ( .I(1'b1), .ZN(n[136]) );
  INVD0 U142 ( .I(1'b1), .ZN(n[140]) );
  INVD0 U144 ( .I(1'b1), .ZN(n[141]) );
  INVD0 U146 ( .I(1'b1), .ZN(n[143]) );
  INVD0 U148 ( .I(1'b1), .ZN(n[144]) );
  INVD0 U150 ( .I(1'b1), .ZN(n[147]) );
  INVD0 U152 ( .I(1'b1), .ZN(n[148]) );
  INVD0 U154 ( .I(1'b1), .ZN(n[150]) );
  INVD0 U156 ( .I(1'b1), .ZN(n[151]) );
  INVD0 U158 ( .I(1'b1), .ZN(n[156]) );
  INVD0 U160 ( .I(1'b1), .ZN(n[157]) );
  INVD0 U162 ( .I(1'b1), .ZN(n[159]) );
  INVD0 U164 ( .I(1'b1), .ZN(n[160]) );
  INVD0 U166 ( .I(1'b1), .ZN(n[163]) );
  INVD0 U168 ( .I(1'b1), .ZN(n[164]) );
  INVD0 U170 ( .I(1'b1), .ZN(n[166]) );
  INVD0 U172 ( .I(1'b1), .ZN(n[167]) );
  INVD0 U174 ( .I(1'b1), .ZN(n[171]) );
  INVD0 U176 ( .I(1'b1), .ZN(n[172]) );
  INVD0 U178 ( .I(1'b1), .ZN(n[174]) );
  INVD0 U180 ( .I(1'b1), .ZN(n[175]) );
  INVD0 U182 ( .I(1'b1), .ZN(n[178]) );
  INVD0 U184 ( .I(1'b1), .ZN(n[179]) );
  INVD0 U186 ( .I(1'b1), .ZN(n[181]) );
  INVD0 U188 ( .I(1'b1), .ZN(n[182]) );
  INVD0 U190 ( .I(1'b1), .ZN(n[188]) );
  INVD0 U192 ( .I(1'b1), .ZN(n[189]) );
  INVD0 U194 ( .I(1'b1), .ZN(n[191]) );
  INVD0 U196 ( .I(1'b1), .ZN(n[192]) );
  INVD0 U198 ( .I(1'b1), .ZN(n[195]) );
  INVD0 U200 ( .I(1'b1), .ZN(n[196]) );
  INVD0 U202 ( .I(1'b1), .ZN(n[198]) );
  INVD0 U204 ( .I(1'b1), .ZN(n[199]) );
  INVD0 U206 ( .I(1'b1), .ZN(n[203]) );
  INVD0 U208 ( .I(1'b1), .ZN(n[204]) );
  INVD0 U210 ( .I(1'b1), .ZN(n[206]) );
  INVD0 U212 ( .I(1'b1), .ZN(n[207]) );
  INVD0 U214 ( .I(1'b1), .ZN(n[210]) );
  INVD0 U216 ( .I(1'b1), .ZN(n[211]) );
  INVD0 U218 ( .I(1'b1), .ZN(n[213]) );
  INVD0 U220 ( .I(1'b1), .ZN(n[214]) );
  INVD0 U222 ( .I(1'b1), .ZN(n[219]) );
  INVD0 U224 ( .I(1'b1), .ZN(n[220]) );
  INVD0 U226 ( .I(1'b1), .ZN(n[222]) );
  INVD0 U228 ( .I(1'b1), .ZN(n[223]) );
  INVD0 U230 ( .I(1'b1), .ZN(n[226]) );
  INVD0 U232 ( .I(1'b1), .ZN(n[227]) );
  INVD0 U234 ( .I(1'b1), .ZN(n[229]) );
  INVD0 U236 ( .I(1'b1), .ZN(n[230]) );
  INVD0 U238 ( .I(1'b1), .ZN(n[234]) );
  INVD0 U240 ( .I(1'b1), .ZN(n[235]) );
  INVD0 U242 ( .I(1'b1), .ZN(n[237]) );
  INVD0 U244 ( .I(1'b1), .ZN(n[238]) );
  INVD0 U246 ( .I(1'b1), .ZN(n[241]) );
  INVD0 U248 ( .I(1'b1), .ZN(n[242]) );
  INVD0 U250 ( .I(1'b1), .ZN(n[244]) );
  INVD0 U252 ( .I(1'b1), .ZN(n[245]) );
  INVD0 U254 ( .I(1'b1), .ZN(n[253]) );
  INVD0 U256 ( .I(1'b1), .ZN(n[254]) );
  INVD0 U258 ( .I(1'b1), .ZN(n[256]) );
  INVD0 U260 ( .I(1'b1), .ZN(n[257]) );
  INVD0 U262 ( .I(1'b1), .ZN(n[260]) );
  INVD0 U264 ( .I(1'b1), .ZN(n[261]) );
  INVD0 U266 ( .I(1'b1), .ZN(n[263]) );
  INVD0 U268 ( .I(1'b1), .ZN(n[264]) );
  INVD0 U270 ( .I(1'b1), .ZN(n[268]) );
  INVD0 U272 ( .I(1'b1), .ZN(n[269]) );
  INVD0 U274 ( .I(1'b1), .ZN(n[271]) );
  INVD0 U276 ( .I(1'b1), .ZN(n[272]) );
  INVD0 U278 ( .I(1'b1), .ZN(n[275]) );
  INVD0 U280 ( .I(1'b1), .ZN(n[276]) );
  INVD0 U282 ( .I(1'b1), .ZN(n[278]) );
  INVD0 U284 ( .I(1'b1), .ZN(n[279]) );
  INVD0 U286 ( .I(1'b1), .ZN(n[284]) );
  INVD0 U288 ( .I(1'b1), .ZN(n[285]) );
  INVD0 U290 ( .I(1'b1), .ZN(n[287]) );
  INVD0 U292 ( .I(1'b1), .ZN(n[288]) );
  INVD0 U294 ( .I(1'b1), .ZN(n[291]) );
  INVD0 U296 ( .I(1'b1), .ZN(n[292]) );
  INVD0 U298 ( .I(1'b1), .ZN(n[294]) );
  INVD0 U300 ( .I(1'b1), .ZN(n[295]) );
  INVD0 U302 ( .I(1'b1), .ZN(n[299]) );
  INVD0 U304 ( .I(1'b1), .ZN(n[300]) );
  INVD0 U306 ( .I(1'b1), .ZN(n[302]) );
  INVD0 U308 ( .I(1'b1), .ZN(n[303]) );
  INVD0 U310 ( .I(1'b1), .ZN(n[306]) );
  INVD0 U312 ( .I(1'b1), .ZN(n[307]) );
  INVD0 U314 ( .I(1'b1), .ZN(n[309]) );
  INVD0 U316 ( .I(1'b1), .ZN(n[310]) );
  INVD0 U318 ( .I(1'b1), .ZN(n[316]) );
  INVD0 U320 ( .I(1'b1), .ZN(n[317]) );
  INVD0 U322 ( .I(1'b1), .ZN(n[319]) );
  INVD0 U324 ( .I(1'b1), .ZN(n[320]) );
  INVD0 U326 ( .I(1'b1), .ZN(n[323]) );
  INVD0 U328 ( .I(1'b1), .ZN(n[324]) );
  INVD0 U330 ( .I(1'b1), .ZN(n[326]) );
  INVD0 U332 ( .I(1'b1), .ZN(n[327]) );
  INVD0 U334 ( .I(1'b1), .ZN(n[331]) );
  INVD0 U336 ( .I(1'b1), .ZN(n[332]) );
  INVD0 U338 ( .I(1'b1), .ZN(n[334]) );
  INVD0 U340 ( .I(1'b1), .ZN(n[335]) );
  INVD0 U342 ( .I(1'b1), .ZN(n[338]) );
  INVD0 U344 ( .I(1'b1), .ZN(n[339]) );
  INVD0 U346 ( .I(1'b1), .ZN(n[341]) );
  INVD0 U348 ( .I(1'b1), .ZN(n[342]) );
  INVD0 U350 ( .I(1'b1), .ZN(n[347]) );
  INVD0 U352 ( .I(1'b1), .ZN(n[348]) );
  INVD0 U354 ( .I(1'b1), .ZN(n[350]) );
  INVD0 U356 ( .I(1'b1), .ZN(n[351]) );
  INVD0 U358 ( .I(1'b1), .ZN(n[354]) );
  INVD0 U360 ( .I(1'b1), .ZN(n[355]) );
  INVD0 U362 ( .I(1'b1), .ZN(n[357]) );
  INVD0 U364 ( .I(1'b1), .ZN(n[358]) );
  INVD0 U366 ( .I(1'b1), .ZN(n[362]) );
  INVD0 U368 ( .I(1'b1), .ZN(n[363]) );
  INVD0 U370 ( .I(1'b1), .ZN(n[365]) );
  INVD0 U372 ( .I(1'b1), .ZN(n[366]) );
  INVD0 U374 ( .I(1'b1), .ZN(n[369]) );
  INVD0 U376 ( .I(1'b1), .ZN(n[370]) );
  INVD0 U378 ( .I(1'b1), .ZN(n[372]) );
  INVD0 U380 ( .I(1'b1), .ZN(n[373]) );
  INVD0 U382 ( .I(1'b1), .ZN(n[380]) );
  INVD0 U384 ( .I(1'b1), .ZN(n[381]) );
  INVD0 U386 ( .I(1'b1), .ZN(n[383]) );
  INVD0 U388 ( .I(1'b1), .ZN(n[384]) );
  INVD0 U390 ( .I(1'b1), .ZN(n[387]) );
  INVD0 U392 ( .I(1'b1), .ZN(n[388]) );
  INVD0 U394 ( .I(1'b1), .ZN(n[390]) );
  INVD0 U396 ( .I(1'b1), .ZN(n[391]) );
  INVD0 U398 ( .I(1'b1), .ZN(n[395]) );
  INVD0 U400 ( .I(1'b1), .ZN(n[396]) );
  INVD0 U402 ( .I(1'b1), .ZN(n[398]) );
  INVD0 U404 ( .I(1'b1), .ZN(n[399]) );
  INVD0 U406 ( .I(1'b1), .ZN(n[402]) );
  INVD0 U408 ( .I(1'b1), .ZN(n[403]) );
  INVD0 U410 ( .I(1'b1), .ZN(n[405]) );
  INVD0 U412 ( .I(1'b1), .ZN(n[406]) );
  INVD0 U414 ( .I(1'b1), .ZN(n[411]) );
  INVD0 U416 ( .I(1'b1), .ZN(n[412]) );
  INVD0 U418 ( .I(1'b1), .ZN(n[414]) );
  INVD0 U420 ( .I(1'b1), .ZN(n[415]) );
  INVD0 U422 ( .I(1'b1), .ZN(n[418]) );
  INVD0 U424 ( .I(1'b1), .ZN(n[419]) );
  INVD0 U426 ( .I(1'b1), .ZN(n[421]) );
  INVD0 U428 ( .I(1'b1), .ZN(n[422]) );
  INVD0 U430 ( .I(1'b1), .ZN(n[426]) );
  INVD0 U432 ( .I(1'b1), .ZN(n[427]) );
  INVD0 U434 ( .I(1'b1), .ZN(n[429]) );
  INVD0 U436 ( .I(1'b1), .ZN(n[430]) );
  INVD0 U438 ( .I(1'b1), .ZN(n[433]) );
  INVD0 U440 ( .I(1'b1), .ZN(n[434]) );
  INVD0 U442 ( .I(1'b1), .ZN(n[436]) );
  INVD0 U444 ( .I(1'b1), .ZN(n[437]) );
  INVD0 U446 ( .I(1'b1), .ZN(n[443]) );
  INVD0 U448 ( .I(1'b1), .ZN(n[444]) );
  INVD0 U450 ( .I(1'b1), .ZN(n[446]) );
  INVD0 U452 ( .I(1'b1), .ZN(n[447]) );
  INVD0 U454 ( .I(1'b1), .ZN(n[450]) );
  INVD0 U456 ( .I(1'b1), .ZN(n[451]) );
  INVD0 U458 ( .I(1'b1), .ZN(n[453]) );
  INVD0 U460 ( .I(1'b1), .ZN(n[454]) );
  INVD0 U462 ( .I(1'b1), .ZN(n[458]) );
  INVD0 U464 ( .I(1'b1), .ZN(n[459]) );
  INVD0 U466 ( .I(1'b1), .ZN(n[461]) );
  INVD0 U468 ( .I(1'b1), .ZN(n[462]) );
  INVD0 U470 ( .I(1'b1), .ZN(n[465]) );
  INVD0 U472 ( .I(1'b1), .ZN(n[466]) );
  INVD0 U474 ( .I(1'b1), .ZN(n[468]) );
  INVD0 U476 ( .I(1'b1), .ZN(n[469]) );
  INVD0 U478 ( .I(1'b1), .ZN(n[474]) );
  INVD0 U480 ( .I(1'b1), .ZN(n[475]) );
  INVD0 U482 ( .I(1'b1), .ZN(n[477]) );
  INVD0 U484 ( .I(1'b1), .ZN(n[478]) );
  INVD0 U486 ( .I(1'b1), .ZN(n[481]) );
  INVD0 U488 ( .I(1'b1), .ZN(n[482]) );
  INVD0 U490 ( .I(1'b1), .ZN(n[484]) );
  INVD0 U492 ( .I(1'b1), .ZN(n[485]) );
  INVD0 U494 ( .I(1'b1), .ZN(n[489]) );
  INVD0 U496 ( .I(1'b1), .ZN(n[490]) );
  INVD0 U498 ( .I(1'b1), .ZN(n[492]) );
  INVD0 U500 ( .I(1'b1), .ZN(n[493]) );
  INVD0 U502 ( .I(1'b1), .ZN(n[496]) );
  INVD0 U504 ( .I(1'b1), .ZN(n[497]) );
  INVD0 U506 ( .I(1'b1), .ZN(n[499]) );
  INVD0 U508 ( .I(1'b1), .ZN(n[500]) );
  INVD0 U510 ( .I(1'b1), .ZN(n[509]) );
  INVD0 U512 ( .I(1'b1), .ZN(n[510]) );
  INVD0 U514 ( .I(1'b1), .ZN(n[512]) );
  INVD0 U516 ( .I(1'b1), .ZN(n[513]) );
  INVD0 U518 ( .I(1'b1), .ZN(n[516]) );
  INVD0 U520 ( .I(1'b1), .ZN(n[517]) );
  INVD0 U522 ( .I(1'b1), .ZN(n[519]) );
  INVD0 U524 ( .I(1'b1), .ZN(n[520]) );
  INVD0 U526 ( .I(1'b1), .ZN(n[524]) );
  INVD0 U528 ( .I(1'b1), .ZN(n[525]) );
  INVD0 U530 ( .I(1'b1), .ZN(n[527]) );
  INVD0 U532 ( .I(1'b1), .ZN(n[528]) );
  INVD0 U534 ( .I(1'b1), .ZN(n[531]) );
  INVD0 U536 ( .I(1'b1), .ZN(n[532]) );
  INVD0 U538 ( .I(1'b1), .ZN(n[534]) );
  INVD0 U540 ( .I(1'b1), .ZN(n[535]) );
  INVD0 U542 ( .I(1'b1), .ZN(n[540]) );
  INVD0 U544 ( .I(1'b1), .ZN(n[541]) );
  INVD0 U546 ( .I(1'b1), .ZN(n[543]) );
  INVD0 U548 ( .I(1'b1), .ZN(n[544]) );
  INVD0 U550 ( .I(1'b1), .ZN(n[547]) );
  INVD0 U552 ( .I(1'b1), .ZN(n[548]) );
  INVD0 U554 ( .I(1'b1), .ZN(n[550]) );
  INVD0 U556 ( .I(1'b1), .ZN(n[551]) );
  INVD0 U558 ( .I(1'b1), .ZN(n[555]) );
  INVD0 U560 ( .I(1'b1), .ZN(n[556]) );
  INVD0 U562 ( .I(1'b1), .ZN(n[558]) );
  INVD0 U564 ( .I(1'b1), .ZN(n[559]) );
  INVD0 U566 ( .I(1'b1), .ZN(n[562]) );
  INVD0 U568 ( .I(1'b1), .ZN(n[563]) );
  INVD0 U570 ( .I(1'b1), .ZN(n[565]) );
  INVD0 U572 ( .I(1'b1), .ZN(n[566]) );
  INVD0 U574 ( .I(1'b1), .ZN(n[572]) );
  INVD0 U576 ( .I(1'b1), .ZN(n[573]) );
  INVD0 U578 ( .I(1'b1), .ZN(n[575]) );
  INVD0 U580 ( .I(1'b1), .ZN(n[576]) );
  INVD0 U582 ( .I(1'b1), .ZN(n[579]) );
  INVD0 U584 ( .I(1'b1), .ZN(n[580]) );
  INVD0 U586 ( .I(1'b1), .ZN(n[582]) );
  INVD0 U588 ( .I(1'b1), .ZN(n[583]) );
  INVD0 U590 ( .I(1'b1), .ZN(n[587]) );
  INVD0 U592 ( .I(1'b1), .ZN(n[588]) );
  INVD0 U594 ( .I(1'b1), .ZN(n[590]) );
  INVD0 U596 ( .I(1'b1), .ZN(n[591]) );
  INVD0 U598 ( .I(1'b1), .ZN(n[594]) );
  INVD0 U600 ( .I(1'b1), .ZN(n[595]) );
  INVD0 U602 ( .I(1'b1), .ZN(n[597]) );
  INVD0 U604 ( .I(1'b1), .ZN(n[598]) );
  INVD0 U606 ( .I(1'b1), .ZN(n[603]) );
  INVD0 U608 ( .I(1'b1), .ZN(n[604]) );
  INVD0 U610 ( .I(1'b1), .ZN(n[606]) );
  INVD0 U612 ( .I(1'b1), .ZN(n[607]) );
  INVD0 U614 ( .I(1'b1), .ZN(n[610]) );
  INVD0 U616 ( .I(1'b1), .ZN(n[611]) );
  INVD0 U618 ( .I(1'b1), .ZN(n[613]) );
  INVD0 U620 ( .I(1'b1), .ZN(n[614]) );
  INVD0 U622 ( .I(1'b1), .ZN(n[618]) );
  INVD0 U624 ( .I(1'b1), .ZN(n[619]) );
  INVD0 U626 ( .I(1'b1), .ZN(n[621]) );
  INVD0 U628 ( .I(1'b1), .ZN(n[622]) );
  INVD0 U630 ( .I(1'b1), .ZN(n[625]) );
  INVD0 U632 ( .I(1'b1), .ZN(n[626]) );
  INVD0 U634 ( .I(1'b1), .ZN(n[628]) );
  INVD0 U636 ( .I(1'b1), .ZN(n[629]) );
  INVD0 U638 ( .I(1'b1), .ZN(n[636]) );
  INVD0 U640 ( .I(1'b1), .ZN(n[637]) );
  INVD0 U642 ( .I(1'b1), .ZN(n[639]) );
  INVD0 U644 ( .I(1'b1), .ZN(n[640]) );
  INVD0 U646 ( .I(1'b1), .ZN(n[643]) );
  INVD0 U648 ( .I(1'b1), .ZN(n[644]) );
  INVD0 U650 ( .I(1'b1), .ZN(n[646]) );
  INVD0 U652 ( .I(1'b1), .ZN(n[647]) );
  INVD0 U654 ( .I(1'b1), .ZN(n[651]) );
  INVD0 U656 ( .I(1'b1), .ZN(n[652]) );
  INVD0 U658 ( .I(1'b1), .ZN(n[654]) );
  INVD0 U660 ( .I(1'b1), .ZN(n[655]) );
  INVD0 U662 ( .I(1'b1), .ZN(n[658]) );
  INVD0 U664 ( .I(1'b1), .ZN(n[659]) );
  INVD0 U666 ( .I(1'b1), .ZN(n[661]) );
  INVD0 U668 ( .I(1'b1), .ZN(n[662]) );
  INVD0 U670 ( .I(1'b1), .ZN(n[667]) );
  INVD0 U672 ( .I(1'b1), .ZN(n[668]) );
  INVD0 U674 ( .I(1'b1), .ZN(n[670]) );
  INVD0 U676 ( .I(1'b1), .ZN(n[671]) );
  INVD0 U678 ( .I(1'b1), .ZN(n[674]) );
  INVD0 U680 ( .I(1'b1), .ZN(n[675]) );
  INVD0 U682 ( .I(1'b1), .ZN(n[677]) );
  INVD0 U684 ( .I(1'b1), .ZN(n[678]) );
  INVD0 U686 ( .I(1'b1), .ZN(n[682]) );
  INVD0 U688 ( .I(1'b1), .ZN(n[683]) );
  INVD0 U690 ( .I(1'b1), .ZN(n[685]) );
  INVD0 U692 ( .I(1'b1), .ZN(n[686]) );
  INVD0 U694 ( .I(1'b1), .ZN(n[689]) );
  INVD0 U696 ( .I(1'b1), .ZN(n[690]) );
  INVD0 U698 ( .I(1'b1), .ZN(n[692]) );
  INVD0 U700 ( .I(1'b1), .ZN(n[693]) );
  INVD0 U702 ( .I(1'b1), .ZN(n[699]) );
  INVD0 U704 ( .I(1'b1), .ZN(n[700]) );
  INVD0 U706 ( .I(1'b1), .ZN(n[702]) );
  INVD0 U708 ( .I(1'b1), .ZN(n[703]) );
  INVD0 U710 ( .I(1'b1), .ZN(n[706]) );
  INVD0 U712 ( .I(1'b1), .ZN(n[707]) );
  INVD0 U714 ( .I(1'b1), .ZN(n[709]) );
  INVD0 U716 ( .I(1'b1), .ZN(n[710]) );
  INVD0 U718 ( .I(1'b1), .ZN(n[714]) );
  INVD0 U720 ( .I(1'b1), .ZN(n[715]) );
  INVD0 U722 ( .I(1'b1), .ZN(n[717]) );
  INVD0 U724 ( .I(1'b1), .ZN(n[718]) );
  INVD0 U726 ( .I(1'b1), .ZN(n[721]) );
  INVD0 U728 ( .I(1'b1), .ZN(n[722]) );
  INVD0 U730 ( .I(1'b1), .ZN(n[724]) );
  INVD0 U732 ( .I(1'b1), .ZN(n[725]) );
  INVD0 U734 ( .I(1'b1), .ZN(n[730]) );
  INVD0 U736 ( .I(1'b1), .ZN(n[731]) );
  INVD0 U738 ( .I(1'b1), .ZN(n[733]) );
  INVD0 U740 ( .I(1'b1), .ZN(n[734]) );
  INVD0 U742 ( .I(1'b1), .ZN(n[737]) );
  INVD0 U744 ( .I(1'b1), .ZN(n[738]) );
  INVD0 U746 ( .I(1'b1), .ZN(n[740]) );
  INVD0 U748 ( .I(1'b1), .ZN(n[741]) );
  INVD0 U750 ( .I(1'b1), .ZN(n[745]) );
  INVD0 U752 ( .I(1'b1), .ZN(n[746]) );
  INVD0 U754 ( .I(1'b1), .ZN(n[748]) );
  INVD0 U756 ( .I(1'b1), .ZN(n[749]) );
  INVD0 U758 ( .I(1'b1), .ZN(n[752]) );
  INVD0 U760 ( .I(1'b1), .ZN(n[753]) );
  INVD0 U762 ( .I(1'b1), .ZN(n[755]) );
  INVD0 U764 ( .I(1'b1), .ZN(n[756]) );
  INVD0 U766 ( .I(1'b1), .ZN(n[764]) );
  INVD0 U768 ( .I(1'b1), .ZN(n[765]) );
  INVD0 U770 ( .I(1'b1), .ZN(n[767]) );
  INVD0 U772 ( .I(1'b1), .ZN(n[768]) );
  INVD0 U774 ( .I(1'b1), .ZN(n[771]) );
  INVD0 U776 ( .I(1'b1), .ZN(n[772]) );
  INVD0 U778 ( .I(1'b1), .ZN(n[774]) );
  INVD0 U780 ( .I(1'b1), .ZN(n[775]) );
  INVD0 U782 ( .I(1'b1), .ZN(n[779]) );
  INVD0 U784 ( .I(1'b1), .ZN(n[780]) );
  INVD0 U786 ( .I(1'b1), .ZN(n[782]) );
  INVD0 U788 ( .I(1'b1), .ZN(n[783]) );
  INVD0 U790 ( .I(1'b1), .ZN(n[786]) );
  INVD0 U792 ( .I(1'b1), .ZN(n[787]) );
  INVD0 U794 ( .I(1'b1), .ZN(n[789]) );
  INVD0 U796 ( .I(1'b1), .ZN(n[790]) );
  INVD0 U798 ( .I(1'b1), .ZN(n[795]) );
  INVD0 U800 ( .I(1'b1), .ZN(n[796]) );
  INVD0 U802 ( .I(1'b1), .ZN(n[798]) );
  INVD0 U804 ( .I(1'b1), .ZN(n[799]) );
  INVD0 U806 ( .I(1'b1), .ZN(n[802]) );
  INVD0 U808 ( .I(1'b1), .ZN(n[803]) );
  INVD0 U810 ( .I(1'b1), .ZN(n[805]) );
  INVD0 U812 ( .I(1'b1), .ZN(n[806]) );
  INVD0 U814 ( .I(1'b1), .ZN(n[810]) );
  INVD0 U816 ( .I(1'b1), .ZN(n[811]) );
  INVD0 U818 ( .I(1'b1), .ZN(n[813]) );
  INVD0 U820 ( .I(1'b1), .ZN(n[814]) );
  INVD0 U822 ( .I(1'b1), .ZN(n[817]) );
  INVD0 U824 ( .I(1'b1), .ZN(n[818]) );
  INVD0 U826 ( .I(1'b1), .ZN(n[820]) );
  INVD0 U828 ( .I(1'b1), .ZN(n[821]) );
  INVD0 U830 ( .I(1'b1), .ZN(n[827]) );
  INVD0 U832 ( .I(1'b1), .ZN(n[828]) );
  INVD0 U834 ( .I(1'b1), .ZN(n[830]) );
  INVD0 U836 ( .I(1'b1), .ZN(n[831]) );
  INVD0 U838 ( .I(1'b1), .ZN(n[834]) );
  INVD0 U840 ( .I(1'b1), .ZN(n[835]) );
  INVD0 U842 ( .I(1'b1), .ZN(n[837]) );
  INVD0 U844 ( .I(1'b1), .ZN(n[838]) );
  INVD0 U846 ( .I(1'b1), .ZN(n[842]) );
  INVD0 U848 ( .I(1'b1), .ZN(n[843]) );
  INVD0 U850 ( .I(1'b1), .ZN(n[845]) );
  INVD0 U852 ( .I(1'b1), .ZN(n[846]) );
  INVD0 U854 ( .I(1'b1), .ZN(n[849]) );
  INVD0 U856 ( .I(1'b1), .ZN(n[850]) );
  INVD0 U858 ( .I(1'b1), .ZN(n[852]) );
  INVD0 U860 ( .I(1'b1), .ZN(n[853]) );
  INVD0 U862 ( .I(1'b1), .ZN(n[858]) );
  INVD0 U864 ( .I(1'b1), .ZN(n[859]) );
  INVD0 U866 ( .I(1'b1), .ZN(n[861]) );
  INVD0 U868 ( .I(1'b1), .ZN(n[862]) );
  INVD0 U870 ( .I(1'b1), .ZN(n[865]) );
  INVD0 U872 ( .I(1'b1), .ZN(n[866]) );
  INVD0 U874 ( .I(1'b1), .ZN(n[868]) );
  INVD0 U876 ( .I(1'b1), .ZN(n[869]) );
  INVD0 U878 ( .I(1'b1), .ZN(n[873]) );
  INVD0 U880 ( .I(1'b1), .ZN(n[874]) );
  INVD0 U882 ( .I(1'b1), .ZN(n[876]) );
  INVD0 U884 ( .I(1'b1), .ZN(n[877]) );
  INVD0 U886 ( .I(1'b1), .ZN(n[880]) );
  INVD0 U888 ( .I(1'b1), .ZN(n[881]) );
  INVD0 U890 ( .I(1'b1), .ZN(n[883]) );
  INVD0 U892 ( .I(1'b1), .ZN(n[884]) );
  INVD0 U894 ( .I(1'b1), .ZN(n[891]) );
  INVD0 U896 ( .I(1'b1), .ZN(n[892]) );
  INVD0 U898 ( .I(1'b1), .ZN(n[894]) );
  INVD0 U900 ( .I(1'b1), .ZN(n[895]) );
  INVD0 U902 ( .I(1'b1), .ZN(n[898]) );
  INVD0 U904 ( .I(1'b1), .ZN(n[899]) );
  INVD0 U906 ( .I(1'b1), .ZN(n[901]) );
  INVD0 U908 ( .I(1'b1), .ZN(n[902]) );
  INVD0 U910 ( .I(1'b1), .ZN(n[906]) );
  INVD0 U912 ( .I(1'b1), .ZN(n[907]) );
  INVD0 U914 ( .I(1'b1), .ZN(n[909]) );
  INVD0 U916 ( .I(1'b1), .ZN(n[910]) );
  INVD0 U918 ( .I(1'b1), .ZN(n[913]) );
  INVD0 U920 ( .I(1'b1), .ZN(n[914]) );
  INVD0 U922 ( .I(1'b1), .ZN(n[916]) );
  INVD0 U924 ( .I(1'b1), .ZN(n[917]) );
  INVD0 U926 ( .I(1'b1), .ZN(n[922]) );
  INVD0 U928 ( .I(1'b1), .ZN(n[923]) );
  INVD0 U930 ( .I(1'b1), .ZN(n[925]) );
  INVD0 U932 ( .I(1'b1), .ZN(n[926]) );
  INVD0 U934 ( .I(1'b1), .ZN(n[929]) );
  INVD0 U936 ( .I(1'b1), .ZN(n[930]) );
  INVD0 U938 ( .I(1'b1), .ZN(n[932]) );
  INVD0 U940 ( .I(1'b1), .ZN(n[933]) );
  INVD0 U942 ( .I(1'b1), .ZN(n[937]) );
  INVD0 U944 ( .I(1'b1), .ZN(n[938]) );
  INVD0 U946 ( .I(1'b1), .ZN(n[940]) );
  INVD0 U948 ( .I(1'b1), .ZN(n[941]) );
  INVD0 U950 ( .I(1'b1), .ZN(n[944]) );
  INVD0 U952 ( .I(1'b1), .ZN(n[945]) );
  INVD0 U954 ( .I(1'b1), .ZN(n[947]) );
  INVD0 U956 ( .I(1'b1), .ZN(n[948]) );
  INVD0 U958 ( .I(1'b1), .ZN(n[954]) );
  INVD0 U960 ( .I(1'b1), .ZN(n[955]) );
  INVD0 U962 ( .I(1'b1), .ZN(n[957]) );
  INVD0 U964 ( .I(1'b1), .ZN(n[958]) );
  INVD0 U966 ( .I(1'b1), .ZN(n[961]) );
  INVD0 U968 ( .I(1'b1), .ZN(n[962]) );
  INVD0 U970 ( .I(1'b1), .ZN(n[964]) );
  INVD0 U972 ( .I(1'b1), .ZN(n[965]) );
  INVD0 U974 ( .I(1'b1), .ZN(n[969]) );
  INVD0 U976 ( .I(1'b1), .ZN(n[970]) );
  INVD0 U978 ( .I(1'b1), .ZN(n[972]) );
  INVD0 U980 ( .I(1'b1), .ZN(n[973]) );
  INVD0 U982 ( .I(1'b1), .ZN(n[976]) );
  INVD0 U984 ( .I(1'b1), .ZN(n[977]) );
  INVD0 U986 ( .I(1'b1), .ZN(n[979]) );
  INVD0 U988 ( .I(1'b1), .ZN(n[980]) );
  INVD0 U990 ( .I(1'b1), .ZN(n[985]) );
  INVD0 U992 ( .I(1'b1), .ZN(n[986]) );
  INVD0 U994 ( .I(1'b1), .ZN(n[988]) );
  INVD0 U996 ( .I(1'b1), .ZN(n[989]) );
  INVD0 U998 ( .I(1'b1), .ZN(n[992]) );
  INVD0 U1000 ( .I(1'b1), .ZN(n[993]) );
  INVD0 U1002 ( .I(1'b1), .ZN(n[995]) );
  INVD0 U1004 ( .I(1'b1), .ZN(n[996]) );
  INVD0 U1006 ( .I(1'b1), .ZN(n[1000]) );
  INVD0 U1008 ( .I(1'b1), .ZN(n[1001]) );
  INVD0 U1010 ( .I(1'b1), .ZN(n[1003]) );
  INVD0 U1012 ( .I(1'b1), .ZN(n[1004]) );
  INVD0 U1014 ( .I(1'b1), .ZN(n[1007]) );
  INVD0 U1016 ( .I(1'b1), .ZN(n[1008]) );
  INVD0 U1018 ( .I(1'b1), .ZN(n[1010]) );
  INVD0 U1020 ( .I(1'b1), .ZN(n[1011]) );
  INVD0 U1022 ( .I(1'b1), .ZN(n[1021]) );
  INVD0 U1024 ( .I(1'b1), .ZN(n[1022]) );
  INVD0 U1026 ( .I(1'b1), .ZN(n[1024]) );
  INVD0 U1028 ( .I(1'b1), .ZN(n[1025]) );
  INVD0 U1030 ( .I(1'b1), .ZN(n[1028]) );
  INVD0 U1032 ( .I(1'b1), .ZN(n[1029]) );
  INVD0 U1034 ( .I(1'b1), .ZN(n[1031]) );
  INVD0 U1036 ( .I(1'b1), .ZN(n[1032]) );
  INVD0 U1038 ( .I(1'b1), .ZN(n[1036]) );
  INVD0 U1040 ( .I(1'b1), .ZN(n[1037]) );
  INVD0 U1042 ( .I(1'b1), .ZN(n[1039]) );
  INVD0 U1044 ( .I(1'b1), .ZN(n[1040]) );
  INVD0 U1046 ( .I(1'b1), .ZN(n[1043]) );
  INVD0 U1048 ( .I(1'b1), .ZN(n[1044]) );
  INVD0 U1050 ( .I(1'b1), .ZN(n[1046]) );
  INVD0 U1052 ( .I(1'b1), .ZN(n[1047]) );
  INVD0 U1054 ( .I(1'b1), .ZN(n[1052]) );
  INVD0 U1056 ( .I(1'b1), .ZN(n[1053]) );
  INVD0 U1058 ( .I(1'b1), .ZN(n[1055]) );
  INVD0 U1060 ( .I(1'b1), .ZN(n[1056]) );
  INVD0 U1062 ( .I(1'b1), .ZN(n[1059]) );
  INVD0 U1064 ( .I(1'b1), .ZN(n[1060]) );
  INVD0 U1066 ( .I(1'b1), .ZN(n[1062]) );
  INVD0 U1068 ( .I(1'b1), .ZN(n[1063]) );
  INVD0 U1070 ( .I(1'b1), .ZN(n[1067]) );
  INVD0 U1072 ( .I(1'b1), .ZN(n[1068]) );
  INVD0 U1074 ( .I(1'b1), .ZN(n[1070]) );
  INVD0 U1076 ( .I(1'b1), .ZN(n[1071]) );
  INVD0 U1078 ( .I(1'b1), .ZN(n[1074]) );
  INVD0 U1080 ( .I(1'b1), .ZN(n[1075]) );
  INVD0 U1082 ( .I(1'b1), .ZN(n[1077]) );
  INVD0 U1084 ( .I(1'b1), .ZN(n[1078]) );
  INVD0 U1086 ( .I(1'b1), .ZN(n[1084]) );
  INVD0 U1088 ( .I(1'b1), .ZN(n[1085]) );
  INVD0 U1090 ( .I(1'b1), .ZN(n[1087]) );
  INVD0 U1092 ( .I(1'b1), .ZN(n[1088]) );
  INVD0 U1094 ( .I(1'b1), .ZN(n[1091]) );
  INVD0 U1096 ( .I(1'b1), .ZN(n[1092]) );
  INVD0 U1098 ( .I(1'b1), .ZN(n[1094]) );
  INVD0 U1100 ( .I(1'b1), .ZN(n[1095]) );
  INVD0 U1102 ( .I(1'b1), .ZN(n[1099]) );
  INVD0 U1104 ( .I(1'b1), .ZN(n[1100]) );
  INVD0 U1106 ( .I(1'b1), .ZN(n[1102]) );
  INVD0 U1108 ( .I(1'b1), .ZN(n[1103]) );
  INVD0 U1110 ( .I(1'b1), .ZN(n[1106]) );
  INVD0 U1112 ( .I(1'b1), .ZN(n[1107]) );
  INVD0 U1114 ( .I(1'b1), .ZN(n[1109]) );
  INVD0 U1116 ( .I(1'b1), .ZN(n[1110]) );
  INVD0 U1118 ( .I(1'b1), .ZN(n[1115]) );
  INVD0 U1120 ( .I(1'b1), .ZN(n[1116]) );
  INVD0 U1122 ( .I(1'b1), .ZN(n[1118]) );
  INVD0 U1124 ( .I(1'b1), .ZN(n[1119]) );
  INVD0 U1126 ( .I(1'b1), .ZN(n[1122]) );
  INVD0 U1128 ( .I(1'b1), .ZN(n[1123]) );
  INVD0 U1130 ( .I(1'b1), .ZN(n[1125]) );
  INVD0 U1132 ( .I(1'b1), .ZN(n[1126]) );
  INVD0 U1134 ( .I(1'b1), .ZN(n[1130]) );
  INVD0 U1136 ( .I(1'b1), .ZN(n[1131]) );
  INVD0 U1138 ( .I(1'b1), .ZN(n[1133]) );
  INVD0 U1140 ( .I(1'b1), .ZN(n[1134]) );
  INVD0 U1142 ( .I(1'b1), .ZN(n[1137]) );
  INVD0 U1144 ( .I(1'b1), .ZN(n[1138]) );
  INVD0 U1146 ( .I(1'b1), .ZN(n[1140]) );
  INVD0 U1148 ( .I(1'b1), .ZN(n[1141]) );
  INVD0 U1150 ( .I(1'b1), .ZN(n[1148]) );
  INVD0 U1152 ( .I(1'b1), .ZN(n[1149]) );
  INVD0 U1154 ( .I(1'b1), .ZN(n[1151]) );
  INVD0 U1156 ( .I(1'b1), .ZN(n[1152]) );
  INVD0 U1158 ( .I(1'b1), .ZN(n[1155]) );
  INVD0 U1160 ( .I(1'b1), .ZN(n[1156]) );
  INVD0 U1162 ( .I(1'b1), .ZN(n[1158]) );
  INVD0 U1164 ( .I(1'b1), .ZN(n[1159]) );
  INVD0 U1166 ( .I(1'b1), .ZN(n[1163]) );
  INVD0 U1168 ( .I(1'b1), .ZN(n[1164]) );
  INVD0 U1170 ( .I(1'b1), .ZN(n[1166]) );
  INVD0 U1172 ( .I(1'b1), .ZN(n[1167]) );
  INVD0 U1174 ( .I(1'b1), .ZN(n[1170]) );
  INVD0 U1176 ( .I(1'b1), .ZN(n[1171]) );
  INVD0 U1178 ( .I(1'b1), .ZN(n[1173]) );
  INVD0 U1180 ( .I(1'b1), .ZN(n[1174]) );
  INVD0 U1182 ( .I(1'b1), .ZN(n[1179]) );
  INVD0 U1184 ( .I(1'b1), .ZN(n[1180]) );
  INVD0 U1186 ( .I(1'b1), .ZN(n[1182]) );
  INVD0 U1188 ( .I(1'b1), .ZN(n[1183]) );
  INVD0 U1190 ( .I(1'b1), .ZN(n[1186]) );
  INVD0 U1192 ( .I(1'b1), .ZN(n[1187]) );
  INVD0 U1194 ( .I(1'b1), .ZN(n[1189]) );
  INVD0 U1196 ( .I(1'b1), .ZN(n[1190]) );
  INVD0 U1198 ( .I(1'b1), .ZN(n[1194]) );
  INVD0 U1200 ( .I(1'b1), .ZN(n[1195]) );
  INVD0 U1202 ( .I(1'b1), .ZN(n[1197]) );
  INVD0 U1204 ( .I(1'b1), .ZN(n[1198]) );
  INVD0 U1206 ( .I(1'b1), .ZN(n[1201]) );
  INVD0 U1208 ( .I(1'b1), .ZN(n[1202]) );
  INVD0 U1210 ( .I(1'b1), .ZN(n[1204]) );
  INVD0 U1212 ( .I(1'b1), .ZN(n[1205]) );
  INVD0 U1214 ( .I(1'b1), .ZN(n[1211]) );
  INVD0 U1216 ( .I(1'b1), .ZN(n[1212]) );
  INVD0 U1218 ( .I(1'b1), .ZN(n[1214]) );
  INVD0 U1220 ( .I(1'b1), .ZN(n[1215]) );
  INVD0 U1222 ( .I(1'b1), .ZN(n[1218]) );
  INVD0 U1224 ( .I(1'b1), .ZN(n[1219]) );
  INVD0 U1226 ( .I(1'b1), .ZN(n[1221]) );
  INVD0 U1228 ( .I(1'b1), .ZN(n[1222]) );
  INVD0 U1230 ( .I(1'b1), .ZN(n[1226]) );
  INVD0 U1232 ( .I(1'b1), .ZN(n[1227]) );
  INVD0 U1234 ( .I(1'b1), .ZN(n[1229]) );
  INVD0 U1236 ( .I(1'b1), .ZN(n[1230]) );
  INVD0 U1238 ( .I(1'b1), .ZN(n[1233]) );
  INVD0 U1240 ( .I(1'b1), .ZN(n[1234]) );
  INVD0 U1242 ( .I(1'b1), .ZN(n[1236]) );
  INVD0 U1244 ( .I(1'b1), .ZN(n[1237]) );
  INVD0 U1246 ( .I(1'b1), .ZN(n[1242]) );
  INVD0 U1248 ( .I(1'b1), .ZN(n[1243]) );
  INVD0 U1250 ( .I(1'b1), .ZN(n[1245]) );
  INVD0 U1252 ( .I(1'b1), .ZN(n[1246]) );
  INVD0 U1254 ( .I(1'b1), .ZN(n[1249]) );
  INVD0 U1256 ( .I(1'b1), .ZN(n[1250]) );
  INVD0 U1258 ( .I(1'b1), .ZN(n[1252]) );
  INVD0 U1260 ( .I(1'b1), .ZN(n[1253]) );
  INVD0 U1262 ( .I(1'b1), .ZN(n[1257]) );
  INVD0 U1264 ( .I(1'b1), .ZN(n[1258]) );
  INVD0 U1266 ( .I(1'b1), .ZN(n[1260]) );
  INVD0 U1268 ( .I(1'b1), .ZN(n[1261]) );
  INVD0 U1270 ( .I(1'b1), .ZN(n[1264]) );
  INVD0 U1272 ( .I(1'b1), .ZN(n[1265]) );
  INVD0 U1274 ( .I(1'b1), .ZN(n[1267]) );
  INVD0 U1276 ( .I(1'b1), .ZN(n[1268]) );
  INVD0 U1278 ( .I(1'b1), .ZN(n[1276]) );
  INVD0 U1280 ( .I(1'b1), .ZN(n[1277]) );
  INVD0 U1282 ( .I(1'b1), .ZN(n[1279]) );
  INVD0 U1284 ( .I(1'b1), .ZN(n[1280]) );
  INVD0 U1286 ( .I(1'b1), .ZN(n[1283]) );
  INVD0 U1288 ( .I(1'b1), .ZN(n[1284]) );
  INVD0 U1290 ( .I(1'b1), .ZN(n[1286]) );
  INVD0 U1292 ( .I(1'b1), .ZN(n[1287]) );
  INVD0 U1294 ( .I(1'b1), .ZN(n[1291]) );
  INVD0 U1296 ( .I(1'b1), .ZN(n[1292]) );
  INVD0 U1298 ( .I(1'b1), .ZN(n[1294]) );
  INVD0 U1300 ( .I(1'b1), .ZN(n[1295]) );
  INVD0 U1302 ( .I(1'b1), .ZN(n[1298]) );
  INVD0 U1304 ( .I(1'b1), .ZN(n[1299]) );
  INVD0 U1306 ( .I(1'b1), .ZN(n[1301]) );
  INVD0 U1308 ( .I(1'b1), .ZN(n[1302]) );
  INVD0 U1310 ( .I(1'b1), .ZN(n[1307]) );
  INVD0 U1312 ( .I(1'b1), .ZN(n[1308]) );
  INVD0 U1314 ( .I(1'b1), .ZN(n[1310]) );
  INVD0 U1316 ( .I(1'b1), .ZN(n[1311]) );
  INVD0 U1318 ( .I(1'b1), .ZN(n[1314]) );
  INVD0 U1320 ( .I(1'b1), .ZN(n[1315]) );
  INVD0 U1322 ( .I(1'b1), .ZN(n[1317]) );
  INVD0 U1324 ( .I(1'b1), .ZN(n[1318]) );
  INVD0 U1326 ( .I(1'b1), .ZN(n[1322]) );
  INVD0 U1328 ( .I(1'b1), .ZN(n[1323]) );
  INVD0 U1330 ( .I(1'b1), .ZN(n[1325]) );
  INVD0 U1332 ( .I(1'b1), .ZN(n[1326]) );
  INVD0 U1334 ( .I(1'b1), .ZN(n[1329]) );
  INVD0 U1336 ( .I(1'b1), .ZN(n[1330]) );
  INVD0 U1338 ( .I(1'b1), .ZN(n[1332]) );
  INVD0 U1340 ( .I(1'b1), .ZN(n[1333]) );
  INVD0 U1342 ( .I(1'b1), .ZN(n[1339]) );
  INVD0 U1344 ( .I(1'b1), .ZN(n[1340]) );
  INVD0 U1346 ( .I(1'b1), .ZN(n[1342]) );
  INVD0 U1348 ( .I(1'b1), .ZN(n[1343]) );
  INVD0 U1350 ( .I(1'b1), .ZN(n[1346]) );
  INVD0 U1352 ( .I(1'b1), .ZN(n[1347]) );
  INVD0 U1354 ( .I(1'b1), .ZN(n[1349]) );
  INVD0 U1356 ( .I(1'b1), .ZN(n[1350]) );
  INVD0 U1358 ( .I(1'b1), .ZN(n[1354]) );
  INVD0 U1360 ( .I(1'b1), .ZN(n[1355]) );
  INVD0 U1362 ( .I(1'b1), .ZN(n[1357]) );
  INVD0 U1364 ( .I(1'b1), .ZN(n[1358]) );
  INVD0 U1366 ( .I(1'b1), .ZN(n[1361]) );
  INVD0 U1368 ( .I(1'b1), .ZN(n[1362]) );
  INVD0 U1370 ( .I(1'b1), .ZN(n[1364]) );
  INVD0 U1372 ( .I(1'b1), .ZN(n[1365]) );
  INVD0 U1374 ( .I(1'b1), .ZN(n[1370]) );
  INVD0 U1376 ( .I(1'b1), .ZN(n[1371]) );
  INVD0 U1378 ( .I(1'b1), .ZN(n[1373]) );
  INVD0 U1380 ( .I(1'b1), .ZN(n[1374]) );
  INVD0 U1382 ( .I(1'b1), .ZN(n[1377]) );
  INVD0 U1384 ( .I(1'b1), .ZN(n[1378]) );
  INVD0 U1386 ( .I(1'b1), .ZN(n[1380]) );
  INVD0 U1388 ( .I(1'b1), .ZN(n[1381]) );
  INVD0 U1390 ( .I(1'b1), .ZN(n[1385]) );
  INVD0 U1392 ( .I(1'b1), .ZN(n[1386]) );
  INVD0 U1394 ( .I(1'b1), .ZN(n[1388]) );
  INVD0 U1396 ( .I(1'b1), .ZN(n[1389]) );
  INVD0 U1398 ( .I(1'b1), .ZN(n[1392]) );
  INVD0 U1400 ( .I(1'b1), .ZN(n[1393]) );
  INVD0 U1402 ( .I(1'b1), .ZN(n[1395]) );
  INVD0 U1404 ( .I(1'b1), .ZN(n[1396]) );
  INVD0 U1406 ( .I(1'b1), .ZN(n[1403]) );
  INVD0 U1408 ( .I(1'b1), .ZN(n[1404]) );
  INVD0 U1410 ( .I(1'b1), .ZN(n[1406]) );
  INVD0 U1412 ( .I(1'b1), .ZN(n[1407]) );
  INVD0 U1414 ( .I(1'b1), .ZN(n[1410]) );
  INVD0 U1416 ( .I(1'b1), .ZN(n[1411]) );
  INVD0 U1418 ( .I(1'b1), .ZN(n[1413]) );
  INVD0 U1420 ( .I(1'b1), .ZN(n[1414]) );
  INVD0 U1422 ( .I(1'b1), .ZN(n[1418]) );
  INVD0 U1424 ( .I(1'b1), .ZN(n[1419]) );
  INVD0 U1426 ( .I(1'b1), .ZN(n[1421]) );
  INVD0 U1428 ( .I(1'b1), .ZN(n[1422]) );
  INVD0 U1430 ( .I(1'b1), .ZN(n[1425]) );
  INVD0 U1432 ( .I(1'b1), .ZN(n[1426]) );
  INVD0 U1434 ( .I(1'b1), .ZN(n[1428]) );
  INVD0 U1436 ( .I(1'b1), .ZN(n[1429]) );
  INVD0 U1438 ( .I(1'b1), .ZN(n[1434]) );
  INVD0 U1440 ( .I(1'b1), .ZN(n[1435]) );
  INVD0 U1442 ( .I(1'b1), .ZN(n[1437]) );
  INVD0 U1444 ( .I(1'b1), .ZN(n[1438]) );
  INVD0 U1446 ( .I(1'b1), .ZN(n[1441]) );
  INVD0 U1448 ( .I(1'b1), .ZN(n[1442]) );
  INVD0 U1450 ( .I(1'b1), .ZN(n[1444]) );
  INVD0 U1452 ( .I(1'b1), .ZN(n[1445]) );
  INVD0 U1454 ( .I(1'b1), .ZN(n[1449]) );
  INVD0 U1456 ( .I(1'b1), .ZN(n[1450]) );
  INVD0 U1458 ( .I(1'b1), .ZN(n[1452]) );
  INVD0 U1460 ( .I(1'b1), .ZN(n[1453]) );
  INVD0 U1462 ( .I(1'b1), .ZN(n[1456]) );
  INVD0 U1464 ( .I(1'b1), .ZN(n[1457]) );
  INVD0 U1466 ( .I(1'b1), .ZN(n[1459]) );
  INVD0 U1468 ( .I(1'b1), .ZN(n[1460]) );
  INVD0 U1470 ( .I(1'b1), .ZN(n[1466]) );
  INVD0 U1472 ( .I(1'b1), .ZN(n[1467]) );
  INVD0 U1474 ( .I(1'b1), .ZN(n[1469]) );
  INVD0 U1476 ( .I(1'b1), .ZN(n[1470]) );
  INVD0 U1478 ( .I(1'b1), .ZN(n[1473]) );
  INVD0 U1480 ( .I(1'b1), .ZN(n[1474]) );
  INVD0 U1482 ( .I(1'b1), .ZN(n[1476]) );
  INVD0 U1484 ( .I(1'b1), .ZN(n[1477]) );
  INVD0 U1486 ( .I(1'b1), .ZN(n[1481]) );
  INVD0 U1488 ( .I(1'b1), .ZN(n[1482]) );
  INVD0 U1490 ( .I(1'b1), .ZN(n[1484]) );
  INVD0 U1492 ( .I(1'b1), .ZN(n[1485]) );
  INVD0 U1494 ( .I(1'b1), .ZN(n[1488]) );
  INVD0 U1496 ( .I(1'b1), .ZN(n[1489]) );
  INVD0 U1498 ( .I(1'b1), .ZN(n[1491]) );
  INVD0 U1500 ( .I(1'b1), .ZN(n[1492]) );
  INVD0 U1502 ( .I(1'b1), .ZN(n[1497]) );
  INVD0 U1504 ( .I(1'b1), .ZN(n[1498]) );
  INVD0 U1506 ( .I(1'b1), .ZN(n[1500]) );
  INVD0 U1508 ( .I(1'b1), .ZN(n[1501]) );
  INVD0 U1510 ( .I(1'b1), .ZN(n[1504]) );
  INVD0 U1512 ( .I(1'b1), .ZN(n[1505]) );
  INVD0 U1514 ( .I(1'b1), .ZN(n[1507]) );
  INVD0 U1516 ( .I(1'b1), .ZN(n[1508]) );
  INVD0 U1518 ( .I(1'b1), .ZN(n[1512]) );
  INVD0 U1520 ( .I(1'b1), .ZN(n[1513]) );
  INVD0 U1522 ( .I(1'b1), .ZN(n[1515]) );
  INVD0 U1524 ( .I(1'b1), .ZN(n[1516]) );
  INVD0 U1526 ( .I(1'b1), .ZN(n[1519]) );
  INVD0 U1528 ( .I(1'b1), .ZN(n[1520]) );
  INVD0 U1530 ( .I(1'b1), .ZN(n[1522]) );
  INVD0 U1532 ( .I(1'b1), .ZN(n[1523]) );
  INVD0 U1534 ( .I(1'b1), .ZN(n[1532]) );
  INVD0 U1536 ( .I(1'b1), .ZN(n[1533]) );
  INVD0 U1538 ( .I(1'b1), .ZN(n[1535]) );
  INVD0 U1540 ( .I(1'b1), .ZN(n[1536]) );
  INVD0 U1542 ( .I(1'b1), .ZN(n[1539]) );
  INVD0 U1544 ( .I(1'b1), .ZN(n[1540]) );
  INVD0 U1546 ( .I(1'b1), .ZN(n[1542]) );
  INVD0 U1548 ( .I(1'b1), .ZN(n[1543]) );
  INVD0 U1550 ( .I(1'b1), .ZN(n[1547]) );
  INVD0 U1552 ( .I(1'b1), .ZN(n[1548]) );
  INVD0 U1554 ( .I(1'b1), .ZN(n[1550]) );
  INVD0 U1556 ( .I(1'b1), .ZN(n[1551]) );
  INVD0 U1558 ( .I(1'b1), .ZN(n[1554]) );
  INVD0 U1560 ( .I(1'b1), .ZN(n[1555]) );
  INVD0 U1562 ( .I(1'b1), .ZN(n[1557]) );
  INVD0 U1564 ( .I(1'b1), .ZN(n[1558]) );
  INVD0 U1566 ( .I(1'b1), .ZN(n[1563]) );
  INVD0 U1568 ( .I(1'b1), .ZN(n[1564]) );
  INVD0 U1570 ( .I(1'b1), .ZN(n[1566]) );
  INVD0 U1572 ( .I(1'b1), .ZN(n[1567]) );
  INVD0 U1574 ( .I(1'b1), .ZN(n[1570]) );
  INVD0 U1576 ( .I(1'b1), .ZN(n[1571]) );
  INVD0 U1578 ( .I(1'b1), .ZN(n[1573]) );
  INVD0 U1580 ( .I(1'b1), .ZN(n[1574]) );
  INVD0 U1582 ( .I(1'b1), .ZN(n[1578]) );
  INVD0 U1584 ( .I(1'b1), .ZN(n[1579]) );
  INVD0 U1586 ( .I(1'b1), .ZN(n[1581]) );
  INVD0 U1588 ( .I(1'b1), .ZN(n[1582]) );
  INVD0 U1590 ( .I(1'b1), .ZN(n[1585]) );
  INVD0 U1592 ( .I(1'b1), .ZN(n[1586]) );
  INVD0 U1594 ( .I(1'b1), .ZN(n[1588]) );
  INVD0 U1596 ( .I(1'b1), .ZN(n[1589]) );
  INVD0 U1598 ( .I(1'b1), .ZN(n[1595]) );
  INVD0 U1600 ( .I(1'b1), .ZN(n[1596]) );
  INVD0 U1602 ( .I(1'b1), .ZN(n[1598]) );
  INVD0 U1604 ( .I(1'b1), .ZN(n[1599]) );
  INVD0 U1606 ( .I(1'b1), .ZN(n[1602]) );
  INVD0 U1608 ( .I(1'b1), .ZN(n[1603]) );
  INVD0 U1610 ( .I(1'b1), .ZN(n[1605]) );
  INVD0 U1612 ( .I(1'b1), .ZN(n[1606]) );
  INVD0 U1614 ( .I(1'b1), .ZN(n[1610]) );
  INVD0 U1616 ( .I(1'b1), .ZN(n[1611]) );
  INVD0 U1618 ( .I(1'b1), .ZN(n[1613]) );
  INVD0 U1620 ( .I(1'b1), .ZN(n[1614]) );
  INVD0 U1622 ( .I(1'b1), .ZN(n[1617]) );
  INVD0 U1624 ( .I(1'b1), .ZN(n[1618]) );
  INVD0 U1626 ( .I(1'b1), .ZN(n[1620]) );
  INVD0 U1628 ( .I(1'b1), .ZN(n[1621]) );
  INVD0 U1630 ( .I(1'b1), .ZN(n[1626]) );
  INVD0 U1632 ( .I(1'b1), .ZN(n[1627]) );
  INVD0 U1634 ( .I(1'b1), .ZN(n[1629]) );
  INVD0 U1636 ( .I(1'b1), .ZN(n[1630]) );
  INVD0 U1638 ( .I(1'b1), .ZN(n[1633]) );
  INVD0 U1640 ( .I(1'b1), .ZN(n[1634]) );
  INVD0 U1642 ( .I(1'b1), .ZN(n[1636]) );
  INVD0 U1644 ( .I(1'b1), .ZN(n[1637]) );
  INVD0 U1646 ( .I(1'b1), .ZN(n[1641]) );
  INVD0 U1648 ( .I(1'b1), .ZN(n[1642]) );
  INVD0 U1650 ( .I(1'b1), .ZN(n[1644]) );
  INVD0 U1652 ( .I(1'b1), .ZN(n[1645]) );
  INVD0 U1654 ( .I(1'b1), .ZN(n[1648]) );
  INVD0 U1656 ( .I(1'b1), .ZN(n[1649]) );
  INVD0 U1658 ( .I(1'b1), .ZN(n[1651]) );
  INVD0 U1660 ( .I(1'b1), .ZN(n[1652]) );
  INVD0 U1662 ( .I(1'b1), .ZN(n[1659]) );
  INVD0 U1664 ( .I(1'b1), .ZN(n[1660]) );
  INVD0 U1666 ( .I(1'b1), .ZN(n[1662]) );
  INVD0 U1668 ( .I(1'b1), .ZN(n[1663]) );
  INVD0 U1670 ( .I(1'b1), .ZN(n[1666]) );
  INVD0 U1672 ( .I(1'b1), .ZN(n[1667]) );
  INVD0 U1674 ( .I(1'b1), .ZN(n[1669]) );
  INVD0 U1676 ( .I(1'b1), .ZN(n[1670]) );
  INVD0 U1678 ( .I(1'b1), .ZN(n[1674]) );
  INVD0 U1680 ( .I(1'b1), .ZN(n[1675]) );
  INVD0 U1682 ( .I(1'b1), .ZN(n[1677]) );
  INVD0 U1684 ( .I(1'b1), .ZN(n[1678]) );
  INVD0 U1686 ( .I(1'b1), .ZN(n[1681]) );
  INVD0 U1688 ( .I(1'b1), .ZN(n[1682]) );
  INVD0 U1690 ( .I(1'b1), .ZN(n[1684]) );
  INVD0 U1692 ( .I(1'b1), .ZN(n[1685]) );
  INVD0 U1694 ( .I(1'b1), .ZN(n[1690]) );
  INVD0 U1696 ( .I(1'b1), .ZN(n[1691]) );
  INVD0 U1698 ( .I(1'b1), .ZN(n[1693]) );
  INVD0 U1700 ( .I(1'b1), .ZN(n[1694]) );
  INVD0 U1702 ( .I(1'b1), .ZN(n[1697]) );
  INVD0 U1704 ( .I(1'b1), .ZN(n[1698]) );
  INVD0 U1706 ( .I(1'b1), .ZN(n[1700]) );
  INVD0 U1708 ( .I(1'b1), .ZN(n[1701]) );
  INVD0 U1710 ( .I(1'b1), .ZN(n[1705]) );
  INVD0 U1712 ( .I(1'b1), .ZN(n[1706]) );
  INVD0 U1714 ( .I(1'b1), .ZN(n[1708]) );
  INVD0 U1716 ( .I(1'b1), .ZN(n[1709]) );
  INVD0 U1718 ( .I(1'b1), .ZN(n[1712]) );
  INVD0 U1720 ( .I(1'b1), .ZN(n[1713]) );
  INVD0 U1722 ( .I(1'b1), .ZN(n[1715]) );
  INVD0 U1724 ( .I(1'b1), .ZN(n[1716]) );
  INVD0 U1726 ( .I(1'b1), .ZN(n[1722]) );
  INVD0 U1728 ( .I(1'b1), .ZN(n[1723]) );
  INVD0 U1730 ( .I(1'b1), .ZN(n[1725]) );
  INVD0 U1732 ( .I(1'b1), .ZN(n[1726]) );
  INVD0 U1734 ( .I(1'b1), .ZN(n[1729]) );
  INVD0 U1736 ( .I(1'b1), .ZN(n[1730]) );
  INVD0 U1738 ( .I(1'b1), .ZN(n[1732]) );
  INVD0 U1740 ( .I(1'b1), .ZN(n[1733]) );
  INVD0 U1742 ( .I(1'b1), .ZN(n[1737]) );
  INVD0 U1744 ( .I(1'b1), .ZN(n[1738]) );
  INVD0 U1746 ( .I(1'b1), .ZN(n[1740]) );
  INVD0 U1748 ( .I(1'b1), .ZN(n[1741]) );
  INVD0 U1750 ( .I(1'b1), .ZN(n[1744]) );
  INVD0 U1752 ( .I(1'b1), .ZN(n[1745]) );
  INVD0 U1754 ( .I(1'b1), .ZN(n[1747]) );
  INVD0 U1756 ( .I(1'b1), .ZN(n[1748]) );
  INVD0 U1758 ( .I(1'b1), .ZN(n[1753]) );
  INVD0 U1760 ( .I(1'b1), .ZN(n[1754]) );
  INVD0 U1762 ( .I(1'b1), .ZN(n[1756]) );
  INVD0 U1764 ( .I(1'b1), .ZN(n[1757]) );
  INVD0 U1766 ( .I(1'b1), .ZN(n[1760]) );
  INVD0 U1768 ( .I(1'b1), .ZN(n[1761]) );
  INVD0 U1770 ( .I(1'b1), .ZN(n[1763]) );
  INVD0 U1772 ( .I(1'b1), .ZN(n[1764]) );
  INVD0 U1774 ( .I(1'b1), .ZN(n[1768]) );
  INVD0 U1776 ( .I(1'b1), .ZN(n[1769]) );
  INVD0 U1778 ( .I(1'b1), .ZN(n[1771]) );
  INVD0 U1780 ( .I(1'b1), .ZN(n[1772]) );
  INVD0 U1782 ( .I(1'b1), .ZN(n[1775]) );
  INVD0 U1784 ( .I(1'b1), .ZN(n[1776]) );
  INVD0 U1786 ( .I(1'b1), .ZN(n[1778]) );
  INVD0 U1788 ( .I(1'b1), .ZN(n[1779]) );
  INVD0 U1790 ( .I(1'b1), .ZN(n[1787]) );
  INVD0 U1792 ( .I(1'b1), .ZN(n[1788]) );
  INVD0 U1794 ( .I(1'b1), .ZN(n[1790]) );
  INVD0 U1796 ( .I(1'b1), .ZN(n[1791]) );
  INVD0 U1798 ( .I(1'b1), .ZN(n[1794]) );
  INVD0 U1800 ( .I(1'b1), .ZN(n[1795]) );
  INVD0 U1802 ( .I(1'b1), .ZN(n[1797]) );
  INVD0 U1804 ( .I(1'b1), .ZN(n[1798]) );
  INVD0 U1806 ( .I(1'b1), .ZN(n[1802]) );
  INVD0 U1808 ( .I(1'b1), .ZN(n[1803]) );
  INVD0 U1810 ( .I(1'b1), .ZN(n[1805]) );
  INVD0 U1812 ( .I(1'b1), .ZN(n[1806]) );
  INVD0 U1814 ( .I(1'b1), .ZN(n[1809]) );
  INVD0 U1816 ( .I(1'b1), .ZN(n[1810]) );
  INVD0 U1818 ( .I(1'b1), .ZN(n[1812]) );
  INVD0 U1820 ( .I(1'b1), .ZN(n[1813]) );
  INVD0 U1822 ( .I(1'b1), .ZN(n[1818]) );
  INVD0 U1824 ( .I(1'b1), .ZN(n[1819]) );
  INVD0 U1826 ( .I(1'b1), .ZN(n[1821]) );
  INVD0 U1828 ( .I(1'b1), .ZN(n[1822]) );
  INVD0 U1830 ( .I(1'b1), .ZN(n[1825]) );
  INVD0 U1832 ( .I(1'b1), .ZN(n[1826]) );
  INVD0 U1834 ( .I(1'b1), .ZN(n[1828]) );
  INVD0 U1836 ( .I(1'b1), .ZN(n[1829]) );
  INVD0 U1838 ( .I(1'b1), .ZN(n[1833]) );
  INVD0 U1840 ( .I(1'b1), .ZN(n[1834]) );
  INVD0 U1842 ( .I(1'b1), .ZN(n[1836]) );
  INVD0 U1844 ( .I(1'b1), .ZN(n[1837]) );
  INVD0 U1846 ( .I(1'b1), .ZN(n[1840]) );
  INVD0 U1848 ( .I(1'b1), .ZN(n[1841]) );
  INVD0 U1850 ( .I(1'b1), .ZN(n[1843]) );
  INVD0 U1852 ( .I(1'b1), .ZN(n[1844]) );
  INVD0 U1854 ( .I(1'b1), .ZN(n[1850]) );
  INVD0 U1856 ( .I(1'b1), .ZN(n[1851]) );
  INVD0 U1858 ( .I(1'b1), .ZN(n[1853]) );
  INVD0 U1860 ( .I(1'b1), .ZN(n[1854]) );
  INVD0 U1862 ( .I(1'b1), .ZN(n[1857]) );
  INVD0 U1864 ( .I(1'b1), .ZN(n[1858]) );
  INVD0 U1866 ( .I(1'b1), .ZN(n[1860]) );
  INVD0 U1868 ( .I(1'b1), .ZN(n[1861]) );
  INVD0 U1870 ( .I(1'b1), .ZN(n[1865]) );
  INVD0 U1872 ( .I(1'b1), .ZN(n[1866]) );
  INVD0 U1874 ( .I(1'b1), .ZN(n[1868]) );
  INVD0 U1876 ( .I(1'b1), .ZN(n[1869]) );
  INVD0 U1878 ( .I(1'b1), .ZN(n[1872]) );
  INVD0 U1880 ( .I(1'b1), .ZN(n[1873]) );
  INVD0 U1882 ( .I(1'b1), .ZN(n[1875]) );
  INVD0 U1884 ( .I(1'b1), .ZN(n[1876]) );
  INVD0 U1886 ( .I(1'b1), .ZN(n[1881]) );
  INVD0 U1888 ( .I(1'b1), .ZN(n[1882]) );
  INVD0 U1890 ( .I(1'b1), .ZN(n[1884]) );
  INVD0 U1892 ( .I(1'b1), .ZN(n[1885]) );
  INVD0 U1894 ( .I(1'b1), .ZN(n[1888]) );
  INVD0 U1896 ( .I(1'b1), .ZN(n[1889]) );
  INVD0 U1898 ( .I(1'b1), .ZN(n[1891]) );
  INVD0 U1900 ( .I(1'b1), .ZN(n[1892]) );
  INVD0 U1902 ( .I(1'b1), .ZN(n[1896]) );
  INVD0 U1904 ( .I(1'b1), .ZN(n[1897]) );
  INVD0 U1906 ( .I(1'b1), .ZN(n[1899]) );
  INVD0 U1908 ( .I(1'b1), .ZN(n[1900]) );
  INVD0 U1910 ( .I(1'b1), .ZN(n[1903]) );
  INVD0 U1912 ( .I(1'b1), .ZN(n[1904]) );
  INVD0 U1914 ( .I(1'b1), .ZN(n[1906]) );
  INVD0 U1916 ( .I(1'b1), .ZN(n[1907]) );
  INVD0 U1918 ( .I(1'b1), .ZN(n[1914]) );
  INVD0 U1920 ( .I(1'b1), .ZN(n[1915]) );
  INVD0 U1922 ( .I(1'b1), .ZN(n[1917]) );
  INVD0 U1924 ( .I(1'b1), .ZN(n[1918]) );
  INVD0 U1926 ( .I(1'b1), .ZN(n[1921]) );
  INVD0 U1928 ( .I(1'b1), .ZN(n[1922]) );
  INVD0 U1930 ( .I(1'b1), .ZN(n[1924]) );
  INVD0 U1932 ( .I(1'b1), .ZN(n[1925]) );
  INVD0 U1934 ( .I(1'b1), .ZN(n[1929]) );
  INVD0 U1936 ( .I(1'b1), .ZN(n[1930]) );
  INVD0 U1938 ( .I(1'b1), .ZN(n[1932]) );
  INVD0 U1940 ( .I(1'b1), .ZN(n[1933]) );
  INVD0 U1942 ( .I(1'b1), .ZN(n[1936]) );
  INVD0 U1944 ( .I(1'b1), .ZN(n[1937]) );
  INVD0 U1946 ( .I(1'b1), .ZN(n[1939]) );
  INVD0 U1948 ( .I(1'b1), .ZN(n[1940]) );
  INVD0 U1950 ( .I(1'b1), .ZN(n[1945]) );
  INVD0 U1952 ( .I(1'b1), .ZN(n[1946]) );
  INVD0 U1954 ( .I(1'b1), .ZN(n[1948]) );
  INVD0 U1956 ( .I(1'b1), .ZN(n[1949]) );
  INVD0 U1958 ( .I(1'b1), .ZN(n[1952]) );
  INVD0 U1960 ( .I(1'b1), .ZN(n[1953]) );
  INVD0 U1962 ( .I(1'b1), .ZN(n[1955]) );
  INVD0 U1964 ( .I(1'b1), .ZN(n[1956]) );
  INVD0 U1966 ( .I(1'b1), .ZN(n[1960]) );
  INVD0 U1968 ( .I(1'b1), .ZN(n[1961]) );
  INVD0 U1970 ( .I(1'b1), .ZN(n[1963]) );
  INVD0 U1972 ( .I(1'b1), .ZN(n[1964]) );
  INVD0 U1974 ( .I(1'b1), .ZN(n[1967]) );
  INVD0 U1976 ( .I(1'b1), .ZN(n[1968]) );
  INVD0 U1978 ( .I(1'b1), .ZN(n[1970]) );
  INVD0 U1980 ( .I(1'b1), .ZN(n[1971]) );
  INVD0 U1982 ( .I(1'b1), .ZN(n[1977]) );
  INVD0 U1984 ( .I(1'b1), .ZN(n[1978]) );
  INVD0 U1986 ( .I(1'b1), .ZN(n[1980]) );
  INVD0 U1988 ( .I(1'b1), .ZN(n[1981]) );
  INVD0 U1990 ( .I(1'b1), .ZN(n[1984]) );
  INVD0 U1992 ( .I(1'b1), .ZN(n[1985]) );
  INVD0 U1994 ( .I(1'b1), .ZN(n[1987]) );
  INVD0 U1996 ( .I(1'b1), .ZN(n[1988]) );
  INVD0 U1998 ( .I(1'b1), .ZN(n[1992]) );
  INVD0 U2000 ( .I(1'b1), .ZN(n[1993]) );
  INVD0 U2002 ( .I(1'b1), .ZN(n[1995]) );
  INVD0 U2004 ( .I(1'b1), .ZN(n[1996]) );
  INVD0 U2006 ( .I(1'b1), .ZN(n[1999]) );
  INVD0 U2008 ( .I(1'b1), .ZN(n[2000]) );
  INVD0 U2010 ( .I(1'b1), .ZN(n[2002]) );
  INVD0 U2012 ( .I(1'b1), .ZN(n[2003]) );
  INVD0 U2014 ( .I(1'b1), .ZN(n[2008]) );
  INVD0 U2016 ( .I(1'b1), .ZN(n[2009]) );
  INVD0 U2018 ( .I(1'b1), .ZN(n[2011]) );
  INVD0 U2020 ( .I(1'b1), .ZN(n[2012]) );
  INVD0 U2022 ( .I(1'b1), .ZN(n[2015]) );
  INVD0 U2024 ( .I(1'b1), .ZN(n[2016]) );
  INVD0 U2026 ( .I(1'b1), .ZN(n[2018]) );
  INVD0 U2028 ( .I(1'b1), .ZN(n[2019]) );
  INVD0 U2030 ( .I(1'b1), .ZN(n[2023]) );
  INVD0 U2032 ( .I(1'b1), .ZN(n[2024]) );
  INVD0 U2034 ( .I(1'b1), .ZN(n[2026]) );
  INVD0 U2036 ( .I(1'b1), .ZN(n[2027]) );
  INVD0 U2039 ( .I(1'b1), .ZN(n[2030]) );
  INVD0 U2041 ( .I(1'b1), .ZN(n[2031]) );
  INVD0 U2043 ( .I(1'b1), .ZN(n[2033]) );
  INVD0 U2045 ( .I(1'b1), .ZN(n[2034]) );
  INVD0 U2047 ( .I(1'b1), .ZN(n[2045]) );
  INVD0 U2049 ( .I(1'b1), .ZN(n[2046]) );
  INVD0 U2051 ( .I(1'b1), .ZN(n[2048]) );
  INVD0 U2053 ( .I(1'b1), .ZN(n[2049]) );
  INVD0 U2055 ( .I(1'b1), .ZN(n[2052]) );
  INVD0 U2057 ( .I(1'b1), .ZN(n[2053]) );
  INVD0 U2059 ( .I(1'b1), .ZN(n[2055]) );
  INVD0 U2061 ( .I(1'b1), .ZN(n[2056]) );
  INVD0 U2063 ( .I(1'b1), .ZN(n[2060]) );
  INVD0 U2065 ( .I(1'b1), .ZN(n[2061]) );
  INVD0 U2067 ( .I(1'b1), .ZN(n[2063]) );
  INVD0 U2069 ( .I(1'b1), .ZN(n[2064]) );
  INVD0 U2071 ( .I(1'b1), .ZN(n[2067]) );
  INVD0 U2073 ( .I(1'b1), .ZN(n[2068]) );
  INVD0 U2075 ( .I(1'b1), .ZN(n[2070]) );
  INVD0 U2077 ( .I(1'b1), .ZN(n[2071]) );
  INVD0 U2079 ( .I(1'b1), .ZN(n[2076]) );
  INVD0 U2081 ( .I(1'b1), .ZN(n[2077]) );
  INVD0 U2083 ( .I(1'b1), .ZN(n[2079]) );
  INVD0 U2085 ( .I(1'b1), .ZN(n[2080]) );
  INVD0 U2087 ( .I(1'b1), .ZN(n[2083]) );
  INVD0 U2089 ( .I(1'b1), .ZN(n[2084]) );
  INVD0 U2091 ( .I(1'b1), .ZN(n[2086]) );
  INVD0 U2093 ( .I(1'b1), .ZN(n[2087]) );
  INVD0 U2095 ( .I(1'b1), .ZN(n[2091]) );
  INVD0 U2097 ( .I(1'b1), .ZN(n[2092]) );
  INVD0 U2099 ( .I(1'b1), .ZN(n[2094]) );
  INVD0 U2101 ( .I(1'b1), .ZN(n[2095]) );
  INVD0 U2103 ( .I(1'b1), .ZN(n[2098]) );
  INVD0 U2105 ( .I(1'b1), .ZN(n[2099]) );
  INVD0 U2107 ( .I(1'b1), .ZN(n[2101]) );
  INVD0 U2109 ( .I(1'b1), .ZN(n[2102]) );
  INVD0 U2111 ( .I(1'b1), .ZN(n[2108]) );
  INVD0 U2113 ( .I(1'b1), .ZN(n[2109]) );
  INVD0 U2115 ( .I(1'b1), .ZN(n[2111]) );
  INVD0 U2117 ( .I(1'b1), .ZN(n[2112]) );
  INVD0 U2119 ( .I(1'b1), .ZN(n[2115]) );
  INVD0 U2121 ( .I(1'b1), .ZN(n[2116]) );
  INVD0 U2123 ( .I(1'b1), .ZN(n[2118]) );
  INVD0 U2125 ( .I(1'b1), .ZN(n[2119]) );
  INVD0 U2127 ( .I(1'b1), .ZN(n[2123]) );
  INVD0 U2129 ( .I(1'b1), .ZN(n[2124]) );
  INVD0 U2131 ( .I(1'b1), .ZN(n[2126]) );
  INVD0 U2133 ( .I(1'b1), .ZN(n[2127]) );
  INVD0 U2135 ( .I(1'b1), .ZN(n[2130]) );
  INVD0 U2137 ( .I(1'b1), .ZN(n[2131]) );
  INVD0 U2139 ( .I(1'b1), .ZN(n[2133]) );
  INVD0 U2141 ( .I(1'b1), .ZN(n[2134]) );
  INVD0 U2143 ( .I(1'b1), .ZN(n[2139]) );
  INVD0 U2145 ( .I(1'b1), .ZN(n[2140]) );
  INVD0 U2147 ( .I(1'b1), .ZN(n[2142]) );
  INVD0 U2149 ( .I(1'b1), .ZN(n[2143]) );
  INVD0 U2151 ( .I(1'b1), .ZN(n[2146]) );
  INVD0 U2153 ( .I(1'b1), .ZN(n[2147]) );
  INVD0 U2155 ( .I(1'b1), .ZN(n[2149]) );
  INVD0 U2157 ( .I(1'b1), .ZN(n[2150]) );
  INVD0 U2159 ( .I(1'b1), .ZN(n[2154]) );
  INVD0 U2161 ( .I(1'b1), .ZN(n[2155]) );
  INVD0 U2163 ( .I(1'b1), .ZN(n[2157]) );
  INVD0 U2165 ( .I(1'b1), .ZN(n[2158]) );
  INVD0 U2167 ( .I(1'b1), .ZN(n[2161]) );
  INVD0 U2169 ( .I(1'b1), .ZN(n[2162]) );
  INVD0 U2171 ( .I(1'b1), .ZN(n[2164]) );
  INVD0 U2173 ( .I(1'b1), .ZN(n[2165]) );
  INVD0 U2175 ( .I(1'b1), .ZN(n[2172]) );
  INVD0 U2177 ( .I(1'b1), .ZN(n[2173]) );
  INVD0 U2179 ( .I(1'b1), .ZN(n[2175]) );
  INVD0 U2181 ( .I(1'b1), .ZN(n[2176]) );
  INVD0 U2183 ( .I(1'b1), .ZN(n[2179]) );
  INVD0 U2185 ( .I(1'b1), .ZN(n[2180]) );
  INVD0 U2187 ( .I(1'b1), .ZN(n[2182]) );
  INVD0 U2189 ( .I(1'b1), .ZN(n[2183]) );
  INVD0 U2191 ( .I(1'b1), .ZN(n[2187]) );
  INVD0 U2193 ( .I(1'b1), .ZN(n[2188]) );
  INVD0 U2195 ( .I(1'b1), .ZN(n[2190]) );
  INVD0 U2197 ( .I(1'b1), .ZN(n[2191]) );
  INVD0 U2199 ( .I(1'b1), .ZN(n[2194]) );
  INVD0 U2201 ( .I(1'b1), .ZN(n[2195]) );
  INVD0 U2203 ( .I(1'b1), .ZN(n[2197]) );
  INVD0 U2205 ( .I(1'b1), .ZN(n[2198]) );
  INVD0 U2207 ( .I(1'b1), .ZN(n[2203]) );
  INVD0 U2209 ( .I(1'b1), .ZN(n[2204]) );
  INVD0 U2211 ( .I(1'b1), .ZN(n[2206]) );
  INVD0 U2213 ( .I(1'b1), .ZN(n[2207]) );
  INVD0 U2215 ( .I(1'b1), .ZN(n[2210]) );
  INVD0 U2217 ( .I(1'b1), .ZN(n[2211]) );
  INVD0 U2219 ( .I(1'b1), .ZN(n[2213]) );
  INVD0 U2221 ( .I(1'b1), .ZN(n[2214]) );
  INVD0 U2223 ( .I(1'b1), .ZN(n[2218]) );
  INVD0 U2225 ( .I(1'b1), .ZN(n[2219]) );
  INVD0 U2227 ( .I(1'b1), .ZN(n[2221]) );
  INVD0 U2229 ( .I(1'b1), .ZN(n[2222]) );
  INVD0 U2231 ( .I(1'b1), .ZN(n[2225]) );
  INVD0 U2233 ( .I(1'b1), .ZN(n[2226]) );
  INVD0 U2235 ( .I(1'b1), .ZN(n[2228]) );
  INVD0 U2237 ( .I(1'b1), .ZN(n[2229]) );
  INVD0 U2239 ( .I(1'b1), .ZN(n[2235]) );
  INVD0 U2241 ( .I(1'b1), .ZN(n[2236]) );
  INVD0 U2243 ( .I(1'b1), .ZN(n[2238]) );
  INVD0 U2245 ( .I(1'b1), .ZN(n[2239]) );
  INVD0 U2247 ( .I(1'b1), .ZN(n[2242]) );
  INVD0 U2249 ( .I(1'b1), .ZN(n[2243]) );
  INVD0 U2251 ( .I(1'b1), .ZN(n[2245]) );
  INVD0 U2253 ( .I(1'b1), .ZN(n[2246]) );
  INVD0 U2255 ( .I(1'b1), .ZN(n[2250]) );
  INVD0 U2257 ( .I(1'b1), .ZN(n[2251]) );
  INVD0 U2259 ( .I(1'b1), .ZN(n[2253]) );
  INVD0 U2261 ( .I(1'b1), .ZN(n[2254]) );
  INVD0 U2263 ( .I(1'b1), .ZN(n[2257]) );
  INVD0 U2265 ( .I(1'b1), .ZN(n[2258]) );
  INVD0 U2267 ( .I(1'b1), .ZN(n[2260]) );
  INVD0 U2269 ( .I(1'b1), .ZN(n[2261]) );
  INVD0 U2271 ( .I(1'b1), .ZN(n[2266]) );
  INVD0 U2273 ( .I(1'b1), .ZN(n[2267]) );
  INVD0 U2275 ( .I(1'b1), .ZN(n[2269]) );
  INVD0 U2277 ( .I(1'b1), .ZN(n[2270]) );
  INVD0 U2279 ( .I(1'b1), .ZN(n[2273]) );
  INVD0 U2281 ( .I(1'b1), .ZN(n[2274]) );
  INVD0 U2283 ( .I(1'b1), .ZN(n[2276]) );
  INVD0 U2285 ( .I(1'b1), .ZN(n[2277]) );
  INVD0 U2287 ( .I(1'b1), .ZN(n[2281]) );
  INVD0 U2289 ( .I(1'b1), .ZN(n[2282]) );
  INVD0 U2291 ( .I(1'b1), .ZN(n[2284]) );
  INVD0 U2293 ( .I(1'b1), .ZN(n[2285]) );
  INVD0 U2295 ( .I(1'b1), .ZN(n[2288]) );
  INVD0 U2297 ( .I(1'b1), .ZN(n[2289]) );
  INVD0 U2299 ( .I(1'b1), .ZN(n[2291]) );
  INVD0 U2301 ( .I(1'b1), .ZN(n[2292]) );
  INVD0 U2303 ( .I(1'b1), .ZN(n[2300]) );
  INVD0 U2305 ( .I(1'b1), .ZN(n[2301]) );
  INVD0 U2307 ( .I(1'b1), .ZN(n[2303]) );
  INVD0 U2309 ( .I(1'b1), .ZN(n[2304]) );
  INVD0 U2311 ( .I(1'b1), .ZN(n[2307]) );
  INVD0 U2313 ( .I(1'b1), .ZN(n[2308]) );
  INVD0 U2315 ( .I(1'b1), .ZN(n[2310]) );
  INVD0 U2317 ( .I(1'b1), .ZN(n[2311]) );
  INVD0 U2319 ( .I(1'b1), .ZN(n[2315]) );
  INVD0 U2321 ( .I(1'b1), .ZN(n[2316]) );
  INVD0 U2323 ( .I(1'b1), .ZN(n[2318]) );
  INVD0 U2325 ( .I(1'b1), .ZN(n[2319]) );
  INVD0 U2327 ( .I(1'b1), .ZN(n[2322]) );
  INVD0 U2329 ( .I(1'b1), .ZN(n[2323]) );
  INVD0 U2331 ( .I(1'b1), .ZN(n[2325]) );
  INVD0 U2333 ( .I(1'b1), .ZN(n[2326]) );
  INVD0 U2335 ( .I(1'b1), .ZN(n[2331]) );
  INVD0 U2337 ( .I(1'b1), .ZN(n[2332]) );
  INVD0 U2339 ( .I(1'b1), .ZN(n[2334]) );
  INVD0 U2341 ( .I(1'b1), .ZN(n[2335]) );
  INVD0 U2343 ( .I(1'b1), .ZN(n[2338]) );
  INVD0 U2345 ( .I(1'b1), .ZN(n[2339]) );
  INVD0 U2347 ( .I(1'b1), .ZN(n[2341]) );
  INVD0 U2349 ( .I(1'b1), .ZN(n[2342]) );
  INVD0 U2351 ( .I(1'b1), .ZN(n[2346]) );
  INVD0 U2353 ( .I(1'b1), .ZN(n[2347]) );
  INVD0 U2355 ( .I(1'b1), .ZN(n[2349]) );
  INVD0 U2357 ( .I(1'b1), .ZN(n[2350]) );
  INVD0 U2359 ( .I(1'b1), .ZN(n[2353]) );
  INVD0 U2361 ( .I(1'b1), .ZN(n[2354]) );
  INVD0 U2363 ( .I(1'b1), .ZN(n[2356]) );
  INVD0 U2365 ( .I(1'b1), .ZN(n[2357]) );
  INVD0 U2367 ( .I(1'b1), .ZN(n[2363]) );
  INVD0 U2369 ( .I(1'b1), .ZN(n[2364]) );
  INVD0 U2371 ( .I(1'b1), .ZN(n[2366]) );
  INVD0 U2373 ( .I(1'b1), .ZN(n[2367]) );
  INVD0 U2375 ( .I(1'b1), .ZN(n[2370]) );
  INVD0 U2377 ( .I(1'b1), .ZN(n[2371]) );
  INVD0 U2379 ( .I(1'b1), .ZN(n[2373]) );
  INVD0 U2381 ( .I(1'b1), .ZN(n[2374]) );
  INVD0 U2383 ( .I(1'b1), .ZN(n[2378]) );
  INVD0 U2385 ( .I(1'b1), .ZN(n[2379]) );
  INVD0 U2387 ( .I(1'b1), .ZN(n[2381]) );
  INVD0 U2389 ( .I(1'b1), .ZN(n[2382]) );
  INVD0 U2391 ( .I(1'b1), .ZN(n[2385]) );
  INVD0 U2393 ( .I(1'b1), .ZN(n[2386]) );
  INVD0 U2395 ( .I(1'b1), .ZN(n[2388]) );
  INVD0 U2397 ( .I(1'b1), .ZN(n[2389]) );
  INVD0 U2399 ( .I(1'b1), .ZN(n[2394]) );
  INVD0 U2401 ( .I(1'b1), .ZN(n[2395]) );
  INVD0 U2403 ( .I(1'b1), .ZN(n[2397]) );
  INVD0 U2405 ( .I(1'b1), .ZN(n[2398]) );
  INVD0 U2407 ( .I(1'b1), .ZN(n[2401]) );
  INVD0 U2409 ( .I(1'b1), .ZN(n[2402]) );
  INVD0 U2411 ( .I(1'b1), .ZN(n[2404]) );
  INVD0 U2413 ( .I(1'b1), .ZN(n[2405]) );
  INVD0 U2415 ( .I(1'b1), .ZN(n[2409]) );
  INVD0 U2417 ( .I(1'b1), .ZN(n[2410]) );
  INVD0 U2419 ( .I(1'b1), .ZN(n[2412]) );
  INVD0 U2421 ( .I(1'b1), .ZN(n[2413]) );
  INVD0 U2423 ( .I(1'b1), .ZN(n[2416]) );
  INVD0 U2425 ( .I(1'b1), .ZN(n[2417]) );
  INVD0 U2427 ( .I(1'b1), .ZN(n[2419]) );
  INVD0 U2429 ( .I(1'b1), .ZN(n[2420]) );
  INVD0 U2431 ( .I(1'b1), .ZN(n[2427]) );
  INVD0 U2433 ( .I(1'b1), .ZN(n[2428]) );
  INVD0 U2435 ( .I(1'b1), .ZN(n[2430]) );
  INVD0 U2437 ( .I(1'b1), .ZN(n[2431]) );
  INVD0 U2439 ( .I(1'b1), .ZN(n[2434]) );
  INVD0 U2441 ( .I(1'b1), .ZN(n[2435]) );
  INVD0 U2443 ( .I(1'b1), .ZN(n[2437]) );
  INVD0 U2445 ( .I(1'b1), .ZN(n[2438]) );
  INVD0 U2447 ( .I(1'b1), .ZN(n[2442]) );
  INVD0 U2449 ( .I(1'b1), .ZN(n[2443]) );
  INVD0 U2451 ( .I(1'b1), .ZN(n[2445]) );
  INVD0 U2453 ( .I(1'b1), .ZN(n[2446]) );
  INVD0 U2455 ( .I(1'b1), .ZN(n[2449]) );
  INVD0 U2457 ( .I(1'b1), .ZN(n[2450]) );
  INVD0 U2459 ( .I(1'b1), .ZN(n[2452]) );
  INVD0 U2461 ( .I(1'b1), .ZN(n[2453]) );
  INVD0 U2463 ( .I(1'b1), .ZN(n[2458]) );
  INVD0 U2465 ( .I(1'b1), .ZN(n[2459]) );
  INVD0 U2467 ( .I(1'b1), .ZN(n[2461]) );
  INVD0 U2469 ( .I(1'b1), .ZN(n[2462]) );
  INVD0 U2471 ( .I(1'b1), .ZN(n[2465]) );
  INVD0 U2473 ( .I(1'b1), .ZN(n[2466]) );
  INVD0 U2475 ( .I(1'b1), .ZN(n[2468]) );
  INVD0 U2477 ( .I(1'b1), .ZN(n[2469]) );
  INVD0 U2479 ( .I(1'b1), .ZN(n[2473]) );
  INVD0 U2481 ( .I(1'b1), .ZN(n[2474]) );
  INVD0 U2483 ( .I(1'b1), .ZN(n[2476]) );
  INVD0 U2485 ( .I(1'b1), .ZN(n[2477]) );
  INVD0 U2487 ( .I(1'b1), .ZN(n[2480]) );
  INVD0 U2489 ( .I(1'b1), .ZN(n[2481]) );
  INVD0 U2491 ( .I(1'b1), .ZN(n[2483]) );
  INVD0 U2493 ( .I(1'b1), .ZN(n[2484]) );
  INVD0 U2495 ( .I(1'b1), .ZN(n[2490]) );
  INVD0 U2497 ( .I(1'b1), .ZN(n[2491]) );
  INVD0 U2499 ( .I(1'b1), .ZN(n[2493]) );
  INVD0 U2501 ( .I(1'b1), .ZN(n[2494]) );
  INVD0 U2503 ( .I(1'b1), .ZN(n[2497]) );
  INVD0 U2505 ( .I(1'b1), .ZN(n[2498]) );
  INVD0 U2507 ( .I(1'b1), .ZN(n[2500]) );
  INVD0 U2509 ( .I(1'b1), .ZN(n[2501]) );
  INVD0 U2511 ( .I(1'b1), .ZN(n[2505]) );
  INVD0 U2513 ( .I(1'b1), .ZN(n[2506]) );
  INVD0 U2515 ( .I(1'b1), .ZN(n[2508]) );
  INVD0 U2517 ( .I(1'b1), .ZN(n[2509]) );
  INVD0 U2519 ( .I(1'b1), .ZN(n[2512]) );
  INVD0 U2521 ( .I(1'b1), .ZN(n[2513]) );
  INVD0 U2523 ( .I(1'b1), .ZN(n[2515]) );
  INVD0 U2525 ( .I(1'b1), .ZN(n[2516]) );
  INVD0 U2527 ( .I(1'b1), .ZN(n[2521]) );
  INVD0 U2529 ( .I(1'b1), .ZN(n[2522]) );
  INVD0 U2531 ( .I(1'b1), .ZN(n[2524]) );
  INVD0 U2533 ( .I(1'b1), .ZN(n[2525]) );
  INVD0 U2535 ( .I(1'b1), .ZN(n[2528]) );
  INVD0 U2537 ( .I(1'b1), .ZN(n[2529]) );
  INVD0 U2539 ( .I(1'b1), .ZN(n[2531]) );
  INVD0 U2541 ( .I(1'b1), .ZN(n[2532]) );
  INVD0 U2543 ( .I(1'b1), .ZN(n[2536]) );
  INVD0 U2545 ( .I(1'b1), .ZN(n[2537]) );
  INVD0 U2547 ( .I(1'b1), .ZN(n[2539]) );
  INVD0 U2549 ( .I(1'b1), .ZN(n[2540]) );
  INVD0 U2551 ( .I(1'b1), .ZN(n[2543]) );
  INVD0 U2553 ( .I(1'b1), .ZN(n[2544]) );
  INVD0 U2555 ( .I(1'b1), .ZN(n[2546]) );
  INVD0 U2557 ( .I(1'b1), .ZN(n[2547]) );
  INVD0 U2559 ( .I(1'b1), .ZN(n[2556]) );
  INVD0 U2561 ( .I(1'b1), .ZN(n[2557]) );
  INVD0 U2563 ( .I(1'b1), .ZN(n[2559]) );
  INVD0 U2565 ( .I(1'b1), .ZN(n[2560]) );
  INVD0 U2567 ( .I(1'b1), .ZN(n[2563]) );
  INVD0 U2569 ( .I(1'b1), .ZN(n[2564]) );
  INVD0 U2571 ( .I(1'b1), .ZN(n[2566]) );
  INVD0 U2573 ( .I(1'b1), .ZN(n[2567]) );
  INVD0 U2575 ( .I(1'b1), .ZN(n[2571]) );
  INVD0 U2577 ( .I(1'b1), .ZN(n[2572]) );
  INVD0 U2579 ( .I(1'b1), .ZN(n[2574]) );
  INVD0 U2581 ( .I(1'b1), .ZN(n[2575]) );
  INVD0 U2583 ( .I(1'b1), .ZN(n[2578]) );
  INVD0 U2585 ( .I(1'b1), .ZN(n[2579]) );
  INVD0 U2587 ( .I(1'b1), .ZN(n[2581]) );
  INVD0 U2589 ( .I(1'b1), .ZN(n[2582]) );
  INVD0 U2591 ( .I(1'b1), .ZN(n[2587]) );
  INVD0 U2593 ( .I(1'b1), .ZN(n[2588]) );
  INVD0 U2595 ( .I(1'b1), .ZN(n[2590]) );
  INVD0 U2597 ( .I(1'b1), .ZN(n[2591]) );
  INVD0 U2599 ( .I(1'b1), .ZN(n[2594]) );
  INVD0 U2601 ( .I(1'b1), .ZN(n[2595]) );
  INVD0 U2603 ( .I(1'b1), .ZN(n[2597]) );
  INVD0 U2605 ( .I(1'b1), .ZN(n[2598]) );
  INVD0 U2607 ( .I(1'b1), .ZN(n[2602]) );
  INVD0 U2609 ( .I(1'b1), .ZN(n[2603]) );
  INVD0 U2611 ( .I(1'b1), .ZN(n[2605]) );
  INVD0 U2613 ( .I(1'b1), .ZN(n[2606]) );
  INVD0 U2615 ( .I(1'b1), .ZN(n[2609]) );
  INVD0 U2617 ( .I(1'b1), .ZN(n[2610]) );
  INVD0 U2619 ( .I(1'b1), .ZN(n[2612]) );
  INVD0 U2621 ( .I(1'b1), .ZN(n[2613]) );
  INVD0 U2623 ( .I(1'b1), .ZN(n[2619]) );
  INVD0 U2625 ( .I(1'b1), .ZN(n[2620]) );
  INVD0 U2627 ( .I(1'b1), .ZN(n[2622]) );
  INVD0 U2629 ( .I(1'b1), .ZN(n[2623]) );
  INVD0 U2631 ( .I(1'b1), .ZN(n[2626]) );
  INVD0 U2633 ( .I(1'b1), .ZN(n[2627]) );
  INVD0 U2635 ( .I(1'b1), .ZN(n[2629]) );
  INVD0 U2637 ( .I(1'b1), .ZN(n[2630]) );
  INVD0 U2639 ( .I(1'b1), .ZN(n[2634]) );
  INVD0 U2641 ( .I(1'b1), .ZN(n[2635]) );
  INVD0 U2643 ( .I(1'b1), .ZN(n[2637]) );
  INVD0 U2645 ( .I(1'b1), .ZN(n[2638]) );
  INVD0 U2647 ( .I(1'b1), .ZN(n[2641]) );
  INVD0 U2649 ( .I(1'b1), .ZN(n[2642]) );
  INVD0 U2651 ( .I(1'b1), .ZN(n[2644]) );
  INVD0 U2653 ( .I(1'b1), .ZN(n[2645]) );
  INVD0 U2655 ( .I(1'b1), .ZN(n[2650]) );
  INVD0 U2657 ( .I(1'b1), .ZN(n[2651]) );
  INVD0 U2659 ( .I(1'b1), .ZN(n[2653]) );
  INVD0 U2661 ( .I(1'b1), .ZN(n[2654]) );
  INVD0 U2663 ( .I(1'b1), .ZN(n[2657]) );
  INVD0 U2665 ( .I(1'b1), .ZN(n[2658]) );
  INVD0 U2667 ( .I(1'b1), .ZN(n[2660]) );
  INVD0 U2669 ( .I(1'b1), .ZN(n[2661]) );
  INVD0 U2671 ( .I(1'b1), .ZN(n[2665]) );
  INVD0 U2673 ( .I(1'b1), .ZN(n[2666]) );
  INVD0 U2675 ( .I(1'b1), .ZN(n[2668]) );
  INVD0 U2677 ( .I(1'b1), .ZN(n[2669]) );
  INVD0 U2679 ( .I(1'b1), .ZN(n[2672]) );
  INVD0 U2681 ( .I(1'b1), .ZN(n[2673]) );
  INVD0 U2683 ( .I(1'b1), .ZN(n[2675]) );
  INVD0 U2685 ( .I(1'b1), .ZN(n[2676]) );
  INVD0 U2687 ( .I(1'b1), .ZN(n[2683]) );
  INVD0 U2689 ( .I(1'b1), .ZN(n[2684]) );
  INVD0 U2691 ( .I(1'b1), .ZN(n[2686]) );
  INVD0 U2693 ( .I(1'b1), .ZN(n[2687]) );
  INVD0 U2695 ( .I(1'b1), .ZN(n[2690]) );
  INVD0 U2697 ( .I(1'b1), .ZN(n[2691]) );
  INVD0 U2699 ( .I(1'b1), .ZN(n[2693]) );
  INVD0 U2701 ( .I(1'b1), .ZN(n[2694]) );
  INVD0 U2703 ( .I(1'b1), .ZN(n[2698]) );
  INVD0 U2705 ( .I(1'b1), .ZN(n[2699]) );
  INVD0 U2707 ( .I(1'b1), .ZN(n[2701]) );
  INVD0 U2709 ( .I(1'b1), .ZN(n[2702]) );
  INVD0 U2711 ( .I(1'b1), .ZN(n[2705]) );
  INVD0 U2713 ( .I(1'b1), .ZN(n[2706]) );
  INVD0 U2715 ( .I(1'b1), .ZN(n[2708]) );
  INVD0 U2717 ( .I(1'b1), .ZN(n[2709]) );
  INVD0 U2719 ( .I(1'b1), .ZN(n[2714]) );
  INVD0 U2721 ( .I(1'b1), .ZN(n[2715]) );
  INVD0 U2723 ( .I(1'b1), .ZN(n[2717]) );
  INVD0 U2725 ( .I(1'b1), .ZN(n[2718]) );
  INVD0 U2727 ( .I(1'b1), .ZN(n[2721]) );
  INVD0 U2729 ( .I(1'b1), .ZN(n[2722]) );
  INVD0 U2731 ( .I(1'b1), .ZN(n[2724]) );
  INVD0 U2733 ( .I(1'b1), .ZN(n[2725]) );
  INVD0 U2735 ( .I(1'b1), .ZN(n[2729]) );
  INVD0 U2737 ( .I(1'b1), .ZN(n[2730]) );
  INVD0 U2739 ( .I(1'b1), .ZN(n[2732]) );
  INVD0 U2741 ( .I(1'b1), .ZN(n[2733]) );
  INVD0 U2743 ( .I(1'b1), .ZN(n[2736]) );
  INVD0 U2745 ( .I(1'b1), .ZN(n[2737]) );
  INVD0 U2747 ( .I(1'b1), .ZN(n[2739]) );
  INVD0 U2749 ( .I(1'b1), .ZN(n[2740]) );
  INVD0 U2751 ( .I(1'b1), .ZN(n[2746]) );
  INVD0 U2753 ( .I(1'b1), .ZN(n[2747]) );
  INVD0 U2755 ( .I(1'b1), .ZN(n[2749]) );
  INVD0 U2757 ( .I(1'b1), .ZN(n[2750]) );
  INVD0 U2759 ( .I(1'b1), .ZN(n[2753]) );
  INVD0 U2761 ( .I(1'b1), .ZN(n[2754]) );
  INVD0 U2763 ( .I(1'b1), .ZN(n[2756]) );
  INVD0 U2765 ( .I(1'b1), .ZN(n[2757]) );
  INVD0 U2767 ( .I(1'b1), .ZN(n[2761]) );
  INVD0 U2769 ( .I(1'b1), .ZN(n[2762]) );
  INVD0 U2771 ( .I(1'b1), .ZN(n[2764]) );
  INVD0 U2773 ( .I(1'b1), .ZN(n[2765]) );
  INVD0 U2775 ( .I(1'b1), .ZN(n[2768]) );
  INVD0 U2777 ( .I(1'b1), .ZN(n[2769]) );
  INVD0 U2779 ( .I(1'b1), .ZN(n[2771]) );
  INVD0 U2781 ( .I(1'b1), .ZN(n[2772]) );
  INVD0 U2783 ( .I(1'b1), .ZN(n[2777]) );
  INVD0 U2785 ( .I(1'b1), .ZN(n[2778]) );
  INVD0 U2787 ( .I(1'b1), .ZN(n[2780]) );
  INVD0 U2789 ( .I(1'b1), .ZN(n[2781]) );
  INVD0 U2791 ( .I(1'b1), .ZN(n[2784]) );
  INVD0 U2793 ( .I(1'b1), .ZN(n[2785]) );
  INVD0 U2795 ( .I(1'b1), .ZN(n[2787]) );
  INVD0 U2797 ( .I(1'b1), .ZN(n[2788]) );
  INVD0 U2799 ( .I(1'b1), .ZN(n[2792]) );
  INVD0 U2801 ( .I(1'b1), .ZN(n[2793]) );
  INVD0 U2803 ( .I(1'b1), .ZN(n[2795]) );
  INVD0 U2805 ( .I(1'b1), .ZN(n[2796]) );
  INVD0 U2807 ( .I(1'b1), .ZN(n[2799]) );
  INVD0 U2809 ( .I(1'b1), .ZN(n[2800]) );
  INVD0 U2811 ( .I(1'b1), .ZN(n[2802]) );
  INVD0 U2813 ( .I(1'b1), .ZN(n[2803]) );
  INVD0 U2815 ( .I(1'b1), .ZN(n[2811]) );
  INVD0 U2817 ( .I(1'b1), .ZN(n[2812]) );
  INVD0 U2819 ( .I(1'b1), .ZN(n[2814]) );
  INVD0 U2821 ( .I(1'b1), .ZN(n[2815]) );
  INVD0 U2823 ( .I(1'b1), .ZN(n[2818]) );
  INVD0 U2825 ( .I(1'b1), .ZN(n[2819]) );
  INVD0 U2827 ( .I(1'b1), .ZN(n[2821]) );
  INVD0 U2829 ( .I(1'b1), .ZN(n[2822]) );
  INVD0 U2831 ( .I(1'b1), .ZN(n[2826]) );
  INVD0 U2833 ( .I(1'b1), .ZN(n[2827]) );
  INVD0 U2835 ( .I(1'b1), .ZN(n[2829]) );
  INVD0 U2837 ( .I(1'b1), .ZN(n[2830]) );
  INVD0 U2839 ( .I(1'b1), .ZN(n[2833]) );
  INVD0 U2841 ( .I(1'b1), .ZN(n[2834]) );
  INVD0 U2843 ( .I(1'b1), .ZN(n[2836]) );
  INVD0 U2845 ( .I(1'b1), .ZN(n[2837]) );
  INVD0 U2847 ( .I(1'b1), .ZN(n[2842]) );
  INVD0 U2849 ( .I(1'b1), .ZN(n[2843]) );
  INVD0 U2851 ( .I(1'b1), .ZN(n[2845]) );
  INVD0 U2853 ( .I(1'b1), .ZN(n[2846]) );
  INVD0 U2855 ( .I(1'b1), .ZN(n[2849]) );
  INVD0 U2857 ( .I(1'b1), .ZN(n[2850]) );
  INVD0 U2859 ( .I(1'b1), .ZN(n[2852]) );
  INVD0 U2861 ( .I(1'b1), .ZN(n[2853]) );
  INVD0 U2863 ( .I(1'b1), .ZN(n[2857]) );
  INVD0 U2865 ( .I(1'b1), .ZN(n[2858]) );
  INVD0 U2867 ( .I(1'b1), .ZN(n[2860]) );
  INVD0 U2869 ( .I(1'b1), .ZN(n[2861]) );
  INVD0 U2871 ( .I(1'b1), .ZN(n[2864]) );
  INVD0 U2873 ( .I(1'b1), .ZN(n[2865]) );
  INVD0 U2875 ( .I(1'b1), .ZN(n[2867]) );
  INVD0 U2877 ( .I(1'b1), .ZN(n[2868]) );
  INVD0 U2879 ( .I(1'b1), .ZN(n[2874]) );
  INVD0 U2881 ( .I(1'b1), .ZN(n[2875]) );
  INVD0 U2883 ( .I(1'b1), .ZN(n[2877]) );
  INVD0 U2885 ( .I(1'b1), .ZN(n[2878]) );
  INVD0 U2887 ( .I(1'b1), .ZN(n[2881]) );
  INVD0 U2889 ( .I(1'b1), .ZN(n[2882]) );
  INVD0 U2891 ( .I(1'b1), .ZN(n[2884]) );
  INVD0 U2893 ( .I(1'b1), .ZN(n[2885]) );
  INVD0 U2895 ( .I(1'b1), .ZN(n[2889]) );
  INVD0 U2897 ( .I(1'b1), .ZN(n[2890]) );
  INVD0 U2899 ( .I(1'b1), .ZN(n[2892]) );
  INVD0 U2901 ( .I(1'b1), .ZN(n[2893]) );
  INVD0 U2903 ( .I(1'b1), .ZN(n[2896]) );
  INVD0 U2905 ( .I(1'b1), .ZN(n[2897]) );
  INVD0 U2907 ( .I(1'b1), .ZN(n[2899]) );
  INVD0 U2909 ( .I(1'b1), .ZN(n[2900]) );
  INVD0 U2911 ( .I(1'b1), .ZN(n[2905]) );
  INVD0 U2913 ( .I(1'b1), .ZN(n[2906]) );
  INVD0 U2915 ( .I(1'b1), .ZN(n[2908]) );
  INVD0 U2917 ( .I(1'b1), .ZN(n[2909]) );
  INVD0 U2919 ( .I(1'b1), .ZN(n[2912]) );
  INVD0 U2921 ( .I(1'b1), .ZN(n[2913]) );
  INVD0 U2923 ( .I(1'b1), .ZN(n[2915]) );
  INVD0 U2925 ( .I(1'b1), .ZN(n[2916]) );
  INVD0 U2927 ( .I(1'b1), .ZN(n[2920]) );
  INVD0 U2929 ( .I(1'b1), .ZN(n[2921]) );
  INVD0 U2931 ( .I(1'b1), .ZN(n[2923]) );
  INVD0 U2933 ( .I(1'b1), .ZN(n[2924]) );
  INVD0 U2935 ( .I(1'b1), .ZN(n[2927]) );
  INVD0 U2937 ( .I(1'b1), .ZN(n[2928]) );
  INVD0 U2939 ( .I(1'b1), .ZN(n[2930]) );
  INVD0 U2941 ( .I(1'b1), .ZN(n[2931]) );
  INVD0 U2943 ( .I(1'b1), .ZN(n[2938]) );
  INVD0 U2945 ( .I(1'b1), .ZN(n[2939]) );
  INVD0 U2947 ( .I(1'b1), .ZN(n[2941]) );
  INVD0 U2949 ( .I(1'b1), .ZN(n[2942]) );
  INVD0 U2951 ( .I(1'b1), .ZN(n[2945]) );
  INVD0 U2953 ( .I(1'b1), .ZN(n[2946]) );
  INVD0 U2955 ( .I(1'b1), .ZN(n[2948]) );
  INVD0 U2957 ( .I(1'b1), .ZN(n[2949]) );
  INVD0 U2959 ( .I(1'b1), .ZN(n[2953]) );
  INVD0 U2961 ( .I(1'b1), .ZN(n[2954]) );
  INVD0 U2963 ( .I(1'b1), .ZN(n[2956]) );
  INVD0 U2965 ( .I(1'b1), .ZN(n[2957]) );
  INVD0 U2967 ( .I(1'b1), .ZN(n[2960]) );
  INVD0 U2969 ( .I(1'b1), .ZN(n[2961]) );
  INVD0 U2971 ( .I(1'b1), .ZN(n[2963]) );
  INVD0 U2973 ( .I(1'b1), .ZN(n[2964]) );
  INVD0 U2975 ( .I(1'b1), .ZN(n[2969]) );
  INVD0 U2977 ( .I(1'b1), .ZN(n[2970]) );
  INVD0 U2979 ( .I(1'b1), .ZN(n[2972]) );
  INVD0 U2981 ( .I(1'b1), .ZN(n[2973]) );
  INVD0 U2983 ( .I(1'b1), .ZN(n[2976]) );
  INVD0 U2985 ( .I(1'b1), .ZN(n[2977]) );
  INVD0 U2987 ( .I(1'b1), .ZN(n[2979]) );
  INVD0 U2989 ( .I(1'b1), .ZN(n[2980]) );
  INVD0 U2991 ( .I(1'b1), .ZN(n[2984]) );
  INVD0 U2993 ( .I(1'b1), .ZN(n[2985]) );
  INVD0 U2995 ( .I(1'b1), .ZN(n[2987]) );
  INVD0 U2997 ( .I(1'b1), .ZN(n[2988]) );
  INVD0 U2999 ( .I(1'b1), .ZN(n[2991]) );
  INVD0 U3001 ( .I(1'b1), .ZN(n[2992]) );
  INVD0 U3003 ( .I(1'b1), .ZN(n[2994]) );
  INVD0 U3005 ( .I(1'b1), .ZN(n[2995]) );
  INVD0 U3007 ( .I(1'b1), .ZN(n[3001]) );
  INVD0 U3009 ( .I(1'b1), .ZN(n[3002]) );
  INVD0 U3011 ( .I(1'b1), .ZN(n[3004]) );
  INVD0 U3013 ( .I(1'b1), .ZN(n[3005]) );
  INVD0 U3015 ( .I(1'b1), .ZN(n[3008]) );
  INVD0 U3017 ( .I(1'b1), .ZN(n[3009]) );
  INVD0 U3019 ( .I(1'b1), .ZN(n[3011]) );
  INVD0 U3021 ( .I(1'b1), .ZN(n[3012]) );
  INVD0 U3023 ( .I(1'b1), .ZN(n[3016]) );
  INVD0 U3025 ( .I(1'b1), .ZN(n[3017]) );
  INVD0 U3027 ( .I(1'b1), .ZN(n[3019]) );
  INVD0 U3029 ( .I(1'b1), .ZN(n[3020]) );
  INVD0 U3031 ( .I(1'b1), .ZN(n[3023]) );
  INVD0 U3033 ( .I(1'b1), .ZN(n[3024]) );
  INVD0 U3035 ( .I(1'b1), .ZN(n[3026]) );
  INVD0 U3037 ( .I(1'b1), .ZN(n[3027]) );
  INVD0 U3039 ( .I(1'b1), .ZN(n[3032]) );
  INVD0 U3041 ( .I(1'b1), .ZN(n[3033]) );
  INVD0 U3043 ( .I(1'b1), .ZN(n[3035]) );
  INVD0 U3045 ( .I(1'b1), .ZN(n[3036]) );
  INVD0 U3047 ( .I(1'b1), .ZN(n[3039]) );
  INVD0 U3049 ( .I(1'b1), .ZN(n[3040]) );
  INVD0 U3051 ( .I(1'b1), .ZN(n[3042]) );
  INVD0 U3053 ( .I(1'b1), .ZN(n[3043]) );
  INVD0 U3055 ( .I(1'b1), .ZN(n[3047]) );
  INVD0 U3057 ( .I(1'b1), .ZN(n[3048]) );
  INVD0 U3059 ( .I(1'b1), .ZN(n[3050]) );
  INVD0 U3061 ( .I(1'b1), .ZN(n[3051]) );
  INVD0 U3063 ( .I(1'b1), .ZN(n[3054]) );
  INVD0 U3065 ( .I(1'b1), .ZN(n[3055]) );
  INVD0 U3067 ( .I(1'b1), .ZN(n[3057]) );
  INVD0 U3069 ( .I(1'b1), .ZN(n[3058]) );
  INVD0 U3071 ( .I(1'b1), .ZN(n[3068]) );
  INVD0 U3073 ( .I(1'b1), .ZN(n[3069]) );
  INVD0 U3075 ( .I(1'b1), .ZN(n[3071]) );
  INVD0 U3077 ( .I(1'b1), .ZN(n[3072]) );
  INVD0 U3079 ( .I(1'b1), .ZN(n[3075]) );
  INVD0 U3081 ( .I(1'b1), .ZN(n[3076]) );
  INVD0 U3083 ( .I(1'b1), .ZN(n[3078]) );
  INVD0 U3085 ( .I(1'b1), .ZN(n[3079]) );
  INVD0 U3087 ( .I(1'b1), .ZN(n[3083]) );
  INVD0 U3089 ( .I(1'b1), .ZN(n[3084]) );
  INVD0 U3091 ( .I(1'b1), .ZN(n[3086]) );
  INVD0 U3093 ( .I(1'b1), .ZN(n[3087]) );
  INVD0 U3095 ( .I(1'b1), .ZN(n[3090]) );
  INVD0 U3097 ( .I(1'b1), .ZN(n[3091]) );
  INVD0 U3099 ( .I(1'b1), .ZN(n[3093]) );
  INVD0 U3101 ( .I(1'b1), .ZN(n[3094]) );
  INVD0 U3103 ( .I(1'b1), .ZN(n[3099]) );
  INVD0 U3105 ( .I(1'b1), .ZN(n[3100]) );
  INVD0 U3107 ( .I(1'b1), .ZN(n[3102]) );
  INVD0 U3109 ( .I(1'b1), .ZN(n[3103]) );
  INVD0 U3111 ( .I(1'b1), .ZN(n[3106]) );
  INVD0 U3113 ( .I(1'b1), .ZN(n[3107]) );
  INVD0 U3115 ( .I(1'b1), .ZN(n[3109]) );
  INVD0 U3117 ( .I(1'b1), .ZN(n[3110]) );
  INVD0 U3119 ( .I(1'b1), .ZN(n[3114]) );
  INVD0 U3121 ( .I(1'b1), .ZN(n[3115]) );
  INVD0 U3123 ( .I(1'b1), .ZN(n[3117]) );
  INVD0 U3125 ( .I(1'b1), .ZN(n[3118]) );
  INVD0 U3127 ( .I(1'b1), .ZN(n[3121]) );
  INVD0 U3129 ( .I(1'b1), .ZN(n[3122]) );
  INVD0 U3131 ( .I(1'b1), .ZN(n[3124]) );
  INVD0 U3133 ( .I(1'b1), .ZN(n[3125]) );
  INVD0 U3135 ( .I(1'b1), .ZN(n[3131]) );
  INVD0 U3137 ( .I(1'b1), .ZN(n[3132]) );
  INVD0 U3139 ( .I(1'b1), .ZN(n[3134]) );
  INVD0 U3141 ( .I(1'b1), .ZN(n[3135]) );
  INVD0 U3143 ( .I(1'b1), .ZN(n[3138]) );
  INVD0 U3145 ( .I(1'b1), .ZN(n[3139]) );
  INVD0 U3147 ( .I(1'b1), .ZN(n[3141]) );
  INVD0 U3149 ( .I(1'b1), .ZN(n[3142]) );
  INVD0 U3151 ( .I(1'b1), .ZN(n[3146]) );
  INVD0 U3153 ( .I(1'b1), .ZN(n[3147]) );
  INVD0 U3155 ( .I(1'b1), .ZN(n[3149]) );
  INVD0 U3157 ( .I(1'b1), .ZN(n[3150]) );
  INVD0 U3159 ( .I(1'b1), .ZN(n[3153]) );
  INVD0 U3161 ( .I(1'b1), .ZN(n[3154]) );
  INVD0 U3163 ( .I(1'b1), .ZN(n[3156]) );
  INVD0 U3165 ( .I(1'b1), .ZN(n[3157]) );
  INVD0 U3167 ( .I(1'b1), .ZN(n[3162]) );
  INVD0 U3169 ( .I(1'b1), .ZN(n[3163]) );
  INVD0 U3171 ( .I(1'b1), .ZN(n[3165]) );
  INVD0 U3173 ( .I(1'b1), .ZN(n[3166]) );
  INVD0 U3175 ( .I(1'b1), .ZN(n[3169]) );
  INVD0 U3177 ( .I(1'b1), .ZN(n[3170]) );
  INVD0 U3179 ( .I(1'b1), .ZN(n[3172]) );
  INVD0 U3181 ( .I(1'b1), .ZN(n[3173]) );
  INVD0 U3183 ( .I(1'b1), .ZN(n[3177]) );
  INVD0 U3185 ( .I(1'b1), .ZN(n[3178]) );
  INVD0 U3187 ( .I(1'b1), .ZN(n[3180]) );
  INVD0 U3189 ( .I(1'b1), .ZN(n[3181]) );
  INVD0 U3191 ( .I(1'b1), .ZN(n[3184]) );
  INVD0 U3193 ( .I(1'b1), .ZN(n[3185]) );
  INVD0 U3195 ( .I(1'b1), .ZN(n[3187]) );
  INVD0 U3197 ( .I(1'b1), .ZN(n[3188]) );
  INVD0 U3199 ( .I(1'b1), .ZN(n[3195]) );
  INVD0 U3201 ( .I(1'b1), .ZN(n[3196]) );
  INVD0 U3203 ( .I(1'b1), .ZN(n[3198]) );
  INVD0 U3205 ( .I(1'b1), .ZN(n[3199]) );
  INVD0 U3207 ( .I(1'b1), .ZN(n[3202]) );
  INVD0 U3209 ( .I(1'b1), .ZN(n[3203]) );
  INVD0 U3211 ( .I(1'b1), .ZN(n[3205]) );
  INVD0 U3213 ( .I(1'b1), .ZN(n[3206]) );
  INVD0 U3215 ( .I(1'b1), .ZN(n[3210]) );
  INVD0 U3217 ( .I(1'b1), .ZN(n[3211]) );
  INVD0 U3219 ( .I(1'b1), .ZN(n[3213]) );
  INVD0 U3221 ( .I(1'b1), .ZN(n[3214]) );
  INVD0 U3223 ( .I(1'b1), .ZN(n[3217]) );
  INVD0 U3225 ( .I(1'b1), .ZN(n[3218]) );
  INVD0 U3227 ( .I(1'b1), .ZN(n[3220]) );
  INVD0 U3229 ( .I(1'b1), .ZN(n[3221]) );
  INVD0 U3231 ( .I(1'b1), .ZN(n[3226]) );
  INVD0 U3233 ( .I(1'b1), .ZN(n[3227]) );
  INVD0 U3235 ( .I(1'b1), .ZN(n[3229]) );
  INVD0 U3237 ( .I(1'b1), .ZN(n[3230]) );
  INVD0 U3239 ( .I(1'b1), .ZN(n[3233]) );
  INVD0 U3241 ( .I(1'b1), .ZN(n[3234]) );
  INVD0 U3243 ( .I(1'b1), .ZN(n[3236]) );
  INVD0 U3245 ( .I(1'b1), .ZN(n[3237]) );
  INVD0 U3247 ( .I(1'b1), .ZN(n[3241]) );
  INVD0 U3249 ( .I(1'b1), .ZN(n[3242]) );
  INVD0 U3251 ( .I(1'b1), .ZN(n[3244]) );
  INVD0 U3253 ( .I(1'b1), .ZN(n[3245]) );
  INVD0 U3255 ( .I(1'b1), .ZN(n[3248]) );
  INVD0 U3257 ( .I(1'b1), .ZN(n[3249]) );
  INVD0 U3259 ( .I(1'b1), .ZN(n[3251]) );
  INVD0 U3261 ( .I(1'b1), .ZN(n[3252]) );
  INVD0 U3263 ( .I(1'b1), .ZN(n[3258]) );
  INVD0 U3265 ( .I(1'b1), .ZN(n[3259]) );
  INVD0 U3267 ( .I(1'b1), .ZN(n[3261]) );
  INVD0 U3269 ( .I(1'b1), .ZN(n[3262]) );
  INVD0 U3271 ( .I(1'b1), .ZN(n[3265]) );
  INVD0 U3273 ( .I(1'b1), .ZN(n[3266]) );
  INVD0 U3275 ( .I(1'b1), .ZN(n[3268]) );
  INVD0 U3277 ( .I(1'b1), .ZN(n[3269]) );
  INVD0 U3279 ( .I(1'b1), .ZN(n[3273]) );
  INVD0 U3281 ( .I(1'b1), .ZN(n[3274]) );
  INVD0 U3283 ( .I(1'b1), .ZN(n[3276]) );
  INVD0 U3285 ( .I(1'b1), .ZN(n[3277]) );
  INVD0 U3287 ( .I(1'b1), .ZN(n[3280]) );
  INVD0 U3289 ( .I(1'b1), .ZN(n[3281]) );
  INVD0 U3291 ( .I(1'b1), .ZN(n[3283]) );
  INVD0 U3293 ( .I(1'b1), .ZN(n[3284]) );
  INVD0 U3295 ( .I(1'b1), .ZN(n[3289]) );
  INVD0 U3297 ( .I(1'b1), .ZN(n[3290]) );
  INVD0 U3299 ( .I(1'b1), .ZN(n[3292]) );
  INVD0 U3301 ( .I(1'b1), .ZN(n[3293]) );
  INVD0 U3303 ( .I(1'b1), .ZN(n[3296]) );
  INVD0 U3305 ( .I(1'b1), .ZN(n[3297]) );
  INVD0 U3307 ( .I(1'b1), .ZN(n[3299]) );
  INVD0 U3309 ( .I(1'b1), .ZN(n[3300]) );
  INVD0 U3311 ( .I(1'b1), .ZN(n[3304]) );
  INVD0 U3313 ( .I(1'b1), .ZN(n[3305]) );
  INVD0 U3315 ( .I(1'b1), .ZN(n[3307]) );
  INVD0 U3317 ( .I(1'b1), .ZN(n[3308]) );
  INVD0 U3319 ( .I(1'b1), .ZN(n[3311]) );
  INVD0 U3321 ( .I(1'b1), .ZN(n[3312]) );
  INVD0 U3323 ( .I(1'b1), .ZN(n[3314]) );
  INVD0 U3325 ( .I(1'b1), .ZN(n[3315]) );
  INVD0 U3327 ( .I(1'b1), .ZN(n[3323]) );
  INVD0 U3329 ( .I(1'b1), .ZN(n[3324]) );
  INVD0 U3331 ( .I(1'b1), .ZN(n[3326]) );
  INVD0 U3333 ( .I(1'b1), .ZN(n[3327]) );
  INVD0 U3335 ( .I(1'b1), .ZN(n[3330]) );
  INVD0 U3337 ( .I(1'b1), .ZN(n[3331]) );
  INVD0 U3339 ( .I(1'b1), .ZN(n[3333]) );
  INVD0 U3341 ( .I(1'b1), .ZN(n[3334]) );
  INVD0 U3343 ( .I(1'b1), .ZN(n[3338]) );
  INVD0 U3345 ( .I(1'b1), .ZN(n[3339]) );
  INVD0 U3347 ( .I(1'b1), .ZN(n[3341]) );
  INVD0 U3349 ( .I(1'b1), .ZN(n[3342]) );
  INVD0 U3351 ( .I(1'b1), .ZN(n[3345]) );
  INVD0 U3353 ( .I(1'b1), .ZN(n[3346]) );
  INVD0 U3355 ( .I(1'b1), .ZN(n[3348]) );
  INVD0 U3357 ( .I(1'b1), .ZN(n[3349]) );
  INVD0 U3359 ( .I(1'b1), .ZN(n[3354]) );
  INVD0 U3361 ( .I(1'b1), .ZN(n[3355]) );
  INVD0 U3363 ( .I(1'b1), .ZN(n[3357]) );
  INVD0 U3365 ( .I(1'b1), .ZN(n[3358]) );
  INVD0 U3367 ( .I(1'b1), .ZN(n[3361]) );
  INVD0 U3369 ( .I(1'b1), .ZN(n[3362]) );
  INVD0 U3371 ( .I(1'b1), .ZN(n[3364]) );
  INVD0 U3373 ( .I(1'b1), .ZN(n[3365]) );
  INVD0 U3375 ( .I(1'b1), .ZN(n[3369]) );
  INVD0 U3377 ( .I(1'b1), .ZN(n[3370]) );
  INVD0 U3379 ( .I(1'b1), .ZN(n[3372]) );
  INVD0 U3381 ( .I(1'b1), .ZN(n[3373]) );
  INVD0 U3383 ( .I(1'b1), .ZN(n[3376]) );
  INVD0 U3385 ( .I(1'b1), .ZN(n[3377]) );
  INVD0 U3387 ( .I(1'b1), .ZN(n[3379]) );
  INVD0 U3389 ( .I(1'b1), .ZN(n[3380]) );
  INVD0 U3391 ( .I(1'b1), .ZN(n[3386]) );
  INVD0 U3393 ( .I(1'b1), .ZN(n[3387]) );
  INVD0 U3395 ( .I(1'b1), .ZN(n[3389]) );
  INVD0 U3397 ( .I(1'b1), .ZN(n[3390]) );
  INVD0 U3399 ( .I(1'b1), .ZN(n[3393]) );
  INVD0 U3401 ( .I(1'b1), .ZN(n[3394]) );
  INVD0 U3403 ( .I(1'b1), .ZN(n[3396]) );
  INVD0 U3405 ( .I(1'b1), .ZN(n[3397]) );
  INVD0 U3407 ( .I(1'b1), .ZN(n[3401]) );
  INVD0 U3409 ( .I(1'b1), .ZN(n[3402]) );
  INVD0 U3411 ( .I(1'b1), .ZN(n[3404]) );
  INVD0 U3413 ( .I(1'b1), .ZN(n[3405]) );
  INVD0 U3415 ( .I(1'b1), .ZN(n[3408]) );
  INVD0 U3417 ( .I(1'b1), .ZN(n[3409]) );
  INVD0 U3419 ( .I(1'b1), .ZN(n[3411]) );
  INVD0 U3421 ( .I(1'b1), .ZN(n[3412]) );
  INVD0 U3423 ( .I(1'b1), .ZN(n[3417]) );
  INVD0 U3425 ( .I(1'b1), .ZN(n[3418]) );
  INVD0 U3427 ( .I(1'b1), .ZN(n[3420]) );
  INVD0 U3429 ( .I(1'b1), .ZN(n[3421]) );
  INVD0 U3431 ( .I(1'b1), .ZN(n[3424]) );
  INVD0 U3433 ( .I(1'b1), .ZN(n[3425]) );
  INVD0 U3435 ( .I(1'b1), .ZN(n[3427]) );
  INVD0 U3437 ( .I(1'b1), .ZN(n[3428]) );
  INVD0 U3439 ( .I(1'b1), .ZN(n[3432]) );
  INVD0 U3441 ( .I(1'b1), .ZN(n[3433]) );
  INVD0 U3443 ( .I(1'b1), .ZN(n[3435]) );
  INVD0 U3445 ( .I(1'b1), .ZN(n[3436]) );
  INVD0 U3447 ( .I(1'b1), .ZN(n[3439]) );
  INVD0 U3449 ( .I(1'b1), .ZN(n[3440]) );
  INVD0 U3451 ( .I(1'b1), .ZN(n[3442]) );
  INVD0 U3453 ( .I(1'b1), .ZN(n[3443]) );
  INVD0 U3455 ( .I(1'b1), .ZN(n[3450]) );
  INVD0 U3457 ( .I(1'b1), .ZN(n[3451]) );
  INVD0 U3459 ( .I(1'b1), .ZN(n[3453]) );
  INVD0 U3461 ( .I(1'b1), .ZN(n[3454]) );
  INVD0 U3463 ( .I(1'b1), .ZN(n[3457]) );
  INVD0 U3465 ( .I(1'b1), .ZN(n[3458]) );
  INVD0 U3467 ( .I(1'b1), .ZN(n[3460]) );
  INVD0 U3469 ( .I(1'b1), .ZN(n[3461]) );
  INVD0 U3471 ( .I(1'b1), .ZN(n[3465]) );
  INVD0 U3473 ( .I(1'b1), .ZN(n[3466]) );
  INVD0 U3475 ( .I(1'b1), .ZN(n[3468]) );
  INVD0 U3477 ( .I(1'b1), .ZN(n[3469]) );
  INVD0 U3479 ( .I(1'b1), .ZN(n[3472]) );
  INVD0 U3481 ( .I(1'b1), .ZN(n[3473]) );
  INVD0 U3483 ( .I(1'b1), .ZN(n[3475]) );
  INVD0 U3485 ( .I(1'b1), .ZN(n[3476]) );
  INVD0 U3487 ( .I(1'b1), .ZN(n[3481]) );
  INVD0 U3489 ( .I(1'b1), .ZN(n[3482]) );
  INVD0 U3491 ( .I(1'b1), .ZN(n[3484]) );
  INVD0 U3493 ( .I(1'b1), .ZN(n[3485]) );
  INVD0 U3495 ( .I(1'b1), .ZN(n[3488]) );
  INVD0 U3497 ( .I(1'b1), .ZN(n[3489]) );
  INVD0 U3499 ( .I(1'b1), .ZN(n[3491]) );
  INVD0 U3501 ( .I(1'b1), .ZN(n[3492]) );
  INVD0 U3503 ( .I(1'b1), .ZN(n[3496]) );
  INVD0 U3505 ( .I(1'b1), .ZN(n[3497]) );
  INVD0 U3507 ( .I(1'b1), .ZN(n[3499]) );
  INVD0 U3509 ( .I(1'b1), .ZN(n[3500]) );
  INVD0 U3511 ( .I(1'b1), .ZN(n[3503]) );
  INVD0 U3513 ( .I(1'b1), .ZN(n[3504]) );
  INVD0 U3515 ( .I(1'b1), .ZN(n[3506]) );
  INVD0 U3517 ( .I(1'b1), .ZN(n[3507]) );
  INVD0 U3519 ( .I(1'b1), .ZN(n[3513]) );
  INVD0 U3521 ( .I(1'b1), .ZN(n[3514]) );
  INVD0 U3523 ( .I(1'b1), .ZN(n[3516]) );
  INVD0 U3525 ( .I(1'b1), .ZN(n[3517]) );
  INVD0 U3527 ( .I(1'b1), .ZN(n[3520]) );
  INVD0 U3529 ( .I(1'b1), .ZN(n[3521]) );
  INVD0 U3531 ( .I(1'b1), .ZN(n[3523]) );
  INVD0 U3533 ( .I(1'b1), .ZN(n[3524]) );
  INVD0 U3535 ( .I(1'b1), .ZN(n[3528]) );
  INVD0 U3537 ( .I(1'b1), .ZN(n[3529]) );
  INVD0 U3539 ( .I(1'b1), .ZN(n[3531]) );
  INVD0 U3541 ( .I(1'b1), .ZN(n[3532]) );
  INVD0 U3543 ( .I(1'b1), .ZN(n[3535]) );
  INVD0 U3545 ( .I(1'b1), .ZN(n[3536]) );
  INVD0 U3547 ( .I(1'b1), .ZN(n[3538]) );
  INVD0 U3549 ( .I(1'b1), .ZN(n[3539]) );
  INVD0 U3551 ( .I(1'b1), .ZN(n[3544]) );
  INVD0 U3553 ( .I(1'b1), .ZN(n[3545]) );
  INVD0 U3555 ( .I(1'b1), .ZN(n[3547]) );
  INVD0 U3557 ( .I(1'b1), .ZN(n[3548]) );
  INVD0 U3559 ( .I(1'b1), .ZN(n[3551]) );
  INVD0 U3561 ( .I(1'b1), .ZN(n[3552]) );
  INVD0 U3563 ( .I(1'b1), .ZN(n[3554]) );
  INVD0 U3565 ( .I(1'b1), .ZN(n[3555]) );
  INVD0 U3567 ( .I(1'b1), .ZN(n[3559]) );
  INVD0 U3569 ( .I(1'b1), .ZN(n[3560]) );
  INVD0 U3571 ( .I(1'b1), .ZN(n[3562]) );
  INVD0 U3573 ( .I(1'b1), .ZN(n[3563]) );
  INVD0 U3575 ( .I(1'b1), .ZN(n[3566]) );
  INVD0 U3577 ( .I(1'b1), .ZN(n[3567]) );
  INVD0 U3579 ( .I(1'b1), .ZN(n[3569]) );
  INVD0 U3581 ( .I(1'b1), .ZN(n[3570]) );
  INVD0 U3583 ( .I(1'b1), .ZN(n[3579]) );
  INVD0 U3585 ( .I(1'b1), .ZN(n[3580]) );
  INVD0 U3587 ( .I(1'b1), .ZN(n[3582]) );
  INVD0 U3589 ( .I(1'b1), .ZN(n[3583]) );
  INVD0 U3591 ( .I(1'b1), .ZN(n[3586]) );
  INVD0 U3593 ( .I(1'b1), .ZN(n[3587]) );
  INVD0 U3595 ( .I(1'b1), .ZN(n[3589]) );
  INVD0 U3597 ( .I(1'b1), .ZN(n[3590]) );
  INVD0 U3599 ( .I(1'b1), .ZN(n[3594]) );
  INVD0 U3601 ( .I(1'b1), .ZN(n[3595]) );
  INVD0 U3603 ( .I(1'b1), .ZN(n[3597]) );
  INVD0 U3605 ( .I(1'b1), .ZN(n[3598]) );
  INVD0 U3607 ( .I(1'b1), .ZN(n[3601]) );
  INVD0 U3609 ( .I(1'b1), .ZN(n[3602]) );
  INVD0 U3611 ( .I(1'b1), .ZN(n[3604]) );
  INVD0 U3613 ( .I(1'b1), .ZN(n[3605]) );
  INVD0 U3615 ( .I(1'b1), .ZN(n[3610]) );
  INVD0 U3617 ( .I(1'b1), .ZN(n[3611]) );
  INVD0 U3619 ( .I(1'b1), .ZN(n[3613]) );
  INVD0 U3621 ( .I(1'b1), .ZN(n[3614]) );
  INVD0 U3623 ( .I(1'b1), .ZN(n[3617]) );
  INVD0 U3625 ( .I(1'b1), .ZN(n[3618]) );
  INVD0 U3627 ( .I(1'b1), .ZN(n[3620]) );
  INVD0 U3629 ( .I(1'b1), .ZN(n[3621]) );
  INVD0 U3631 ( .I(1'b1), .ZN(n[3625]) );
  INVD0 U3633 ( .I(1'b1), .ZN(n[3626]) );
  INVD0 U3635 ( .I(1'b1), .ZN(n[3628]) );
  INVD0 U3637 ( .I(1'b1), .ZN(n[3629]) );
  INVD0 U3639 ( .I(1'b1), .ZN(n[3632]) );
  INVD0 U3641 ( .I(1'b1), .ZN(n[3633]) );
  INVD0 U3643 ( .I(1'b1), .ZN(n[3635]) );
  INVD0 U3645 ( .I(1'b1), .ZN(n[3636]) );
  INVD0 U3647 ( .I(1'b1), .ZN(n[3642]) );
  INVD0 U3649 ( .I(1'b1), .ZN(n[3643]) );
  INVD0 U3651 ( .I(1'b1), .ZN(n[3645]) );
  INVD0 U3653 ( .I(1'b1), .ZN(n[3646]) );
  INVD0 U3655 ( .I(1'b1), .ZN(n[3649]) );
  INVD0 U3657 ( .I(1'b1), .ZN(n[3650]) );
  INVD0 U3659 ( .I(1'b1), .ZN(n[3652]) );
  INVD0 U3661 ( .I(1'b1), .ZN(n[3653]) );
  INVD0 U3663 ( .I(1'b1), .ZN(n[3657]) );
  INVD0 U3665 ( .I(1'b1), .ZN(n[3658]) );
  INVD0 U3667 ( .I(1'b1), .ZN(n[3660]) );
  INVD0 U3669 ( .I(1'b1), .ZN(n[3661]) );
  INVD0 U3671 ( .I(1'b1), .ZN(n[3664]) );
  INVD0 U3673 ( .I(1'b1), .ZN(n[3665]) );
  INVD0 U3675 ( .I(1'b1), .ZN(n[3667]) );
  INVD0 U3677 ( .I(1'b1), .ZN(n[3668]) );
  INVD0 U3679 ( .I(1'b1), .ZN(n[3673]) );
  INVD0 U3681 ( .I(1'b1), .ZN(n[3674]) );
  INVD0 U3683 ( .I(1'b1), .ZN(n[3676]) );
  INVD0 U3685 ( .I(1'b1), .ZN(n[3677]) );
  INVD0 U3687 ( .I(1'b1), .ZN(n[3680]) );
  INVD0 U3689 ( .I(1'b1), .ZN(n[3681]) );
  INVD0 U3691 ( .I(1'b1), .ZN(n[3683]) );
  INVD0 U3693 ( .I(1'b1), .ZN(n[3684]) );
  INVD0 U3695 ( .I(1'b1), .ZN(n[3688]) );
  INVD0 U3697 ( .I(1'b1), .ZN(n[3689]) );
  INVD0 U3699 ( .I(1'b1), .ZN(n[3691]) );
  INVD0 U3701 ( .I(1'b1), .ZN(n[3692]) );
  INVD0 U3703 ( .I(1'b1), .ZN(n[3695]) );
  INVD0 U3705 ( .I(1'b1), .ZN(n[3696]) );
  INVD0 U3707 ( .I(1'b1), .ZN(n[3698]) );
  INVD0 U3709 ( .I(1'b1), .ZN(n[3699]) );
  INVD0 U3711 ( .I(1'b1), .ZN(n[3706]) );
  INVD0 U3713 ( .I(1'b1), .ZN(n[3707]) );
  INVD0 U3715 ( .I(1'b1), .ZN(n[3709]) );
  INVD0 U3717 ( .I(1'b1), .ZN(n[3710]) );
  INVD0 U3719 ( .I(1'b1), .ZN(n[3713]) );
  INVD0 U3721 ( .I(1'b1), .ZN(n[3714]) );
  INVD0 U3723 ( .I(1'b1), .ZN(n[3716]) );
  INVD0 U3725 ( .I(1'b1), .ZN(n[3717]) );
  INVD0 U3727 ( .I(1'b1), .ZN(n[3721]) );
  INVD0 U3729 ( .I(1'b1), .ZN(n[3722]) );
  INVD0 U3731 ( .I(1'b1), .ZN(n[3724]) );
  INVD0 U3733 ( .I(1'b1), .ZN(n[3725]) );
  INVD0 U3735 ( .I(1'b1), .ZN(n[3728]) );
  INVD0 U3737 ( .I(1'b1), .ZN(n[3729]) );
  INVD0 U3739 ( .I(1'b1), .ZN(n[3731]) );
  INVD0 U3741 ( .I(1'b1), .ZN(n[3732]) );
  INVD0 U3743 ( .I(1'b1), .ZN(n[3737]) );
  INVD0 U3745 ( .I(1'b1), .ZN(n[3738]) );
  INVD0 U3747 ( .I(1'b1), .ZN(n[3740]) );
  INVD0 U3749 ( .I(1'b1), .ZN(n[3741]) );
  INVD0 U3751 ( .I(1'b1), .ZN(n[3744]) );
  INVD0 U3753 ( .I(1'b1), .ZN(n[3745]) );
  INVD0 U3755 ( .I(1'b1), .ZN(n[3747]) );
  INVD0 U3757 ( .I(1'b1), .ZN(n[3748]) );
  INVD0 U3759 ( .I(1'b1), .ZN(n[3752]) );
  INVD0 U3761 ( .I(1'b1), .ZN(n[3753]) );
  INVD0 U3763 ( .I(1'b1), .ZN(n[3755]) );
  INVD0 U3765 ( .I(1'b1), .ZN(n[3756]) );
  INVD0 U3767 ( .I(1'b1), .ZN(n[3759]) );
  INVD0 U3769 ( .I(1'b1), .ZN(n[3760]) );
  INVD0 U3771 ( .I(1'b1), .ZN(n[3762]) );
  INVD0 U3773 ( .I(1'b1), .ZN(n[3763]) );
  INVD0 U3775 ( .I(1'b1), .ZN(n[3769]) );
  INVD0 U3777 ( .I(1'b1), .ZN(n[3770]) );
  INVD0 U3779 ( .I(1'b1), .ZN(n[3772]) );
  INVD0 U3781 ( .I(1'b1), .ZN(n[3773]) );
  INVD0 U3783 ( .I(1'b1), .ZN(n[3776]) );
  INVD0 U3785 ( .I(1'b1), .ZN(n[3777]) );
  INVD0 U3787 ( .I(1'b1), .ZN(n[3779]) );
  INVD0 U3789 ( .I(1'b1), .ZN(n[3780]) );
  INVD0 U3791 ( .I(1'b1), .ZN(n[3784]) );
  INVD0 U3793 ( .I(1'b1), .ZN(n[3785]) );
  INVD0 U3795 ( .I(1'b1), .ZN(n[3787]) );
  INVD0 U3797 ( .I(1'b1), .ZN(n[3788]) );
  INVD0 U3799 ( .I(1'b1), .ZN(n[3791]) );
  INVD0 U3801 ( .I(1'b1), .ZN(n[3792]) );
  INVD0 U3803 ( .I(1'b1), .ZN(n[3794]) );
  INVD0 U3805 ( .I(1'b1), .ZN(n[3795]) );
  INVD0 U3807 ( .I(1'b1), .ZN(n[3800]) );
  INVD0 U3809 ( .I(1'b1), .ZN(n[3801]) );
  INVD0 U3811 ( .I(1'b1), .ZN(n[3803]) );
  INVD0 U3813 ( .I(1'b1), .ZN(n[3804]) );
  INVD0 U3815 ( .I(1'b1), .ZN(n[3807]) );
  INVD0 U3817 ( .I(1'b1), .ZN(n[3808]) );
  INVD0 U3819 ( .I(1'b1), .ZN(n[3810]) );
  INVD0 U3821 ( .I(1'b1), .ZN(n[3811]) );
  INVD0 U3823 ( .I(1'b1), .ZN(n[3815]) );
  INVD0 U3825 ( .I(1'b1), .ZN(n[3816]) );
  INVD0 U3827 ( .I(1'b1), .ZN(n[3818]) );
  INVD0 U3829 ( .I(1'b1), .ZN(n[3819]) );
  INVD0 U3831 ( .I(1'b1), .ZN(n[3822]) );
  INVD0 U3833 ( .I(1'b1), .ZN(n[3823]) );
  INVD0 U3835 ( .I(1'b1), .ZN(n[3825]) );
  INVD0 U3837 ( .I(1'b1), .ZN(n[3826]) );
  INVD0 U3839 ( .I(1'b1), .ZN(n[3834]) );
  INVD0 U3841 ( .I(1'b1), .ZN(n[3835]) );
  INVD0 U3843 ( .I(1'b1), .ZN(n[3837]) );
  INVD0 U3845 ( .I(1'b1), .ZN(n[3838]) );
  INVD0 U3847 ( .I(1'b1), .ZN(n[3841]) );
  INVD0 U3849 ( .I(1'b1), .ZN(n[3842]) );
  INVD0 U3851 ( .I(1'b1), .ZN(n[3844]) );
  INVD0 U3853 ( .I(1'b1), .ZN(n[3845]) );
  INVD0 U3855 ( .I(1'b1), .ZN(n[3849]) );
  INVD0 U3857 ( .I(1'b1), .ZN(n[3850]) );
  INVD0 U3859 ( .I(1'b1), .ZN(n[3852]) );
  INVD0 U3861 ( .I(1'b1), .ZN(n[3853]) );
  INVD0 U3863 ( .I(1'b1), .ZN(n[3856]) );
  INVD0 U3865 ( .I(1'b1), .ZN(n[3857]) );
  INVD0 U3867 ( .I(1'b1), .ZN(n[3859]) );
  INVD0 U3869 ( .I(1'b1), .ZN(n[3860]) );
  INVD0 U3871 ( .I(1'b1), .ZN(n[3865]) );
  INVD0 U3873 ( .I(1'b1), .ZN(n[3866]) );
  INVD0 U3875 ( .I(1'b1), .ZN(n[3868]) );
  INVD0 U3877 ( .I(1'b1), .ZN(n[3869]) );
  INVD0 U3879 ( .I(1'b1), .ZN(n[3872]) );
  INVD0 U3881 ( .I(1'b1), .ZN(n[3873]) );
  INVD0 U3883 ( .I(1'b1), .ZN(n[3875]) );
  INVD0 U3885 ( .I(1'b1), .ZN(n[3876]) );
  INVD0 U3887 ( .I(1'b1), .ZN(n[3880]) );
  INVD0 U3889 ( .I(1'b1), .ZN(n[3881]) );
  INVD0 U3891 ( .I(1'b1), .ZN(n[3883]) );
  INVD0 U3893 ( .I(1'b1), .ZN(n[3884]) );
  INVD0 U3895 ( .I(1'b1), .ZN(n[3887]) );
  INVD0 U3897 ( .I(1'b1), .ZN(n[3888]) );
  INVD0 U3899 ( .I(1'b1), .ZN(n[3890]) );
  INVD0 U3901 ( .I(1'b1), .ZN(n[3891]) );
  INVD0 U3903 ( .I(1'b1), .ZN(n[3897]) );
  INVD0 U3905 ( .I(1'b1), .ZN(n[3898]) );
  INVD0 U3907 ( .I(1'b1), .ZN(n[3900]) );
  INVD0 U3909 ( .I(1'b1), .ZN(n[3901]) );
  INVD0 U3911 ( .I(1'b1), .ZN(n[3904]) );
  INVD0 U3913 ( .I(1'b1), .ZN(n[3905]) );
  INVD0 U3915 ( .I(1'b1), .ZN(n[3907]) );
  INVD0 U3917 ( .I(1'b1), .ZN(n[3908]) );
  INVD0 U3919 ( .I(1'b1), .ZN(n[3912]) );
  INVD0 U3921 ( .I(1'b1), .ZN(n[3913]) );
  INVD0 U3923 ( .I(1'b1), .ZN(n[3915]) );
  INVD0 U3925 ( .I(1'b1), .ZN(n[3916]) );
  INVD0 U3927 ( .I(1'b1), .ZN(n[3919]) );
  INVD0 U3929 ( .I(1'b1), .ZN(n[3920]) );
  INVD0 U3931 ( .I(1'b1), .ZN(n[3922]) );
  INVD0 U3933 ( .I(1'b1), .ZN(n[3923]) );
  INVD0 U3935 ( .I(1'b1), .ZN(n[3928]) );
  INVD0 U3937 ( .I(1'b1), .ZN(n[3929]) );
  INVD0 U3939 ( .I(1'b1), .ZN(n[3931]) );
  INVD0 U3941 ( .I(1'b1), .ZN(n[3932]) );
  INVD0 U3943 ( .I(1'b1), .ZN(n[3935]) );
  INVD0 U3945 ( .I(1'b1), .ZN(n[3936]) );
  INVD0 U3947 ( .I(1'b1), .ZN(n[3938]) );
  INVD0 U3949 ( .I(1'b1), .ZN(n[3939]) );
  INVD0 U3951 ( .I(1'b1), .ZN(n[3943]) );
  INVD0 U3953 ( .I(1'b1), .ZN(n[3944]) );
  INVD0 U3955 ( .I(1'b1), .ZN(n[3946]) );
  INVD0 U3957 ( .I(1'b1), .ZN(n[3947]) );
  INVD0 U3959 ( .I(1'b1), .ZN(n[3950]) );
  INVD0 U3961 ( .I(1'b1), .ZN(n[3951]) );
  INVD0 U3963 ( .I(1'b1), .ZN(n[3953]) );
  INVD0 U3965 ( .I(1'b1), .ZN(n[3954]) );
  INVD0 U3967 ( .I(1'b1), .ZN(n[3961]) );
  INVD0 U3969 ( .I(1'b1), .ZN(n[3962]) );
  INVD0 U3971 ( .I(1'b1), .ZN(n[3964]) );
  INVD0 U3973 ( .I(1'b1), .ZN(n[3965]) );
  INVD0 U3975 ( .I(1'b1), .ZN(n[3968]) );
  INVD0 U3977 ( .I(1'b1), .ZN(n[3969]) );
  INVD0 U3979 ( .I(1'b1), .ZN(n[3971]) );
  INVD0 U3981 ( .I(1'b1), .ZN(n[3972]) );
  INVD0 U3983 ( .I(1'b1), .ZN(n[3976]) );
  INVD0 U3985 ( .I(1'b1), .ZN(n[3977]) );
  INVD0 U3987 ( .I(1'b1), .ZN(n[3979]) );
  INVD0 U3989 ( .I(1'b1), .ZN(n[3980]) );
  INVD0 U3991 ( .I(1'b1), .ZN(n[3983]) );
  INVD0 U3993 ( .I(1'b1), .ZN(n[3984]) );
  INVD0 U3995 ( .I(1'b1), .ZN(n[3986]) );
  INVD0 U3997 ( .I(1'b1), .ZN(n[3987]) );
  INVD0 U3999 ( .I(1'b1), .ZN(n[3992]) );
  INVD0 U4001 ( .I(1'b1), .ZN(n[3993]) );
  INVD0 U4003 ( .I(1'b1), .ZN(n[3995]) );
  INVD0 U4005 ( .I(1'b1), .ZN(n[3996]) );
  INVD0 U4007 ( .I(1'b1), .ZN(n[3999]) );
  INVD0 U4009 ( .I(1'b1), .ZN(n[4000]) );
  INVD0 U4011 ( .I(1'b1), .ZN(n[4002]) );
  INVD0 U4013 ( .I(1'b1), .ZN(n[4003]) );
  INVD0 U4015 ( .I(1'b1), .ZN(n[4007]) );
  INVD0 U4017 ( .I(1'b1), .ZN(n[4008]) );
  INVD0 U4019 ( .I(1'b1), .ZN(n[4010]) );
  INVD0 U4021 ( .I(1'b1), .ZN(n[4011]) );
  INVD0 U4023 ( .I(1'b1), .ZN(n[4014]) );
  INVD0 U4025 ( .I(1'b1), .ZN(n[4015]) );
  INVD0 U4027 ( .I(1'b1), .ZN(n[4017]) );
  INVD0 U4029 ( .I(1'b1), .ZN(n[4018]) );
  INVD0 U4031 ( .I(1'b1), .ZN(n[4024]) );
  INVD0 U4033 ( .I(1'b1), .ZN(n[4025]) );
  INVD0 U4035 ( .I(1'b1), .ZN(n[4027]) );
  INVD0 U4037 ( .I(1'b1), .ZN(n[4028]) );
  INVD0 U4039 ( .I(1'b1), .ZN(n[4031]) );
  INVD0 U4041 ( .I(1'b1), .ZN(n[4032]) );
  INVD0 U4043 ( .I(1'b1), .ZN(n[4034]) );
  INVD0 U4045 ( .I(1'b1), .ZN(n[4035]) );
  INVD0 U4047 ( .I(1'b1), .ZN(n[4039]) );
  INVD0 U4049 ( .I(1'b1), .ZN(n[4040]) );
  INVD0 U4051 ( .I(1'b1), .ZN(n[4042]) );
  INVD0 U4053 ( .I(1'b1), .ZN(n[4043]) );
  INVD0 U4055 ( .I(1'b1), .ZN(n[4046]) );
  INVD0 U4057 ( .I(1'b1), .ZN(n[4047]) );
  INVD0 U4059 ( .I(1'b1), .ZN(n[4049]) );
  INVD0 U4061 ( .I(1'b1), .ZN(n[4050]) );
  INVD0 U4063 ( .I(1'b1), .ZN(n[4055]) );
  INVD0 U4065 ( .I(1'b1), .ZN(n[4056]) );
  INVD0 U4067 ( .I(1'b1), .ZN(n[4058]) );
  INVD0 U4069 ( .I(1'b1), .ZN(n[4059]) );
  INVD0 U4071 ( .I(1'b1), .ZN(n[4062]) );
  INVD0 U4073 ( .I(1'b1), .ZN(n[4063]) );
  INVD0 U4075 ( .I(1'b1), .ZN(n[4065]) );
  INVD0 U4077 ( .I(1'b1), .ZN(n[4066]) );
  INVD0 U4079 ( .I(1'b1), .ZN(n[4070]) );
  INVD0 U4081 ( .I(1'b1), .ZN(n[4071]) );
  INVD0 U4083 ( .I(1'b1), .ZN(n[4073]) );
  INVD0 U4085 ( .I(1'b1), .ZN(n[4074]) );
  INVD0 U4087 ( .I(1'b1), .ZN(n[4077]) );
  INVD0 U4089 ( .I(1'b1), .ZN(n[4078]) );
  INVD0 U4091 ( .I(1'b1), .ZN(n[4080]) );
  INVD0 U4093 ( .I(1'b1), .ZN(n[4081]) );
  AN2D0 U4095 ( .A1(b[9]), .A2(n[2032]), .Z(n[4079]) );
  AN2D0 U4096 ( .A1(n[2029]), .A2(b[9]), .Z(n[4076]) );
  AN2D0 U4097 ( .A1(n[2028]), .A2(b[9]), .Z(n[4075]) );
  AN2D0 U4098 ( .A1(n[2025]), .A2(b[9]), .Z(n[4072]) );
  AN2D0 U4099 ( .A1(n[2022]), .A2(b[9]), .Z(n[4069]) );
  AN2D0 U4100 ( .A1(n[2021]), .A2(b[9]), .Z(n[4068]) );
  AN2D0 U4101 ( .A1(n[2020]), .A2(b[9]), .Z(n[4067]) );
  AN2D0 U4102 ( .A1(n[2017]), .A2(b[9]), .Z(n[4064]) );
  AN2D0 U4103 ( .A1(n[2014]), .A2(b[9]), .Z(n[4061]) );
  AN2D0 U4104 ( .A1(n[2013]), .A2(b[9]), .Z(n[4060]) );
  AN2D0 U4105 ( .A1(n[2010]), .A2(b[9]), .Z(n[4057]) );
  AN2D0 U4106 ( .A1(n[2007]), .A2(b[9]), .Z(n[4054]) );
  AN2D0 U4107 ( .A1(n[2006]), .A2(b[9]), .Z(n[4053]) );
  AN2D0 U4108 ( .A1(n[2005]), .A2(b[9]), .Z(n[4052]) );
  AN2D0 U4109 ( .A1(n[2004]), .A2(b[9]), .Z(n[4051]) );
  AN2D0 U4110 ( .A1(n[2001]), .A2(b[9]), .Z(n[4048]) );
  AN2D0 U4111 ( .A1(n[1998]), .A2(b[9]), .Z(n[4045]) );
  AN2D0 U4112 ( .A1(n[1997]), .A2(b[9]), .Z(n[4044]) );
  AN2D0 U4113 ( .A1(n[1994]), .A2(b[9]), .Z(n[4041]) );
  AN2D0 U4114 ( .A1(n[1991]), .A2(b[9]), .Z(n[4038]) );
  AN2D0 U4115 ( .A1(n[1990]), .A2(b[9]), .Z(n[4037]) );
  AN2D0 U4116 ( .A1(n[1989]), .A2(b[9]), .Z(n[4036]) );
  AN2D0 U4117 ( .A1(n[1986]), .A2(b[9]), .Z(n[4033]) );
  AN2D0 U4118 ( .A1(n[1983]), .A2(b[9]), .Z(n[4030]) );
  AN2D0 U4119 ( .A1(n[1982]), .A2(b[9]), .Z(n[4029]) );
  AN2D0 U4120 ( .A1(n[1979]), .A2(b[9]), .Z(n[4026]) );
  AN2D0 U4121 ( .A1(n[1976]), .A2(b[9]), .Z(n[4023]) );
  AN2D0 U4122 ( .A1(n[1975]), .A2(b[9]), .Z(n[4022]) );
  AN2D0 U4123 ( .A1(n[1974]), .A2(b[9]), .Z(n[4021]) );
  AN2D0 U4124 ( .A1(n[1973]), .A2(b[9]), .Z(n[4020]) );
  AN2D0 U4125 ( .A1(n[1972]), .A2(b[9]), .Z(n[4019]) );
  AN2D0 U4126 ( .A1(n[1969]), .A2(b[9]), .Z(n[4016]) );
  AN2D0 U4127 ( .A1(n[1966]), .A2(b[9]), .Z(n[4013]) );
  AN2D0 U4128 ( .A1(n[1965]), .A2(b[9]), .Z(n[4012]) );
  AN2D0 U4129 ( .A1(n[1962]), .A2(b[9]), .Z(n[4009]) );
  AN2D0 U4130 ( .A1(n[1959]), .A2(b[9]), .Z(n[4006]) );
  AN2D0 U4131 ( .A1(n[1958]), .A2(b[9]), .Z(n[4005]) );
  AN2D0 U4132 ( .A1(n[1957]), .A2(b[9]), .Z(n[4004]) );
  AN2D0 U4133 ( .A1(n[1954]), .A2(b[9]), .Z(n[4001]) );
  AN2D0 U4134 ( .A1(n[1951]), .A2(b[9]), .Z(n[3998]) );
  AN2D0 U4135 ( .A1(n[1950]), .A2(b[9]), .Z(n[3997]) );
  AN2D0 U4136 ( .A1(n[1947]), .A2(b[9]), .Z(n[3994]) );
  AN2D0 U4137 ( .A1(n[1944]), .A2(b[9]), .Z(n[3991]) );
  AN2D0 U4138 ( .A1(n[1943]), .A2(b[9]), .Z(n[3990]) );
  AN2D0 U4139 ( .A1(n[1942]), .A2(b[9]), .Z(n[3989]) );
  AN2D0 U4140 ( .A1(n[1941]), .A2(b[9]), .Z(n[3988]) );
  AN2D0 U4141 ( .A1(n[1938]), .A2(b[9]), .Z(n[3985]) );
  AN2D0 U4142 ( .A1(n[1935]), .A2(b[9]), .Z(n[3982]) );
  AN2D0 U4143 ( .A1(n[1934]), .A2(b[9]), .Z(n[3981]) );
  AN2D0 U4144 ( .A1(n[1931]), .A2(b[9]), .Z(n[3978]) );
  AN2D0 U4145 ( .A1(n[1928]), .A2(b[9]), .Z(n[3975]) );
  AN2D0 U4146 ( .A1(n[1927]), .A2(b[9]), .Z(n[3974]) );
  AN2D0 U4147 ( .A1(n[1926]), .A2(b[9]), .Z(n[3973]) );
  AN2D0 U4148 ( .A1(n[1923]), .A2(b[9]), .Z(n[3970]) );
  AN2D0 U4149 ( .A1(n[1920]), .A2(b[9]), .Z(n[3967]) );
  AN2D0 U4150 ( .A1(n[1919]), .A2(b[9]), .Z(n[3966]) );
  AN2D0 U4151 ( .A1(n[1916]), .A2(b[9]), .Z(n[3963]) );
  AN2D0 U4152 ( .A1(n[1913]), .A2(b[9]), .Z(n[3960]) );
  AN2D0 U4153 ( .A1(n[1912]), .A2(b[9]), .Z(n[3959]) );
  AN2D0 U4154 ( .A1(n[1911]), .A2(b[9]), .Z(n[3958]) );
  AN2D0 U4155 ( .A1(n[1910]), .A2(b[9]), .Z(n[3957]) );
  AN2D0 U4156 ( .A1(n[1909]), .A2(b[9]), .Z(n[3956]) );
  AN2D0 U4157 ( .A1(n[1908]), .A2(b[9]), .Z(n[3955]) );
  AN2D0 U4158 ( .A1(n[1905]), .A2(b[9]), .Z(n[3952]) );
  AN2D0 U4159 ( .A1(n[1902]), .A2(b[9]), .Z(n[3949]) );
  AN2D0 U4160 ( .A1(n[1901]), .A2(b[9]), .Z(n[3948]) );
  AN2D0 U4161 ( .A1(n[1898]), .A2(b[9]), .Z(n[3945]) );
  AN2D0 U4162 ( .A1(n[1895]), .A2(b[9]), .Z(n[3942]) );
  AN2D0 U4163 ( .A1(n[1894]), .A2(b[9]), .Z(n[3941]) );
  AN2D0 U4164 ( .A1(n[1893]), .A2(b[9]), .Z(n[3940]) );
  AN2D0 U4165 ( .A1(n[1890]), .A2(b[9]), .Z(n[3937]) );
  AN2D0 U4166 ( .A1(n[1887]), .A2(b[9]), .Z(n[3934]) );
  AN2D0 U4167 ( .A1(n[1886]), .A2(b[9]), .Z(n[3933]) );
  AN2D0 U4168 ( .A1(n[1883]), .A2(b[9]), .Z(n[3930]) );
  AN2D0 U4169 ( .A1(n[1880]), .A2(b[9]), .Z(n[3927]) );
  AN2D0 U4170 ( .A1(n[1879]), .A2(b[9]), .Z(n[3926]) );
  AN2D0 U4171 ( .A1(n[1878]), .A2(b[9]), .Z(n[3925]) );
  AN2D0 U4172 ( .A1(n[1877]), .A2(b[9]), .Z(n[3924]) );
  AN2D0 U4173 ( .A1(n[1874]), .A2(b[9]), .Z(n[3921]) );
  AN2D0 U4174 ( .A1(n[1871]), .A2(b[9]), .Z(n[3918]) );
  AN2D0 U4175 ( .A1(n[1870]), .A2(b[9]), .Z(n[3917]) );
  AN2D0 U4176 ( .A1(n[1867]), .A2(b[9]), .Z(n[3914]) );
  AN2D0 U4177 ( .A1(n[1864]), .A2(b[9]), .Z(n[3911]) );
  AN2D0 U4178 ( .A1(n[1863]), .A2(b[9]), .Z(n[3910]) );
  AN2D0 U4179 ( .A1(n[1862]), .A2(b[9]), .Z(n[3909]) );
  AN2D0 U4180 ( .A1(n[1859]), .A2(b[9]), .Z(n[3906]) );
  AN2D0 U4181 ( .A1(n[1856]), .A2(b[9]), .Z(n[3903]) );
  AN2D0 U4182 ( .A1(n[1855]), .A2(b[9]), .Z(n[3902]) );
  AN2D0 U4183 ( .A1(n[1852]), .A2(b[9]), .Z(n[3899]) );
  AN2D0 U4184 ( .A1(n[1849]), .A2(b[9]), .Z(n[3896]) );
  AN2D0 U4185 ( .A1(n[1848]), .A2(b[9]), .Z(n[3895]) );
  AN2D0 U4186 ( .A1(n[1847]), .A2(b[9]), .Z(n[3894]) );
  AN2D0 U4187 ( .A1(n[1846]), .A2(b[9]), .Z(n[3893]) );
  AN2D0 U4188 ( .A1(n[1845]), .A2(b[9]), .Z(n[3892]) );
  AN2D0 U4189 ( .A1(n[1842]), .A2(b[9]), .Z(n[3889]) );
  AN2D0 U4190 ( .A1(n[1839]), .A2(b[9]), .Z(n[3886]) );
  AN2D0 U4191 ( .A1(n[1838]), .A2(b[9]), .Z(n[3885]) );
  AN2D0 U4192 ( .A1(n[1835]), .A2(b[9]), .Z(n[3882]) );
  AN2D0 U4193 ( .A1(n[1832]), .A2(b[9]), .Z(n[3879]) );
  AN2D0 U4194 ( .A1(n[1831]), .A2(b[9]), .Z(n[3878]) );
  AN2D0 U4195 ( .A1(n[1830]), .A2(b[9]), .Z(n[3877]) );
  AN2D0 U4196 ( .A1(n[1827]), .A2(b[9]), .Z(n[3874]) );
  AN2D0 U4197 ( .A1(n[1824]), .A2(b[9]), .Z(n[3871]) );
  AN2D0 U4198 ( .A1(n[1823]), .A2(b[9]), .Z(n[3870]) );
  AN2D0 U4199 ( .A1(n[1820]), .A2(b[9]), .Z(n[3867]) );
  AN2D0 U4200 ( .A1(n[1817]), .A2(b[9]), .Z(n[3864]) );
  AN2D0 U4201 ( .A1(n[1816]), .A2(b[9]), .Z(n[3863]) );
  AN2D0 U4202 ( .A1(n[1815]), .A2(b[9]), .Z(n[3862]) );
  AN2D0 U4203 ( .A1(n[1814]), .A2(b[9]), .Z(n[3861]) );
  AN2D0 U4204 ( .A1(n[1811]), .A2(b[9]), .Z(n[3858]) );
  AN2D0 U4205 ( .A1(n[1808]), .A2(b[9]), .Z(n[3855]) );
  AN2D0 U4206 ( .A1(n[1807]), .A2(b[9]), .Z(n[3854]) );
  AN2D0 U4207 ( .A1(n[1804]), .A2(b[9]), .Z(n[3851]) );
  AN2D0 U4208 ( .A1(n[1801]), .A2(b[9]), .Z(n[3848]) );
  AN2D0 U4209 ( .A1(n[1800]), .A2(b[9]), .Z(n[3847]) );
  AN2D0 U4210 ( .A1(n[1799]), .A2(b[9]), .Z(n[3846]) );
  AN2D0 U4211 ( .A1(n[1796]), .A2(b[9]), .Z(n[3843]) );
  AN2D0 U4212 ( .A1(n[1793]), .A2(b[9]), .Z(n[3840]) );
  AN2D0 U4213 ( .A1(n[1792]), .A2(b[9]), .Z(n[3839]) );
  AN2D0 U4214 ( .A1(n[1789]), .A2(b[9]), .Z(n[3836]) );
  AN2D0 U4215 ( .A1(n[1786]), .A2(b[9]), .Z(n[3833]) );
  AN2D0 U4216 ( .A1(n[1785]), .A2(b[9]), .Z(n[3832]) );
  AN2D0 U4217 ( .A1(n[1784]), .A2(b[9]), .Z(n[3831]) );
  AN2D0 U4218 ( .A1(n[1783]), .A2(b[9]), .Z(n[3830]) );
  AN2D0 U4219 ( .A1(n[1782]), .A2(b[9]), .Z(n[3829]) );
  AN2D0 U4220 ( .A1(n[1781]), .A2(b[9]), .Z(n[3828]) );
  AN2D0 U4221 ( .A1(n[1780]), .A2(b[9]), .Z(n[3827]) );
  AN2D0 U4222 ( .A1(n[1777]), .A2(b[9]), .Z(n[3824]) );
  AN2D0 U4223 ( .A1(n[1774]), .A2(b[9]), .Z(n[3821]) );
  AN2D0 U4224 ( .A1(n[1773]), .A2(b[9]), .Z(n[3820]) );
  AN2D0 U4225 ( .A1(n[1770]), .A2(b[9]), .Z(n[3817]) );
  AN2D0 U4226 ( .A1(n[1767]), .A2(b[9]), .Z(n[3814]) );
  AN2D0 U4227 ( .A1(n[1766]), .A2(b[9]), .Z(n[3813]) );
  AN2D0 U4228 ( .A1(n[1765]), .A2(b[9]), .Z(n[3812]) );
  AN2D0 U4229 ( .A1(n[1762]), .A2(b[9]), .Z(n[3809]) );
  AN2D0 U4230 ( .A1(n[1759]), .A2(b[9]), .Z(n[3806]) );
  AN2D0 U4231 ( .A1(n[1758]), .A2(b[9]), .Z(n[3805]) );
  AN2D0 U4232 ( .A1(n[1755]), .A2(b[9]), .Z(n[3802]) );
  AN2D0 U4233 ( .A1(n[1752]), .A2(b[9]), .Z(n[3799]) );
  AN2D0 U4234 ( .A1(n[1751]), .A2(b[9]), .Z(n[3798]) );
  AN2D0 U4235 ( .A1(n[1750]), .A2(b[9]), .Z(n[3797]) );
  AN2D0 U4236 ( .A1(n[1749]), .A2(b[9]), .Z(n[3796]) );
  AN2D0 U4237 ( .A1(n[1746]), .A2(b[9]), .Z(n[3793]) );
  AN2D0 U4238 ( .A1(n[1743]), .A2(b[9]), .Z(n[3790]) );
  AN2D0 U4239 ( .A1(n[1742]), .A2(b[9]), .Z(n[3789]) );
  AN2D0 U4240 ( .A1(n[1739]), .A2(b[9]), .Z(n[3786]) );
  AN2D0 U4241 ( .A1(n[1736]), .A2(b[9]), .Z(n[3783]) );
  AN2D0 U4242 ( .A1(n[1735]), .A2(b[9]), .Z(n[3782]) );
  AN2D0 U4243 ( .A1(n[1734]), .A2(b[9]), .Z(n[3781]) );
  AN2D0 U4244 ( .A1(n[1731]), .A2(b[9]), .Z(n[3778]) );
  AN2D0 U4245 ( .A1(n[1728]), .A2(b[9]), .Z(n[3775]) );
  AN2D0 U4246 ( .A1(n[1727]), .A2(b[9]), .Z(n[3774]) );
  AN2D0 U4247 ( .A1(n[1724]), .A2(b[9]), .Z(n[3771]) );
  AN2D0 U4248 ( .A1(n[1721]), .A2(b[9]), .Z(n[3768]) );
  AN2D0 U4249 ( .A1(n[1720]), .A2(b[9]), .Z(n[3767]) );
  AN2D0 U4250 ( .A1(n[1719]), .A2(b[9]), .Z(n[3766]) );
  AN2D0 U4251 ( .A1(n[1718]), .A2(b[9]), .Z(n[3765]) );
  AN2D0 U4252 ( .A1(n[1717]), .A2(b[9]), .Z(n[3764]) );
  AN2D0 U4253 ( .A1(n[1714]), .A2(b[9]), .Z(n[3761]) );
  AN2D0 U4254 ( .A1(n[1711]), .A2(b[9]), .Z(n[3758]) );
  AN2D0 U4255 ( .A1(n[1710]), .A2(b[9]), .Z(n[3757]) );
  AN2D0 U4256 ( .A1(n[1707]), .A2(b[9]), .Z(n[3754]) );
  AN2D0 U4257 ( .A1(n[1704]), .A2(b[9]), .Z(n[3751]) );
  AN2D0 U4258 ( .A1(n[1703]), .A2(b[9]), .Z(n[3750]) );
  AN2D0 U4259 ( .A1(n[1702]), .A2(b[9]), .Z(n[3749]) );
  AN2D0 U4260 ( .A1(n[1699]), .A2(b[9]), .Z(n[3746]) );
  AN2D0 U4261 ( .A1(n[1696]), .A2(b[9]), .Z(n[3743]) );
  AN2D0 U4262 ( .A1(n[1695]), .A2(b[9]), .Z(n[3742]) );
  AN2D0 U4263 ( .A1(n[1692]), .A2(b[9]), .Z(n[3739]) );
  AN2D0 U4264 ( .A1(n[1689]), .A2(b[9]), .Z(n[3736]) );
  AN2D0 U4265 ( .A1(n[1688]), .A2(b[9]), .Z(n[3735]) );
  AN2D0 U4266 ( .A1(n[1687]), .A2(b[9]), .Z(n[3734]) );
  AN2D0 U4267 ( .A1(n[1686]), .A2(b[9]), .Z(n[3733]) );
  AN2D0 U4268 ( .A1(n[1683]), .A2(b[9]), .Z(n[3730]) );
  AN2D0 U4269 ( .A1(n[1680]), .A2(b[9]), .Z(n[3727]) );
  AN2D0 U4270 ( .A1(n[1679]), .A2(b[9]), .Z(n[3726]) );
  AN2D0 U4271 ( .A1(n[1676]), .A2(b[9]), .Z(n[3723]) );
  AN2D0 U4272 ( .A1(n[1673]), .A2(b[9]), .Z(n[3720]) );
  AN2D0 U4273 ( .A1(n[1672]), .A2(b[9]), .Z(n[3719]) );
  AN2D0 U4274 ( .A1(n[1671]), .A2(b[9]), .Z(n[3718]) );
  AN2D0 U4275 ( .A1(n[1668]), .A2(b[9]), .Z(n[3715]) );
  AN2D0 U4276 ( .A1(n[1665]), .A2(b[9]), .Z(n[3712]) );
  AN2D0 U4277 ( .A1(n[1664]), .A2(b[9]), .Z(n[3711]) );
  AN2D0 U4278 ( .A1(n[1661]), .A2(b[9]), .Z(n[3708]) );
  AN2D0 U4279 ( .A1(n[1658]), .A2(b[9]), .Z(n[3705]) );
  AN2D0 U4280 ( .A1(n[1657]), .A2(b[9]), .Z(n[3704]) );
  AN2D0 U4281 ( .A1(n[1656]), .A2(b[9]), .Z(n[3703]) );
  AN2D0 U4282 ( .A1(n[1655]), .A2(b[9]), .Z(n[3702]) );
  AN2D0 U4283 ( .A1(n[1654]), .A2(b[9]), .Z(n[3701]) );
  AN2D0 U4284 ( .A1(n[1653]), .A2(b[9]), .Z(n[3700]) );
  AN2D0 U4285 ( .A1(n[1650]), .A2(b[9]), .Z(n[3697]) );
  AN2D0 U4286 ( .A1(n[1647]), .A2(b[9]), .Z(n[3694]) );
  AN2D0 U4287 ( .A1(n[1646]), .A2(b[9]), .Z(n[3693]) );
  AN2D0 U4288 ( .A1(n[1643]), .A2(b[9]), .Z(n[3690]) );
  AN2D0 U4289 ( .A1(n[1640]), .A2(b[9]), .Z(n[3687]) );
  AN2D0 U4290 ( .A1(n[1639]), .A2(b[9]), .Z(n[3686]) );
  AN2D0 U4291 ( .A1(n[1638]), .A2(b[9]), .Z(n[3685]) );
  AN2D0 U4292 ( .A1(n[1635]), .A2(b[9]), .Z(n[3682]) );
  AN2D0 U4293 ( .A1(n[1632]), .A2(b[9]), .Z(n[3679]) );
  AN2D0 U4294 ( .A1(n[1631]), .A2(b[9]), .Z(n[3678]) );
  AN2D0 U4295 ( .A1(n[1628]), .A2(b[9]), .Z(n[3675]) );
  AN2D0 U4296 ( .A1(n[1625]), .A2(b[9]), .Z(n[3672]) );
  AN2D0 U4297 ( .A1(n[1624]), .A2(b[9]), .Z(n[3671]) );
  AN2D0 U4298 ( .A1(n[1623]), .A2(b[9]), .Z(n[3670]) );
  AN2D0 U4299 ( .A1(n[1622]), .A2(b[9]), .Z(n[3669]) );
  AN2D0 U4300 ( .A1(n[1619]), .A2(b[9]), .Z(n[3666]) );
  AN2D0 U4301 ( .A1(n[1616]), .A2(b[9]), .Z(n[3663]) );
  AN2D0 U4302 ( .A1(n[1615]), .A2(b[9]), .Z(n[3662]) );
  AN2D0 U4303 ( .A1(n[1612]), .A2(b[9]), .Z(n[3659]) );
  AN2D0 U4304 ( .A1(n[1609]), .A2(b[9]), .Z(n[3656]) );
  AN2D0 U4305 ( .A1(n[1608]), .A2(b[9]), .Z(n[3655]) );
  AN2D0 U4306 ( .A1(n[1607]), .A2(b[9]), .Z(n[3654]) );
  AN2D0 U4307 ( .A1(n[1604]), .A2(b[9]), .Z(n[3651]) );
  AN2D0 U4308 ( .A1(n[1601]), .A2(b[9]), .Z(n[3648]) );
  AN2D0 U4309 ( .A1(n[1600]), .A2(b[9]), .Z(n[3647]) );
  AN2D0 U4310 ( .A1(n[1597]), .A2(b[9]), .Z(n[3644]) );
  AN2D0 U4311 ( .A1(n[1594]), .A2(b[9]), .Z(n[3641]) );
  AN2D0 U4312 ( .A1(n[1593]), .A2(b[9]), .Z(n[3640]) );
  AN2D0 U4313 ( .A1(n[1592]), .A2(b[9]), .Z(n[3639]) );
  AN2D0 U4314 ( .A1(n[1591]), .A2(b[9]), .Z(n[3638]) );
  AN2D0 U4315 ( .A1(n[1590]), .A2(b[9]), .Z(n[3637]) );
  AN2D0 U4316 ( .A1(n[1587]), .A2(b[9]), .Z(n[3634]) );
  AN2D0 U4317 ( .A1(n[1584]), .A2(b[9]), .Z(n[3631]) );
  AN2D0 U4318 ( .A1(n[1583]), .A2(b[9]), .Z(n[3630]) );
  AN2D0 U4319 ( .A1(n[1580]), .A2(b[9]), .Z(n[3627]) );
  AN2D0 U4320 ( .A1(n[1577]), .A2(b[9]), .Z(n[3624]) );
  AN2D0 U4321 ( .A1(n[1576]), .A2(b[9]), .Z(n[3623]) );
  AN2D0 U4322 ( .A1(n[1575]), .A2(b[9]), .Z(n[3622]) );
  AN2D0 U4323 ( .A1(n[1572]), .A2(b[9]), .Z(n[3619]) );
  AN2D0 U4324 ( .A1(n[1569]), .A2(b[9]), .Z(n[3616]) );
  AN2D0 U4325 ( .A1(n[1568]), .A2(b[9]), .Z(n[3615]) );
  AN2D0 U4326 ( .A1(n[1565]), .A2(b[9]), .Z(n[3612]) );
  AN2D0 U4327 ( .A1(n[1562]), .A2(b[9]), .Z(n[3609]) );
  AN2D0 U4328 ( .A1(n[1561]), .A2(b[9]), .Z(n[3608]) );
  AN2D0 U4329 ( .A1(n[1560]), .A2(b[9]), .Z(n[3607]) );
  AN2D0 U4330 ( .A1(n[1559]), .A2(b[9]), .Z(n[3606]) );
  AN2D0 U4331 ( .A1(n[1556]), .A2(b[9]), .Z(n[3603]) );
  AN2D0 U4332 ( .A1(n[1553]), .A2(b[9]), .Z(n[3600]) );
  AN2D0 U4333 ( .A1(n[1552]), .A2(b[9]), .Z(n[3599]) );
  AN2D0 U4334 ( .A1(n[1549]), .A2(b[9]), .Z(n[3596]) );
  AN2D0 U4335 ( .A1(n[1546]), .A2(b[9]), .Z(n[3593]) );
  AN2D0 U4336 ( .A1(n[1545]), .A2(b[9]), .Z(n[3592]) );
  AN2D0 U4337 ( .A1(n[1544]), .A2(b[9]), .Z(n[3591]) );
  AN2D0 U4338 ( .A1(n[1541]), .A2(b[9]), .Z(n[3588]) );
  AN2D0 U4339 ( .A1(n[1538]), .A2(b[9]), .Z(n[3585]) );
  AN2D0 U4340 ( .A1(n[1537]), .A2(b[9]), .Z(n[3584]) );
  AN2D0 U4341 ( .A1(n[1534]), .A2(b[9]), .Z(n[3581]) );
  AN2D0 U4342 ( .A1(n[1531]), .A2(b[9]), .Z(n[3578]) );
  AN2D0 U4343 ( .A1(n[1530]), .A2(b[9]), .Z(n[3577]) );
  AN2D0 U4344 ( .A1(n[1529]), .A2(b[9]), .Z(n[3576]) );
  AN2D0 U4345 ( .A1(n[1528]), .A2(b[9]), .Z(n[3575]) );
  AN2D0 U4346 ( .A1(n[1527]), .A2(b[9]), .Z(n[3574]) );
  AN2D0 U4347 ( .A1(n[1526]), .A2(b[9]), .Z(n[3573]) );
  AN2D0 U4348 ( .A1(n[1525]), .A2(b[9]), .Z(n[3572]) );
  AN2D0 U4349 ( .A1(n[1524]), .A2(b[9]), .Z(n[3571]) );
  AN2D0 U4350 ( .A1(n[1521]), .A2(b[9]), .Z(n[3568]) );
  AN2D0 U4351 ( .A1(n[1518]), .A2(b[9]), .Z(n[3565]) );
  AN2D0 U4352 ( .A1(n[1517]), .A2(b[9]), .Z(n[3564]) );
  AN2D0 U4353 ( .A1(n[1514]), .A2(b[9]), .Z(n[3561]) );
  AN2D0 U4354 ( .A1(n[1511]), .A2(b[9]), .Z(n[3558]) );
  AN2D0 U4355 ( .A1(n[1510]), .A2(b[9]), .Z(n[3557]) );
  AN2D0 U4356 ( .A1(n[1509]), .A2(b[9]), .Z(n[3556]) );
  AN2D0 U4357 ( .A1(n[1506]), .A2(b[9]), .Z(n[3553]) );
  AN2D0 U4358 ( .A1(n[1503]), .A2(b[9]), .Z(n[3550]) );
  AN2D0 U4359 ( .A1(n[1502]), .A2(b[9]), .Z(n[3549]) );
  AN2D0 U4360 ( .A1(n[1499]), .A2(b[9]), .Z(n[3546]) );
  AN2D0 U4361 ( .A1(n[1496]), .A2(b[9]), .Z(n[3543]) );
  AN2D0 U4362 ( .A1(n[1495]), .A2(b[9]), .Z(n[3542]) );
  AN2D0 U4363 ( .A1(n[1494]), .A2(b[9]), .Z(n[3541]) );
  AN2D0 U4364 ( .A1(n[1493]), .A2(b[9]), .Z(n[3540]) );
  AN2D0 U4365 ( .A1(n[1490]), .A2(b[9]), .Z(n[3537]) );
  AN2D0 U4366 ( .A1(n[1487]), .A2(b[9]), .Z(n[3534]) );
  AN2D0 U4367 ( .A1(n[1486]), .A2(b[9]), .Z(n[3533]) );
  AN2D0 U4368 ( .A1(n[1483]), .A2(b[9]), .Z(n[3530]) );
  AN2D0 U4369 ( .A1(n[1480]), .A2(b[9]), .Z(n[3527]) );
  AN2D0 U4370 ( .A1(n[1479]), .A2(b[9]), .Z(n[3526]) );
  AN2D0 U4371 ( .A1(n[1478]), .A2(b[9]), .Z(n[3525]) );
  AN2D0 U4372 ( .A1(n[1475]), .A2(b[9]), .Z(n[3522]) );
  AN2D0 U4373 ( .A1(n[1472]), .A2(b[9]), .Z(n[3519]) );
  AN2D0 U4374 ( .A1(n[1471]), .A2(b[9]), .Z(n[3518]) );
  AN2D0 U4375 ( .A1(n[1468]), .A2(b[9]), .Z(n[3515]) );
  AN2D0 U4376 ( .A1(n[1465]), .A2(b[9]), .Z(n[3512]) );
  AN2D0 U4377 ( .A1(n[1464]), .A2(b[9]), .Z(n[3511]) );
  AN2D0 U4378 ( .A1(n[1463]), .A2(b[9]), .Z(n[3510]) );
  AN2D0 U4379 ( .A1(n[1462]), .A2(b[9]), .Z(n[3509]) );
  AN2D0 U4380 ( .A1(n[1461]), .A2(b[9]), .Z(n[3508]) );
  AN2D0 U4381 ( .A1(n[1458]), .A2(b[9]), .Z(n[3505]) );
  AN2D0 U4382 ( .A1(n[1455]), .A2(b[9]), .Z(n[3502]) );
  AN2D0 U4383 ( .A1(n[1454]), .A2(b[9]), .Z(n[3501]) );
  AN2D0 U4384 ( .A1(n[1451]), .A2(b[9]), .Z(n[3498]) );
  AN2D0 U4385 ( .A1(n[1448]), .A2(b[9]), .Z(n[3495]) );
  AN2D0 U4386 ( .A1(n[1447]), .A2(b[9]), .Z(n[3494]) );
  AN2D0 U4387 ( .A1(n[1446]), .A2(b[9]), .Z(n[3493]) );
  AN2D0 U4388 ( .A1(n[1443]), .A2(b[9]), .Z(n[3490]) );
  AN2D0 U4389 ( .A1(n[1440]), .A2(b[9]), .Z(n[3487]) );
  AN2D0 U4390 ( .A1(n[1439]), .A2(b[9]), .Z(n[3486]) );
  AN2D0 U4391 ( .A1(n[1436]), .A2(b[9]), .Z(n[3483]) );
  AN2D0 U4392 ( .A1(n[1433]), .A2(b[9]), .Z(n[3480]) );
  AN2D0 U4393 ( .A1(n[1432]), .A2(b[9]), .Z(n[3479]) );
  AN2D0 U4394 ( .A1(n[1431]), .A2(b[9]), .Z(n[3478]) );
  AN2D0 U4395 ( .A1(n[1430]), .A2(b[9]), .Z(n[3477]) );
  AN2D0 U4396 ( .A1(n[1427]), .A2(b[9]), .Z(n[3474]) );
  AN2D0 U4397 ( .A1(n[1424]), .A2(b[9]), .Z(n[3471]) );
  AN2D0 U4398 ( .A1(n[1423]), .A2(b[9]), .Z(n[3470]) );
  AN2D0 U4399 ( .A1(n[1420]), .A2(b[9]), .Z(n[3467]) );
  AN2D0 U4400 ( .A1(n[1417]), .A2(b[9]), .Z(n[3464]) );
  AN2D0 U4401 ( .A1(n[1416]), .A2(b[9]), .Z(n[3463]) );
  AN2D0 U4402 ( .A1(n[1415]), .A2(b[9]), .Z(n[3462]) );
  AN2D0 U4403 ( .A1(n[1412]), .A2(b[9]), .Z(n[3459]) );
  AN2D0 U4404 ( .A1(n[1409]), .A2(b[9]), .Z(n[3456]) );
  AN2D0 U4405 ( .A1(n[1408]), .A2(b[9]), .Z(n[3455]) );
  AN2D0 U4406 ( .A1(n[1405]), .A2(b[9]), .Z(n[3452]) );
  AN2D0 U4407 ( .A1(n[1402]), .A2(b[9]), .Z(n[3449]) );
  AN2D0 U4408 ( .A1(n[1401]), .A2(b[9]), .Z(n[3448]) );
  AN2D0 U4409 ( .A1(n[1400]), .A2(b[9]), .Z(n[3447]) );
  AN2D0 U4410 ( .A1(n[1399]), .A2(b[9]), .Z(n[3446]) );
  AN2D0 U4411 ( .A1(n[1398]), .A2(b[9]), .Z(n[3445]) );
  AN2D0 U4412 ( .A1(n[1397]), .A2(b[9]), .Z(n[3444]) );
  AN2D0 U4413 ( .A1(n[1394]), .A2(b[9]), .Z(n[3441]) );
  AN2D0 U4414 ( .A1(n[1391]), .A2(b[9]), .Z(n[3438]) );
  AN2D0 U4415 ( .A1(n[1390]), .A2(b[9]), .Z(n[3437]) );
  AN2D0 U4416 ( .A1(n[1387]), .A2(b[9]), .Z(n[3434]) );
  AN2D0 U4417 ( .A1(n[1384]), .A2(b[9]), .Z(n[3431]) );
  AN2D0 U4418 ( .A1(n[1383]), .A2(b[9]), .Z(n[3430]) );
  AN2D0 U4419 ( .A1(n[1382]), .A2(b[9]), .Z(n[3429]) );
  AN2D0 U4420 ( .A1(n[1379]), .A2(b[9]), .Z(n[3426]) );
  AN2D0 U4421 ( .A1(n[1376]), .A2(b[9]), .Z(n[3423]) );
  AN2D0 U4422 ( .A1(n[1375]), .A2(b[9]), .Z(n[3422]) );
  AN2D0 U4423 ( .A1(n[1372]), .A2(b[9]), .Z(n[3419]) );
  AN2D0 U4424 ( .A1(n[1369]), .A2(b[9]), .Z(n[3416]) );
  AN2D0 U4425 ( .A1(n[1368]), .A2(b[9]), .Z(n[3415]) );
  AN2D0 U4426 ( .A1(n[1367]), .A2(b[9]), .Z(n[3414]) );
  AN2D0 U4427 ( .A1(n[1366]), .A2(b[9]), .Z(n[3413]) );
  AN2D0 U4428 ( .A1(n[1363]), .A2(b[9]), .Z(n[3410]) );
  AN2D0 U4429 ( .A1(n[1360]), .A2(b[9]), .Z(n[3407]) );
  AN2D0 U4430 ( .A1(n[1359]), .A2(b[9]), .Z(n[3406]) );
  AN2D0 U4431 ( .A1(n[1356]), .A2(b[9]), .Z(n[3403]) );
  AN2D0 U4432 ( .A1(n[1353]), .A2(b[9]), .Z(n[3400]) );
  AN2D0 U4433 ( .A1(n[1352]), .A2(b[9]), .Z(n[3399]) );
  AN2D0 U4434 ( .A1(n[1351]), .A2(b[9]), .Z(n[3398]) );
  AN2D0 U4435 ( .A1(n[1348]), .A2(b[9]), .Z(n[3395]) );
  AN2D0 U4436 ( .A1(n[1345]), .A2(b[9]), .Z(n[3392]) );
  AN2D0 U4437 ( .A1(n[1344]), .A2(b[9]), .Z(n[3391]) );
  AN2D0 U4438 ( .A1(n[1341]), .A2(b[9]), .Z(n[3388]) );
  AN2D0 U4439 ( .A1(n[1338]), .A2(b[9]), .Z(n[3385]) );
  AN2D0 U4440 ( .A1(n[1337]), .A2(b[9]), .Z(n[3384]) );
  AN2D0 U4441 ( .A1(n[1336]), .A2(b[9]), .Z(n[3383]) );
  AN2D0 U4442 ( .A1(n[1335]), .A2(b[9]), .Z(n[3382]) );
  AN2D0 U4443 ( .A1(n[1334]), .A2(b[9]), .Z(n[3381]) );
  AN2D0 U4444 ( .A1(n[1331]), .A2(b[9]), .Z(n[3378]) );
  AN2D0 U4445 ( .A1(n[1328]), .A2(b[9]), .Z(n[3375]) );
  AN2D0 U4446 ( .A1(n[1327]), .A2(b[9]), .Z(n[3374]) );
  AN2D0 U4447 ( .A1(n[1324]), .A2(b[9]), .Z(n[3371]) );
  AN2D0 U4448 ( .A1(n[1321]), .A2(b[9]), .Z(n[3368]) );
  AN2D0 U4449 ( .A1(n[1320]), .A2(b[9]), .Z(n[3367]) );
  AN2D0 U4450 ( .A1(n[1319]), .A2(b[9]), .Z(n[3366]) );
  AN2D0 U4451 ( .A1(n[1316]), .A2(b[9]), .Z(n[3363]) );
  AN2D0 U4452 ( .A1(n[1313]), .A2(b[9]), .Z(n[3360]) );
  AN2D0 U4453 ( .A1(n[1312]), .A2(b[9]), .Z(n[3359]) );
  AN2D0 U4454 ( .A1(n[1309]), .A2(b[9]), .Z(n[3356]) );
  AN2D0 U4455 ( .A1(n[1306]), .A2(b[9]), .Z(n[3353]) );
  AN2D0 U4456 ( .A1(n[1305]), .A2(b[9]), .Z(n[3352]) );
  AN2D0 U4457 ( .A1(n[1304]), .A2(b[9]), .Z(n[3351]) );
  AN2D0 U4458 ( .A1(n[1303]), .A2(b[9]), .Z(n[3350]) );
  AN2D0 U4459 ( .A1(n[1300]), .A2(b[9]), .Z(n[3347]) );
  AN2D0 U4460 ( .A1(n[1297]), .A2(b[9]), .Z(n[3344]) );
  AN2D0 U4461 ( .A1(n[1296]), .A2(b[9]), .Z(n[3343]) );
  AN2D0 U4462 ( .A1(n[1293]), .A2(b[9]), .Z(n[3340]) );
  AN2D0 U4463 ( .A1(n[1290]), .A2(b[9]), .Z(n[3337]) );
  AN2D0 U4464 ( .A1(n[1289]), .A2(b[9]), .Z(n[3336]) );
  AN2D0 U4465 ( .A1(n[1288]), .A2(b[9]), .Z(n[3335]) );
  AN2D0 U4466 ( .A1(n[1285]), .A2(b[9]), .Z(n[3332]) );
  AN2D0 U4467 ( .A1(n[1282]), .A2(b[9]), .Z(n[3329]) );
  AN2D0 U4468 ( .A1(n[1281]), .A2(b[9]), .Z(n[3328]) );
  AN2D0 U4469 ( .A1(n[1278]), .A2(b[9]), .Z(n[3325]) );
  AN2D0 U4470 ( .A1(n[1275]), .A2(b[9]), .Z(n[3322]) );
  AN2D0 U4471 ( .A1(n[1274]), .A2(b[9]), .Z(n[3321]) );
  AN2D0 U4472 ( .A1(n[1273]), .A2(b[9]), .Z(n[3320]) );
  AN2D0 U4473 ( .A1(n[1272]), .A2(b[9]), .Z(n[3319]) );
  AN2D0 U4474 ( .A1(n[1271]), .A2(b[9]), .Z(n[3318]) );
  AN2D0 U4475 ( .A1(n[1270]), .A2(b[9]), .Z(n[3317]) );
  AN2D0 U4476 ( .A1(n[1269]), .A2(b[9]), .Z(n[3316]) );
  AN2D0 U4477 ( .A1(n[1266]), .A2(b[9]), .Z(n[3313]) );
  AN2D0 U4478 ( .A1(n[1263]), .A2(b[9]), .Z(n[3310]) );
  AN2D0 U4479 ( .A1(n[1262]), .A2(b[9]), .Z(n[3309]) );
  AN2D0 U4480 ( .A1(n[1259]), .A2(b[9]), .Z(n[3306]) );
  AN2D0 U4481 ( .A1(n[1256]), .A2(b[9]), .Z(n[3303]) );
  AN2D0 U4482 ( .A1(n[1255]), .A2(b[9]), .Z(n[3302]) );
  AN2D0 U4483 ( .A1(n[1254]), .A2(b[9]), .Z(n[3301]) );
  AN2D0 U4484 ( .A1(n[1251]), .A2(b[9]), .Z(n[3298]) );
  AN2D0 U4485 ( .A1(n[1248]), .A2(b[9]), .Z(n[3295]) );
  AN2D0 U4486 ( .A1(n[1247]), .A2(b[9]), .Z(n[3294]) );
  AN2D0 U4487 ( .A1(n[1244]), .A2(b[9]), .Z(n[3291]) );
  AN2D0 U4488 ( .A1(n[1241]), .A2(b[9]), .Z(n[3288]) );
  AN2D0 U4489 ( .A1(n[1240]), .A2(b[9]), .Z(n[3287]) );
  AN2D0 U4490 ( .A1(n[1239]), .A2(b[9]), .Z(n[3286]) );
  AN2D0 U4491 ( .A1(n[1238]), .A2(b[9]), .Z(n[3285]) );
  AN2D0 U4492 ( .A1(n[1235]), .A2(b[9]), .Z(n[3282]) );
  AN2D0 U4493 ( .A1(n[1232]), .A2(b[9]), .Z(n[3279]) );
  AN2D0 U4494 ( .A1(n[1231]), .A2(b[9]), .Z(n[3278]) );
  AN2D0 U4495 ( .A1(n[1228]), .A2(b[9]), .Z(n[3275]) );
  AN2D0 U4496 ( .A1(n[1225]), .A2(b[9]), .Z(n[3272]) );
  AN2D0 U4497 ( .A1(n[1224]), .A2(b[9]), .Z(n[3271]) );
  AN2D0 U4498 ( .A1(n[1223]), .A2(b[9]), .Z(n[3270]) );
  AN2D0 U4499 ( .A1(n[1220]), .A2(b[9]), .Z(n[3267]) );
  AN2D0 U4500 ( .A1(n[1217]), .A2(b[9]), .Z(n[3264]) );
  AN2D0 U4501 ( .A1(n[1216]), .A2(b[9]), .Z(n[3263]) );
  AN2D0 U4502 ( .A1(n[1213]), .A2(b[9]), .Z(n[3260]) );
  AN2D0 U4503 ( .A1(n[1210]), .A2(b[9]), .Z(n[3257]) );
  AN2D0 U4504 ( .A1(n[1209]), .A2(b[9]), .Z(n[3256]) );
  AN2D0 U4505 ( .A1(n[1208]), .A2(b[9]), .Z(n[3255]) );
  AN2D0 U4506 ( .A1(n[1207]), .A2(b[9]), .Z(n[3254]) );
  AN2D0 U4507 ( .A1(n[1206]), .A2(b[9]), .Z(n[3253]) );
  AN2D0 U4508 ( .A1(n[1203]), .A2(b[9]), .Z(n[3250]) );
  AN2D0 U4509 ( .A1(n[1200]), .A2(b[9]), .Z(n[3247]) );
  AN2D0 U4510 ( .A1(n[1199]), .A2(b[9]), .Z(n[3246]) );
  AN2D0 U4511 ( .A1(n[1196]), .A2(b[9]), .Z(n[3243]) );
  AN2D0 U4512 ( .A1(n[1193]), .A2(b[9]), .Z(n[3240]) );
  AN2D0 U4513 ( .A1(n[1192]), .A2(b[9]), .Z(n[3239]) );
  AN2D0 U4514 ( .A1(n[1191]), .A2(b[9]), .Z(n[3238]) );
  AN2D0 U4515 ( .A1(n[1188]), .A2(b[9]), .Z(n[3235]) );
  AN2D0 U4516 ( .A1(n[1185]), .A2(b[9]), .Z(n[3232]) );
  AN2D0 U4517 ( .A1(n[1184]), .A2(b[9]), .Z(n[3231]) );
  AN2D0 U4518 ( .A1(n[1181]), .A2(b[9]), .Z(n[3228]) );
  AN2D0 U4519 ( .A1(n[1178]), .A2(b[9]), .Z(n[3225]) );
  AN2D0 U4520 ( .A1(n[1177]), .A2(b[9]), .Z(n[3224]) );
  AN2D0 U4521 ( .A1(n[1176]), .A2(b[9]), .Z(n[3223]) );
  AN2D0 U4522 ( .A1(n[1175]), .A2(b[9]), .Z(n[3222]) );
  AN2D0 U4523 ( .A1(n[1172]), .A2(b[9]), .Z(n[3219]) );
  AN2D0 U4524 ( .A1(n[1169]), .A2(b[9]), .Z(n[3216]) );
  AN2D0 U4525 ( .A1(n[1168]), .A2(b[9]), .Z(n[3215]) );
  AN2D0 U4526 ( .A1(n[1165]), .A2(b[9]), .Z(n[3212]) );
  AN2D0 U4527 ( .A1(n[1162]), .A2(b[9]), .Z(n[3209]) );
  AN2D0 U4528 ( .A1(n[1161]), .A2(b[9]), .Z(n[3208]) );
  AN2D0 U4529 ( .A1(n[1160]), .A2(b[9]), .Z(n[3207]) );
  AN2D0 U4530 ( .A1(n[1157]), .A2(b[9]), .Z(n[3204]) );
  AN2D0 U4531 ( .A1(n[1154]), .A2(b[9]), .Z(n[3201]) );
  AN2D0 U4532 ( .A1(n[1153]), .A2(b[9]), .Z(n[3200]) );
  AN2D0 U4533 ( .A1(n[1150]), .A2(b[9]), .Z(n[3197]) );
  AN2D0 U4534 ( .A1(n[1147]), .A2(b[9]), .Z(n[3194]) );
  AN2D0 U4535 ( .A1(n[1146]), .A2(b[9]), .Z(n[3193]) );
  AN2D0 U4536 ( .A1(n[1145]), .A2(b[9]), .Z(n[3192]) );
  AN2D0 U4537 ( .A1(n[1144]), .A2(b[9]), .Z(n[3191]) );
  AN2D0 U4538 ( .A1(n[1143]), .A2(b[9]), .Z(n[3190]) );
  AN2D0 U4539 ( .A1(n[1142]), .A2(b[9]), .Z(n[3189]) );
  AN2D0 U4540 ( .A1(n[1139]), .A2(b[9]), .Z(n[3186]) );
  AN2D0 U4541 ( .A1(n[1136]), .A2(b[9]), .Z(n[3183]) );
  AN2D0 U4542 ( .A1(n[1135]), .A2(b[9]), .Z(n[3182]) );
  AN2D0 U4543 ( .A1(n[1132]), .A2(b[9]), .Z(n[3179]) );
  AN2D0 U4544 ( .A1(n[1129]), .A2(b[9]), .Z(n[3176]) );
  AN2D0 U4545 ( .A1(n[1128]), .A2(b[9]), .Z(n[3175]) );
  AN2D0 U4546 ( .A1(n[1127]), .A2(b[9]), .Z(n[3174]) );
  AN2D0 U4547 ( .A1(n[1124]), .A2(b[9]), .Z(n[3171]) );
  AN2D0 U4548 ( .A1(n[1121]), .A2(b[9]), .Z(n[3168]) );
  AN2D0 U4549 ( .A1(n[1120]), .A2(b[9]), .Z(n[3167]) );
  AN2D0 U4550 ( .A1(n[1117]), .A2(b[9]), .Z(n[3164]) );
  AN2D0 U4551 ( .A1(n[1114]), .A2(b[9]), .Z(n[3161]) );
  AN2D0 U4552 ( .A1(n[1113]), .A2(b[9]), .Z(n[3160]) );
  AN2D0 U4553 ( .A1(n[1112]), .A2(b[9]), .Z(n[3159]) );
  AN2D0 U4554 ( .A1(n[1111]), .A2(b[9]), .Z(n[3158]) );
  AN2D0 U4555 ( .A1(n[1108]), .A2(b[9]), .Z(n[3155]) );
  AN2D0 U4556 ( .A1(n[1105]), .A2(b[9]), .Z(n[3152]) );
  AN2D0 U4557 ( .A1(n[1104]), .A2(b[9]), .Z(n[3151]) );
  AN2D0 U4558 ( .A1(n[1101]), .A2(b[9]), .Z(n[3148]) );
  AN2D0 U4559 ( .A1(n[1098]), .A2(b[9]), .Z(n[3145]) );
  AN2D0 U4560 ( .A1(n[1097]), .A2(b[9]), .Z(n[3144]) );
  AN2D0 U4561 ( .A1(n[1096]), .A2(b[9]), .Z(n[3143]) );
  AN2D0 U4562 ( .A1(n[1093]), .A2(b[9]), .Z(n[3140]) );
  AN2D0 U4563 ( .A1(n[1090]), .A2(b[9]), .Z(n[3137]) );
  AN2D0 U4564 ( .A1(n[1089]), .A2(b[9]), .Z(n[3136]) );
  AN2D0 U4565 ( .A1(n[1086]), .A2(b[9]), .Z(n[3133]) );
  AN2D0 U4566 ( .A1(n[1083]), .A2(b[9]), .Z(n[3130]) );
  AN2D0 U4567 ( .A1(n[1082]), .A2(b[9]), .Z(n[3129]) );
  AN2D0 U4568 ( .A1(n[1081]), .A2(b[9]), .Z(n[3128]) );
  AN2D0 U4569 ( .A1(n[1080]), .A2(b[9]), .Z(n[3127]) );
  AN2D0 U4570 ( .A1(n[1079]), .A2(b[9]), .Z(n[3126]) );
  AN2D0 U4571 ( .A1(n[1076]), .A2(b[9]), .Z(n[3123]) );
  AN2D0 U4572 ( .A1(n[1073]), .A2(b[9]), .Z(n[3120]) );
  AN2D0 U4573 ( .A1(n[1072]), .A2(b[9]), .Z(n[3119]) );
  AN2D0 U4574 ( .A1(n[1069]), .A2(b[9]), .Z(n[3116]) );
  AN2D0 U4575 ( .A1(n[1066]), .A2(b[9]), .Z(n[3113]) );
  AN2D0 U4576 ( .A1(n[1065]), .A2(b[9]), .Z(n[3112]) );
  AN2D0 U4577 ( .A1(n[1064]), .A2(b[9]), .Z(n[3111]) );
  AN2D0 U4578 ( .A1(n[1061]), .A2(b[9]), .Z(n[3108]) );
  AN2D0 U4579 ( .A1(n[1058]), .A2(b[9]), .Z(n[3105]) );
  AN2D0 U4580 ( .A1(n[1057]), .A2(b[9]), .Z(n[3104]) );
  AN2D0 U4581 ( .A1(n[1054]), .A2(b[9]), .Z(n[3101]) );
  AN2D0 U4582 ( .A1(n[1051]), .A2(b[9]), .Z(n[3098]) );
  AN2D0 U4583 ( .A1(n[1050]), .A2(b[9]), .Z(n[3097]) );
  AN2D0 U4584 ( .A1(n[1049]), .A2(b[9]), .Z(n[3096]) );
  AN2D0 U4585 ( .A1(n[1048]), .A2(b[9]), .Z(n[3095]) );
  AN2D0 U4586 ( .A1(n[1045]), .A2(b[9]), .Z(n[3092]) );
  AN2D0 U4587 ( .A1(n[1042]), .A2(b[9]), .Z(n[3089]) );
  AN2D0 U4588 ( .A1(n[1041]), .A2(b[9]), .Z(n[3088]) );
  AN2D0 U4589 ( .A1(n[1038]), .A2(b[9]), .Z(n[3085]) );
  AN2D0 U4590 ( .A1(n[1035]), .A2(b[9]), .Z(n[3082]) );
  AN2D0 U4591 ( .A1(n[1034]), .A2(b[9]), .Z(n[3081]) );
  AN2D0 U4592 ( .A1(n[1033]), .A2(b[9]), .Z(n[3080]) );
  AN2D0 U4593 ( .A1(n[1030]), .A2(b[9]), .Z(n[3077]) );
  AN2D0 U4594 ( .A1(n[1027]), .A2(b[9]), .Z(n[3074]) );
  AN2D0 U4595 ( .A1(n[1026]), .A2(b[9]), .Z(n[3073]) );
  AN2D0 U4596 ( .A1(n[1023]), .A2(b[9]), .Z(n[3070]) );
  AN2D0 U4597 ( .A1(n[1020]), .A2(b[9]), .Z(n[3067]) );
  AN2D0 U4598 ( .A1(n[1019]), .A2(b[9]), .Z(n[3066]) );
  AN2D0 U4599 ( .A1(n[1018]), .A2(b[9]), .Z(n[3065]) );
  AN2D0 U4600 ( .A1(n[1017]), .A2(b[9]), .Z(n[3064]) );
  AN2D0 U4601 ( .A1(n[1016]), .A2(b[9]), .Z(n[3063]) );
  AN2D0 U4602 ( .A1(n[1015]), .A2(b[9]), .Z(n[3062]) );
  AN2D0 U4603 ( .A1(n[1014]), .A2(b[9]), .Z(n[3061]) );
  AN2D0 U4604 ( .A1(n[1013]), .A2(b[9]), .Z(n[3060]) );
  AN2D0 U4605 ( .A1(n[1012]), .A2(b[9]), .Z(n[3059]) );
  AN2D0 U4606 ( .A1(a[9]), .A2(n[2032]), .Z(n[3056]) );
  AN2D0 U4607 ( .A1(a[9]), .A2(n[2029]), .Z(n[3053]) );
  AN2D0 U4608 ( .A1(a[9]), .A2(n[2028]), .Z(n[3052]) );
  AN2D0 U4609 ( .A1(a[9]), .A2(n[2025]), .Z(n[3049]) );
  AN2D0 U4610 ( .A1(a[9]), .A2(n[2022]), .Z(n[3046]) );
  AN2D0 U4611 ( .A1(a[9]), .A2(n[2021]), .Z(n[3045]) );
  AN2D0 U4612 ( .A1(a[9]), .A2(n[2020]), .Z(n[3044]) );
  AN2D0 U4613 ( .A1(a[9]), .A2(n[2017]), .Z(n[3041]) );
  AN2D0 U4614 ( .A1(a[9]), .A2(n[2014]), .Z(n[3038]) );
  AN2D0 U4615 ( .A1(a[9]), .A2(n[2013]), .Z(n[3037]) );
  AN2D0 U4616 ( .A1(a[9]), .A2(n[2010]), .Z(n[3034]) );
  AN2D0 U4617 ( .A1(a[9]), .A2(n[2007]), .Z(n[3031]) );
  AN2D0 U4618 ( .A1(a[9]), .A2(n[2006]), .Z(n[3030]) );
  AN2D0 U4619 ( .A1(a[9]), .A2(n[2005]), .Z(n[3029]) );
  AN2D0 U4620 ( .A1(a[9]), .A2(n[2004]), .Z(n[3028]) );
  AN2D0 U4621 ( .A1(a[9]), .A2(n[2001]), .Z(n[3025]) );
  AN2D0 U4622 ( .A1(a[9]), .A2(n[1998]), .Z(n[3022]) );
  AN2D0 U4623 ( .A1(a[9]), .A2(n[1997]), .Z(n[3021]) );
  AN2D0 U4624 ( .A1(a[9]), .A2(n[1994]), .Z(n[3018]) );
  AN2D0 U4625 ( .A1(a[9]), .A2(n[1991]), .Z(n[3015]) );
  AN2D0 U4626 ( .A1(a[9]), .A2(n[1990]), .Z(n[3014]) );
  AN2D0 U4627 ( .A1(a[9]), .A2(n[1989]), .Z(n[3013]) );
  AN2D0 U4628 ( .A1(a[9]), .A2(n[1986]), .Z(n[3010]) );
  AN2D0 U4629 ( .A1(a[9]), .A2(n[1983]), .Z(n[3007]) );
  AN2D0 U4630 ( .A1(a[9]), .A2(n[1982]), .Z(n[3006]) );
  AN2D0 U4631 ( .A1(a[9]), .A2(n[1979]), .Z(n[3003]) );
  AN2D0 U4632 ( .A1(a[9]), .A2(n[1976]), .Z(n[3000]) );
  AN2D0 U4633 ( .A1(a[9]), .A2(n[1975]), .Z(n[2999]) );
  AN2D0 U4634 ( .A1(a[9]), .A2(n[1974]), .Z(n[2998]) );
  AN2D0 U4635 ( .A1(a[9]), .A2(n[1973]), .Z(n[2997]) );
  AN2D0 U4636 ( .A1(a[9]), .A2(n[1972]), .Z(n[2996]) );
  AN2D0 U4637 ( .A1(a[9]), .A2(n[1969]), .Z(n[2993]) );
  AN2D0 U4638 ( .A1(a[9]), .A2(n[1966]), .Z(n[2990]) );
  AN2D0 U4639 ( .A1(a[9]), .A2(n[1965]), .Z(n[2989]) );
  AN2D0 U4640 ( .A1(a[9]), .A2(n[1962]), .Z(n[2986]) );
  AN2D0 U4641 ( .A1(a[9]), .A2(n[1959]), .Z(n[2983]) );
  AN2D0 U4642 ( .A1(a[9]), .A2(n[1958]), .Z(n[2982]) );
  AN2D0 U4643 ( .A1(a[9]), .A2(n[1957]), .Z(n[2981]) );
  AN2D0 U4644 ( .A1(a[9]), .A2(n[1954]), .Z(n[2978]) );
  AN2D0 U4645 ( .A1(a[9]), .A2(n[1951]), .Z(n[2975]) );
  AN2D0 U4646 ( .A1(a[9]), .A2(n[1950]), .Z(n[2974]) );
  AN2D0 U4647 ( .A1(a[9]), .A2(n[1947]), .Z(n[2971]) );
  AN2D0 U4648 ( .A1(a[9]), .A2(n[1944]), .Z(n[2968]) );
  AN2D0 U4649 ( .A1(a[9]), .A2(n[1943]), .Z(n[2967]) );
  AN2D0 U4650 ( .A1(a[9]), .A2(n[1942]), .Z(n[2966]) );
  AN2D0 U4651 ( .A1(a[9]), .A2(n[1941]), .Z(n[2965]) );
  AN2D0 U4652 ( .A1(a[9]), .A2(n[1938]), .Z(n[2962]) );
  AN2D0 U4653 ( .A1(a[9]), .A2(n[1935]), .Z(n[2959]) );
  AN2D0 U4654 ( .A1(a[9]), .A2(n[1934]), .Z(n[2958]) );
  AN2D0 U4655 ( .A1(a[9]), .A2(n[1931]), .Z(n[2955]) );
  AN2D0 U4656 ( .A1(a[9]), .A2(n[1928]), .Z(n[2952]) );
  AN2D0 U4657 ( .A1(a[9]), .A2(n[1927]), .Z(n[2951]) );
  AN2D0 U4658 ( .A1(a[9]), .A2(n[1926]), .Z(n[2950]) );
  AN2D0 U4659 ( .A1(a[9]), .A2(n[1923]), .Z(n[2947]) );
  AN2D0 U4660 ( .A1(a[9]), .A2(n[1920]), .Z(n[2944]) );
  AN2D0 U4661 ( .A1(a[9]), .A2(n[1919]), .Z(n[2943]) );
  AN2D0 U4662 ( .A1(a[9]), .A2(n[1916]), .Z(n[2940]) );
  AN2D0 U4663 ( .A1(a[9]), .A2(n[1913]), .Z(n[2937]) );
  AN2D0 U4664 ( .A1(a[9]), .A2(n[1912]), .Z(n[2936]) );
  AN2D0 U4665 ( .A1(a[9]), .A2(n[1911]), .Z(n[2935]) );
  AN2D0 U4666 ( .A1(a[9]), .A2(n[1910]), .Z(n[2934]) );
  AN2D0 U4667 ( .A1(a[9]), .A2(n[1909]), .Z(n[2933]) );
  AN2D0 U4668 ( .A1(a[9]), .A2(n[1908]), .Z(n[2932]) );
  AN2D0 U4669 ( .A1(a[9]), .A2(n[1905]), .Z(n[2929]) );
  AN2D0 U4670 ( .A1(a[9]), .A2(n[1902]), .Z(n[2926]) );
  AN2D0 U4671 ( .A1(a[9]), .A2(n[1901]), .Z(n[2925]) );
  AN2D0 U4672 ( .A1(a[9]), .A2(n[1898]), .Z(n[2922]) );
  AN2D0 U4673 ( .A1(a[9]), .A2(n[1895]), .Z(n[2919]) );
  AN2D0 U4674 ( .A1(a[9]), .A2(n[1894]), .Z(n[2918]) );
  AN2D0 U4675 ( .A1(a[9]), .A2(n[1893]), .Z(n[2917]) );
  AN2D0 U4676 ( .A1(a[9]), .A2(n[1890]), .Z(n[2914]) );
  AN2D0 U4677 ( .A1(a[9]), .A2(n[1887]), .Z(n[2911]) );
  AN2D0 U4678 ( .A1(a[9]), .A2(n[1886]), .Z(n[2910]) );
  AN2D0 U4679 ( .A1(a[9]), .A2(n[1883]), .Z(n[2907]) );
  AN2D0 U4680 ( .A1(a[9]), .A2(n[1880]), .Z(n[2904]) );
  AN2D0 U4681 ( .A1(a[9]), .A2(n[1879]), .Z(n[2903]) );
  AN2D0 U4682 ( .A1(a[9]), .A2(n[1878]), .Z(n[2902]) );
  AN2D0 U4683 ( .A1(a[9]), .A2(n[1877]), .Z(n[2901]) );
  AN2D0 U4684 ( .A1(a[9]), .A2(n[1874]), .Z(n[2898]) );
  AN2D0 U4685 ( .A1(a[9]), .A2(n[1871]), .Z(n[2895]) );
  AN2D0 U4686 ( .A1(a[9]), .A2(n[1870]), .Z(n[2894]) );
  AN2D0 U4687 ( .A1(a[9]), .A2(n[1867]), .Z(n[2891]) );
  AN2D0 U4688 ( .A1(a[9]), .A2(n[1864]), .Z(n[2888]) );
  AN2D0 U4689 ( .A1(a[9]), .A2(n[1863]), .Z(n[2887]) );
  AN2D0 U4690 ( .A1(a[9]), .A2(n[1862]), .Z(n[2886]) );
  AN2D0 U4691 ( .A1(a[9]), .A2(n[1859]), .Z(n[2883]) );
  AN2D0 U4692 ( .A1(a[9]), .A2(n[1856]), .Z(n[2880]) );
  AN2D0 U4693 ( .A1(a[9]), .A2(n[1855]), .Z(n[2879]) );
  AN2D0 U4694 ( .A1(a[9]), .A2(n[1852]), .Z(n[2876]) );
  AN2D0 U4695 ( .A1(a[9]), .A2(n[1849]), .Z(n[2873]) );
  AN2D0 U4696 ( .A1(a[9]), .A2(n[1848]), .Z(n[2872]) );
  AN2D0 U4697 ( .A1(a[9]), .A2(n[1847]), .Z(n[2871]) );
  AN2D0 U4698 ( .A1(a[9]), .A2(n[1846]), .Z(n[2870]) );
  AN2D0 U4699 ( .A1(a[9]), .A2(n[1845]), .Z(n[2869]) );
  AN2D0 U4700 ( .A1(a[9]), .A2(n[1842]), .Z(n[2866]) );
  AN2D0 U4701 ( .A1(a[9]), .A2(n[1839]), .Z(n[2863]) );
  AN2D0 U4702 ( .A1(a[9]), .A2(n[1838]), .Z(n[2862]) );
  AN2D0 U4703 ( .A1(a[9]), .A2(n[1835]), .Z(n[2859]) );
  AN2D0 U4704 ( .A1(a[9]), .A2(n[1832]), .Z(n[2856]) );
  AN2D0 U4705 ( .A1(a[9]), .A2(n[1831]), .Z(n[2855]) );
  AN2D0 U4706 ( .A1(a[9]), .A2(n[1830]), .Z(n[2854]) );
  AN2D0 U4707 ( .A1(a[9]), .A2(n[1827]), .Z(n[2851]) );
  AN2D0 U4708 ( .A1(a[9]), .A2(n[1824]), .Z(n[2848]) );
  AN2D0 U4709 ( .A1(a[9]), .A2(n[1823]), .Z(n[2847]) );
  AN2D0 U4710 ( .A1(a[9]), .A2(n[1820]), .Z(n[2844]) );
  AN2D0 U4711 ( .A1(a[9]), .A2(n[1817]), .Z(n[2841]) );
  AN2D0 U4712 ( .A1(a[9]), .A2(n[1816]), .Z(n[2840]) );
  AN2D0 U4713 ( .A1(a[9]), .A2(n[1815]), .Z(n[2839]) );
  AN2D0 U4714 ( .A1(a[9]), .A2(n[1814]), .Z(n[2838]) );
  AN2D0 U4715 ( .A1(a[9]), .A2(n[1811]), .Z(n[2835]) );
  AN2D0 U4716 ( .A1(a[9]), .A2(n[1808]), .Z(n[2832]) );
  AN2D0 U4717 ( .A1(a[9]), .A2(n[1807]), .Z(n[2831]) );
  AN2D0 U4718 ( .A1(a[9]), .A2(n[1804]), .Z(n[2828]) );
  AN2D0 U4719 ( .A1(a[9]), .A2(n[1801]), .Z(n[2825]) );
  AN2D0 U4720 ( .A1(a[9]), .A2(n[1800]), .Z(n[2824]) );
  AN2D0 U4721 ( .A1(a[9]), .A2(n[1799]), .Z(n[2823]) );
  AN2D0 U4722 ( .A1(a[9]), .A2(n[1796]), .Z(n[2820]) );
  AN2D0 U4723 ( .A1(a[9]), .A2(n[1793]), .Z(n[2817]) );
  AN2D0 U4724 ( .A1(a[9]), .A2(n[1792]), .Z(n[2816]) );
  AN2D0 U4725 ( .A1(a[9]), .A2(n[1789]), .Z(n[2813]) );
  AN2D0 U4726 ( .A1(a[9]), .A2(n[1786]), .Z(n[2810]) );
  AN2D0 U4727 ( .A1(a[9]), .A2(n[1785]), .Z(n[2809]) );
  AN2D0 U4728 ( .A1(a[9]), .A2(n[1784]), .Z(n[2808]) );
  AN2D0 U4729 ( .A1(a[9]), .A2(n[1783]), .Z(n[2807]) );
  AN2D0 U4730 ( .A1(a[9]), .A2(n[1782]), .Z(n[2806]) );
  AN2D0 U4731 ( .A1(a[9]), .A2(n[1781]), .Z(n[2805]) );
  AN2D0 U4732 ( .A1(a[9]), .A2(n[1780]), .Z(n[2804]) );
  AN2D0 U4733 ( .A1(a[9]), .A2(n[1777]), .Z(n[2801]) );
  AN2D0 U4734 ( .A1(a[9]), .A2(n[1774]), .Z(n[2798]) );
  AN2D0 U4735 ( .A1(a[9]), .A2(n[1773]), .Z(n[2797]) );
  AN2D0 U4736 ( .A1(a[9]), .A2(n[1770]), .Z(n[2794]) );
  AN2D0 U4737 ( .A1(a[9]), .A2(n[1767]), .Z(n[2791]) );
  AN2D0 U4738 ( .A1(a[9]), .A2(n[1766]), .Z(n[2790]) );
  AN2D0 U4739 ( .A1(a[9]), .A2(n[1765]), .Z(n[2789]) );
  AN2D0 U4740 ( .A1(a[9]), .A2(n[1762]), .Z(n[2786]) );
  AN2D0 U4741 ( .A1(a[9]), .A2(n[1759]), .Z(n[2783]) );
  AN2D0 U4742 ( .A1(a[9]), .A2(n[1758]), .Z(n[2782]) );
  AN2D0 U4743 ( .A1(a[9]), .A2(n[1755]), .Z(n[2779]) );
  AN2D0 U4744 ( .A1(a[9]), .A2(n[1752]), .Z(n[2776]) );
  AN2D0 U4745 ( .A1(a[9]), .A2(n[1751]), .Z(n[2775]) );
  AN2D0 U4746 ( .A1(a[9]), .A2(n[1750]), .Z(n[2774]) );
  AN2D0 U4747 ( .A1(a[9]), .A2(n[1749]), .Z(n[2773]) );
  AN2D0 U4748 ( .A1(a[9]), .A2(n[1746]), .Z(n[2770]) );
  AN2D0 U4749 ( .A1(a[9]), .A2(n[1743]), .Z(n[2767]) );
  AN2D0 U4750 ( .A1(a[9]), .A2(n[1742]), .Z(n[2766]) );
  AN2D0 U4751 ( .A1(a[9]), .A2(n[1739]), .Z(n[2763]) );
  AN2D0 U4752 ( .A1(a[9]), .A2(n[1736]), .Z(n[2760]) );
  AN2D0 U4753 ( .A1(a[9]), .A2(n[1735]), .Z(n[2759]) );
  AN2D0 U4754 ( .A1(a[9]), .A2(n[1734]), .Z(n[2758]) );
  AN2D0 U4755 ( .A1(a[9]), .A2(n[1731]), .Z(n[2755]) );
  AN2D0 U4756 ( .A1(a[9]), .A2(n[1728]), .Z(n[2752]) );
  AN2D0 U4757 ( .A1(a[9]), .A2(n[1727]), .Z(n[2751]) );
  AN2D0 U4758 ( .A1(a[9]), .A2(n[1724]), .Z(n[2748]) );
  AN2D0 U4759 ( .A1(a[9]), .A2(n[1721]), .Z(n[2745]) );
  AN2D0 U4760 ( .A1(a[9]), .A2(n[1720]), .Z(n[2744]) );
  AN2D0 U4761 ( .A1(a[9]), .A2(n[1719]), .Z(n[2743]) );
  AN2D0 U4762 ( .A1(a[9]), .A2(n[1718]), .Z(n[2742]) );
  AN2D0 U4763 ( .A1(a[9]), .A2(n[1717]), .Z(n[2741]) );
  AN2D0 U4764 ( .A1(a[9]), .A2(n[1714]), .Z(n[2738]) );
  AN2D0 U4765 ( .A1(a[9]), .A2(n[1711]), .Z(n[2735]) );
  AN2D0 U4766 ( .A1(a[9]), .A2(n[1710]), .Z(n[2734]) );
  AN2D0 U4767 ( .A1(a[9]), .A2(n[1707]), .Z(n[2731]) );
  AN2D0 U4768 ( .A1(a[9]), .A2(n[1704]), .Z(n[2728]) );
  AN2D0 U4769 ( .A1(a[9]), .A2(n[1703]), .Z(n[2727]) );
  AN2D0 U4770 ( .A1(a[9]), .A2(n[1702]), .Z(n[2726]) );
  AN2D0 U4771 ( .A1(a[9]), .A2(n[1699]), .Z(n[2723]) );
  AN2D0 U4772 ( .A1(a[9]), .A2(n[1696]), .Z(n[2720]) );
  AN2D0 U4773 ( .A1(a[9]), .A2(n[1695]), .Z(n[2719]) );
  AN2D0 U4774 ( .A1(a[9]), .A2(n[1692]), .Z(n[2716]) );
  AN2D0 U4775 ( .A1(a[9]), .A2(n[1689]), .Z(n[2713]) );
  AN2D0 U4776 ( .A1(a[9]), .A2(n[1688]), .Z(n[2712]) );
  AN2D0 U4777 ( .A1(a[9]), .A2(n[1687]), .Z(n[2711]) );
  AN2D0 U4778 ( .A1(a[9]), .A2(n[1686]), .Z(n[2710]) );
  AN2D0 U4779 ( .A1(a[9]), .A2(n[1683]), .Z(n[2707]) );
  AN2D0 U4780 ( .A1(a[9]), .A2(n[1680]), .Z(n[2704]) );
  AN2D0 U4781 ( .A1(a[9]), .A2(n[1679]), .Z(n[2703]) );
  AN2D0 U4782 ( .A1(a[9]), .A2(n[1676]), .Z(n[2700]) );
  AN2D0 U4783 ( .A1(a[9]), .A2(n[1673]), .Z(n[2697]) );
  AN2D0 U4784 ( .A1(a[9]), .A2(n[1672]), .Z(n[2696]) );
  AN2D0 U4785 ( .A1(a[9]), .A2(n[1671]), .Z(n[2695]) );
  AN2D0 U4786 ( .A1(a[9]), .A2(n[1668]), .Z(n[2692]) );
  AN2D0 U4787 ( .A1(a[9]), .A2(n[1665]), .Z(n[2689]) );
  AN2D0 U4788 ( .A1(a[9]), .A2(n[1664]), .Z(n[2688]) );
  AN2D0 U4789 ( .A1(a[9]), .A2(n[1661]), .Z(n[2685]) );
  AN2D0 U4790 ( .A1(a[9]), .A2(n[1658]), .Z(n[2682]) );
  AN2D0 U4791 ( .A1(a[9]), .A2(n[1657]), .Z(n[2681]) );
  AN2D0 U4792 ( .A1(a[9]), .A2(n[1656]), .Z(n[2680]) );
  AN2D0 U4793 ( .A1(a[9]), .A2(n[1655]), .Z(n[2679]) );
  AN2D0 U4794 ( .A1(a[9]), .A2(n[1654]), .Z(n[2678]) );
  AN2D0 U4795 ( .A1(a[9]), .A2(n[1653]), .Z(n[2677]) );
  AN2D0 U4796 ( .A1(a[9]), .A2(n[1650]), .Z(n[2674]) );
  AN2D0 U4797 ( .A1(a[9]), .A2(n[1647]), .Z(n[2671]) );
  AN2D0 U4798 ( .A1(a[9]), .A2(n[1646]), .Z(n[2670]) );
  AN2D0 U4799 ( .A1(a[9]), .A2(n[1643]), .Z(n[2667]) );
  AN2D0 U4800 ( .A1(a[9]), .A2(n[1640]), .Z(n[2664]) );
  AN2D0 U4801 ( .A1(a[9]), .A2(n[1639]), .Z(n[2663]) );
  AN2D0 U4802 ( .A1(a[9]), .A2(n[1638]), .Z(n[2662]) );
  AN2D0 U4803 ( .A1(a[9]), .A2(n[1635]), .Z(n[2659]) );
  AN2D0 U4804 ( .A1(a[9]), .A2(n[1632]), .Z(n[2656]) );
  AN2D0 U4805 ( .A1(a[9]), .A2(n[1631]), .Z(n[2655]) );
  AN2D0 U4806 ( .A1(a[9]), .A2(n[1628]), .Z(n[2652]) );
  AN2D0 U4807 ( .A1(a[9]), .A2(n[1625]), .Z(n[2649]) );
  AN2D0 U4808 ( .A1(a[9]), .A2(n[1624]), .Z(n[2648]) );
  AN2D0 U4809 ( .A1(a[9]), .A2(n[1623]), .Z(n[2647]) );
  AN2D0 U4810 ( .A1(a[9]), .A2(n[1622]), .Z(n[2646]) );
  AN2D0 U4811 ( .A1(a[9]), .A2(n[1619]), .Z(n[2643]) );
  AN2D0 U4812 ( .A1(a[9]), .A2(n[1616]), .Z(n[2640]) );
  AN2D0 U4813 ( .A1(a[9]), .A2(n[1615]), .Z(n[2639]) );
  AN2D0 U4814 ( .A1(a[9]), .A2(n[1612]), .Z(n[2636]) );
  AN2D0 U4815 ( .A1(a[9]), .A2(n[1609]), .Z(n[2633]) );
  AN2D0 U4816 ( .A1(a[9]), .A2(n[1608]), .Z(n[2632]) );
  AN2D0 U4817 ( .A1(a[9]), .A2(n[1607]), .Z(n[2631]) );
  AN2D0 U4818 ( .A1(a[9]), .A2(n[1604]), .Z(n[2628]) );
  AN2D0 U4819 ( .A1(a[9]), .A2(n[1601]), .Z(n[2625]) );
  AN2D0 U4820 ( .A1(a[9]), .A2(n[1600]), .Z(n[2624]) );
  AN2D0 U4821 ( .A1(a[9]), .A2(n[1597]), .Z(n[2621]) );
  AN2D0 U4822 ( .A1(a[9]), .A2(n[1594]), .Z(n[2618]) );
  AN2D0 U4823 ( .A1(a[9]), .A2(n[1593]), .Z(n[2617]) );
  AN2D0 U4824 ( .A1(a[9]), .A2(n[1592]), .Z(n[2616]) );
  AN2D0 U4825 ( .A1(a[9]), .A2(n[1591]), .Z(n[2615]) );
  AN2D0 U4826 ( .A1(a[9]), .A2(n[1590]), .Z(n[2614]) );
  AN2D0 U4827 ( .A1(a[9]), .A2(n[1587]), .Z(n[2611]) );
  AN2D0 U4828 ( .A1(a[9]), .A2(n[1584]), .Z(n[2608]) );
  AN2D0 U4829 ( .A1(a[9]), .A2(n[1583]), .Z(n[2607]) );
  AN2D0 U4830 ( .A1(a[9]), .A2(n[1580]), .Z(n[2604]) );
  AN2D0 U4831 ( .A1(a[9]), .A2(n[1577]), .Z(n[2601]) );
  AN2D0 U4832 ( .A1(a[9]), .A2(n[1576]), .Z(n[2600]) );
  AN2D0 U4833 ( .A1(a[9]), .A2(n[1575]), .Z(n[2599]) );
  AN2D0 U4834 ( .A1(a[9]), .A2(n[1572]), .Z(n[2596]) );
  AN2D0 U4835 ( .A1(a[9]), .A2(n[1569]), .Z(n[2593]) );
  AN2D0 U4836 ( .A1(a[9]), .A2(n[1568]), .Z(n[2592]) );
  AN2D0 U4837 ( .A1(a[9]), .A2(n[1565]), .Z(n[2589]) );
  AN2D0 U4838 ( .A1(a[9]), .A2(n[1562]), .Z(n[2586]) );
  AN2D0 U4839 ( .A1(a[9]), .A2(n[1561]), .Z(n[2585]) );
  AN2D0 U4840 ( .A1(a[9]), .A2(n[1560]), .Z(n[2584]) );
  AN2D0 U4841 ( .A1(a[9]), .A2(n[1559]), .Z(n[2583]) );
  AN2D0 U4842 ( .A1(a[9]), .A2(n[1556]), .Z(n[2580]) );
  AN2D0 U4843 ( .A1(a[9]), .A2(n[1553]), .Z(n[2577]) );
  AN2D0 U4844 ( .A1(a[9]), .A2(n[1552]), .Z(n[2576]) );
  AN2D0 U4845 ( .A1(a[9]), .A2(n[1549]), .Z(n[2573]) );
  AN2D0 U4846 ( .A1(a[9]), .A2(n[1546]), .Z(n[2570]) );
  AN2D0 U4847 ( .A1(a[9]), .A2(n[1545]), .Z(n[2569]) );
  AN2D0 U4848 ( .A1(a[9]), .A2(n[1544]), .Z(n[2568]) );
  AN2D0 U4849 ( .A1(a[9]), .A2(n[1541]), .Z(n[2565]) );
  AN2D0 U4850 ( .A1(a[9]), .A2(n[1538]), .Z(n[2562]) );
  AN2D0 U4851 ( .A1(a[9]), .A2(n[1537]), .Z(n[2561]) );
  AN2D0 U4852 ( .A1(a[9]), .A2(n[1534]), .Z(n[2558]) );
  AN2D0 U4853 ( .A1(a[9]), .A2(n[1531]), .Z(n[2555]) );
  AN2D0 U4854 ( .A1(a[9]), .A2(n[1530]), .Z(n[2554]) );
  AN2D0 U4855 ( .A1(a[9]), .A2(n[1529]), .Z(n[2553]) );
  AN2D0 U4856 ( .A1(a[9]), .A2(n[1528]), .Z(n[2552]) );
  AN2D0 U4857 ( .A1(a[9]), .A2(n[1527]), .Z(n[2551]) );
  AN2D0 U4858 ( .A1(a[9]), .A2(n[1526]), .Z(n[2550]) );
  AN2D0 U4859 ( .A1(a[9]), .A2(n[1525]), .Z(n[2549]) );
  AN2D0 U4860 ( .A1(a[9]), .A2(n[1524]), .Z(n[2548]) );
  AN2D0 U4861 ( .A1(a[9]), .A2(n[1521]), .Z(n[2545]) );
  AN2D0 U4862 ( .A1(a[9]), .A2(n[1518]), .Z(n[2542]) );
  AN2D0 U4863 ( .A1(a[9]), .A2(n[1517]), .Z(n[2541]) );
  AN2D0 U4864 ( .A1(a[9]), .A2(n[1514]), .Z(n[2538]) );
  AN2D0 U4865 ( .A1(a[9]), .A2(n[1511]), .Z(n[2535]) );
  AN2D0 U4866 ( .A1(a[9]), .A2(n[1510]), .Z(n[2534]) );
  AN2D0 U4867 ( .A1(a[9]), .A2(n[1509]), .Z(n[2533]) );
  AN2D0 U4868 ( .A1(a[9]), .A2(n[1506]), .Z(n[2530]) );
  AN2D0 U4869 ( .A1(a[9]), .A2(n[1503]), .Z(n[2527]) );
  AN2D0 U4870 ( .A1(a[9]), .A2(n[1502]), .Z(n[2526]) );
  AN2D0 U4871 ( .A1(a[9]), .A2(n[1499]), .Z(n[2523]) );
  AN2D0 U4872 ( .A1(a[9]), .A2(n[1496]), .Z(n[2520]) );
  AN2D0 U4873 ( .A1(a[9]), .A2(n[1495]), .Z(n[2519]) );
  AN2D0 U4874 ( .A1(a[9]), .A2(n[1494]), .Z(n[2518]) );
  AN2D0 U4875 ( .A1(a[9]), .A2(n[1493]), .Z(n[2517]) );
  AN2D0 U4876 ( .A1(a[9]), .A2(n[1490]), .Z(n[2514]) );
  AN2D0 U4877 ( .A1(a[9]), .A2(n[1487]), .Z(n[2511]) );
  AN2D0 U4878 ( .A1(a[9]), .A2(n[1486]), .Z(n[2510]) );
  AN2D0 U4879 ( .A1(a[9]), .A2(n[1483]), .Z(n[2507]) );
  AN2D0 U4880 ( .A1(a[9]), .A2(n[1480]), .Z(n[2504]) );
  AN2D0 U4881 ( .A1(a[9]), .A2(n[1479]), .Z(n[2503]) );
  AN2D0 U4882 ( .A1(a[9]), .A2(n[1478]), .Z(n[2502]) );
  AN2D0 U4883 ( .A1(a[9]), .A2(n[1475]), .Z(n[2499]) );
  AN2D0 U4884 ( .A1(a[9]), .A2(n[1472]), .Z(n[2496]) );
  AN2D0 U4885 ( .A1(a[9]), .A2(n[1471]), .Z(n[2495]) );
  AN2D0 U4886 ( .A1(a[9]), .A2(n[1468]), .Z(n[2492]) );
  AN2D0 U4887 ( .A1(a[9]), .A2(n[1465]), .Z(n[2489]) );
  AN2D0 U4888 ( .A1(a[9]), .A2(n[1464]), .Z(n[2488]) );
  AN2D0 U4889 ( .A1(a[9]), .A2(n[1463]), .Z(n[2487]) );
  AN2D0 U4890 ( .A1(a[9]), .A2(n[1462]), .Z(n[2486]) );
  AN2D0 U4891 ( .A1(a[9]), .A2(n[1461]), .Z(n[2485]) );
  AN2D0 U4892 ( .A1(a[9]), .A2(n[1458]), .Z(n[2482]) );
  AN2D0 U4893 ( .A1(a[9]), .A2(n[1455]), .Z(n[2479]) );
  AN2D0 U4894 ( .A1(a[9]), .A2(n[1454]), .Z(n[2478]) );
  AN2D0 U4895 ( .A1(a[9]), .A2(n[1451]), .Z(n[2475]) );
  AN2D0 U4896 ( .A1(a[9]), .A2(n[1448]), .Z(n[2472]) );
  AN2D0 U4897 ( .A1(a[9]), .A2(n[1447]), .Z(n[2471]) );
  AN2D0 U4898 ( .A1(a[9]), .A2(n[1446]), .Z(n[2470]) );
  AN2D0 U4899 ( .A1(a[9]), .A2(n[1443]), .Z(n[2467]) );
  AN2D0 U4900 ( .A1(a[9]), .A2(n[1440]), .Z(n[2464]) );
  AN2D0 U4901 ( .A1(a[9]), .A2(n[1439]), .Z(n[2463]) );
  AN2D0 U4902 ( .A1(a[9]), .A2(n[1436]), .Z(n[2460]) );
  AN2D0 U4903 ( .A1(a[9]), .A2(n[1433]), .Z(n[2457]) );
  AN2D0 U4904 ( .A1(a[9]), .A2(n[1432]), .Z(n[2456]) );
  AN2D0 U4905 ( .A1(a[9]), .A2(n[1431]), .Z(n[2455]) );
  AN2D0 U4906 ( .A1(a[9]), .A2(n[1430]), .Z(n[2454]) );
  AN2D0 U4907 ( .A1(a[9]), .A2(n[1427]), .Z(n[2451]) );
  AN2D0 U4908 ( .A1(a[9]), .A2(n[1424]), .Z(n[2448]) );
  AN2D0 U4909 ( .A1(a[9]), .A2(n[1423]), .Z(n[2447]) );
  AN2D0 U4910 ( .A1(a[9]), .A2(n[1420]), .Z(n[2444]) );
  AN2D0 U4911 ( .A1(a[9]), .A2(n[1417]), .Z(n[2441]) );
  AN2D0 U4912 ( .A1(a[9]), .A2(n[1416]), .Z(n[2440]) );
  AN2D0 U4913 ( .A1(a[9]), .A2(n[1415]), .Z(n[2439]) );
  AN2D0 U4914 ( .A1(a[9]), .A2(n[1412]), .Z(n[2436]) );
  AN2D0 U4915 ( .A1(a[9]), .A2(n[1409]), .Z(n[2433]) );
  AN2D0 U4916 ( .A1(a[9]), .A2(n[1408]), .Z(n[2432]) );
  AN2D0 U4917 ( .A1(a[9]), .A2(n[1405]), .Z(n[2429]) );
  AN2D0 U4918 ( .A1(a[9]), .A2(n[1402]), .Z(n[2426]) );
  AN2D0 U4919 ( .A1(a[9]), .A2(n[1401]), .Z(n[2425]) );
  AN2D0 U4920 ( .A1(a[9]), .A2(n[1400]), .Z(n[2424]) );
  AN2D0 U4921 ( .A1(a[9]), .A2(n[1399]), .Z(n[2423]) );
  AN2D0 U4922 ( .A1(a[9]), .A2(n[1398]), .Z(n[2422]) );
  AN2D0 U4923 ( .A1(a[9]), .A2(n[1397]), .Z(n[2421]) );
  AN2D0 U4924 ( .A1(a[9]), .A2(n[1394]), .Z(n[2418]) );
  AN2D0 U4925 ( .A1(a[9]), .A2(n[1391]), .Z(n[2415]) );
  AN2D0 U4926 ( .A1(a[9]), .A2(n[1390]), .Z(n[2414]) );
  AN2D0 U4927 ( .A1(a[9]), .A2(n[1387]), .Z(n[2411]) );
  AN2D0 U4928 ( .A1(a[9]), .A2(n[1384]), .Z(n[2408]) );
  AN2D0 U4929 ( .A1(a[9]), .A2(n[1383]), .Z(n[2407]) );
  AN2D0 U4930 ( .A1(a[9]), .A2(n[1382]), .Z(n[2406]) );
  AN2D0 U4931 ( .A1(a[9]), .A2(n[1379]), .Z(n[2403]) );
  AN2D0 U4932 ( .A1(a[9]), .A2(n[1376]), .Z(n[2400]) );
  AN2D0 U4933 ( .A1(a[9]), .A2(n[1375]), .Z(n[2399]) );
  AN2D0 U4934 ( .A1(a[9]), .A2(n[1372]), .Z(n[2396]) );
  AN2D0 U4935 ( .A1(a[9]), .A2(n[1369]), .Z(n[2393]) );
  AN2D0 U4936 ( .A1(a[9]), .A2(n[1368]), .Z(n[2392]) );
  AN2D0 U4937 ( .A1(a[9]), .A2(n[1367]), .Z(n[2391]) );
  AN2D0 U4938 ( .A1(a[9]), .A2(n[1366]), .Z(n[2390]) );
  AN2D0 U4939 ( .A1(a[9]), .A2(n[1363]), .Z(n[2387]) );
  AN2D0 U4940 ( .A1(a[9]), .A2(n[1360]), .Z(n[2384]) );
  AN2D0 U4941 ( .A1(a[9]), .A2(n[1359]), .Z(n[2383]) );
  AN2D0 U4942 ( .A1(a[9]), .A2(n[1356]), .Z(n[2380]) );
  AN2D0 U4943 ( .A1(a[9]), .A2(n[1353]), .Z(n[2377]) );
  AN2D0 U4944 ( .A1(a[9]), .A2(n[1352]), .Z(n[2376]) );
  AN2D0 U4945 ( .A1(a[9]), .A2(n[1351]), .Z(n[2375]) );
  AN2D0 U4946 ( .A1(a[9]), .A2(n[1348]), .Z(n[2372]) );
  AN2D0 U4947 ( .A1(a[9]), .A2(n[1345]), .Z(n[2369]) );
  AN2D0 U4948 ( .A1(a[9]), .A2(n[1344]), .Z(n[2368]) );
  AN2D0 U4949 ( .A1(a[9]), .A2(n[1341]), .Z(n[2365]) );
  AN2D0 U4950 ( .A1(a[9]), .A2(n[1338]), .Z(n[2362]) );
  AN2D0 U4951 ( .A1(a[9]), .A2(n[1337]), .Z(n[2361]) );
  AN2D0 U4952 ( .A1(a[9]), .A2(n[1336]), .Z(n[2360]) );
  AN2D0 U4953 ( .A1(a[9]), .A2(n[1335]), .Z(n[2359]) );
  AN2D0 U4954 ( .A1(a[9]), .A2(n[1334]), .Z(n[2358]) );
  AN2D0 U4955 ( .A1(a[9]), .A2(n[1331]), .Z(n[2355]) );
  AN2D0 U4956 ( .A1(a[9]), .A2(n[1328]), .Z(n[2352]) );
  AN2D0 U4957 ( .A1(a[9]), .A2(n[1327]), .Z(n[2351]) );
  AN2D0 U4958 ( .A1(a[9]), .A2(n[1324]), .Z(n[2348]) );
  AN2D0 U4959 ( .A1(a[9]), .A2(n[1321]), .Z(n[2345]) );
  AN2D0 U4960 ( .A1(a[9]), .A2(n[1320]), .Z(n[2344]) );
  AN2D0 U4961 ( .A1(a[9]), .A2(n[1319]), .Z(n[2343]) );
  AN2D0 U4962 ( .A1(a[9]), .A2(n[1316]), .Z(n[2340]) );
  AN2D0 U4963 ( .A1(a[9]), .A2(n[1313]), .Z(n[2337]) );
  AN2D0 U4964 ( .A1(a[9]), .A2(n[1312]), .Z(n[2336]) );
  AN2D0 U4965 ( .A1(a[9]), .A2(n[1309]), .Z(n[2333]) );
  AN2D0 U4966 ( .A1(a[9]), .A2(n[1306]), .Z(n[2330]) );
  AN2D0 U4967 ( .A1(a[9]), .A2(n[1305]), .Z(n[2329]) );
  AN2D0 U4968 ( .A1(a[9]), .A2(n[1304]), .Z(n[2328]) );
  AN2D0 U4969 ( .A1(a[9]), .A2(n[1303]), .Z(n[2327]) );
  AN2D0 U4970 ( .A1(a[9]), .A2(n[1300]), .Z(n[2324]) );
  AN2D0 U4971 ( .A1(a[9]), .A2(n[1297]), .Z(n[2321]) );
  AN2D0 U4972 ( .A1(a[9]), .A2(n[1296]), .Z(n[2320]) );
  AN2D0 U4973 ( .A1(a[9]), .A2(n[1293]), .Z(n[2317]) );
  AN2D0 U4974 ( .A1(a[9]), .A2(n[1290]), .Z(n[2314]) );
  AN2D0 U4975 ( .A1(a[9]), .A2(n[1289]), .Z(n[2313]) );
  AN2D0 U4976 ( .A1(a[9]), .A2(n[1288]), .Z(n[2312]) );
  AN2D0 U4977 ( .A1(a[9]), .A2(n[1285]), .Z(n[2309]) );
  AN2D0 U4978 ( .A1(a[9]), .A2(n[1282]), .Z(n[2306]) );
  AN2D0 U4979 ( .A1(a[9]), .A2(n[1281]), .Z(n[2305]) );
  AN2D0 U4980 ( .A1(a[9]), .A2(n[1278]), .Z(n[2302]) );
  AN2D0 U4981 ( .A1(a[9]), .A2(n[1275]), .Z(n[2299]) );
  AN2D0 U4982 ( .A1(a[9]), .A2(n[1274]), .Z(n[2298]) );
  AN2D0 U4983 ( .A1(a[9]), .A2(n[1273]), .Z(n[2297]) );
  AN2D0 U4984 ( .A1(a[9]), .A2(n[1272]), .Z(n[2296]) );
  AN2D0 U4985 ( .A1(a[9]), .A2(n[1271]), .Z(n[2295]) );
  AN2D0 U4986 ( .A1(a[9]), .A2(n[1270]), .Z(n[2294]) );
  AN2D0 U4987 ( .A1(a[9]), .A2(n[1269]), .Z(n[2293]) );
  AN2D0 U4988 ( .A1(a[9]), .A2(n[1266]), .Z(n[2290]) );
  AN2D0 U4989 ( .A1(a[9]), .A2(n[1263]), .Z(n[2287]) );
  AN2D0 U4990 ( .A1(a[9]), .A2(n[1262]), .Z(n[2286]) );
  AN2D0 U4991 ( .A1(a[9]), .A2(n[1259]), .Z(n[2283]) );
  AN2D0 U4992 ( .A1(a[9]), .A2(n[1256]), .Z(n[2280]) );
  AN2D0 U4993 ( .A1(a[9]), .A2(n[1255]), .Z(n[2279]) );
  AN2D0 U4994 ( .A1(a[9]), .A2(n[1254]), .Z(n[2278]) );
  AN2D0 U4995 ( .A1(a[9]), .A2(n[1251]), .Z(n[2275]) );
  AN2D0 U4996 ( .A1(a[9]), .A2(n[1248]), .Z(n[2272]) );
  AN2D0 U4997 ( .A1(a[9]), .A2(n[1247]), .Z(n[2271]) );
  AN2D0 U4998 ( .A1(a[9]), .A2(n[1244]), .Z(n[2268]) );
  AN2D0 U4999 ( .A1(a[9]), .A2(n[1241]), .Z(n[2265]) );
  AN2D0 U5000 ( .A1(a[9]), .A2(n[1240]), .Z(n[2264]) );
  AN2D0 U5001 ( .A1(a[9]), .A2(n[1239]), .Z(n[2263]) );
  AN2D0 U5002 ( .A1(a[9]), .A2(n[1238]), .Z(n[2262]) );
  AN2D0 U5003 ( .A1(a[9]), .A2(n[1235]), .Z(n[2259]) );
  AN2D0 U5004 ( .A1(a[9]), .A2(n[1232]), .Z(n[2256]) );
  AN2D0 U5005 ( .A1(a[9]), .A2(n[1231]), .Z(n[2255]) );
  AN2D0 U5006 ( .A1(a[9]), .A2(n[1228]), .Z(n[2252]) );
  AN2D0 U5007 ( .A1(a[9]), .A2(n[1225]), .Z(n[2249]) );
  AN2D0 U5008 ( .A1(a[9]), .A2(n[1224]), .Z(n[2248]) );
  AN2D0 U5009 ( .A1(a[9]), .A2(n[1223]), .Z(n[2247]) );
  AN2D0 U5010 ( .A1(a[9]), .A2(n[1220]), .Z(n[2244]) );
  AN2D0 U5011 ( .A1(a[9]), .A2(n[1217]), .Z(n[2241]) );
  AN2D0 U5012 ( .A1(a[9]), .A2(n[1216]), .Z(n[2240]) );
  AN2D0 U5013 ( .A1(a[9]), .A2(n[1213]), .Z(n[2237]) );
  AN2D0 U5014 ( .A1(a[9]), .A2(n[1210]), .Z(n[2234]) );
  AN2D0 U5015 ( .A1(a[9]), .A2(n[1209]), .Z(n[2233]) );
  AN2D0 U5016 ( .A1(a[9]), .A2(n[1208]), .Z(n[2232]) );
  AN2D0 U5017 ( .A1(a[9]), .A2(n[1207]), .Z(n[2231]) );
  AN2D0 U5018 ( .A1(a[9]), .A2(n[1206]), .Z(n[2230]) );
  AN2D0 U5019 ( .A1(a[9]), .A2(n[1203]), .Z(n[2227]) );
  AN2D0 U5020 ( .A1(a[9]), .A2(n[1200]), .Z(n[2224]) );
  AN2D0 U5021 ( .A1(a[9]), .A2(n[1199]), .Z(n[2223]) );
  AN2D0 U5022 ( .A1(a[9]), .A2(n[1196]), .Z(n[2220]) );
  AN2D0 U5023 ( .A1(a[9]), .A2(n[1193]), .Z(n[2217]) );
  AN2D0 U5024 ( .A1(a[9]), .A2(n[1192]), .Z(n[2216]) );
  AN2D0 U5025 ( .A1(a[9]), .A2(n[1191]), .Z(n[2215]) );
  AN2D0 U5026 ( .A1(a[9]), .A2(n[1188]), .Z(n[2212]) );
  AN2D0 U5027 ( .A1(a[9]), .A2(n[1185]), .Z(n[2209]) );
  AN2D0 U5028 ( .A1(a[9]), .A2(n[1184]), .Z(n[2208]) );
  AN2D0 U5029 ( .A1(a[9]), .A2(n[1181]), .Z(n[2205]) );
  AN2D0 U5030 ( .A1(a[9]), .A2(n[1178]), .Z(n[2202]) );
  AN2D0 U5031 ( .A1(a[9]), .A2(n[1177]), .Z(n[2201]) );
  AN2D0 U5032 ( .A1(a[9]), .A2(n[1176]), .Z(n[2200]) );
  AN2D0 U5033 ( .A1(a[9]), .A2(n[1175]), .Z(n[2199]) );
  AN2D0 U5034 ( .A1(a[9]), .A2(n[1172]), .Z(n[2196]) );
  AN2D0 U5035 ( .A1(a[9]), .A2(n[1169]), .Z(n[2193]) );
  AN2D0 U5036 ( .A1(a[9]), .A2(n[1168]), .Z(n[2192]) );
  AN2D0 U5037 ( .A1(a[9]), .A2(n[1165]), .Z(n[2189]) );
  AN2D0 U5038 ( .A1(a[9]), .A2(n[1162]), .Z(n[2186]) );
  AN2D0 U5039 ( .A1(a[9]), .A2(n[1161]), .Z(n[2185]) );
  AN2D0 U5040 ( .A1(a[9]), .A2(n[1160]), .Z(n[2184]) );
  AN2D0 U5041 ( .A1(a[9]), .A2(n[1157]), .Z(n[2181]) );
  AN2D0 U5042 ( .A1(a[9]), .A2(n[1154]), .Z(n[2178]) );
  AN2D0 U5043 ( .A1(a[9]), .A2(n[1153]), .Z(n[2177]) );
  AN2D0 U5044 ( .A1(a[9]), .A2(n[1150]), .Z(n[2174]) );
  AN2D0 U5045 ( .A1(a[9]), .A2(n[1147]), .Z(n[2171]) );
  AN2D0 U5046 ( .A1(a[9]), .A2(n[1146]), .Z(n[2170]) );
  AN2D0 U5047 ( .A1(a[9]), .A2(n[1145]), .Z(n[2169]) );
  AN2D0 U5048 ( .A1(a[9]), .A2(n[1144]), .Z(n[2168]) );
  AN2D0 U5049 ( .A1(a[9]), .A2(n[1143]), .Z(n[2167]) );
  AN2D0 U5050 ( .A1(a[9]), .A2(n[1142]), .Z(n[2166]) );
  AN2D0 U5051 ( .A1(a[9]), .A2(n[1139]), .Z(n[2163]) );
  AN2D0 U5052 ( .A1(a[9]), .A2(n[1136]), .Z(n[2160]) );
  AN2D0 U5053 ( .A1(a[9]), .A2(n[1135]), .Z(n[2159]) );
  AN2D0 U5054 ( .A1(a[9]), .A2(n[1132]), .Z(n[2156]) );
  AN2D0 U5055 ( .A1(a[9]), .A2(n[1129]), .Z(n[2153]) );
  AN2D0 U5056 ( .A1(a[9]), .A2(n[1128]), .Z(n[2152]) );
  AN2D0 U5057 ( .A1(a[9]), .A2(n[1127]), .Z(n[2151]) );
  AN2D0 U5058 ( .A1(a[9]), .A2(n[1124]), .Z(n[2148]) );
  AN2D0 U5059 ( .A1(a[9]), .A2(n[1121]), .Z(n[2145]) );
  AN2D0 U5060 ( .A1(a[9]), .A2(n[1120]), .Z(n[2144]) );
  AN2D0 U5061 ( .A1(a[9]), .A2(n[1117]), .Z(n[2141]) );
  AN2D0 U5062 ( .A1(a[9]), .A2(n[1114]), .Z(n[2138]) );
  AN2D0 U5063 ( .A1(a[9]), .A2(n[1113]), .Z(n[2137]) );
  AN2D0 U5064 ( .A1(a[9]), .A2(n[1112]), .Z(n[2136]) );
  AN2D0 U5065 ( .A1(a[9]), .A2(n[1111]), .Z(n[2135]) );
  AN2D0 U5066 ( .A1(a[9]), .A2(n[1108]), .Z(n[2132]) );
  AN2D0 U5067 ( .A1(a[9]), .A2(n[1105]), .Z(n[2129]) );
  AN2D0 U5068 ( .A1(a[9]), .A2(n[1104]), .Z(n[2128]) );
  AN2D0 U5069 ( .A1(a[9]), .A2(n[1101]), .Z(n[2125]) );
  AN2D0 U5070 ( .A1(a[9]), .A2(n[1098]), .Z(n[2122]) );
  AN2D0 U5071 ( .A1(a[9]), .A2(n[1097]), .Z(n[2121]) );
  AN2D0 U5072 ( .A1(a[9]), .A2(n[1096]), .Z(n[2120]) );
  AN2D0 U5073 ( .A1(a[9]), .A2(n[1093]), .Z(n[2117]) );
  AN2D0 U5074 ( .A1(a[9]), .A2(n[1090]), .Z(n[2114]) );
  AN2D0 U5075 ( .A1(a[9]), .A2(n[1089]), .Z(n[2113]) );
  AN2D0 U5076 ( .A1(a[9]), .A2(n[1086]), .Z(n[2110]) );
  AN2D0 U5077 ( .A1(a[9]), .A2(n[1083]), .Z(n[2107]) );
  AN2D0 U5078 ( .A1(a[9]), .A2(n[1082]), .Z(n[2106]) );
  AN2D0 U5079 ( .A1(a[9]), .A2(n[1081]), .Z(n[2105]) );
  AN2D0 U5080 ( .A1(a[9]), .A2(n[1080]), .Z(n[2104]) );
  AN2D0 U5081 ( .A1(a[9]), .A2(n[1079]), .Z(n[2103]) );
  AN2D0 U5082 ( .A1(a[9]), .A2(n[1076]), .Z(n[2100]) );
  AN2D0 U5083 ( .A1(a[9]), .A2(n[1073]), .Z(n[2097]) );
  AN2D0 U5084 ( .A1(a[9]), .A2(n[1072]), .Z(n[2096]) );
  AN2D0 U5085 ( .A1(a[9]), .A2(n[1069]), .Z(n[2093]) );
  AN2D0 U5086 ( .A1(a[9]), .A2(n[1066]), .Z(n[2090]) );
  AN2D0 U5087 ( .A1(a[9]), .A2(n[1065]), .Z(n[2089]) );
  AN2D0 U5088 ( .A1(a[9]), .A2(n[1064]), .Z(n[2088]) );
  AN2D0 U5089 ( .A1(a[9]), .A2(n[1061]), .Z(n[2085]) );
  AN2D0 U5090 ( .A1(a[9]), .A2(n[1058]), .Z(n[2082]) );
  AN2D0 U5091 ( .A1(a[9]), .A2(n[1057]), .Z(n[2081]) );
  AN2D0 U5092 ( .A1(a[9]), .A2(n[1054]), .Z(n[2078]) );
  AN2D0 U5093 ( .A1(a[9]), .A2(n[1051]), .Z(n[2075]) );
  AN2D0 U5094 ( .A1(a[9]), .A2(n[1050]), .Z(n[2074]) );
  AN2D0 U5095 ( .A1(a[9]), .A2(n[1049]), .Z(n[2073]) );
  AN2D0 U5096 ( .A1(a[9]), .A2(n[1048]), .Z(n[2072]) );
  AN2D0 U5097 ( .A1(a[9]), .A2(n[1045]), .Z(n[2069]) );
  AN2D0 U5098 ( .A1(a[9]), .A2(n[1042]), .Z(n[2066]) );
  AN2D0 U5099 ( .A1(a[9]), .A2(n[1041]), .Z(n[2065]) );
  AN2D0 U5100 ( .A1(a[9]), .A2(n[1038]), .Z(n[2062]) );
  AN2D0 U5101 ( .A1(a[9]), .A2(n[1035]), .Z(n[2059]) );
  AN2D0 U5102 ( .A1(a[9]), .A2(n[1034]), .Z(n[2058]) );
  AN2D0 U5103 ( .A1(a[9]), .A2(n[1033]), .Z(n[2057]) );
  AN2D0 U5104 ( .A1(a[9]), .A2(n[1030]), .Z(n[2054]) );
  AN2D0 U5105 ( .A1(a[9]), .A2(n[1027]), .Z(n[2051]) );
  AN2D0 U5106 ( .A1(a[9]), .A2(n[1026]), .Z(n[2050]) );
  AN2D0 U5107 ( .A1(a[9]), .A2(n[1023]), .Z(n[2047]) );
  AN2D0 U5108 ( .A1(a[9]), .A2(n[1020]), .Z(n[2044]) );
  AN2D0 U5109 ( .A1(a[9]), .A2(n[1019]), .Z(n[2043]) );
  AN2D0 U5110 ( .A1(a[9]), .A2(n[1018]), .Z(n[2042]) );
  AN2D0 U5111 ( .A1(a[9]), .A2(n[1017]), .Z(n[2041]) );
  AN2D0 U5112 ( .A1(a[9]), .A2(n[1016]), .Z(n[2040]) );
  AN2D0 U5113 ( .A1(a[9]), .A2(n[1015]), .Z(n[2039]) );
  AN2D0 U5114 ( .A1(a[9]), .A2(n[1014]), .Z(n[2038]) );
  AN2D0 U5115 ( .A1(a[9]), .A2(n[1013]), .Z(n[2037]) );
  AN2D0 U5116 ( .A1(a[9]), .A2(n[1012]), .Z(n[2036]) );
  AN2D0 U5117 ( .A1(a[9]), .A2(b[9]), .Z(n[2035]) );
  AN2D0 U5118 ( .A1(n[1009]), .A2(b[8]), .Z(n[2032]) );
  AN2D0 U5119 ( .A1(b[8]), .A2(n[1006]), .Z(n[2029]) );
  AN2D0 U5120 ( .A1(b[8]), .A2(n[1005]), .Z(n[2028]) );
  AN2D0 U5121 ( .A1(b[8]), .A2(n[1002]), .Z(n[2025]) );
  AN2D0 U5122 ( .A1(b[8]), .A2(n[999]), .Z(n[2022]) );
  AN2D0 U5123 ( .A1(b[8]), .A2(n[998]), .Z(n[2021]) );
  AN2D0 U5124 ( .A1(b[8]), .A2(n[997]), .Z(n[2020]) );
  AN2D0 U5125 ( .A1(b[8]), .A2(n[994]), .Z(n[2017]) );
  AN2D0 U5126 ( .A1(b[8]), .A2(n[991]), .Z(n[2014]) );
  AN2D0 U5127 ( .A1(b[8]), .A2(n[990]), .Z(n[2013]) );
  AN2D0 U5128 ( .A1(b[8]), .A2(n[987]), .Z(n[2010]) );
  AN2D0 U5129 ( .A1(b[8]), .A2(n[984]), .Z(n[2007]) );
  AN2D0 U5130 ( .A1(b[8]), .A2(n[983]), .Z(n[2006]) );
  AN2D0 U5131 ( .A1(b[8]), .A2(n[982]), .Z(n[2005]) );
  AN2D0 U5132 ( .A1(b[8]), .A2(n[981]), .Z(n[2004]) );
  AN2D0 U5133 ( .A1(b[8]), .A2(n[978]), .Z(n[2001]) );
  AN2D0 U5134 ( .A1(b[8]), .A2(n[975]), .Z(n[1998]) );
  AN2D0 U5135 ( .A1(b[8]), .A2(n[974]), .Z(n[1997]) );
  AN2D0 U5136 ( .A1(b[8]), .A2(n[971]), .Z(n[1994]) );
  AN2D0 U5137 ( .A1(b[8]), .A2(n[968]), .Z(n[1991]) );
  AN2D0 U5138 ( .A1(b[8]), .A2(n[967]), .Z(n[1990]) );
  AN2D0 U5139 ( .A1(b[8]), .A2(n[966]), .Z(n[1989]) );
  AN2D0 U5140 ( .A1(b[8]), .A2(n[963]), .Z(n[1986]) );
  AN2D0 U5141 ( .A1(b[8]), .A2(n[960]), .Z(n[1983]) );
  AN2D0 U5142 ( .A1(b[8]), .A2(n[959]), .Z(n[1982]) );
  AN2D0 U5143 ( .A1(b[8]), .A2(n[956]), .Z(n[1979]) );
  AN2D0 U5144 ( .A1(b[8]), .A2(n[953]), .Z(n[1976]) );
  AN2D0 U5145 ( .A1(b[8]), .A2(n[952]), .Z(n[1975]) );
  AN2D0 U5146 ( .A1(b[8]), .A2(n[951]), .Z(n[1974]) );
  AN2D0 U5147 ( .A1(b[8]), .A2(n[950]), .Z(n[1973]) );
  AN2D0 U5148 ( .A1(b[8]), .A2(n[949]), .Z(n[1972]) );
  AN2D0 U5149 ( .A1(b[8]), .A2(n[946]), .Z(n[1969]) );
  AN2D0 U5150 ( .A1(b[8]), .A2(n[943]), .Z(n[1966]) );
  AN2D0 U5151 ( .A1(b[8]), .A2(n[942]), .Z(n[1965]) );
  AN2D0 U5152 ( .A1(b[8]), .A2(n[939]), .Z(n[1962]) );
  AN2D0 U5153 ( .A1(b[8]), .A2(n[936]), .Z(n[1959]) );
  AN2D0 U5154 ( .A1(b[8]), .A2(n[935]), .Z(n[1958]) );
  AN2D0 U5155 ( .A1(b[8]), .A2(n[934]), .Z(n[1957]) );
  AN2D0 U5156 ( .A1(b[8]), .A2(n[931]), .Z(n[1954]) );
  AN2D0 U5157 ( .A1(b[8]), .A2(n[928]), .Z(n[1951]) );
  AN2D0 U5158 ( .A1(b[8]), .A2(n[927]), .Z(n[1950]) );
  AN2D0 U5159 ( .A1(b[8]), .A2(n[924]), .Z(n[1947]) );
  AN2D0 U5160 ( .A1(b[8]), .A2(n[921]), .Z(n[1944]) );
  AN2D0 U5161 ( .A1(b[8]), .A2(n[920]), .Z(n[1943]) );
  AN2D0 U5162 ( .A1(b[8]), .A2(n[919]), .Z(n[1942]) );
  AN2D0 U5163 ( .A1(b[8]), .A2(n[918]), .Z(n[1941]) );
  AN2D0 U5164 ( .A1(b[8]), .A2(n[915]), .Z(n[1938]) );
  AN2D0 U5165 ( .A1(b[8]), .A2(n[912]), .Z(n[1935]) );
  AN2D0 U5166 ( .A1(b[8]), .A2(n[911]), .Z(n[1934]) );
  AN2D0 U5167 ( .A1(b[8]), .A2(n[908]), .Z(n[1931]) );
  AN2D0 U5168 ( .A1(b[8]), .A2(n[905]), .Z(n[1928]) );
  AN2D0 U5169 ( .A1(b[8]), .A2(n[904]), .Z(n[1927]) );
  AN2D0 U5170 ( .A1(b[8]), .A2(n[903]), .Z(n[1926]) );
  AN2D0 U5171 ( .A1(b[8]), .A2(n[900]), .Z(n[1923]) );
  AN2D0 U5172 ( .A1(b[8]), .A2(n[897]), .Z(n[1920]) );
  AN2D0 U5173 ( .A1(b[8]), .A2(n[896]), .Z(n[1919]) );
  AN2D0 U5174 ( .A1(b[8]), .A2(n[893]), .Z(n[1916]) );
  AN2D0 U5175 ( .A1(b[8]), .A2(n[890]), .Z(n[1913]) );
  AN2D0 U5176 ( .A1(b[8]), .A2(n[889]), .Z(n[1912]) );
  AN2D0 U5177 ( .A1(b[8]), .A2(n[888]), .Z(n[1911]) );
  AN2D0 U5178 ( .A1(b[8]), .A2(n[887]), .Z(n[1910]) );
  AN2D0 U5179 ( .A1(b[8]), .A2(n[886]), .Z(n[1909]) );
  AN2D0 U5180 ( .A1(b[8]), .A2(n[885]), .Z(n[1908]) );
  AN2D0 U5181 ( .A1(b[8]), .A2(n[882]), .Z(n[1905]) );
  AN2D0 U5182 ( .A1(b[8]), .A2(n[879]), .Z(n[1902]) );
  AN2D0 U5183 ( .A1(b[8]), .A2(n[878]), .Z(n[1901]) );
  AN2D0 U5184 ( .A1(b[8]), .A2(n[875]), .Z(n[1898]) );
  AN2D0 U5185 ( .A1(b[8]), .A2(n[872]), .Z(n[1895]) );
  AN2D0 U5186 ( .A1(b[8]), .A2(n[871]), .Z(n[1894]) );
  AN2D0 U5187 ( .A1(b[8]), .A2(n[870]), .Z(n[1893]) );
  AN2D0 U5188 ( .A1(b[8]), .A2(n[867]), .Z(n[1890]) );
  AN2D0 U5189 ( .A1(b[8]), .A2(n[864]), .Z(n[1887]) );
  AN2D0 U5190 ( .A1(b[8]), .A2(n[863]), .Z(n[1886]) );
  AN2D0 U5191 ( .A1(b[8]), .A2(n[860]), .Z(n[1883]) );
  AN2D0 U5192 ( .A1(b[8]), .A2(n[857]), .Z(n[1880]) );
  AN2D0 U5193 ( .A1(b[8]), .A2(n[856]), .Z(n[1879]) );
  AN2D0 U5194 ( .A1(b[8]), .A2(n[855]), .Z(n[1878]) );
  AN2D0 U5195 ( .A1(b[8]), .A2(n[854]), .Z(n[1877]) );
  AN2D0 U5196 ( .A1(b[8]), .A2(n[851]), .Z(n[1874]) );
  AN2D0 U5197 ( .A1(b[8]), .A2(n[848]), .Z(n[1871]) );
  AN2D0 U5198 ( .A1(b[8]), .A2(n[847]), .Z(n[1870]) );
  AN2D0 U5199 ( .A1(b[8]), .A2(n[844]), .Z(n[1867]) );
  AN2D0 U5200 ( .A1(b[8]), .A2(n[841]), .Z(n[1864]) );
  AN2D0 U5201 ( .A1(b[8]), .A2(n[840]), .Z(n[1863]) );
  AN2D0 U5202 ( .A1(b[8]), .A2(n[839]), .Z(n[1862]) );
  AN2D0 U5203 ( .A1(b[8]), .A2(n[836]), .Z(n[1859]) );
  AN2D0 U5204 ( .A1(b[8]), .A2(n[833]), .Z(n[1856]) );
  AN2D0 U5205 ( .A1(b[8]), .A2(n[832]), .Z(n[1855]) );
  AN2D0 U5206 ( .A1(b[8]), .A2(n[829]), .Z(n[1852]) );
  AN2D0 U5207 ( .A1(b[8]), .A2(n[826]), .Z(n[1849]) );
  AN2D0 U5208 ( .A1(b[8]), .A2(n[825]), .Z(n[1848]) );
  AN2D0 U5209 ( .A1(b[8]), .A2(n[824]), .Z(n[1847]) );
  AN2D0 U5210 ( .A1(b[8]), .A2(n[823]), .Z(n[1846]) );
  AN2D0 U5211 ( .A1(b[8]), .A2(n[822]), .Z(n[1845]) );
  AN2D0 U5212 ( .A1(b[8]), .A2(n[819]), .Z(n[1842]) );
  AN2D0 U5213 ( .A1(b[8]), .A2(n[816]), .Z(n[1839]) );
  AN2D0 U5214 ( .A1(b[8]), .A2(n[815]), .Z(n[1838]) );
  AN2D0 U5215 ( .A1(b[8]), .A2(n[812]), .Z(n[1835]) );
  AN2D0 U5216 ( .A1(b[8]), .A2(n[809]), .Z(n[1832]) );
  AN2D0 U5217 ( .A1(b[8]), .A2(n[808]), .Z(n[1831]) );
  AN2D0 U5218 ( .A1(b[8]), .A2(n[807]), .Z(n[1830]) );
  AN2D0 U5219 ( .A1(b[8]), .A2(n[804]), .Z(n[1827]) );
  AN2D0 U5220 ( .A1(b[8]), .A2(n[801]), .Z(n[1824]) );
  AN2D0 U5221 ( .A1(b[8]), .A2(n[800]), .Z(n[1823]) );
  AN2D0 U5222 ( .A1(b[8]), .A2(n[797]), .Z(n[1820]) );
  AN2D0 U5223 ( .A1(b[8]), .A2(n[794]), .Z(n[1817]) );
  AN2D0 U5224 ( .A1(b[8]), .A2(n[793]), .Z(n[1816]) );
  AN2D0 U5225 ( .A1(b[8]), .A2(n[792]), .Z(n[1815]) );
  AN2D0 U5226 ( .A1(b[8]), .A2(n[791]), .Z(n[1814]) );
  AN2D0 U5227 ( .A1(b[8]), .A2(n[788]), .Z(n[1811]) );
  AN2D0 U5228 ( .A1(b[8]), .A2(n[785]), .Z(n[1808]) );
  AN2D0 U5229 ( .A1(b[8]), .A2(n[784]), .Z(n[1807]) );
  AN2D0 U5230 ( .A1(b[8]), .A2(n[781]), .Z(n[1804]) );
  AN2D0 U5231 ( .A1(b[8]), .A2(n[778]), .Z(n[1801]) );
  AN2D0 U5232 ( .A1(b[8]), .A2(n[777]), .Z(n[1800]) );
  AN2D0 U5233 ( .A1(b[8]), .A2(n[776]), .Z(n[1799]) );
  AN2D0 U5234 ( .A1(b[8]), .A2(n[773]), .Z(n[1796]) );
  AN2D0 U5235 ( .A1(b[8]), .A2(n[770]), .Z(n[1793]) );
  AN2D0 U5236 ( .A1(b[8]), .A2(n[769]), .Z(n[1792]) );
  AN2D0 U5237 ( .A1(b[8]), .A2(n[766]), .Z(n[1789]) );
  AN2D0 U5238 ( .A1(b[8]), .A2(n[763]), .Z(n[1786]) );
  AN2D0 U5239 ( .A1(b[8]), .A2(n[762]), .Z(n[1785]) );
  AN2D0 U5240 ( .A1(b[8]), .A2(n[761]), .Z(n[1784]) );
  AN2D0 U5241 ( .A1(b[8]), .A2(n[760]), .Z(n[1783]) );
  AN2D0 U5242 ( .A1(b[8]), .A2(n[759]), .Z(n[1782]) );
  AN2D0 U5243 ( .A1(b[8]), .A2(n[758]), .Z(n[1781]) );
  AN2D0 U5244 ( .A1(b[8]), .A2(n[757]), .Z(n[1780]) );
  AN2D0 U5245 ( .A1(b[8]), .A2(n[754]), .Z(n[1777]) );
  AN2D0 U5246 ( .A1(b[8]), .A2(n[751]), .Z(n[1774]) );
  AN2D0 U5247 ( .A1(b[8]), .A2(n[750]), .Z(n[1773]) );
  AN2D0 U5248 ( .A1(b[8]), .A2(n[747]), .Z(n[1770]) );
  AN2D0 U5249 ( .A1(b[8]), .A2(n[744]), .Z(n[1767]) );
  AN2D0 U5250 ( .A1(b[8]), .A2(n[743]), .Z(n[1766]) );
  AN2D0 U5251 ( .A1(b[8]), .A2(n[742]), .Z(n[1765]) );
  AN2D0 U5252 ( .A1(b[8]), .A2(n[739]), .Z(n[1762]) );
  AN2D0 U5253 ( .A1(b[8]), .A2(n[736]), .Z(n[1759]) );
  AN2D0 U5254 ( .A1(b[8]), .A2(n[735]), .Z(n[1758]) );
  AN2D0 U5255 ( .A1(b[8]), .A2(n[732]), .Z(n[1755]) );
  AN2D0 U5256 ( .A1(b[8]), .A2(n[729]), .Z(n[1752]) );
  AN2D0 U5257 ( .A1(b[8]), .A2(n[728]), .Z(n[1751]) );
  AN2D0 U5258 ( .A1(b[8]), .A2(n[727]), .Z(n[1750]) );
  AN2D0 U5259 ( .A1(b[8]), .A2(n[726]), .Z(n[1749]) );
  AN2D0 U5260 ( .A1(b[8]), .A2(n[723]), .Z(n[1746]) );
  AN2D0 U5261 ( .A1(b[8]), .A2(n[720]), .Z(n[1743]) );
  AN2D0 U5262 ( .A1(b[8]), .A2(n[719]), .Z(n[1742]) );
  AN2D0 U5263 ( .A1(b[8]), .A2(n[716]), .Z(n[1739]) );
  AN2D0 U5264 ( .A1(b[8]), .A2(n[713]), .Z(n[1736]) );
  AN2D0 U5265 ( .A1(b[8]), .A2(n[712]), .Z(n[1735]) );
  AN2D0 U5266 ( .A1(b[8]), .A2(n[711]), .Z(n[1734]) );
  AN2D0 U5267 ( .A1(b[8]), .A2(n[708]), .Z(n[1731]) );
  AN2D0 U5268 ( .A1(b[8]), .A2(n[705]), .Z(n[1728]) );
  AN2D0 U5269 ( .A1(b[8]), .A2(n[704]), .Z(n[1727]) );
  AN2D0 U5270 ( .A1(b[8]), .A2(n[701]), .Z(n[1724]) );
  AN2D0 U5271 ( .A1(b[8]), .A2(n[698]), .Z(n[1721]) );
  AN2D0 U5272 ( .A1(b[8]), .A2(n[697]), .Z(n[1720]) );
  AN2D0 U5273 ( .A1(b[8]), .A2(n[696]), .Z(n[1719]) );
  AN2D0 U5274 ( .A1(b[8]), .A2(n[695]), .Z(n[1718]) );
  AN2D0 U5275 ( .A1(b[8]), .A2(n[694]), .Z(n[1717]) );
  AN2D0 U5276 ( .A1(b[8]), .A2(n[691]), .Z(n[1714]) );
  AN2D0 U5277 ( .A1(b[8]), .A2(n[688]), .Z(n[1711]) );
  AN2D0 U5278 ( .A1(b[8]), .A2(n[687]), .Z(n[1710]) );
  AN2D0 U5279 ( .A1(b[8]), .A2(n[684]), .Z(n[1707]) );
  AN2D0 U5280 ( .A1(b[8]), .A2(n[681]), .Z(n[1704]) );
  AN2D0 U5281 ( .A1(b[8]), .A2(n[680]), .Z(n[1703]) );
  AN2D0 U5282 ( .A1(b[8]), .A2(n[679]), .Z(n[1702]) );
  AN2D0 U5283 ( .A1(b[8]), .A2(n[676]), .Z(n[1699]) );
  AN2D0 U5284 ( .A1(b[8]), .A2(n[673]), .Z(n[1696]) );
  AN2D0 U5285 ( .A1(b[8]), .A2(n[672]), .Z(n[1695]) );
  AN2D0 U5286 ( .A1(b[8]), .A2(n[669]), .Z(n[1692]) );
  AN2D0 U5287 ( .A1(b[8]), .A2(n[666]), .Z(n[1689]) );
  AN2D0 U5288 ( .A1(b[8]), .A2(n[665]), .Z(n[1688]) );
  AN2D0 U5289 ( .A1(b[8]), .A2(n[664]), .Z(n[1687]) );
  AN2D0 U5290 ( .A1(b[8]), .A2(n[663]), .Z(n[1686]) );
  AN2D0 U5291 ( .A1(b[8]), .A2(n[660]), .Z(n[1683]) );
  AN2D0 U5292 ( .A1(b[8]), .A2(n[657]), .Z(n[1680]) );
  AN2D0 U5293 ( .A1(b[8]), .A2(n[656]), .Z(n[1679]) );
  AN2D0 U5294 ( .A1(b[8]), .A2(n[653]), .Z(n[1676]) );
  AN2D0 U5295 ( .A1(b[8]), .A2(n[650]), .Z(n[1673]) );
  AN2D0 U5296 ( .A1(b[8]), .A2(n[649]), .Z(n[1672]) );
  AN2D0 U5297 ( .A1(b[8]), .A2(n[648]), .Z(n[1671]) );
  AN2D0 U5298 ( .A1(b[8]), .A2(n[645]), .Z(n[1668]) );
  AN2D0 U5299 ( .A1(b[8]), .A2(n[642]), .Z(n[1665]) );
  AN2D0 U5300 ( .A1(b[8]), .A2(n[641]), .Z(n[1664]) );
  AN2D0 U5301 ( .A1(b[8]), .A2(n[638]), .Z(n[1661]) );
  AN2D0 U5302 ( .A1(b[8]), .A2(n[635]), .Z(n[1658]) );
  AN2D0 U5303 ( .A1(b[8]), .A2(n[634]), .Z(n[1657]) );
  AN2D0 U5304 ( .A1(b[8]), .A2(n[633]), .Z(n[1656]) );
  AN2D0 U5305 ( .A1(b[8]), .A2(n[632]), .Z(n[1655]) );
  AN2D0 U5306 ( .A1(b[8]), .A2(n[631]), .Z(n[1654]) );
  AN2D0 U5307 ( .A1(b[8]), .A2(n[630]), .Z(n[1653]) );
  AN2D0 U5308 ( .A1(b[8]), .A2(n[627]), .Z(n[1650]) );
  AN2D0 U5309 ( .A1(b[8]), .A2(n[624]), .Z(n[1647]) );
  AN2D0 U5310 ( .A1(b[8]), .A2(n[623]), .Z(n[1646]) );
  AN2D0 U5311 ( .A1(b[8]), .A2(n[620]), .Z(n[1643]) );
  AN2D0 U5312 ( .A1(b[8]), .A2(n[617]), .Z(n[1640]) );
  AN2D0 U5313 ( .A1(b[8]), .A2(n[616]), .Z(n[1639]) );
  AN2D0 U5314 ( .A1(b[8]), .A2(n[615]), .Z(n[1638]) );
  AN2D0 U5315 ( .A1(b[8]), .A2(n[612]), .Z(n[1635]) );
  AN2D0 U5316 ( .A1(b[8]), .A2(n[609]), .Z(n[1632]) );
  AN2D0 U5317 ( .A1(b[8]), .A2(n[608]), .Z(n[1631]) );
  AN2D0 U5318 ( .A1(b[8]), .A2(n[605]), .Z(n[1628]) );
  AN2D0 U5319 ( .A1(b[8]), .A2(n[602]), .Z(n[1625]) );
  AN2D0 U5320 ( .A1(b[8]), .A2(n[601]), .Z(n[1624]) );
  AN2D0 U5321 ( .A1(b[8]), .A2(n[600]), .Z(n[1623]) );
  AN2D0 U5322 ( .A1(b[8]), .A2(n[599]), .Z(n[1622]) );
  AN2D0 U5323 ( .A1(b[8]), .A2(n[596]), .Z(n[1619]) );
  AN2D0 U5324 ( .A1(b[8]), .A2(n[593]), .Z(n[1616]) );
  AN2D0 U5325 ( .A1(b[8]), .A2(n[592]), .Z(n[1615]) );
  AN2D0 U5326 ( .A1(b[8]), .A2(n[589]), .Z(n[1612]) );
  AN2D0 U5327 ( .A1(b[8]), .A2(n[586]), .Z(n[1609]) );
  AN2D0 U5328 ( .A1(b[8]), .A2(n[585]), .Z(n[1608]) );
  AN2D0 U5329 ( .A1(b[8]), .A2(n[584]), .Z(n[1607]) );
  AN2D0 U5330 ( .A1(b[8]), .A2(n[581]), .Z(n[1604]) );
  AN2D0 U5331 ( .A1(b[8]), .A2(n[578]), .Z(n[1601]) );
  AN2D0 U5332 ( .A1(b[8]), .A2(n[577]), .Z(n[1600]) );
  AN2D0 U5333 ( .A1(b[8]), .A2(n[574]), .Z(n[1597]) );
  AN2D0 U5334 ( .A1(b[8]), .A2(n[571]), .Z(n[1594]) );
  AN2D0 U5335 ( .A1(b[8]), .A2(n[570]), .Z(n[1593]) );
  AN2D0 U5336 ( .A1(b[8]), .A2(n[569]), .Z(n[1592]) );
  AN2D0 U5337 ( .A1(b[8]), .A2(n[568]), .Z(n[1591]) );
  AN2D0 U5338 ( .A1(b[8]), .A2(n[567]), .Z(n[1590]) );
  AN2D0 U5339 ( .A1(b[8]), .A2(n[564]), .Z(n[1587]) );
  AN2D0 U5340 ( .A1(b[8]), .A2(n[561]), .Z(n[1584]) );
  AN2D0 U5341 ( .A1(b[8]), .A2(n[560]), .Z(n[1583]) );
  AN2D0 U5342 ( .A1(b[8]), .A2(n[557]), .Z(n[1580]) );
  AN2D0 U5343 ( .A1(b[8]), .A2(n[554]), .Z(n[1577]) );
  AN2D0 U5344 ( .A1(b[8]), .A2(n[553]), .Z(n[1576]) );
  AN2D0 U5345 ( .A1(b[8]), .A2(n[552]), .Z(n[1575]) );
  AN2D0 U5346 ( .A1(b[8]), .A2(n[549]), .Z(n[1572]) );
  AN2D0 U5347 ( .A1(b[8]), .A2(n[546]), .Z(n[1569]) );
  AN2D0 U5348 ( .A1(b[8]), .A2(n[545]), .Z(n[1568]) );
  AN2D0 U5349 ( .A1(b[8]), .A2(n[542]), .Z(n[1565]) );
  AN2D0 U5350 ( .A1(b[8]), .A2(n[539]), .Z(n[1562]) );
  AN2D0 U5351 ( .A1(b[8]), .A2(n[538]), .Z(n[1561]) );
  AN2D0 U5352 ( .A1(b[8]), .A2(n[537]), .Z(n[1560]) );
  AN2D0 U5353 ( .A1(b[8]), .A2(n[536]), .Z(n[1559]) );
  AN2D0 U5354 ( .A1(b[8]), .A2(n[533]), .Z(n[1556]) );
  AN2D0 U5355 ( .A1(b[8]), .A2(n[530]), .Z(n[1553]) );
  AN2D0 U5356 ( .A1(b[8]), .A2(n[529]), .Z(n[1552]) );
  AN2D0 U5357 ( .A1(b[8]), .A2(n[526]), .Z(n[1549]) );
  AN2D0 U5358 ( .A1(b[8]), .A2(n[523]), .Z(n[1546]) );
  AN2D0 U5359 ( .A1(b[8]), .A2(n[522]), .Z(n[1545]) );
  AN2D0 U5360 ( .A1(b[8]), .A2(n[521]), .Z(n[1544]) );
  AN2D0 U5361 ( .A1(b[8]), .A2(n[518]), .Z(n[1541]) );
  AN2D0 U5362 ( .A1(b[8]), .A2(n[515]), .Z(n[1538]) );
  AN2D0 U5363 ( .A1(b[8]), .A2(n[514]), .Z(n[1537]) );
  AN2D0 U5364 ( .A1(b[8]), .A2(n[511]), .Z(n[1534]) );
  AN2D0 U5365 ( .A1(b[8]), .A2(n[508]), .Z(n[1531]) );
  AN2D0 U5366 ( .A1(b[8]), .A2(n[507]), .Z(n[1530]) );
  AN2D0 U5367 ( .A1(b[8]), .A2(n[506]), .Z(n[1529]) );
  AN2D0 U5368 ( .A1(b[8]), .A2(n[505]), .Z(n[1528]) );
  AN2D0 U5369 ( .A1(b[8]), .A2(n[504]), .Z(n[1527]) );
  AN2D0 U5370 ( .A1(b[8]), .A2(n[503]), .Z(n[1526]) );
  AN2D0 U5371 ( .A1(b[8]), .A2(n[502]), .Z(n[1525]) );
  AN2D0 U5372 ( .A1(b[8]), .A2(n[501]), .Z(n[1524]) );
  AN2D0 U5373 ( .A1(n[1009]), .A2(a[8]), .Z(n[1521]) );
  AN2D0 U5374 ( .A1(n[1006]), .A2(a[8]), .Z(n[1518]) );
  AN2D0 U5375 ( .A1(n[1005]), .A2(a[8]), .Z(n[1517]) );
  AN2D0 U5376 ( .A1(n[1002]), .A2(a[8]), .Z(n[1514]) );
  AN2D0 U5377 ( .A1(n[999]), .A2(a[8]), .Z(n[1511]) );
  AN2D0 U5378 ( .A1(n[488]), .A2(b[7]), .Z(n[999]) );
  AN2D0 U5379 ( .A1(n[998]), .A2(a[8]), .Z(n[1510]) );
  AN2D0 U5380 ( .A1(b[7]), .A2(n[487]), .Z(n[998]) );
  AN2D0 U5381 ( .A1(n[997]), .A2(a[8]), .Z(n[1509]) );
  AN2D0 U5382 ( .A1(b[7]), .A2(n[486]), .Z(n[997]) );
  AN2D0 U5383 ( .A1(n[994]), .A2(a[8]), .Z(n[1506]) );
  AN2D0 U5384 ( .A1(b[7]), .A2(n[483]), .Z(n[994]) );
  AN2D0 U5385 ( .A1(n[991]), .A2(a[8]), .Z(n[1503]) );
  AN2D0 U5386 ( .A1(b[7]), .A2(n[480]), .Z(n[991]) );
  AN2D0 U5387 ( .A1(n[990]), .A2(a[8]), .Z(n[1502]) );
  AN2D0 U5388 ( .A1(b[7]), .A2(n[479]), .Z(n[990]) );
  AN2D0 U5389 ( .A1(n[987]), .A2(a[8]), .Z(n[1499]) );
  AN2D0 U5390 ( .A1(b[7]), .A2(n[476]), .Z(n[987]) );
  AN2D0 U5391 ( .A1(n[984]), .A2(a[8]), .Z(n[1496]) );
  AN2D0 U5392 ( .A1(b[7]), .A2(n[473]), .Z(n[984]) );
  AN2D0 U5393 ( .A1(n[983]), .A2(a[8]), .Z(n[1495]) );
  AN2D0 U5394 ( .A1(b[7]), .A2(n[472]), .Z(n[983]) );
  AN2D0 U5395 ( .A1(n[982]), .A2(a[8]), .Z(n[1494]) );
  AN2D0 U5396 ( .A1(b[7]), .A2(n[471]), .Z(n[982]) );
  AN2D0 U5397 ( .A1(n[981]), .A2(a[8]), .Z(n[1493]) );
  AN2D0 U5398 ( .A1(b[7]), .A2(n[470]), .Z(n[981]) );
  AN2D0 U5399 ( .A1(n[978]), .A2(a[8]), .Z(n[1490]) );
  AN2D0 U5400 ( .A1(b[7]), .A2(n[467]), .Z(n[978]) );
  AN2D0 U5401 ( .A1(n[975]), .A2(a[8]), .Z(n[1487]) );
  AN2D0 U5402 ( .A1(b[7]), .A2(n[464]), .Z(n[975]) );
  AN2D0 U5403 ( .A1(n[974]), .A2(a[8]), .Z(n[1486]) );
  AN2D0 U5404 ( .A1(b[7]), .A2(n[463]), .Z(n[974]) );
  AN2D0 U5405 ( .A1(n[971]), .A2(a[8]), .Z(n[1483]) );
  AN2D0 U5406 ( .A1(b[7]), .A2(n[460]), .Z(n[971]) );
  AN2D0 U5407 ( .A1(n[968]), .A2(a[8]), .Z(n[1480]) );
  AN2D0 U5408 ( .A1(b[7]), .A2(n[457]), .Z(n[968]) );
  AN2D0 U5409 ( .A1(n[967]), .A2(a[8]), .Z(n[1479]) );
  AN2D0 U5410 ( .A1(b[7]), .A2(n[456]), .Z(n[967]) );
  AN2D0 U5411 ( .A1(n[966]), .A2(a[8]), .Z(n[1478]) );
  AN2D0 U5412 ( .A1(b[7]), .A2(n[455]), .Z(n[966]) );
  AN2D0 U5413 ( .A1(n[963]), .A2(a[8]), .Z(n[1475]) );
  AN2D0 U5414 ( .A1(b[7]), .A2(n[452]), .Z(n[963]) );
  AN2D0 U5415 ( .A1(n[960]), .A2(a[8]), .Z(n[1472]) );
  AN2D0 U5416 ( .A1(b[7]), .A2(n[449]), .Z(n[960]) );
  AN2D0 U5417 ( .A1(n[959]), .A2(a[8]), .Z(n[1471]) );
  AN2D0 U5418 ( .A1(b[7]), .A2(n[448]), .Z(n[959]) );
  AN2D0 U5419 ( .A1(n[956]), .A2(a[8]), .Z(n[1468]) );
  AN2D0 U5420 ( .A1(b[7]), .A2(n[445]), .Z(n[956]) );
  AN2D0 U5421 ( .A1(n[953]), .A2(a[8]), .Z(n[1465]) );
  AN2D0 U5422 ( .A1(b[7]), .A2(n[442]), .Z(n[953]) );
  AN2D0 U5423 ( .A1(n[952]), .A2(a[8]), .Z(n[1464]) );
  AN2D0 U5424 ( .A1(b[7]), .A2(n[441]), .Z(n[952]) );
  AN2D0 U5425 ( .A1(n[951]), .A2(a[8]), .Z(n[1463]) );
  AN2D0 U5426 ( .A1(b[7]), .A2(n[440]), .Z(n[951]) );
  AN2D0 U5427 ( .A1(n[950]), .A2(a[8]), .Z(n[1462]) );
  AN2D0 U5428 ( .A1(b[7]), .A2(n[439]), .Z(n[950]) );
  AN2D0 U5429 ( .A1(n[949]), .A2(a[8]), .Z(n[1461]) );
  AN2D0 U5430 ( .A1(b[7]), .A2(n[438]), .Z(n[949]) );
  AN2D0 U5431 ( .A1(n[946]), .A2(a[8]), .Z(n[1458]) );
  AN2D0 U5432 ( .A1(b[7]), .A2(n[435]), .Z(n[946]) );
  AN2D0 U5433 ( .A1(n[943]), .A2(a[8]), .Z(n[1455]) );
  AN2D0 U5434 ( .A1(b[7]), .A2(n[432]), .Z(n[943]) );
  AN2D0 U5435 ( .A1(n[942]), .A2(a[8]), .Z(n[1454]) );
  AN2D0 U5436 ( .A1(b[7]), .A2(n[431]), .Z(n[942]) );
  AN2D0 U5437 ( .A1(n[939]), .A2(a[8]), .Z(n[1451]) );
  AN2D0 U5438 ( .A1(b[7]), .A2(n[428]), .Z(n[939]) );
  AN2D0 U5439 ( .A1(n[936]), .A2(a[8]), .Z(n[1448]) );
  AN2D0 U5440 ( .A1(b[7]), .A2(n[425]), .Z(n[936]) );
  AN2D0 U5441 ( .A1(n[935]), .A2(a[8]), .Z(n[1447]) );
  AN2D0 U5442 ( .A1(b[7]), .A2(n[424]), .Z(n[935]) );
  AN2D0 U5443 ( .A1(n[934]), .A2(a[8]), .Z(n[1446]) );
  AN2D0 U5444 ( .A1(b[7]), .A2(n[423]), .Z(n[934]) );
  AN2D0 U5445 ( .A1(n[931]), .A2(a[8]), .Z(n[1443]) );
  AN2D0 U5446 ( .A1(b[7]), .A2(n[420]), .Z(n[931]) );
  AN2D0 U5447 ( .A1(n[928]), .A2(a[8]), .Z(n[1440]) );
  AN2D0 U5448 ( .A1(b[7]), .A2(n[417]), .Z(n[928]) );
  AN2D0 U5449 ( .A1(n[927]), .A2(a[8]), .Z(n[1439]) );
  AN2D0 U5450 ( .A1(b[7]), .A2(n[416]), .Z(n[927]) );
  AN2D0 U5451 ( .A1(n[924]), .A2(a[8]), .Z(n[1436]) );
  AN2D0 U5452 ( .A1(b[7]), .A2(n[413]), .Z(n[924]) );
  AN2D0 U5453 ( .A1(n[921]), .A2(a[8]), .Z(n[1433]) );
  AN2D0 U5454 ( .A1(b[7]), .A2(n[410]), .Z(n[921]) );
  AN2D0 U5455 ( .A1(n[920]), .A2(a[8]), .Z(n[1432]) );
  AN2D0 U5456 ( .A1(b[7]), .A2(n[409]), .Z(n[920]) );
  AN2D0 U5457 ( .A1(n[919]), .A2(a[8]), .Z(n[1431]) );
  AN2D0 U5458 ( .A1(b[7]), .A2(n[408]), .Z(n[919]) );
  AN2D0 U5459 ( .A1(n[918]), .A2(a[8]), .Z(n[1430]) );
  AN2D0 U5460 ( .A1(b[7]), .A2(n[407]), .Z(n[918]) );
  AN2D0 U5461 ( .A1(n[915]), .A2(a[8]), .Z(n[1427]) );
  AN2D0 U5462 ( .A1(b[7]), .A2(n[404]), .Z(n[915]) );
  AN2D0 U5463 ( .A1(n[912]), .A2(a[8]), .Z(n[1424]) );
  AN2D0 U5464 ( .A1(b[7]), .A2(n[401]), .Z(n[912]) );
  AN2D0 U5465 ( .A1(n[911]), .A2(a[8]), .Z(n[1423]) );
  AN2D0 U5466 ( .A1(b[7]), .A2(n[400]), .Z(n[911]) );
  AN2D0 U5467 ( .A1(n[908]), .A2(a[8]), .Z(n[1420]) );
  AN2D0 U5468 ( .A1(b[7]), .A2(n[397]), .Z(n[908]) );
  AN2D0 U5469 ( .A1(n[905]), .A2(a[8]), .Z(n[1417]) );
  AN2D0 U5470 ( .A1(b[7]), .A2(n[394]), .Z(n[905]) );
  AN2D0 U5471 ( .A1(n[904]), .A2(a[8]), .Z(n[1416]) );
  AN2D0 U5472 ( .A1(b[7]), .A2(n[393]), .Z(n[904]) );
  AN2D0 U5473 ( .A1(n[903]), .A2(a[8]), .Z(n[1415]) );
  AN2D0 U5474 ( .A1(b[7]), .A2(n[392]), .Z(n[903]) );
  AN2D0 U5475 ( .A1(n[900]), .A2(a[8]), .Z(n[1412]) );
  AN2D0 U5476 ( .A1(b[7]), .A2(n[389]), .Z(n[900]) );
  AN2D0 U5477 ( .A1(n[897]), .A2(a[8]), .Z(n[1409]) );
  AN2D0 U5478 ( .A1(b[7]), .A2(n[386]), .Z(n[897]) );
  AN2D0 U5479 ( .A1(n[896]), .A2(a[8]), .Z(n[1408]) );
  AN2D0 U5480 ( .A1(b[7]), .A2(n[385]), .Z(n[896]) );
  AN2D0 U5481 ( .A1(n[893]), .A2(a[8]), .Z(n[1405]) );
  AN2D0 U5482 ( .A1(b[7]), .A2(n[382]), .Z(n[893]) );
  AN2D0 U5483 ( .A1(n[890]), .A2(a[8]), .Z(n[1402]) );
  AN2D0 U5484 ( .A1(b[7]), .A2(n[379]), .Z(n[890]) );
  AN2D0 U5485 ( .A1(n[889]), .A2(a[8]), .Z(n[1401]) );
  AN2D0 U5486 ( .A1(b[7]), .A2(n[378]), .Z(n[889]) );
  AN2D0 U5487 ( .A1(n[888]), .A2(a[8]), .Z(n[1400]) );
  AN2D0 U5488 ( .A1(b[7]), .A2(n[377]), .Z(n[888]) );
  AN2D0 U5489 ( .A1(n[887]), .A2(a[8]), .Z(n[1399]) );
  AN2D0 U5490 ( .A1(b[7]), .A2(n[376]), .Z(n[887]) );
  AN2D0 U5491 ( .A1(n[886]), .A2(a[8]), .Z(n[1398]) );
  AN2D0 U5492 ( .A1(b[7]), .A2(n[375]), .Z(n[886]) );
  AN2D0 U5493 ( .A1(n[885]), .A2(a[8]), .Z(n[1397]) );
  AN2D0 U5494 ( .A1(b[7]), .A2(n[374]), .Z(n[885]) );
  AN2D0 U5495 ( .A1(n[882]), .A2(a[8]), .Z(n[1394]) );
  AN2D0 U5496 ( .A1(b[7]), .A2(n[371]), .Z(n[882]) );
  AN2D0 U5497 ( .A1(n[879]), .A2(a[8]), .Z(n[1391]) );
  AN2D0 U5498 ( .A1(b[7]), .A2(n[368]), .Z(n[879]) );
  AN2D0 U5499 ( .A1(n[878]), .A2(a[8]), .Z(n[1390]) );
  AN2D0 U5500 ( .A1(b[7]), .A2(n[367]), .Z(n[878]) );
  AN2D0 U5501 ( .A1(n[875]), .A2(a[8]), .Z(n[1387]) );
  AN2D0 U5502 ( .A1(b[7]), .A2(n[364]), .Z(n[875]) );
  AN2D0 U5503 ( .A1(n[872]), .A2(a[8]), .Z(n[1384]) );
  AN2D0 U5504 ( .A1(b[7]), .A2(n[361]), .Z(n[872]) );
  AN2D0 U5505 ( .A1(n[871]), .A2(a[8]), .Z(n[1383]) );
  AN2D0 U5506 ( .A1(b[7]), .A2(n[360]), .Z(n[871]) );
  AN2D0 U5507 ( .A1(n[870]), .A2(a[8]), .Z(n[1382]) );
  AN2D0 U5508 ( .A1(b[7]), .A2(n[359]), .Z(n[870]) );
  AN2D0 U5509 ( .A1(n[867]), .A2(a[8]), .Z(n[1379]) );
  AN2D0 U5510 ( .A1(b[7]), .A2(n[356]), .Z(n[867]) );
  AN2D0 U5511 ( .A1(n[864]), .A2(a[8]), .Z(n[1376]) );
  AN2D0 U5512 ( .A1(b[7]), .A2(n[353]), .Z(n[864]) );
  AN2D0 U5513 ( .A1(n[863]), .A2(a[8]), .Z(n[1375]) );
  AN2D0 U5514 ( .A1(b[7]), .A2(n[352]), .Z(n[863]) );
  AN2D0 U5515 ( .A1(n[860]), .A2(a[8]), .Z(n[1372]) );
  AN2D0 U5516 ( .A1(b[7]), .A2(n[349]), .Z(n[860]) );
  AN2D0 U5517 ( .A1(n[857]), .A2(a[8]), .Z(n[1369]) );
  AN2D0 U5518 ( .A1(b[7]), .A2(n[346]), .Z(n[857]) );
  AN2D0 U5519 ( .A1(n[856]), .A2(a[8]), .Z(n[1368]) );
  AN2D0 U5520 ( .A1(b[7]), .A2(n[345]), .Z(n[856]) );
  AN2D0 U5521 ( .A1(n[855]), .A2(a[8]), .Z(n[1367]) );
  AN2D0 U5522 ( .A1(b[7]), .A2(n[344]), .Z(n[855]) );
  AN2D0 U5523 ( .A1(n[854]), .A2(a[8]), .Z(n[1366]) );
  AN2D0 U5524 ( .A1(b[7]), .A2(n[343]), .Z(n[854]) );
  AN2D0 U5525 ( .A1(n[851]), .A2(a[8]), .Z(n[1363]) );
  AN2D0 U5526 ( .A1(b[7]), .A2(n[340]), .Z(n[851]) );
  AN2D0 U5527 ( .A1(n[848]), .A2(a[8]), .Z(n[1360]) );
  AN2D0 U5528 ( .A1(b[7]), .A2(n[337]), .Z(n[848]) );
  AN2D0 U5529 ( .A1(n[847]), .A2(a[8]), .Z(n[1359]) );
  AN2D0 U5530 ( .A1(b[7]), .A2(n[336]), .Z(n[847]) );
  AN2D0 U5531 ( .A1(n[844]), .A2(a[8]), .Z(n[1356]) );
  AN2D0 U5532 ( .A1(b[7]), .A2(n[333]), .Z(n[844]) );
  AN2D0 U5533 ( .A1(n[841]), .A2(a[8]), .Z(n[1353]) );
  AN2D0 U5534 ( .A1(b[7]), .A2(n[330]), .Z(n[841]) );
  AN2D0 U5535 ( .A1(n[840]), .A2(a[8]), .Z(n[1352]) );
  AN2D0 U5536 ( .A1(b[7]), .A2(n[329]), .Z(n[840]) );
  AN2D0 U5537 ( .A1(n[839]), .A2(a[8]), .Z(n[1351]) );
  AN2D0 U5538 ( .A1(b[7]), .A2(n[328]), .Z(n[839]) );
  AN2D0 U5539 ( .A1(n[836]), .A2(a[8]), .Z(n[1348]) );
  AN2D0 U5540 ( .A1(b[7]), .A2(n[325]), .Z(n[836]) );
  AN2D0 U5541 ( .A1(n[833]), .A2(a[8]), .Z(n[1345]) );
  AN2D0 U5542 ( .A1(b[7]), .A2(n[322]), .Z(n[833]) );
  AN2D0 U5543 ( .A1(n[832]), .A2(a[8]), .Z(n[1344]) );
  AN2D0 U5544 ( .A1(b[7]), .A2(n[321]), .Z(n[832]) );
  AN2D0 U5545 ( .A1(n[829]), .A2(a[8]), .Z(n[1341]) );
  AN2D0 U5546 ( .A1(b[7]), .A2(n[318]), .Z(n[829]) );
  AN2D0 U5547 ( .A1(n[826]), .A2(a[8]), .Z(n[1338]) );
  AN2D0 U5548 ( .A1(b[7]), .A2(n[315]), .Z(n[826]) );
  AN2D0 U5549 ( .A1(n[825]), .A2(a[8]), .Z(n[1337]) );
  AN2D0 U5550 ( .A1(b[7]), .A2(n[314]), .Z(n[825]) );
  AN2D0 U5551 ( .A1(n[824]), .A2(a[8]), .Z(n[1336]) );
  AN2D0 U5552 ( .A1(b[7]), .A2(n[313]), .Z(n[824]) );
  AN2D0 U5553 ( .A1(n[823]), .A2(a[8]), .Z(n[1335]) );
  AN2D0 U5554 ( .A1(b[7]), .A2(n[312]), .Z(n[823]) );
  AN2D0 U5555 ( .A1(n[822]), .A2(a[8]), .Z(n[1334]) );
  AN2D0 U5556 ( .A1(b[7]), .A2(n[311]), .Z(n[822]) );
  AN2D0 U5557 ( .A1(n[819]), .A2(a[8]), .Z(n[1331]) );
  AN2D0 U5558 ( .A1(b[7]), .A2(n[308]), .Z(n[819]) );
  AN2D0 U5559 ( .A1(n[816]), .A2(a[8]), .Z(n[1328]) );
  AN2D0 U5560 ( .A1(b[7]), .A2(n[305]), .Z(n[816]) );
  AN2D0 U5561 ( .A1(n[815]), .A2(a[8]), .Z(n[1327]) );
  AN2D0 U5562 ( .A1(b[7]), .A2(n[304]), .Z(n[815]) );
  AN2D0 U5563 ( .A1(n[812]), .A2(a[8]), .Z(n[1324]) );
  AN2D0 U5564 ( .A1(b[7]), .A2(n[301]), .Z(n[812]) );
  AN2D0 U5565 ( .A1(n[809]), .A2(a[8]), .Z(n[1321]) );
  AN2D0 U5566 ( .A1(b[7]), .A2(n[298]), .Z(n[809]) );
  AN2D0 U5567 ( .A1(n[808]), .A2(a[8]), .Z(n[1320]) );
  AN2D0 U5568 ( .A1(b[7]), .A2(n[297]), .Z(n[808]) );
  AN2D0 U5569 ( .A1(n[807]), .A2(a[8]), .Z(n[1319]) );
  AN2D0 U5570 ( .A1(b[7]), .A2(n[296]), .Z(n[807]) );
  AN2D0 U5571 ( .A1(n[804]), .A2(a[8]), .Z(n[1316]) );
  AN2D0 U5572 ( .A1(b[7]), .A2(n[293]), .Z(n[804]) );
  AN2D0 U5573 ( .A1(n[801]), .A2(a[8]), .Z(n[1313]) );
  AN2D0 U5574 ( .A1(b[7]), .A2(n[290]), .Z(n[801]) );
  AN2D0 U5575 ( .A1(n[800]), .A2(a[8]), .Z(n[1312]) );
  AN2D0 U5576 ( .A1(b[7]), .A2(n[289]), .Z(n[800]) );
  AN2D0 U5577 ( .A1(n[797]), .A2(a[8]), .Z(n[1309]) );
  AN2D0 U5578 ( .A1(b[7]), .A2(n[286]), .Z(n[797]) );
  AN2D0 U5579 ( .A1(n[794]), .A2(a[8]), .Z(n[1306]) );
  AN2D0 U5580 ( .A1(b[7]), .A2(n[283]), .Z(n[794]) );
  AN2D0 U5581 ( .A1(n[793]), .A2(a[8]), .Z(n[1305]) );
  AN2D0 U5582 ( .A1(b[7]), .A2(n[282]), .Z(n[793]) );
  AN2D0 U5583 ( .A1(n[792]), .A2(a[8]), .Z(n[1304]) );
  AN2D0 U5584 ( .A1(b[7]), .A2(n[281]), .Z(n[792]) );
  AN2D0 U5585 ( .A1(n[791]), .A2(a[8]), .Z(n[1303]) );
  AN2D0 U5586 ( .A1(b[7]), .A2(n[280]), .Z(n[791]) );
  AN2D0 U5587 ( .A1(n[788]), .A2(a[8]), .Z(n[1300]) );
  AN2D0 U5588 ( .A1(b[7]), .A2(n[277]), .Z(n[788]) );
  AN2D0 U5589 ( .A1(n[785]), .A2(a[8]), .Z(n[1297]) );
  AN2D0 U5590 ( .A1(b[7]), .A2(n[274]), .Z(n[785]) );
  AN2D0 U5591 ( .A1(n[784]), .A2(a[8]), .Z(n[1296]) );
  AN2D0 U5592 ( .A1(b[7]), .A2(n[273]), .Z(n[784]) );
  AN2D0 U5593 ( .A1(n[781]), .A2(a[8]), .Z(n[1293]) );
  AN2D0 U5594 ( .A1(b[7]), .A2(n[270]), .Z(n[781]) );
  AN2D0 U5595 ( .A1(n[778]), .A2(a[8]), .Z(n[1290]) );
  AN2D0 U5596 ( .A1(b[7]), .A2(n[267]), .Z(n[778]) );
  AN2D0 U5597 ( .A1(n[777]), .A2(a[8]), .Z(n[1289]) );
  AN2D0 U5598 ( .A1(b[7]), .A2(n[266]), .Z(n[777]) );
  AN2D0 U5599 ( .A1(n[776]), .A2(a[8]), .Z(n[1288]) );
  AN2D0 U5600 ( .A1(b[7]), .A2(n[265]), .Z(n[776]) );
  AN2D0 U5601 ( .A1(n[773]), .A2(a[8]), .Z(n[1285]) );
  AN2D0 U5602 ( .A1(b[7]), .A2(n[262]), .Z(n[773]) );
  AN2D0 U5603 ( .A1(n[770]), .A2(a[8]), .Z(n[1282]) );
  AN2D0 U5604 ( .A1(b[7]), .A2(n[259]), .Z(n[770]) );
  AN2D0 U5605 ( .A1(n[769]), .A2(a[8]), .Z(n[1281]) );
  AN2D0 U5606 ( .A1(b[7]), .A2(n[258]), .Z(n[769]) );
  AN2D0 U5607 ( .A1(n[766]), .A2(a[8]), .Z(n[1278]) );
  AN2D0 U5608 ( .A1(b[7]), .A2(n[255]), .Z(n[766]) );
  AN2D0 U5609 ( .A1(n[763]), .A2(a[8]), .Z(n[1275]) );
  AN2D0 U5610 ( .A1(b[7]), .A2(n[252]), .Z(n[763]) );
  AN2D0 U5611 ( .A1(n[762]), .A2(a[8]), .Z(n[1274]) );
  AN2D0 U5612 ( .A1(b[7]), .A2(n[251]), .Z(n[762]) );
  AN2D0 U5613 ( .A1(n[761]), .A2(a[8]), .Z(n[1273]) );
  AN2D0 U5614 ( .A1(b[7]), .A2(n[250]), .Z(n[761]) );
  AN2D0 U5615 ( .A1(n[760]), .A2(a[8]), .Z(n[1272]) );
  AN2D0 U5616 ( .A1(b[7]), .A2(n[249]), .Z(n[760]) );
  AN2D0 U5617 ( .A1(n[759]), .A2(a[8]), .Z(n[1271]) );
  AN2D0 U5618 ( .A1(b[7]), .A2(n[248]), .Z(n[759]) );
  AN2D0 U5619 ( .A1(n[758]), .A2(a[8]), .Z(n[1270]) );
  AN2D0 U5620 ( .A1(b[7]), .A2(n[247]), .Z(n[758]) );
  AN2D0 U5621 ( .A1(n[757]), .A2(a[8]), .Z(n[1269]) );
  AN2D0 U5622 ( .A1(b[7]), .A2(n[246]), .Z(n[757]) );
  AN2D0 U5623 ( .A1(n[754]), .A2(a[8]), .Z(n[1266]) );
  AN2D0 U5624 ( .A1(n[498]), .A2(a[7]), .Z(n[754]) );
  AN2D0 U5625 ( .A1(n[751]), .A2(a[8]), .Z(n[1263]) );
  AN2D0 U5626 ( .A1(a[7]), .A2(n[495]), .Z(n[751]) );
  AN2D0 U5627 ( .A1(n[750]), .A2(a[8]), .Z(n[1262]) );
  AN2D0 U5628 ( .A1(a[7]), .A2(n[494]), .Z(n[750]) );
  AN2D0 U5629 ( .A1(n[747]), .A2(a[8]), .Z(n[1259]) );
  AN2D0 U5630 ( .A1(a[7]), .A2(n[491]), .Z(n[747]) );
  AN2D0 U5631 ( .A1(n[744]), .A2(a[8]), .Z(n[1256]) );
  AN2D0 U5632 ( .A1(n[488]), .A2(a[7]), .Z(n[744]) );
  AN2D0 U5633 ( .A1(n[233]), .A2(b[6]), .Z(n[488]) );
  AN2D0 U5634 ( .A1(n[743]), .A2(a[8]), .Z(n[1255]) );
  AN2D0 U5635 ( .A1(n[487]), .A2(a[7]), .Z(n[743]) );
  AN2D0 U5636 ( .A1(b[6]), .A2(n[232]), .Z(n[487]) );
  AN2D0 U5637 ( .A1(n[742]), .A2(a[8]), .Z(n[1254]) );
  AN2D0 U5638 ( .A1(n[486]), .A2(a[7]), .Z(n[742]) );
  AN2D0 U5639 ( .A1(b[6]), .A2(n[231]), .Z(n[486]) );
  AN2D0 U5640 ( .A1(n[739]), .A2(a[8]), .Z(n[1251]) );
  AN2D0 U5641 ( .A1(n[483]), .A2(a[7]), .Z(n[739]) );
  AN2D0 U5642 ( .A1(b[6]), .A2(n[228]), .Z(n[483]) );
  AN2D0 U5643 ( .A1(n[736]), .A2(a[8]), .Z(n[1248]) );
  AN2D0 U5644 ( .A1(n[480]), .A2(a[7]), .Z(n[736]) );
  AN2D0 U5645 ( .A1(b[6]), .A2(n[225]), .Z(n[480]) );
  AN2D0 U5646 ( .A1(n[735]), .A2(a[8]), .Z(n[1247]) );
  AN2D0 U5647 ( .A1(n[479]), .A2(a[7]), .Z(n[735]) );
  AN2D0 U5648 ( .A1(b[6]), .A2(n[224]), .Z(n[479]) );
  AN2D0 U5649 ( .A1(n[732]), .A2(a[8]), .Z(n[1244]) );
  AN2D0 U5650 ( .A1(n[476]), .A2(a[7]), .Z(n[732]) );
  AN2D0 U5651 ( .A1(b[6]), .A2(n[221]), .Z(n[476]) );
  AN2D0 U5652 ( .A1(n[729]), .A2(a[8]), .Z(n[1241]) );
  AN2D0 U5653 ( .A1(n[473]), .A2(a[7]), .Z(n[729]) );
  AN2D0 U5654 ( .A1(b[6]), .A2(n[218]), .Z(n[473]) );
  AN2D0 U5655 ( .A1(n[728]), .A2(a[8]), .Z(n[1240]) );
  AN2D0 U5656 ( .A1(n[472]), .A2(a[7]), .Z(n[728]) );
  AN2D0 U5657 ( .A1(b[6]), .A2(n[217]), .Z(n[472]) );
  AN2D0 U5658 ( .A1(n[727]), .A2(a[8]), .Z(n[1239]) );
  AN2D0 U5659 ( .A1(n[471]), .A2(a[7]), .Z(n[727]) );
  AN2D0 U5660 ( .A1(b[6]), .A2(n[216]), .Z(n[471]) );
  AN2D0 U5661 ( .A1(n[726]), .A2(a[8]), .Z(n[1238]) );
  AN2D0 U5662 ( .A1(n[470]), .A2(a[7]), .Z(n[726]) );
  AN2D0 U5663 ( .A1(b[6]), .A2(n[215]), .Z(n[470]) );
  AN2D0 U5664 ( .A1(n[723]), .A2(a[8]), .Z(n[1235]) );
  AN2D0 U5665 ( .A1(n[467]), .A2(a[7]), .Z(n[723]) );
  AN2D0 U5666 ( .A1(b[6]), .A2(n[212]), .Z(n[467]) );
  AN2D0 U5667 ( .A1(n[720]), .A2(a[8]), .Z(n[1232]) );
  AN2D0 U5668 ( .A1(n[464]), .A2(a[7]), .Z(n[720]) );
  AN2D0 U5669 ( .A1(b[6]), .A2(n[209]), .Z(n[464]) );
  AN2D0 U5670 ( .A1(n[719]), .A2(a[8]), .Z(n[1231]) );
  AN2D0 U5671 ( .A1(n[463]), .A2(a[7]), .Z(n[719]) );
  AN2D0 U5672 ( .A1(b[6]), .A2(n[208]), .Z(n[463]) );
  AN2D0 U5673 ( .A1(n[716]), .A2(a[8]), .Z(n[1228]) );
  AN2D0 U5674 ( .A1(n[460]), .A2(a[7]), .Z(n[716]) );
  AN2D0 U5675 ( .A1(b[6]), .A2(n[205]), .Z(n[460]) );
  AN2D0 U5676 ( .A1(n[713]), .A2(a[8]), .Z(n[1225]) );
  AN2D0 U5677 ( .A1(n[457]), .A2(a[7]), .Z(n[713]) );
  AN2D0 U5678 ( .A1(b[6]), .A2(n[202]), .Z(n[457]) );
  AN2D0 U5679 ( .A1(n[712]), .A2(a[8]), .Z(n[1224]) );
  AN2D0 U5680 ( .A1(n[456]), .A2(a[7]), .Z(n[712]) );
  AN2D0 U5681 ( .A1(b[6]), .A2(n[201]), .Z(n[456]) );
  AN2D0 U5682 ( .A1(n[711]), .A2(a[8]), .Z(n[1223]) );
  AN2D0 U5683 ( .A1(n[455]), .A2(a[7]), .Z(n[711]) );
  AN2D0 U5684 ( .A1(b[6]), .A2(n[200]), .Z(n[455]) );
  AN2D0 U5685 ( .A1(n[708]), .A2(a[8]), .Z(n[1220]) );
  AN2D0 U5686 ( .A1(n[452]), .A2(a[7]), .Z(n[708]) );
  AN2D0 U5687 ( .A1(b[6]), .A2(n[197]), .Z(n[452]) );
  AN2D0 U5688 ( .A1(n[705]), .A2(a[8]), .Z(n[1217]) );
  AN2D0 U5689 ( .A1(n[449]), .A2(a[7]), .Z(n[705]) );
  AN2D0 U5690 ( .A1(b[6]), .A2(n[194]), .Z(n[449]) );
  AN2D0 U5691 ( .A1(n[704]), .A2(a[8]), .Z(n[1216]) );
  AN2D0 U5692 ( .A1(n[448]), .A2(a[7]), .Z(n[704]) );
  AN2D0 U5693 ( .A1(b[6]), .A2(n[193]), .Z(n[448]) );
  AN2D0 U5694 ( .A1(n[701]), .A2(a[8]), .Z(n[1213]) );
  AN2D0 U5695 ( .A1(n[445]), .A2(a[7]), .Z(n[701]) );
  AN2D0 U5696 ( .A1(b[6]), .A2(n[190]), .Z(n[445]) );
  AN2D0 U5697 ( .A1(n[698]), .A2(a[8]), .Z(n[1210]) );
  AN2D0 U5698 ( .A1(n[442]), .A2(a[7]), .Z(n[698]) );
  AN2D0 U5699 ( .A1(b[6]), .A2(n[187]), .Z(n[442]) );
  AN2D0 U5700 ( .A1(n[697]), .A2(a[8]), .Z(n[1209]) );
  AN2D0 U5701 ( .A1(n[441]), .A2(a[7]), .Z(n[697]) );
  AN2D0 U5702 ( .A1(b[6]), .A2(n[186]), .Z(n[441]) );
  AN2D0 U5703 ( .A1(n[696]), .A2(a[8]), .Z(n[1208]) );
  AN2D0 U5704 ( .A1(n[440]), .A2(a[7]), .Z(n[696]) );
  AN2D0 U5705 ( .A1(b[6]), .A2(n[185]), .Z(n[440]) );
  AN2D0 U5706 ( .A1(n[695]), .A2(a[8]), .Z(n[1207]) );
  AN2D0 U5707 ( .A1(n[439]), .A2(a[7]), .Z(n[695]) );
  AN2D0 U5708 ( .A1(b[6]), .A2(n[184]), .Z(n[439]) );
  AN2D0 U5709 ( .A1(n[694]), .A2(a[8]), .Z(n[1206]) );
  AN2D0 U5710 ( .A1(n[438]), .A2(a[7]), .Z(n[694]) );
  AN2D0 U5711 ( .A1(b[6]), .A2(n[183]), .Z(n[438]) );
  AN2D0 U5712 ( .A1(n[691]), .A2(a[8]), .Z(n[1203]) );
  AN2D0 U5713 ( .A1(n[435]), .A2(a[7]), .Z(n[691]) );
  AN2D0 U5714 ( .A1(b[6]), .A2(n[180]), .Z(n[435]) );
  AN2D0 U5715 ( .A1(n[688]), .A2(a[8]), .Z(n[1200]) );
  AN2D0 U5716 ( .A1(n[432]), .A2(a[7]), .Z(n[688]) );
  AN2D0 U5717 ( .A1(b[6]), .A2(n[177]), .Z(n[432]) );
  AN2D0 U5718 ( .A1(n[687]), .A2(a[8]), .Z(n[1199]) );
  AN2D0 U5719 ( .A1(n[431]), .A2(a[7]), .Z(n[687]) );
  AN2D0 U5720 ( .A1(b[6]), .A2(n[176]), .Z(n[431]) );
  AN2D0 U5721 ( .A1(n[684]), .A2(a[8]), .Z(n[1196]) );
  AN2D0 U5722 ( .A1(n[428]), .A2(a[7]), .Z(n[684]) );
  AN2D0 U5723 ( .A1(b[6]), .A2(n[173]), .Z(n[428]) );
  AN2D0 U5724 ( .A1(n[681]), .A2(a[8]), .Z(n[1193]) );
  AN2D0 U5725 ( .A1(n[425]), .A2(a[7]), .Z(n[681]) );
  AN2D0 U5726 ( .A1(b[6]), .A2(n[170]), .Z(n[425]) );
  AN2D0 U5727 ( .A1(n[680]), .A2(a[8]), .Z(n[1192]) );
  AN2D0 U5728 ( .A1(n[424]), .A2(a[7]), .Z(n[680]) );
  AN2D0 U5729 ( .A1(b[6]), .A2(n[169]), .Z(n[424]) );
  AN2D0 U5730 ( .A1(n[679]), .A2(a[8]), .Z(n[1191]) );
  AN2D0 U5731 ( .A1(n[423]), .A2(a[7]), .Z(n[679]) );
  AN2D0 U5732 ( .A1(b[6]), .A2(n[168]), .Z(n[423]) );
  AN2D0 U5733 ( .A1(n[676]), .A2(a[8]), .Z(n[1188]) );
  AN2D0 U5734 ( .A1(n[420]), .A2(a[7]), .Z(n[676]) );
  AN2D0 U5735 ( .A1(b[6]), .A2(n[165]), .Z(n[420]) );
  AN2D0 U5736 ( .A1(n[673]), .A2(a[8]), .Z(n[1185]) );
  AN2D0 U5737 ( .A1(n[417]), .A2(a[7]), .Z(n[673]) );
  AN2D0 U5738 ( .A1(b[6]), .A2(n[162]), .Z(n[417]) );
  AN2D0 U5739 ( .A1(n[672]), .A2(a[8]), .Z(n[1184]) );
  AN2D0 U5740 ( .A1(n[416]), .A2(a[7]), .Z(n[672]) );
  AN2D0 U5741 ( .A1(b[6]), .A2(n[161]), .Z(n[416]) );
  AN2D0 U5742 ( .A1(n[669]), .A2(a[8]), .Z(n[1181]) );
  AN2D0 U5743 ( .A1(n[413]), .A2(a[7]), .Z(n[669]) );
  AN2D0 U5744 ( .A1(b[6]), .A2(n[158]), .Z(n[413]) );
  AN2D0 U5745 ( .A1(n[666]), .A2(a[8]), .Z(n[1178]) );
  AN2D0 U5746 ( .A1(n[410]), .A2(a[7]), .Z(n[666]) );
  AN2D0 U5747 ( .A1(b[6]), .A2(n[155]), .Z(n[410]) );
  AN2D0 U5748 ( .A1(n[665]), .A2(a[8]), .Z(n[1177]) );
  AN2D0 U5749 ( .A1(n[409]), .A2(a[7]), .Z(n[665]) );
  AN2D0 U5750 ( .A1(b[6]), .A2(n[154]), .Z(n[409]) );
  AN2D0 U5751 ( .A1(n[664]), .A2(a[8]), .Z(n[1176]) );
  AN2D0 U5752 ( .A1(n[408]), .A2(a[7]), .Z(n[664]) );
  AN2D0 U5753 ( .A1(b[6]), .A2(n[153]), .Z(n[408]) );
  AN2D0 U5754 ( .A1(n[663]), .A2(a[8]), .Z(n[1175]) );
  AN2D0 U5755 ( .A1(n[407]), .A2(a[7]), .Z(n[663]) );
  AN2D0 U5756 ( .A1(b[6]), .A2(n[152]), .Z(n[407]) );
  AN2D0 U5757 ( .A1(n[660]), .A2(a[8]), .Z(n[1172]) );
  AN2D0 U5758 ( .A1(n[404]), .A2(a[7]), .Z(n[660]) );
  AN2D0 U5759 ( .A1(b[6]), .A2(n[149]), .Z(n[404]) );
  AN2D0 U5760 ( .A1(n[657]), .A2(a[8]), .Z(n[1169]) );
  AN2D0 U5761 ( .A1(n[401]), .A2(a[7]), .Z(n[657]) );
  AN2D0 U5762 ( .A1(b[6]), .A2(n[146]), .Z(n[401]) );
  AN2D0 U5763 ( .A1(n[656]), .A2(a[8]), .Z(n[1168]) );
  AN2D0 U5764 ( .A1(n[400]), .A2(a[7]), .Z(n[656]) );
  AN2D0 U5765 ( .A1(b[6]), .A2(n[145]), .Z(n[400]) );
  AN2D0 U5766 ( .A1(n[653]), .A2(a[8]), .Z(n[1165]) );
  AN2D0 U5767 ( .A1(n[397]), .A2(a[7]), .Z(n[653]) );
  AN2D0 U5768 ( .A1(b[6]), .A2(n[142]), .Z(n[397]) );
  AN2D0 U5769 ( .A1(n[650]), .A2(a[8]), .Z(n[1162]) );
  AN2D0 U5770 ( .A1(n[394]), .A2(a[7]), .Z(n[650]) );
  AN2D0 U5771 ( .A1(b[6]), .A2(n[139]), .Z(n[394]) );
  AN2D0 U5772 ( .A1(n[649]), .A2(a[8]), .Z(n[1161]) );
  AN2D0 U5773 ( .A1(n[393]), .A2(a[7]), .Z(n[649]) );
  AN2D0 U5774 ( .A1(b[6]), .A2(n[138]), .Z(n[393]) );
  AN2D0 U5775 ( .A1(n[648]), .A2(a[8]), .Z(n[1160]) );
  AN2D0 U5776 ( .A1(n[392]), .A2(a[7]), .Z(n[648]) );
  AN2D0 U5777 ( .A1(b[6]), .A2(n[137]), .Z(n[392]) );
  AN2D0 U5778 ( .A1(n[645]), .A2(a[8]), .Z(n[1157]) );
  AN2D0 U5779 ( .A1(n[389]), .A2(a[7]), .Z(n[645]) );
  AN2D0 U5780 ( .A1(b[6]), .A2(n[134]), .Z(n[389]) );
  AN2D0 U5781 ( .A1(n[642]), .A2(a[8]), .Z(n[1154]) );
  AN2D0 U5782 ( .A1(n[386]), .A2(a[7]), .Z(n[642]) );
  AN2D0 U5783 ( .A1(b[6]), .A2(n[131]), .Z(n[386]) );
  AN2D0 U5784 ( .A1(n[641]), .A2(a[8]), .Z(n[1153]) );
  AN2D0 U5785 ( .A1(n[385]), .A2(a[7]), .Z(n[641]) );
  AN2D0 U5786 ( .A1(b[6]), .A2(n[130]), .Z(n[385]) );
  AN2D0 U5787 ( .A1(n[638]), .A2(a[8]), .Z(n[1150]) );
  AN2D0 U5788 ( .A1(n[382]), .A2(a[7]), .Z(n[638]) );
  AN2D0 U5789 ( .A1(b[6]), .A2(n[127]), .Z(n[382]) );
  AN2D0 U5790 ( .A1(n[635]), .A2(a[8]), .Z(n[1147]) );
  AN2D0 U5791 ( .A1(n[379]), .A2(a[7]), .Z(n[635]) );
  AN2D0 U5792 ( .A1(b[6]), .A2(n[124]), .Z(n[379]) );
  AN2D0 U5793 ( .A1(n[634]), .A2(a[8]), .Z(n[1146]) );
  AN2D0 U5794 ( .A1(n[378]), .A2(a[7]), .Z(n[634]) );
  AN2D0 U5795 ( .A1(b[6]), .A2(n[123]), .Z(n[378]) );
  AN2D0 U5796 ( .A1(n[633]), .A2(a[8]), .Z(n[1145]) );
  AN2D0 U5797 ( .A1(n[377]), .A2(a[7]), .Z(n[633]) );
  AN2D0 U5798 ( .A1(b[6]), .A2(n[122]), .Z(n[377]) );
  AN2D0 U5799 ( .A1(n[632]), .A2(a[8]), .Z(n[1144]) );
  AN2D0 U5800 ( .A1(n[376]), .A2(a[7]), .Z(n[632]) );
  AN2D0 U5801 ( .A1(b[6]), .A2(n[121]), .Z(n[376]) );
  AN2D0 U5802 ( .A1(n[631]), .A2(a[8]), .Z(n[1143]) );
  AN2D0 U5803 ( .A1(n[375]), .A2(a[7]), .Z(n[631]) );
  AN2D0 U5804 ( .A1(b[6]), .A2(n[120]), .Z(n[375]) );
  AN2D0 U5805 ( .A1(n[630]), .A2(a[8]), .Z(n[1142]) );
  AN2D0 U5806 ( .A1(n[374]), .A2(a[7]), .Z(n[630]) );
  AN2D0 U5807 ( .A1(b[6]), .A2(n[119]), .Z(n[374]) );
  AN2D0 U5808 ( .A1(n[627]), .A2(a[8]), .Z(n[1139]) );
  AN2D0 U5809 ( .A1(n[371]), .A2(a[7]), .Z(n[627]) );
  AN2D0 U5810 ( .A1(n[243]), .A2(a[6]), .Z(n[371]) );
  AN2D0 U5811 ( .A1(n[624]), .A2(a[8]), .Z(n[1136]) );
  AN2D0 U5812 ( .A1(n[368]), .A2(a[7]), .Z(n[624]) );
  AN2D0 U5813 ( .A1(a[6]), .A2(n[240]), .Z(n[368]) );
  AN2D0 U5814 ( .A1(n[623]), .A2(a[8]), .Z(n[1135]) );
  AN2D0 U5815 ( .A1(n[367]), .A2(a[7]), .Z(n[623]) );
  AN2D0 U5816 ( .A1(a[6]), .A2(n[239]), .Z(n[367]) );
  AN2D0 U5817 ( .A1(n[620]), .A2(a[8]), .Z(n[1132]) );
  AN2D0 U5818 ( .A1(n[364]), .A2(a[7]), .Z(n[620]) );
  AN2D0 U5819 ( .A1(a[6]), .A2(n[236]), .Z(n[364]) );
  AN2D0 U5820 ( .A1(n[617]), .A2(a[8]), .Z(n[1129]) );
  AN2D0 U5821 ( .A1(n[361]), .A2(a[7]), .Z(n[617]) );
  AN2D0 U5822 ( .A1(n[233]), .A2(a[6]), .Z(n[361]) );
  AN2D0 U5823 ( .A1(n[106]), .A2(b[5]), .Z(n[233]) );
  AN2D0 U5824 ( .A1(n[616]), .A2(a[8]), .Z(n[1128]) );
  AN2D0 U5825 ( .A1(n[360]), .A2(a[7]), .Z(n[616]) );
  AN2D0 U5826 ( .A1(n[232]), .A2(a[6]), .Z(n[360]) );
  AN2D0 U5827 ( .A1(b[5]), .A2(n[105]), .Z(n[232]) );
  AN2D0 U5828 ( .A1(n[615]), .A2(a[8]), .Z(n[1127]) );
  AN2D0 U5829 ( .A1(n[359]), .A2(a[7]), .Z(n[615]) );
  AN2D0 U5830 ( .A1(n[231]), .A2(a[6]), .Z(n[359]) );
  AN2D0 U5831 ( .A1(b[5]), .A2(n[104]), .Z(n[231]) );
  AN2D0 U5832 ( .A1(n[612]), .A2(a[8]), .Z(n[1124]) );
  AN2D0 U5833 ( .A1(n[356]), .A2(a[7]), .Z(n[612]) );
  AN2D0 U5834 ( .A1(n[228]), .A2(a[6]), .Z(n[356]) );
  AN2D0 U5835 ( .A1(b[5]), .A2(n[101]), .Z(n[228]) );
  AN2D0 U5836 ( .A1(n[609]), .A2(a[8]), .Z(n[1121]) );
  AN2D0 U5837 ( .A1(n[353]), .A2(a[7]), .Z(n[609]) );
  AN2D0 U5838 ( .A1(n[225]), .A2(a[6]), .Z(n[353]) );
  AN2D0 U5839 ( .A1(b[5]), .A2(n[98]), .Z(n[225]) );
  AN2D0 U5840 ( .A1(n[608]), .A2(a[8]), .Z(n[1120]) );
  AN2D0 U5841 ( .A1(n[352]), .A2(a[7]), .Z(n[608]) );
  AN2D0 U5842 ( .A1(n[224]), .A2(a[6]), .Z(n[352]) );
  AN2D0 U5843 ( .A1(b[5]), .A2(n[97]), .Z(n[224]) );
  AN2D0 U5844 ( .A1(n[605]), .A2(a[8]), .Z(n[1117]) );
  AN2D0 U5845 ( .A1(n[349]), .A2(a[7]), .Z(n[605]) );
  AN2D0 U5846 ( .A1(n[221]), .A2(a[6]), .Z(n[349]) );
  AN2D0 U5847 ( .A1(b[5]), .A2(n[94]), .Z(n[221]) );
  AN2D0 U5848 ( .A1(n[602]), .A2(a[8]), .Z(n[1114]) );
  AN2D0 U5849 ( .A1(n[346]), .A2(a[7]), .Z(n[602]) );
  AN2D0 U5850 ( .A1(n[218]), .A2(a[6]), .Z(n[346]) );
  AN2D0 U5851 ( .A1(b[5]), .A2(n[91]), .Z(n[218]) );
  AN2D0 U5852 ( .A1(n[601]), .A2(a[8]), .Z(n[1113]) );
  AN2D0 U5853 ( .A1(n[345]), .A2(a[7]), .Z(n[601]) );
  AN2D0 U5854 ( .A1(n[217]), .A2(a[6]), .Z(n[345]) );
  AN2D0 U5855 ( .A1(b[5]), .A2(n[90]), .Z(n[217]) );
  AN2D0 U5856 ( .A1(n[600]), .A2(a[8]), .Z(n[1112]) );
  AN2D0 U5857 ( .A1(n[344]), .A2(a[7]), .Z(n[600]) );
  AN2D0 U5858 ( .A1(n[216]), .A2(a[6]), .Z(n[344]) );
  AN2D0 U5859 ( .A1(b[5]), .A2(n[89]), .Z(n[216]) );
  AN2D0 U5860 ( .A1(n[599]), .A2(a[8]), .Z(n[1111]) );
  AN2D0 U5861 ( .A1(n[343]), .A2(a[7]), .Z(n[599]) );
  AN2D0 U5862 ( .A1(n[215]), .A2(a[6]), .Z(n[343]) );
  AN2D0 U5863 ( .A1(b[5]), .A2(n[88]), .Z(n[215]) );
  AN2D0 U5864 ( .A1(n[596]), .A2(a[8]), .Z(n[1108]) );
  AN2D0 U5865 ( .A1(n[340]), .A2(a[7]), .Z(n[596]) );
  AN2D0 U5866 ( .A1(n[212]), .A2(a[6]), .Z(n[340]) );
  AN2D0 U5867 ( .A1(b[5]), .A2(n[85]), .Z(n[212]) );
  AN2D0 U5868 ( .A1(n[593]), .A2(a[8]), .Z(n[1105]) );
  AN2D0 U5869 ( .A1(n[337]), .A2(a[7]), .Z(n[593]) );
  AN2D0 U5870 ( .A1(n[209]), .A2(a[6]), .Z(n[337]) );
  AN2D0 U5871 ( .A1(b[5]), .A2(n[82]), .Z(n[209]) );
  AN2D0 U5872 ( .A1(n[592]), .A2(a[8]), .Z(n[1104]) );
  AN2D0 U5873 ( .A1(n[336]), .A2(a[7]), .Z(n[592]) );
  AN2D0 U5874 ( .A1(n[208]), .A2(a[6]), .Z(n[336]) );
  AN2D0 U5875 ( .A1(b[5]), .A2(n[81]), .Z(n[208]) );
  AN2D0 U5876 ( .A1(n[589]), .A2(a[8]), .Z(n[1101]) );
  AN2D0 U5877 ( .A1(n[333]), .A2(a[7]), .Z(n[589]) );
  AN2D0 U5878 ( .A1(n[205]), .A2(a[6]), .Z(n[333]) );
  AN2D0 U5879 ( .A1(b[5]), .A2(n[78]), .Z(n[205]) );
  AN2D0 U5880 ( .A1(n[586]), .A2(a[8]), .Z(n[1098]) );
  AN2D0 U5881 ( .A1(n[330]), .A2(a[7]), .Z(n[586]) );
  AN2D0 U5882 ( .A1(n[202]), .A2(a[6]), .Z(n[330]) );
  AN2D0 U5883 ( .A1(b[5]), .A2(n[75]), .Z(n[202]) );
  AN2D0 U5884 ( .A1(n[585]), .A2(a[8]), .Z(n[1097]) );
  AN2D0 U5885 ( .A1(n[329]), .A2(a[7]), .Z(n[585]) );
  AN2D0 U5886 ( .A1(n[201]), .A2(a[6]), .Z(n[329]) );
  AN2D0 U5887 ( .A1(b[5]), .A2(n[74]), .Z(n[201]) );
  AN2D0 U5888 ( .A1(n[584]), .A2(a[8]), .Z(n[1096]) );
  AN2D0 U5889 ( .A1(n[328]), .A2(a[7]), .Z(n[584]) );
  AN2D0 U5890 ( .A1(n[200]), .A2(a[6]), .Z(n[328]) );
  AN2D0 U5891 ( .A1(b[5]), .A2(n[73]), .Z(n[200]) );
  AN2D0 U5892 ( .A1(n[581]), .A2(a[8]), .Z(n[1093]) );
  AN2D0 U5893 ( .A1(n[325]), .A2(a[7]), .Z(n[581]) );
  AN2D0 U5894 ( .A1(n[197]), .A2(a[6]), .Z(n[325]) );
  AN2D0 U5895 ( .A1(b[5]), .A2(n[70]), .Z(n[197]) );
  AN2D0 U5896 ( .A1(n[578]), .A2(a[8]), .Z(n[1090]) );
  AN2D0 U5897 ( .A1(n[322]), .A2(a[7]), .Z(n[578]) );
  AN2D0 U5898 ( .A1(n[194]), .A2(a[6]), .Z(n[322]) );
  AN2D0 U5899 ( .A1(b[5]), .A2(n[67]), .Z(n[194]) );
  AN2D0 U5900 ( .A1(n[577]), .A2(a[8]), .Z(n[1089]) );
  AN2D0 U5901 ( .A1(n[321]), .A2(a[7]), .Z(n[577]) );
  AN2D0 U5902 ( .A1(n[193]), .A2(a[6]), .Z(n[321]) );
  AN2D0 U5903 ( .A1(b[5]), .A2(n[66]), .Z(n[193]) );
  AN2D0 U5904 ( .A1(n[574]), .A2(a[8]), .Z(n[1086]) );
  AN2D0 U5905 ( .A1(n[318]), .A2(a[7]), .Z(n[574]) );
  AN2D0 U5906 ( .A1(n[190]), .A2(a[6]), .Z(n[318]) );
  AN2D0 U5907 ( .A1(b[5]), .A2(n[63]), .Z(n[190]) );
  AN2D0 U5908 ( .A1(n[571]), .A2(a[8]), .Z(n[1083]) );
  AN2D0 U5909 ( .A1(n[315]), .A2(a[7]), .Z(n[571]) );
  AN2D0 U5910 ( .A1(n[187]), .A2(a[6]), .Z(n[315]) );
  AN2D0 U5911 ( .A1(b[5]), .A2(n[60]), .Z(n[187]) );
  AN2D0 U5912 ( .A1(n[570]), .A2(a[8]), .Z(n[1082]) );
  AN2D0 U5913 ( .A1(n[314]), .A2(a[7]), .Z(n[570]) );
  AN2D0 U5914 ( .A1(n[186]), .A2(a[6]), .Z(n[314]) );
  AN2D0 U5915 ( .A1(b[5]), .A2(n[59]), .Z(n[186]) );
  AN2D0 U5916 ( .A1(n[569]), .A2(a[8]), .Z(n[1081]) );
  AN2D0 U5917 ( .A1(n[313]), .A2(a[7]), .Z(n[569]) );
  AN2D0 U5918 ( .A1(n[185]), .A2(a[6]), .Z(n[313]) );
  AN2D0 U5919 ( .A1(b[5]), .A2(n[58]), .Z(n[185]) );
  AN2D0 U5920 ( .A1(n[568]), .A2(a[8]), .Z(n[1080]) );
  AN2D0 U5921 ( .A1(n[312]), .A2(a[7]), .Z(n[568]) );
  AN2D0 U5922 ( .A1(n[184]), .A2(a[6]), .Z(n[312]) );
  AN2D0 U5923 ( .A1(b[5]), .A2(n[57]), .Z(n[184]) );
  AN2D0 U5924 ( .A1(n[567]), .A2(a[8]), .Z(n[1079]) );
  AN2D0 U5925 ( .A1(n[311]), .A2(a[7]), .Z(n[567]) );
  AN2D0 U5926 ( .A1(n[183]), .A2(a[6]), .Z(n[311]) );
  AN2D0 U5927 ( .A1(b[5]), .A2(n[56]), .Z(n[183]) );
  AN2D0 U5928 ( .A1(n[564]), .A2(a[8]), .Z(n[1076]) );
  AN2D0 U5929 ( .A1(n[308]), .A2(a[7]), .Z(n[564]) );
  AN2D0 U5930 ( .A1(n[180]), .A2(a[6]), .Z(n[308]) );
  AN2D0 U5931 ( .A1(n[116]), .A2(a[5]), .Z(n[180]) );
  AN2D0 U5932 ( .A1(n[561]), .A2(a[8]), .Z(n[1073]) );
  AN2D0 U5933 ( .A1(n[305]), .A2(a[7]), .Z(n[561]) );
  AN2D0 U5934 ( .A1(n[177]), .A2(a[6]), .Z(n[305]) );
  AN2D0 U5935 ( .A1(a[5]), .A2(n[113]), .Z(n[177]) );
  AN2D0 U5936 ( .A1(n[560]), .A2(a[8]), .Z(n[1072]) );
  AN2D0 U5937 ( .A1(n[304]), .A2(a[7]), .Z(n[560]) );
  AN2D0 U5938 ( .A1(n[176]), .A2(a[6]), .Z(n[304]) );
  AN2D0 U5939 ( .A1(a[5]), .A2(n[112]), .Z(n[176]) );
  AN2D0 U5940 ( .A1(n[557]), .A2(a[8]), .Z(n[1069]) );
  AN2D0 U5941 ( .A1(n[301]), .A2(a[7]), .Z(n[557]) );
  AN2D0 U5942 ( .A1(n[173]), .A2(a[6]), .Z(n[301]) );
  AN2D0 U5943 ( .A1(a[5]), .A2(n[109]), .Z(n[173]) );
  AN2D0 U5944 ( .A1(n[554]), .A2(a[8]), .Z(n[1066]) );
  AN2D0 U5945 ( .A1(n[298]), .A2(a[7]), .Z(n[554]) );
  AN2D0 U5946 ( .A1(n[170]), .A2(a[6]), .Z(n[298]) );
  AN2D0 U5947 ( .A1(n[106]), .A2(a[5]), .Z(n[170]) );
  AN2D0 U5948 ( .A1(n[43]), .A2(b[4]), .Z(n[106]) );
  AN2D0 U5949 ( .A1(n[553]), .A2(a[8]), .Z(n[1065]) );
  AN2D0 U5950 ( .A1(n[297]), .A2(a[7]), .Z(n[553]) );
  AN2D0 U5951 ( .A1(n[169]), .A2(a[6]), .Z(n[297]) );
  AN2D0 U5952 ( .A1(n[105]), .A2(a[5]), .Z(n[169]) );
  AN2D0 U5953 ( .A1(n[552]), .A2(a[8]), .Z(n[1064]) );
  AN2D0 U5954 ( .A1(n[296]), .A2(a[7]), .Z(n[552]) );
  AN2D0 U5955 ( .A1(n[168]), .A2(a[6]), .Z(n[296]) );
  AN2D0 U5956 ( .A1(n[104]), .A2(a[5]), .Z(n[168]) );
  AN2D0 U5957 ( .A1(n[549]), .A2(a[8]), .Z(n[1061]) );
  AN2D0 U5958 ( .A1(n[293]), .A2(a[7]), .Z(n[549]) );
  AN2D0 U5959 ( .A1(n[165]), .A2(a[6]), .Z(n[293]) );
  AN2D0 U5960 ( .A1(n[101]), .A2(a[5]), .Z(n[165]) );
  AN2D0 U5961 ( .A1(b[4]), .A2(n[42]), .Z(n[105]) );
  AN2D0 U5962 ( .A1(n[546]), .A2(a[8]), .Z(n[1058]) );
  AN2D0 U5963 ( .A1(n[290]), .A2(a[7]), .Z(n[546]) );
  AN2D0 U5964 ( .A1(n[162]), .A2(a[6]), .Z(n[290]) );
  AN2D0 U5965 ( .A1(n[98]), .A2(a[5]), .Z(n[162]) );
  AN2D0 U5966 ( .A1(b[4]), .A2(n[35]), .Z(n[98]) );
  AN2D0 U5967 ( .A1(n[545]), .A2(a[8]), .Z(n[1057]) );
  AN2D0 U5968 ( .A1(n[289]), .A2(a[7]), .Z(n[545]) );
  AN2D0 U5969 ( .A1(n[161]), .A2(a[6]), .Z(n[289]) );
  AN2D0 U5970 ( .A1(n[97]), .A2(a[5]), .Z(n[161]) );
  AN2D0 U5971 ( .A1(b[4]), .A2(n[34]), .Z(n[97]) );
  AN2D0 U5972 ( .A1(n[542]), .A2(a[8]), .Z(n[1054]) );
  AN2D0 U5973 ( .A1(n[286]), .A2(a[7]), .Z(n[542]) );
  AN2D0 U5974 ( .A1(n[158]), .A2(a[6]), .Z(n[286]) );
  AN2D0 U5975 ( .A1(n[94]), .A2(a[5]), .Z(n[158]) );
  AN2D0 U5976 ( .A1(b[4]), .A2(n[31]), .Z(n[94]) );
  AN2D0 U5977 ( .A1(n[539]), .A2(a[8]), .Z(n[1051]) );
  AN2D0 U5978 ( .A1(n[283]), .A2(a[7]), .Z(n[539]) );
  AN2D0 U5979 ( .A1(n[155]), .A2(a[6]), .Z(n[283]) );
  AN2D0 U5980 ( .A1(n[91]), .A2(a[5]), .Z(n[155]) );
  AN2D0 U5981 ( .A1(b[4]), .A2(n[28]), .Z(n[91]) );
  AN2D0 U5982 ( .A1(n[538]), .A2(a[8]), .Z(n[1050]) );
  AN2D0 U5983 ( .A1(n[282]), .A2(a[7]), .Z(n[538]) );
  AN2D0 U5984 ( .A1(n[154]), .A2(a[6]), .Z(n[282]) );
  AN2D0 U5985 ( .A1(n[90]), .A2(a[5]), .Z(n[154]) );
  AN2D0 U5986 ( .A1(b[4]), .A2(n[27]), .Z(n[90]) );
  AN2D0 U5987 ( .A1(b[4]), .A2(n[41]), .Z(n[104]) );
  AN2D0 U5988 ( .A1(n[537]), .A2(a[8]), .Z(n[1049]) );
  AN2D0 U5989 ( .A1(n[281]), .A2(a[7]), .Z(n[537]) );
  AN2D0 U5990 ( .A1(n[153]), .A2(a[6]), .Z(n[281]) );
  AN2D0 U5991 ( .A1(n[89]), .A2(a[5]), .Z(n[153]) );
  AN2D0 U5992 ( .A1(b[4]), .A2(n[26]), .Z(n[89]) );
  AN2D0 U5993 ( .A1(n[536]), .A2(a[8]), .Z(n[1048]) );
  AN2D0 U5994 ( .A1(n[280]), .A2(a[7]), .Z(n[536]) );
  AN2D0 U5995 ( .A1(n[152]), .A2(a[6]), .Z(n[280]) );
  AN2D0 U5996 ( .A1(n[88]), .A2(a[5]), .Z(n[152]) );
  AN2D0 U5997 ( .A1(b[4]), .A2(n[25]), .Z(n[88]) );
  AN2D0 U5998 ( .A1(n[533]), .A2(a[8]), .Z(n[1045]) );
  AN2D0 U5999 ( .A1(n[277]), .A2(a[7]), .Z(n[533]) );
  AN2D0 U6000 ( .A1(n[149]), .A2(a[6]), .Z(n[277]) );
  AN2D0 U6001 ( .A1(n[85]), .A2(a[5]), .Z(n[149]) );
  AN2D0 U6002 ( .A1(n[53]), .A2(a[4]), .Z(n[85]) );
  AN2D0 U6003 ( .A1(n[530]), .A2(a[8]), .Z(n[1042]) );
  AN2D0 U6004 ( .A1(n[274]), .A2(a[7]), .Z(n[530]) );
  AN2D0 U6005 ( .A1(n[146]), .A2(a[6]), .Z(n[274]) );
  AN2D0 U6006 ( .A1(n[82]), .A2(a[5]), .Z(n[146]) );
  AN2D0 U6007 ( .A1(a[4]), .A2(n[50]), .Z(n[82]) );
  AN2D0 U6008 ( .A1(n[529]), .A2(a[8]), .Z(n[1041]) );
  AN2D0 U6009 ( .A1(n[273]), .A2(a[7]), .Z(n[529]) );
  AN2D0 U6010 ( .A1(n[145]), .A2(a[6]), .Z(n[273]) );
  AN2D0 U6011 ( .A1(n[81]), .A2(a[5]), .Z(n[145]) );
  AN2D0 U6012 ( .A1(a[4]), .A2(n[49]), .Z(n[81]) );
  AN2D0 U6013 ( .A1(n[526]), .A2(a[8]), .Z(n[1038]) );
  AN2D0 U6014 ( .A1(n[270]), .A2(a[7]), .Z(n[526]) );
  AN2D0 U6015 ( .A1(n[142]), .A2(a[6]), .Z(n[270]) );
  AN2D0 U6016 ( .A1(n[78]), .A2(a[5]), .Z(n[142]) );
  AN2D0 U6017 ( .A1(a[4]), .A2(n[46]), .Z(n[78]) );
  AN2D0 U6018 ( .A1(n[523]), .A2(a[8]), .Z(n[1035]) );
  AN2D0 U6019 ( .A1(n[267]), .A2(a[7]), .Z(n[523]) );
  AN2D0 U6020 ( .A1(n[139]), .A2(a[6]), .Z(n[267]) );
  AN2D0 U6021 ( .A1(n[75]), .A2(a[5]), .Z(n[139]) );
  AN2D0 U6022 ( .A1(n[43]), .A2(a[4]), .Z(n[75]) );
  AN2D0 U6023 ( .A1(n[12]), .A2(b[3]), .Z(n[43]) );
  AN2D0 U6024 ( .A1(n[522]), .A2(a[8]), .Z(n[1034]) );
  AN2D0 U6025 ( .A1(n[266]), .A2(a[7]), .Z(n[522]) );
  AN2D0 U6026 ( .A1(n[138]), .A2(a[6]), .Z(n[266]) );
  AN2D0 U6027 ( .A1(n[74]), .A2(a[5]), .Z(n[138]) );
  AN2D0 U6028 ( .A1(n[42]), .A2(a[4]), .Z(n[74]) );
  AN2D0 U6029 ( .A1(b[3]), .A2(n[11]), .Z(n[42]) );
  AN2D0 U6030 ( .A1(n[521]), .A2(a[8]), .Z(n[1033]) );
  AN2D0 U6031 ( .A1(n[265]), .A2(a[7]), .Z(n[521]) );
  AN2D0 U6032 ( .A1(n[137]), .A2(a[6]), .Z(n[265]) );
  AN2D0 U6033 ( .A1(n[73]), .A2(a[5]), .Z(n[137]) );
  AN2D0 U6034 ( .A1(n[41]), .A2(a[4]), .Z(n[73]) );
  AN2D0 U6035 ( .A1(b[3]), .A2(n[10]), .Z(n[41]) );
  AN2D0 U6036 ( .A1(n[518]), .A2(a[8]), .Z(n[1030]) );
  AN2D0 U6037 ( .A1(n[262]), .A2(a[7]), .Z(n[518]) );
  AN2D0 U6038 ( .A1(n[134]), .A2(a[6]), .Z(n[262]) );
  AN2D0 U6039 ( .A1(n[70]), .A2(a[5]), .Z(n[134]) );
  AN2D0 U6040 ( .A1(n[38]), .A2(a[4]), .Z(n[70]) );
  AN2D0 U6041 ( .A1(n[515]), .A2(a[8]), .Z(n[1027]) );
  AN2D0 U6042 ( .A1(n[259]), .A2(a[7]), .Z(n[515]) );
  AN2D0 U6043 ( .A1(n[131]), .A2(a[6]), .Z(n[259]) );
  AN2D0 U6044 ( .A1(n[67]), .A2(a[5]), .Z(n[131]) );
  AN2D0 U6045 ( .A1(n[35]), .A2(a[4]), .Z(n[67]) );
  AN2D0 U6046 ( .A1(a[3]), .A2(n[19]), .Z(n[35]) );
  AN2D0 U6047 ( .A1(n[514]), .A2(a[8]), .Z(n[1026]) );
  AN2D0 U6048 ( .A1(n[258]), .A2(a[7]), .Z(n[514]) );
  AN2D0 U6049 ( .A1(n[130]), .A2(a[6]), .Z(n[258]) );
  AN2D0 U6050 ( .A1(n[66]), .A2(a[5]), .Z(n[130]) );
  AN2D0 U6051 ( .A1(n[34]), .A2(a[4]), .Z(n[66]) );
  AN2D0 U6052 ( .A1(a[3]), .A2(n[18]), .Z(n[34]) );
  AN2D0 U6053 ( .A1(n[511]), .A2(a[8]), .Z(n[1023]) );
  AN2D0 U6054 ( .A1(n[255]), .A2(a[7]), .Z(n[511]) );
  AN2D0 U6055 ( .A1(n[127]), .A2(a[6]), .Z(n[255]) );
  AN2D0 U6056 ( .A1(n[63]), .A2(a[5]), .Z(n[127]) );
  AN2D0 U6057 ( .A1(n[31]), .A2(a[4]), .Z(n[63]) );
  AN2D0 U6058 ( .A1(a[3]), .A2(n[15]), .Z(n[31]) );
  AN2D0 U6059 ( .A1(n[508]), .A2(a[8]), .Z(n[1020]) );
  AN2D0 U6060 ( .A1(n[252]), .A2(a[7]), .Z(n[508]) );
  AN2D0 U6061 ( .A1(n[124]), .A2(a[6]), .Z(n[252]) );
  AN2D0 U6062 ( .A1(n[60]), .A2(a[5]), .Z(n[124]) );
  AN2D0 U6063 ( .A1(n[28]), .A2(a[4]), .Z(n[60]) );
  AN2D0 U6064 ( .A1(n[12]), .A2(a[3]), .Z(n[28]) );
  AN2D0 U6065 ( .A1(n[4]), .A2(a[2]), .Z(n[12]) );
  AN2D0 U6066 ( .A1(b[4]), .A2(n[38]), .Z(n[101]) );
  AN2D0 U6067 ( .A1(n[22]), .A2(a[3]), .Z(n[38]) );
  AN2D0 U6068 ( .A1(n[507]), .A2(a[8]), .Z(n[1019]) );
  AN2D0 U6069 ( .A1(n[251]), .A2(a[7]), .Z(n[507]) );
  AN2D0 U6070 ( .A1(n[123]), .A2(a[6]), .Z(n[251]) );
  AN2D0 U6071 ( .A1(n[59]), .A2(a[5]), .Z(n[123]) );
  AN2D0 U6072 ( .A1(n[27]), .A2(a[4]), .Z(n[59]) );
  AN2D0 U6073 ( .A1(n[11]), .A2(a[3]), .Z(n[27]) );
  AN2D0 U6074 ( .A1(a[2]), .A2(n[3]), .Z(n[11]) );
  AN2D0 U6075 ( .A1(n[506]), .A2(a[8]), .Z(n[1018]) );
  AN2D0 U6076 ( .A1(n[250]), .A2(a[7]), .Z(n[506]) );
  AN2D0 U6077 ( .A1(n[122]), .A2(a[6]), .Z(n[250]) );
  AN2D0 U6078 ( .A1(n[58]), .A2(a[5]), .Z(n[122]) );
  AN2D0 U6079 ( .A1(n[26]), .A2(a[4]), .Z(n[58]) );
  AN2D0 U6080 ( .A1(n[10]), .A2(a[3]), .Z(n[26]) );
  AN2D0 U6081 ( .A1(a[2]), .A2(b[2]), .Z(n[10]) );
  AN2D0 U6082 ( .A1(n[505]), .A2(a[8]), .Z(n[1017]) );
  AN2D0 U6083 ( .A1(n[249]), .A2(a[7]), .Z(n[505]) );
  AN2D0 U6084 ( .A1(n[121]), .A2(a[6]), .Z(n[249]) );
  AN2D0 U6085 ( .A1(n[57]), .A2(a[5]), .Z(n[121]) );
  AN2D0 U6086 ( .A1(n[25]), .A2(a[4]), .Z(n[57]) );
  AN2D0 U6087 ( .A1(b[3]), .A2(a[3]), .Z(n[25]) );
  AN2D0 U6088 ( .A1(n[504]), .A2(a[8]), .Z(n[1016]) );
  AN2D0 U6089 ( .A1(n[248]), .A2(a[7]), .Z(n[504]) );
  AN2D0 U6090 ( .A1(n[120]), .A2(a[6]), .Z(n[248]) );
  AN2D0 U6091 ( .A1(n[56]), .A2(a[5]), .Z(n[120]) );
  AN2D0 U6092 ( .A1(b[4]), .A2(a[4]), .Z(n[56]) );
  AN2D0 U6093 ( .A1(n[503]), .A2(a[8]), .Z(n[1015]) );
  AN2D0 U6094 ( .A1(n[247]), .A2(a[7]), .Z(n[503]) );
  AN2D0 U6095 ( .A1(n[119]), .A2(a[6]), .Z(n[247]) );
  AN2D0 U6096 ( .A1(b[5]), .A2(a[5]), .Z(n[119]) );
  AN2D0 U6097 ( .A1(n[502]), .A2(a[8]), .Z(n[1014]) );
  AN2D0 U6098 ( .A1(n[246]), .A2(a[7]), .Z(n[502]) );
  AN2D0 U6099 ( .A1(b[6]), .A2(a[6]), .Z(n[246]) );
  AN2D0 U6100 ( .A1(n[501]), .A2(a[8]), .Z(n[1013]) );
  AN2D0 U6101 ( .A1(b[7]), .A2(a[7]), .Z(n[501]) );
  AN2D0 U6102 ( .A1(b[8]), .A2(a[8]), .Z(n[1012]) );
  AN2D0 U6103 ( .A1(b[7]), .A2(n[498]), .Z(n[1009]) );
  AN2D0 U6104 ( .A1(b[6]), .A2(n[243]), .Z(n[498]) );
  AN2D0 U6105 ( .A1(b[5]), .A2(n[116]), .Z(n[243]) );
  AN2D0 U6106 ( .A1(b[4]), .A2(n[53]), .Z(n[116]) );
  AN2D0 U6107 ( .A1(b[3]), .A2(n[22]), .Z(n[53]) );
  AN2D0 U6108 ( .A1(b[2]), .A2(n[7]), .Z(n[22]) );
  AN2D0 U6109 ( .A1(b[7]), .A2(n[495]), .Z(n[1006]) );
  AN2D0 U6110 ( .A1(b[6]), .A2(n[240]), .Z(n[495]) );
  AN2D0 U6111 ( .A1(b[5]), .A2(n[113]), .Z(n[240]) );
  AN2D0 U6112 ( .A1(b[4]), .A2(n[50]), .Z(n[113]) );
  AN2D0 U6113 ( .A1(b[3]), .A2(n[19]), .Z(n[50]) );
  AN2D0 U6114 ( .A1(n[4]), .A2(b[2]), .Z(n[19]) );
  AN2D0 U6115 ( .A1(n[0]), .A2(a[1]), .Z(n[4]) );
  AN2D0 U6116 ( .A1(b[7]), .A2(n[494]), .Z(n[1005]) );
  AN2D0 U6117 ( .A1(b[6]), .A2(n[239]), .Z(n[494]) );
  AN2D0 U6118 ( .A1(b[5]), .A2(n[112]), .Z(n[239]) );
  AN2D0 U6119 ( .A1(b[4]), .A2(n[49]), .Z(n[112]) );
  AN2D0 U6120 ( .A1(b[3]), .A2(n[18]), .Z(n[49]) );
  AN2D0 U6121 ( .A1(n[3]), .A2(b[2]), .Z(n[18]) );
  AN2D0 U6122 ( .A1(a[1]), .A2(b[1]), .Z(n[3]) );
  AN2D0 U6123 ( .A1(b[7]), .A2(n[491]), .Z(n[1002]) );
  AN2D0 U6124 ( .A1(b[6]), .A2(n[236]), .Z(n[491]) );
  AN2D0 U6125 ( .A1(b[5]), .A2(n[109]), .Z(n[236]) );
  AN2D0 U6126 ( .A1(b[4]), .A2(n[46]), .Z(n[109]) );
  AN2D0 U6127 ( .A1(b[3]), .A2(n[15]), .Z(n[46]) );
  AN2D0 U6128 ( .A1(a[2]), .A2(n[7]), .Z(n[15]) );
  AN2D0 U6129 ( .A1(n[0]), .A2(b[1]), .Z(n[7]) );
  AN2D0 U6130 ( .A1(b[0]), .A2(a[0]), .Z(n[0]) );
endmodule


module gen_cla_decomposed ( a, b, s );
  input [10:0] a;
  input [10:0] b;
  output [10:0] s;

  wire   [4081:0] n;

  gen_nonlinear_part NLIN ( .a(a), .b(b), .n(n) );
  gen_linear_part LIN ( .a(a), .b(b), .n({1'b0, 1'b0, n[4079], 1'b0, 1'b0, 
        n[4076:4075], 1'b0, 1'b0, n[4072], 1'b0, 1'b0, n[4069:4067], 1'b0, 
        1'b0, n[4064], 1'b0, 1'b0, n[4061:4060], 1'b0, 1'b0, n[4057], 1'b0, 
        1'b0, n[4054:4051], 1'b0, 1'b0, n[4048], 1'b0, 1'b0, n[4045:4044], 
        1'b0, 1'b0, n[4041], 1'b0, 1'b0, n[4038:4036], 1'b0, 1'b0, n[4033], 
        1'b0, 1'b0, n[4030:4029], 1'b0, 1'b0, n[4026], 1'b0, 1'b0, 
        n[4023:4019], 1'b0, 1'b0, n[4016], 1'b0, 1'b0, n[4013:4012], 1'b0, 
        1'b0, n[4009], 1'b0, 1'b0, n[4006:4004], 1'b0, 1'b0, n[4001], 1'b0, 
        1'b0, n[3998:3997], 1'b0, 1'b0, n[3994], 1'b0, 1'b0, n[3991:3988], 
        1'b0, 1'b0, n[3985], 1'b0, 1'b0, n[3982:3981], 1'b0, 1'b0, n[3978], 
        1'b0, 1'b0, n[3975:3973], 1'b0, 1'b0, n[3970], 1'b0, 1'b0, 
        n[3967:3966], 1'b0, 1'b0, n[3963], 1'b0, 1'b0, n[3960:3955], 1'b0, 
        1'b0, n[3952], 1'b0, 1'b0, n[3949:3948], 1'b0, 1'b0, n[3945], 1'b0, 
        1'b0, n[3942:3940], 1'b0, 1'b0, n[3937], 1'b0, 1'b0, n[3934:3933], 
        1'b0, 1'b0, n[3930], 1'b0, 1'b0, n[3927:3924], 1'b0, 1'b0, n[3921], 
        1'b0, 1'b0, n[3918:3917], 1'b0, 1'b0, n[3914], 1'b0, 1'b0, 
        n[3911:3909], 1'b0, 1'b0, n[3906], 1'b0, 1'b0, n[3903:3902], 1'b0, 
        1'b0, n[3899], 1'b0, 1'b0, n[3896:3892], 1'b0, 1'b0, n[3889], 1'b0, 
        1'b0, n[3886:3885], 1'b0, 1'b0, n[3882], 1'b0, 1'b0, n[3879:3877], 
        1'b0, 1'b0, n[3874], 1'b0, 1'b0, n[3871:3870], 1'b0, 1'b0, n[3867], 
        1'b0, 1'b0, n[3864:3861], 1'b0, 1'b0, n[3858], 1'b0, 1'b0, 
        n[3855:3854], 1'b0, 1'b0, n[3851], 1'b0, 1'b0, n[3848:3846], 1'b0, 
        1'b0, n[3843], 1'b0, 1'b0, n[3840:3839], 1'b0, 1'b0, n[3836], 1'b0, 
        1'b0, n[3833:3827], 1'b0, 1'b0, n[3824], 1'b0, 1'b0, n[3821:3820], 
        1'b0, 1'b0, n[3817], 1'b0, 1'b0, n[3814:3812], 1'b0, 1'b0, n[3809], 
        1'b0, 1'b0, n[3806:3805], 1'b0, 1'b0, n[3802], 1'b0, 1'b0, 
        n[3799:3796], 1'b0, 1'b0, n[3793], 1'b0, 1'b0, n[3790:3789], 1'b0, 
        1'b0, n[3786], 1'b0, 1'b0, n[3783:3781], 1'b0, 1'b0, n[3778], 1'b0, 
        1'b0, n[3775:3774], 1'b0, 1'b0, n[3771], 1'b0, 1'b0, n[3768:3764], 
        1'b0, 1'b0, n[3761], 1'b0, 1'b0, n[3758:3757], 1'b0, 1'b0, n[3754], 
        1'b0, 1'b0, n[3751:3749], 1'b0, 1'b0, n[3746], 1'b0, 1'b0, 
        n[3743:3742], 1'b0, 1'b0, n[3739], 1'b0, 1'b0, n[3736:3733], 1'b0, 
        1'b0, n[3730], 1'b0, 1'b0, n[3727:3726], 1'b0, 1'b0, n[3723], 1'b0, 
        1'b0, n[3720:3718], 1'b0, 1'b0, n[3715], 1'b0, 1'b0, n[3712:3711], 
        1'b0, 1'b0, n[3708], 1'b0, 1'b0, n[3705:3700], 1'b0, 1'b0, n[3697], 
        1'b0, 1'b0, n[3694:3693], 1'b0, 1'b0, n[3690], 1'b0, 1'b0, 
        n[3687:3685], 1'b0, 1'b0, n[3682], 1'b0, 1'b0, n[3679:3678], 1'b0, 
        1'b0, n[3675], 1'b0, 1'b0, n[3672:3669], 1'b0, 1'b0, n[3666], 1'b0, 
        1'b0, n[3663:3662], 1'b0, 1'b0, n[3659], 1'b0, 1'b0, n[3656:3654], 
        1'b0, 1'b0, n[3651], 1'b0, 1'b0, n[3648:3647], 1'b0, 1'b0, n[3644], 
        1'b0, 1'b0, n[3641:3637], 1'b0, 1'b0, n[3634], 1'b0, 1'b0, 
        n[3631:3630], 1'b0, 1'b0, n[3627], 1'b0, 1'b0, n[3624:3622], 1'b0, 
        1'b0, n[3619], 1'b0, 1'b0, n[3616:3615], 1'b0, 1'b0, n[3612], 1'b0, 
        1'b0, n[3609:3606], 1'b0, 1'b0, n[3603], 1'b0, 1'b0, n[3600:3599], 
        1'b0, 1'b0, n[3596], 1'b0, 1'b0, n[3593:3591], 1'b0, 1'b0, n[3588], 
        1'b0, 1'b0, n[3585:3584], 1'b0, 1'b0, n[3581], 1'b0, 1'b0, 
        n[3578:3571], 1'b0, 1'b0, n[3568], 1'b0, 1'b0, n[3565:3564], 1'b0, 
        1'b0, n[3561], 1'b0, 1'b0, n[3558:3556], 1'b0, 1'b0, n[3553], 1'b0, 
        1'b0, n[3550:3549], 1'b0, 1'b0, n[3546], 1'b0, 1'b0, n[3543:3540], 
        1'b0, 1'b0, n[3537], 1'b0, 1'b0, n[3534:3533], 1'b0, 1'b0, n[3530], 
        1'b0, 1'b0, n[3527:3525], 1'b0, 1'b0, n[3522], 1'b0, 1'b0, 
        n[3519:3518], 1'b0, 1'b0, n[3515], 1'b0, 1'b0, n[3512:3508], 1'b0, 
        1'b0, n[3505], 1'b0, 1'b0, n[3502:3501], 1'b0, 1'b0, n[3498], 1'b0, 
        1'b0, n[3495:3493], 1'b0, 1'b0, n[3490], 1'b0, 1'b0, n[3487:3486], 
        1'b0, 1'b0, n[3483], 1'b0, 1'b0, n[3480:3477], 1'b0, 1'b0, n[3474], 
        1'b0, 1'b0, n[3471:3470], 1'b0, 1'b0, n[3467], 1'b0, 1'b0, 
        n[3464:3462], 1'b0, 1'b0, n[3459], 1'b0, 1'b0, n[3456:3455], 1'b0, 
        1'b0, n[3452], 1'b0, 1'b0, n[3449:3444], 1'b0, 1'b0, n[3441], 1'b0, 
        1'b0, n[3438:3437], 1'b0, 1'b0, n[3434], 1'b0, 1'b0, n[3431:3429], 
        1'b0, 1'b0, n[3426], 1'b0, 1'b0, n[3423:3422], 1'b0, 1'b0, n[3419], 
        1'b0, 1'b0, n[3416:3413], 1'b0, 1'b0, n[3410], 1'b0, 1'b0, 
        n[3407:3406], 1'b0, 1'b0, n[3403], 1'b0, 1'b0, n[3400:3398], 1'b0, 
        1'b0, n[3395], 1'b0, 1'b0, n[3392:3391], 1'b0, 1'b0, n[3388], 1'b0, 
        1'b0, n[3385:3381], 1'b0, 1'b0, n[3378], 1'b0, 1'b0, n[3375:3374], 
        1'b0, 1'b0, n[3371], 1'b0, 1'b0, n[3368:3366], 1'b0, 1'b0, n[3363], 
        1'b0, 1'b0, n[3360:3359], 1'b0, 1'b0, n[3356], 1'b0, 1'b0, 
        n[3353:3350], 1'b0, 1'b0, n[3347], 1'b0, 1'b0, n[3344:3343], 1'b0, 
        1'b0, n[3340], 1'b0, 1'b0, n[3337:3335], 1'b0, 1'b0, n[3332], 1'b0, 
        1'b0, n[3329:3328], 1'b0, 1'b0, n[3325], 1'b0, 1'b0, n[3322:3316], 
        1'b0, 1'b0, n[3313], 1'b0, 1'b0, n[3310:3309], 1'b0, 1'b0, n[3306], 
        1'b0, 1'b0, n[3303:3301], 1'b0, 1'b0, n[3298], 1'b0, 1'b0, 
        n[3295:3294], 1'b0, 1'b0, n[3291], 1'b0, 1'b0, n[3288:3285], 1'b0, 
        1'b0, n[3282], 1'b0, 1'b0, n[3279:3278], 1'b0, 1'b0, n[3275], 1'b0, 
        1'b0, n[3272:3270], 1'b0, 1'b0, n[3267], 1'b0, 1'b0, n[3264:3263], 
        1'b0, 1'b0, n[3260], 1'b0, 1'b0, n[3257:3253], 1'b0, 1'b0, n[3250], 
        1'b0, 1'b0, n[3247:3246], 1'b0, 1'b0, n[3243], 1'b0, 1'b0, 
        n[3240:3238], 1'b0, 1'b0, n[3235], 1'b0, 1'b0, n[3232:3231], 1'b0, 
        1'b0, n[3228], 1'b0, 1'b0, n[3225:3222], 1'b0, 1'b0, n[3219], 1'b0, 
        1'b0, n[3216:3215], 1'b0, 1'b0, n[3212], 1'b0, 1'b0, n[3209:3207], 
        1'b0, 1'b0, n[3204], 1'b0, 1'b0, n[3201:3200], 1'b0, 1'b0, n[3197], 
        1'b0, 1'b0, n[3194:3189], 1'b0, 1'b0, n[3186], 1'b0, 1'b0, 
        n[3183:3182], 1'b0, 1'b0, n[3179], 1'b0, 1'b0, n[3176:3174], 1'b0, 
        1'b0, n[3171], 1'b0, 1'b0, n[3168:3167], 1'b0, 1'b0, n[3164], 1'b0, 
        1'b0, n[3161:3158], 1'b0, 1'b0, n[3155], 1'b0, 1'b0, n[3152:3151], 
        1'b0, 1'b0, n[3148], 1'b0, 1'b0, n[3145:3143], 1'b0, 1'b0, n[3140], 
        1'b0, 1'b0, n[3137:3136], 1'b0, 1'b0, n[3133], 1'b0, 1'b0, 
        n[3130:3126], 1'b0, 1'b0, n[3123], 1'b0, 1'b0, n[3120:3119], 1'b0, 
        1'b0, n[3116], 1'b0, 1'b0, n[3113:3111], 1'b0, 1'b0, n[3108], 1'b0, 
        1'b0, n[3105:3104], 1'b0, 1'b0, n[3101], 1'b0, 1'b0, n[3098:3095], 
        1'b0, 1'b0, n[3092], 1'b0, 1'b0, n[3089:3088], 1'b0, 1'b0, n[3085], 
        1'b0, 1'b0, n[3082:3080], 1'b0, 1'b0, n[3077], 1'b0, 1'b0, 
        n[3074:3073], 1'b0, 1'b0, n[3070], 1'b0, 1'b0, n[3067:3059], 1'b0, 
        1'b0, n[3056], 1'b0, 1'b0, n[3053:3052], 1'b0, 1'b0, n[3049], 1'b0, 
        1'b0, n[3046:3044], 1'b0, 1'b0, n[3041], 1'b0, 1'b0, n[3038:3037], 
        1'b0, 1'b0, n[3034], 1'b0, 1'b0, n[3031:3028], 1'b0, 1'b0, n[3025], 
        1'b0, 1'b0, n[3022:3021], 1'b0, 1'b0, n[3018], 1'b0, 1'b0, 
        n[3015:3013], 1'b0, 1'b0, n[3010], 1'b0, 1'b0, n[3007:3006], 1'b0, 
        1'b0, n[3003], 1'b0, 1'b0, n[3000:2996], 1'b0, 1'b0, n[2993], 1'b0, 
        1'b0, n[2990:2989], 1'b0, 1'b0, n[2986], 1'b0, 1'b0, n[2983:2981], 
        1'b0, 1'b0, n[2978], 1'b0, 1'b0, n[2975:2974], 1'b0, 1'b0, n[2971], 
        1'b0, 1'b0, n[2968:2965], 1'b0, 1'b0, n[2962], 1'b0, 1'b0, 
        n[2959:2958], 1'b0, 1'b0, n[2955], 1'b0, 1'b0, n[2952:2950], 1'b0, 
        1'b0, n[2947], 1'b0, 1'b0, n[2944:2943], 1'b0, 1'b0, n[2940], 1'b0, 
        1'b0, n[2937:2932], 1'b0, 1'b0, n[2929], 1'b0, 1'b0, n[2926:2925], 
        1'b0, 1'b0, n[2922], 1'b0, 1'b0, n[2919:2917], 1'b0, 1'b0, n[2914], 
        1'b0, 1'b0, n[2911:2910], 1'b0, 1'b0, n[2907], 1'b0, 1'b0, 
        n[2904:2901], 1'b0, 1'b0, n[2898], 1'b0, 1'b0, n[2895:2894], 1'b0, 
        1'b0, n[2891], 1'b0, 1'b0, n[2888:2886], 1'b0, 1'b0, n[2883], 1'b0, 
        1'b0, n[2880:2879], 1'b0, 1'b0, n[2876], 1'b0, 1'b0, n[2873:2869], 
        1'b0, 1'b0, n[2866], 1'b0, 1'b0, n[2863:2862], 1'b0, 1'b0, n[2859], 
        1'b0, 1'b0, n[2856:2854], 1'b0, 1'b0, n[2851], 1'b0, 1'b0, 
        n[2848:2847], 1'b0, 1'b0, n[2844], 1'b0, 1'b0, n[2841:2838], 1'b0, 
        1'b0, n[2835], 1'b0, 1'b0, n[2832:2831], 1'b0, 1'b0, n[2828], 1'b0, 
        1'b0, n[2825:2823], 1'b0, 1'b0, n[2820], 1'b0, 1'b0, n[2817:2816], 
        1'b0, 1'b0, n[2813], 1'b0, 1'b0, n[2810:2804], 1'b0, 1'b0, n[2801], 
        1'b0, 1'b0, n[2798:2797], 1'b0, 1'b0, n[2794], 1'b0, 1'b0, 
        n[2791:2789], 1'b0, 1'b0, n[2786], 1'b0, 1'b0, n[2783:2782], 1'b0, 
        1'b0, n[2779], 1'b0, 1'b0, n[2776:2773], 1'b0, 1'b0, n[2770], 1'b0, 
        1'b0, n[2767:2766], 1'b0, 1'b0, n[2763], 1'b0, 1'b0, n[2760:2758], 
        1'b0, 1'b0, n[2755], 1'b0, 1'b0, n[2752:2751], 1'b0, 1'b0, n[2748], 
        1'b0, 1'b0, n[2745:2741], 1'b0, 1'b0, n[2738], 1'b0, 1'b0, 
        n[2735:2734], 1'b0, 1'b0, n[2731], 1'b0, 1'b0, n[2728:2726], 1'b0, 
        1'b0, n[2723], 1'b0, 1'b0, n[2720:2719], 1'b0, 1'b0, n[2716], 1'b0, 
        1'b0, n[2713:2710], 1'b0, 1'b0, n[2707], 1'b0, 1'b0, n[2704:2703], 
        1'b0, 1'b0, n[2700], 1'b0, 1'b0, n[2697:2695], 1'b0, 1'b0, n[2692], 
        1'b0, 1'b0, n[2689:2688], 1'b0, 1'b0, n[2685], 1'b0, 1'b0, 
        n[2682:2677], 1'b0, 1'b0, n[2674], 1'b0, 1'b0, n[2671:2670], 1'b0, 
        1'b0, n[2667], 1'b0, 1'b0, n[2664:2662], 1'b0, 1'b0, n[2659], 1'b0, 
        1'b0, n[2656:2655], 1'b0, 1'b0, n[2652], 1'b0, 1'b0, n[2649:2646], 
        1'b0, 1'b0, n[2643], 1'b0, 1'b0, n[2640:2639], 1'b0, 1'b0, n[2636], 
        1'b0, 1'b0, n[2633:2631], 1'b0, 1'b0, n[2628], 1'b0, 1'b0, 
        n[2625:2624], 1'b0, 1'b0, n[2621], 1'b0, 1'b0, n[2618:2614], 1'b0, 
        1'b0, n[2611], 1'b0, 1'b0, n[2608:2607], 1'b0, 1'b0, n[2604], 1'b0, 
        1'b0, n[2601:2599], 1'b0, 1'b0, n[2596], 1'b0, 1'b0, n[2593:2592], 
        1'b0, 1'b0, n[2589], 1'b0, 1'b0, n[2586:2583], 1'b0, 1'b0, n[2580], 
        1'b0, 1'b0, n[2577:2576], 1'b0, 1'b0, n[2573], 1'b0, 1'b0, 
        n[2570:2568], 1'b0, 1'b0, n[2565], 1'b0, 1'b0, n[2562:2561], 1'b0, 
        1'b0, n[2558], 1'b0, 1'b0, n[2555:2548], 1'b0, 1'b0, n[2545], 1'b0, 
        1'b0, n[2542:2541], 1'b0, 1'b0, n[2538], 1'b0, 1'b0, n[2535:2533], 
        1'b0, 1'b0, n[2530], 1'b0, 1'b0, n[2527:2526], 1'b0, 1'b0, n[2523], 
        1'b0, 1'b0, n[2520:2517], 1'b0, 1'b0, n[2514], 1'b0, 1'b0, 
        n[2511:2510], 1'b0, 1'b0, n[2507], 1'b0, 1'b0, n[2504:2502], 1'b0, 
        1'b0, n[2499], 1'b0, 1'b0, n[2496:2495], 1'b0, 1'b0, n[2492], 1'b0, 
        1'b0, n[2489:2485], 1'b0, 1'b0, n[2482], 1'b0, 1'b0, n[2479:2478], 
        1'b0, 1'b0, n[2475], 1'b0, 1'b0, n[2472:2470], 1'b0, 1'b0, n[2467], 
        1'b0, 1'b0, n[2464:2463], 1'b0, 1'b0, n[2460], 1'b0, 1'b0, 
        n[2457:2454], 1'b0, 1'b0, n[2451], 1'b0, 1'b0, n[2448:2447], 1'b0, 
        1'b0, n[2444], 1'b0, 1'b0, n[2441:2439], 1'b0, 1'b0, n[2436], 1'b0, 
        1'b0, n[2433:2432], 1'b0, 1'b0, n[2429], 1'b0, 1'b0, n[2426:2421], 
        1'b0, 1'b0, n[2418], 1'b0, 1'b0, n[2415:2414], 1'b0, 1'b0, n[2411], 
        1'b0, 1'b0, n[2408:2406], 1'b0, 1'b0, n[2403], 1'b0, 1'b0, 
        n[2400:2399], 1'b0, 1'b0, n[2396], 1'b0, 1'b0, n[2393:2390], 1'b0, 
        1'b0, n[2387], 1'b0, 1'b0, n[2384:2383], 1'b0, 1'b0, n[2380], 1'b0, 
        1'b0, n[2377:2375], 1'b0, 1'b0, n[2372], 1'b0, 1'b0, n[2369:2368], 
        1'b0, 1'b0, n[2365], 1'b0, 1'b0, n[2362:2358], 1'b0, 1'b0, n[2355], 
        1'b0, 1'b0, n[2352:2351], 1'b0, 1'b0, n[2348], 1'b0, 1'b0, 
        n[2345:2343], 1'b0, 1'b0, n[2340], 1'b0, 1'b0, n[2337:2336], 1'b0, 
        1'b0, n[2333], 1'b0, 1'b0, n[2330:2327], 1'b0, 1'b0, n[2324], 1'b0, 
        1'b0, n[2321:2320], 1'b0, 1'b0, n[2317], 1'b0, 1'b0, n[2314:2312], 
        1'b0, 1'b0, n[2309], 1'b0, 1'b0, n[2306:2305], 1'b0, 1'b0, n[2302], 
        1'b0, 1'b0, n[2299:2293], 1'b0, 1'b0, n[2290], 1'b0, 1'b0, 
        n[2287:2286], 1'b0, 1'b0, n[2283], 1'b0, 1'b0, n[2280:2278], 1'b0, 
        1'b0, n[2275], 1'b0, 1'b0, n[2272:2271], 1'b0, 1'b0, n[2268], 1'b0, 
        1'b0, n[2265:2262], 1'b0, 1'b0, n[2259], 1'b0, 1'b0, n[2256:2255], 
        1'b0, 1'b0, n[2252], 1'b0, 1'b0, n[2249:2247], 1'b0, 1'b0, n[2244], 
        1'b0, 1'b0, n[2241:2240], 1'b0, 1'b0, n[2237], 1'b0, 1'b0, 
        n[2234:2230], 1'b0, 1'b0, n[2227], 1'b0, 1'b0, n[2224:2223], 1'b0, 
        1'b0, n[2220], 1'b0, 1'b0, n[2217:2215], 1'b0, 1'b0, n[2212], 1'b0, 
        1'b0, n[2209:2208], 1'b0, 1'b0, n[2205], 1'b0, 1'b0, n[2202:2199], 
        1'b0, 1'b0, n[2196], 1'b0, 1'b0, n[2193:2192], 1'b0, 1'b0, n[2189], 
        1'b0, 1'b0, n[2186:2184], 1'b0, 1'b0, n[2181], 1'b0, 1'b0, 
        n[2178:2177], 1'b0, 1'b0, n[2174], 1'b0, 1'b0, n[2171:2166], 1'b0, 
        1'b0, n[2163], 1'b0, 1'b0, n[2160:2159], 1'b0, 1'b0, n[2156], 1'b0, 
        1'b0, n[2153:2151], 1'b0, 1'b0, n[2148], 1'b0, 1'b0, n[2145:2144], 
        1'b0, 1'b0, n[2141], 1'b0, 1'b0, n[2138:2135], 1'b0, 1'b0, n[2132], 
        1'b0, 1'b0, n[2129:2128], 1'b0, 1'b0, n[2125], 1'b0, 1'b0, 
        n[2122:2120], 1'b0, 1'b0, n[2117], 1'b0, 1'b0, n[2114:2113], 1'b0, 
        1'b0, n[2110], 1'b0, 1'b0, n[2107:2103], 1'b0, 1'b0, n[2100], 1'b0, 
        1'b0, n[2097:2096], 1'b0, 1'b0, n[2093], 1'b0, 1'b0, n[2090:2088], 
        1'b0, 1'b0, n[2085], 1'b0, 1'b0, n[2082:2081], 1'b0, 1'b0, n[2078], 
        1'b0, 1'b0, n[2075:2072], 1'b0, 1'b0, n[2069], 1'b0, 1'b0, 
        n[2066:2065], 1'b0, 1'b0, n[2062], 1'b0, 1'b0, n[2059:2057], 1'b0, 
        1'b0, n[2054], 1'b0, 1'b0, n[2051:2050], 1'b0, 1'b0, n[2047], 1'b0, 
        1'b0, n[2044:2035], 1'b0, 1'b0, n[2032], 1'b0, 1'b0, n[2029:2028], 
        1'b0, 1'b0, n[2025], 1'b0, 1'b0, n[2022:2020], 1'b0, 1'b0, n[2017], 
        1'b0, 1'b0, n[2014:2013], 1'b0, 1'b0, n[2010], 1'b0, 1'b0, 
        n[2007:2004], 1'b0, 1'b0, n[2001], 1'b0, 1'b0, n[1998:1997], 1'b0, 
        1'b0, n[1994], 1'b0, 1'b0, n[1991:1989], 1'b0, 1'b0, n[1986], 1'b0, 
        1'b0, n[1983:1982], 1'b0, 1'b0, n[1979], 1'b0, 1'b0, n[1976:1972], 
        1'b0, 1'b0, n[1969], 1'b0, 1'b0, n[1966:1965], 1'b0, 1'b0, n[1962], 
        1'b0, 1'b0, n[1959:1957], 1'b0, 1'b0, n[1954], 1'b0, 1'b0, 
        n[1951:1950], 1'b0, 1'b0, n[1947], 1'b0, 1'b0, n[1944:1941], 1'b0, 
        1'b0, n[1938], 1'b0, 1'b0, n[1935:1934], 1'b0, 1'b0, n[1931], 1'b0, 
        1'b0, n[1928:1926], 1'b0, 1'b0, n[1923], 1'b0, 1'b0, n[1920:1919], 
        1'b0, 1'b0, n[1916], 1'b0, 1'b0, n[1913:1908], 1'b0, 1'b0, n[1905], 
        1'b0, 1'b0, n[1902:1901], 1'b0, 1'b0, n[1898], 1'b0, 1'b0, 
        n[1895:1893], 1'b0, 1'b0, n[1890], 1'b0, 1'b0, n[1887:1886], 1'b0, 
        1'b0, n[1883], 1'b0, 1'b0, n[1880:1877], 1'b0, 1'b0, n[1874], 1'b0, 
        1'b0, n[1871:1870], 1'b0, 1'b0, n[1867], 1'b0, 1'b0, n[1864:1862], 
        1'b0, 1'b0, n[1859], 1'b0, 1'b0, n[1856:1855], 1'b0, 1'b0, n[1852], 
        1'b0, 1'b0, n[1849:1845], 1'b0, 1'b0, n[1842], 1'b0, 1'b0, 
        n[1839:1838], 1'b0, 1'b0, n[1835], 1'b0, 1'b0, n[1832:1830], 1'b0, 
        1'b0, n[1827], 1'b0, 1'b0, n[1824:1823], 1'b0, 1'b0, n[1820], 1'b0, 
        1'b0, n[1817:1814], 1'b0, 1'b0, n[1811], 1'b0, 1'b0, n[1808:1807], 
        1'b0, 1'b0, n[1804], 1'b0, 1'b0, n[1801:1799], 1'b0, 1'b0, n[1796], 
        1'b0, 1'b0, n[1793:1792], 1'b0, 1'b0, n[1789], 1'b0, 1'b0, 
        n[1786:1780], 1'b0, 1'b0, n[1777], 1'b0, 1'b0, n[1774:1773], 1'b0, 
        1'b0, n[1770], 1'b0, 1'b0, n[1767:1765], 1'b0, 1'b0, n[1762], 1'b0, 
        1'b0, n[1759:1758], 1'b0, 1'b0, n[1755], 1'b0, 1'b0, n[1752:1749], 
        1'b0, 1'b0, n[1746], 1'b0, 1'b0, n[1743:1742], 1'b0, 1'b0, n[1739], 
        1'b0, 1'b0, n[1736:1734], 1'b0, 1'b0, n[1731], 1'b0, 1'b0, 
        n[1728:1727], 1'b0, 1'b0, n[1724], 1'b0, 1'b0, n[1721:1717], 1'b0, 
        1'b0, n[1714], 1'b0, 1'b0, n[1711:1710], 1'b0, 1'b0, n[1707], 1'b0, 
        1'b0, n[1704:1702], 1'b0, 1'b0, n[1699], 1'b0, 1'b0, n[1696:1695], 
        1'b0, 1'b0, n[1692], 1'b0, 1'b0, n[1689:1686], 1'b0, 1'b0, n[1683], 
        1'b0, 1'b0, n[1680:1679], 1'b0, 1'b0, n[1676], 1'b0, 1'b0, 
        n[1673:1671], 1'b0, 1'b0, n[1668], 1'b0, 1'b0, n[1665:1664], 1'b0, 
        1'b0, n[1661], 1'b0, 1'b0, n[1658:1653], 1'b0, 1'b0, n[1650], 1'b0, 
        1'b0, n[1647:1646], 1'b0, 1'b0, n[1643], 1'b0, 1'b0, n[1640:1638], 
        1'b0, 1'b0, n[1635], 1'b0, 1'b0, n[1632:1631], 1'b0, 1'b0, n[1628], 
        1'b0, 1'b0, n[1625:1622], 1'b0, 1'b0, n[1619], 1'b0, 1'b0, 
        n[1616:1615], 1'b0, 1'b0, n[1612], 1'b0, 1'b0, n[1609:1607], 1'b0, 
        1'b0, n[1604], 1'b0, 1'b0, n[1601:1600], 1'b0, 1'b0, n[1597], 1'b0, 
        1'b0, n[1594:1590], 1'b0, 1'b0, n[1587], 1'b0, 1'b0, n[1584:1583], 
        1'b0, 1'b0, n[1580], 1'b0, 1'b0, n[1577:1575], 1'b0, 1'b0, n[1572], 
        1'b0, 1'b0, n[1569:1568], 1'b0, 1'b0, n[1565], 1'b0, 1'b0, 
        n[1562:1559], 1'b0, 1'b0, n[1556], 1'b0, 1'b0, n[1553:1552], 1'b0, 
        1'b0, n[1549], 1'b0, 1'b0, n[1546:1544], 1'b0, 1'b0, n[1541], 1'b0, 
        1'b0, n[1538:1537], 1'b0, 1'b0, n[1534], 1'b0, 1'b0, n[1531:1524], 
        1'b0, 1'b0, n[1521], 1'b0, 1'b0, n[1518:1517], 1'b0, 1'b0, n[1514], 
        1'b0, 1'b0, n[1511:1509], 1'b0, 1'b0, n[1506], 1'b0, 1'b0, 
        n[1503:1502], 1'b0, 1'b0, n[1499], 1'b0, 1'b0, n[1496:1493], 1'b0, 
        1'b0, n[1490], 1'b0, 1'b0, n[1487:1486], 1'b0, 1'b0, n[1483], 1'b0, 
        1'b0, n[1480:1478], 1'b0, 1'b0, n[1475], 1'b0, 1'b0, n[1472:1471], 
        1'b0, 1'b0, n[1468], 1'b0, 1'b0, n[1465:1461], 1'b0, 1'b0, n[1458], 
        1'b0, 1'b0, n[1455:1454], 1'b0, 1'b0, n[1451], 1'b0, 1'b0, 
        n[1448:1446], 1'b0, 1'b0, n[1443], 1'b0, 1'b0, n[1440:1439], 1'b0, 
        1'b0, n[1436], 1'b0, 1'b0, n[1433:1430], 1'b0, 1'b0, n[1427], 1'b0, 
        1'b0, n[1424:1423], 1'b0, 1'b0, n[1420], 1'b0, 1'b0, n[1417:1415], 
        1'b0, 1'b0, n[1412], 1'b0, 1'b0, n[1409:1408], 1'b0, 1'b0, n[1405], 
        1'b0, 1'b0, n[1402:1397], 1'b0, 1'b0, n[1394], 1'b0, 1'b0, 
        n[1391:1390], 1'b0, 1'b0, n[1387], 1'b0, 1'b0, n[1384:1382], 1'b0, 
        1'b0, n[1379], 1'b0, 1'b0, n[1376:1375], 1'b0, 1'b0, n[1372], 1'b0, 
        1'b0, n[1369:1366], 1'b0, 1'b0, n[1363], 1'b0, 1'b0, n[1360:1359], 
        1'b0, 1'b0, n[1356], 1'b0, 1'b0, n[1353:1351], 1'b0, 1'b0, n[1348], 
        1'b0, 1'b0, n[1345:1344], 1'b0, 1'b0, n[1341], 1'b0, 1'b0, 
        n[1338:1334], 1'b0, 1'b0, n[1331], 1'b0, 1'b0, n[1328:1327], 1'b0, 
        1'b0, n[1324], 1'b0, 1'b0, n[1321:1319], 1'b0, 1'b0, n[1316], 1'b0, 
        1'b0, n[1313:1312], 1'b0, 1'b0, n[1309], 1'b0, 1'b0, n[1306:1303], 
        1'b0, 1'b0, n[1300], 1'b0, 1'b0, n[1297:1296], 1'b0, 1'b0, n[1293], 
        1'b0, 1'b0, n[1290:1288], 1'b0, 1'b0, n[1285], 1'b0, 1'b0, 
        n[1282:1281], 1'b0, 1'b0, n[1278], 1'b0, 1'b0, n[1275:1269], 1'b0, 
        1'b0, n[1266], 1'b0, 1'b0, n[1263:1262], 1'b0, 1'b0, n[1259], 1'b0, 
        1'b0, n[1256:1254], 1'b0, 1'b0, n[1251], 1'b0, 1'b0, n[1248:1247], 
        1'b0, 1'b0, n[1244], 1'b0, 1'b0, n[1241:1238], 1'b0, 1'b0, n[1235], 
        1'b0, 1'b0, n[1232:1231], 1'b0, 1'b0, n[1228], 1'b0, 1'b0, 
        n[1225:1223], 1'b0, 1'b0, n[1220], 1'b0, 1'b0, n[1217:1216], 1'b0, 
        1'b0, n[1213], 1'b0, 1'b0, n[1210:1206], 1'b0, 1'b0, n[1203], 1'b0, 
        1'b0, n[1200:1199], 1'b0, 1'b0, n[1196], 1'b0, 1'b0, n[1193:1191], 
        1'b0, 1'b0, n[1188], 1'b0, 1'b0, n[1185:1184], 1'b0, 1'b0, n[1181], 
        1'b0, 1'b0, n[1178:1175], 1'b0, 1'b0, n[1172], 1'b0, 1'b0, 
        n[1169:1168], 1'b0, 1'b0, n[1165], 1'b0, 1'b0, n[1162:1160], 1'b0, 
        1'b0, n[1157], 1'b0, 1'b0, n[1154:1153], 1'b0, 1'b0, n[1150], 1'b0, 
        1'b0, n[1147:1142], 1'b0, 1'b0, n[1139], 1'b0, 1'b0, n[1136:1135], 
        1'b0, 1'b0, n[1132], 1'b0, 1'b0, n[1129:1127], 1'b0, 1'b0, n[1124], 
        1'b0, 1'b0, n[1121:1120], 1'b0, 1'b0, n[1117], 1'b0, 1'b0, 
        n[1114:1111], 1'b0, 1'b0, n[1108], 1'b0, 1'b0, n[1105:1104], 1'b0, 
        1'b0, n[1101], 1'b0, 1'b0, n[1098:1096], 1'b0, 1'b0, n[1093], 1'b0, 
        1'b0, n[1090:1089], 1'b0, 1'b0, n[1086], 1'b0, 1'b0, n[1083:1079], 
        1'b0, 1'b0, n[1076], 1'b0, 1'b0, n[1073:1072], 1'b0, 1'b0, n[1069], 
        1'b0, 1'b0, n[1066:1064], 1'b0, 1'b0, n[1061], 1'b0, 1'b0, 
        n[1058:1057], 1'b0, 1'b0, n[1054], 1'b0, 1'b0, n[1051:1048], 1'b0, 
        1'b0, n[1045], 1'b0, 1'b0, n[1042:1041], 1'b0, 1'b0, n[1038], 1'b0, 
        1'b0, n[1035:1033], 1'b0, 1'b0, n[1030], 1'b0, 1'b0, n[1027:1026], 
        1'b0, 1'b0, n[1023], 1'b0, 1'b0, n[1020:1012], 1'b0, 1'b0, n[1009], 
        1'b0, 1'b0, n[1006:1005], 1'b0, 1'b0, n[1002], 1'b0, 1'b0, n[999:997], 
        1'b0, 1'b0, n[994], 1'b0, 1'b0, n[991:990], 1'b0, 1'b0, n[987], 1'b0, 
        1'b0, n[984:981], 1'b0, 1'b0, n[978], 1'b0, 1'b0, n[975:974], 1'b0, 
        1'b0, n[971], 1'b0, 1'b0, n[968:966], 1'b0, 1'b0, n[963], 1'b0, 1'b0, 
        n[960:959], 1'b0, 1'b0, n[956], 1'b0, 1'b0, n[953:949], 1'b0, 1'b0, 
        n[946], 1'b0, 1'b0, n[943:942], 1'b0, 1'b0, n[939], 1'b0, 1'b0, 
        n[936:934], 1'b0, 1'b0, n[931], 1'b0, 1'b0, n[928:927], 1'b0, 1'b0, 
        n[924], 1'b0, 1'b0, n[921:918], 1'b0, 1'b0, n[915], 1'b0, 1'b0, 
        n[912:911], 1'b0, 1'b0, n[908], 1'b0, 1'b0, n[905:903], 1'b0, 1'b0, 
        n[900], 1'b0, 1'b0, n[897:896], 1'b0, 1'b0, n[893], 1'b0, 1'b0, 
        n[890:885], 1'b0, 1'b0, n[882], 1'b0, 1'b0, n[879:878], 1'b0, 1'b0, 
        n[875], 1'b0, 1'b0, n[872:870], 1'b0, 1'b0, n[867], 1'b0, 1'b0, 
        n[864:863], 1'b0, 1'b0, n[860], 1'b0, 1'b0, n[857:854], 1'b0, 1'b0, 
        n[851], 1'b0, 1'b0, n[848:847], 1'b0, 1'b0, n[844], 1'b0, 1'b0, 
        n[841:839], 1'b0, 1'b0, n[836], 1'b0, 1'b0, n[833:832], 1'b0, 1'b0, 
        n[829], 1'b0, 1'b0, n[826:822], 1'b0, 1'b0, n[819], 1'b0, 1'b0, 
        n[816:815], 1'b0, 1'b0, n[812], 1'b0, 1'b0, n[809:807], 1'b0, 1'b0, 
        n[804], 1'b0, 1'b0, n[801:800], 1'b0, 1'b0, n[797], 1'b0, 1'b0, 
        n[794:791], 1'b0, 1'b0, n[788], 1'b0, 1'b0, n[785:784], 1'b0, 1'b0, 
        n[781], 1'b0, 1'b0, n[778:776], 1'b0, 1'b0, n[773], 1'b0, 1'b0, 
        n[770:769], 1'b0, 1'b0, n[766], 1'b0, 1'b0, n[763:757], 1'b0, 1'b0, 
        n[754], 1'b0, 1'b0, n[751:750], 1'b0, 1'b0, n[747], 1'b0, 1'b0, 
        n[744:742], 1'b0, 1'b0, n[739], 1'b0, 1'b0, n[736:735], 1'b0, 1'b0, 
        n[732], 1'b0, 1'b0, n[729:726], 1'b0, 1'b0, n[723], 1'b0, 1'b0, 
        n[720:719], 1'b0, 1'b0, n[716], 1'b0, 1'b0, n[713:711], 1'b0, 1'b0, 
        n[708], 1'b0, 1'b0, n[705:704], 1'b0, 1'b0, n[701], 1'b0, 1'b0, 
        n[698:694], 1'b0, 1'b0, n[691], 1'b0, 1'b0, n[688:687], 1'b0, 1'b0, 
        n[684], 1'b0, 1'b0, n[681:679], 1'b0, 1'b0, n[676], 1'b0, 1'b0, 
        n[673:672], 1'b0, 1'b0, n[669], 1'b0, 1'b0, n[666:663], 1'b0, 1'b0, 
        n[660], 1'b0, 1'b0, n[657:656], 1'b0, 1'b0, n[653], 1'b0, 1'b0, 
        n[650:648], 1'b0, 1'b0, n[645], 1'b0, 1'b0, n[642:641], 1'b0, 1'b0, 
        n[638], 1'b0, 1'b0, n[635:630], 1'b0, 1'b0, n[627], 1'b0, 1'b0, 
        n[624:623], 1'b0, 1'b0, n[620], 1'b0, 1'b0, n[617:615], 1'b0, 1'b0, 
        n[612], 1'b0, 1'b0, n[609:608], 1'b0, 1'b0, n[605], 1'b0, 1'b0, 
        n[602:599], 1'b0, 1'b0, n[596], 1'b0, 1'b0, n[593:592], 1'b0, 1'b0, 
        n[589], 1'b0, 1'b0, n[586:584], 1'b0, 1'b0, n[581], 1'b0, 1'b0, 
        n[578:577], 1'b0, 1'b0, n[574], 1'b0, 1'b0, n[571:567], 1'b0, 1'b0, 
        n[564], 1'b0, 1'b0, n[561:560], 1'b0, 1'b0, n[557], 1'b0, 1'b0, 
        n[554:552], 1'b0, 1'b0, n[549], 1'b0, 1'b0, n[546:545], 1'b0, 1'b0, 
        n[542], 1'b0, 1'b0, n[539:536], 1'b0, 1'b0, n[533], 1'b0, 1'b0, 
        n[530:529], 1'b0, 1'b0, n[526], 1'b0, 1'b0, n[523:521], 1'b0, 1'b0, 
        n[518], 1'b0, 1'b0, n[515:514], 1'b0, 1'b0, n[511], 1'b0, 1'b0, 
        n[508:501], 1'b0, 1'b0, n[498], 1'b0, 1'b0, n[495:494], 1'b0, 1'b0, 
        n[491], 1'b0, 1'b0, n[488:486], 1'b0, 1'b0, n[483], 1'b0, 1'b0, 
        n[480:479], 1'b0, 1'b0, n[476], 1'b0, 1'b0, n[473:470], 1'b0, 1'b0, 
        n[467], 1'b0, 1'b0, n[464:463], 1'b0, 1'b0, n[460], 1'b0, 1'b0, 
        n[457:455], 1'b0, 1'b0, n[452], 1'b0, 1'b0, n[449:448], 1'b0, 1'b0, 
        n[445], 1'b0, 1'b0, n[442:438], 1'b0, 1'b0, n[435], 1'b0, 1'b0, 
        n[432:431], 1'b0, 1'b0, n[428], 1'b0, 1'b0, n[425:423], 1'b0, 1'b0, 
        n[420], 1'b0, 1'b0, n[417:416], 1'b0, 1'b0, n[413], 1'b0, 1'b0, 
        n[410:407], 1'b0, 1'b0, n[404], 1'b0, 1'b0, n[401:400], 1'b0, 1'b0, 
        n[397], 1'b0, 1'b0, n[394:392], 1'b0, 1'b0, n[389], 1'b0, 1'b0, 
        n[386:385], 1'b0, 1'b0, n[382], 1'b0, 1'b0, n[379:374], 1'b0, 1'b0, 
        n[371], 1'b0, 1'b0, n[368:367], 1'b0, 1'b0, n[364], 1'b0, 1'b0, 
        n[361:359], 1'b0, 1'b0, n[356], 1'b0, 1'b0, n[353:352], 1'b0, 1'b0, 
        n[349], 1'b0, 1'b0, n[346:343], 1'b0, 1'b0, n[340], 1'b0, 1'b0, 
        n[337:336], 1'b0, 1'b0, n[333], 1'b0, 1'b0, n[330:328], 1'b0, 1'b0, 
        n[325], 1'b0, 1'b0, n[322:321], 1'b0, 1'b0, n[318], 1'b0, 1'b0, 
        n[315:311], 1'b0, 1'b0, n[308], 1'b0, 1'b0, n[305:304], 1'b0, 1'b0, 
        n[301], 1'b0, 1'b0, n[298:296], 1'b0, 1'b0, n[293], 1'b0, 1'b0, 
        n[290:289], 1'b0, 1'b0, n[286], 1'b0, 1'b0, n[283:280], 1'b0, 1'b0, 
        n[277], 1'b0, 1'b0, n[274:273], 1'b0, 1'b0, n[270], 1'b0, 1'b0, 
        n[267:265], 1'b0, 1'b0, n[262], 1'b0, 1'b0, n[259:258], 1'b0, 1'b0, 
        n[255], 1'b0, 1'b0, n[252:246], 1'b0, 1'b0, n[243], 1'b0, 1'b0, 
        n[240:239], 1'b0, 1'b0, n[236], 1'b0, 1'b0, n[233:231], 1'b0, 1'b0, 
        n[228], 1'b0, 1'b0, n[225:224], 1'b0, 1'b0, n[221], 1'b0, 1'b0, 
        n[218:215], 1'b0, 1'b0, n[212], 1'b0, 1'b0, n[209:208], 1'b0, 1'b0, 
        n[205], 1'b0, 1'b0, n[202:200], 1'b0, 1'b0, n[197], 1'b0, 1'b0, 
        n[194:193], 1'b0, 1'b0, n[190], 1'b0, 1'b0, n[187:183], 1'b0, 1'b0, 
        n[180], 1'b0, 1'b0, n[177:176], 1'b0, 1'b0, n[173], 1'b0, 1'b0, 
        n[170:168], 1'b0, 1'b0, n[165], 1'b0, 1'b0, n[162:161], 1'b0, 1'b0, 
        n[158], 1'b0, 1'b0, n[155:152], 1'b0, 1'b0, n[149], 1'b0, 1'b0, 
        n[146:145], 1'b0, 1'b0, n[142], 1'b0, 1'b0, n[139:137], 1'b0, 1'b0, 
        n[134], 1'b0, 1'b0, n[131:130], 1'b0, 1'b0, n[127], 1'b0, 1'b0, 
        n[124:119], 1'b0, 1'b0, n[116], 1'b0, 1'b0, n[113:112], 1'b0, 1'b0, 
        n[109], 1'b0, 1'b0, n[106:104], 1'b0, 1'b0, n[101], 1'b0, 1'b0, 
        n[98:97], 1'b0, 1'b0, n[94], 1'b0, 1'b0, n[91:88], 1'b0, 1'b0, n[85], 
        1'b0, 1'b0, n[82:81], 1'b0, 1'b0, n[78], 1'b0, 1'b0, n[75:73], 1'b0, 
        1'b0, n[70], 1'b0, 1'b0, n[67:66], 1'b0, 1'b0, n[63], 1'b0, 1'b0, 
        n[60:56], 1'b0, 1'b0, n[53], 1'b0, 1'b0, n[50:49], 1'b0, 1'b0, n[46], 
        1'b0, 1'b0, n[43:41], 1'b0, 1'b0, n[38], 1'b0, 1'b0, n[35:34], 1'b0, 
        1'b0, n[31], 1'b0, 1'b0, n[28:25], 1'b0, 1'b0, n[22], 1'b0, 1'b0, 
        n[19:18], 1'b0, 1'b0, n[15], 1'b0, 1'b0, n[12:10], 1'b0, 1'b0, n[7], 
        1'b0, 1'b0, n[4:3], 1'b0, 1'b0, n[0]}), .s(s) );
endmodule

