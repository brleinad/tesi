
module gen_linear_part ( a, b, n, s );
  input [7:0] a;
  input [7:0] b;
  input [500:0] n;
  output [7:0] s;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177;

  XOR4D0 U1 ( .A1(n1), .A2(n[495]), .A3(n2), .A4(n3), .Z(s[7]) );
  XOR4D0 U2 ( .A1(n[492]), .A2(b[7]), .A3(n4), .A4(a[7]), .Z(n3) );
  XOR4D0 U3 ( .A1(n[487]), .A2(n[486]), .A3(n5), .A4(n6), .Z(n4) );
  XOR3D0 U4 ( .A1(n[485]), .A2(n7), .A3(n8), .Z(n6) );
  XOR4D0 U5 ( .A1(n[480]), .A2(n[479]), .A3(n9), .A4(n[478]), .Z(n8) );
  XOR4D0 U6 ( .A1(n[473]), .A2(n[472]), .A3(n10), .A4(n11), .Z(n9) );
  XOR3D0 U7 ( .A1(n[471]), .A2(n12), .A3(n13), .Z(n11) );
  XOR4D0 U8 ( .A1(n[466]), .A2(n[465]), .A3(n14), .A4(n[464]), .Z(n13) );
  XOR4D0 U9 ( .A1(n[459]), .A2(n[458]), .A3(n15), .A4(n16), .Z(n14) );
  XOR3D0 U10 ( .A1(n[457]), .A2(n17), .A3(n18), .Z(n16) );
  XOR4D0 U11 ( .A1(n[452]), .A2(n[451]), .A3(n19), .A4(n[450]), .Z(n18) );
  XOR4D0 U12 ( .A1(n[445]), .A2(n[444]), .A3(n20), .A4(n21), .Z(n19) );
  XOR3D0 U13 ( .A1(n[443]), .A2(n22), .A3(n23), .Z(n21) );
  XOR4D0 U14 ( .A1(n[438]), .A2(n[437]), .A3(n24), .A4(n[436]), .Z(n23) );
  XOR4D0 U15 ( .A1(n[431]), .A2(n[430]), .A3(n25), .A4(n26), .Z(n24) );
  XOR3D0 U16 ( .A1(n[429]), .A2(n27), .A3(n28), .Z(n26) );
  XOR4D0 U17 ( .A1(n[424]), .A2(n[423]), .A3(n29), .A4(n[422]), .Z(n28) );
  XOR4D0 U18 ( .A1(n[417]), .A2(n[416]), .A3(n30), .A4(n31), .Z(n29) );
  XOR3D0 U19 ( .A1(n[415]), .A2(n32), .A3(n33), .Z(n31) );
  XOR4D0 U20 ( .A1(n[410]), .A2(n[409]), .A3(n34), .A4(n[408]), .Z(n33) );
  XOR4D0 U21 ( .A1(n[403]), .A2(n[402]), .A3(n35), .A4(n36), .Z(n34) );
  XOR3D0 U22 ( .A1(n[401]), .A2(n37), .A3(n38), .Z(n36) );
  XOR4D0 U23 ( .A1(n[396]), .A2(n[395]), .A3(n39), .A4(n[394]), .Z(n38) );
  XOR4D0 U24 ( .A1(n[389]), .A2(n[388]), .A3(n40), .A4(n41), .Z(n39) );
  XOR3D0 U25 ( .A1(n[387]), .A2(n42), .A3(n43), .Z(n41) );
  XOR4D0 U26 ( .A1(n[382]), .A2(n[381]), .A3(n44), .A4(n[380]), .Z(n43) );
  XOR4D0 U27 ( .A1(n[375]), .A2(n[374]), .A3(n45), .A4(n46), .Z(n44) );
  XOR3D0 U28 ( .A1(n[373]), .A2(n47), .A3(n48), .Z(n46) );
  XOR4D0 U29 ( .A1(n[368]), .A2(n[367]), .A3(n49), .A4(n[366]), .Z(n48) );
  XOR4D0 U30 ( .A1(n[361]), .A2(n[360]), .A3(n50), .A4(n51), .Z(n49) );
  XOR3D0 U31 ( .A1(n[359]), .A2(n52), .A3(n53), .Z(n51) );
  XOR4D0 U32 ( .A1(n[354]), .A2(n[353]), .A3(n54), .A4(n[352]), .Z(n53) );
  XOR4D0 U33 ( .A1(n[347]), .A2(n[346]), .A3(n55), .A4(n56), .Z(n54) );
  XOR3D0 U34 ( .A1(n[345]), .A2(n57), .A3(n58), .Z(n56) );
  XOR4D0 U35 ( .A1(n[340]), .A2(n[339]), .A3(n59), .A4(n[338]), .Z(n58) );
  XOR4D0 U36 ( .A1(n[333]), .A2(n[332]), .A3(n60), .A4(n61), .Z(n59) );
  XOR3D0 U37 ( .A1(n[331]), .A2(n62), .A3(n63), .Z(n61) );
  XOR4D0 U38 ( .A1(n[326]), .A2(n[325]), .A3(n64), .A4(n[324]), .Z(n63) );
  XOR4D0 U39 ( .A1(n[319]), .A2(n[318]), .A3(n65), .A4(n66), .Z(n64) );
  XOR3D0 U40 ( .A1(n[317]), .A2(n67), .A3(n68), .Z(n66) );
  XOR4D0 U41 ( .A1(n[312]), .A2(n[311]), .A3(n69), .A4(n[310]), .Z(n68) );
  XOR4D0 U42 ( .A1(n[305]), .A2(n[304]), .A3(n70), .A4(n71), .Z(n69) );
  XOR3D0 U43 ( .A1(n[303]), .A2(n72), .A3(n73), .Z(n71) );
  XOR4D0 U44 ( .A1(n[298]), .A2(n[297]), .A3(n74), .A4(n[296]), .Z(n73) );
  XOR4D0 U45 ( .A1(n[291]), .A2(n[290]), .A3(n75), .A4(n76), .Z(n74) );
  XOR3D0 U46 ( .A1(n[289]), .A2(n77), .A3(n78), .Z(n76) );
  XOR4D0 U47 ( .A1(n[284]), .A2(n[283]), .A3(n79), .A4(n[282]), .Z(n78) );
  XOR4D0 U48 ( .A1(n[277]), .A2(n[276]), .A3(n80), .A4(n81), .Z(n79) );
  XOR3D0 U49 ( .A1(n[275]), .A2(n82), .A3(n83), .Z(n81) );
  XOR3D0 U50 ( .A1(n[270]), .A2(n[269]), .A3(n84), .Z(n83) );
  XOR3D0 U51 ( .A1(n85), .A2(n[268]), .A3(n86), .Z(n84) );
  XOR4D0 U52 ( .A1(n[263]), .A2(n[262]), .A3(n87), .A4(n[261]), .Z(n86) );
  XOR4D0 U53 ( .A1(n[256]), .A2(n[255]), .A3(n88), .A4(n89), .Z(n87) );
  XOR3D0 U54 ( .A1(n[254]), .A2(n90), .A3(n91), .Z(n89) );
  XNR4D0 U55 ( .A1(n[247]), .A2(n[246]), .A3(n[249]), .A4(n[248]), .ZN(n91) );
  XNR4D0 U56 ( .A1(n[251]), .A2(n[250]), .A3(n[253]), .A4(n[252]), .ZN(n90) );
  XNR4D0 U57 ( .A1(n[258]), .A2(n[257]), .A3(n[260]), .A4(n[259]), .ZN(n88) );
  XOR4D0 U58 ( .A1(n[265]), .A2(n[264]), .A3(n[267]), .A4(n[266]), .Z(n85) );
  XNR4D0 U59 ( .A1(n[272]), .A2(n[271]), .A3(n[274]), .A4(n[273]), .ZN(n82) );
  XNR4D0 U60 ( .A1(n[279]), .A2(n[278]), .A3(n[281]), .A4(n[280]), .ZN(n80) );
  XNR4D0 U61 ( .A1(n[286]), .A2(n[285]), .A3(n[288]), .A4(n[287]), .ZN(n77) );
  XNR4D0 U62 ( .A1(n[293]), .A2(n[292]), .A3(n[295]), .A4(n[294]), .ZN(n75) );
  XNR4D0 U63 ( .A1(n[300]), .A2(n[299]), .A3(n[302]), .A4(n[301]), .ZN(n72) );
  XNR4D0 U64 ( .A1(n[307]), .A2(n[306]), .A3(n[309]), .A4(n[308]), .ZN(n70) );
  XNR4D0 U65 ( .A1(n[314]), .A2(n[313]), .A3(n[316]), .A4(n[315]), .ZN(n67) );
  XNR4D0 U66 ( .A1(n[321]), .A2(n[320]), .A3(n[323]), .A4(n[322]), .ZN(n65) );
  XNR4D0 U67 ( .A1(n[328]), .A2(n[327]), .A3(n[330]), .A4(n[329]), .ZN(n62) );
  XNR4D0 U68 ( .A1(n[335]), .A2(n[334]), .A3(n[337]), .A4(n[336]), .ZN(n60) );
  XNR4D0 U69 ( .A1(n[342]), .A2(n[341]), .A3(n[344]), .A4(n[343]), .ZN(n57) );
  XNR4D0 U70 ( .A1(n[349]), .A2(n[348]), .A3(n[351]), .A4(n[350]), .ZN(n55) );
  XNR4D0 U71 ( .A1(n[356]), .A2(n[355]), .A3(n[358]), .A4(n[357]), .ZN(n52) );
  XNR4D0 U72 ( .A1(n[363]), .A2(n[362]), .A3(n[365]), .A4(n[364]), .ZN(n50) );
  XNR4D0 U73 ( .A1(n[370]), .A2(n[369]), .A3(n[372]), .A4(n[371]), .ZN(n47) );
  XNR4D0 U74 ( .A1(n[377]), .A2(n[376]), .A3(n[379]), .A4(n[378]), .ZN(n45) );
  XNR4D0 U75 ( .A1(n[384]), .A2(n[383]), .A3(n[386]), .A4(n[385]), .ZN(n42) );
  XNR4D0 U76 ( .A1(n[391]), .A2(n[390]), .A3(n[393]), .A4(n[392]), .ZN(n40) );
  XNR4D0 U77 ( .A1(n[398]), .A2(n[397]), .A3(n[400]), .A4(n[399]), .ZN(n37) );
  XNR4D0 U78 ( .A1(n[405]), .A2(n[404]), .A3(n[407]), .A4(n[406]), .ZN(n35) );
  XNR4D0 U79 ( .A1(n[412]), .A2(n[411]), .A3(n[414]), .A4(n[413]), .ZN(n32) );
  XNR4D0 U80 ( .A1(n[419]), .A2(n[418]), .A3(n[421]), .A4(n[420]), .ZN(n30) );
  XNR4D0 U81 ( .A1(n[426]), .A2(n[425]), .A3(n[428]), .A4(n[427]), .ZN(n27) );
  XNR4D0 U82 ( .A1(n[433]), .A2(n[432]), .A3(n[435]), .A4(n[434]), .ZN(n25) );
  XNR4D0 U83 ( .A1(n[440]), .A2(n[439]), .A3(n[442]), .A4(n[441]), .ZN(n22) );
  XNR4D0 U84 ( .A1(n[447]), .A2(n[446]), .A3(n[449]), .A4(n[448]), .ZN(n20) );
  XNR4D0 U85 ( .A1(n[454]), .A2(n[453]), .A3(n[456]), .A4(n[455]), .ZN(n17) );
  XNR4D0 U86 ( .A1(n[461]), .A2(n[460]), .A3(n[463]), .A4(n[462]), .ZN(n15) );
  XNR4D0 U87 ( .A1(n[468]), .A2(n[467]), .A3(n[470]), .A4(n[469]), .ZN(n12) );
  XNR4D0 U88 ( .A1(n[475]), .A2(n[474]), .A3(n[477]), .A4(n[476]), .ZN(n10) );
  XNR4D0 U89 ( .A1(n[482]), .A2(n[481]), .A3(n[484]), .A4(n[483]), .ZN(n7) );
  XNR4D0 U90 ( .A1(n[489]), .A2(n[488]), .A3(n[491]), .A4(n[490]), .ZN(n5) );
  XNR3D0 U91 ( .A1(n[498]), .A2(n[497]), .A3(n[496]), .ZN(n2) );
  XOR4D0 U92 ( .A1(n[494]), .A2(n[493]), .A3(n[500]), .A4(n[499]), .Z(n1) );
  XOR4D0 U93 ( .A1(b[6]), .A2(a[6]), .A3(n92), .A4(n93), .Z(s[6]) );
  XOR4D0 U94 ( .A1(n[241]), .A2(n[240]), .A3(n94), .A4(n[239]), .Z(n93) );
  XOR4D0 U95 ( .A1(n[234]), .A2(n[233]), .A3(n95), .A4(n96), .Z(n94) );
  XOR3D0 U96 ( .A1(n[232]), .A2(n97), .A3(n98), .Z(n96) );
  XOR4D0 U97 ( .A1(n[227]), .A2(n[226]), .A3(n99), .A4(n[225]), .Z(n98) );
  XOR4D0 U98 ( .A1(n[220]), .A2(n[219]), .A3(n100), .A4(n101), .Z(n99) );
  XOR3D0 U99 ( .A1(n[218]), .A2(n102), .A3(n103), .Z(n101) );
  XOR4D0 U100 ( .A1(n[213]), .A2(n[212]), .A3(n104), .A4(n[211]), .Z(n103) );
  XOR4D0 U101 ( .A1(n[206]), .A2(n[205]), .A3(n105), .A4(n106), .Z(n104) );
  XOR3D0 U102 ( .A1(n[204]), .A2(n107), .A3(n108), .Z(n106) );
  XOR4D0 U103 ( .A1(n[199]), .A2(n[198]), .A3(n109), .A4(n[197]), .Z(n108) );
  XOR4D0 U104 ( .A1(n[192]), .A2(n[191]), .A3(n110), .A4(n111), .Z(n109) );
  XOR3D0 U105 ( .A1(n[190]), .A2(n112), .A3(n113), .Z(n111) );
  XOR4D0 U106 ( .A1(n[185]), .A2(n[184]), .A3(n114), .A4(n[183]), .Z(n113) );
  XOR4D0 U107 ( .A1(n[178]), .A2(n[177]), .A3(n115), .A4(n116), .Z(n114) );
  XOR3D0 U108 ( .A1(n[176]), .A2(n117), .A3(n118), .Z(n116) );
  XOR4D0 U109 ( .A1(n[171]), .A2(n[170]), .A3(n119), .A4(n[169]), .Z(n118) );
  XOR4D0 U110 ( .A1(n[164]), .A2(n[163]), .A3(n120), .A4(n121), .Z(n119) );
  XOR3D0 U111 ( .A1(n[162]), .A2(n122), .A3(n123), .Z(n121) );
  XOR4D0 U112 ( .A1(n[157]), .A2(n[156]), .A3(n124), .A4(n[155]), .Z(n123) );
  XOR4D0 U113 ( .A1(n[150]), .A2(n[149]), .A3(n125), .A4(n126), .Z(n124) );
  XOR3D0 U114 ( .A1(n[148]), .A2(n127), .A3(n128), .Z(n126) );
  XOR3D0 U115 ( .A1(n[143]), .A2(n[142]), .A3(n129), .Z(n128) );
  XOR3D0 U116 ( .A1(n130), .A2(n[141]), .A3(n131), .Z(n129) );
  XOR4D0 U117 ( .A1(n[136]), .A2(n[135]), .A3(n132), .A4(n[134]), .Z(n131) );
  XOR4D0 U118 ( .A1(n[129]), .A2(n[128]), .A3(n133), .A4(n134), .Z(n132) );
  XOR3D0 U119 ( .A1(n[127]), .A2(n135), .A3(n136), .Z(n134) );
  XNR4D0 U120 ( .A1(n[120]), .A2(n[119]), .A3(n[122]), .A4(n[121]), .ZN(n136)
         );
  XNR4D0 U121 ( .A1(n[124]), .A2(n[123]), .A3(n[126]), .A4(n[125]), .ZN(n135)
         );
  XNR4D0 U122 ( .A1(n[131]), .A2(n[130]), .A3(n[133]), .A4(n[132]), .ZN(n133)
         );
  XOR4D0 U123 ( .A1(n[138]), .A2(n[137]), .A3(n[140]), .A4(n[139]), .Z(n130)
         );
  XNR4D0 U124 ( .A1(n[145]), .A2(n[144]), .A3(n[147]), .A4(n[146]), .ZN(n127)
         );
  XNR4D0 U125 ( .A1(n[152]), .A2(n[151]), .A3(n[154]), .A4(n[153]), .ZN(n125)
         );
  XNR4D0 U126 ( .A1(n[159]), .A2(n[158]), .A3(n[161]), .A4(n[160]), .ZN(n122)
         );
  XNR4D0 U127 ( .A1(n[166]), .A2(n[165]), .A3(n[168]), .A4(n[167]), .ZN(n120)
         );
  XNR4D0 U128 ( .A1(n[173]), .A2(n[172]), .A3(n[175]), .A4(n[174]), .ZN(n117)
         );
  XNR4D0 U129 ( .A1(n[180]), .A2(n[179]), .A3(n[182]), .A4(n[181]), .ZN(n115)
         );
  XNR4D0 U130 ( .A1(n[187]), .A2(n[186]), .A3(n[189]), .A4(n[188]), .ZN(n112)
         );
  XNR4D0 U131 ( .A1(n[194]), .A2(n[193]), .A3(n[196]), .A4(n[195]), .ZN(n110)
         );
  XNR4D0 U132 ( .A1(n[201]), .A2(n[200]), .A3(n[203]), .A4(n[202]), .ZN(n107)
         );
  XNR4D0 U133 ( .A1(n[208]), .A2(n[207]), .A3(n[210]), .A4(n[209]), .ZN(n105)
         );
  XNR4D0 U134 ( .A1(n[215]), .A2(n[214]), .A3(n[217]), .A4(n[216]), .ZN(n102)
         );
  XNR4D0 U135 ( .A1(n[222]), .A2(n[221]), .A3(n[224]), .A4(n[223]), .ZN(n100)
         );
  XNR4D0 U136 ( .A1(n[229]), .A2(n[228]), .A3(n[231]), .A4(n[230]), .ZN(n97)
         );
  XNR4D0 U137 ( .A1(n[236]), .A2(n[235]), .A3(n[238]), .A4(n[237]), .ZN(n95)
         );
  XNR4D0 U138 ( .A1(n[243]), .A2(n[242]), .A3(n[245]), .A4(n[244]), .ZN(n92)
         );
  XOR3D0 U139 ( .A1(n[118]), .A2(n137), .A3(n138), .Z(s[5]) );
  XOR4D0 U140 ( .A1(n[113]), .A2(b[5]), .A3(n139), .A4(a[5]), .Z(n138) );
  XOR4D0 U141 ( .A1(n[108]), .A2(n[107]), .A3(n140), .A4(n141), .Z(n139) );
  XOR3D0 U142 ( .A1(n[106]), .A2(n142), .A3(n143), .Z(n141) );
  XOR4D0 U143 ( .A1(n[102]), .A2(n[101]), .A3(n144), .A4(n[100]), .Z(n143) );
  XOR4D0 U144 ( .A1(n[94]), .A2(n[93]), .A3(n145), .A4(n146), .Z(n144) );
  XOR3D0 U145 ( .A1(n[92]), .A2(n147), .A3(n148), .Z(n146) );
  XOR4D0 U146 ( .A1(n[87]), .A2(n[86]), .A3(n149), .A4(n[85]), .Z(n148) );
  XOR4D0 U147 ( .A1(n[80]), .A2(n[79]), .A3(n150), .A4(n151), .Z(n149) );
  XOR3D0 U148 ( .A1(n[78]), .A2(n152), .A3(n153), .Z(n151) );
  XOR4D0 U149 ( .A1(n[73]), .A2(n[72]), .A3(n154), .A4(n[71]), .Z(n153) );
  XOR4D0 U150 ( .A1(n[66]), .A2(n[65]), .A3(n155), .A4(n156), .Z(n154) );
  XOR3D0 U151 ( .A1(n[64]), .A2(n157), .A3(n158), .Z(n156) );
  XNR4D0 U152 ( .A1(n[57]), .A2(n[56]), .A3(n[59]), .A4(n[58]), .ZN(n158) );
  XNR4D0 U153 ( .A1(n[61]), .A2(n[60]), .A3(n[63]), .A4(n[62]), .ZN(n157) );
  XNR4D0 U154 ( .A1(n[68]), .A2(n[67]), .A3(n[70]), .A4(n[69]), .ZN(n155) );
  XNR4D0 U155 ( .A1(n[75]), .A2(n[74]), .A3(n[77]), .A4(n[76]), .ZN(n152) );
  XNR4D0 U156 ( .A1(n[82]), .A2(n[81]), .A3(n[84]), .A4(n[83]), .ZN(n150) );
  XNR4D0 U157 ( .A1(n[89]), .A2(n[88]), .A3(n[91]), .A4(n[90]), .ZN(n147) );
  XNR4D0 U158 ( .A1(n[96]), .A2(n[95]), .A3(n[98]), .A4(n[97]), .ZN(n145) );
  XNR4D0 U159 ( .A1(n[104]), .A2(n[103]), .A3(n[99]), .A4(n[105]), .ZN(n142)
         );
  XNR4D0 U160 ( .A1(n[110]), .A2(n[109]), .A3(n[112]), .A4(n[111]), .ZN(n140)
         );
  XNR4D0 U161 ( .A1(n[115]), .A2(n[114]), .A3(n[117]), .A4(n[116]), .ZN(n137)
         );
  XOR4D0 U162 ( .A1(n159), .A2(n[50]), .A3(n160), .A4(n161), .Z(s[4]) );
  XOR3D0 U163 ( .A1(n[47]), .A2(b[4]), .A3(n162), .Z(n161) );
  XOR3D0 U164 ( .A1(n163), .A2(a[4]), .A3(n164), .Z(n162) );
  XOR4D0 U165 ( .A1(n[42]), .A2(n[41]), .A3(n165), .A4(n[40]), .Z(n164) );
  XOR4D0 U166 ( .A1(n[35]), .A2(n[34]), .A3(n166), .A4(n167), .Z(n165) );
  XOR3D0 U167 ( .A1(n[33]), .A2(n168), .A3(n169), .Z(n167) );
  XNR4D0 U168 ( .A1(n[26]), .A2(n[25]), .A3(n[28]), .A4(n[27]), .ZN(n169) );
  XNR4D0 U169 ( .A1(n[30]), .A2(n[29]), .A3(n[32]), .A4(n[31]), .ZN(n168) );
  XNR4D0 U170 ( .A1(n[37]), .A2(n[36]), .A3(n[39]), .A4(n[38]), .ZN(n166) );
  XOR4D0 U171 ( .A1(n[44]), .A2(n[43]), .A3(n[46]), .A4(n[45]), .Z(n163) );
  XNR3D0 U172 ( .A1(n[53]), .A2(n[52]), .A3(n[51]), .ZN(n160) );
  XOR4D0 U173 ( .A1(n[49]), .A2(n[48]), .A3(n[55]), .A4(n[54]), .Z(n159) );
  XOR4D0 U174 ( .A1(b[3]), .A2(a[3]), .A3(n170), .A4(n171), .Z(s[3]) );
  XOR3D0 U175 ( .A1(n[20]), .A2(n[19]), .A3(n172), .Z(n171) );
  XOR3D0 U176 ( .A1(n[18]), .A2(n173), .A3(n174), .Z(n172) );
  XNR4D0 U177 ( .A1(n[11]), .A2(n[10]), .A3(n[13]), .A4(n[12]), .ZN(n174) );
  XNR4D0 U178 ( .A1(n[15]), .A2(n[14]), .A3(n[17]), .A4(n[16]), .ZN(n173) );
  XOR4D0 U179 ( .A1(n[22]), .A2(n[21]), .A3(n[24]), .A4(n[23]), .Z(n170) );
  XOR3D0 U180 ( .A1(n[9]), .A2(n175), .A3(n176), .Z(s[2]) );
  XNR4D0 U181 ( .A1(b[2]), .A2(a[2]), .A3(n[4]), .A4(n[3]), .ZN(n176) );
  XNR4D0 U182 ( .A1(n[6]), .A2(n[5]), .A3(n[8]), .A4(n[7]), .ZN(n175) );
  XOR3D0 U183 ( .A1(b[1]), .A2(a[1]), .A3(n177), .Z(s[1]) );
  XOR3D0 U184 ( .A1(n[2]), .A2(n[1]), .A3(n[0]), .Z(n177) );
  CKXOR2D0 U185 ( .A1(b[0]), .A2(a[0]), .Z(s[0]) );
endmodule


module gen_nonlinear_part ( a, b, n );
  input [7:0] a;
  input [7:0] b;
  output [500:0] n;
  wire   n2, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320;

  TIEH U2 ( .Z(n2) );
  INVD1 U3 ( .I(n2), .ZN(n[1]) );
  INVD1 U4 ( .I(n2), .ZN(n[2]) );
  INVD1 U5 ( .I(n2), .ZN(n[5]) );
  INVD1 U6 ( .I(n2), .ZN(n[6]) );
  INVD1 U7 ( .I(n2), .ZN(n[8]) );
  INVD1 U8 ( .I(n2), .ZN(n[9]) );
  INVD1 U9 ( .I(n2), .ZN(n[13]) );
  INVD1 U10 ( .I(n2), .ZN(n[14]) );
  INVD1 U11 ( .I(n2), .ZN(n[16]) );
  INVD1 U12 ( .I(n2), .ZN(n[17]) );
  INVD1 U13 ( .I(n2), .ZN(n[20]) );
  INVD1 U14 ( .I(n2), .ZN(n[21]) );
  INVD1 U15 ( .I(n2), .ZN(n[23]) );
  INVD1 U16 ( .I(n2), .ZN(n[24]) );
  INVD1 U17 ( .I(n2), .ZN(n[29]) );
  INVD1 U18 ( .I(n2), .ZN(n[30]) );
  INVD1 U19 ( .I(n2), .ZN(n[32]) );
  INVD1 U20 ( .I(n2), .ZN(n[33]) );
  INVD1 U21 ( .I(n2), .ZN(n[36]) );
  INVD1 U22 ( .I(n2), .ZN(n[37]) );
  INVD1 U23 ( .I(n2), .ZN(n[39]) );
  INVD1 U24 ( .I(n2), .ZN(n[40]) );
  INVD1 U25 ( .I(n2), .ZN(n[44]) );
  INVD1 U26 ( .I(n2), .ZN(n[45]) );
  INVD1 U27 ( .I(n2), .ZN(n[47]) );
  INVD1 U28 ( .I(n2), .ZN(n[48]) );
  INVD1 U29 ( .I(n2), .ZN(n[51]) );
  INVD1 U30 ( .I(n2), .ZN(n[52]) );
  INVD1 U31 ( .I(n2), .ZN(n[54]) );
  INVD1 U32 ( .I(n2), .ZN(n[55]) );
  INVD1 U33 ( .I(n2), .ZN(n[61]) );
  INVD1 U34 ( .I(n2), .ZN(n[62]) );
  INVD1 U35 ( .I(n2), .ZN(n[64]) );
  INVD1 U36 ( .I(n2), .ZN(n[65]) );
  INVD1 U37 ( .I(n2), .ZN(n[68]) );
  INVD1 U38 ( .I(n2), .ZN(n[69]) );
  INVD1 U39 ( .I(n2), .ZN(n[71]) );
  INVD1 U40 ( .I(n2), .ZN(n[72]) );
  INVD1 U41 ( .I(n2), .ZN(n[76]) );
  INVD1 U42 ( .I(n2), .ZN(n[77]) );
  INVD1 U43 ( .I(n2), .ZN(n[79]) );
  INVD1 U44 ( .I(n2), .ZN(n[80]) );
  INVD1 U45 ( .I(n2), .ZN(n[83]) );
  INVD1 U46 ( .I(n2), .ZN(n[84]) );
  INVD1 U47 ( .I(n2), .ZN(n[86]) );
  INVD1 U48 ( .I(n2), .ZN(n[87]) );
  INVD1 U49 ( .I(n2), .ZN(n[92]) );
  INVD1 U50 ( .I(n2), .ZN(n[93]) );
  INVD1 U51 ( .I(n2), .ZN(n[95]) );
  INVD1 U52 ( .I(n2), .ZN(n[96]) );
  INVD1 U53 ( .I(n2), .ZN(n[99]) );
  INVD1 U54 ( .I(n2), .ZN(n[100]) );
  INVD1 U55 ( .I(n2), .ZN(n[102]) );
  INVD1 U56 ( .I(n2), .ZN(n[103]) );
  INVD1 U57 ( .I(n2), .ZN(n[107]) );
  INVD1 U58 ( .I(n2), .ZN(n[108]) );
  INVD1 U59 ( .I(n2), .ZN(n[110]) );
  INVD1 U60 ( .I(n2), .ZN(n[111]) );
  INVD1 U61 ( .I(n2), .ZN(n[114]) );
  INVD1 U62 ( .I(n2), .ZN(n[115]) );
  INVD1 U63 ( .I(n2), .ZN(n[117]) );
  INVD1 U64 ( .I(n2), .ZN(n[118]) );
  INVD1 U65 ( .I(n2), .ZN(n[125]) );
  INVD1 U66 ( .I(n2), .ZN(n[126]) );
  INVD1 U67 ( .I(n2), .ZN(n[128]) );
  INVD1 U68 ( .I(n2), .ZN(n[129]) );
  INVD1 U69 ( .I(n2), .ZN(n[132]) );
  INVD1 U70 ( .I(n2), .ZN(n[133]) );
  INVD1 U71 ( .I(n2), .ZN(n[135]) );
  INVD1 U72 ( .I(n2), .ZN(n[136]) );
  INVD1 U73 ( .I(n2), .ZN(n[140]) );
  INVD1 U74 ( .I(n2), .ZN(n[141]) );
  INVD1 U75 ( .I(n2), .ZN(n[143]) );
  INVD1 U76 ( .I(n2), .ZN(n[144]) );
  INVD1 U77 ( .I(n2), .ZN(n[147]) );
  INVD1 U78 ( .I(n2), .ZN(n[148]) );
  INVD1 U79 ( .I(n2), .ZN(n[150]) );
  INVD1 U80 ( .I(n2), .ZN(n[151]) );
  INVD1 U81 ( .I(n2), .ZN(n[156]) );
  INVD1 U82 ( .I(n2), .ZN(n[157]) );
  INVD1 U83 ( .I(n2), .ZN(n[159]) );
  INVD1 U84 ( .I(n2), .ZN(n[160]) );
  INVD1 U85 ( .I(n2), .ZN(n[163]) );
  INVD1 U86 ( .I(n2), .ZN(n[164]) );
  INVD1 U87 ( .I(n2), .ZN(n[166]) );
  INVD1 U88 ( .I(n2), .ZN(n[167]) );
  INVD1 U89 ( .I(n2), .ZN(n[171]) );
  INVD1 U90 ( .I(n2), .ZN(n[172]) );
  INVD1 U91 ( .I(n2), .ZN(n[174]) );
  INVD1 U92 ( .I(n2), .ZN(n[175]) );
  INVD1 U93 ( .I(n2), .ZN(n[178]) );
  INVD1 U94 ( .I(n2), .ZN(n[179]) );
  INVD1 U95 ( .I(n2), .ZN(n[181]) );
  INVD1 U96 ( .I(n2), .ZN(n[182]) );
  INVD1 U97 ( .I(n2), .ZN(n[188]) );
  INVD1 U98 ( .I(n2), .ZN(n[189]) );
  INVD1 U99 ( .I(n2), .ZN(n[191]) );
  INVD1 U100 ( .I(n2), .ZN(n[192]) );
  INVD1 U101 ( .I(n2), .ZN(n[195]) );
  INVD1 U102 ( .I(n2), .ZN(n[196]) );
  INVD1 U103 ( .I(n2), .ZN(n[198]) );
  INVD1 U104 ( .I(n2), .ZN(n[199]) );
  INVD1 U105 ( .I(n2), .ZN(n[203]) );
  INVD1 U106 ( .I(n2), .ZN(n[204]) );
  INVD1 U107 ( .I(n2), .ZN(n[206]) );
  INVD1 U108 ( .I(n2), .ZN(n[207]) );
  INVD1 U109 ( .I(n2), .ZN(n[210]) );
  INVD1 U110 ( .I(n2), .ZN(n[211]) );
  INVD1 U111 ( .I(n2), .ZN(n[213]) );
  INVD1 U112 ( .I(n2), .ZN(n[214]) );
  INVD1 U113 ( .I(n2), .ZN(n[219]) );
  INVD1 U114 ( .I(n2), .ZN(n[220]) );
  INVD1 U115 ( .I(n2), .ZN(n[222]) );
  INVD1 U116 ( .I(n2), .ZN(n[223]) );
  INVD1 U117 ( .I(n2), .ZN(n[226]) );
  INVD1 U118 ( .I(n2), .ZN(n[227]) );
  INVD1 U119 ( .I(n2), .ZN(n[229]) );
  INVD1 U120 ( .I(n2), .ZN(n[230]) );
  INVD1 U121 ( .I(n2), .ZN(n[234]) );
  INVD1 U122 ( .I(n2), .ZN(n[235]) );
  INVD1 U123 ( .I(n2), .ZN(n[237]) );
  INVD1 U124 ( .I(n2), .ZN(n[238]) );
  INVD1 U125 ( .I(n2), .ZN(n[241]) );
  INVD1 U126 ( .I(n2), .ZN(n[242]) );
  INVD1 U127 ( .I(n2), .ZN(n[244]) );
  INVD1 U128 ( .I(n2), .ZN(n[245]) );
  INVD1 U129 ( .I(n2), .ZN(n[253]) );
  INVD1 U130 ( .I(n2), .ZN(n[254]) );
  INVD1 U131 ( .I(n2), .ZN(n[256]) );
  INVD1 U132 ( .I(n2), .ZN(n[257]) );
  INVD1 U133 ( .I(n2), .ZN(n[260]) );
  INVD1 U134 ( .I(n2), .ZN(n[261]) );
  INVD1 U135 ( .I(n2), .ZN(n[263]) );
  INVD1 U136 ( .I(n2), .ZN(n[264]) );
  INVD1 U137 ( .I(n2), .ZN(n[268]) );
  INVD1 U138 ( .I(n2), .ZN(n[269]) );
  INVD1 U139 ( .I(n2), .ZN(n[271]) );
  INVD1 U140 ( .I(n2), .ZN(n[272]) );
  INVD1 U141 ( .I(n2), .ZN(n[275]) );
  INVD1 U142 ( .I(n2), .ZN(n[276]) );
  INVD1 U143 ( .I(n2), .ZN(n[278]) );
  INVD1 U144 ( .I(n2), .ZN(n[279]) );
  INVD1 U145 ( .I(n2), .ZN(n[284]) );
  INVD1 U146 ( .I(n2), .ZN(n[285]) );
  INVD1 U147 ( .I(n2), .ZN(n[287]) );
  INVD1 U148 ( .I(n2), .ZN(n[288]) );
  INVD1 U149 ( .I(n2), .ZN(n[291]) );
  INVD1 U150 ( .I(n2), .ZN(n[292]) );
  INVD1 U151 ( .I(n2), .ZN(n[294]) );
  INVD1 U152 ( .I(n2), .ZN(n[295]) );
  INVD1 U153 ( .I(n2), .ZN(n[299]) );
  INVD1 U154 ( .I(n2), .ZN(n[300]) );
  INVD1 U155 ( .I(n2), .ZN(n[302]) );
  INVD1 U156 ( .I(n2), .ZN(n[303]) );
  INVD1 U157 ( .I(n2), .ZN(n[306]) );
  INVD1 U158 ( .I(n2), .ZN(n[307]) );
  INVD1 U159 ( .I(n2), .ZN(n[309]) );
  INVD1 U160 ( .I(n2), .ZN(n[310]) );
  INVD1 U161 ( .I(n2), .ZN(n[316]) );
  INVD1 U162 ( .I(n2), .ZN(n[317]) );
  INVD1 U163 ( .I(n2), .ZN(n[319]) );
  INVD1 U164 ( .I(n2), .ZN(n[320]) );
  INVD1 U165 ( .I(n2), .ZN(n[323]) );
  INVD1 U166 ( .I(n2), .ZN(n[324]) );
  INVD1 U167 ( .I(n2), .ZN(n[326]) );
  INVD1 U168 ( .I(n2), .ZN(n[327]) );
  INVD1 U169 ( .I(n2), .ZN(n[331]) );
  INVD1 U170 ( .I(n2), .ZN(n[332]) );
  INVD1 U171 ( .I(n2), .ZN(n[334]) );
  INVD1 U172 ( .I(n2), .ZN(n[335]) );
  INVD1 U173 ( .I(n2), .ZN(n[338]) );
  INVD1 U174 ( .I(n2), .ZN(n[339]) );
  INVD1 U175 ( .I(n2), .ZN(n[341]) );
  INVD1 U176 ( .I(n2), .ZN(n[342]) );
  INVD1 U177 ( .I(n2), .ZN(n[347]) );
  INVD1 U178 ( .I(n2), .ZN(n[348]) );
  INVD1 U179 ( .I(n2), .ZN(n[350]) );
  INVD1 U180 ( .I(n2), .ZN(n[351]) );
  INVD1 U181 ( .I(n2), .ZN(n[354]) );
  INVD1 U182 ( .I(n2), .ZN(n[355]) );
  INVD1 U183 ( .I(n2), .ZN(n[357]) );
  INVD1 U184 ( .I(n2), .ZN(n[358]) );
  INVD1 U185 ( .I(n2), .ZN(n[362]) );
  INVD1 U186 ( .I(n2), .ZN(n[363]) );
  INVD1 U187 ( .I(n2), .ZN(n[365]) );
  INVD1 U188 ( .I(n2), .ZN(n[366]) );
  INVD1 U189 ( .I(n2), .ZN(n[369]) );
  INVD1 U190 ( .I(n2), .ZN(n[370]) );
  INVD1 U191 ( .I(n2), .ZN(n[372]) );
  INVD1 U192 ( .I(n2), .ZN(n[373]) );
  INVD1 U193 ( .I(n2), .ZN(n[380]) );
  INVD1 U194 ( .I(n2), .ZN(n[381]) );
  INVD1 U195 ( .I(n2), .ZN(n[383]) );
  INVD1 U196 ( .I(n2), .ZN(n[384]) );
  INVD1 U197 ( .I(n2), .ZN(n[387]) );
  INVD1 U198 ( .I(n2), .ZN(n[388]) );
  INVD1 U199 ( .I(n2), .ZN(n[390]) );
  INVD1 U200 ( .I(n2), .ZN(n[391]) );
  INVD1 U201 ( .I(n2), .ZN(n[395]) );
  INVD1 U202 ( .I(n2), .ZN(n[396]) );
  INVD1 U203 ( .I(n2), .ZN(n[398]) );
  INVD1 U204 ( .I(n2), .ZN(n[399]) );
  INVD1 U205 ( .I(n2), .ZN(n[402]) );
  INVD1 U206 ( .I(n2), .ZN(n[403]) );
  INVD1 U207 ( .I(n2), .ZN(n[405]) );
  INVD1 U208 ( .I(n2), .ZN(n[406]) );
  INVD1 U209 ( .I(n2), .ZN(n[411]) );
  INVD1 U210 ( .I(n2), .ZN(n[412]) );
  INVD1 U211 ( .I(n2), .ZN(n[414]) );
  INVD1 U212 ( .I(n2), .ZN(n[415]) );
  INVD1 U213 ( .I(n2), .ZN(n[418]) );
  INVD1 U214 ( .I(n2), .ZN(n[419]) );
  INVD1 U215 ( .I(n2), .ZN(n[421]) );
  INVD1 U216 ( .I(n2), .ZN(n[422]) );
  INVD1 U217 ( .I(n2), .ZN(n[426]) );
  INVD1 U218 ( .I(n2), .ZN(n[427]) );
  INVD1 U219 ( .I(n2), .ZN(n[429]) );
  INVD1 U220 ( .I(n2), .ZN(n[430]) );
  INVD1 U221 ( .I(n2), .ZN(n[433]) );
  INVD1 U222 ( .I(n2), .ZN(n[434]) );
  INVD1 U223 ( .I(n2), .ZN(n[436]) );
  INVD1 U224 ( .I(n2), .ZN(n[437]) );
  INVD1 U225 ( .I(n2), .ZN(n[443]) );
  INVD1 U226 ( .I(n2), .ZN(n[444]) );
  INVD1 U227 ( .I(n2), .ZN(n[446]) );
  INVD1 U228 ( .I(n2), .ZN(n[447]) );
  INVD1 U229 ( .I(n2), .ZN(n[450]) );
  INVD1 U230 ( .I(n2), .ZN(n[451]) );
  INVD1 U231 ( .I(n2), .ZN(n[453]) );
  INVD1 U232 ( .I(n2), .ZN(n[454]) );
  INVD1 U233 ( .I(n2), .ZN(n[458]) );
  INVD1 U234 ( .I(n2), .ZN(n[459]) );
  INVD1 U235 ( .I(n2), .ZN(n[461]) );
  INVD1 U236 ( .I(n2), .ZN(n[462]) );
  INVD1 U237 ( .I(n2), .ZN(n[465]) );
  INVD1 U238 ( .I(n2), .ZN(n[466]) );
  INVD1 U239 ( .I(n2), .ZN(n[468]) );
  INVD1 U240 ( .I(n2), .ZN(n[469]) );
  INVD1 U241 ( .I(n2), .ZN(n[474]) );
  INVD1 U242 ( .I(n2), .ZN(n[475]) );
  INVD1 U243 ( .I(n2), .ZN(n[477]) );
  INVD1 U244 ( .I(n2), .ZN(n[478]) );
  INVD1 U245 ( .I(n2), .ZN(n[481]) );
  INVD1 U246 ( .I(n2), .ZN(n[482]) );
  INVD1 U247 ( .I(n2), .ZN(n[484]) );
  INVD1 U248 ( .I(n2), .ZN(n[485]) );
  INVD1 U249 ( .I(n2), .ZN(n[489]) );
  INVD1 U250 ( .I(n2), .ZN(n[490]) );
  INVD1 U251 ( .I(n2), .ZN(n[492]) );
  INVD1 U252 ( .I(n2), .ZN(n[493]) );
  INVD1 U253 ( .I(n2), .ZN(n[496]) );
  INVD1 U254 ( .I(n2), .ZN(n[497]) );
  INVD1 U255 ( .I(n2), .ZN(n[499]) );
  INVD1 U256 ( .I(n2), .ZN(n[500]) );
  INVD1 U257 ( .I(a[6]), .ZN(n320) );
  INVD1 U258 ( .I(b[6]), .ZN(n257) );
  NR2D0 U259 ( .A1(n256), .A2(n257), .ZN(n[498]) );
  NR2D0 U260 ( .A1(n257), .A2(n258), .ZN(n[495]) );
  NR2D0 U261 ( .A1(n257), .A2(n259), .ZN(n[494]) );
  NR2D0 U262 ( .A1(n257), .A2(n260), .ZN(n[491]) );
  NR2D0 U263 ( .A1(n257), .A2(n261), .ZN(n[488]) );
  NR2D0 U264 ( .A1(n257), .A2(n262), .ZN(n[487]) );
  NR2D0 U265 ( .A1(n257), .A2(n263), .ZN(n[486]) );
  NR2D0 U266 ( .A1(n257), .A2(n264), .ZN(n[483]) );
  NR2D0 U267 ( .A1(n257), .A2(n265), .ZN(n[480]) );
  NR2D0 U268 ( .A1(n257), .A2(n266), .ZN(n[479]) );
  NR2D0 U269 ( .A1(n257), .A2(n267), .ZN(n[476]) );
  NR2D0 U270 ( .A1(n257), .A2(n268), .ZN(n[473]) );
  NR2D0 U271 ( .A1(n257), .A2(n269), .ZN(n[472]) );
  NR2D0 U272 ( .A1(n257), .A2(n270), .ZN(n[471]) );
  NR2D0 U273 ( .A1(n257), .A2(n271), .ZN(n[470]) );
  NR2D0 U274 ( .A1(n257), .A2(n272), .ZN(n[467]) );
  NR2D0 U275 ( .A1(n257), .A2(n273), .ZN(n[464]) );
  NR2D0 U276 ( .A1(n257), .A2(n274), .ZN(n[463]) );
  NR2D0 U277 ( .A1(n257), .A2(n275), .ZN(n[460]) );
  NR2D0 U278 ( .A1(n257), .A2(n276), .ZN(n[457]) );
  NR2D0 U279 ( .A1(n257), .A2(n277), .ZN(n[456]) );
  NR2D0 U280 ( .A1(n257), .A2(n278), .ZN(n[455]) );
  NR2D0 U281 ( .A1(n257), .A2(n279), .ZN(n[452]) );
  NR2D0 U282 ( .A1(n257), .A2(n280), .ZN(n[449]) );
  NR2D0 U283 ( .A1(n257), .A2(n281), .ZN(n[448]) );
  NR2D0 U284 ( .A1(n257), .A2(n282), .ZN(n[445]) );
  NR2D0 U285 ( .A1(n257), .A2(n283), .ZN(n[442]) );
  NR2D0 U286 ( .A1(n257), .A2(n284), .ZN(n[441]) );
  NR2D0 U287 ( .A1(n257), .A2(n285), .ZN(n[440]) );
  NR2D0 U288 ( .A1(n257), .A2(n286), .ZN(n[439]) );
  NR2D0 U289 ( .A1(n257), .A2(n287), .ZN(n[438]) );
  NR2D0 U290 ( .A1(n257), .A2(n288), .ZN(n[435]) );
  NR2D0 U291 ( .A1(n257), .A2(n289), .ZN(n[432]) );
  NR2D0 U292 ( .A1(n257), .A2(n290), .ZN(n[431]) );
  NR2D0 U293 ( .A1(n257), .A2(n291), .ZN(n[428]) );
  NR2D0 U294 ( .A1(n257), .A2(n292), .ZN(n[425]) );
  NR2D0 U295 ( .A1(n257), .A2(n293), .ZN(n[424]) );
  NR2D0 U296 ( .A1(n257), .A2(n294), .ZN(n[423]) );
  NR2D0 U297 ( .A1(n257), .A2(n295), .ZN(n[420]) );
  NR2D0 U298 ( .A1(n257), .A2(n296), .ZN(n[417]) );
  NR2D0 U299 ( .A1(n257), .A2(n297), .ZN(n[416]) );
  NR2D0 U300 ( .A1(n257), .A2(n298), .ZN(n[413]) );
  NR2D0 U301 ( .A1(n257), .A2(n299), .ZN(n[410]) );
  NR2D0 U302 ( .A1(n257), .A2(n300), .ZN(n[409]) );
  NR2D0 U303 ( .A1(n257), .A2(n301), .ZN(n[408]) );
  NR2D0 U304 ( .A1(n257), .A2(n302), .ZN(n[407]) );
  NR2D0 U305 ( .A1(n257), .A2(n303), .ZN(n[404]) );
  NR2D0 U306 ( .A1(n257), .A2(n304), .ZN(n[401]) );
  NR2D0 U307 ( .A1(n257), .A2(n305), .ZN(n[400]) );
  NR2D0 U308 ( .A1(n257), .A2(n306), .ZN(n[397]) );
  NR2D0 U309 ( .A1(n257), .A2(n307), .ZN(n[394]) );
  NR2D0 U310 ( .A1(n257), .A2(n308), .ZN(n[393]) );
  NR2D0 U311 ( .A1(n257), .A2(n309), .ZN(n[392]) );
  NR2D0 U312 ( .A1(n257), .A2(n310), .ZN(n[389]) );
  NR2D0 U313 ( .A1(n257), .A2(n311), .ZN(n[386]) );
  NR2D0 U314 ( .A1(n257), .A2(n312), .ZN(n[385]) );
  NR2D0 U315 ( .A1(n257), .A2(n313), .ZN(n[382]) );
  NR2D0 U316 ( .A1(n257), .A2(n314), .ZN(n[379]) );
  NR2D0 U317 ( .A1(n257), .A2(n315), .ZN(n[378]) );
  NR2D0 U318 ( .A1(n257), .A2(n316), .ZN(n[377]) );
  NR2D0 U319 ( .A1(n257), .A2(n317), .ZN(n[376]) );
  NR2D0 U320 ( .A1(n257), .A2(n318), .ZN(n[375]) );
  NR2D0 U321 ( .A1(n257), .A2(n319), .ZN(n[374]) );
  NR2D0 U322 ( .A1(n256), .A2(n320), .ZN(n[371]) );
  NR2D0 U323 ( .A1(n258), .A2(n320), .ZN(n[368]) );
  NR2D0 U324 ( .A1(n259), .A2(n320), .ZN(n[367]) );
  NR2D0 U325 ( .A1(n260), .A2(n320), .ZN(n[364]) );
  NR2D0 U326 ( .A1(n261), .A2(n320), .ZN(n[361]) );
  NR2D0 U327 ( .A1(n262), .A2(n320), .ZN(n[360]) );
  NR2D0 U328 ( .A1(n263), .A2(n320), .ZN(n[359]) );
  NR2D0 U329 ( .A1(n264), .A2(n320), .ZN(n[356]) );
  NR2D0 U330 ( .A1(n265), .A2(n320), .ZN(n[353]) );
  NR2D0 U331 ( .A1(n266), .A2(n320), .ZN(n[352]) );
  NR2D0 U332 ( .A1(n267), .A2(n320), .ZN(n[349]) );
  NR2D0 U333 ( .A1(n268), .A2(n320), .ZN(n[346]) );
  NR2D0 U334 ( .A1(n269), .A2(n320), .ZN(n[345]) );
  NR2D0 U335 ( .A1(n270), .A2(n320), .ZN(n[344]) );
  NR2D0 U336 ( .A1(n271), .A2(n320), .ZN(n[343]) );
  NR2D0 U337 ( .A1(n272), .A2(n320), .ZN(n[340]) );
  NR2D0 U338 ( .A1(n273), .A2(n320), .ZN(n[337]) );
  NR2D0 U339 ( .A1(n274), .A2(n320), .ZN(n[336]) );
  NR2D0 U340 ( .A1(n275), .A2(n320), .ZN(n[333]) );
  NR2D0 U341 ( .A1(n276), .A2(n320), .ZN(n[330]) );
  NR2D0 U342 ( .A1(n277), .A2(n320), .ZN(n[329]) );
  NR2D0 U343 ( .A1(n278), .A2(n320), .ZN(n[328]) );
  NR2D0 U344 ( .A1(n279), .A2(n320), .ZN(n[325]) );
  NR2D0 U345 ( .A1(n280), .A2(n320), .ZN(n[322]) );
  NR2D0 U346 ( .A1(n281), .A2(n320), .ZN(n[321]) );
  NR2D0 U347 ( .A1(n282), .A2(n320), .ZN(n[318]) );
  NR2D0 U348 ( .A1(n283), .A2(n320), .ZN(n[315]) );
  NR2D0 U349 ( .A1(n284), .A2(n320), .ZN(n[314]) );
  NR2D0 U350 ( .A1(n285), .A2(n320), .ZN(n[313]) );
  NR2D0 U351 ( .A1(n286), .A2(n320), .ZN(n[312]) );
  NR2D0 U352 ( .A1(n287), .A2(n320), .ZN(n[311]) );
  NR2D0 U353 ( .A1(n288), .A2(n320), .ZN(n[308]) );
  NR2D0 U354 ( .A1(n289), .A2(n320), .ZN(n[305]) );
  NR2D0 U355 ( .A1(n290), .A2(n320), .ZN(n[304]) );
  NR2D0 U356 ( .A1(n291), .A2(n320), .ZN(n[301]) );
  NR2D0 U357 ( .A1(n292), .A2(n320), .ZN(n[298]) );
  NR2D0 U358 ( .A1(n293), .A2(n320), .ZN(n[297]) );
  NR2D0 U359 ( .A1(n294), .A2(n320), .ZN(n[296]) );
  NR2D0 U360 ( .A1(n295), .A2(n320), .ZN(n[293]) );
  NR2D0 U361 ( .A1(n296), .A2(n320), .ZN(n[290]) );
  NR2D0 U362 ( .A1(n297), .A2(n320), .ZN(n[289]) );
  NR2D0 U363 ( .A1(n298), .A2(n320), .ZN(n[286]) );
  NR2D0 U364 ( .A1(n299), .A2(n320), .ZN(n[283]) );
  NR2D0 U365 ( .A1(n300), .A2(n320), .ZN(n[282]) );
  NR2D0 U366 ( .A1(n301), .A2(n320), .ZN(n[281]) );
  NR2D0 U367 ( .A1(n302), .A2(n320), .ZN(n[280]) );
  NR2D0 U368 ( .A1(n303), .A2(n320), .ZN(n[277]) );
  NR2D0 U369 ( .A1(n304), .A2(n320), .ZN(n[274]) );
  NR2D0 U370 ( .A1(n305), .A2(n320), .ZN(n[273]) );
  NR2D0 U371 ( .A1(n306), .A2(n320), .ZN(n[270]) );
  NR2D0 U372 ( .A1(n307), .A2(n320), .ZN(n[267]) );
  NR2D0 U373 ( .A1(n308), .A2(n320), .ZN(n[266]) );
  NR2D0 U374 ( .A1(n309), .A2(n320), .ZN(n[265]) );
  NR2D0 U375 ( .A1(n310), .A2(n320), .ZN(n[262]) );
  NR2D0 U376 ( .A1(n311), .A2(n320), .ZN(n[259]) );
  NR2D0 U377 ( .A1(n312), .A2(n320), .ZN(n[258]) );
  NR2D0 U378 ( .A1(n313), .A2(n320), .ZN(n[255]) );
  NR2D0 U379 ( .A1(n314), .A2(n320), .ZN(n[252]) );
  NR2D0 U380 ( .A1(n315), .A2(n320), .ZN(n[251]) );
  NR2D0 U381 ( .A1(n316), .A2(n320), .ZN(n[250]) );
  NR2D0 U382 ( .A1(n317), .A2(n320), .ZN(n[249]) );
  NR2D0 U383 ( .A1(n318), .A2(n320), .ZN(n[248]) );
  NR2D0 U384 ( .A1(n319), .A2(n320), .ZN(n[247]) );
  NR2D0 U385 ( .A1(n257), .A2(n320), .ZN(n[246]) );
  CKND0 U386 ( .I(n256), .ZN(n[243]) );
  CKND2D0 U387 ( .A1(b[5]), .A2(n[116]), .ZN(n256) );
  CKND0 U388 ( .I(n258), .ZN(n[240]) );
  CKND2D0 U389 ( .A1(n[113]), .A2(b[5]), .ZN(n258) );
  CKND0 U390 ( .I(n259), .ZN(n[239]) );
  CKND2D0 U391 ( .A1(n[112]), .A2(b[5]), .ZN(n259) );
  CKND0 U392 ( .I(n260), .ZN(n[236]) );
  CKND2D0 U393 ( .A1(n[109]), .A2(b[5]), .ZN(n260) );
  CKND0 U394 ( .I(n261), .ZN(n[233]) );
  CKND2D0 U395 ( .A1(n[106]), .A2(b[5]), .ZN(n261) );
  CKND0 U396 ( .I(n262), .ZN(n[232]) );
  CKND2D0 U397 ( .A1(n[105]), .A2(b[5]), .ZN(n262) );
  CKND0 U398 ( .I(n263), .ZN(n[231]) );
  CKND2D0 U399 ( .A1(n[104]), .A2(b[5]), .ZN(n263) );
  CKND0 U400 ( .I(n264), .ZN(n[228]) );
  CKND2D0 U401 ( .A1(n[101]), .A2(b[5]), .ZN(n264) );
  CKND0 U402 ( .I(n265), .ZN(n[225]) );
  CKND2D0 U403 ( .A1(n[98]), .A2(b[5]), .ZN(n265) );
  CKND0 U404 ( .I(n266), .ZN(n[224]) );
  CKND2D0 U405 ( .A1(n[97]), .A2(b[5]), .ZN(n266) );
  CKND0 U406 ( .I(n267), .ZN(n[221]) );
  CKND2D0 U407 ( .A1(n[94]), .A2(b[5]), .ZN(n267) );
  CKND0 U408 ( .I(n268), .ZN(n[218]) );
  CKND2D0 U409 ( .A1(n[91]), .A2(b[5]), .ZN(n268) );
  CKND0 U410 ( .I(n269), .ZN(n[217]) );
  CKND2D0 U411 ( .A1(n[90]), .A2(b[5]), .ZN(n269) );
  CKND0 U412 ( .I(n270), .ZN(n[216]) );
  CKND2D0 U413 ( .A1(n[89]), .A2(b[5]), .ZN(n270) );
  CKND0 U414 ( .I(n271), .ZN(n[215]) );
  CKND2D0 U415 ( .A1(n[88]), .A2(b[5]), .ZN(n271) );
  CKND0 U416 ( .I(n272), .ZN(n[212]) );
  CKND2D0 U417 ( .A1(n[85]), .A2(b[5]), .ZN(n272) );
  CKND0 U418 ( .I(n273), .ZN(n[209]) );
  CKND2D0 U419 ( .A1(n[82]), .A2(b[5]), .ZN(n273) );
  CKND0 U420 ( .I(n274), .ZN(n[208]) );
  CKND2D0 U421 ( .A1(n[81]), .A2(b[5]), .ZN(n274) );
  CKND0 U422 ( .I(n275), .ZN(n[205]) );
  CKND2D0 U423 ( .A1(n[78]), .A2(b[5]), .ZN(n275) );
  CKND0 U424 ( .I(n276), .ZN(n[202]) );
  CKND2D0 U425 ( .A1(n[75]), .A2(b[5]), .ZN(n276) );
  CKND0 U426 ( .I(n277), .ZN(n[201]) );
  CKND2D0 U427 ( .A1(n[74]), .A2(b[5]), .ZN(n277) );
  CKND0 U428 ( .I(n278), .ZN(n[200]) );
  CKND2D0 U429 ( .A1(n[73]), .A2(b[5]), .ZN(n278) );
  CKND0 U430 ( .I(n279), .ZN(n[197]) );
  CKND2D0 U431 ( .A1(n[70]), .A2(b[5]), .ZN(n279) );
  CKND0 U432 ( .I(n280), .ZN(n[194]) );
  CKND2D0 U433 ( .A1(n[67]), .A2(b[5]), .ZN(n280) );
  CKND0 U434 ( .I(n281), .ZN(n[193]) );
  CKND2D0 U435 ( .A1(n[66]), .A2(b[5]), .ZN(n281) );
  CKND0 U436 ( .I(n282), .ZN(n[190]) );
  CKND2D0 U437 ( .A1(n[63]), .A2(b[5]), .ZN(n282) );
  CKND0 U438 ( .I(n283), .ZN(n[187]) );
  CKND2D0 U439 ( .A1(n[60]), .A2(b[5]), .ZN(n283) );
  CKND0 U440 ( .I(n284), .ZN(n[186]) );
  CKND2D0 U441 ( .A1(n[59]), .A2(b[5]), .ZN(n284) );
  CKND0 U442 ( .I(n285), .ZN(n[185]) );
  CKND2D0 U443 ( .A1(n[58]), .A2(b[5]), .ZN(n285) );
  CKND0 U444 ( .I(n286), .ZN(n[184]) );
  CKND2D0 U445 ( .A1(n[57]), .A2(b[5]), .ZN(n286) );
  CKND0 U446 ( .I(n287), .ZN(n[183]) );
  CKND2D0 U447 ( .A1(n[56]), .A2(b[5]), .ZN(n287) );
  CKND0 U448 ( .I(n288), .ZN(n[180]) );
  CKND2D0 U449 ( .A1(a[5]), .A2(n[116]), .ZN(n288) );
  CKND0 U450 ( .I(n289), .ZN(n[177]) );
  CKND2D0 U451 ( .A1(a[5]), .A2(n[113]), .ZN(n289) );
  CKND0 U452 ( .I(n290), .ZN(n[176]) );
  CKND2D0 U453 ( .A1(a[5]), .A2(n[112]), .ZN(n290) );
  CKND0 U454 ( .I(n291), .ZN(n[173]) );
  CKND2D0 U455 ( .A1(a[5]), .A2(n[109]), .ZN(n291) );
  CKND0 U456 ( .I(n292), .ZN(n[170]) );
  CKND2D0 U457 ( .A1(a[5]), .A2(n[106]), .ZN(n292) );
  CKND0 U458 ( .I(n293), .ZN(n[169]) );
  CKND2D0 U459 ( .A1(a[5]), .A2(n[105]), .ZN(n293) );
  CKND0 U460 ( .I(n294), .ZN(n[168]) );
  CKND2D0 U461 ( .A1(a[5]), .A2(n[104]), .ZN(n294) );
  CKND0 U462 ( .I(n295), .ZN(n[165]) );
  CKND2D0 U463 ( .A1(a[5]), .A2(n[101]), .ZN(n295) );
  CKND0 U464 ( .I(n296), .ZN(n[162]) );
  CKND2D0 U465 ( .A1(a[5]), .A2(n[98]), .ZN(n296) );
  AN2D0 U466 ( .A1(b[4]), .A2(n[35]), .Z(n[98]) );
  CKND0 U467 ( .I(n297), .ZN(n[161]) );
  CKND2D0 U468 ( .A1(a[5]), .A2(n[97]), .ZN(n297) );
  AN2D0 U469 ( .A1(n[34]), .A2(b[4]), .Z(n[97]) );
  CKND0 U470 ( .I(n298), .ZN(n[158]) );
  CKND2D0 U471 ( .A1(a[5]), .A2(n[94]), .ZN(n298) );
  AN2D0 U472 ( .A1(n[31]), .A2(b[4]), .Z(n[94]) );
  CKND0 U473 ( .I(n299), .ZN(n[155]) );
  CKND2D0 U474 ( .A1(a[5]), .A2(n[91]), .ZN(n299) );
  AN2D0 U475 ( .A1(n[28]), .A2(b[4]), .Z(n[91]) );
  CKND0 U476 ( .I(n300), .ZN(n[154]) );
  CKND2D0 U477 ( .A1(a[5]), .A2(n[90]), .ZN(n300) );
  AN2D0 U478 ( .A1(n[27]), .A2(b[4]), .Z(n[90]) );
  CKND0 U479 ( .I(n301), .ZN(n[153]) );
  CKND2D0 U480 ( .A1(a[5]), .A2(n[89]), .ZN(n301) );
  AN2D0 U481 ( .A1(n[26]), .A2(b[4]), .Z(n[89]) );
  CKND0 U482 ( .I(n302), .ZN(n[152]) );
  CKND2D0 U483 ( .A1(a[5]), .A2(n[88]), .ZN(n302) );
  AN2D0 U484 ( .A1(n[25]), .A2(b[4]), .Z(n[88]) );
  CKND0 U485 ( .I(n303), .ZN(n[149]) );
  CKND2D0 U486 ( .A1(a[5]), .A2(n[85]), .ZN(n303) );
  AN2D0 U487 ( .A1(a[4]), .A2(n[53]), .Z(n[85]) );
  CKND0 U488 ( .I(n304), .ZN(n[146]) );
  CKND2D0 U489 ( .A1(a[5]), .A2(n[82]), .ZN(n304) );
  AN2D0 U490 ( .A1(n[50]), .A2(a[4]), .Z(n[82]) );
  CKND0 U491 ( .I(n305), .ZN(n[145]) );
  CKND2D0 U492 ( .A1(a[5]), .A2(n[81]), .ZN(n305) );
  AN2D0 U493 ( .A1(n[49]), .A2(a[4]), .Z(n[81]) );
  CKND0 U494 ( .I(n306), .ZN(n[142]) );
  CKND2D0 U495 ( .A1(a[5]), .A2(n[78]), .ZN(n306) );
  AN2D0 U496 ( .A1(n[46]), .A2(a[4]), .Z(n[78]) );
  CKND0 U497 ( .I(n307), .ZN(n[139]) );
  CKND2D0 U498 ( .A1(a[5]), .A2(n[75]), .ZN(n307) );
  AN2D0 U499 ( .A1(n[43]), .A2(a[4]), .Z(n[75]) );
  CKND0 U500 ( .I(n308), .ZN(n[138]) );
  CKND2D0 U501 ( .A1(a[5]), .A2(n[74]), .ZN(n308) );
  AN2D0 U502 ( .A1(n[42]), .A2(a[4]), .Z(n[74]) );
  CKND0 U503 ( .I(n309), .ZN(n[137]) );
  CKND2D0 U504 ( .A1(a[5]), .A2(n[73]), .ZN(n309) );
  AN2D0 U505 ( .A1(n[41]), .A2(a[4]), .Z(n[73]) );
  CKND0 U506 ( .I(n310), .ZN(n[134]) );
  CKND2D0 U507 ( .A1(a[5]), .A2(n[70]), .ZN(n310) );
  AN2D0 U508 ( .A1(n[38]), .A2(a[4]), .Z(n[70]) );
  CKND0 U509 ( .I(n311), .ZN(n[131]) );
  CKND2D0 U510 ( .A1(a[5]), .A2(n[67]), .ZN(n311) );
  AN2D0 U511 ( .A1(a[4]), .A2(n[35]), .Z(n[67]) );
  AN2D0 U512 ( .A1(a[3]), .A2(n[19]), .Z(n[35]) );
  CKND0 U513 ( .I(n312), .ZN(n[130]) );
  CKND2D0 U514 ( .A1(a[5]), .A2(n[66]), .ZN(n312) );
  AN2D0 U515 ( .A1(a[4]), .A2(n[34]), .Z(n[66]) );
  AN2D0 U516 ( .A1(n[18]), .A2(a[3]), .Z(n[34]) );
  CKND0 U517 ( .I(n313), .ZN(n[127]) );
  CKND2D0 U518 ( .A1(a[5]), .A2(n[63]), .ZN(n313) );
  AN2D0 U519 ( .A1(a[4]), .A2(n[31]), .Z(n[63]) );
  AN2D0 U520 ( .A1(n[15]), .A2(a[3]), .Z(n[31]) );
  CKND0 U521 ( .I(n314), .ZN(n[124]) );
  CKND2D0 U522 ( .A1(a[5]), .A2(n[60]), .ZN(n314) );
  AN2D0 U523 ( .A1(a[4]), .A2(n[28]), .Z(n[60]) );
  AN2D0 U524 ( .A1(n[12]), .A2(a[3]), .Z(n[28]) );
  CKND0 U525 ( .I(n315), .ZN(n[123]) );
  CKND2D0 U526 ( .A1(a[5]), .A2(n[59]), .ZN(n315) );
  AN2D0 U527 ( .A1(a[4]), .A2(n[27]), .Z(n[59]) );
  AN2D0 U528 ( .A1(n[11]), .A2(a[3]), .Z(n[27]) );
  CKND0 U529 ( .I(n316), .ZN(n[122]) );
  CKND2D0 U530 ( .A1(a[5]), .A2(n[58]), .ZN(n316) );
  AN2D0 U531 ( .A1(a[4]), .A2(n[26]), .Z(n[58]) );
  AN2D0 U532 ( .A1(n[10]), .A2(a[3]), .Z(n[26]) );
  CKND0 U533 ( .I(n317), .ZN(n[121]) );
  CKND2D0 U534 ( .A1(a[5]), .A2(n[57]), .ZN(n317) );
  AN2D0 U535 ( .A1(a[4]), .A2(n[25]), .Z(n[57]) );
  AN2D0 U536 ( .A1(b[3]), .A2(a[3]), .Z(n[25]) );
  CKND0 U537 ( .I(n318), .ZN(n[120]) );
  CKND2D0 U538 ( .A1(a[5]), .A2(n[56]), .ZN(n318) );
  AN2D0 U539 ( .A1(a[4]), .A2(b[4]), .Z(n[56]) );
  CKND0 U540 ( .I(n319), .ZN(n[119]) );
  CKND2D0 U541 ( .A1(a[5]), .A2(b[5]), .ZN(n319) );
  AN2D0 U542 ( .A1(n[53]), .A2(b[4]), .Z(n[116]) );
  AN2D0 U543 ( .A1(n[22]), .A2(b[3]), .Z(n[53]) );
  AN2D0 U544 ( .A1(n[50]), .A2(b[4]), .Z(n[113]) );
  AN2D0 U545 ( .A1(b[3]), .A2(n[19]), .Z(n[50]) );
  AN2D0 U546 ( .A1(b[2]), .A2(n[4]), .Z(n[19]) );
  AN2D0 U547 ( .A1(n[49]), .A2(b[4]), .Z(n[112]) );
  AN2D0 U548 ( .A1(b[3]), .A2(n[18]), .Z(n[49]) );
  AN2D0 U549 ( .A1(n[3]), .A2(b[2]), .Z(n[18]) );
  AN2D0 U550 ( .A1(n[46]), .A2(b[4]), .Z(n[109]) );
  AN2D0 U551 ( .A1(b[3]), .A2(n[15]), .Z(n[46]) );
  AN2D0 U552 ( .A1(a[2]), .A2(n[7]), .Z(n[15]) );
  AN2D0 U553 ( .A1(n[43]), .A2(b[4]), .Z(n[106]) );
  AN2D0 U554 ( .A1(b[3]), .A2(n[12]), .Z(n[43]) );
  AN2D0 U555 ( .A1(a[2]), .A2(n[4]), .Z(n[12]) );
  AN2D0 U556 ( .A1(a[1]), .A2(n[0]), .Z(n[4]) );
  AN2D0 U557 ( .A1(n[42]), .A2(b[4]), .Z(n[105]) );
  AN2D0 U558 ( .A1(b[3]), .A2(n[11]), .Z(n[42]) );
  AN2D0 U559 ( .A1(a[2]), .A2(n[3]), .Z(n[11]) );
  AN2D0 U560 ( .A1(b[1]), .A2(a[1]), .Z(n[3]) );
  AN2D0 U561 ( .A1(n[41]), .A2(b[4]), .Z(n[104]) );
  AN2D0 U562 ( .A1(b[3]), .A2(n[10]), .Z(n[41]) );
  AN2D0 U563 ( .A1(a[2]), .A2(b[2]), .Z(n[10]) );
  AN2D0 U564 ( .A1(n[38]), .A2(b[4]), .Z(n[101]) );
  AN2D0 U565 ( .A1(n[22]), .A2(a[3]), .Z(n[38]) );
  AN2D0 U566 ( .A1(n[7]), .A2(b[2]), .Z(n[22]) );
  AN2D0 U567 ( .A1(b[1]), .A2(n[0]), .Z(n[7]) );
  AN2D0 U568 ( .A1(b[0]), .A2(a[0]), .Z(n[0]) );
endmodule


module gen_cla_decomposed ( a, b, s );
  input [7:0] a;
  input [7:0] b;
  output [7:0] s;
  wire   n1;
  wire   [500:0] n;

  gen_nonlinear_part NLIN ( .a(a), .b(b), .n(n) );
  gen_linear_part LIN ( .a(a), .b(b), .n({n1, n1, n[498], n1, n1, n[495:494], 
        n1, n1, n[491], n1, n1, n[488:486], n1, n1, n[483], n1, n1, n[480:479], 
        n1, n1, n[476], n1, n1, n[473:470], n1, n1, n[467], n1, n1, n[464:463], 
        n1, n1, n[460], n1, n1, n[457:455], n1, n1, n[452], n1, n1, n[449:448], 
        n1, n1, n[445], n1, n1, n[442:438], n1, n1, n[435], n1, n1, n[432:431], 
        n1, n1, n[428], n1, n1, n[425:423], n1, n1, n[420], n1, n1, n[417:416], 
        n1, n1, n[413], n1, n1, n[410:407], n1, n1, n[404], n1, n1, n[401:400], 
        n1, n1, n[397], n1, n1, n[394:392], n1, n1, n[389], n1, n1, n[386:385], 
        n1, n1, n[382], n1, n1, n[379:374], n1, n1, n[371], n1, n1, n[368:367], 
        n1, n1, n[364], n1, n1, n[361:359], n1, n1, n[356], n1, n1, n[353:352], 
        n1, n1, n[349], n1, n1, n[346:343], n1, n1, n[340], n1, n1, n[337:336], 
        n1, n1, n[333], n1, n1, n[330:328], n1, n1, n[325], n1, n1, n[322:321], 
        n1, n1, n[318], n1, n1, n[315:311], n1, n1, n[308], n1, n1, n[305:304], 
        n1, n1, n[301], n1, n1, n[298:296], n1, n1, n[293], n1, n1, n[290:289], 
        n1, n1, n[286], n1, n1, n[283:280], n1, n1, n[277], n1, n1, n[274:273], 
        n1, n1, n[270], n1, n1, n[267:265], n1, n1, n[262], n1, n1, n[259:258], 
        n1, n1, n[255], n1, n1, n[252:246], n1, n1, n[243], n1, n1, n[240:239], 
        n1, n1, n[236], n1, n1, n[233:231], n1, n1, n[228], n1, n1, n[225:224], 
        n1, n1, n[221], n1, n1, n[218:215], n1, n1, n[212], n1, n1, n[209:208], 
        n1, n1, n[205], n1, n1, n[202:200], n1, n1, n[197], n1, n1, n[194:193], 
        n1, n1, n[190], n1, n1, n[187:183], n1, n1, n[180], n1, n1, n[177:176], 
        n1, n1, n[173], n1, n1, n[170:168], n1, n1, n[165], n1, n1, n[162:161], 
        n1, n1, n[158], n1, n1, n[155:152], n1, n1, n[149], n1, n1, n[146:145], 
        n1, n1, n[142], n1, n1, n[139:137], n1, n1, n[134], n1, n1, n[131:130], 
        n1, n1, n[127], n1, n1, n[124:119], n1, n1, n[116], n1, n1, n[113:112], 
        n1, n1, n[109], n1, n1, n[106:104], n1, n1, n[101], n1, n1, n[98:97], 
        n1, n1, n[94], n1, n1, n[91:88], n1, n1, n[85], n1, n1, n[82:81], n1, 
        n1, n[78], n1, n1, n[75:73], n1, n1, n[70], n1, n1, n[67:66], n1, n1, 
        n[63], n1, n1, n[60:56], n1, n1, n[53], n1, n1, n[50:49], n1, n1, 
        n[46], n1, n1, n[43:41], n1, n1, n[38], n1, n1, n[35:34], n1, n1, 
        n[31], n1, n1, n[28:25], n1, n1, n[22], n1, n1, n[19:18], n1, n1, 
        n[15], n1, n1, n[12:10], n1, n1, n[7], n1, n1, n[4:3], n1, n1, n[0]}), 
        .s(s) );
  TIEL U1 ( .ZN(n1) );
endmodule

