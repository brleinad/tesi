//Inlcude file for the global parameters

//'ifndef _glogals_vh
//'define _globals_vh

'define N 128

//'endif

