
module cla_adder ( a, b, s, cin, cout );
  input [127:0] a;
  input [127:0] b;
  output [127:0] s;
  input cin;
  output cout;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126;
  wire   [126:0] g;
  wire   [127:0] p;
  wire   [127:1] c;

  XOR2D0 C1154 ( .A1(p[0]), .A2(cin), .Z(s[0]) );
  XOR2D0 C1153 ( .A1(p[1]), .A2(c[1]), .Z(s[1]) );
  XOR2D0 C1152 ( .A1(p[2]), .A2(c[2]), .Z(s[2]) );
  XOR2D0 C1151 ( .A1(p[3]), .A2(c[3]), .Z(s[3]) );
  XOR2D0 C1150 ( .A1(p[4]), .A2(c[4]), .Z(s[4]) );
  XOR2D0 C1149 ( .A1(p[5]), .A2(c[5]), .Z(s[5]) );
  XOR2D0 C1148 ( .A1(p[6]), .A2(c[6]), .Z(s[6]) );
  XOR2D0 C1147 ( .A1(p[7]), .A2(c[7]), .Z(s[7]) );
  XOR2D0 C1146 ( .A1(p[8]), .A2(c[8]), .Z(s[8]) );
  XOR2D0 C1145 ( .A1(p[9]), .A2(c[9]), .Z(s[9]) );
  XOR2D0 C1144 ( .A1(p[10]), .A2(c[10]), .Z(s[10]) );
  XOR2D0 C1143 ( .A1(p[11]), .A2(c[11]), .Z(s[11]) );
  XOR2D0 C1142 ( .A1(p[12]), .A2(c[12]), .Z(s[12]) );
  XOR2D0 C1141 ( .A1(p[13]), .A2(c[13]), .Z(s[13]) );
  XOR2D0 C1140 ( .A1(p[14]), .A2(c[14]), .Z(s[14]) );
  XOR2D0 C1139 ( .A1(p[15]), .A2(c[15]), .Z(s[15]) );
  XOR2D0 C1138 ( .A1(p[16]), .A2(c[16]), .Z(s[16]) );
  XOR2D0 C1137 ( .A1(p[17]), .A2(c[17]), .Z(s[17]) );
  XOR2D0 C1136 ( .A1(p[18]), .A2(c[18]), .Z(s[18]) );
  XOR2D0 C1135 ( .A1(p[19]), .A2(c[19]), .Z(s[19]) );
  XOR2D0 C1134 ( .A1(p[20]), .A2(c[20]), .Z(s[20]) );
  XOR2D0 C1133 ( .A1(p[21]), .A2(c[21]), .Z(s[21]) );
  XOR2D0 C1132 ( .A1(p[22]), .A2(c[22]), .Z(s[22]) );
  XOR2D0 C1131 ( .A1(p[23]), .A2(c[23]), .Z(s[23]) );
  XOR2D0 C1130 ( .A1(p[24]), .A2(c[24]), .Z(s[24]) );
  XOR2D0 C1129 ( .A1(p[25]), .A2(c[25]), .Z(s[25]) );
  XOR2D0 C1128 ( .A1(p[26]), .A2(c[26]), .Z(s[26]) );
  XOR2D0 C1127 ( .A1(p[27]), .A2(c[27]), .Z(s[27]) );
  XOR2D0 C1126 ( .A1(p[28]), .A2(c[28]), .Z(s[28]) );
  XOR2D0 C1125 ( .A1(p[29]), .A2(c[29]), .Z(s[29]) );
  XOR2D0 C1124 ( .A1(p[30]), .A2(c[30]), .Z(s[30]) );
  XOR2D0 C1123 ( .A1(p[31]), .A2(c[31]), .Z(s[31]) );
  XOR2D0 C1122 ( .A1(p[32]), .A2(c[32]), .Z(s[32]) );
  XOR2D0 C1121 ( .A1(p[33]), .A2(c[33]), .Z(s[33]) );
  XOR2D0 C1120 ( .A1(p[34]), .A2(c[34]), .Z(s[34]) );
  XOR2D0 C1119 ( .A1(p[35]), .A2(c[35]), .Z(s[35]) );
  XOR2D0 C1118 ( .A1(p[36]), .A2(c[36]), .Z(s[36]) );
  XOR2D0 C1117 ( .A1(p[37]), .A2(c[37]), .Z(s[37]) );
  XOR2D0 C1116 ( .A1(p[38]), .A2(c[38]), .Z(s[38]) );
  XOR2D0 C1115 ( .A1(p[39]), .A2(c[39]), .Z(s[39]) );
  XOR2D0 C1114 ( .A1(p[40]), .A2(c[40]), .Z(s[40]) );
  XOR2D0 C1113 ( .A1(p[41]), .A2(c[41]), .Z(s[41]) );
  XOR2D0 C1112 ( .A1(p[42]), .A2(c[42]), .Z(s[42]) );
  XOR2D0 C1111 ( .A1(p[43]), .A2(c[43]), .Z(s[43]) );
  XOR2D0 C1110 ( .A1(p[44]), .A2(c[44]), .Z(s[44]) );
  XOR2D0 C1109 ( .A1(p[45]), .A2(c[45]), .Z(s[45]) );
  XOR2D0 C1108 ( .A1(p[46]), .A2(c[46]), .Z(s[46]) );
  XOR2D0 C1107 ( .A1(p[47]), .A2(c[47]), .Z(s[47]) );
  XOR2D0 C1106 ( .A1(p[48]), .A2(c[48]), .Z(s[48]) );
  XOR2D0 C1105 ( .A1(p[49]), .A2(c[49]), .Z(s[49]) );
  XOR2D0 C1104 ( .A1(p[50]), .A2(c[50]), .Z(s[50]) );
  XOR2D0 C1103 ( .A1(p[51]), .A2(c[51]), .Z(s[51]) );
  XOR2D0 C1102 ( .A1(p[52]), .A2(c[52]), .Z(s[52]) );
  XOR2D0 C1101 ( .A1(p[53]), .A2(c[53]), .Z(s[53]) );
  XOR2D0 C1100 ( .A1(p[54]), .A2(c[54]), .Z(s[54]) );
  XOR2D0 C1099 ( .A1(p[55]), .A2(c[55]), .Z(s[55]) );
  XOR2D0 C1098 ( .A1(p[56]), .A2(c[56]), .Z(s[56]) );
  XOR2D0 C1097 ( .A1(p[57]), .A2(c[57]), .Z(s[57]) );
  XOR2D0 C1096 ( .A1(p[58]), .A2(c[58]), .Z(s[58]) );
  XOR2D0 C1095 ( .A1(p[59]), .A2(c[59]), .Z(s[59]) );
  XOR2D0 C1094 ( .A1(p[60]), .A2(c[60]), .Z(s[60]) );
  XOR2D0 C1093 ( .A1(p[61]), .A2(c[61]), .Z(s[61]) );
  XOR2D0 C1092 ( .A1(p[62]), .A2(c[62]), .Z(s[62]) );
  XOR2D0 C1091 ( .A1(p[63]), .A2(c[63]), .Z(s[63]) );
  XOR2D0 C1090 ( .A1(p[64]), .A2(c[64]), .Z(s[64]) );
  XOR2D0 C1089 ( .A1(p[65]), .A2(c[65]), .Z(s[65]) );
  XOR2D0 C1088 ( .A1(p[66]), .A2(c[66]), .Z(s[66]) );
  XOR2D0 C1087 ( .A1(p[67]), .A2(c[67]), .Z(s[67]) );
  XOR2D0 C1086 ( .A1(p[68]), .A2(c[68]), .Z(s[68]) );
  XOR2D0 C1085 ( .A1(p[69]), .A2(c[69]), .Z(s[69]) );
  XOR2D0 C1084 ( .A1(p[70]), .A2(c[70]), .Z(s[70]) );
  XOR2D0 C1083 ( .A1(p[71]), .A2(c[71]), .Z(s[71]) );
  XOR2D0 C1082 ( .A1(p[72]), .A2(c[72]), .Z(s[72]) );
  XOR2D0 C1081 ( .A1(p[73]), .A2(c[73]), .Z(s[73]) );
  XOR2D0 C1080 ( .A1(p[74]), .A2(c[74]), .Z(s[74]) );
  XOR2D0 C1079 ( .A1(p[75]), .A2(c[75]), .Z(s[75]) );
  XOR2D0 C1078 ( .A1(p[76]), .A2(c[76]), .Z(s[76]) );
  XOR2D0 C1077 ( .A1(p[77]), .A2(c[77]), .Z(s[77]) );
  XOR2D0 C1076 ( .A1(p[78]), .A2(c[78]), .Z(s[78]) );
  XOR2D0 C1075 ( .A1(p[79]), .A2(c[79]), .Z(s[79]) );
  XOR2D0 C1074 ( .A1(p[80]), .A2(c[80]), .Z(s[80]) );
  XOR2D0 C1073 ( .A1(p[81]), .A2(c[81]), .Z(s[81]) );
  XOR2D0 C1072 ( .A1(p[82]), .A2(c[82]), .Z(s[82]) );
  XOR2D0 C1071 ( .A1(p[83]), .A2(c[83]), .Z(s[83]) );
  XOR2D0 C1070 ( .A1(p[84]), .A2(c[84]), .Z(s[84]) );
  XOR2D0 C1069 ( .A1(p[85]), .A2(c[85]), .Z(s[85]) );
  XOR2D0 C1068 ( .A1(p[86]), .A2(c[86]), .Z(s[86]) );
  XOR2D0 C1067 ( .A1(p[87]), .A2(c[87]), .Z(s[87]) );
  XOR2D0 C1066 ( .A1(p[88]), .A2(c[88]), .Z(s[88]) );
  XOR2D0 C1065 ( .A1(p[89]), .A2(c[89]), .Z(s[89]) );
  XOR2D0 C1064 ( .A1(p[90]), .A2(c[90]), .Z(s[90]) );
  XOR2D0 C1063 ( .A1(p[91]), .A2(c[91]), .Z(s[91]) );
  XOR2D0 C1062 ( .A1(p[92]), .A2(c[92]), .Z(s[92]) );
  XOR2D0 C1061 ( .A1(p[93]), .A2(c[93]), .Z(s[93]) );
  XOR2D0 C1060 ( .A1(p[94]), .A2(c[94]), .Z(s[94]) );
  XOR2D0 C1059 ( .A1(p[95]), .A2(c[95]), .Z(s[95]) );
  XOR2D0 C1058 ( .A1(p[96]), .A2(c[96]), .Z(s[96]) );
  XOR2D0 C1057 ( .A1(p[97]), .A2(c[97]), .Z(s[97]) );
  XOR2D0 C1056 ( .A1(p[98]), .A2(c[98]), .Z(s[98]) );
  XOR2D0 C1055 ( .A1(p[99]), .A2(c[99]), .Z(s[99]) );
  XOR2D0 C1054 ( .A1(p[100]), .A2(c[100]), .Z(s[100]) );
  XOR2D0 C1053 ( .A1(p[101]), .A2(c[101]), .Z(s[101]) );
  XOR2D0 C1052 ( .A1(p[102]), .A2(c[102]), .Z(s[102]) );
  XOR2D0 C1051 ( .A1(p[103]), .A2(c[103]), .Z(s[103]) );
  XOR2D0 C1050 ( .A1(p[104]), .A2(c[104]), .Z(s[104]) );
  XOR2D0 C1049 ( .A1(p[105]), .A2(c[105]), .Z(s[105]) );
  XOR2D0 C1048 ( .A1(p[106]), .A2(c[106]), .Z(s[106]) );
  XOR2D0 C1047 ( .A1(p[107]), .A2(c[107]), .Z(s[107]) );
  XOR2D0 C1046 ( .A1(p[108]), .A2(c[108]), .Z(s[108]) );
  XOR2D0 C1045 ( .A1(p[109]), .A2(c[109]), .Z(s[109]) );
  XOR2D0 C1044 ( .A1(p[110]), .A2(c[110]), .Z(s[110]) );
  XOR2D0 C1043 ( .A1(p[111]), .A2(c[111]), .Z(s[111]) );
  XOR2D0 C1042 ( .A1(p[112]), .A2(c[112]), .Z(s[112]) );
  XOR2D0 C1041 ( .A1(p[113]), .A2(c[113]), .Z(s[113]) );
  XOR2D0 C1040 ( .A1(p[114]), .A2(c[114]), .Z(s[114]) );
  XOR2D0 C1039 ( .A1(p[115]), .A2(c[115]), .Z(s[115]) );
  XOR2D0 C1038 ( .A1(p[116]), .A2(c[116]), .Z(s[116]) );
  XOR2D0 C1037 ( .A1(p[117]), .A2(c[117]), .Z(s[117]) );
  XOR2D0 C1036 ( .A1(p[118]), .A2(c[118]), .Z(s[118]) );
  XOR2D0 C1035 ( .A1(p[119]), .A2(c[119]), .Z(s[119]) );
  XOR2D0 C1034 ( .A1(p[120]), .A2(c[120]), .Z(s[120]) );
  XOR2D0 C1033 ( .A1(p[121]), .A2(c[121]), .Z(s[121]) );
  XOR2D0 C1032 ( .A1(p[122]), .A2(c[122]), .Z(s[122]) );
  XOR2D0 C1031 ( .A1(p[123]), .A2(c[123]), .Z(s[123]) );
  XOR2D0 C1030 ( .A1(p[124]), .A2(c[124]), .Z(s[124]) );
  XOR2D0 C1029 ( .A1(p[125]), .A2(c[125]), .Z(s[125]) );
  XOR2D0 C1028 ( .A1(p[126]), .A2(c[126]), .Z(s[126]) );
  XOR2D0 C1027 ( .A1(p[127]), .A2(c[127]), .Z(s[127]) );
  AN2D0 C1026 ( .A1(p[126]), .A2(c[126]), .Z(N126) );
  OR2D0 C1025 ( .A1(g[126]), .A2(N126), .Z(c[127]) );
  AN2D0 C1024 ( .A1(p[125]), .A2(c[125]), .Z(N125) );
  OR2D0 C1023 ( .A1(g[125]), .A2(N125), .Z(c[126]) );
  AN2D0 C1022 ( .A1(p[124]), .A2(c[124]), .Z(N124) );
  OR2D0 C1021 ( .A1(g[124]), .A2(N124), .Z(c[125]) );
  AN2D0 C1020 ( .A1(p[123]), .A2(c[123]), .Z(N123) );
  OR2D0 C1019 ( .A1(g[123]), .A2(N123), .Z(c[124]) );
  AN2D0 C1018 ( .A1(p[122]), .A2(c[122]), .Z(N122) );
  OR2D0 C1017 ( .A1(g[122]), .A2(N122), .Z(c[123]) );
  AN2D0 C1016 ( .A1(p[121]), .A2(c[121]), .Z(N121) );
  OR2D0 C1015 ( .A1(g[121]), .A2(N121), .Z(c[122]) );
  AN2D0 C1014 ( .A1(p[120]), .A2(c[120]), .Z(N120) );
  OR2D0 C1013 ( .A1(g[120]), .A2(N120), .Z(c[121]) );
  AN2D0 C1012 ( .A1(p[119]), .A2(c[119]), .Z(N119) );
  OR2D0 C1011 ( .A1(g[119]), .A2(N119), .Z(c[120]) );
  AN2D0 C1010 ( .A1(p[118]), .A2(c[118]), .Z(N118) );
  OR2D0 C1009 ( .A1(g[118]), .A2(N118), .Z(c[119]) );
  AN2D0 C1008 ( .A1(p[117]), .A2(c[117]), .Z(N117) );
  OR2D0 C1007 ( .A1(g[117]), .A2(N117), .Z(c[118]) );
  AN2D0 C1006 ( .A1(p[116]), .A2(c[116]), .Z(N116) );
  OR2D0 C1005 ( .A1(g[116]), .A2(N116), .Z(c[117]) );
  AN2D0 C1004 ( .A1(p[115]), .A2(c[115]), .Z(N115) );
  OR2D0 C1003 ( .A1(g[115]), .A2(N115), .Z(c[116]) );
  AN2D0 C1002 ( .A1(p[114]), .A2(c[114]), .Z(N114) );
  OR2D0 C1001 ( .A1(g[114]), .A2(N114), .Z(c[115]) );
  AN2D0 C1000 ( .A1(p[113]), .A2(c[113]), .Z(N113) );
  OR2D0 C999 ( .A1(g[113]), .A2(N113), .Z(c[114]) );
  AN2D0 C998 ( .A1(p[112]), .A2(c[112]), .Z(N112) );
  OR2D0 C997 ( .A1(g[112]), .A2(N112), .Z(c[113]) );
  AN2D0 C996 ( .A1(p[111]), .A2(c[111]), .Z(N111) );
  OR2D0 C995 ( .A1(g[111]), .A2(N111), .Z(c[112]) );
  AN2D0 C994 ( .A1(p[110]), .A2(c[110]), .Z(N110) );
  OR2D0 C993 ( .A1(g[110]), .A2(N110), .Z(c[111]) );
  AN2D0 C992 ( .A1(p[109]), .A2(c[109]), .Z(N109) );
  OR2D0 C991 ( .A1(g[109]), .A2(N109), .Z(c[110]) );
  AN2D0 C990 ( .A1(p[108]), .A2(c[108]), .Z(N108) );
  OR2D0 C989 ( .A1(g[108]), .A2(N108), .Z(c[109]) );
  AN2D0 C988 ( .A1(p[107]), .A2(c[107]), .Z(N107) );
  OR2D0 C987 ( .A1(g[107]), .A2(N107), .Z(c[108]) );
  AN2D0 C986 ( .A1(p[106]), .A2(c[106]), .Z(N106) );
  OR2D0 C985 ( .A1(g[106]), .A2(N106), .Z(c[107]) );
  AN2D0 C984 ( .A1(p[105]), .A2(c[105]), .Z(N105) );
  OR2D0 C983 ( .A1(g[105]), .A2(N105), .Z(c[106]) );
  AN2D0 C982 ( .A1(p[104]), .A2(c[104]), .Z(N104) );
  OR2D0 C981 ( .A1(g[104]), .A2(N104), .Z(c[105]) );
  AN2D0 C980 ( .A1(p[103]), .A2(c[103]), .Z(N103) );
  OR2D0 C979 ( .A1(g[103]), .A2(N103), .Z(c[104]) );
  AN2D0 C978 ( .A1(p[102]), .A2(c[102]), .Z(N102) );
  OR2D0 C977 ( .A1(g[102]), .A2(N102), .Z(c[103]) );
  AN2D0 C976 ( .A1(p[101]), .A2(c[101]), .Z(N101) );
  OR2D0 C975 ( .A1(g[101]), .A2(N101), .Z(c[102]) );
  AN2D0 C974 ( .A1(p[100]), .A2(c[100]), .Z(N100) );
  OR2D0 C973 ( .A1(g[100]), .A2(N100), .Z(c[101]) );
  AN2D0 C972 ( .A1(p[99]), .A2(c[99]), .Z(N99) );
  OR2D0 C971 ( .A1(g[99]), .A2(N99), .Z(c[100]) );
  AN2D0 C970 ( .A1(p[98]), .A2(c[98]), .Z(N98) );
  OR2D0 C969 ( .A1(g[98]), .A2(N98), .Z(c[99]) );
  AN2D0 C968 ( .A1(p[97]), .A2(c[97]), .Z(N97) );
  OR2D0 C967 ( .A1(g[97]), .A2(N97), .Z(c[98]) );
  AN2D0 C966 ( .A1(p[96]), .A2(c[96]), .Z(N96) );
  OR2D0 C965 ( .A1(g[96]), .A2(N96), .Z(c[97]) );
  AN2D0 C964 ( .A1(p[95]), .A2(c[95]), .Z(N95) );
  OR2D0 C963 ( .A1(g[95]), .A2(N95), .Z(c[96]) );
  AN2D0 C962 ( .A1(p[94]), .A2(c[94]), .Z(N94) );
  OR2D0 C961 ( .A1(g[94]), .A2(N94), .Z(c[95]) );
  AN2D0 C960 ( .A1(p[93]), .A2(c[93]), .Z(N93) );
  OR2D0 C959 ( .A1(g[93]), .A2(N93), .Z(c[94]) );
  AN2D0 C958 ( .A1(p[92]), .A2(c[92]), .Z(N92) );
  OR2D0 C957 ( .A1(g[92]), .A2(N92), .Z(c[93]) );
  AN2D0 C956 ( .A1(p[91]), .A2(c[91]), .Z(N91) );
  OR2D0 C955 ( .A1(g[91]), .A2(N91), .Z(c[92]) );
  AN2D0 C954 ( .A1(p[90]), .A2(c[90]), .Z(N90) );
  OR2D0 C953 ( .A1(g[90]), .A2(N90), .Z(c[91]) );
  AN2D0 C952 ( .A1(p[89]), .A2(c[89]), .Z(N89) );
  OR2D0 C951 ( .A1(g[89]), .A2(N89), .Z(c[90]) );
  AN2D0 C950 ( .A1(p[88]), .A2(c[88]), .Z(N88) );
  OR2D0 C949 ( .A1(g[88]), .A2(N88), .Z(c[89]) );
  AN2D0 C948 ( .A1(p[87]), .A2(c[87]), .Z(N87) );
  OR2D0 C947 ( .A1(g[87]), .A2(N87), .Z(c[88]) );
  AN2D0 C946 ( .A1(p[86]), .A2(c[86]), .Z(N86) );
  OR2D0 C945 ( .A1(g[86]), .A2(N86), .Z(c[87]) );
  AN2D0 C944 ( .A1(p[85]), .A2(c[85]), .Z(N85) );
  OR2D0 C943 ( .A1(g[85]), .A2(N85), .Z(c[86]) );
  AN2D0 C942 ( .A1(p[84]), .A2(c[84]), .Z(N84) );
  OR2D0 C941 ( .A1(g[84]), .A2(N84), .Z(c[85]) );
  AN2D0 C940 ( .A1(p[83]), .A2(c[83]), .Z(N83) );
  OR2D0 C939 ( .A1(g[83]), .A2(N83), .Z(c[84]) );
  AN2D0 C938 ( .A1(p[82]), .A2(c[82]), .Z(N82) );
  OR2D0 C937 ( .A1(g[82]), .A2(N82), .Z(c[83]) );
  AN2D0 C936 ( .A1(p[81]), .A2(c[81]), .Z(N81) );
  OR2D0 C935 ( .A1(g[81]), .A2(N81), .Z(c[82]) );
  AN2D0 C934 ( .A1(p[80]), .A2(c[80]), .Z(N80) );
  OR2D0 C933 ( .A1(g[80]), .A2(N80), .Z(c[81]) );
  AN2D0 C932 ( .A1(p[79]), .A2(c[79]), .Z(N79) );
  OR2D0 C931 ( .A1(g[79]), .A2(N79), .Z(c[80]) );
  AN2D0 C930 ( .A1(p[78]), .A2(c[78]), .Z(N78) );
  OR2D0 C929 ( .A1(g[78]), .A2(N78), .Z(c[79]) );
  AN2D0 C928 ( .A1(p[77]), .A2(c[77]), .Z(N77) );
  OR2D0 C927 ( .A1(g[77]), .A2(N77), .Z(c[78]) );
  AN2D0 C926 ( .A1(p[76]), .A2(c[76]), .Z(N76) );
  OR2D0 C925 ( .A1(g[76]), .A2(N76), .Z(c[77]) );
  AN2D0 C924 ( .A1(p[75]), .A2(c[75]), .Z(N75) );
  OR2D0 C923 ( .A1(g[75]), .A2(N75), .Z(c[76]) );
  AN2D0 C922 ( .A1(p[74]), .A2(c[74]), .Z(N74) );
  OR2D0 C921 ( .A1(g[74]), .A2(N74), .Z(c[75]) );
  AN2D0 C920 ( .A1(p[73]), .A2(c[73]), .Z(N73) );
  OR2D0 C919 ( .A1(g[73]), .A2(N73), .Z(c[74]) );
  AN2D0 C918 ( .A1(p[72]), .A2(c[72]), .Z(N72) );
  OR2D0 C917 ( .A1(g[72]), .A2(N72), .Z(c[73]) );
  AN2D0 C916 ( .A1(p[71]), .A2(c[71]), .Z(N71) );
  OR2D0 C915 ( .A1(g[71]), .A2(N71), .Z(c[72]) );
  AN2D0 C914 ( .A1(p[70]), .A2(c[70]), .Z(N70) );
  OR2D0 C913 ( .A1(g[70]), .A2(N70), .Z(c[71]) );
  AN2D0 C912 ( .A1(p[69]), .A2(c[69]), .Z(N69) );
  OR2D0 C911 ( .A1(g[69]), .A2(N69), .Z(c[70]) );
  AN2D0 C910 ( .A1(p[68]), .A2(c[68]), .Z(N68) );
  OR2D0 C909 ( .A1(g[68]), .A2(N68), .Z(c[69]) );
  AN2D0 C908 ( .A1(p[67]), .A2(c[67]), .Z(N67) );
  OR2D0 C907 ( .A1(g[67]), .A2(N67), .Z(c[68]) );
  AN2D0 C906 ( .A1(p[66]), .A2(c[66]), .Z(N66) );
  OR2D0 C905 ( .A1(g[66]), .A2(N66), .Z(c[67]) );
  AN2D0 C904 ( .A1(p[65]), .A2(c[65]), .Z(N65) );
  OR2D0 C903 ( .A1(g[65]), .A2(N65), .Z(c[66]) );
  AN2D0 C902 ( .A1(p[64]), .A2(c[64]), .Z(N64) );
  OR2D0 C901 ( .A1(g[64]), .A2(N64), .Z(c[65]) );
  AN2D0 C900 ( .A1(p[63]), .A2(c[63]), .Z(N63) );
  OR2D0 C899 ( .A1(g[63]), .A2(N63), .Z(c[64]) );
  AN2D0 C898 ( .A1(p[62]), .A2(c[62]), .Z(N62) );
  OR2D0 C897 ( .A1(g[62]), .A2(N62), .Z(c[63]) );
  AN2D0 C896 ( .A1(p[61]), .A2(c[61]), .Z(N61) );
  OR2D0 C895 ( .A1(g[61]), .A2(N61), .Z(c[62]) );
  AN2D0 C894 ( .A1(p[60]), .A2(c[60]), .Z(N60) );
  OR2D0 C893 ( .A1(g[60]), .A2(N60), .Z(c[61]) );
  AN2D0 C892 ( .A1(p[59]), .A2(c[59]), .Z(N59) );
  OR2D0 C891 ( .A1(g[59]), .A2(N59), .Z(c[60]) );
  AN2D0 C890 ( .A1(p[58]), .A2(c[58]), .Z(N58) );
  OR2D0 C889 ( .A1(g[58]), .A2(N58), .Z(c[59]) );
  AN2D0 C888 ( .A1(p[57]), .A2(c[57]), .Z(N57) );
  OR2D0 C887 ( .A1(g[57]), .A2(N57), .Z(c[58]) );
  AN2D0 C886 ( .A1(p[56]), .A2(c[56]), .Z(N56) );
  OR2D0 C885 ( .A1(g[56]), .A2(N56), .Z(c[57]) );
  AN2D0 C884 ( .A1(p[55]), .A2(c[55]), .Z(N55) );
  OR2D0 C883 ( .A1(g[55]), .A2(N55), .Z(c[56]) );
  AN2D0 C882 ( .A1(p[54]), .A2(c[54]), .Z(N54) );
  OR2D0 C881 ( .A1(g[54]), .A2(N54), .Z(c[55]) );
  AN2D0 C880 ( .A1(p[53]), .A2(c[53]), .Z(N53) );
  OR2D0 C879 ( .A1(g[53]), .A2(N53), .Z(c[54]) );
  AN2D0 C878 ( .A1(p[52]), .A2(c[52]), .Z(N52) );
  OR2D0 C877 ( .A1(g[52]), .A2(N52), .Z(c[53]) );
  AN2D0 C876 ( .A1(p[51]), .A2(c[51]), .Z(N51) );
  OR2D0 C875 ( .A1(g[51]), .A2(N51), .Z(c[52]) );
  AN2D0 C874 ( .A1(p[50]), .A2(c[50]), .Z(N50) );
  OR2D0 C873 ( .A1(g[50]), .A2(N50), .Z(c[51]) );
  AN2D0 C872 ( .A1(p[49]), .A2(c[49]), .Z(N49) );
  OR2D0 C871 ( .A1(g[49]), .A2(N49), .Z(c[50]) );
  AN2D0 C870 ( .A1(p[48]), .A2(c[48]), .Z(N48) );
  OR2D0 C869 ( .A1(g[48]), .A2(N48), .Z(c[49]) );
  AN2D0 C868 ( .A1(p[47]), .A2(c[47]), .Z(N47) );
  OR2D0 C867 ( .A1(g[47]), .A2(N47), .Z(c[48]) );
  AN2D0 C866 ( .A1(p[46]), .A2(c[46]), .Z(N46) );
  OR2D0 C865 ( .A1(g[46]), .A2(N46), .Z(c[47]) );
  AN2D0 C864 ( .A1(p[45]), .A2(c[45]), .Z(N45) );
  OR2D0 C863 ( .A1(g[45]), .A2(N45), .Z(c[46]) );
  AN2D0 C862 ( .A1(p[44]), .A2(c[44]), .Z(N44) );
  OR2D0 C861 ( .A1(g[44]), .A2(N44), .Z(c[45]) );
  AN2D0 C860 ( .A1(p[43]), .A2(c[43]), .Z(N43) );
  OR2D0 C859 ( .A1(g[43]), .A2(N43), .Z(c[44]) );
  AN2D0 C858 ( .A1(p[42]), .A2(c[42]), .Z(N42) );
  OR2D0 C857 ( .A1(g[42]), .A2(N42), .Z(c[43]) );
  AN2D0 C856 ( .A1(p[41]), .A2(c[41]), .Z(N41) );
  OR2D0 C855 ( .A1(g[41]), .A2(N41), .Z(c[42]) );
  AN2D0 C854 ( .A1(p[40]), .A2(c[40]), .Z(N40) );
  OR2D0 C853 ( .A1(g[40]), .A2(N40), .Z(c[41]) );
  AN2D0 C852 ( .A1(p[39]), .A2(c[39]), .Z(N39) );
  OR2D0 C851 ( .A1(g[39]), .A2(N39), .Z(c[40]) );
  AN2D0 C850 ( .A1(p[38]), .A2(c[38]), .Z(N38) );
  OR2D0 C849 ( .A1(g[38]), .A2(N38), .Z(c[39]) );
  AN2D0 C848 ( .A1(p[37]), .A2(c[37]), .Z(N37) );
  OR2D0 C847 ( .A1(g[37]), .A2(N37), .Z(c[38]) );
  AN2D0 C846 ( .A1(p[36]), .A2(c[36]), .Z(N36) );
  OR2D0 C845 ( .A1(g[36]), .A2(N36), .Z(c[37]) );
  AN2D0 C844 ( .A1(p[35]), .A2(c[35]), .Z(N35) );
  OR2D0 C843 ( .A1(g[35]), .A2(N35), .Z(c[36]) );
  AN2D0 C842 ( .A1(p[34]), .A2(c[34]), .Z(N34) );
  OR2D0 C841 ( .A1(g[34]), .A2(N34), .Z(c[35]) );
  AN2D0 C840 ( .A1(p[33]), .A2(c[33]), .Z(N33) );
  OR2D0 C839 ( .A1(g[33]), .A2(N33), .Z(c[34]) );
  AN2D0 C838 ( .A1(p[32]), .A2(c[32]), .Z(N32) );
  OR2D0 C837 ( .A1(g[32]), .A2(N32), .Z(c[33]) );
  AN2D0 C836 ( .A1(p[31]), .A2(c[31]), .Z(N31) );
  OR2D0 C835 ( .A1(g[31]), .A2(N31), .Z(c[32]) );
  AN2D0 C834 ( .A1(p[30]), .A2(c[30]), .Z(N30) );
  OR2D0 C833 ( .A1(g[30]), .A2(N30), .Z(c[31]) );
  AN2D0 C832 ( .A1(p[29]), .A2(c[29]), .Z(N29) );
  OR2D0 C831 ( .A1(g[29]), .A2(N29), .Z(c[30]) );
  AN2D0 C830 ( .A1(p[28]), .A2(c[28]), .Z(N28) );
  OR2D0 C829 ( .A1(g[28]), .A2(N28), .Z(c[29]) );
  AN2D0 C828 ( .A1(p[27]), .A2(c[27]), .Z(N27) );
  OR2D0 C827 ( .A1(g[27]), .A2(N27), .Z(c[28]) );
  AN2D0 C826 ( .A1(p[26]), .A2(c[26]), .Z(N26) );
  OR2D0 C825 ( .A1(g[26]), .A2(N26), .Z(c[27]) );
  AN2D0 C824 ( .A1(p[25]), .A2(c[25]), .Z(N25) );
  OR2D0 C823 ( .A1(g[25]), .A2(N25), .Z(c[26]) );
  AN2D0 C822 ( .A1(p[24]), .A2(c[24]), .Z(N24) );
  OR2D0 C821 ( .A1(g[24]), .A2(N24), .Z(c[25]) );
  AN2D0 C820 ( .A1(p[23]), .A2(c[23]), .Z(N23) );
  OR2D0 C819 ( .A1(g[23]), .A2(N23), .Z(c[24]) );
  AN2D0 C818 ( .A1(p[22]), .A2(c[22]), .Z(N22) );
  OR2D0 C817 ( .A1(g[22]), .A2(N22), .Z(c[23]) );
  AN2D0 C816 ( .A1(p[21]), .A2(c[21]), .Z(N21) );
  OR2D0 C815 ( .A1(g[21]), .A2(N21), .Z(c[22]) );
  AN2D0 C814 ( .A1(p[20]), .A2(c[20]), .Z(N20) );
  OR2D0 C813 ( .A1(g[20]), .A2(N20), .Z(c[21]) );
  AN2D0 C812 ( .A1(p[19]), .A2(c[19]), .Z(N19) );
  OR2D0 C811 ( .A1(g[19]), .A2(N19), .Z(c[20]) );
  AN2D0 C810 ( .A1(p[18]), .A2(c[18]), .Z(N18) );
  OR2D0 C809 ( .A1(g[18]), .A2(N18), .Z(c[19]) );
  AN2D0 C808 ( .A1(p[17]), .A2(c[17]), .Z(N17) );
  OR2D0 C807 ( .A1(g[17]), .A2(N17), .Z(c[18]) );
  AN2D0 C806 ( .A1(p[16]), .A2(c[16]), .Z(N16) );
  OR2D0 C805 ( .A1(g[16]), .A2(N16), .Z(c[17]) );
  AN2D0 C804 ( .A1(p[15]), .A2(c[15]), .Z(N15) );
  OR2D0 C803 ( .A1(g[15]), .A2(N15), .Z(c[16]) );
  AN2D0 C802 ( .A1(p[14]), .A2(c[14]), .Z(N14) );
  OR2D0 C801 ( .A1(g[14]), .A2(N14), .Z(c[15]) );
  AN2D0 C800 ( .A1(p[13]), .A2(c[13]), .Z(N13) );
  OR2D0 C799 ( .A1(g[13]), .A2(N13), .Z(c[14]) );
  AN2D0 C798 ( .A1(p[12]), .A2(c[12]), .Z(N12) );
  OR2D0 C797 ( .A1(g[12]), .A2(N12), .Z(c[13]) );
  AN2D0 C796 ( .A1(p[11]), .A2(c[11]), .Z(N11) );
  OR2D0 C795 ( .A1(g[11]), .A2(N11), .Z(c[12]) );
  AN2D0 C794 ( .A1(p[10]), .A2(c[10]), .Z(N10) );
  OR2D0 C793 ( .A1(g[10]), .A2(N10), .Z(c[11]) );
  AN2D0 C792 ( .A1(p[9]), .A2(c[9]), .Z(N9) );
  OR2D0 C791 ( .A1(g[9]), .A2(N9), .Z(c[10]) );
  AN2D0 C790 ( .A1(p[8]), .A2(c[8]), .Z(N8) );
  OR2D0 C789 ( .A1(g[8]), .A2(N8), .Z(c[9]) );
  AN2D0 C788 ( .A1(p[7]), .A2(c[7]), .Z(N7) );
  OR2D0 C787 ( .A1(g[7]), .A2(N7), .Z(c[8]) );
  AN2D0 C786 ( .A1(p[6]), .A2(c[6]), .Z(N6) );
  OR2D0 C785 ( .A1(g[6]), .A2(N6), .Z(c[7]) );
  AN2D0 C784 ( .A1(p[5]), .A2(c[5]), .Z(N5) );
  OR2D0 C783 ( .A1(g[5]), .A2(N5), .Z(c[6]) );
  AN2D0 C782 ( .A1(p[4]), .A2(c[4]), .Z(N4) );
  OR2D0 C781 ( .A1(g[4]), .A2(N4), .Z(c[5]) );
  AN2D0 C780 ( .A1(p[3]), .A2(c[3]), .Z(N3) );
  OR2D0 C779 ( .A1(g[3]), .A2(N3), .Z(c[4]) );
  AN2D0 C778 ( .A1(p[2]), .A2(c[2]), .Z(N2) );
  OR2D0 C777 ( .A1(g[2]), .A2(N2), .Z(c[3]) );
  AN2D0 C776 ( .A1(p[1]), .A2(c[1]), .Z(N1) );
  OR2D0 C775 ( .A1(g[1]), .A2(N1), .Z(c[2]) );
  AN2D0 C774 ( .A1(p[0]), .A2(cin), .Z(N0) );
  OR2D0 C773 ( .A1(g[0]), .A2(N0), .Z(c[1]) );
  XOR2D0 C772 ( .A1(a[0]), .A2(b[0]), .Z(p[0]) );
  XOR2D0 C771 ( .A1(a[1]), .A2(b[1]), .Z(p[1]) );
  XOR2D0 C770 ( .A1(a[2]), .A2(b[2]), .Z(p[2]) );
  XOR2D0 C769 ( .A1(a[3]), .A2(b[3]), .Z(p[3]) );
  XOR2D0 C768 ( .A1(a[4]), .A2(b[4]), .Z(p[4]) );
  XOR2D0 C767 ( .A1(a[5]), .A2(b[5]), .Z(p[5]) );
  XOR2D0 C766 ( .A1(a[6]), .A2(b[6]), .Z(p[6]) );
  XOR2D0 C765 ( .A1(a[7]), .A2(b[7]), .Z(p[7]) );
  XOR2D0 C764 ( .A1(a[8]), .A2(b[8]), .Z(p[8]) );
  XOR2D0 C763 ( .A1(a[9]), .A2(b[9]), .Z(p[9]) );
  XOR2D0 C762 ( .A1(a[10]), .A2(b[10]), .Z(p[10]) );
  XOR2D0 C761 ( .A1(a[11]), .A2(b[11]), .Z(p[11]) );
  XOR2D0 C760 ( .A1(a[12]), .A2(b[12]), .Z(p[12]) );
  XOR2D0 C759 ( .A1(a[13]), .A2(b[13]), .Z(p[13]) );
  XOR2D0 C758 ( .A1(a[14]), .A2(b[14]), .Z(p[14]) );
  XOR2D0 C757 ( .A1(a[15]), .A2(b[15]), .Z(p[15]) );
  XOR2D0 C756 ( .A1(a[16]), .A2(b[16]), .Z(p[16]) );
  XOR2D0 C755 ( .A1(a[17]), .A2(b[17]), .Z(p[17]) );
  XOR2D0 C754 ( .A1(a[18]), .A2(b[18]), .Z(p[18]) );
  XOR2D0 C753 ( .A1(a[19]), .A2(b[19]), .Z(p[19]) );
  XOR2D0 C752 ( .A1(a[20]), .A2(b[20]), .Z(p[20]) );
  XOR2D0 C751 ( .A1(a[21]), .A2(b[21]), .Z(p[21]) );
  XOR2D0 C750 ( .A1(a[22]), .A2(b[22]), .Z(p[22]) );
  XOR2D0 C749 ( .A1(a[23]), .A2(b[23]), .Z(p[23]) );
  XOR2D0 C748 ( .A1(a[24]), .A2(b[24]), .Z(p[24]) );
  XOR2D0 C747 ( .A1(a[25]), .A2(b[25]), .Z(p[25]) );
  XOR2D0 C746 ( .A1(a[26]), .A2(b[26]), .Z(p[26]) );
  XOR2D0 C745 ( .A1(a[27]), .A2(b[27]), .Z(p[27]) );
  XOR2D0 C744 ( .A1(a[28]), .A2(b[28]), .Z(p[28]) );
  XOR2D0 C743 ( .A1(a[29]), .A2(b[29]), .Z(p[29]) );
  XOR2D0 C742 ( .A1(a[30]), .A2(b[30]), .Z(p[30]) );
  XOR2D0 C741 ( .A1(a[31]), .A2(b[31]), .Z(p[31]) );
  XOR2D0 C740 ( .A1(a[32]), .A2(b[32]), .Z(p[32]) );
  XOR2D0 C739 ( .A1(a[33]), .A2(b[33]), .Z(p[33]) );
  XOR2D0 C738 ( .A1(a[34]), .A2(b[34]), .Z(p[34]) );
  XOR2D0 C737 ( .A1(a[35]), .A2(b[35]), .Z(p[35]) );
  XOR2D0 C736 ( .A1(a[36]), .A2(b[36]), .Z(p[36]) );
  XOR2D0 C735 ( .A1(a[37]), .A2(b[37]), .Z(p[37]) );
  XOR2D0 C734 ( .A1(a[38]), .A2(b[38]), .Z(p[38]) );
  XOR2D0 C733 ( .A1(a[39]), .A2(b[39]), .Z(p[39]) );
  XOR2D0 C732 ( .A1(a[40]), .A2(b[40]), .Z(p[40]) );
  XOR2D0 C731 ( .A1(a[41]), .A2(b[41]), .Z(p[41]) );
  XOR2D0 C730 ( .A1(a[42]), .A2(b[42]), .Z(p[42]) );
  XOR2D0 C729 ( .A1(a[43]), .A2(b[43]), .Z(p[43]) );
  XOR2D0 C728 ( .A1(a[44]), .A2(b[44]), .Z(p[44]) );
  XOR2D0 C727 ( .A1(a[45]), .A2(b[45]), .Z(p[45]) );
  XOR2D0 C726 ( .A1(a[46]), .A2(b[46]), .Z(p[46]) );
  XOR2D0 C725 ( .A1(a[47]), .A2(b[47]), .Z(p[47]) );
  XOR2D0 C724 ( .A1(a[48]), .A2(b[48]), .Z(p[48]) );
  XOR2D0 C723 ( .A1(a[49]), .A2(b[49]), .Z(p[49]) );
  XOR2D0 C722 ( .A1(a[50]), .A2(b[50]), .Z(p[50]) );
  XOR2D0 C721 ( .A1(a[51]), .A2(b[51]), .Z(p[51]) );
  XOR2D0 C720 ( .A1(a[52]), .A2(b[52]), .Z(p[52]) );
  XOR2D0 C719 ( .A1(a[53]), .A2(b[53]), .Z(p[53]) );
  XOR2D0 C718 ( .A1(a[54]), .A2(b[54]), .Z(p[54]) );
  XOR2D0 C717 ( .A1(a[55]), .A2(b[55]), .Z(p[55]) );
  XOR2D0 C716 ( .A1(a[56]), .A2(b[56]), .Z(p[56]) );
  XOR2D0 C715 ( .A1(a[57]), .A2(b[57]), .Z(p[57]) );
  XOR2D0 C714 ( .A1(a[58]), .A2(b[58]), .Z(p[58]) );
  XOR2D0 C713 ( .A1(a[59]), .A2(b[59]), .Z(p[59]) );
  XOR2D0 C712 ( .A1(a[60]), .A2(b[60]), .Z(p[60]) );
  XOR2D0 C711 ( .A1(a[61]), .A2(b[61]), .Z(p[61]) );
  XOR2D0 C710 ( .A1(a[62]), .A2(b[62]), .Z(p[62]) );
  XOR2D0 C709 ( .A1(a[63]), .A2(b[63]), .Z(p[63]) );
  XOR2D0 C708 ( .A1(a[64]), .A2(b[64]), .Z(p[64]) );
  XOR2D0 C707 ( .A1(a[65]), .A2(b[65]), .Z(p[65]) );
  XOR2D0 C706 ( .A1(a[66]), .A2(b[66]), .Z(p[66]) );
  XOR2D0 C705 ( .A1(a[67]), .A2(b[67]), .Z(p[67]) );
  XOR2D0 C704 ( .A1(a[68]), .A2(b[68]), .Z(p[68]) );
  XOR2D0 C703 ( .A1(a[69]), .A2(b[69]), .Z(p[69]) );
  XOR2D0 C702 ( .A1(a[70]), .A2(b[70]), .Z(p[70]) );
  XOR2D0 C701 ( .A1(a[71]), .A2(b[71]), .Z(p[71]) );
  XOR2D0 C700 ( .A1(a[72]), .A2(b[72]), .Z(p[72]) );
  XOR2D0 C699 ( .A1(a[73]), .A2(b[73]), .Z(p[73]) );
  XOR2D0 C698 ( .A1(a[74]), .A2(b[74]), .Z(p[74]) );
  XOR2D0 C697 ( .A1(a[75]), .A2(b[75]), .Z(p[75]) );
  XOR2D0 C696 ( .A1(a[76]), .A2(b[76]), .Z(p[76]) );
  XOR2D0 C695 ( .A1(a[77]), .A2(b[77]), .Z(p[77]) );
  XOR2D0 C694 ( .A1(a[78]), .A2(b[78]), .Z(p[78]) );
  XOR2D0 C693 ( .A1(a[79]), .A2(b[79]), .Z(p[79]) );
  XOR2D0 C692 ( .A1(a[80]), .A2(b[80]), .Z(p[80]) );
  XOR2D0 C691 ( .A1(a[81]), .A2(b[81]), .Z(p[81]) );
  XOR2D0 C690 ( .A1(a[82]), .A2(b[82]), .Z(p[82]) );
  XOR2D0 C689 ( .A1(a[83]), .A2(b[83]), .Z(p[83]) );
  XOR2D0 C688 ( .A1(a[84]), .A2(b[84]), .Z(p[84]) );
  XOR2D0 C687 ( .A1(a[85]), .A2(b[85]), .Z(p[85]) );
  XOR2D0 C686 ( .A1(a[86]), .A2(b[86]), .Z(p[86]) );
  XOR2D0 C685 ( .A1(a[87]), .A2(b[87]), .Z(p[87]) );
  XOR2D0 C684 ( .A1(a[88]), .A2(b[88]), .Z(p[88]) );
  XOR2D0 C683 ( .A1(a[89]), .A2(b[89]), .Z(p[89]) );
  XOR2D0 C682 ( .A1(a[90]), .A2(b[90]), .Z(p[90]) );
  XOR2D0 C681 ( .A1(a[91]), .A2(b[91]), .Z(p[91]) );
  XOR2D0 C680 ( .A1(a[92]), .A2(b[92]), .Z(p[92]) );
  XOR2D0 C679 ( .A1(a[93]), .A2(b[93]), .Z(p[93]) );
  XOR2D0 C678 ( .A1(a[94]), .A2(b[94]), .Z(p[94]) );
  XOR2D0 C677 ( .A1(a[95]), .A2(b[95]), .Z(p[95]) );
  XOR2D0 C676 ( .A1(a[96]), .A2(b[96]), .Z(p[96]) );
  XOR2D0 C675 ( .A1(a[97]), .A2(b[97]), .Z(p[97]) );
  XOR2D0 C674 ( .A1(a[98]), .A2(b[98]), .Z(p[98]) );
  XOR2D0 C673 ( .A1(a[99]), .A2(b[99]), .Z(p[99]) );
  XOR2D0 C672 ( .A1(a[100]), .A2(b[100]), .Z(p[100]) );
  XOR2D0 C671 ( .A1(a[101]), .A2(b[101]), .Z(p[101]) );
  XOR2D0 C670 ( .A1(a[102]), .A2(b[102]), .Z(p[102]) );
  XOR2D0 C669 ( .A1(a[103]), .A2(b[103]), .Z(p[103]) );
  XOR2D0 C668 ( .A1(a[104]), .A2(b[104]), .Z(p[104]) );
  XOR2D0 C667 ( .A1(a[105]), .A2(b[105]), .Z(p[105]) );
  XOR2D0 C666 ( .A1(a[106]), .A2(b[106]), .Z(p[106]) );
  XOR2D0 C665 ( .A1(a[107]), .A2(b[107]), .Z(p[107]) );
  XOR2D0 C664 ( .A1(a[108]), .A2(b[108]), .Z(p[108]) );
  XOR2D0 C663 ( .A1(a[109]), .A2(b[109]), .Z(p[109]) );
  XOR2D0 C662 ( .A1(a[110]), .A2(b[110]), .Z(p[110]) );
  XOR2D0 C661 ( .A1(a[111]), .A2(b[111]), .Z(p[111]) );
  XOR2D0 C660 ( .A1(a[112]), .A2(b[112]), .Z(p[112]) );
  XOR2D0 C659 ( .A1(a[113]), .A2(b[113]), .Z(p[113]) );
  XOR2D0 C658 ( .A1(a[114]), .A2(b[114]), .Z(p[114]) );
  XOR2D0 C657 ( .A1(a[115]), .A2(b[115]), .Z(p[115]) );
  XOR2D0 C656 ( .A1(a[116]), .A2(b[116]), .Z(p[116]) );
  XOR2D0 C655 ( .A1(a[117]), .A2(b[117]), .Z(p[117]) );
  XOR2D0 C654 ( .A1(a[118]), .A2(b[118]), .Z(p[118]) );
  XOR2D0 C653 ( .A1(a[119]), .A2(b[119]), .Z(p[119]) );
  XOR2D0 C652 ( .A1(a[120]), .A2(b[120]), .Z(p[120]) );
  XOR2D0 C651 ( .A1(a[121]), .A2(b[121]), .Z(p[121]) );
  XOR2D0 C650 ( .A1(a[122]), .A2(b[122]), .Z(p[122]) );
  XOR2D0 C649 ( .A1(a[123]), .A2(b[123]), .Z(p[123]) );
  XOR2D0 C648 ( .A1(a[124]), .A2(b[124]), .Z(p[124]) );
  XOR2D0 C647 ( .A1(a[125]), .A2(b[125]), .Z(p[125]) );
  XOR2D0 C646 ( .A1(a[126]), .A2(b[126]), .Z(p[126]) );
  XOR2D0 C645 ( .A1(a[127]), .A2(b[127]), .Z(p[127]) );
  AN2D0 C644 ( .A1(a[0]), .A2(b[0]), .Z(g[0]) );
  AN2D0 C643 ( .A1(a[1]), .A2(b[1]), .Z(g[1]) );
  AN2D0 C642 ( .A1(a[2]), .A2(b[2]), .Z(g[2]) );
  AN2D0 C641 ( .A1(a[3]), .A2(b[3]), .Z(g[3]) );
  AN2D0 C640 ( .A1(a[4]), .A2(b[4]), .Z(g[4]) );
  AN2D0 C639 ( .A1(a[5]), .A2(b[5]), .Z(g[5]) );
  AN2D0 C638 ( .A1(a[6]), .A2(b[6]), .Z(g[6]) );
  AN2D0 C637 ( .A1(a[7]), .A2(b[7]), .Z(g[7]) );
  AN2D0 C636 ( .A1(a[8]), .A2(b[8]), .Z(g[8]) );
  AN2D0 C635 ( .A1(a[9]), .A2(b[9]), .Z(g[9]) );
  AN2D0 C634 ( .A1(a[10]), .A2(b[10]), .Z(g[10]) );
  AN2D0 C633 ( .A1(a[11]), .A2(b[11]), .Z(g[11]) );
  AN2D0 C632 ( .A1(a[12]), .A2(b[12]), .Z(g[12]) );
  AN2D0 C631 ( .A1(a[13]), .A2(b[13]), .Z(g[13]) );
  AN2D0 C630 ( .A1(a[14]), .A2(b[14]), .Z(g[14]) );
  AN2D0 C629 ( .A1(a[15]), .A2(b[15]), .Z(g[15]) );
  AN2D0 C628 ( .A1(a[16]), .A2(b[16]), .Z(g[16]) );
  AN2D0 C627 ( .A1(a[17]), .A2(b[17]), .Z(g[17]) );
  AN2D0 C626 ( .A1(a[18]), .A2(b[18]), .Z(g[18]) );
  AN2D0 C625 ( .A1(a[19]), .A2(b[19]), .Z(g[19]) );
  AN2D0 C624 ( .A1(a[20]), .A2(b[20]), .Z(g[20]) );
  AN2D0 C623 ( .A1(a[21]), .A2(b[21]), .Z(g[21]) );
  AN2D0 C622 ( .A1(a[22]), .A2(b[22]), .Z(g[22]) );
  AN2D0 C621 ( .A1(a[23]), .A2(b[23]), .Z(g[23]) );
  AN2D0 C620 ( .A1(a[24]), .A2(b[24]), .Z(g[24]) );
  AN2D0 C619 ( .A1(a[25]), .A2(b[25]), .Z(g[25]) );
  AN2D0 C618 ( .A1(a[26]), .A2(b[26]), .Z(g[26]) );
  AN2D0 C617 ( .A1(a[27]), .A2(b[27]), .Z(g[27]) );
  AN2D0 C616 ( .A1(a[28]), .A2(b[28]), .Z(g[28]) );
  AN2D0 C615 ( .A1(a[29]), .A2(b[29]), .Z(g[29]) );
  AN2D0 C614 ( .A1(a[30]), .A2(b[30]), .Z(g[30]) );
  AN2D0 C613 ( .A1(a[31]), .A2(b[31]), .Z(g[31]) );
  AN2D0 C612 ( .A1(a[32]), .A2(b[32]), .Z(g[32]) );
  AN2D0 C611 ( .A1(a[33]), .A2(b[33]), .Z(g[33]) );
  AN2D0 C610 ( .A1(a[34]), .A2(b[34]), .Z(g[34]) );
  AN2D0 C609 ( .A1(a[35]), .A2(b[35]), .Z(g[35]) );
  AN2D0 C608 ( .A1(a[36]), .A2(b[36]), .Z(g[36]) );
  AN2D0 C607 ( .A1(a[37]), .A2(b[37]), .Z(g[37]) );
  AN2D0 C606 ( .A1(a[38]), .A2(b[38]), .Z(g[38]) );
  AN2D0 C605 ( .A1(a[39]), .A2(b[39]), .Z(g[39]) );
  AN2D0 C604 ( .A1(a[40]), .A2(b[40]), .Z(g[40]) );
  AN2D0 C603 ( .A1(a[41]), .A2(b[41]), .Z(g[41]) );
  AN2D0 C602 ( .A1(a[42]), .A2(b[42]), .Z(g[42]) );
  AN2D0 C601 ( .A1(a[43]), .A2(b[43]), .Z(g[43]) );
  AN2D0 C600 ( .A1(a[44]), .A2(b[44]), .Z(g[44]) );
  AN2D0 C599 ( .A1(a[45]), .A2(b[45]), .Z(g[45]) );
  AN2D0 C598 ( .A1(a[46]), .A2(b[46]), .Z(g[46]) );
  AN2D0 C597 ( .A1(a[47]), .A2(b[47]), .Z(g[47]) );
  AN2D0 C596 ( .A1(a[48]), .A2(b[48]), .Z(g[48]) );
  AN2D0 C595 ( .A1(a[49]), .A2(b[49]), .Z(g[49]) );
  AN2D0 C594 ( .A1(a[50]), .A2(b[50]), .Z(g[50]) );
  AN2D0 C593 ( .A1(a[51]), .A2(b[51]), .Z(g[51]) );
  AN2D0 C592 ( .A1(a[52]), .A2(b[52]), .Z(g[52]) );
  AN2D0 C591 ( .A1(a[53]), .A2(b[53]), .Z(g[53]) );
  AN2D0 C590 ( .A1(a[54]), .A2(b[54]), .Z(g[54]) );
  AN2D0 C589 ( .A1(a[55]), .A2(b[55]), .Z(g[55]) );
  AN2D0 C588 ( .A1(a[56]), .A2(b[56]), .Z(g[56]) );
  AN2D0 C587 ( .A1(a[57]), .A2(b[57]), .Z(g[57]) );
  AN2D0 C586 ( .A1(a[58]), .A2(b[58]), .Z(g[58]) );
  AN2D0 C585 ( .A1(a[59]), .A2(b[59]), .Z(g[59]) );
  AN2D0 C584 ( .A1(a[60]), .A2(b[60]), .Z(g[60]) );
  AN2D0 C583 ( .A1(a[61]), .A2(b[61]), .Z(g[61]) );
  AN2D0 C582 ( .A1(a[62]), .A2(b[62]), .Z(g[62]) );
  AN2D0 C581 ( .A1(a[63]), .A2(b[63]), .Z(g[63]) );
  AN2D0 C580 ( .A1(a[64]), .A2(b[64]), .Z(g[64]) );
  AN2D0 C579 ( .A1(a[65]), .A2(b[65]), .Z(g[65]) );
  AN2D0 C578 ( .A1(a[66]), .A2(b[66]), .Z(g[66]) );
  AN2D0 C577 ( .A1(a[67]), .A2(b[67]), .Z(g[67]) );
  AN2D0 C576 ( .A1(a[68]), .A2(b[68]), .Z(g[68]) );
  AN2D0 C575 ( .A1(a[69]), .A2(b[69]), .Z(g[69]) );
  AN2D0 C574 ( .A1(a[70]), .A2(b[70]), .Z(g[70]) );
  AN2D0 C573 ( .A1(a[71]), .A2(b[71]), .Z(g[71]) );
  AN2D0 C572 ( .A1(a[72]), .A2(b[72]), .Z(g[72]) );
  AN2D0 C571 ( .A1(a[73]), .A2(b[73]), .Z(g[73]) );
  AN2D0 C570 ( .A1(a[74]), .A2(b[74]), .Z(g[74]) );
  AN2D0 C569 ( .A1(a[75]), .A2(b[75]), .Z(g[75]) );
  AN2D0 C568 ( .A1(a[76]), .A2(b[76]), .Z(g[76]) );
  AN2D0 C567 ( .A1(a[77]), .A2(b[77]), .Z(g[77]) );
  AN2D0 C566 ( .A1(a[78]), .A2(b[78]), .Z(g[78]) );
  AN2D0 C565 ( .A1(a[79]), .A2(b[79]), .Z(g[79]) );
  AN2D0 C564 ( .A1(a[80]), .A2(b[80]), .Z(g[80]) );
  AN2D0 C563 ( .A1(a[81]), .A2(b[81]), .Z(g[81]) );
  AN2D0 C562 ( .A1(a[82]), .A2(b[82]), .Z(g[82]) );
  AN2D0 C561 ( .A1(a[83]), .A2(b[83]), .Z(g[83]) );
  AN2D0 C560 ( .A1(a[84]), .A2(b[84]), .Z(g[84]) );
  AN2D0 C559 ( .A1(a[85]), .A2(b[85]), .Z(g[85]) );
  AN2D0 C558 ( .A1(a[86]), .A2(b[86]), .Z(g[86]) );
  AN2D0 C557 ( .A1(a[87]), .A2(b[87]), .Z(g[87]) );
  AN2D0 C556 ( .A1(a[88]), .A2(b[88]), .Z(g[88]) );
  AN2D0 C555 ( .A1(a[89]), .A2(b[89]), .Z(g[89]) );
  AN2D0 C554 ( .A1(a[90]), .A2(b[90]), .Z(g[90]) );
  AN2D0 C553 ( .A1(a[91]), .A2(b[91]), .Z(g[91]) );
  AN2D0 C552 ( .A1(a[92]), .A2(b[92]), .Z(g[92]) );
  AN2D0 C551 ( .A1(a[93]), .A2(b[93]), .Z(g[93]) );
  AN2D0 C550 ( .A1(a[94]), .A2(b[94]), .Z(g[94]) );
  AN2D0 C549 ( .A1(a[95]), .A2(b[95]), .Z(g[95]) );
  AN2D0 C548 ( .A1(a[96]), .A2(b[96]), .Z(g[96]) );
  AN2D0 C547 ( .A1(a[97]), .A2(b[97]), .Z(g[97]) );
  AN2D0 C546 ( .A1(a[98]), .A2(b[98]), .Z(g[98]) );
  AN2D0 C545 ( .A1(a[99]), .A2(b[99]), .Z(g[99]) );
  AN2D0 C544 ( .A1(a[100]), .A2(b[100]), .Z(g[100]) );
  AN2D0 C543 ( .A1(a[101]), .A2(b[101]), .Z(g[101]) );
  AN2D0 C542 ( .A1(a[102]), .A2(b[102]), .Z(g[102]) );
  AN2D0 C541 ( .A1(a[103]), .A2(b[103]), .Z(g[103]) );
  AN2D0 C540 ( .A1(a[104]), .A2(b[104]), .Z(g[104]) );
  AN2D0 C539 ( .A1(a[105]), .A2(b[105]), .Z(g[105]) );
  AN2D0 C538 ( .A1(a[106]), .A2(b[106]), .Z(g[106]) );
  AN2D0 C537 ( .A1(a[107]), .A2(b[107]), .Z(g[107]) );
  AN2D0 C536 ( .A1(a[108]), .A2(b[108]), .Z(g[108]) );
  AN2D0 C535 ( .A1(a[109]), .A2(b[109]), .Z(g[109]) );
  AN2D0 C534 ( .A1(a[110]), .A2(b[110]), .Z(g[110]) );
  AN2D0 C533 ( .A1(a[111]), .A2(b[111]), .Z(g[111]) );
  AN2D0 C532 ( .A1(a[112]), .A2(b[112]), .Z(g[112]) );
  AN2D0 C531 ( .A1(a[113]), .A2(b[113]), .Z(g[113]) );
  AN2D0 C530 ( .A1(a[114]), .A2(b[114]), .Z(g[114]) );
  AN2D0 C529 ( .A1(a[115]), .A2(b[115]), .Z(g[115]) );
  AN2D0 C528 ( .A1(a[116]), .A2(b[116]), .Z(g[116]) );
  AN2D0 C527 ( .A1(a[117]), .A2(b[117]), .Z(g[117]) );
  AN2D0 C526 ( .A1(a[118]), .A2(b[118]), .Z(g[118]) );
  AN2D0 C525 ( .A1(a[119]), .A2(b[119]), .Z(g[119]) );
  AN2D0 C524 ( .A1(a[120]), .A2(b[120]), .Z(g[120]) );
  AN2D0 C523 ( .A1(a[121]), .A2(b[121]), .Z(g[121]) );
  AN2D0 C522 ( .A1(a[122]), .A2(b[122]), .Z(g[122]) );
  AN2D0 C521 ( .A1(a[123]), .A2(b[123]), .Z(g[123]) );
  AN2D0 C520 ( .A1(a[124]), .A2(b[124]), .Z(g[124]) );
  AN2D0 C519 ( .A1(a[125]), .A2(b[125]), .Z(g[125]) );
  AN2D0 C518 ( .A1(a[126]), .A2(b[126]), .Z(g[126]) );
endmodule

