module gen_nonlinear_part(a,b,n);
input  [15:0] a, b; //adder inputs
output [65518:0] n; // non-linear outputs

wire [65518:0] g; 

assign n = g; //assign outputs

//Assigning outputs for input bit 1
assign g[0] = a[0] & b[0];
//Assigning outputs for input bit 2
assign g[1] = a[1] & b[1];
assign g[2] = a[1] & g[0];
assign g[3] = b[1] & g[0];
//Assigning outputs for input bit 3
assign g[4] = a[2] & b[2];
assign g[5] = a[2] & g[1];
assign g[8] = b[2] & g[1];
assign g[6] = a[2] & g[2];
assign g[9] = b[2] & g[2];
assign g[7] = a[2] & g[3];
assign g[10] = b[2] & g[3];
//Assigning outputs for input bit 4
assign g[11] = a[3] & b[3];
assign g[12] = a[3] & g[4];
assign g[19] = b[3] & g[4];
assign g[13] = a[3] & g[5];
assign g[20] = b[3] & g[5];
assign g[14] = a[3] & g[6];
assign g[21] = b[3] & g[6];
assign g[15] = a[3] & g[7];
assign g[22] = b[3] & g[7];
assign g[16] = a[3] & g[8];
assign g[23] = b[3] & g[8];
assign g[17] = a[3] & g[9];
assign g[24] = b[3] & g[9];
assign g[18] = a[3] & g[10];
assign g[25] = b[3] & g[10];
//Assigning outputs for input bit 5
assign g[26] = a[4] & b[4];
assign g[27] = a[4] & g[11];
assign g[42] = b[4] & g[11];
assign g[28] = a[4] & g[12];
assign g[43] = b[4] & g[12];
assign g[29] = a[4] & g[13];
assign g[44] = b[4] & g[13];
assign g[30] = a[4] & g[14];
assign g[45] = b[4] & g[14];
assign g[31] = a[4] & g[15];
assign g[46] = b[4] & g[15];
assign g[32] = a[4] & g[16];
assign g[47] = b[4] & g[16];
assign g[33] = a[4] & g[17];
assign g[48] = b[4] & g[17];
assign g[34] = a[4] & g[18];
assign g[49] = b[4] & g[18];
assign g[35] = a[4] & g[19];
assign g[50] = b[4] & g[19];
assign g[36] = a[4] & g[20];
assign g[51] = b[4] & g[20];
assign g[37] = a[4] & g[21];
assign g[52] = b[4] & g[21];
assign g[38] = a[4] & g[22];
assign g[53] = b[4] & g[22];
assign g[39] = a[4] & g[23];
assign g[54] = b[4] & g[23];
assign g[40] = a[4] & g[24];
assign g[55] = b[4] & g[24];
assign g[41] = a[4] & g[25];
assign g[56] = b[4] & g[25];
//Assigning outputs for input bit 6
assign g[57] = a[5] & b[5];
assign g[58] = a[5] & g[26];
assign g[89] = b[5] & g[26];
assign g[59] = a[5] & g[27];
assign g[90] = b[5] & g[27];
assign g[60] = a[5] & g[28];
assign g[91] = b[5] & g[28];
assign g[61] = a[5] & g[29];
assign g[92] = b[5] & g[29];
assign g[62] = a[5] & g[30];
assign g[93] = b[5] & g[30];
assign g[63] = a[5] & g[31];
assign g[94] = b[5] & g[31];
assign g[64] = a[5] & g[32];
assign g[95] = b[5] & g[32];
assign g[65] = a[5] & g[33];
assign g[96] = b[5] & g[33];
assign g[66] = a[5] & g[34];
assign g[97] = b[5] & g[34];
assign g[67] = a[5] & g[35];
assign g[98] = b[5] & g[35];
assign g[68] = a[5] & g[36];
assign g[99] = b[5] & g[36];
assign g[69] = a[5] & g[37];
assign g[100] = b[5] & g[37];
assign g[70] = a[5] & g[38];
assign g[101] = b[5] & g[38];
assign g[71] = a[5] & g[39];
assign g[102] = b[5] & g[39];
assign g[72] = a[5] & g[40];
assign g[103] = b[5] & g[40];
assign g[73] = a[5] & g[41];
assign g[104] = b[5] & g[41];
assign g[74] = a[5] & g[42];
assign g[105] = b[5] & g[42];
assign g[75] = a[5] & g[43];
assign g[106] = b[5] & g[43];
assign g[76] = a[5] & g[44];
assign g[107] = b[5] & g[44];
assign g[77] = a[5] & g[45];
assign g[108] = b[5] & g[45];
assign g[78] = a[5] & g[46];
assign g[109] = b[5] & g[46];
assign g[79] = a[5] & g[47];
assign g[110] = b[5] & g[47];
assign g[80] = a[5] & g[48];
assign g[111] = b[5] & g[48];
assign g[81] = a[5] & g[49];
assign g[112] = b[5] & g[49];
assign g[82] = a[5] & g[50];
assign g[113] = b[5] & g[50];
assign g[83] = a[5] & g[51];
assign g[114] = b[5] & g[51];
assign g[84] = a[5] & g[52];
assign g[115] = b[5] & g[52];
assign g[85] = a[5] & g[53];
assign g[116] = b[5] & g[53];
assign g[86] = a[5] & g[54];
assign g[117] = b[5] & g[54];
assign g[87] = a[5] & g[55];
assign g[118] = b[5] & g[55];
assign g[88] = a[5] & g[56];
assign g[119] = b[5] & g[56];
//Assigning outputs for input bit 7
assign g[120] = a[6] & b[6];
assign g[121] = a[6] & g[57];
assign g[184] = b[6] & g[57];
assign g[122] = a[6] & g[58];
assign g[185] = b[6] & g[58];
assign g[123] = a[6] & g[59];
assign g[186] = b[6] & g[59];
assign g[124] = a[6] & g[60];
assign g[187] = b[6] & g[60];
assign g[125] = a[6] & g[61];
assign g[188] = b[6] & g[61];
assign g[126] = a[6] & g[62];
assign g[189] = b[6] & g[62];
assign g[127] = a[6] & g[63];
assign g[190] = b[6] & g[63];
assign g[128] = a[6] & g[64];
assign g[191] = b[6] & g[64];
assign g[129] = a[6] & g[65];
assign g[192] = b[6] & g[65];
assign g[130] = a[6] & g[66];
assign g[193] = b[6] & g[66];
assign g[131] = a[6] & g[67];
assign g[194] = b[6] & g[67];
assign g[132] = a[6] & g[68];
assign g[195] = b[6] & g[68];
assign g[133] = a[6] & g[69];
assign g[196] = b[6] & g[69];
assign g[134] = a[6] & g[70];
assign g[197] = b[6] & g[70];
assign g[135] = a[6] & g[71];
assign g[198] = b[6] & g[71];
assign g[136] = a[6] & g[72];
assign g[199] = b[6] & g[72];
assign g[137] = a[6] & g[73];
assign g[200] = b[6] & g[73];
assign g[138] = a[6] & g[74];
assign g[201] = b[6] & g[74];
assign g[139] = a[6] & g[75];
assign g[202] = b[6] & g[75];
assign g[140] = a[6] & g[76];
assign g[203] = b[6] & g[76];
assign g[141] = a[6] & g[77];
assign g[204] = b[6] & g[77];
assign g[142] = a[6] & g[78];
assign g[205] = b[6] & g[78];
assign g[143] = a[6] & g[79];
assign g[206] = b[6] & g[79];
assign g[144] = a[6] & g[80];
assign g[207] = b[6] & g[80];
assign g[145] = a[6] & g[81];
assign g[208] = b[6] & g[81];
assign g[146] = a[6] & g[82];
assign g[209] = b[6] & g[82];
assign g[147] = a[6] & g[83];
assign g[210] = b[6] & g[83];
assign g[148] = a[6] & g[84];
assign g[211] = b[6] & g[84];
assign g[149] = a[6] & g[85];
assign g[212] = b[6] & g[85];
assign g[150] = a[6] & g[86];
assign g[213] = b[6] & g[86];
assign g[151] = a[6] & g[87];
assign g[214] = b[6] & g[87];
assign g[152] = a[6] & g[88];
assign g[215] = b[6] & g[88];
assign g[153] = a[6] & g[89];
assign g[216] = b[6] & g[89];
assign g[154] = a[6] & g[90];
assign g[217] = b[6] & g[90];
assign g[155] = a[6] & g[91];
assign g[218] = b[6] & g[91];
assign g[156] = a[6] & g[92];
assign g[219] = b[6] & g[92];
assign g[157] = a[6] & g[93];
assign g[220] = b[6] & g[93];
assign g[158] = a[6] & g[94];
assign g[221] = b[6] & g[94];
assign g[159] = a[6] & g[95];
assign g[222] = b[6] & g[95];
assign g[160] = a[6] & g[96];
assign g[223] = b[6] & g[96];
assign g[161] = a[6] & g[97];
assign g[224] = b[6] & g[97];
assign g[162] = a[6] & g[98];
assign g[225] = b[6] & g[98];
assign g[163] = a[6] & g[99];
assign g[226] = b[6] & g[99];
assign g[164] = a[6] & g[100];
assign g[227] = b[6] & g[100];
assign g[165] = a[6] & g[101];
assign g[228] = b[6] & g[101];
assign g[166] = a[6] & g[102];
assign g[229] = b[6] & g[102];
assign g[167] = a[6] & g[103];
assign g[230] = b[6] & g[103];
assign g[168] = a[6] & g[104];
assign g[231] = b[6] & g[104];
assign g[169] = a[6] & g[105];
assign g[232] = b[6] & g[105];
assign g[170] = a[6] & g[106];
assign g[233] = b[6] & g[106];
assign g[171] = a[6] & g[107];
assign g[234] = b[6] & g[107];
assign g[172] = a[6] & g[108];
assign g[235] = b[6] & g[108];
assign g[173] = a[6] & g[109];
assign g[236] = b[6] & g[109];
assign g[174] = a[6] & g[110];
assign g[237] = b[6] & g[110];
assign g[175] = a[6] & g[111];
assign g[238] = b[6] & g[111];
assign g[176] = a[6] & g[112];
assign g[239] = b[6] & g[112];
assign g[177] = a[6] & g[113];
assign g[240] = b[6] & g[113];
assign g[178] = a[6] & g[114];
assign g[241] = b[6] & g[114];
assign g[179] = a[6] & g[115];
assign g[242] = b[6] & g[115];
assign g[180] = a[6] & g[116];
assign g[243] = b[6] & g[116];
assign g[181] = a[6] & g[117];
assign g[244] = b[6] & g[117];
assign g[182] = a[6] & g[118];
assign g[245] = b[6] & g[118];
assign g[183] = a[6] & g[119];
assign g[246] = b[6] & g[119];
//Assigning outputs for input bit 8
assign g[247] = a[7] & b[7];
assign g[248] = a[7] & g[120];
assign g[375] = b[7] & g[120];
assign g[249] = a[7] & g[121];
assign g[376] = b[7] & g[121];
assign g[250] = a[7] & g[122];
assign g[377] = b[7] & g[122];
assign g[251] = a[7] & g[123];
assign g[378] = b[7] & g[123];
assign g[252] = a[7] & g[124];
assign g[379] = b[7] & g[124];
assign g[253] = a[7] & g[125];
assign g[380] = b[7] & g[125];
assign g[254] = a[7] & g[126];
assign g[381] = b[7] & g[126];
assign g[255] = a[7] & g[127];
assign g[382] = b[7] & g[127];
assign g[256] = a[7] & g[128];
assign g[383] = b[7] & g[128];
assign g[257] = a[7] & g[129];
assign g[384] = b[7] & g[129];
assign g[258] = a[7] & g[130];
assign g[385] = b[7] & g[130];
assign g[259] = a[7] & g[131];
assign g[386] = b[7] & g[131];
assign g[260] = a[7] & g[132];
assign g[387] = b[7] & g[132];
assign g[261] = a[7] & g[133];
assign g[388] = b[7] & g[133];
assign g[262] = a[7] & g[134];
assign g[389] = b[7] & g[134];
assign g[263] = a[7] & g[135];
assign g[390] = b[7] & g[135];
assign g[264] = a[7] & g[136];
assign g[391] = b[7] & g[136];
assign g[265] = a[7] & g[137];
assign g[392] = b[7] & g[137];
assign g[266] = a[7] & g[138];
assign g[393] = b[7] & g[138];
assign g[267] = a[7] & g[139];
assign g[394] = b[7] & g[139];
assign g[268] = a[7] & g[140];
assign g[395] = b[7] & g[140];
assign g[269] = a[7] & g[141];
assign g[396] = b[7] & g[141];
assign g[270] = a[7] & g[142];
assign g[397] = b[7] & g[142];
assign g[271] = a[7] & g[143];
assign g[398] = b[7] & g[143];
assign g[272] = a[7] & g[144];
assign g[399] = b[7] & g[144];
assign g[273] = a[7] & g[145];
assign g[400] = b[7] & g[145];
assign g[274] = a[7] & g[146];
assign g[401] = b[7] & g[146];
assign g[275] = a[7] & g[147];
assign g[402] = b[7] & g[147];
assign g[276] = a[7] & g[148];
assign g[403] = b[7] & g[148];
assign g[277] = a[7] & g[149];
assign g[404] = b[7] & g[149];
assign g[278] = a[7] & g[150];
assign g[405] = b[7] & g[150];
assign g[279] = a[7] & g[151];
assign g[406] = b[7] & g[151];
assign g[280] = a[7] & g[152];
assign g[407] = b[7] & g[152];
assign g[281] = a[7] & g[153];
assign g[408] = b[7] & g[153];
assign g[282] = a[7] & g[154];
assign g[409] = b[7] & g[154];
assign g[283] = a[7] & g[155];
assign g[410] = b[7] & g[155];
assign g[284] = a[7] & g[156];
assign g[411] = b[7] & g[156];
assign g[285] = a[7] & g[157];
assign g[412] = b[7] & g[157];
assign g[286] = a[7] & g[158];
assign g[413] = b[7] & g[158];
assign g[287] = a[7] & g[159];
assign g[414] = b[7] & g[159];
assign g[288] = a[7] & g[160];
assign g[415] = b[7] & g[160];
assign g[289] = a[7] & g[161];
assign g[416] = b[7] & g[161];
assign g[290] = a[7] & g[162];
assign g[417] = b[7] & g[162];
assign g[291] = a[7] & g[163];
assign g[418] = b[7] & g[163];
assign g[292] = a[7] & g[164];
assign g[419] = b[7] & g[164];
assign g[293] = a[7] & g[165];
assign g[420] = b[7] & g[165];
assign g[294] = a[7] & g[166];
assign g[421] = b[7] & g[166];
assign g[295] = a[7] & g[167];
assign g[422] = b[7] & g[167];
assign g[296] = a[7] & g[168];
assign g[423] = b[7] & g[168];
assign g[297] = a[7] & g[169];
assign g[424] = b[7] & g[169];
assign g[298] = a[7] & g[170];
assign g[425] = b[7] & g[170];
assign g[299] = a[7] & g[171];
assign g[426] = b[7] & g[171];
assign g[300] = a[7] & g[172];
assign g[427] = b[7] & g[172];
assign g[301] = a[7] & g[173];
assign g[428] = b[7] & g[173];
assign g[302] = a[7] & g[174];
assign g[429] = b[7] & g[174];
assign g[303] = a[7] & g[175];
assign g[430] = b[7] & g[175];
assign g[304] = a[7] & g[176];
assign g[431] = b[7] & g[176];
assign g[305] = a[7] & g[177];
assign g[432] = b[7] & g[177];
assign g[306] = a[7] & g[178];
assign g[433] = b[7] & g[178];
assign g[307] = a[7] & g[179];
assign g[434] = b[7] & g[179];
assign g[308] = a[7] & g[180];
assign g[435] = b[7] & g[180];
assign g[309] = a[7] & g[181];
assign g[436] = b[7] & g[181];
assign g[310] = a[7] & g[182];
assign g[437] = b[7] & g[182];
assign g[311] = a[7] & g[183];
assign g[438] = b[7] & g[183];
assign g[312] = a[7] & g[184];
assign g[439] = b[7] & g[184];
assign g[313] = a[7] & g[185];
assign g[440] = b[7] & g[185];
assign g[314] = a[7] & g[186];
assign g[441] = b[7] & g[186];
assign g[315] = a[7] & g[187];
assign g[442] = b[7] & g[187];
assign g[316] = a[7] & g[188];
assign g[443] = b[7] & g[188];
assign g[317] = a[7] & g[189];
assign g[444] = b[7] & g[189];
assign g[318] = a[7] & g[190];
assign g[445] = b[7] & g[190];
assign g[319] = a[7] & g[191];
assign g[446] = b[7] & g[191];
assign g[320] = a[7] & g[192];
assign g[447] = b[7] & g[192];
assign g[321] = a[7] & g[193];
assign g[448] = b[7] & g[193];
assign g[322] = a[7] & g[194];
assign g[449] = b[7] & g[194];
assign g[323] = a[7] & g[195];
assign g[450] = b[7] & g[195];
assign g[324] = a[7] & g[196];
assign g[451] = b[7] & g[196];
assign g[325] = a[7] & g[197];
assign g[452] = b[7] & g[197];
assign g[326] = a[7] & g[198];
assign g[453] = b[7] & g[198];
assign g[327] = a[7] & g[199];
assign g[454] = b[7] & g[199];
assign g[328] = a[7] & g[200];
assign g[455] = b[7] & g[200];
assign g[329] = a[7] & g[201];
assign g[456] = b[7] & g[201];
assign g[330] = a[7] & g[202];
assign g[457] = b[7] & g[202];
assign g[331] = a[7] & g[203];
assign g[458] = b[7] & g[203];
assign g[332] = a[7] & g[204];
assign g[459] = b[7] & g[204];
assign g[333] = a[7] & g[205];
assign g[460] = b[7] & g[205];
assign g[334] = a[7] & g[206];
assign g[461] = b[7] & g[206];
assign g[335] = a[7] & g[207];
assign g[462] = b[7] & g[207];
assign g[336] = a[7] & g[208];
assign g[463] = b[7] & g[208];
assign g[337] = a[7] & g[209];
assign g[464] = b[7] & g[209];
assign g[338] = a[7] & g[210];
assign g[465] = b[7] & g[210];
assign g[339] = a[7] & g[211];
assign g[466] = b[7] & g[211];
assign g[340] = a[7] & g[212];
assign g[467] = b[7] & g[212];
assign g[341] = a[7] & g[213];
assign g[468] = b[7] & g[213];
assign g[342] = a[7] & g[214];
assign g[469] = b[7] & g[214];
assign g[343] = a[7] & g[215];
assign g[470] = b[7] & g[215];
assign g[344] = a[7] & g[216];
assign g[471] = b[7] & g[216];
assign g[345] = a[7] & g[217];
assign g[472] = b[7] & g[217];
assign g[346] = a[7] & g[218];
assign g[473] = b[7] & g[218];
assign g[347] = a[7] & g[219];
assign g[474] = b[7] & g[219];
assign g[348] = a[7] & g[220];
assign g[475] = b[7] & g[220];
assign g[349] = a[7] & g[221];
assign g[476] = b[7] & g[221];
assign g[350] = a[7] & g[222];
assign g[477] = b[7] & g[222];
assign g[351] = a[7] & g[223];
assign g[478] = b[7] & g[223];
assign g[352] = a[7] & g[224];
assign g[479] = b[7] & g[224];
assign g[353] = a[7] & g[225];
assign g[480] = b[7] & g[225];
assign g[354] = a[7] & g[226];
assign g[481] = b[7] & g[226];
assign g[355] = a[7] & g[227];
assign g[482] = b[7] & g[227];
assign g[356] = a[7] & g[228];
assign g[483] = b[7] & g[228];
assign g[357] = a[7] & g[229];
assign g[484] = b[7] & g[229];
assign g[358] = a[7] & g[230];
assign g[485] = b[7] & g[230];
assign g[359] = a[7] & g[231];
assign g[486] = b[7] & g[231];
assign g[360] = a[7] & g[232];
assign g[487] = b[7] & g[232];
assign g[361] = a[7] & g[233];
assign g[488] = b[7] & g[233];
assign g[362] = a[7] & g[234];
assign g[489] = b[7] & g[234];
assign g[363] = a[7] & g[235];
assign g[490] = b[7] & g[235];
assign g[364] = a[7] & g[236];
assign g[491] = b[7] & g[236];
assign g[365] = a[7] & g[237];
assign g[492] = b[7] & g[237];
assign g[366] = a[7] & g[238];
assign g[493] = b[7] & g[238];
assign g[367] = a[7] & g[239];
assign g[494] = b[7] & g[239];
assign g[368] = a[7] & g[240];
assign g[495] = b[7] & g[240];
assign g[369] = a[7] & g[241];
assign g[496] = b[7] & g[241];
assign g[370] = a[7] & g[242];
assign g[497] = b[7] & g[242];
assign g[371] = a[7] & g[243];
assign g[498] = b[7] & g[243];
assign g[372] = a[7] & g[244];
assign g[499] = b[7] & g[244];
assign g[373] = a[7] & g[245];
assign g[500] = b[7] & g[245];
assign g[374] = a[7] & g[246];
assign g[501] = b[7] & g[246];
//Assigning outputs for input bit 9
assign g[502] = a[8] & b[8];
assign g[503] = a[8] & g[247];
assign g[758] = b[8] & g[247];
assign g[504] = a[8] & g[248];
assign g[759] = b[8] & g[248];
assign g[505] = a[8] & g[249];
assign g[760] = b[8] & g[249];
assign g[506] = a[8] & g[250];
assign g[761] = b[8] & g[250];
assign g[507] = a[8] & g[251];
assign g[762] = b[8] & g[251];
assign g[508] = a[8] & g[252];
assign g[763] = b[8] & g[252];
assign g[509] = a[8] & g[253];
assign g[764] = b[8] & g[253];
assign g[510] = a[8] & g[254];
assign g[765] = b[8] & g[254];
assign g[511] = a[8] & g[255];
assign g[766] = b[8] & g[255];
assign g[512] = a[8] & g[256];
assign g[767] = b[8] & g[256];
assign g[513] = a[8] & g[257];
assign g[768] = b[8] & g[257];
assign g[514] = a[8] & g[258];
assign g[769] = b[8] & g[258];
assign g[515] = a[8] & g[259];
assign g[770] = b[8] & g[259];
assign g[516] = a[8] & g[260];
assign g[771] = b[8] & g[260];
assign g[517] = a[8] & g[261];
assign g[772] = b[8] & g[261];
assign g[518] = a[8] & g[262];
assign g[773] = b[8] & g[262];
assign g[519] = a[8] & g[263];
assign g[774] = b[8] & g[263];
assign g[520] = a[8] & g[264];
assign g[775] = b[8] & g[264];
assign g[521] = a[8] & g[265];
assign g[776] = b[8] & g[265];
assign g[522] = a[8] & g[266];
assign g[777] = b[8] & g[266];
assign g[523] = a[8] & g[267];
assign g[778] = b[8] & g[267];
assign g[524] = a[8] & g[268];
assign g[779] = b[8] & g[268];
assign g[525] = a[8] & g[269];
assign g[780] = b[8] & g[269];
assign g[526] = a[8] & g[270];
assign g[781] = b[8] & g[270];
assign g[527] = a[8] & g[271];
assign g[782] = b[8] & g[271];
assign g[528] = a[8] & g[272];
assign g[783] = b[8] & g[272];
assign g[529] = a[8] & g[273];
assign g[784] = b[8] & g[273];
assign g[530] = a[8] & g[274];
assign g[785] = b[8] & g[274];
assign g[531] = a[8] & g[275];
assign g[786] = b[8] & g[275];
assign g[532] = a[8] & g[276];
assign g[787] = b[8] & g[276];
assign g[533] = a[8] & g[277];
assign g[788] = b[8] & g[277];
assign g[534] = a[8] & g[278];
assign g[789] = b[8] & g[278];
assign g[535] = a[8] & g[279];
assign g[790] = b[8] & g[279];
assign g[536] = a[8] & g[280];
assign g[791] = b[8] & g[280];
assign g[537] = a[8] & g[281];
assign g[792] = b[8] & g[281];
assign g[538] = a[8] & g[282];
assign g[793] = b[8] & g[282];
assign g[539] = a[8] & g[283];
assign g[794] = b[8] & g[283];
assign g[540] = a[8] & g[284];
assign g[795] = b[8] & g[284];
assign g[541] = a[8] & g[285];
assign g[796] = b[8] & g[285];
assign g[542] = a[8] & g[286];
assign g[797] = b[8] & g[286];
assign g[543] = a[8] & g[287];
assign g[798] = b[8] & g[287];
assign g[544] = a[8] & g[288];
assign g[799] = b[8] & g[288];
assign g[545] = a[8] & g[289];
assign g[800] = b[8] & g[289];
assign g[546] = a[8] & g[290];
assign g[801] = b[8] & g[290];
assign g[547] = a[8] & g[291];
assign g[802] = b[8] & g[291];
assign g[548] = a[8] & g[292];
assign g[803] = b[8] & g[292];
assign g[549] = a[8] & g[293];
assign g[804] = b[8] & g[293];
assign g[550] = a[8] & g[294];
assign g[805] = b[8] & g[294];
assign g[551] = a[8] & g[295];
assign g[806] = b[8] & g[295];
assign g[552] = a[8] & g[296];
assign g[807] = b[8] & g[296];
assign g[553] = a[8] & g[297];
assign g[808] = b[8] & g[297];
assign g[554] = a[8] & g[298];
assign g[809] = b[8] & g[298];
assign g[555] = a[8] & g[299];
assign g[810] = b[8] & g[299];
assign g[556] = a[8] & g[300];
assign g[811] = b[8] & g[300];
assign g[557] = a[8] & g[301];
assign g[812] = b[8] & g[301];
assign g[558] = a[8] & g[302];
assign g[813] = b[8] & g[302];
assign g[559] = a[8] & g[303];
assign g[814] = b[8] & g[303];
assign g[560] = a[8] & g[304];
assign g[815] = b[8] & g[304];
assign g[561] = a[8] & g[305];
assign g[816] = b[8] & g[305];
assign g[562] = a[8] & g[306];
assign g[817] = b[8] & g[306];
assign g[563] = a[8] & g[307];
assign g[818] = b[8] & g[307];
assign g[564] = a[8] & g[308];
assign g[819] = b[8] & g[308];
assign g[565] = a[8] & g[309];
assign g[820] = b[8] & g[309];
assign g[566] = a[8] & g[310];
assign g[821] = b[8] & g[310];
assign g[567] = a[8] & g[311];
assign g[822] = b[8] & g[311];
assign g[568] = a[8] & g[312];
assign g[823] = b[8] & g[312];
assign g[569] = a[8] & g[313];
assign g[824] = b[8] & g[313];
assign g[570] = a[8] & g[314];
assign g[825] = b[8] & g[314];
assign g[571] = a[8] & g[315];
assign g[826] = b[8] & g[315];
assign g[572] = a[8] & g[316];
assign g[827] = b[8] & g[316];
assign g[573] = a[8] & g[317];
assign g[828] = b[8] & g[317];
assign g[574] = a[8] & g[318];
assign g[829] = b[8] & g[318];
assign g[575] = a[8] & g[319];
assign g[830] = b[8] & g[319];
assign g[576] = a[8] & g[320];
assign g[831] = b[8] & g[320];
assign g[577] = a[8] & g[321];
assign g[832] = b[8] & g[321];
assign g[578] = a[8] & g[322];
assign g[833] = b[8] & g[322];
assign g[579] = a[8] & g[323];
assign g[834] = b[8] & g[323];
assign g[580] = a[8] & g[324];
assign g[835] = b[8] & g[324];
assign g[581] = a[8] & g[325];
assign g[836] = b[8] & g[325];
assign g[582] = a[8] & g[326];
assign g[837] = b[8] & g[326];
assign g[583] = a[8] & g[327];
assign g[838] = b[8] & g[327];
assign g[584] = a[8] & g[328];
assign g[839] = b[8] & g[328];
assign g[585] = a[8] & g[329];
assign g[840] = b[8] & g[329];
assign g[586] = a[8] & g[330];
assign g[841] = b[8] & g[330];
assign g[587] = a[8] & g[331];
assign g[842] = b[8] & g[331];
assign g[588] = a[8] & g[332];
assign g[843] = b[8] & g[332];
assign g[589] = a[8] & g[333];
assign g[844] = b[8] & g[333];
assign g[590] = a[8] & g[334];
assign g[845] = b[8] & g[334];
assign g[591] = a[8] & g[335];
assign g[846] = b[8] & g[335];
assign g[592] = a[8] & g[336];
assign g[847] = b[8] & g[336];
assign g[593] = a[8] & g[337];
assign g[848] = b[8] & g[337];
assign g[594] = a[8] & g[338];
assign g[849] = b[8] & g[338];
assign g[595] = a[8] & g[339];
assign g[850] = b[8] & g[339];
assign g[596] = a[8] & g[340];
assign g[851] = b[8] & g[340];
assign g[597] = a[8] & g[341];
assign g[852] = b[8] & g[341];
assign g[598] = a[8] & g[342];
assign g[853] = b[8] & g[342];
assign g[599] = a[8] & g[343];
assign g[854] = b[8] & g[343];
assign g[600] = a[8] & g[344];
assign g[855] = b[8] & g[344];
assign g[601] = a[8] & g[345];
assign g[856] = b[8] & g[345];
assign g[602] = a[8] & g[346];
assign g[857] = b[8] & g[346];
assign g[603] = a[8] & g[347];
assign g[858] = b[8] & g[347];
assign g[604] = a[8] & g[348];
assign g[859] = b[8] & g[348];
assign g[605] = a[8] & g[349];
assign g[860] = b[8] & g[349];
assign g[606] = a[8] & g[350];
assign g[861] = b[8] & g[350];
assign g[607] = a[8] & g[351];
assign g[862] = b[8] & g[351];
assign g[608] = a[8] & g[352];
assign g[863] = b[8] & g[352];
assign g[609] = a[8] & g[353];
assign g[864] = b[8] & g[353];
assign g[610] = a[8] & g[354];
assign g[865] = b[8] & g[354];
assign g[611] = a[8] & g[355];
assign g[866] = b[8] & g[355];
assign g[612] = a[8] & g[356];
assign g[867] = b[8] & g[356];
assign g[613] = a[8] & g[357];
assign g[868] = b[8] & g[357];
assign g[614] = a[8] & g[358];
assign g[869] = b[8] & g[358];
assign g[615] = a[8] & g[359];
assign g[870] = b[8] & g[359];
assign g[616] = a[8] & g[360];
assign g[871] = b[8] & g[360];
assign g[617] = a[8] & g[361];
assign g[872] = b[8] & g[361];
assign g[618] = a[8] & g[362];
assign g[873] = b[8] & g[362];
assign g[619] = a[8] & g[363];
assign g[874] = b[8] & g[363];
assign g[620] = a[8] & g[364];
assign g[875] = b[8] & g[364];
assign g[621] = a[8] & g[365];
assign g[876] = b[8] & g[365];
assign g[622] = a[8] & g[366];
assign g[877] = b[8] & g[366];
assign g[623] = a[8] & g[367];
assign g[878] = b[8] & g[367];
assign g[624] = a[8] & g[368];
assign g[879] = b[8] & g[368];
assign g[625] = a[8] & g[369];
assign g[880] = b[8] & g[369];
assign g[626] = a[8] & g[370];
assign g[881] = b[8] & g[370];
assign g[627] = a[8] & g[371];
assign g[882] = b[8] & g[371];
assign g[628] = a[8] & g[372];
assign g[883] = b[8] & g[372];
assign g[629] = a[8] & g[373];
assign g[884] = b[8] & g[373];
assign g[630] = a[8] & g[374];
assign g[885] = b[8] & g[374];
assign g[631] = a[8] & g[375];
assign g[886] = b[8] & g[375];
assign g[632] = a[8] & g[376];
assign g[887] = b[8] & g[376];
assign g[633] = a[8] & g[377];
assign g[888] = b[8] & g[377];
assign g[634] = a[8] & g[378];
assign g[889] = b[8] & g[378];
assign g[635] = a[8] & g[379];
assign g[890] = b[8] & g[379];
assign g[636] = a[8] & g[380];
assign g[891] = b[8] & g[380];
assign g[637] = a[8] & g[381];
assign g[892] = b[8] & g[381];
assign g[638] = a[8] & g[382];
assign g[893] = b[8] & g[382];
assign g[639] = a[8] & g[383];
assign g[894] = b[8] & g[383];
assign g[640] = a[8] & g[384];
assign g[895] = b[8] & g[384];
assign g[641] = a[8] & g[385];
assign g[896] = b[8] & g[385];
assign g[642] = a[8] & g[386];
assign g[897] = b[8] & g[386];
assign g[643] = a[8] & g[387];
assign g[898] = b[8] & g[387];
assign g[644] = a[8] & g[388];
assign g[899] = b[8] & g[388];
assign g[645] = a[8] & g[389];
assign g[900] = b[8] & g[389];
assign g[646] = a[8] & g[390];
assign g[901] = b[8] & g[390];
assign g[647] = a[8] & g[391];
assign g[902] = b[8] & g[391];
assign g[648] = a[8] & g[392];
assign g[903] = b[8] & g[392];
assign g[649] = a[8] & g[393];
assign g[904] = b[8] & g[393];
assign g[650] = a[8] & g[394];
assign g[905] = b[8] & g[394];
assign g[651] = a[8] & g[395];
assign g[906] = b[8] & g[395];
assign g[652] = a[8] & g[396];
assign g[907] = b[8] & g[396];
assign g[653] = a[8] & g[397];
assign g[908] = b[8] & g[397];
assign g[654] = a[8] & g[398];
assign g[909] = b[8] & g[398];
assign g[655] = a[8] & g[399];
assign g[910] = b[8] & g[399];
assign g[656] = a[8] & g[400];
assign g[911] = b[8] & g[400];
assign g[657] = a[8] & g[401];
assign g[912] = b[8] & g[401];
assign g[658] = a[8] & g[402];
assign g[913] = b[8] & g[402];
assign g[659] = a[8] & g[403];
assign g[914] = b[8] & g[403];
assign g[660] = a[8] & g[404];
assign g[915] = b[8] & g[404];
assign g[661] = a[8] & g[405];
assign g[916] = b[8] & g[405];
assign g[662] = a[8] & g[406];
assign g[917] = b[8] & g[406];
assign g[663] = a[8] & g[407];
assign g[918] = b[8] & g[407];
assign g[664] = a[8] & g[408];
assign g[919] = b[8] & g[408];
assign g[665] = a[8] & g[409];
assign g[920] = b[8] & g[409];
assign g[666] = a[8] & g[410];
assign g[921] = b[8] & g[410];
assign g[667] = a[8] & g[411];
assign g[922] = b[8] & g[411];
assign g[668] = a[8] & g[412];
assign g[923] = b[8] & g[412];
assign g[669] = a[8] & g[413];
assign g[924] = b[8] & g[413];
assign g[670] = a[8] & g[414];
assign g[925] = b[8] & g[414];
assign g[671] = a[8] & g[415];
assign g[926] = b[8] & g[415];
assign g[672] = a[8] & g[416];
assign g[927] = b[8] & g[416];
assign g[673] = a[8] & g[417];
assign g[928] = b[8] & g[417];
assign g[674] = a[8] & g[418];
assign g[929] = b[8] & g[418];
assign g[675] = a[8] & g[419];
assign g[930] = b[8] & g[419];
assign g[676] = a[8] & g[420];
assign g[931] = b[8] & g[420];
assign g[677] = a[8] & g[421];
assign g[932] = b[8] & g[421];
assign g[678] = a[8] & g[422];
assign g[933] = b[8] & g[422];
assign g[679] = a[8] & g[423];
assign g[934] = b[8] & g[423];
assign g[680] = a[8] & g[424];
assign g[935] = b[8] & g[424];
assign g[681] = a[8] & g[425];
assign g[936] = b[8] & g[425];
assign g[682] = a[8] & g[426];
assign g[937] = b[8] & g[426];
assign g[683] = a[8] & g[427];
assign g[938] = b[8] & g[427];
assign g[684] = a[8] & g[428];
assign g[939] = b[8] & g[428];
assign g[685] = a[8] & g[429];
assign g[940] = b[8] & g[429];
assign g[686] = a[8] & g[430];
assign g[941] = b[8] & g[430];
assign g[687] = a[8] & g[431];
assign g[942] = b[8] & g[431];
assign g[688] = a[8] & g[432];
assign g[943] = b[8] & g[432];
assign g[689] = a[8] & g[433];
assign g[944] = b[8] & g[433];
assign g[690] = a[8] & g[434];
assign g[945] = b[8] & g[434];
assign g[691] = a[8] & g[435];
assign g[946] = b[8] & g[435];
assign g[692] = a[8] & g[436];
assign g[947] = b[8] & g[436];
assign g[693] = a[8] & g[437];
assign g[948] = b[8] & g[437];
assign g[694] = a[8] & g[438];
assign g[949] = b[8] & g[438];
assign g[695] = a[8] & g[439];
assign g[950] = b[8] & g[439];
assign g[696] = a[8] & g[440];
assign g[951] = b[8] & g[440];
assign g[697] = a[8] & g[441];
assign g[952] = b[8] & g[441];
assign g[698] = a[8] & g[442];
assign g[953] = b[8] & g[442];
assign g[699] = a[8] & g[443];
assign g[954] = b[8] & g[443];
assign g[700] = a[8] & g[444];
assign g[955] = b[8] & g[444];
assign g[701] = a[8] & g[445];
assign g[956] = b[8] & g[445];
assign g[702] = a[8] & g[446];
assign g[957] = b[8] & g[446];
assign g[703] = a[8] & g[447];
assign g[958] = b[8] & g[447];
assign g[704] = a[8] & g[448];
assign g[959] = b[8] & g[448];
assign g[705] = a[8] & g[449];
assign g[960] = b[8] & g[449];
assign g[706] = a[8] & g[450];
assign g[961] = b[8] & g[450];
assign g[707] = a[8] & g[451];
assign g[962] = b[8] & g[451];
assign g[708] = a[8] & g[452];
assign g[963] = b[8] & g[452];
assign g[709] = a[8] & g[453];
assign g[964] = b[8] & g[453];
assign g[710] = a[8] & g[454];
assign g[965] = b[8] & g[454];
assign g[711] = a[8] & g[455];
assign g[966] = b[8] & g[455];
assign g[712] = a[8] & g[456];
assign g[967] = b[8] & g[456];
assign g[713] = a[8] & g[457];
assign g[968] = b[8] & g[457];
assign g[714] = a[8] & g[458];
assign g[969] = b[8] & g[458];
assign g[715] = a[8] & g[459];
assign g[970] = b[8] & g[459];
assign g[716] = a[8] & g[460];
assign g[971] = b[8] & g[460];
assign g[717] = a[8] & g[461];
assign g[972] = b[8] & g[461];
assign g[718] = a[8] & g[462];
assign g[973] = b[8] & g[462];
assign g[719] = a[8] & g[463];
assign g[974] = b[8] & g[463];
assign g[720] = a[8] & g[464];
assign g[975] = b[8] & g[464];
assign g[721] = a[8] & g[465];
assign g[976] = b[8] & g[465];
assign g[722] = a[8] & g[466];
assign g[977] = b[8] & g[466];
assign g[723] = a[8] & g[467];
assign g[978] = b[8] & g[467];
assign g[724] = a[8] & g[468];
assign g[979] = b[8] & g[468];
assign g[725] = a[8] & g[469];
assign g[980] = b[8] & g[469];
assign g[726] = a[8] & g[470];
assign g[981] = b[8] & g[470];
assign g[727] = a[8] & g[471];
assign g[982] = b[8] & g[471];
assign g[728] = a[8] & g[472];
assign g[983] = b[8] & g[472];
assign g[729] = a[8] & g[473];
assign g[984] = b[8] & g[473];
assign g[730] = a[8] & g[474];
assign g[985] = b[8] & g[474];
assign g[731] = a[8] & g[475];
assign g[986] = b[8] & g[475];
assign g[732] = a[8] & g[476];
assign g[987] = b[8] & g[476];
assign g[733] = a[8] & g[477];
assign g[988] = b[8] & g[477];
assign g[734] = a[8] & g[478];
assign g[989] = b[8] & g[478];
assign g[735] = a[8] & g[479];
assign g[990] = b[8] & g[479];
assign g[736] = a[8] & g[480];
assign g[991] = b[8] & g[480];
assign g[737] = a[8] & g[481];
assign g[992] = b[8] & g[481];
assign g[738] = a[8] & g[482];
assign g[993] = b[8] & g[482];
assign g[739] = a[8] & g[483];
assign g[994] = b[8] & g[483];
assign g[740] = a[8] & g[484];
assign g[995] = b[8] & g[484];
assign g[741] = a[8] & g[485];
assign g[996] = b[8] & g[485];
assign g[742] = a[8] & g[486];
assign g[997] = b[8] & g[486];
assign g[743] = a[8] & g[487];
assign g[998] = b[8] & g[487];
assign g[744] = a[8] & g[488];
assign g[999] = b[8] & g[488];
assign g[745] = a[8] & g[489];
assign g[1000] = b[8] & g[489];
assign g[746] = a[8] & g[490];
assign g[1001] = b[8] & g[490];
assign g[747] = a[8] & g[491];
assign g[1002] = b[8] & g[491];
assign g[748] = a[8] & g[492];
assign g[1003] = b[8] & g[492];
assign g[749] = a[8] & g[493];
assign g[1004] = b[8] & g[493];
assign g[750] = a[8] & g[494];
assign g[1005] = b[8] & g[494];
assign g[751] = a[8] & g[495];
assign g[1006] = b[8] & g[495];
assign g[752] = a[8] & g[496];
assign g[1007] = b[8] & g[496];
assign g[753] = a[8] & g[497];
assign g[1008] = b[8] & g[497];
assign g[754] = a[8] & g[498];
assign g[1009] = b[8] & g[498];
assign g[755] = a[8] & g[499];
assign g[1010] = b[8] & g[499];
assign g[756] = a[8] & g[500];
assign g[1011] = b[8] & g[500];
assign g[757] = a[8] & g[501];
assign g[1012] = b[8] & g[501];
//Assigning outputs for input bit 10
assign g[1013] = a[9] & b[9];
assign g[1014] = a[9] & g[502];
assign g[1525] = b[9] & g[502];
assign g[1015] = a[9] & g[503];
assign g[1526] = b[9] & g[503];
assign g[1016] = a[9] & g[504];
assign g[1527] = b[9] & g[504];
assign g[1017] = a[9] & g[505];
assign g[1528] = b[9] & g[505];
assign g[1018] = a[9] & g[506];
assign g[1529] = b[9] & g[506];
assign g[1019] = a[9] & g[507];
assign g[1530] = b[9] & g[507];
assign g[1020] = a[9] & g[508];
assign g[1531] = b[9] & g[508];
assign g[1021] = a[9] & g[509];
assign g[1532] = b[9] & g[509];
assign g[1022] = a[9] & g[510];
assign g[1533] = b[9] & g[510];
assign g[1023] = a[9] & g[511];
assign g[1534] = b[9] & g[511];
assign g[1024] = a[9] & g[512];
assign g[1535] = b[9] & g[512];
assign g[1025] = a[9] & g[513];
assign g[1536] = b[9] & g[513];
assign g[1026] = a[9] & g[514];
assign g[1537] = b[9] & g[514];
assign g[1027] = a[9] & g[515];
assign g[1538] = b[9] & g[515];
assign g[1028] = a[9] & g[516];
assign g[1539] = b[9] & g[516];
assign g[1029] = a[9] & g[517];
assign g[1540] = b[9] & g[517];
assign g[1030] = a[9] & g[518];
assign g[1541] = b[9] & g[518];
assign g[1031] = a[9] & g[519];
assign g[1542] = b[9] & g[519];
assign g[1032] = a[9] & g[520];
assign g[1543] = b[9] & g[520];
assign g[1033] = a[9] & g[521];
assign g[1544] = b[9] & g[521];
assign g[1034] = a[9] & g[522];
assign g[1545] = b[9] & g[522];
assign g[1035] = a[9] & g[523];
assign g[1546] = b[9] & g[523];
assign g[1036] = a[9] & g[524];
assign g[1547] = b[9] & g[524];
assign g[1037] = a[9] & g[525];
assign g[1548] = b[9] & g[525];
assign g[1038] = a[9] & g[526];
assign g[1549] = b[9] & g[526];
assign g[1039] = a[9] & g[527];
assign g[1550] = b[9] & g[527];
assign g[1040] = a[9] & g[528];
assign g[1551] = b[9] & g[528];
assign g[1041] = a[9] & g[529];
assign g[1552] = b[9] & g[529];
assign g[1042] = a[9] & g[530];
assign g[1553] = b[9] & g[530];
assign g[1043] = a[9] & g[531];
assign g[1554] = b[9] & g[531];
assign g[1044] = a[9] & g[532];
assign g[1555] = b[9] & g[532];
assign g[1045] = a[9] & g[533];
assign g[1556] = b[9] & g[533];
assign g[1046] = a[9] & g[534];
assign g[1557] = b[9] & g[534];
assign g[1047] = a[9] & g[535];
assign g[1558] = b[9] & g[535];
assign g[1048] = a[9] & g[536];
assign g[1559] = b[9] & g[536];
assign g[1049] = a[9] & g[537];
assign g[1560] = b[9] & g[537];
assign g[1050] = a[9] & g[538];
assign g[1561] = b[9] & g[538];
assign g[1051] = a[9] & g[539];
assign g[1562] = b[9] & g[539];
assign g[1052] = a[9] & g[540];
assign g[1563] = b[9] & g[540];
assign g[1053] = a[9] & g[541];
assign g[1564] = b[9] & g[541];
assign g[1054] = a[9] & g[542];
assign g[1565] = b[9] & g[542];
assign g[1055] = a[9] & g[543];
assign g[1566] = b[9] & g[543];
assign g[1056] = a[9] & g[544];
assign g[1567] = b[9] & g[544];
assign g[1057] = a[9] & g[545];
assign g[1568] = b[9] & g[545];
assign g[1058] = a[9] & g[546];
assign g[1569] = b[9] & g[546];
assign g[1059] = a[9] & g[547];
assign g[1570] = b[9] & g[547];
assign g[1060] = a[9] & g[548];
assign g[1571] = b[9] & g[548];
assign g[1061] = a[9] & g[549];
assign g[1572] = b[9] & g[549];
assign g[1062] = a[9] & g[550];
assign g[1573] = b[9] & g[550];
assign g[1063] = a[9] & g[551];
assign g[1574] = b[9] & g[551];
assign g[1064] = a[9] & g[552];
assign g[1575] = b[9] & g[552];
assign g[1065] = a[9] & g[553];
assign g[1576] = b[9] & g[553];
assign g[1066] = a[9] & g[554];
assign g[1577] = b[9] & g[554];
assign g[1067] = a[9] & g[555];
assign g[1578] = b[9] & g[555];
assign g[1068] = a[9] & g[556];
assign g[1579] = b[9] & g[556];
assign g[1069] = a[9] & g[557];
assign g[1580] = b[9] & g[557];
assign g[1070] = a[9] & g[558];
assign g[1581] = b[9] & g[558];
assign g[1071] = a[9] & g[559];
assign g[1582] = b[9] & g[559];
assign g[1072] = a[9] & g[560];
assign g[1583] = b[9] & g[560];
assign g[1073] = a[9] & g[561];
assign g[1584] = b[9] & g[561];
assign g[1074] = a[9] & g[562];
assign g[1585] = b[9] & g[562];
assign g[1075] = a[9] & g[563];
assign g[1586] = b[9] & g[563];
assign g[1076] = a[9] & g[564];
assign g[1587] = b[9] & g[564];
assign g[1077] = a[9] & g[565];
assign g[1588] = b[9] & g[565];
assign g[1078] = a[9] & g[566];
assign g[1589] = b[9] & g[566];
assign g[1079] = a[9] & g[567];
assign g[1590] = b[9] & g[567];
assign g[1080] = a[9] & g[568];
assign g[1591] = b[9] & g[568];
assign g[1081] = a[9] & g[569];
assign g[1592] = b[9] & g[569];
assign g[1082] = a[9] & g[570];
assign g[1593] = b[9] & g[570];
assign g[1083] = a[9] & g[571];
assign g[1594] = b[9] & g[571];
assign g[1084] = a[9] & g[572];
assign g[1595] = b[9] & g[572];
assign g[1085] = a[9] & g[573];
assign g[1596] = b[9] & g[573];
assign g[1086] = a[9] & g[574];
assign g[1597] = b[9] & g[574];
assign g[1087] = a[9] & g[575];
assign g[1598] = b[9] & g[575];
assign g[1088] = a[9] & g[576];
assign g[1599] = b[9] & g[576];
assign g[1089] = a[9] & g[577];
assign g[1600] = b[9] & g[577];
assign g[1090] = a[9] & g[578];
assign g[1601] = b[9] & g[578];
assign g[1091] = a[9] & g[579];
assign g[1602] = b[9] & g[579];
assign g[1092] = a[9] & g[580];
assign g[1603] = b[9] & g[580];
assign g[1093] = a[9] & g[581];
assign g[1604] = b[9] & g[581];
assign g[1094] = a[9] & g[582];
assign g[1605] = b[9] & g[582];
assign g[1095] = a[9] & g[583];
assign g[1606] = b[9] & g[583];
assign g[1096] = a[9] & g[584];
assign g[1607] = b[9] & g[584];
assign g[1097] = a[9] & g[585];
assign g[1608] = b[9] & g[585];
assign g[1098] = a[9] & g[586];
assign g[1609] = b[9] & g[586];
assign g[1099] = a[9] & g[587];
assign g[1610] = b[9] & g[587];
assign g[1100] = a[9] & g[588];
assign g[1611] = b[9] & g[588];
assign g[1101] = a[9] & g[589];
assign g[1612] = b[9] & g[589];
assign g[1102] = a[9] & g[590];
assign g[1613] = b[9] & g[590];
assign g[1103] = a[9] & g[591];
assign g[1614] = b[9] & g[591];
assign g[1104] = a[9] & g[592];
assign g[1615] = b[9] & g[592];
assign g[1105] = a[9] & g[593];
assign g[1616] = b[9] & g[593];
assign g[1106] = a[9] & g[594];
assign g[1617] = b[9] & g[594];
assign g[1107] = a[9] & g[595];
assign g[1618] = b[9] & g[595];
assign g[1108] = a[9] & g[596];
assign g[1619] = b[9] & g[596];
assign g[1109] = a[9] & g[597];
assign g[1620] = b[9] & g[597];
assign g[1110] = a[9] & g[598];
assign g[1621] = b[9] & g[598];
assign g[1111] = a[9] & g[599];
assign g[1622] = b[9] & g[599];
assign g[1112] = a[9] & g[600];
assign g[1623] = b[9] & g[600];
assign g[1113] = a[9] & g[601];
assign g[1624] = b[9] & g[601];
assign g[1114] = a[9] & g[602];
assign g[1625] = b[9] & g[602];
assign g[1115] = a[9] & g[603];
assign g[1626] = b[9] & g[603];
assign g[1116] = a[9] & g[604];
assign g[1627] = b[9] & g[604];
assign g[1117] = a[9] & g[605];
assign g[1628] = b[9] & g[605];
assign g[1118] = a[9] & g[606];
assign g[1629] = b[9] & g[606];
assign g[1119] = a[9] & g[607];
assign g[1630] = b[9] & g[607];
assign g[1120] = a[9] & g[608];
assign g[1631] = b[9] & g[608];
assign g[1121] = a[9] & g[609];
assign g[1632] = b[9] & g[609];
assign g[1122] = a[9] & g[610];
assign g[1633] = b[9] & g[610];
assign g[1123] = a[9] & g[611];
assign g[1634] = b[9] & g[611];
assign g[1124] = a[9] & g[612];
assign g[1635] = b[9] & g[612];
assign g[1125] = a[9] & g[613];
assign g[1636] = b[9] & g[613];
assign g[1126] = a[9] & g[614];
assign g[1637] = b[9] & g[614];
assign g[1127] = a[9] & g[615];
assign g[1638] = b[9] & g[615];
assign g[1128] = a[9] & g[616];
assign g[1639] = b[9] & g[616];
assign g[1129] = a[9] & g[617];
assign g[1640] = b[9] & g[617];
assign g[1130] = a[9] & g[618];
assign g[1641] = b[9] & g[618];
assign g[1131] = a[9] & g[619];
assign g[1642] = b[9] & g[619];
assign g[1132] = a[9] & g[620];
assign g[1643] = b[9] & g[620];
assign g[1133] = a[9] & g[621];
assign g[1644] = b[9] & g[621];
assign g[1134] = a[9] & g[622];
assign g[1645] = b[9] & g[622];
assign g[1135] = a[9] & g[623];
assign g[1646] = b[9] & g[623];
assign g[1136] = a[9] & g[624];
assign g[1647] = b[9] & g[624];
assign g[1137] = a[9] & g[625];
assign g[1648] = b[9] & g[625];
assign g[1138] = a[9] & g[626];
assign g[1649] = b[9] & g[626];
assign g[1139] = a[9] & g[627];
assign g[1650] = b[9] & g[627];
assign g[1140] = a[9] & g[628];
assign g[1651] = b[9] & g[628];
assign g[1141] = a[9] & g[629];
assign g[1652] = b[9] & g[629];
assign g[1142] = a[9] & g[630];
assign g[1653] = b[9] & g[630];
assign g[1143] = a[9] & g[631];
assign g[1654] = b[9] & g[631];
assign g[1144] = a[9] & g[632];
assign g[1655] = b[9] & g[632];
assign g[1145] = a[9] & g[633];
assign g[1656] = b[9] & g[633];
assign g[1146] = a[9] & g[634];
assign g[1657] = b[9] & g[634];
assign g[1147] = a[9] & g[635];
assign g[1658] = b[9] & g[635];
assign g[1148] = a[9] & g[636];
assign g[1659] = b[9] & g[636];
assign g[1149] = a[9] & g[637];
assign g[1660] = b[9] & g[637];
assign g[1150] = a[9] & g[638];
assign g[1661] = b[9] & g[638];
assign g[1151] = a[9] & g[639];
assign g[1662] = b[9] & g[639];
assign g[1152] = a[9] & g[640];
assign g[1663] = b[9] & g[640];
assign g[1153] = a[9] & g[641];
assign g[1664] = b[9] & g[641];
assign g[1154] = a[9] & g[642];
assign g[1665] = b[9] & g[642];
assign g[1155] = a[9] & g[643];
assign g[1666] = b[9] & g[643];
assign g[1156] = a[9] & g[644];
assign g[1667] = b[9] & g[644];
assign g[1157] = a[9] & g[645];
assign g[1668] = b[9] & g[645];
assign g[1158] = a[9] & g[646];
assign g[1669] = b[9] & g[646];
assign g[1159] = a[9] & g[647];
assign g[1670] = b[9] & g[647];
assign g[1160] = a[9] & g[648];
assign g[1671] = b[9] & g[648];
assign g[1161] = a[9] & g[649];
assign g[1672] = b[9] & g[649];
assign g[1162] = a[9] & g[650];
assign g[1673] = b[9] & g[650];
assign g[1163] = a[9] & g[651];
assign g[1674] = b[9] & g[651];
assign g[1164] = a[9] & g[652];
assign g[1675] = b[9] & g[652];
assign g[1165] = a[9] & g[653];
assign g[1676] = b[9] & g[653];
assign g[1166] = a[9] & g[654];
assign g[1677] = b[9] & g[654];
assign g[1167] = a[9] & g[655];
assign g[1678] = b[9] & g[655];
assign g[1168] = a[9] & g[656];
assign g[1679] = b[9] & g[656];
assign g[1169] = a[9] & g[657];
assign g[1680] = b[9] & g[657];
assign g[1170] = a[9] & g[658];
assign g[1681] = b[9] & g[658];
assign g[1171] = a[9] & g[659];
assign g[1682] = b[9] & g[659];
assign g[1172] = a[9] & g[660];
assign g[1683] = b[9] & g[660];
assign g[1173] = a[9] & g[661];
assign g[1684] = b[9] & g[661];
assign g[1174] = a[9] & g[662];
assign g[1685] = b[9] & g[662];
assign g[1175] = a[9] & g[663];
assign g[1686] = b[9] & g[663];
assign g[1176] = a[9] & g[664];
assign g[1687] = b[9] & g[664];
assign g[1177] = a[9] & g[665];
assign g[1688] = b[9] & g[665];
assign g[1178] = a[9] & g[666];
assign g[1689] = b[9] & g[666];
assign g[1179] = a[9] & g[667];
assign g[1690] = b[9] & g[667];
assign g[1180] = a[9] & g[668];
assign g[1691] = b[9] & g[668];
assign g[1181] = a[9] & g[669];
assign g[1692] = b[9] & g[669];
assign g[1182] = a[9] & g[670];
assign g[1693] = b[9] & g[670];
assign g[1183] = a[9] & g[671];
assign g[1694] = b[9] & g[671];
assign g[1184] = a[9] & g[672];
assign g[1695] = b[9] & g[672];
assign g[1185] = a[9] & g[673];
assign g[1696] = b[9] & g[673];
assign g[1186] = a[9] & g[674];
assign g[1697] = b[9] & g[674];
assign g[1187] = a[9] & g[675];
assign g[1698] = b[9] & g[675];
assign g[1188] = a[9] & g[676];
assign g[1699] = b[9] & g[676];
assign g[1189] = a[9] & g[677];
assign g[1700] = b[9] & g[677];
assign g[1190] = a[9] & g[678];
assign g[1701] = b[9] & g[678];
assign g[1191] = a[9] & g[679];
assign g[1702] = b[9] & g[679];
assign g[1192] = a[9] & g[680];
assign g[1703] = b[9] & g[680];
assign g[1193] = a[9] & g[681];
assign g[1704] = b[9] & g[681];
assign g[1194] = a[9] & g[682];
assign g[1705] = b[9] & g[682];
assign g[1195] = a[9] & g[683];
assign g[1706] = b[9] & g[683];
assign g[1196] = a[9] & g[684];
assign g[1707] = b[9] & g[684];
assign g[1197] = a[9] & g[685];
assign g[1708] = b[9] & g[685];
assign g[1198] = a[9] & g[686];
assign g[1709] = b[9] & g[686];
assign g[1199] = a[9] & g[687];
assign g[1710] = b[9] & g[687];
assign g[1200] = a[9] & g[688];
assign g[1711] = b[9] & g[688];
assign g[1201] = a[9] & g[689];
assign g[1712] = b[9] & g[689];
assign g[1202] = a[9] & g[690];
assign g[1713] = b[9] & g[690];
assign g[1203] = a[9] & g[691];
assign g[1714] = b[9] & g[691];
assign g[1204] = a[9] & g[692];
assign g[1715] = b[9] & g[692];
assign g[1205] = a[9] & g[693];
assign g[1716] = b[9] & g[693];
assign g[1206] = a[9] & g[694];
assign g[1717] = b[9] & g[694];
assign g[1207] = a[9] & g[695];
assign g[1718] = b[9] & g[695];
assign g[1208] = a[9] & g[696];
assign g[1719] = b[9] & g[696];
assign g[1209] = a[9] & g[697];
assign g[1720] = b[9] & g[697];
assign g[1210] = a[9] & g[698];
assign g[1721] = b[9] & g[698];
assign g[1211] = a[9] & g[699];
assign g[1722] = b[9] & g[699];
assign g[1212] = a[9] & g[700];
assign g[1723] = b[9] & g[700];
assign g[1213] = a[9] & g[701];
assign g[1724] = b[9] & g[701];
assign g[1214] = a[9] & g[702];
assign g[1725] = b[9] & g[702];
assign g[1215] = a[9] & g[703];
assign g[1726] = b[9] & g[703];
assign g[1216] = a[9] & g[704];
assign g[1727] = b[9] & g[704];
assign g[1217] = a[9] & g[705];
assign g[1728] = b[9] & g[705];
assign g[1218] = a[9] & g[706];
assign g[1729] = b[9] & g[706];
assign g[1219] = a[9] & g[707];
assign g[1730] = b[9] & g[707];
assign g[1220] = a[9] & g[708];
assign g[1731] = b[9] & g[708];
assign g[1221] = a[9] & g[709];
assign g[1732] = b[9] & g[709];
assign g[1222] = a[9] & g[710];
assign g[1733] = b[9] & g[710];
assign g[1223] = a[9] & g[711];
assign g[1734] = b[9] & g[711];
assign g[1224] = a[9] & g[712];
assign g[1735] = b[9] & g[712];
assign g[1225] = a[9] & g[713];
assign g[1736] = b[9] & g[713];
assign g[1226] = a[9] & g[714];
assign g[1737] = b[9] & g[714];
assign g[1227] = a[9] & g[715];
assign g[1738] = b[9] & g[715];
assign g[1228] = a[9] & g[716];
assign g[1739] = b[9] & g[716];
assign g[1229] = a[9] & g[717];
assign g[1740] = b[9] & g[717];
assign g[1230] = a[9] & g[718];
assign g[1741] = b[9] & g[718];
assign g[1231] = a[9] & g[719];
assign g[1742] = b[9] & g[719];
assign g[1232] = a[9] & g[720];
assign g[1743] = b[9] & g[720];
assign g[1233] = a[9] & g[721];
assign g[1744] = b[9] & g[721];
assign g[1234] = a[9] & g[722];
assign g[1745] = b[9] & g[722];
assign g[1235] = a[9] & g[723];
assign g[1746] = b[9] & g[723];
assign g[1236] = a[9] & g[724];
assign g[1747] = b[9] & g[724];
assign g[1237] = a[9] & g[725];
assign g[1748] = b[9] & g[725];
assign g[1238] = a[9] & g[726];
assign g[1749] = b[9] & g[726];
assign g[1239] = a[9] & g[727];
assign g[1750] = b[9] & g[727];
assign g[1240] = a[9] & g[728];
assign g[1751] = b[9] & g[728];
assign g[1241] = a[9] & g[729];
assign g[1752] = b[9] & g[729];
assign g[1242] = a[9] & g[730];
assign g[1753] = b[9] & g[730];
assign g[1243] = a[9] & g[731];
assign g[1754] = b[9] & g[731];
assign g[1244] = a[9] & g[732];
assign g[1755] = b[9] & g[732];
assign g[1245] = a[9] & g[733];
assign g[1756] = b[9] & g[733];
assign g[1246] = a[9] & g[734];
assign g[1757] = b[9] & g[734];
assign g[1247] = a[9] & g[735];
assign g[1758] = b[9] & g[735];
assign g[1248] = a[9] & g[736];
assign g[1759] = b[9] & g[736];
assign g[1249] = a[9] & g[737];
assign g[1760] = b[9] & g[737];
assign g[1250] = a[9] & g[738];
assign g[1761] = b[9] & g[738];
assign g[1251] = a[9] & g[739];
assign g[1762] = b[9] & g[739];
assign g[1252] = a[9] & g[740];
assign g[1763] = b[9] & g[740];
assign g[1253] = a[9] & g[741];
assign g[1764] = b[9] & g[741];
assign g[1254] = a[9] & g[742];
assign g[1765] = b[9] & g[742];
assign g[1255] = a[9] & g[743];
assign g[1766] = b[9] & g[743];
assign g[1256] = a[9] & g[744];
assign g[1767] = b[9] & g[744];
assign g[1257] = a[9] & g[745];
assign g[1768] = b[9] & g[745];
assign g[1258] = a[9] & g[746];
assign g[1769] = b[9] & g[746];
assign g[1259] = a[9] & g[747];
assign g[1770] = b[9] & g[747];
assign g[1260] = a[9] & g[748];
assign g[1771] = b[9] & g[748];
assign g[1261] = a[9] & g[749];
assign g[1772] = b[9] & g[749];
assign g[1262] = a[9] & g[750];
assign g[1773] = b[9] & g[750];
assign g[1263] = a[9] & g[751];
assign g[1774] = b[9] & g[751];
assign g[1264] = a[9] & g[752];
assign g[1775] = b[9] & g[752];
assign g[1265] = a[9] & g[753];
assign g[1776] = b[9] & g[753];
assign g[1266] = a[9] & g[754];
assign g[1777] = b[9] & g[754];
assign g[1267] = a[9] & g[755];
assign g[1778] = b[9] & g[755];
assign g[1268] = a[9] & g[756];
assign g[1779] = b[9] & g[756];
assign g[1269] = a[9] & g[757];
assign g[1780] = b[9] & g[757];
assign g[1270] = a[9] & g[758];
assign g[1781] = b[9] & g[758];
assign g[1271] = a[9] & g[759];
assign g[1782] = b[9] & g[759];
assign g[1272] = a[9] & g[760];
assign g[1783] = b[9] & g[760];
assign g[1273] = a[9] & g[761];
assign g[1784] = b[9] & g[761];
assign g[1274] = a[9] & g[762];
assign g[1785] = b[9] & g[762];
assign g[1275] = a[9] & g[763];
assign g[1786] = b[9] & g[763];
assign g[1276] = a[9] & g[764];
assign g[1787] = b[9] & g[764];
assign g[1277] = a[9] & g[765];
assign g[1788] = b[9] & g[765];
assign g[1278] = a[9] & g[766];
assign g[1789] = b[9] & g[766];
assign g[1279] = a[9] & g[767];
assign g[1790] = b[9] & g[767];
assign g[1280] = a[9] & g[768];
assign g[1791] = b[9] & g[768];
assign g[1281] = a[9] & g[769];
assign g[1792] = b[9] & g[769];
assign g[1282] = a[9] & g[770];
assign g[1793] = b[9] & g[770];
assign g[1283] = a[9] & g[771];
assign g[1794] = b[9] & g[771];
assign g[1284] = a[9] & g[772];
assign g[1795] = b[9] & g[772];
assign g[1285] = a[9] & g[773];
assign g[1796] = b[9] & g[773];
assign g[1286] = a[9] & g[774];
assign g[1797] = b[9] & g[774];
assign g[1287] = a[9] & g[775];
assign g[1798] = b[9] & g[775];
assign g[1288] = a[9] & g[776];
assign g[1799] = b[9] & g[776];
assign g[1289] = a[9] & g[777];
assign g[1800] = b[9] & g[777];
assign g[1290] = a[9] & g[778];
assign g[1801] = b[9] & g[778];
assign g[1291] = a[9] & g[779];
assign g[1802] = b[9] & g[779];
assign g[1292] = a[9] & g[780];
assign g[1803] = b[9] & g[780];
assign g[1293] = a[9] & g[781];
assign g[1804] = b[9] & g[781];
assign g[1294] = a[9] & g[782];
assign g[1805] = b[9] & g[782];
assign g[1295] = a[9] & g[783];
assign g[1806] = b[9] & g[783];
assign g[1296] = a[9] & g[784];
assign g[1807] = b[9] & g[784];
assign g[1297] = a[9] & g[785];
assign g[1808] = b[9] & g[785];
assign g[1298] = a[9] & g[786];
assign g[1809] = b[9] & g[786];
assign g[1299] = a[9] & g[787];
assign g[1810] = b[9] & g[787];
assign g[1300] = a[9] & g[788];
assign g[1811] = b[9] & g[788];
assign g[1301] = a[9] & g[789];
assign g[1812] = b[9] & g[789];
assign g[1302] = a[9] & g[790];
assign g[1813] = b[9] & g[790];
assign g[1303] = a[9] & g[791];
assign g[1814] = b[9] & g[791];
assign g[1304] = a[9] & g[792];
assign g[1815] = b[9] & g[792];
assign g[1305] = a[9] & g[793];
assign g[1816] = b[9] & g[793];
assign g[1306] = a[9] & g[794];
assign g[1817] = b[9] & g[794];
assign g[1307] = a[9] & g[795];
assign g[1818] = b[9] & g[795];
assign g[1308] = a[9] & g[796];
assign g[1819] = b[9] & g[796];
assign g[1309] = a[9] & g[797];
assign g[1820] = b[9] & g[797];
assign g[1310] = a[9] & g[798];
assign g[1821] = b[9] & g[798];
assign g[1311] = a[9] & g[799];
assign g[1822] = b[9] & g[799];
assign g[1312] = a[9] & g[800];
assign g[1823] = b[9] & g[800];
assign g[1313] = a[9] & g[801];
assign g[1824] = b[9] & g[801];
assign g[1314] = a[9] & g[802];
assign g[1825] = b[9] & g[802];
assign g[1315] = a[9] & g[803];
assign g[1826] = b[9] & g[803];
assign g[1316] = a[9] & g[804];
assign g[1827] = b[9] & g[804];
assign g[1317] = a[9] & g[805];
assign g[1828] = b[9] & g[805];
assign g[1318] = a[9] & g[806];
assign g[1829] = b[9] & g[806];
assign g[1319] = a[9] & g[807];
assign g[1830] = b[9] & g[807];
assign g[1320] = a[9] & g[808];
assign g[1831] = b[9] & g[808];
assign g[1321] = a[9] & g[809];
assign g[1832] = b[9] & g[809];
assign g[1322] = a[9] & g[810];
assign g[1833] = b[9] & g[810];
assign g[1323] = a[9] & g[811];
assign g[1834] = b[9] & g[811];
assign g[1324] = a[9] & g[812];
assign g[1835] = b[9] & g[812];
assign g[1325] = a[9] & g[813];
assign g[1836] = b[9] & g[813];
assign g[1326] = a[9] & g[814];
assign g[1837] = b[9] & g[814];
assign g[1327] = a[9] & g[815];
assign g[1838] = b[9] & g[815];
assign g[1328] = a[9] & g[816];
assign g[1839] = b[9] & g[816];
assign g[1329] = a[9] & g[817];
assign g[1840] = b[9] & g[817];
assign g[1330] = a[9] & g[818];
assign g[1841] = b[9] & g[818];
assign g[1331] = a[9] & g[819];
assign g[1842] = b[9] & g[819];
assign g[1332] = a[9] & g[820];
assign g[1843] = b[9] & g[820];
assign g[1333] = a[9] & g[821];
assign g[1844] = b[9] & g[821];
assign g[1334] = a[9] & g[822];
assign g[1845] = b[9] & g[822];
assign g[1335] = a[9] & g[823];
assign g[1846] = b[9] & g[823];
assign g[1336] = a[9] & g[824];
assign g[1847] = b[9] & g[824];
assign g[1337] = a[9] & g[825];
assign g[1848] = b[9] & g[825];
assign g[1338] = a[9] & g[826];
assign g[1849] = b[9] & g[826];
assign g[1339] = a[9] & g[827];
assign g[1850] = b[9] & g[827];
assign g[1340] = a[9] & g[828];
assign g[1851] = b[9] & g[828];
assign g[1341] = a[9] & g[829];
assign g[1852] = b[9] & g[829];
assign g[1342] = a[9] & g[830];
assign g[1853] = b[9] & g[830];
assign g[1343] = a[9] & g[831];
assign g[1854] = b[9] & g[831];
assign g[1344] = a[9] & g[832];
assign g[1855] = b[9] & g[832];
assign g[1345] = a[9] & g[833];
assign g[1856] = b[9] & g[833];
assign g[1346] = a[9] & g[834];
assign g[1857] = b[9] & g[834];
assign g[1347] = a[9] & g[835];
assign g[1858] = b[9] & g[835];
assign g[1348] = a[9] & g[836];
assign g[1859] = b[9] & g[836];
assign g[1349] = a[9] & g[837];
assign g[1860] = b[9] & g[837];
assign g[1350] = a[9] & g[838];
assign g[1861] = b[9] & g[838];
assign g[1351] = a[9] & g[839];
assign g[1862] = b[9] & g[839];
assign g[1352] = a[9] & g[840];
assign g[1863] = b[9] & g[840];
assign g[1353] = a[9] & g[841];
assign g[1864] = b[9] & g[841];
assign g[1354] = a[9] & g[842];
assign g[1865] = b[9] & g[842];
assign g[1355] = a[9] & g[843];
assign g[1866] = b[9] & g[843];
assign g[1356] = a[9] & g[844];
assign g[1867] = b[9] & g[844];
assign g[1357] = a[9] & g[845];
assign g[1868] = b[9] & g[845];
assign g[1358] = a[9] & g[846];
assign g[1869] = b[9] & g[846];
assign g[1359] = a[9] & g[847];
assign g[1870] = b[9] & g[847];
assign g[1360] = a[9] & g[848];
assign g[1871] = b[9] & g[848];
assign g[1361] = a[9] & g[849];
assign g[1872] = b[9] & g[849];
assign g[1362] = a[9] & g[850];
assign g[1873] = b[9] & g[850];
assign g[1363] = a[9] & g[851];
assign g[1874] = b[9] & g[851];
assign g[1364] = a[9] & g[852];
assign g[1875] = b[9] & g[852];
assign g[1365] = a[9] & g[853];
assign g[1876] = b[9] & g[853];
assign g[1366] = a[9] & g[854];
assign g[1877] = b[9] & g[854];
assign g[1367] = a[9] & g[855];
assign g[1878] = b[9] & g[855];
assign g[1368] = a[9] & g[856];
assign g[1879] = b[9] & g[856];
assign g[1369] = a[9] & g[857];
assign g[1880] = b[9] & g[857];
assign g[1370] = a[9] & g[858];
assign g[1881] = b[9] & g[858];
assign g[1371] = a[9] & g[859];
assign g[1882] = b[9] & g[859];
assign g[1372] = a[9] & g[860];
assign g[1883] = b[9] & g[860];
assign g[1373] = a[9] & g[861];
assign g[1884] = b[9] & g[861];
assign g[1374] = a[9] & g[862];
assign g[1885] = b[9] & g[862];
assign g[1375] = a[9] & g[863];
assign g[1886] = b[9] & g[863];
assign g[1376] = a[9] & g[864];
assign g[1887] = b[9] & g[864];
assign g[1377] = a[9] & g[865];
assign g[1888] = b[9] & g[865];
assign g[1378] = a[9] & g[866];
assign g[1889] = b[9] & g[866];
assign g[1379] = a[9] & g[867];
assign g[1890] = b[9] & g[867];
assign g[1380] = a[9] & g[868];
assign g[1891] = b[9] & g[868];
assign g[1381] = a[9] & g[869];
assign g[1892] = b[9] & g[869];
assign g[1382] = a[9] & g[870];
assign g[1893] = b[9] & g[870];
assign g[1383] = a[9] & g[871];
assign g[1894] = b[9] & g[871];
assign g[1384] = a[9] & g[872];
assign g[1895] = b[9] & g[872];
assign g[1385] = a[9] & g[873];
assign g[1896] = b[9] & g[873];
assign g[1386] = a[9] & g[874];
assign g[1897] = b[9] & g[874];
assign g[1387] = a[9] & g[875];
assign g[1898] = b[9] & g[875];
assign g[1388] = a[9] & g[876];
assign g[1899] = b[9] & g[876];
assign g[1389] = a[9] & g[877];
assign g[1900] = b[9] & g[877];
assign g[1390] = a[9] & g[878];
assign g[1901] = b[9] & g[878];
assign g[1391] = a[9] & g[879];
assign g[1902] = b[9] & g[879];
assign g[1392] = a[9] & g[880];
assign g[1903] = b[9] & g[880];
assign g[1393] = a[9] & g[881];
assign g[1904] = b[9] & g[881];
assign g[1394] = a[9] & g[882];
assign g[1905] = b[9] & g[882];
assign g[1395] = a[9] & g[883];
assign g[1906] = b[9] & g[883];
assign g[1396] = a[9] & g[884];
assign g[1907] = b[9] & g[884];
assign g[1397] = a[9] & g[885];
assign g[1908] = b[9] & g[885];
assign g[1398] = a[9] & g[886];
assign g[1909] = b[9] & g[886];
assign g[1399] = a[9] & g[887];
assign g[1910] = b[9] & g[887];
assign g[1400] = a[9] & g[888];
assign g[1911] = b[9] & g[888];
assign g[1401] = a[9] & g[889];
assign g[1912] = b[9] & g[889];
assign g[1402] = a[9] & g[890];
assign g[1913] = b[9] & g[890];
assign g[1403] = a[9] & g[891];
assign g[1914] = b[9] & g[891];
assign g[1404] = a[9] & g[892];
assign g[1915] = b[9] & g[892];
assign g[1405] = a[9] & g[893];
assign g[1916] = b[9] & g[893];
assign g[1406] = a[9] & g[894];
assign g[1917] = b[9] & g[894];
assign g[1407] = a[9] & g[895];
assign g[1918] = b[9] & g[895];
assign g[1408] = a[9] & g[896];
assign g[1919] = b[9] & g[896];
assign g[1409] = a[9] & g[897];
assign g[1920] = b[9] & g[897];
assign g[1410] = a[9] & g[898];
assign g[1921] = b[9] & g[898];
assign g[1411] = a[9] & g[899];
assign g[1922] = b[9] & g[899];
assign g[1412] = a[9] & g[900];
assign g[1923] = b[9] & g[900];
assign g[1413] = a[9] & g[901];
assign g[1924] = b[9] & g[901];
assign g[1414] = a[9] & g[902];
assign g[1925] = b[9] & g[902];
assign g[1415] = a[9] & g[903];
assign g[1926] = b[9] & g[903];
assign g[1416] = a[9] & g[904];
assign g[1927] = b[9] & g[904];
assign g[1417] = a[9] & g[905];
assign g[1928] = b[9] & g[905];
assign g[1418] = a[9] & g[906];
assign g[1929] = b[9] & g[906];
assign g[1419] = a[9] & g[907];
assign g[1930] = b[9] & g[907];
assign g[1420] = a[9] & g[908];
assign g[1931] = b[9] & g[908];
assign g[1421] = a[9] & g[909];
assign g[1932] = b[9] & g[909];
assign g[1422] = a[9] & g[910];
assign g[1933] = b[9] & g[910];
assign g[1423] = a[9] & g[911];
assign g[1934] = b[9] & g[911];
assign g[1424] = a[9] & g[912];
assign g[1935] = b[9] & g[912];
assign g[1425] = a[9] & g[913];
assign g[1936] = b[9] & g[913];
assign g[1426] = a[9] & g[914];
assign g[1937] = b[9] & g[914];
assign g[1427] = a[9] & g[915];
assign g[1938] = b[9] & g[915];
assign g[1428] = a[9] & g[916];
assign g[1939] = b[9] & g[916];
assign g[1429] = a[9] & g[917];
assign g[1940] = b[9] & g[917];
assign g[1430] = a[9] & g[918];
assign g[1941] = b[9] & g[918];
assign g[1431] = a[9] & g[919];
assign g[1942] = b[9] & g[919];
assign g[1432] = a[9] & g[920];
assign g[1943] = b[9] & g[920];
assign g[1433] = a[9] & g[921];
assign g[1944] = b[9] & g[921];
assign g[1434] = a[9] & g[922];
assign g[1945] = b[9] & g[922];
assign g[1435] = a[9] & g[923];
assign g[1946] = b[9] & g[923];
assign g[1436] = a[9] & g[924];
assign g[1947] = b[9] & g[924];
assign g[1437] = a[9] & g[925];
assign g[1948] = b[9] & g[925];
assign g[1438] = a[9] & g[926];
assign g[1949] = b[9] & g[926];
assign g[1439] = a[9] & g[927];
assign g[1950] = b[9] & g[927];
assign g[1440] = a[9] & g[928];
assign g[1951] = b[9] & g[928];
assign g[1441] = a[9] & g[929];
assign g[1952] = b[9] & g[929];
assign g[1442] = a[9] & g[930];
assign g[1953] = b[9] & g[930];
assign g[1443] = a[9] & g[931];
assign g[1954] = b[9] & g[931];
assign g[1444] = a[9] & g[932];
assign g[1955] = b[9] & g[932];
assign g[1445] = a[9] & g[933];
assign g[1956] = b[9] & g[933];
assign g[1446] = a[9] & g[934];
assign g[1957] = b[9] & g[934];
assign g[1447] = a[9] & g[935];
assign g[1958] = b[9] & g[935];
assign g[1448] = a[9] & g[936];
assign g[1959] = b[9] & g[936];
assign g[1449] = a[9] & g[937];
assign g[1960] = b[9] & g[937];
assign g[1450] = a[9] & g[938];
assign g[1961] = b[9] & g[938];
assign g[1451] = a[9] & g[939];
assign g[1962] = b[9] & g[939];
assign g[1452] = a[9] & g[940];
assign g[1963] = b[9] & g[940];
assign g[1453] = a[9] & g[941];
assign g[1964] = b[9] & g[941];
assign g[1454] = a[9] & g[942];
assign g[1965] = b[9] & g[942];
assign g[1455] = a[9] & g[943];
assign g[1966] = b[9] & g[943];
assign g[1456] = a[9] & g[944];
assign g[1967] = b[9] & g[944];
assign g[1457] = a[9] & g[945];
assign g[1968] = b[9] & g[945];
assign g[1458] = a[9] & g[946];
assign g[1969] = b[9] & g[946];
assign g[1459] = a[9] & g[947];
assign g[1970] = b[9] & g[947];
assign g[1460] = a[9] & g[948];
assign g[1971] = b[9] & g[948];
assign g[1461] = a[9] & g[949];
assign g[1972] = b[9] & g[949];
assign g[1462] = a[9] & g[950];
assign g[1973] = b[9] & g[950];
assign g[1463] = a[9] & g[951];
assign g[1974] = b[9] & g[951];
assign g[1464] = a[9] & g[952];
assign g[1975] = b[9] & g[952];
assign g[1465] = a[9] & g[953];
assign g[1976] = b[9] & g[953];
assign g[1466] = a[9] & g[954];
assign g[1977] = b[9] & g[954];
assign g[1467] = a[9] & g[955];
assign g[1978] = b[9] & g[955];
assign g[1468] = a[9] & g[956];
assign g[1979] = b[9] & g[956];
assign g[1469] = a[9] & g[957];
assign g[1980] = b[9] & g[957];
assign g[1470] = a[9] & g[958];
assign g[1981] = b[9] & g[958];
assign g[1471] = a[9] & g[959];
assign g[1982] = b[9] & g[959];
assign g[1472] = a[9] & g[960];
assign g[1983] = b[9] & g[960];
assign g[1473] = a[9] & g[961];
assign g[1984] = b[9] & g[961];
assign g[1474] = a[9] & g[962];
assign g[1985] = b[9] & g[962];
assign g[1475] = a[9] & g[963];
assign g[1986] = b[9] & g[963];
assign g[1476] = a[9] & g[964];
assign g[1987] = b[9] & g[964];
assign g[1477] = a[9] & g[965];
assign g[1988] = b[9] & g[965];
assign g[1478] = a[9] & g[966];
assign g[1989] = b[9] & g[966];
assign g[1479] = a[9] & g[967];
assign g[1990] = b[9] & g[967];
assign g[1480] = a[9] & g[968];
assign g[1991] = b[9] & g[968];
assign g[1481] = a[9] & g[969];
assign g[1992] = b[9] & g[969];
assign g[1482] = a[9] & g[970];
assign g[1993] = b[9] & g[970];
assign g[1483] = a[9] & g[971];
assign g[1994] = b[9] & g[971];
assign g[1484] = a[9] & g[972];
assign g[1995] = b[9] & g[972];
assign g[1485] = a[9] & g[973];
assign g[1996] = b[9] & g[973];
assign g[1486] = a[9] & g[974];
assign g[1997] = b[9] & g[974];
assign g[1487] = a[9] & g[975];
assign g[1998] = b[9] & g[975];
assign g[1488] = a[9] & g[976];
assign g[1999] = b[9] & g[976];
assign g[1489] = a[9] & g[977];
assign g[2000] = b[9] & g[977];
assign g[1490] = a[9] & g[978];
assign g[2001] = b[9] & g[978];
assign g[1491] = a[9] & g[979];
assign g[2002] = b[9] & g[979];
assign g[1492] = a[9] & g[980];
assign g[2003] = b[9] & g[980];
assign g[1493] = a[9] & g[981];
assign g[2004] = b[9] & g[981];
assign g[1494] = a[9] & g[982];
assign g[2005] = b[9] & g[982];
assign g[1495] = a[9] & g[983];
assign g[2006] = b[9] & g[983];
assign g[1496] = a[9] & g[984];
assign g[2007] = b[9] & g[984];
assign g[1497] = a[9] & g[985];
assign g[2008] = b[9] & g[985];
assign g[1498] = a[9] & g[986];
assign g[2009] = b[9] & g[986];
assign g[1499] = a[9] & g[987];
assign g[2010] = b[9] & g[987];
assign g[1500] = a[9] & g[988];
assign g[2011] = b[9] & g[988];
assign g[1501] = a[9] & g[989];
assign g[2012] = b[9] & g[989];
assign g[1502] = a[9] & g[990];
assign g[2013] = b[9] & g[990];
assign g[1503] = a[9] & g[991];
assign g[2014] = b[9] & g[991];
assign g[1504] = a[9] & g[992];
assign g[2015] = b[9] & g[992];
assign g[1505] = a[9] & g[993];
assign g[2016] = b[9] & g[993];
assign g[1506] = a[9] & g[994];
assign g[2017] = b[9] & g[994];
assign g[1507] = a[9] & g[995];
assign g[2018] = b[9] & g[995];
assign g[1508] = a[9] & g[996];
assign g[2019] = b[9] & g[996];
assign g[1509] = a[9] & g[997];
assign g[2020] = b[9] & g[997];
assign g[1510] = a[9] & g[998];
assign g[2021] = b[9] & g[998];
assign g[1511] = a[9] & g[999];
assign g[2022] = b[9] & g[999];
assign g[1512] = a[9] & g[1000];
assign g[2023] = b[9] & g[1000];
assign g[1513] = a[9] & g[1001];
assign g[2024] = b[9] & g[1001];
assign g[1514] = a[9] & g[1002];
assign g[2025] = b[9] & g[1002];
assign g[1515] = a[9] & g[1003];
assign g[2026] = b[9] & g[1003];
assign g[1516] = a[9] & g[1004];
assign g[2027] = b[9] & g[1004];
assign g[1517] = a[9] & g[1005];
assign g[2028] = b[9] & g[1005];
assign g[1518] = a[9] & g[1006];
assign g[2029] = b[9] & g[1006];
assign g[1519] = a[9] & g[1007];
assign g[2030] = b[9] & g[1007];
assign g[1520] = a[9] & g[1008];
assign g[2031] = b[9] & g[1008];
assign g[1521] = a[9] & g[1009];
assign g[2032] = b[9] & g[1009];
assign g[1522] = a[9] & g[1010];
assign g[2033] = b[9] & g[1010];
assign g[1523] = a[9] & g[1011];
assign g[2034] = b[9] & g[1011];
assign g[1524] = a[9] & g[1012];
assign g[2035] = b[9] & g[1012];
//Assigning outputs for input bit 11
assign g[2036] = a[10] & b[10];
assign g[2037] = a[10] & g[1013];
assign g[3060] = b[10] & g[1013];
assign g[2038] = a[10] & g[1014];
assign g[3061] = b[10] & g[1014];
assign g[2039] = a[10] & g[1015];
assign g[3062] = b[10] & g[1015];
assign g[2040] = a[10] & g[1016];
assign g[3063] = b[10] & g[1016];
assign g[2041] = a[10] & g[1017];
assign g[3064] = b[10] & g[1017];
assign g[2042] = a[10] & g[1018];
assign g[3065] = b[10] & g[1018];
assign g[2043] = a[10] & g[1019];
assign g[3066] = b[10] & g[1019];
assign g[2044] = a[10] & g[1020];
assign g[3067] = b[10] & g[1020];
assign g[2045] = a[10] & g[1021];
assign g[3068] = b[10] & g[1021];
assign g[2046] = a[10] & g[1022];
assign g[3069] = b[10] & g[1022];
assign g[2047] = a[10] & g[1023];
assign g[3070] = b[10] & g[1023];
assign g[2048] = a[10] & g[1024];
assign g[3071] = b[10] & g[1024];
assign g[2049] = a[10] & g[1025];
assign g[3072] = b[10] & g[1025];
assign g[2050] = a[10] & g[1026];
assign g[3073] = b[10] & g[1026];
assign g[2051] = a[10] & g[1027];
assign g[3074] = b[10] & g[1027];
assign g[2052] = a[10] & g[1028];
assign g[3075] = b[10] & g[1028];
assign g[2053] = a[10] & g[1029];
assign g[3076] = b[10] & g[1029];
assign g[2054] = a[10] & g[1030];
assign g[3077] = b[10] & g[1030];
assign g[2055] = a[10] & g[1031];
assign g[3078] = b[10] & g[1031];
assign g[2056] = a[10] & g[1032];
assign g[3079] = b[10] & g[1032];
assign g[2057] = a[10] & g[1033];
assign g[3080] = b[10] & g[1033];
assign g[2058] = a[10] & g[1034];
assign g[3081] = b[10] & g[1034];
assign g[2059] = a[10] & g[1035];
assign g[3082] = b[10] & g[1035];
assign g[2060] = a[10] & g[1036];
assign g[3083] = b[10] & g[1036];
assign g[2061] = a[10] & g[1037];
assign g[3084] = b[10] & g[1037];
assign g[2062] = a[10] & g[1038];
assign g[3085] = b[10] & g[1038];
assign g[2063] = a[10] & g[1039];
assign g[3086] = b[10] & g[1039];
assign g[2064] = a[10] & g[1040];
assign g[3087] = b[10] & g[1040];
assign g[2065] = a[10] & g[1041];
assign g[3088] = b[10] & g[1041];
assign g[2066] = a[10] & g[1042];
assign g[3089] = b[10] & g[1042];
assign g[2067] = a[10] & g[1043];
assign g[3090] = b[10] & g[1043];
assign g[2068] = a[10] & g[1044];
assign g[3091] = b[10] & g[1044];
assign g[2069] = a[10] & g[1045];
assign g[3092] = b[10] & g[1045];
assign g[2070] = a[10] & g[1046];
assign g[3093] = b[10] & g[1046];
assign g[2071] = a[10] & g[1047];
assign g[3094] = b[10] & g[1047];
assign g[2072] = a[10] & g[1048];
assign g[3095] = b[10] & g[1048];
assign g[2073] = a[10] & g[1049];
assign g[3096] = b[10] & g[1049];
assign g[2074] = a[10] & g[1050];
assign g[3097] = b[10] & g[1050];
assign g[2075] = a[10] & g[1051];
assign g[3098] = b[10] & g[1051];
assign g[2076] = a[10] & g[1052];
assign g[3099] = b[10] & g[1052];
assign g[2077] = a[10] & g[1053];
assign g[3100] = b[10] & g[1053];
assign g[2078] = a[10] & g[1054];
assign g[3101] = b[10] & g[1054];
assign g[2079] = a[10] & g[1055];
assign g[3102] = b[10] & g[1055];
assign g[2080] = a[10] & g[1056];
assign g[3103] = b[10] & g[1056];
assign g[2081] = a[10] & g[1057];
assign g[3104] = b[10] & g[1057];
assign g[2082] = a[10] & g[1058];
assign g[3105] = b[10] & g[1058];
assign g[2083] = a[10] & g[1059];
assign g[3106] = b[10] & g[1059];
assign g[2084] = a[10] & g[1060];
assign g[3107] = b[10] & g[1060];
assign g[2085] = a[10] & g[1061];
assign g[3108] = b[10] & g[1061];
assign g[2086] = a[10] & g[1062];
assign g[3109] = b[10] & g[1062];
assign g[2087] = a[10] & g[1063];
assign g[3110] = b[10] & g[1063];
assign g[2088] = a[10] & g[1064];
assign g[3111] = b[10] & g[1064];
assign g[2089] = a[10] & g[1065];
assign g[3112] = b[10] & g[1065];
assign g[2090] = a[10] & g[1066];
assign g[3113] = b[10] & g[1066];
assign g[2091] = a[10] & g[1067];
assign g[3114] = b[10] & g[1067];
assign g[2092] = a[10] & g[1068];
assign g[3115] = b[10] & g[1068];
assign g[2093] = a[10] & g[1069];
assign g[3116] = b[10] & g[1069];
assign g[2094] = a[10] & g[1070];
assign g[3117] = b[10] & g[1070];
assign g[2095] = a[10] & g[1071];
assign g[3118] = b[10] & g[1071];
assign g[2096] = a[10] & g[1072];
assign g[3119] = b[10] & g[1072];
assign g[2097] = a[10] & g[1073];
assign g[3120] = b[10] & g[1073];
assign g[2098] = a[10] & g[1074];
assign g[3121] = b[10] & g[1074];
assign g[2099] = a[10] & g[1075];
assign g[3122] = b[10] & g[1075];
assign g[2100] = a[10] & g[1076];
assign g[3123] = b[10] & g[1076];
assign g[2101] = a[10] & g[1077];
assign g[3124] = b[10] & g[1077];
assign g[2102] = a[10] & g[1078];
assign g[3125] = b[10] & g[1078];
assign g[2103] = a[10] & g[1079];
assign g[3126] = b[10] & g[1079];
assign g[2104] = a[10] & g[1080];
assign g[3127] = b[10] & g[1080];
assign g[2105] = a[10] & g[1081];
assign g[3128] = b[10] & g[1081];
assign g[2106] = a[10] & g[1082];
assign g[3129] = b[10] & g[1082];
assign g[2107] = a[10] & g[1083];
assign g[3130] = b[10] & g[1083];
assign g[2108] = a[10] & g[1084];
assign g[3131] = b[10] & g[1084];
assign g[2109] = a[10] & g[1085];
assign g[3132] = b[10] & g[1085];
assign g[2110] = a[10] & g[1086];
assign g[3133] = b[10] & g[1086];
assign g[2111] = a[10] & g[1087];
assign g[3134] = b[10] & g[1087];
assign g[2112] = a[10] & g[1088];
assign g[3135] = b[10] & g[1088];
assign g[2113] = a[10] & g[1089];
assign g[3136] = b[10] & g[1089];
assign g[2114] = a[10] & g[1090];
assign g[3137] = b[10] & g[1090];
assign g[2115] = a[10] & g[1091];
assign g[3138] = b[10] & g[1091];
assign g[2116] = a[10] & g[1092];
assign g[3139] = b[10] & g[1092];
assign g[2117] = a[10] & g[1093];
assign g[3140] = b[10] & g[1093];
assign g[2118] = a[10] & g[1094];
assign g[3141] = b[10] & g[1094];
assign g[2119] = a[10] & g[1095];
assign g[3142] = b[10] & g[1095];
assign g[2120] = a[10] & g[1096];
assign g[3143] = b[10] & g[1096];
assign g[2121] = a[10] & g[1097];
assign g[3144] = b[10] & g[1097];
assign g[2122] = a[10] & g[1098];
assign g[3145] = b[10] & g[1098];
assign g[2123] = a[10] & g[1099];
assign g[3146] = b[10] & g[1099];
assign g[2124] = a[10] & g[1100];
assign g[3147] = b[10] & g[1100];
assign g[2125] = a[10] & g[1101];
assign g[3148] = b[10] & g[1101];
assign g[2126] = a[10] & g[1102];
assign g[3149] = b[10] & g[1102];
assign g[2127] = a[10] & g[1103];
assign g[3150] = b[10] & g[1103];
assign g[2128] = a[10] & g[1104];
assign g[3151] = b[10] & g[1104];
assign g[2129] = a[10] & g[1105];
assign g[3152] = b[10] & g[1105];
assign g[2130] = a[10] & g[1106];
assign g[3153] = b[10] & g[1106];
assign g[2131] = a[10] & g[1107];
assign g[3154] = b[10] & g[1107];
assign g[2132] = a[10] & g[1108];
assign g[3155] = b[10] & g[1108];
assign g[2133] = a[10] & g[1109];
assign g[3156] = b[10] & g[1109];
assign g[2134] = a[10] & g[1110];
assign g[3157] = b[10] & g[1110];
assign g[2135] = a[10] & g[1111];
assign g[3158] = b[10] & g[1111];
assign g[2136] = a[10] & g[1112];
assign g[3159] = b[10] & g[1112];
assign g[2137] = a[10] & g[1113];
assign g[3160] = b[10] & g[1113];
assign g[2138] = a[10] & g[1114];
assign g[3161] = b[10] & g[1114];
assign g[2139] = a[10] & g[1115];
assign g[3162] = b[10] & g[1115];
assign g[2140] = a[10] & g[1116];
assign g[3163] = b[10] & g[1116];
assign g[2141] = a[10] & g[1117];
assign g[3164] = b[10] & g[1117];
assign g[2142] = a[10] & g[1118];
assign g[3165] = b[10] & g[1118];
assign g[2143] = a[10] & g[1119];
assign g[3166] = b[10] & g[1119];
assign g[2144] = a[10] & g[1120];
assign g[3167] = b[10] & g[1120];
assign g[2145] = a[10] & g[1121];
assign g[3168] = b[10] & g[1121];
assign g[2146] = a[10] & g[1122];
assign g[3169] = b[10] & g[1122];
assign g[2147] = a[10] & g[1123];
assign g[3170] = b[10] & g[1123];
assign g[2148] = a[10] & g[1124];
assign g[3171] = b[10] & g[1124];
assign g[2149] = a[10] & g[1125];
assign g[3172] = b[10] & g[1125];
assign g[2150] = a[10] & g[1126];
assign g[3173] = b[10] & g[1126];
assign g[2151] = a[10] & g[1127];
assign g[3174] = b[10] & g[1127];
assign g[2152] = a[10] & g[1128];
assign g[3175] = b[10] & g[1128];
assign g[2153] = a[10] & g[1129];
assign g[3176] = b[10] & g[1129];
assign g[2154] = a[10] & g[1130];
assign g[3177] = b[10] & g[1130];
assign g[2155] = a[10] & g[1131];
assign g[3178] = b[10] & g[1131];
assign g[2156] = a[10] & g[1132];
assign g[3179] = b[10] & g[1132];
assign g[2157] = a[10] & g[1133];
assign g[3180] = b[10] & g[1133];
assign g[2158] = a[10] & g[1134];
assign g[3181] = b[10] & g[1134];
assign g[2159] = a[10] & g[1135];
assign g[3182] = b[10] & g[1135];
assign g[2160] = a[10] & g[1136];
assign g[3183] = b[10] & g[1136];
assign g[2161] = a[10] & g[1137];
assign g[3184] = b[10] & g[1137];
assign g[2162] = a[10] & g[1138];
assign g[3185] = b[10] & g[1138];
assign g[2163] = a[10] & g[1139];
assign g[3186] = b[10] & g[1139];
assign g[2164] = a[10] & g[1140];
assign g[3187] = b[10] & g[1140];
assign g[2165] = a[10] & g[1141];
assign g[3188] = b[10] & g[1141];
assign g[2166] = a[10] & g[1142];
assign g[3189] = b[10] & g[1142];
assign g[2167] = a[10] & g[1143];
assign g[3190] = b[10] & g[1143];
assign g[2168] = a[10] & g[1144];
assign g[3191] = b[10] & g[1144];
assign g[2169] = a[10] & g[1145];
assign g[3192] = b[10] & g[1145];
assign g[2170] = a[10] & g[1146];
assign g[3193] = b[10] & g[1146];
assign g[2171] = a[10] & g[1147];
assign g[3194] = b[10] & g[1147];
assign g[2172] = a[10] & g[1148];
assign g[3195] = b[10] & g[1148];
assign g[2173] = a[10] & g[1149];
assign g[3196] = b[10] & g[1149];
assign g[2174] = a[10] & g[1150];
assign g[3197] = b[10] & g[1150];
assign g[2175] = a[10] & g[1151];
assign g[3198] = b[10] & g[1151];
assign g[2176] = a[10] & g[1152];
assign g[3199] = b[10] & g[1152];
assign g[2177] = a[10] & g[1153];
assign g[3200] = b[10] & g[1153];
assign g[2178] = a[10] & g[1154];
assign g[3201] = b[10] & g[1154];
assign g[2179] = a[10] & g[1155];
assign g[3202] = b[10] & g[1155];
assign g[2180] = a[10] & g[1156];
assign g[3203] = b[10] & g[1156];
assign g[2181] = a[10] & g[1157];
assign g[3204] = b[10] & g[1157];
assign g[2182] = a[10] & g[1158];
assign g[3205] = b[10] & g[1158];
assign g[2183] = a[10] & g[1159];
assign g[3206] = b[10] & g[1159];
assign g[2184] = a[10] & g[1160];
assign g[3207] = b[10] & g[1160];
assign g[2185] = a[10] & g[1161];
assign g[3208] = b[10] & g[1161];
assign g[2186] = a[10] & g[1162];
assign g[3209] = b[10] & g[1162];
assign g[2187] = a[10] & g[1163];
assign g[3210] = b[10] & g[1163];
assign g[2188] = a[10] & g[1164];
assign g[3211] = b[10] & g[1164];
assign g[2189] = a[10] & g[1165];
assign g[3212] = b[10] & g[1165];
assign g[2190] = a[10] & g[1166];
assign g[3213] = b[10] & g[1166];
assign g[2191] = a[10] & g[1167];
assign g[3214] = b[10] & g[1167];
assign g[2192] = a[10] & g[1168];
assign g[3215] = b[10] & g[1168];
assign g[2193] = a[10] & g[1169];
assign g[3216] = b[10] & g[1169];
assign g[2194] = a[10] & g[1170];
assign g[3217] = b[10] & g[1170];
assign g[2195] = a[10] & g[1171];
assign g[3218] = b[10] & g[1171];
assign g[2196] = a[10] & g[1172];
assign g[3219] = b[10] & g[1172];
assign g[2197] = a[10] & g[1173];
assign g[3220] = b[10] & g[1173];
assign g[2198] = a[10] & g[1174];
assign g[3221] = b[10] & g[1174];
assign g[2199] = a[10] & g[1175];
assign g[3222] = b[10] & g[1175];
assign g[2200] = a[10] & g[1176];
assign g[3223] = b[10] & g[1176];
assign g[2201] = a[10] & g[1177];
assign g[3224] = b[10] & g[1177];
assign g[2202] = a[10] & g[1178];
assign g[3225] = b[10] & g[1178];
assign g[2203] = a[10] & g[1179];
assign g[3226] = b[10] & g[1179];
assign g[2204] = a[10] & g[1180];
assign g[3227] = b[10] & g[1180];
assign g[2205] = a[10] & g[1181];
assign g[3228] = b[10] & g[1181];
assign g[2206] = a[10] & g[1182];
assign g[3229] = b[10] & g[1182];
assign g[2207] = a[10] & g[1183];
assign g[3230] = b[10] & g[1183];
assign g[2208] = a[10] & g[1184];
assign g[3231] = b[10] & g[1184];
assign g[2209] = a[10] & g[1185];
assign g[3232] = b[10] & g[1185];
assign g[2210] = a[10] & g[1186];
assign g[3233] = b[10] & g[1186];
assign g[2211] = a[10] & g[1187];
assign g[3234] = b[10] & g[1187];
assign g[2212] = a[10] & g[1188];
assign g[3235] = b[10] & g[1188];
assign g[2213] = a[10] & g[1189];
assign g[3236] = b[10] & g[1189];
assign g[2214] = a[10] & g[1190];
assign g[3237] = b[10] & g[1190];
assign g[2215] = a[10] & g[1191];
assign g[3238] = b[10] & g[1191];
assign g[2216] = a[10] & g[1192];
assign g[3239] = b[10] & g[1192];
assign g[2217] = a[10] & g[1193];
assign g[3240] = b[10] & g[1193];
assign g[2218] = a[10] & g[1194];
assign g[3241] = b[10] & g[1194];
assign g[2219] = a[10] & g[1195];
assign g[3242] = b[10] & g[1195];
assign g[2220] = a[10] & g[1196];
assign g[3243] = b[10] & g[1196];
assign g[2221] = a[10] & g[1197];
assign g[3244] = b[10] & g[1197];
assign g[2222] = a[10] & g[1198];
assign g[3245] = b[10] & g[1198];
assign g[2223] = a[10] & g[1199];
assign g[3246] = b[10] & g[1199];
assign g[2224] = a[10] & g[1200];
assign g[3247] = b[10] & g[1200];
assign g[2225] = a[10] & g[1201];
assign g[3248] = b[10] & g[1201];
assign g[2226] = a[10] & g[1202];
assign g[3249] = b[10] & g[1202];
assign g[2227] = a[10] & g[1203];
assign g[3250] = b[10] & g[1203];
assign g[2228] = a[10] & g[1204];
assign g[3251] = b[10] & g[1204];
assign g[2229] = a[10] & g[1205];
assign g[3252] = b[10] & g[1205];
assign g[2230] = a[10] & g[1206];
assign g[3253] = b[10] & g[1206];
assign g[2231] = a[10] & g[1207];
assign g[3254] = b[10] & g[1207];
assign g[2232] = a[10] & g[1208];
assign g[3255] = b[10] & g[1208];
assign g[2233] = a[10] & g[1209];
assign g[3256] = b[10] & g[1209];
assign g[2234] = a[10] & g[1210];
assign g[3257] = b[10] & g[1210];
assign g[2235] = a[10] & g[1211];
assign g[3258] = b[10] & g[1211];
assign g[2236] = a[10] & g[1212];
assign g[3259] = b[10] & g[1212];
assign g[2237] = a[10] & g[1213];
assign g[3260] = b[10] & g[1213];
assign g[2238] = a[10] & g[1214];
assign g[3261] = b[10] & g[1214];
assign g[2239] = a[10] & g[1215];
assign g[3262] = b[10] & g[1215];
assign g[2240] = a[10] & g[1216];
assign g[3263] = b[10] & g[1216];
assign g[2241] = a[10] & g[1217];
assign g[3264] = b[10] & g[1217];
assign g[2242] = a[10] & g[1218];
assign g[3265] = b[10] & g[1218];
assign g[2243] = a[10] & g[1219];
assign g[3266] = b[10] & g[1219];
assign g[2244] = a[10] & g[1220];
assign g[3267] = b[10] & g[1220];
assign g[2245] = a[10] & g[1221];
assign g[3268] = b[10] & g[1221];
assign g[2246] = a[10] & g[1222];
assign g[3269] = b[10] & g[1222];
assign g[2247] = a[10] & g[1223];
assign g[3270] = b[10] & g[1223];
assign g[2248] = a[10] & g[1224];
assign g[3271] = b[10] & g[1224];
assign g[2249] = a[10] & g[1225];
assign g[3272] = b[10] & g[1225];
assign g[2250] = a[10] & g[1226];
assign g[3273] = b[10] & g[1226];
assign g[2251] = a[10] & g[1227];
assign g[3274] = b[10] & g[1227];
assign g[2252] = a[10] & g[1228];
assign g[3275] = b[10] & g[1228];
assign g[2253] = a[10] & g[1229];
assign g[3276] = b[10] & g[1229];
assign g[2254] = a[10] & g[1230];
assign g[3277] = b[10] & g[1230];
assign g[2255] = a[10] & g[1231];
assign g[3278] = b[10] & g[1231];
assign g[2256] = a[10] & g[1232];
assign g[3279] = b[10] & g[1232];
assign g[2257] = a[10] & g[1233];
assign g[3280] = b[10] & g[1233];
assign g[2258] = a[10] & g[1234];
assign g[3281] = b[10] & g[1234];
assign g[2259] = a[10] & g[1235];
assign g[3282] = b[10] & g[1235];
assign g[2260] = a[10] & g[1236];
assign g[3283] = b[10] & g[1236];
assign g[2261] = a[10] & g[1237];
assign g[3284] = b[10] & g[1237];
assign g[2262] = a[10] & g[1238];
assign g[3285] = b[10] & g[1238];
assign g[2263] = a[10] & g[1239];
assign g[3286] = b[10] & g[1239];
assign g[2264] = a[10] & g[1240];
assign g[3287] = b[10] & g[1240];
assign g[2265] = a[10] & g[1241];
assign g[3288] = b[10] & g[1241];
assign g[2266] = a[10] & g[1242];
assign g[3289] = b[10] & g[1242];
assign g[2267] = a[10] & g[1243];
assign g[3290] = b[10] & g[1243];
assign g[2268] = a[10] & g[1244];
assign g[3291] = b[10] & g[1244];
assign g[2269] = a[10] & g[1245];
assign g[3292] = b[10] & g[1245];
assign g[2270] = a[10] & g[1246];
assign g[3293] = b[10] & g[1246];
assign g[2271] = a[10] & g[1247];
assign g[3294] = b[10] & g[1247];
assign g[2272] = a[10] & g[1248];
assign g[3295] = b[10] & g[1248];
assign g[2273] = a[10] & g[1249];
assign g[3296] = b[10] & g[1249];
assign g[2274] = a[10] & g[1250];
assign g[3297] = b[10] & g[1250];
assign g[2275] = a[10] & g[1251];
assign g[3298] = b[10] & g[1251];
assign g[2276] = a[10] & g[1252];
assign g[3299] = b[10] & g[1252];
assign g[2277] = a[10] & g[1253];
assign g[3300] = b[10] & g[1253];
assign g[2278] = a[10] & g[1254];
assign g[3301] = b[10] & g[1254];
assign g[2279] = a[10] & g[1255];
assign g[3302] = b[10] & g[1255];
assign g[2280] = a[10] & g[1256];
assign g[3303] = b[10] & g[1256];
assign g[2281] = a[10] & g[1257];
assign g[3304] = b[10] & g[1257];
assign g[2282] = a[10] & g[1258];
assign g[3305] = b[10] & g[1258];
assign g[2283] = a[10] & g[1259];
assign g[3306] = b[10] & g[1259];
assign g[2284] = a[10] & g[1260];
assign g[3307] = b[10] & g[1260];
assign g[2285] = a[10] & g[1261];
assign g[3308] = b[10] & g[1261];
assign g[2286] = a[10] & g[1262];
assign g[3309] = b[10] & g[1262];
assign g[2287] = a[10] & g[1263];
assign g[3310] = b[10] & g[1263];
assign g[2288] = a[10] & g[1264];
assign g[3311] = b[10] & g[1264];
assign g[2289] = a[10] & g[1265];
assign g[3312] = b[10] & g[1265];
assign g[2290] = a[10] & g[1266];
assign g[3313] = b[10] & g[1266];
assign g[2291] = a[10] & g[1267];
assign g[3314] = b[10] & g[1267];
assign g[2292] = a[10] & g[1268];
assign g[3315] = b[10] & g[1268];
assign g[2293] = a[10] & g[1269];
assign g[3316] = b[10] & g[1269];
assign g[2294] = a[10] & g[1270];
assign g[3317] = b[10] & g[1270];
assign g[2295] = a[10] & g[1271];
assign g[3318] = b[10] & g[1271];
assign g[2296] = a[10] & g[1272];
assign g[3319] = b[10] & g[1272];
assign g[2297] = a[10] & g[1273];
assign g[3320] = b[10] & g[1273];
assign g[2298] = a[10] & g[1274];
assign g[3321] = b[10] & g[1274];
assign g[2299] = a[10] & g[1275];
assign g[3322] = b[10] & g[1275];
assign g[2300] = a[10] & g[1276];
assign g[3323] = b[10] & g[1276];
assign g[2301] = a[10] & g[1277];
assign g[3324] = b[10] & g[1277];
assign g[2302] = a[10] & g[1278];
assign g[3325] = b[10] & g[1278];
assign g[2303] = a[10] & g[1279];
assign g[3326] = b[10] & g[1279];
assign g[2304] = a[10] & g[1280];
assign g[3327] = b[10] & g[1280];
assign g[2305] = a[10] & g[1281];
assign g[3328] = b[10] & g[1281];
assign g[2306] = a[10] & g[1282];
assign g[3329] = b[10] & g[1282];
assign g[2307] = a[10] & g[1283];
assign g[3330] = b[10] & g[1283];
assign g[2308] = a[10] & g[1284];
assign g[3331] = b[10] & g[1284];
assign g[2309] = a[10] & g[1285];
assign g[3332] = b[10] & g[1285];
assign g[2310] = a[10] & g[1286];
assign g[3333] = b[10] & g[1286];
assign g[2311] = a[10] & g[1287];
assign g[3334] = b[10] & g[1287];
assign g[2312] = a[10] & g[1288];
assign g[3335] = b[10] & g[1288];
assign g[2313] = a[10] & g[1289];
assign g[3336] = b[10] & g[1289];
assign g[2314] = a[10] & g[1290];
assign g[3337] = b[10] & g[1290];
assign g[2315] = a[10] & g[1291];
assign g[3338] = b[10] & g[1291];
assign g[2316] = a[10] & g[1292];
assign g[3339] = b[10] & g[1292];
assign g[2317] = a[10] & g[1293];
assign g[3340] = b[10] & g[1293];
assign g[2318] = a[10] & g[1294];
assign g[3341] = b[10] & g[1294];
assign g[2319] = a[10] & g[1295];
assign g[3342] = b[10] & g[1295];
assign g[2320] = a[10] & g[1296];
assign g[3343] = b[10] & g[1296];
assign g[2321] = a[10] & g[1297];
assign g[3344] = b[10] & g[1297];
assign g[2322] = a[10] & g[1298];
assign g[3345] = b[10] & g[1298];
assign g[2323] = a[10] & g[1299];
assign g[3346] = b[10] & g[1299];
assign g[2324] = a[10] & g[1300];
assign g[3347] = b[10] & g[1300];
assign g[2325] = a[10] & g[1301];
assign g[3348] = b[10] & g[1301];
assign g[2326] = a[10] & g[1302];
assign g[3349] = b[10] & g[1302];
assign g[2327] = a[10] & g[1303];
assign g[3350] = b[10] & g[1303];
assign g[2328] = a[10] & g[1304];
assign g[3351] = b[10] & g[1304];
assign g[2329] = a[10] & g[1305];
assign g[3352] = b[10] & g[1305];
assign g[2330] = a[10] & g[1306];
assign g[3353] = b[10] & g[1306];
assign g[2331] = a[10] & g[1307];
assign g[3354] = b[10] & g[1307];
assign g[2332] = a[10] & g[1308];
assign g[3355] = b[10] & g[1308];
assign g[2333] = a[10] & g[1309];
assign g[3356] = b[10] & g[1309];
assign g[2334] = a[10] & g[1310];
assign g[3357] = b[10] & g[1310];
assign g[2335] = a[10] & g[1311];
assign g[3358] = b[10] & g[1311];
assign g[2336] = a[10] & g[1312];
assign g[3359] = b[10] & g[1312];
assign g[2337] = a[10] & g[1313];
assign g[3360] = b[10] & g[1313];
assign g[2338] = a[10] & g[1314];
assign g[3361] = b[10] & g[1314];
assign g[2339] = a[10] & g[1315];
assign g[3362] = b[10] & g[1315];
assign g[2340] = a[10] & g[1316];
assign g[3363] = b[10] & g[1316];
assign g[2341] = a[10] & g[1317];
assign g[3364] = b[10] & g[1317];
assign g[2342] = a[10] & g[1318];
assign g[3365] = b[10] & g[1318];
assign g[2343] = a[10] & g[1319];
assign g[3366] = b[10] & g[1319];
assign g[2344] = a[10] & g[1320];
assign g[3367] = b[10] & g[1320];
assign g[2345] = a[10] & g[1321];
assign g[3368] = b[10] & g[1321];
assign g[2346] = a[10] & g[1322];
assign g[3369] = b[10] & g[1322];
assign g[2347] = a[10] & g[1323];
assign g[3370] = b[10] & g[1323];
assign g[2348] = a[10] & g[1324];
assign g[3371] = b[10] & g[1324];
assign g[2349] = a[10] & g[1325];
assign g[3372] = b[10] & g[1325];
assign g[2350] = a[10] & g[1326];
assign g[3373] = b[10] & g[1326];
assign g[2351] = a[10] & g[1327];
assign g[3374] = b[10] & g[1327];
assign g[2352] = a[10] & g[1328];
assign g[3375] = b[10] & g[1328];
assign g[2353] = a[10] & g[1329];
assign g[3376] = b[10] & g[1329];
assign g[2354] = a[10] & g[1330];
assign g[3377] = b[10] & g[1330];
assign g[2355] = a[10] & g[1331];
assign g[3378] = b[10] & g[1331];
assign g[2356] = a[10] & g[1332];
assign g[3379] = b[10] & g[1332];
assign g[2357] = a[10] & g[1333];
assign g[3380] = b[10] & g[1333];
assign g[2358] = a[10] & g[1334];
assign g[3381] = b[10] & g[1334];
assign g[2359] = a[10] & g[1335];
assign g[3382] = b[10] & g[1335];
assign g[2360] = a[10] & g[1336];
assign g[3383] = b[10] & g[1336];
assign g[2361] = a[10] & g[1337];
assign g[3384] = b[10] & g[1337];
assign g[2362] = a[10] & g[1338];
assign g[3385] = b[10] & g[1338];
assign g[2363] = a[10] & g[1339];
assign g[3386] = b[10] & g[1339];
assign g[2364] = a[10] & g[1340];
assign g[3387] = b[10] & g[1340];
assign g[2365] = a[10] & g[1341];
assign g[3388] = b[10] & g[1341];
assign g[2366] = a[10] & g[1342];
assign g[3389] = b[10] & g[1342];
assign g[2367] = a[10] & g[1343];
assign g[3390] = b[10] & g[1343];
assign g[2368] = a[10] & g[1344];
assign g[3391] = b[10] & g[1344];
assign g[2369] = a[10] & g[1345];
assign g[3392] = b[10] & g[1345];
assign g[2370] = a[10] & g[1346];
assign g[3393] = b[10] & g[1346];
assign g[2371] = a[10] & g[1347];
assign g[3394] = b[10] & g[1347];
assign g[2372] = a[10] & g[1348];
assign g[3395] = b[10] & g[1348];
assign g[2373] = a[10] & g[1349];
assign g[3396] = b[10] & g[1349];
assign g[2374] = a[10] & g[1350];
assign g[3397] = b[10] & g[1350];
assign g[2375] = a[10] & g[1351];
assign g[3398] = b[10] & g[1351];
assign g[2376] = a[10] & g[1352];
assign g[3399] = b[10] & g[1352];
assign g[2377] = a[10] & g[1353];
assign g[3400] = b[10] & g[1353];
assign g[2378] = a[10] & g[1354];
assign g[3401] = b[10] & g[1354];
assign g[2379] = a[10] & g[1355];
assign g[3402] = b[10] & g[1355];
assign g[2380] = a[10] & g[1356];
assign g[3403] = b[10] & g[1356];
assign g[2381] = a[10] & g[1357];
assign g[3404] = b[10] & g[1357];
assign g[2382] = a[10] & g[1358];
assign g[3405] = b[10] & g[1358];
assign g[2383] = a[10] & g[1359];
assign g[3406] = b[10] & g[1359];
assign g[2384] = a[10] & g[1360];
assign g[3407] = b[10] & g[1360];
assign g[2385] = a[10] & g[1361];
assign g[3408] = b[10] & g[1361];
assign g[2386] = a[10] & g[1362];
assign g[3409] = b[10] & g[1362];
assign g[2387] = a[10] & g[1363];
assign g[3410] = b[10] & g[1363];
assign g[2388] = a[10] & g[1364];
assign g[3411] = b[10] & g[1364];
assign g[2389] = a[10] & g[1365];
assign g[3412] = b[10] & g[1365];
assign g[2390] = a[10] & g[1366];
assign g[3413] = b[10] & g[1366];
assign g[2391] = a[10] & g[1367];
assign g[3414] = b[10] & g[1367];
assign g[2392] = a[10] & g[1368];
assign g[3415] = b[10] & g[1368];
assign g[2393] = a[10] & g[1369];
assign g[3416] = b[10] & g[1369];
assign g[2394] = a[10] & g[1370];
assign g[3417] = b[10] & g[1370];
assign g[2395] = a[10] & g[1371];
assign g[3418] = b[10] & g[1371];
assign g[2396] = a[10] & g[1372];
assign g[3419] = b[10] & g[1372];
assign g[2397] = a[10] & g[1373];
assign g[3420] = b[10] & g[1373];
assign g[2398] = a[10] & g[1374];
assign g[3421] = b[10] & g[1374];
assign g[2399] = a[10] & g[1375];
assign g[3422] = b[10] & g[1375];
assign g[2400] = a[10] & g[1376];
assign g[3423] = b[10] & g[1376];
assign g[2401] = a[10] & g[1377];
assign g[3424] = b[10] & g[1377];
assign g[2402] = a[10] & g[1378];
assign g[3425] = b[10] & g[1378];
assign g[2403] = a[10] & g[1379];
assign g[3426] = b[10] & g[1379];
assign g[2404] = a[10] & g[1380];
assign g[3427] = b[10] & g[1380];
assign g[2405] = a[10] & g[1381];
assign g[3428] = b[10] & g[1381];
assign g[2406] = a[10] & g[1382];
assign g[3429] = b[10] & g[1382];
assign g[2407] = a[10] & g[1383];
assign g[3430] = b[10] & g[1383];
assign g[2408] = a[10] & g[1384];
assign g[3431] = b[10] & g[1384];
assign g[2409] = a[10] & g[1385];
assign g[3432] = b[10] & g[1385];
assign g[2410] = a[10] & g[1386];
assign g[3433] = b[10] & g[1386];
assign g[2411] = a[10] & g[1387];
assign g[3434] = b[10] & g[1387];
assign g[2412] = a[10] & g[1388];
assign g[3435] = b[10] & g[1388];
assign g[2413] = a[10] & g[1389];
assign g[3436] = b[10] & g[1389];
assign g[2414] = a[10] & g[1390];
assign g[3437] = b[10] & g[1390];
assign g[2415] = a[10] & g[1391];
assign g[3438] = b[10] & g[1391];
assign g[2416] = a[10] & g[1392];
assign g[3439] = b[10] & g[1392];
assign g[2417] = a[10] & g[1393];
assign g[3440] = b[10] & g[1393];
assign g[2418] = a[10] & g[1394];
assign g[3441] = b[10] & g[1394];
assign g[2419] = a[10] & g[1395];
assign g[3442] = b[10] & g[1395];
assign g[2420] = a[10] & g[1396];
assign g[3443] = b[10] & g[1396];
assign g[2421] = a[10] & g[1397];
assign g[3444] = b[10] & g[1397];
assign g[2422] = a[10] & g[1398];
assign g[3445] = b[10] & g[1398];
assign g[2423] = a[10] & g[1399];
assign g[3446] = b[10] & g[1399];
assign g[2424] = a[10] & g[1400];
assign g[3447] = b[10] & g[1400];
assign g[2425] = a[10] & g[1401];
assign g[3448] = b[10] & g[1401];
assign g[2426] = a[10] & g[1402];
assign g[3449] = b[10] & g[1402];
assign g[2427] = a[10] & g[1403];
assign g[3450] = b[10] & g[1403];
assign g[2428] = a[10] & g[1404];
assign g[3451] = b[10] & g[1404];
assign g[2429] = a[10] & g[1405];
assign g[3452] = b[10] & g[1405];
assign g[2430] = a[10] & g[1406];
assign g[3453] = b[10] & g[1406];
assign g[2431] = a[10] & g[1407];
assign g[3454] = b[10] & g[1407];
assign g[2432] = a[10] & g[1408];
assign g[3455] = b[10] & g[1408];
assign g[2433] = a[10] & g[1409];
assign g[3456] = b[10] & g[1409];
assign g[2434] = a[10] & g[1410];
assign g[3457] = b[10] & g[1410];
assign g[2435] = a[10] & g[1411];
assign g[3458] = b[10] & g[1411];
assign g[2436] = a[10] & g[1412];
assign g[3459] = b[10] & g[1412];
assign g[2437] = a[10] & g[1413];
assign g[3460] = b[10] & g[1413];
assign g[2438] = a[10] & g[1414];
assign g[3461] = b[10] & g[1414];
assign g[2439] = a[10] & g[1415];
assign g[3462] = b[10] & g[1415];
assign g[2440] = a[10] & g[1416];
assign g[3463] = b[10] & g[1416];
assign g[2441] = a[10] & g[1417];
assign g[3464] = b[10] & g[1417];
assign g[2442] = a[10] & g[1418];
assign g[3465] = b[10] & g[1418];
assign g[2443] = a[10] & g[1419];
assign g[3466] = b[10] & g[1419];
assign g[2444] = a[10] & g[1420];
assign g[3467] = b[10] & g[1420];
assign g[2445] = a[10] & g[1421];
assign g[3468] = b[10] & g[1421];
assign g[2446] = a[10] & g[1422];
assign g[3469] = b[10] & g[1422];
assign g[2447] = a[10] & g[1423];
assign g[3470] = b[10] & g[1423];
assign g[2448] = a[10] & g[1424];
assign g[3471] = b[10] & g[1424];
assign g[2449] = a[10] & g[1425];
assign g[3472] = b[10] & g[1425];
assign g[2450] = a[10] & g[1426];
assign g[3473] = b[10] & g[1426];
assign g[2451] = a[10] & g[1427];
assign g[3474] = b[10] & g[1427];
assign g[2452] = a[10] & g[1428];
assign g[3475] = b[10] & g[1428];
assign g[2453] = a[10] & g[1429];
assign g[3476] = b[10] & g[1429];
assign g[2454] = a[10] & g[1430];
assign g[3477] = b[10] & g[1430];
assign g[2455] = a[10] & g[1431];
assign g[3478] = b[10] & g[1431];
assign g[2456] = a[10] & g[1432];
assign g[3479] = b[10] & g[1432];
assign g[2457] = a[10] & g[1433];
assign g[3480] = b[10] & g[1433];
assign g[2458] = a[10] & g[1434];
assign g[3481] = b[10] & g[1434];
assign g[2459] = a[10] & g[1435];
assign g[3482] = b[10] & g[1435];
assign g[2460] = a[10] & g[1436];
assign g[3483] = b[10] & g[1436];
assign g[2461] = a[10] & g[1437];
assign g[3484] = b[10] & g[1437];
assign g[2462] = a[10] & g[1438];
assign g[3485] = b[10] & g[1438];
assign g[2463] = a[10] & g[1439];
assign g[3486] = b[10] & g[1439];
assign g[2464] = a[10] & g[1440];
assign g[3487] = b[10] & g[1440];
assign g[2465] = a[10] & g[1441];
assign g[3488] = b[10] & g[1441];
assign g[2466] = a[10] & g[1442];
assign g[3489] = b[10] & g[1442];
assign g[2467] = a[10] & g[1443];
assign g[3490] = b[10] & g[1443];
assign g[2468] = a[10] & g[1444];
assign g[3491] = b[10] & g[1444];
assign g[2469] = a[10] & g[1445];
assign g[3492] = b[10] & g[1445];
assign g[2470] = a[10] & g[1446];
assign g[3493] = b[10] & g[1446];
assign g[2471] = a[10] & g[1447];
assign g[3494] = b[10] & g[1447];
assign g[2472] = a[10] & g[1448];
assign g[3495] = b[10] & g[1448];
assign g[2473] = a[10] & g[1449];
assign g[3496] = b[10] & g[1449];
assign g[2474] = a[10] & g[1450];
assign g[3497] = b[10] & g[1450];
assign g[2475] = a[10] & g[1451];
assign g[3498] = b[10] & g[1451];
assign g[2476] = a[10] & g[1452];
assign g[3499] = b[10] & g[1452];
assign g[2477] = a[10] & g[1453];
assign g[3500] = b[10] & g[1453];
assign g[2478] = a[10] & g[1454];
assign g[3501] = b[10] & g[1454];
assign g[2479] = a[10] & g[1455];
assign g[3502] = b[10] & g[1455];
assign g[2480] = a[10] & g[1456];
assign g[3503] = b[10] & g[1456];
assign g[2481] = a[10] & g[1457];
assign g[3504] = b[10] & g[1457];
assign g[2482] = a[10] & g[1458];
assign g[3505] = b[10] & g[1458];
assign g[2483] = a[10] & g[1459];
assign g[3506] = b[10] & g[1459];
assign g[2484] = a[10] & g[1460];
assign g[3507] = b[10] & g[1460];
assign g[2485] = a[10] & g[1461];
assign g[3508] = b[10] & g[1461];
assign g[2486] = a[10] & g[1462];
assign g[3509] = b[10] & g[1462];
assign g[2487] = a[10] & g[1463];
assign g[3510] = b[10] & g[1463];
assign g[2488] = a[10] & g[1464];
assign g[3511] = b[10] & g[1464];
assign g[2489] = a[10] & g[1465];
assign g[3512] = b[10] & g[1465];
assign g[2490] = a[10] & g[1466];
assign g[3513] = b[10] & g[1466];
assign g[2491] = a[10] & g[1467];
assign g[3514] = b[10] & g[1467];
assign g[2492] = a[10] & g[1468];
assign g[3515] = b[10] & g[1468];
assign g[2493] = a[10] & g[1469];
assign g[3516] = b[10] & g[1469];
assign g[2494] = a[10] & g[1470];
assign g[3517] = b[10] & g[1470];
assign g[2495] = a[10] & g[1471];
assign g[3518] = b[10] & g[1471];
assign g[2496] = a[10] & g[1472];
assign g[3519] = b[10] & g[1472];
assign g[2497] = a[10] & g[1473];
assign g[3520] = b[10] & g[1473];
assign g[2498] = a[10] & g[1474];
assign g[3521] = b[10] & g[1474];
assign g[2499] = a[10] & g[1475];
assign g[3522] = b[10] & g[1475];
assign g[2500] = a[10] & g[1476];
assign g[3523] = b[10] & g[1476];
assign g[2501] = a[10] & g[1477];
assign g[3524] = b[10] & g[1477];
assign g[2502] = a[10] & g[1478];
assign g[3525] = b[10] & g[1478];
assign g[2503] = a[10] & g[1479];
assign g[3526] = b[10] & g[1479];
assign g[2504] = a[10] & g[1480];
assign g[3527] = b[10] & g[1480];
assign g[2505] = a[10] & g[1481];
assign g[3528] = b[10] & g[1481];
assign g[2506] = a[10] & g[1482];
assign g[3529] = b[10] & g[1482];
assign g[2507] = a[10] & g[1483];
assign g[3530] = b[10] & g[1483];
assign g[2508] = a[10] & g[1484];
assign g[3531] = b[10] & g[1484];
assign g[2509] = a[10] & g[1485];
assign g[3532] = b[10] & g[1485];
assign g[2510] = a[10] & g[1486];
assign g[3533] = b[10] & g[1486];
assign g[2511] = a[10] & g[1487];
assign g[3534] = b[10] & g[1487];
assign g[2512] = a[10] & g[1488];
assign g[3535] = b[10] & g[1488];
assign g[2513] = a[10] & g[1489];
assign g[3536] = b[10] & g[1489];
assign g[2514] = a[10] & g[1490];
assign g[3537] = b[10] & g[1490];
assign g[2515] = a[10] & g[1491];
assign g[3538] = b[10] & g[1491];
assign g[2516] = a[10] & g[1492];
assign g[3539] = b[10] & g[1492];
assign g[2517] = a[10] & g[1493];
assign g[3540] = b[10] & g[1493];
assign g[2518] = a[10] & g[1494];
assign g[3541] = b[10] & g[1494];
assign g[2519] = a[10] & g[1495];
assign g[3542] = b[10] & g[1495];
assign g[2520] = a[10] & g[1496];
assign g[3543] = b[10] & g[1496];
assign g[2521] = a[10] & g[1497];
assign g[3544] = b[10] & g[1497];
assign g[2522] = a[10] & g[1498];
assign g[3545] = b[10] & g[1498];
assign g[2523] = a[10] & g[1499];
assign g[3546] = b[10] & g[1499];
assign g[2524] = a[10] & g[1500];
assign g[3547] = b[10] & g[1500];
assign g[2525] = a[10] & g[1501];
assign g[3548] = b[10] & g[1501];
assign g[2526] = a[10] & g[1502];
assign g[3549] = b[10] & g[1502];
assign g[2527] = a[10] & g[1503];
assign g[3550] = b[10] & g[1503];
assign g[2528] = a[10] & g[1504];
assign g[3551] = b[10] & g[1504];
assign g[2529] = a[10] & g[1505];
assign g[3552] = b[10] & g[1505];
assign g[2530] = a[10] & g[1506];
assign g[3553] = b[10] & g[1506];
assign g[2531] = a[10] & g[1507];
assign g[3554] = b[10] & g[1507];
assign g[2532] = a[10] & g[1508];
assign g[3555] = b[10] & g[1508];
assign g[2533] = a[10] & g[1509];
assign g[3556] = b[10] & g[1509];
assign g[2534] = a[10] & g[1510];
assign g[3557] = b[10] & g[1510];
assign g[2535] = a[10] & g[1511];
assign g[3558] = b[10] & g[1511];
assign g[2536] = a[10] & g[1512];
assign g[3559] = b[10] & g[1512];
assign g[2537] = a[10] & g[1513];
assign g[3560] = b[10] & g[1513];
assign g[2538] = a[10] & g[1514];
assign g[3561] = b[10] & g[1514];
assign g[2539] = a[10] & g[1515];
assign g[3562] = b[10] & g[1515];
assign g[2540] = a[10] & g[1516];
assign g[3563] = b[10] & g[1516];
assign g[2541] = a[10] & g[1517];
assign g[3564] = b[10] & g[1517];
assign g[2542] = a[10] & g[1518];
assign g[3565] = b[10] & g[1518];
assign g[2543] = a[10] & g[1519];
assign g[3566] = b[10] & g[1519];
assign g[2544] = a[10] & g[1520];
assign g[3567] = b[10] & g[1520];
assign g[2545] = a[10] & g[1521];
assign g[3568] = b[10] & g[1521];
assign g[2546] = a[10] & g[1522];
assign g[3569] = b[10] & g[1522];
assign g[2547] = a[10] & g[1523];
assign g[3570] = b[10] & g[1523];
assign g[2548] = a[10] & g[1524];
assign g[3571] = b[10] & g[1524];
assign g[2549] = a[10] & g[1525];
assign g[3572] = b[10] & g[1525];
assign g[2550] = a[10] & g[1526];
assign g[3573] = b[10] & g[1526];
assign g[2551] = a[10] & g[1527];
assign g[3574] = b[10] & g[1527];
assign g[2552] = a[10] & g[1528];
assign g[3575] = b[10] & g[1528];
assign g[2553] = a[10] & g[1529];
assign g[3576] = b[10] & g[1529];
assign g[2554] = a[10] & g[1530];
assign g[3577] = b[10] & g[1530];
assign g[2555] = a[10] & g[1531];
assign g[3578] = b[10] & g[1531];
assign g[2556] = a[10] & g[1532];
assign g[3579] = b[10] & g[1532];
assign g[2557] = a[10] & g[1533];
assign g[3580] = b[10] & g[1533];
assign g[2558] = a[10] & g[1534];
assign g[3581] = b[10] & g[1534];
assign g[2559] = a[10] & g[1535];
assign g[3582] = b[10] & g[1535];
assign g[2560] = a[10] & g[1536];
assign g[3583] = b[10] & g[1536];
assign g[2561] = a[10] & g[1537];
assign g[3584] = b[10] & g[1537];
assign g[2562] = a[10] & g[1538];
assign g[3585] = b[10] & g[1538];
assign g[2563] = a[10] & g[1539];
assign g[3586] = b[10] & g[1539];
assign g[2564] = a[10] & g[1540];
assign g[3587] = b[10] & g[1540];
assign g[2565] = a[10] & g[1541];
assign g[3588] = b[10] & g[1541];
assign g[2566] = a[10] & g[1542];
assign g[3589] = b[10] & g[1542];
assign g[2567] = a[10] & g[1543];
assign g[3590] = b[10] & g[1543];
assign g[2568] = a[10] & g[1544];
assign g[3591] = b[10] & g[1544];
assign g[2569] = a[10] & g[1545];
assign g[3592] = b[10] & g[1545];
assign g[2570] = a[10] & g[1546];
assign g[3593] = b[10] & g[1546];
assign g[2571] = a[10] & g[1547];
assign g[3594] = b[10] & g[1547];
assign g[2572] = a[10] & g[1548];
assign g[3595] = b[10] & g[1548];
assign g[2573] = a[10] & g[1549];
assign g[3596] = b[10] & g[1549];
assign g[2574] = a[10] & g[1550];
assign g[3597] = b[10] & g[1550];
assign g[2575] = a[10] & g[1551];
assign g[3598] = b[10] & g[1551];
assign g[2576] = a[10] & g[1552];
assign g[3599] = b[10] & g[1552];
assign g[2577] = a[10] & g[1553];
assign g[3600] = b[10] & g[1553];
assign g[2578] = a[10] & g[1554];
assign g[3601] = b[10] & g[1554];
assign g[2579] = a[10] & g[1555];
assign g[3602] = b[10] & g[1555];
assign g[2580] = a[10] & g[1556];
assign g[3603] = b[10] & g[1556];
assign g[2581] = a[10] & g[1557];
assign g[3604] = b[10] & g[1557];
assign g[2582] = a[10] & g[1558];
assign g[3605] = b[10] & g[1558];
assign g[2583] = a[10] & g[1559];
assign g[3606] = b[10] & g[1559];
assign g[2584] = a[10] & g[1560];
assign g[3607] = b[10] & g[1560];
assign g[2585] = a[10] & g[1561];
assign g[3608] = b[10] & g[1561];
assign g[2586] = a[10] & g[1562];
assign g[3609] = b[10] & g[1562];
assign g[2587] = a[10] & g[1563];
assign g[3610] = b[10] & g[1563];
assign g[2588] = a[10] & g[1564];
assign g[3611] = b[10] & g[1564];
assign g[2589] = a[10] & g[1565];
assign g[3612] = b[10] & g[1565];
assign g[2590] = a[10] & g[1566];
assign g[3613] = b[10] & g[1566];
assign g[2591] = a[10] & g[1567];
assign g[3614] = b[10] & g[1567];
assign g[2592] = a[10] & g[1568];
assign g[3615] = b[10] & g[1568];
assign g[2593] = a[10] & g[1569];
assign g[3616] = b[10] & g[1569];
assign g[2594] = a[10] & g[1570];
assign g[3617] = b[10] & g[1570];
assign g[2595] = a[10] & g[1571];
assign g[3618] = b[10] & g[1571];
assign g[2596] = a[10] & g[1572];
assign g[3619] = b[10] & g[1572];
assign g[2597] = a[10] & g[1573];
assign g[3620] = b[10] & g[1573];
assign g[2598] = a[10] & g[1574];
assign g[3621] = b[10] & g[1574];
assign g[2599] = a[10] & g[1575];
assign g[3622] = b[10] & g[1575];
assign g[2600] = a[10] & g[1576];
assign g[3623] = b[10] & g[1576];
assign g[2601] = a[10] & g[1577];
assign g[3624] = b[10] & g[1577];
assign g[2602] = a[10] & g[1578];
assign g[3625] = b[10] & g[1578];
assign g[2603] = a[10] & g[1579];
assign g[3626] = b[10] & g[1579];
assign g[2604] = a[10] & g[1580];
assign g[3627] = b[10] & g[1580];
assign g[2605] = a[10] & g[1581];
assign g[3628] = b[10] & g[1581];
assign g[2606] = a[10] & g[1582];
assign g[3629] = b[10] & g[1582];
assign g[2607] = a[10] & g[1583];
assign g[3630] = b[10] & g[1583];
assign g[2608] = a[10] & g[1584];
assign g[3631] = b[10] & g[1584];
assign g[2609] = a[10] & g[1585];
assign g[3632] = b[10] & g[1585];
assign g[2610] = a[10] & g[1586];
assign g[3633] = b[10] & g[1586];
assign g[2611] = a[10] & g[1587];
assign g[3634] = b[10] & g[1587];
assign g[2612] = a[10] & g[1588];
assign g[3635] = b[10] & g[1588];
assign g[2613] = a[10] & g[1589];
assign g[3636] = b[10] & g[1589];
assign g[2614] = a[10] & g[1590];
assign g[3637] = b[10] & g[1590];
assign g[2615] = a[10] & g[1591];
assign g[3638] = b[10] & g[1591];
assign g[2616] = a[10] & g[1592];
assign g[3639] = b[10] & g[1592];
assign g[2617] = a[10] & g[1593];
assign g[3640] = b[10] & g[1593];
assign g[2618] = a[10] & g[1594];
assign g[3641] = b[10] & g[1594];
assign g[2619] = a[10] & g[1595];
assign g[3642] = b[10] & g[1595];
assign g[2620] = a[10] & g[1596];
assign g[3643] = b[10] & g[1596];
assign g[2621] = a[10] & g[1597];
assign g[3644] = b[10] & g[1597];
assign g[2622] = a[10] & g[1598];
assign g[3645] = b[10] & g[1598];
assign g[2623] = a[10] & g[1599];
assign g[3646] = b[10] & g[1599];
assign g[2624] = a[10] & g[1600];
assign g[3647] = b[10] & g[1600];
assign g[2625] = a[10] & g[1601];
assign g[3648] = b[10] & g[1601];
assign g[2626] = a[10] & g[1602];
assign g[3649] = b[10] & g[1602];
assign g[2627] = a[10] & g[1603];
assign g[3650] = b[10] & g[1603];
assign g[2628] = a[10] & g[1604];
assign g[3651] = b[10] & g[1604];
assign g[2629] = a[10] & g[1605];
assign g[3652] = b[10] & g[1605];
assign g[2630] = a[10] & g[1606];
assign g[3653] = b[10] & g[1606];
assign g[2631] = a[10] & g[1607];
assign g[3654] = b[10] & g[1607];
assign g[2632] = a[10] & g[1608];
assign g[3655] = b[10] & g[1608];
assign g[2633] = a[10] & g[1609];
assign g[3656] = b[10] & g[1609];
assign g[2634] = a[10] & g[1610];
assign g[3657] = b[10] & g[1610];
assign g[2635] = a[10] & g[1611];
assign g[3658] = b[10] & g[1611];
assign g[2636] = a[10] & g[1612];
assign g[3659] = b[10] & g[1612];
assign g[2637] = a[10] & g[1613];
assign g[3660] = b[10] & g[1613];
assign g[2638] = a[10] & g[1614];
assign g[3661] = b[10] & g[1614];
assign g[2639] = a[10] & g[1615];
assign g[3662] = b[10] & g[1615];
assign g[2640] = a[10] & g[1616];
assign g[3663] = b[10] & g[1616];
assign g[2641] = a[10] & g[1617];
assign g[3664] = b[10] & g[1617];
assign g[2642] = a[10] & g[1618];
assign g[3665] = b[10] & g[1618];
assign g[2643] = a[10] & g[1619];
assign g[3666] = b[10] & g[1619];
assign g[2644] = a[10] & g[1620];
assign g[3667] = b[10] & g[1620];
assign g[2645] = a[10] & g[1621];
assign g[3668] = b[10] & g[1621];
assign g[2646] = a[10] & g[1622];
assign g[3669] = b[10] & g[1622];
assign g[2647] = a[10] & g[1623];
assign g[3670] = b[10] & g[1623];
assign g[2648] = a[10] & g[1624];
assign g[3671] = b[10] & g[1624];
assign g[2649] = a[10] & g[1625];
assign g[3672] = b[10] & g[1625];
assign g[2650] = a[10] & g[1626];
assign g[3673] = b[10] & g[1626];
assign g[2651] = a[10] & g[1627];
assign g[3674] = b[10] & g[1627];
assign g[2652] = a[10] & g[1628];
assign g[3675] = b[10] & g[1628];
assign g[2653] = a[10] & g[1629];
assign g[3676] = b[10] & g[1629];
assign g[2654] = a[10] & g[1630];
assign g[3677] = b[10] & g[1630];
assign g[2655] = a[10] & g[1631];
assign g[3678] = b[10] & g[1631];
assign g[2656] = a[10] & g[1632];
assign g[3679] = b[10] & g[1632];
assign g[2657] = a[10] & g[1633];
assign g[3680] = b[10] & g[1633];
assign g[2658] = a[10] & g[1634];
assign g[3681] = b[10] & g[1634];
assign g[2659] = a[10] & g[1635];
assign g[3682] = b[10] & g[1635];
assign g[2660] = a[10] & g[1636];
assign g[3683] = b[10] & g[1636];
assign g[2661] = a[10] & g[1637];
assign g[3684] = b[10] & g[1637];
assign g[2662] = a[10] & g[1638];
assign g[3685] = b[10] & g[1638];
assign g[2663] = a[10] & g[1639];
assign g[3686] = b[10] & g[1639];
assign g[2664] = a[10] & g[1640];
assign g[3687] = b[10] & g[1640];
assign g[2665] = a[10] & g[1641];
assign g[3688] = b[10] & g[1641];
assign g[2666] = a[10] & g[1642];
assign g[3689] = b[10] & g[1642];
assign g[2667] = a[10] & g[1643];
assign g[3690] = b[10] & g[1643];
assign g[2668] = a[10] & g[1644];
assign g[3691] = b[10] & g[1644];
assign g[2669] = a[10] & g[1645];
assign g[3692] = b[10] & g[1645];
assign g[2670] = a[10] & g[1646];
assign g[3693] = b[10] & g[1646];
assign g[2671] = a[10] & g[1647];
assign g[3694] = b[10] & g[1647];
assign g[2672] = a[10] & g[1648];
assign g[3695] = b[10] & g[1648];
assign g[2673] = a[10] & g[1649];
assign g[3696] = b[10] & g[1649];
assign g[2674] = a[10] & g[1650];
assign g[3697] = b[10] & g[1650];
assign g[2675] = a[10] & g[1651];
assign g[3698] = b[10] & g[1651];
assign g[2676] = a[10] & g[1652];
assign g[3699] = b[10] & g[1652];
assign g[2677] = a[10] & g[1653];
assign g[3700] = b[10] & g[1653];
assign g[2678] = a[10] & g[1654];
assign g[3701] = b[10] & g[1654];
assign g[2679] = a[10] & g[1655];
assign g[3702] = b[10] & g[1655];
assign g[2680] = a[10] & g[1656];
assign g[3703] = b[10] & g[1656];
assign g[2681] = a[10] & g[1657];
assign g[3704] = b[10] & g[1657];
assign g[2682] = a[10] & g[1658];
assign g[3705] = b[10] & g[1658];
assign g[2683] = a[10] & g[1659];
assign g[3706] = b[10] & g[1659];
assign g[2684] = a[10] & g[1660];
assign g[3707] = b[10] & g[1660];
assign g[2685] = a[10] & g[1661];
assign g[3708] = b[10] & g[1661];
assign g[2686] = a[10] & g[1662];
assign g[3709] = b[10] & g[1662];
assign g[2687] = a[10] & g[1663];
assign g[3710] = b[10] & g[1663];
assign g[2688] = a[10] & g[1664];
assign g[3711] = b[10] & g[1664];
assign g[2689] = a[10] & g[1665];
assign g[3712] = b[10] & g[1665];
assign g[2690] = a[10] & g[1666];
assign g[3713] = b[10] & g[1666];
assign g[2691] = a[10] & g[1667];
assign g[3714] = b[10] & g[1667];
assign g[2692] = a[10] & g[1668];
assign g[3715] = b[10] & g[1668];
assign g[2693] = a[10] & g[1669];
assign g[3716] = b[10] & g[1669];
assign g[2694] = a[10] & g[1670];
assign g[3717] = b[10] & g[1670];
assign g[2695] = a[10] & g[1671];
assign g[3718] = b[10] & g[1671];
assign g[2696] = a[10] & g[1672];
assign g[3719] = b[10] & g[1672];
assign g[2697] = a[10] & g[1673];
assign g[3720] = b[10] & g[1673];
assign g[2698] = a[10] & g[1674];
assign g[3721] = b[10] & g[1674];
assign g[2699] = a[10] & g[1675];
assign g[3722] = b[10] & g[1675];
assign g[2700] = a[10] & g[1676];
assign g[3723] = b[10] & g[1676];
assign g[2701] = a[10] & g[1677];
assign g[3724] = b[10] & g[1677];
assign g[2702] = a[10] & g[1678];
assign g[3725] = b[10] & g[1678];
assign g[2703] = a[10] & g[1679];
assign g[3726] = b[10] & g[1679];
assign g[2704] = a[10] & g[1680];
assign g[3727] = b[10] & g[1680];
assign g[2705] = a[10] & g[1681];
assign g[3728] = b[10] & g[1681];
assign g[2706] = a[10] & g[1682];
assign g[3729] = b[10] & g[1682];
assign g[2707] = a[10] & g[1683];
assign g[3730] = b[10] & g[1683];
assign g[2708] = a[10] & g[1684];
assign g[3731] = b[10] & g[1684];
assign g[2709] = a[10] & g[1685];
assign g[3732] = b[10] & g[1685];
assign g[2710] = a[10] & g[1686];
assign g[3733] = b[10] & g[1686];
assign g[2711] = a[10] & g[1687];
assign g[3734] = b[10] & g[1687];
assign g[2712] = a[10] & g[1688];
assign g[3735] = b[10] & g[1688];
assign g[2713] = a[10] & g[1689];
assign g[3736] = b[10] & g[1689];
assign g[2714] = a[10] & g[1690];
assign g[3737] = b[10] & g[1690];
assign g[2715] = a[10] & g[1691];
assign g[3738] = b[10] & g[1691];
assign g[2716] = a[10] & g[1692];
assign g[3739] = b[10] & g[1692];
assign g[2717] = a[10] & g[1693];
assign g[3740] = b[10] & g[1693];
assign g[2718] = a[10] & g[1694];
assign g[3741] = b[10] & g[1694];
assign g[2719] = a[10] & g[1695];
assign g[3742] = b[10] & g[1695];
assign g[2720] = a[10] & g[1696];
assign g[3743] = b[10] & g[1696];
assign g[2721] = a[10] & g[1697];
assign g[3744] = b[10] & g[1697];
assign g[2722] = a[10] & g[1698];
assign g[3745] = b[10] & g[1698];
assign g[2723] = a[10] & g[1699];
assign g[3746] = b[10] & g[1699];
assign g[2724] = a[10] & g[1700];
assign g[3747] = b[10] & g[1700];
assign g[2725] = a[10] & g[1701];
assign g[3748] = b[10] & g[1701];
assign g[2726] = a[10] & g[1702];
assign g[3749] = b[10] & g[1702];
assign g[2727] = a[10] & g[1703];
assign g[3750] = b[10] & g[1703];
assign g[2728] = a[10] & g[1704];
assign g[3751] = b[10] & g[1704];
assign g[2729] = a[10] & g[1705];
assign g[3752] = b[10] & g[1705];
assign g[2730] = a[10] & g[1706];
assign g[3753] = b[10] & g[1706];
assign g[2731] = a[10] & g[1707];
assign g[3754] = b[10] & g[1707];
assign g[2732] = a[10] & g[1708];
assign g[3755] = b[10] & g[1708];
assign g[2733] = a[10] & g[1709];
assign g[3756] = b[10] & g[1709];
assign g[2734] = a[10] & g[1710];
assign g[3757] = b[10] & g[1710];
assign g[2735] = a[10] & g[1711];
assign g[3758] = b[10] & g[1711];
assign g[2736] = a[10] & g[1712];
assign g[3759] = b[10] & g[1712];
assign g[2737] = a[10] & g[1713];
assign g[3760] = b[10] & g[1713];
assign g[2738] = a[10] & g[1714];
assign g[3761] = b[10] & g[1714];
assign g[2739] = a[10] & g[1715];
assign g[3762] = b[10] & g[1715];
assign g[2740] = a[10] & g[1716];
assign g[3763] = b[10] & g[1716];
assign g[2741] = a[10] & g[1717];
assign g[3764] = b[10] & g[1717];
assign g[2742] = a[10] & g[1718];
assign g[3765] = b[10] & g[1718];
assign g[2743] = a[10] & g[1719];
assign g[3766] = b[10] & g[1719];
assign g[2744] = a[10] & g[1720];
assign g[3767] = b[10] & g[1720];
assign g[2745] = a[10] & g[1721];
assign g[3768] = b[10] & g[1721];
assign g[2746] = a[10] & g[1722];
assign g[3769] = b[10] & g[1722];
assign g[2747] = a[10] & g[1723];
assign g[3770] = b[10] & g[1723];
assign g[2748] = a[10] & g[1724];
assign g[3771] = b[10] & g[1724];
assign g[2749] = a[10] & g[1725];
assign g[3772] = b[10] & g[1725];
assign g[2750] = a[10] & g[1726];
assign g[3773] = b[10] & g[1726];
assign g[2751] = a[10] & g[1727];
assign g[3774] = b[10] & g[1727];
assign g[2752] = a[10] & g[1728];
assign g[3775] = b[10] & g[1728];
assign g[2753] = a[10] & g[1729];
assign g[3776] = b[10] & g[1729];
assign g[2754] = a[10] & g[1730];
assign g[3777] = b[10] & g[1730];
assign g[2755] = a[10] & g[1731];
assign g[3778] = b[10] & g[1731];
assign g[2756] = a[10] & g[1732];
assign g[3779] = b[10] & g[1732];
assign g[2757] = a[10] & g[1733];
assign g[3780] = b[10] & g[1733];
assign g[2758] = a[10] & g[1734];
assign g[3781] = b[10] & g[1734];
assign g[2759] = a[10] & g[1735];
assign g[3782] = b[10] & g[1735];
assign g[2760] = a[10] & g[1736];
assign g[3783] = b[10] & g[1736];
assign g[2761] = a[10] & g[1737];
assign g[3784] = b[10] & g[1737];
assign g[2762] = a[10] & g[1738];
assign g[3785] = b[10] & g[1738];
assign g[2763] = a[10] & g[1739];
assign g[3786] = b[10] & g[1739];
assign g[2764] = a[10] & g[1740];
assign g[3787] = b[10] & g[1740];
assign g[2765] = a[10] & g[1741];
assign g[3788] = b[10] & g[1741];
assign g[2766] = a[10] & g[1742];
assign g[3789] = b[10] & g[1742];
assign g[2767] = a[10] & g[1743];
assign g[3790] = b[10] & g[1743];
assign g[2768] = a[10] & g[1744];
assign g[3791] = b[10] & g[1744];
assign g[2769] = a[10] & g[1745];
assign g[3792] = b[10] & g[1745];
assign g[2770] = a[10] & g[1746];
assign g[3793] = b[10] & g[1746];
assign g[2771] = a[10] & g[1747];
assign g[3794] = b[10] & g[1747];
assign g[2772] = a[10] & g[1748];
assign g[3795] = b[10] & g[1748];
assign g[2773] = a[10] & g[1749];
assign g[3796] = b[10] & g[1749];
assign g[2774] = a[10] & g[1750];
assign g[3797] = b[10] & g[1750];
assign g[2775] = a[10] & g[1751];
assign g[3798] = b[10] & g[1751];
assign g[2776] = a[10] & g[1752];
assign g[3799] = b[10] & g[1752];
assign g[2777] = a[10] & g[1753];
assign g[3800] = b[10] & g[1753];
assign g[2778] = a[10] & g[1754];
assign g[3801] = b[10] & g[1754];
assign g[2779] = a[10] & g[1755];
assign g[3802] = b[10] & g[1755];
assign g[2780] = a[10] & g[1756];
assign g[3803] = b[10] & g[1756];
assign g[2781] = a[10] & g[1757];
assign g[3804] = b[10] & g[1757];
assign g[2782] = a[10] & g[1758];
assign g[3805] = b[10] & g[1758];
assign g[2783] = a[10] & g[1759];
assign g[3806] = b[10] & g[1759];
assign g[2784] = a[10] & g[1760];
assign g[3807] = b[10] & g[1760];
assign g[2785] = a[10] & g[1761];
assign g[3808] = b[10] & g[1761];
assign g[2786] = a[10] & g[1762];
assign g[3809] = b[10] & g[1762];
assign g[2787] = a[10] & g[1763];
assign g[3810] = b[10] & g[1763];
assign g[2788] = a[10] & g[1764];
assign g[3811] = b[10] & g[1764];
assign g[2789] = a[10] & g[1765];
assign g[3812] = b[10] & g[1765];
assign g[2790] = a[10] & g[1766];
assign g[3813] = b[10] & g[1766];
assign g[2791] = a[10] & g[1767];
assign g[3814] = b[10] & g[1767];
assign g[2792] = a[10] & g[1768];
assign g[3815] = b[10] & g[1768];
assign g[2793] = a[10] & g[1769];
assign g[3816] = b[10] & g[1769];
assign g[2794] = a[10] & g[1770];
assign g[3817] = b[10] & g[1770];
assign g[2795] = a[10] & g[1771];
assign g[3818] = b[10] & g[1771];
assign g[2796] = a[10] & g[1772];
assign g[3819] = b[10] & g[1772];
assign g[2797] = a[10] & g[1773];
assign g[3820] = b[10] & g[1773];
assign g[2798] = a[10] & g[1774];
assign g[3821] = b[10] & g[1774];
assign g[2799] = a[10] & g[1775];
assign g[3822] = b[10] & g[1775];
assign g[2800] = a[10] & g[1776];
assign g[3823] = b[10] & g[1776];
assign g[2801] = a[10] & g[1777];
assign g[3824] = b[10] & g[1777];
assign g[2802] = a[10] & g[1778];
assign g[3825] = b[10] & g[1778];
assign g[2803] = a[10] & g[1779];
assign g[3826] = b[10] & g[1779];
assign g[2804] = a[10] & g[1780];
assign g[3827] = b[10] & g[1780];
assign g[2805] = a[10] & g[1781];
assign g[3828] = b[10] & g[1781];
assign g[2806] = a[10] & g[1782];
assign g[3829] = b[10] & g[1782];
assign g[2807] = a[10] & g[1783];
assign g[3830] = b[10] & g[1783];
assign g[2808] = a[10] & g[1784];
assign g[3831] = b[10] & g[1784];
assign g[2809] = a[10] & g[1785];
assign g[3832] = b[10] & g[1785];
assign g[2810] = a[10] & g[1786];
assign g[3833] = b[10] & g[1786];
assign g[2811] = a[10] & g[1787];
assign g[3834] = b[10] & g[1787];
assign g[2812] = a[10] & g[1788];
assign g[3835] = b[10] & g[1788];
assign g[2813] = a[10] & g[1789];
assign g[3836] = b[10] & g[1789];
assign g[2814] = a[10] & g[1790];
assign g[3837] = b[10] & g[1790];
assign g[2815] = a[10] & g[1791];
assign g[3838] = b[10] & g[1791];
assign g[2816] = a[10] & g[1792];
assign g[3839] = b[10] & g[1792];
assign g[2817] = a[10] & g[1793];
assign g[3840] = b[10] & g[1793];
assign g[2818] = a[10] & g[1794];
assign g[3841] = b[10] & g[1794];
assign g[2819] = a[10] & g[1795];
assign g[3842] = b[10] & g[1795];
assign g[2820] = a[10] & g[1796];
assign g[3843] = b[10] & g[1796];
assign g[2821] = a[10] & g[1797];
assign g[3844] = b[10] & g[1797];
assign g[2822] = a[10] & g[1798];
assign g[3845] = b[10] & g[1798];
assign g[2823] = a[10] & g[1799];
assign g[3846] = b[10] & g[1799];
assign g[2824] = a[10] & g[1800];
assign g[3847] = b[10] & g[1800];
assign g[2825] = a[10] & g[1801];
assign g[3848] = b[10] & g[1801];
assign g[2826] = a[10] & g[1802];
assign g[3849] = b[10] & g[1802];
assign g[2827] = a[10] & g[1803];
assign g[3850] = b[10] & g[1803];
assign g[2828] = a[10] & g[1804];
assign g[3851] = b[10] & g[1804];
assign g[2829] = a[10] & g[1805];
assign g[3852] = b[10] & g[1805];
assign g[2830] = a[10] & g[1806];
assign g[3853] = b[10] & g[1806];
assign g[2831] = a[10] & g[1807];
assign g[3854] = b[10] & g[1807];
assign g[2832] = a[10] & g[1808];
assign g[3855] = b[10] & g[1808];
assign g[2833] = a[10] & g[1809];
assign g[3856] = b[10] & g[1809];
assign g[2834] = a[10] & g[1810];
assign g[3857] = b[10] & g[1810];
assign g[2835] = a[10] & g[1811];
assign g[3858] = b[10] & g[1811];
assign g[2836] = a[10] & g[1812];
assign g[3859] = b[10] & g[1812];
assign g[2837] = a[10] & g[1813];
assign g[3860] = b[10] & g[1813];
assign g[2838] = a[10] & g[1814];
assign g[3861] = b[10] & g[1814];
assign g[2839] = a[10] & g[1815];
assign g[3862] = b[10] & g[1815];
assign g[2840] = a[10] & g[1816];
assign g[3863] = b[10] & g[1816];
assign g[2841] = a[10] & g[1817];
assign g[3864] = b[10] & g[1817];
assign g[2842] = a[10] & g[1818];
assign g[3865] = b[10] & g[1818];
assign g[2843] = a[10] & g[1819];
assign g[3866] = b[10] & g[1819];
assign g[2844] = a[10] & g[1820];
assign g[3867] = b[10] & g[1820];
assign g[2845] = a[10] & g[1821];
assign g[3868] = b[10] & g[1821];
assign g[2846] = a[10] & g[1822];
assign g[3869] = b[10] & g[1822];
assign g[2847] = a[10] & g[1823];
assign g[3870] = b[10] & g[1823];
assign g[2848] = a[10] & g[1824];
assign g[3871] = b[10] & g[1824];
assign g[2849] = a[10] & g[1825];
assign g[3872] = b[10] & g[1825];
assign g[2850] = a[10] & g[1826];
assign g[3873] = b[10] & g[1826];
assign g[2851] = a[10] & g[1827];
assign g[3874] = b[10] & g[1827];
assign g[2852] = a[10] & g[1828];
assign g[3875] = b[10] & g[1828];
assign g[2853] = a[10] & g[1829];
assign g[3876] = b[10] & g[1829];
assign g[2854] = a[10] & g[1830];
assign g[3877] = b[10] & g[1830];
assign g[2855] = a[10] & g[1831];
assign g[3878] = b[10] & g[1831];
assign g[2856] = a[10] & g[1832];
assign g[3879] = b[10] & g[1832];
assign g[2857] = a[10] & g[1833];
assign g[3880] = b[10] & g[1833];
assign g[2858] = a[10] & g[1834];
assign g[3881] = b[10] & g[1834];
assign g[2859] = a[10] & g[1835];
assign g[3882] = b[10] & g[1835];
assign g[2860] = a[10] & g[1836];
assign g[3883] = b[10] & g[1836];
assign g[2861] = a[10] & g[1837];
assign g[3884] = b[10] & g[1837];
assign g[2862] = a[10] & g[1838];
assign g[3885] = b[10] & g[1838];
assign g[2863] = a[10] & g[1839];
assign g[3886] = b[10] & g[1839];
assign g[2864] = a[10] & g[1840];
assign g[3887] = b[10] & g[1840];
assign g[2865] = a[10] & g[1841];
assign g[3888] = b[10] & g[1841];
assign g[2866] = a[10] & g[1842];
assign g[3889] = b[10] & g[1842];
assign g[2867] = a[10] & g[1843];
assign g[3890] = b[10] & g[1843];
assign g[2868] = a[10] & g[1844];
assign g[3891] = b[10] & g[1844];
assign g[2869] = a[10] & g[1845];
assign g[3892] = b[10] & g[1845];
assign g[2870] = a[10] & g[1846];
assign g[3893] = b[10] & g[1846];
assign g[2871] = a[10] & g[1847];
assign g[3894] = b[10] & g[1847];
assign g[2872] = a[10] & g[1848];
assign g[3895] = b[10] & g[1848];
assign g[2873] = a[10] & g[1849];
assign g[3896] = b[10] & g[1849];
assign g[2874] = a[10] & g[1850];
assign g[3897] = b[10] & g[1850];
assign g[2875] = a[10] & g[1851];
assign g[3898] = b[10] & g[1851];
assign g[2876] = a[10] & g[1852];
assign g[3899] = b[10] & g[1852];
assign g[2877] = a[10] & g[1853];
assign g[3900] = b[10] & g[1853];
assign g[2878] = a[10] & g[1854];
assign g[3901] = b[10] & g[1854];
assign g[2879] = a[10] & g[1855];
assign g[3902] = b[10] & g[1855];
assign g[2880] = a[10] & g[1856];
assign g[3903] = b[10] & g[1856];
assign g[2881] = a[10] & g[1857];
assign g[3904] = b[10] & g[1857];
assign g[2882] = a[10] & g[1858];
assign g[3905] = b[10] & g[1858];
assign g[2883] = a[10] & g[1859];
assign g[3906] = b[10] & g[1859];
assign g[2884] = a[10] & g[1860];
assign g[3907] = b[10] & g[1860];
assign g[2885] = a[10] & g[1861];
assign g[3908] = b[10] & g[1861];
assign g[2886] = a[10] & g[1862];
assign g[3909] = b[10] & g[1862];
assign g[2887] = a[10] & g[1863];
assign g[3910] = b[10] & g[1863];
assign g[2888] = a[10] & g[1864];
assign g[3911] = b[10] & g[1864];
assign g[2889] = a[10] & g[1865];
assign g[3912] = b[10] & g[1865];
assign g[2890] = a[10] & g[1866];
assign g[3913] = b[10] & g[1866];
assign g[2891] = a[10] & g[1867];
assign g[3914] = b[10] & g[1867];
assign g[2892] = a[10] & g[1868];
assign g[3915] = b[10] & g[1868];
assign g[2893] = a[10] & g[1869];
assign g[3916] = b[10] & g[1869];
assign g[2894] = a[10] & g[1870];
assign g[3917] = b[10] & g[1870];
assign g[2895] = a[10] & g[1871];
assign g[3918] = b[10] & g[1871];
assign g[2896] = a[10] & g[1872];
assign g[3919] = b[10] & g[1872];
assign g[2897] = a[10] & g[1873];
assign g[3920] = b[10] & g[1873];
assign g[2898] = a[10] & g[1874];
assign g[3921] = b[10] & g[1874];
assign g[2899] = a[10] & g[1875];
assign g[3922] = b[10] & g[1875];
assign g[2900] = a[10] & g[1876];
assign g[3923] = b[10] & g[1876];
assign g[2901] = a[10] & g[1877];
assign g[3924] = b[10] & g[1877];
assign g[2902] = a[10] & g[1878];
assign g[3925] = b[10] & g[1878];
assign g[2903] = a[10] & g[1879];
assign g[3926] = b[10] & g[1879];
assign g[2904] = a[10] & g[1880];
assign g[3927] = b[10] & g[1880];
assign g[2905] = a[10] & g[1881];
assign g[3928] = b[10] & g[1881];
assign g[2906] = a[10] & g[1882];
assign g[3929] = b[10] & g[1882];
assign g[2907] = a[10] & g[1883];
assign g[3930] = b[10] & g[1883];
assign g[2908] = a[10] & g[1884];
assign g[3931] = b[10] & g[1884];
assign g[2909] = a[10] & g[1885];
assign g[3932] = b[10] & g[1885];
assign g[2910] = a[10] & g[1886];
assign g[3933] = b[10] & g[1886];
assign g[2911] = a[10] & g[1887];
assign g[3934] = b[10] & g[1887];
assign g[2912] = a[10] & g[1888];
assign g[3935] = b[10] & g[1888];
assign g[2913] = a[10] & g[1889];
assign g[3936] = b[10] & g[1889];
assign g[2914] = a[10] & g[1890];
assign g[3937] = b[10] & g[1890];
assign g[2915] = a[10] & g[1891];
assign g[3938] = b[10] & g[1891];
assign g[2916] = a[10] & g[1892];
assign g[3939] = b[10] & g[1892];
assign g[2917] = a[10] & g[1893];
assign g[3940] = b[10] & g[1893];
assign g[2918] = a[10] & g[1894];
assign g[3941] = b[10] & g[1894];
assign g[2919] = a[10] & g[1895];
assign g[3942] = b[10] & g[1895];
assign g[2920] = a[10] & g[1896];
assign g[3943] = b[10] & g[1896];
assign g[2921] = a[10] & g[1897];
assign g[3944] = b[10] & g[1897];
assign g[2922] = a[10] & g[1898];
assign g[3945] = b[10] & g[1898];
assign g[2923] = a[10] & g[1899];
assign g[3946] = b[10] & g[1899];
assign g[2924] = a[10] & g[1900];
assign g[3947] = b[10] & g[1900];
assign g[2925] = a[10] & g[1901];
assign g[3948] = b[10] & g[1901];
assign g[2926] = a[10] & g[1902];
assign g[3949] = b[10] & g[1902];
assign g[2927] = a[10] & g[1903];
assign g[3950] = b[10] & g[1903];
assign g[2928] = a[10] & g[1904];
assign g[3951] = b[10] & g[1904];
assign g[2929] = a[10] & g[1905];
assign g[3952] = b[10] & g[1905];
assign g[2930] = a[10] & g[1906];
assign g[3953] = b[10] & g[1906];
assign g[2931] = a[10] & g[1907];
assign g[3954] = b[10] & g[1907];
assign g[2932] = a[10] & g[1908];
assign g[3955] = b[10] & g[1908];
assign g[2933] = a[10] & g[1909];
assign g[3956] = b[10] & g[1909];
assign g[2934] = a[10] & g[1910];
assign g[3957] = b[10] & g[1910];
assign g[2935] = a[10] & g[1911];
assign g[3958] = b[10] & g[1911];
assign g[2936] = a[10] & g[1912];
assign g[3959] = b[10] & g[1912];
assign g[2937] = a[10] & g[1913];
assign g[3960] = b[10] & g[1913];
assign g[2938] = a[10] & g[1914];
assign g[3961] = b[10] & g[1914];
assign g[2939] = a[10] & g[1915];
assign g[3962] = b[10] & g[1915];
assign g[2940] = a[10] & g[1916];
assign g[3963] = b[10] & g[1916];
assign g[2941] = a[10] & g[1917];
assign g[3964] = b[10] & g[1917];
assign g[2942] = a[10] & g[1918];
assign g[3965] = b[10] & g[1918];
assign g[2943] = a[10] & g[1919];
assign g[3966] = b[10] & g[1919];
assign g[2944] = a[10] & g[1920];
assign g[3967] = b[10] & g[1920];
assign g[2945] = a[10] & g[1921];
assign g[3968] = b[10] & g[1921];
assign g[2946] = a[10] & g[1922];
assign g[3969] = b[10] & g[1922];
assign g[2947] = a[10] & g[1923];
assign g[3970] = b[10] & g[1923];
assign g[2948] = a[10] & g[1924];
assign g[3971] = b[10] & g[1924];
assign g[2949] = a[10] & g[1925];
assign g[3972] = b[10] & g[1925];
assign g[2950] = a[10] & g[1926];
assign g[3973] = b[10] & g[1926];
assign g[2951] = a[10] & g[1927];
assign g[3974] = b[10] & g[1927];
assign g[2952] = a[10] & g[1928];
assign g[3975] = b[10] & g[1928];
assign g[2953] = a[10] & g[1929];
assign g[3976] = b[10] & g[1929];
assign g[2954] = a[10] & g[1930];
assign g[3977] = b[10] & g[1930];
assign g[2955] = a[10] & g[1931];
assign g[3978] = b[10] & g[1931];
assign g[2956] = a[10] & g[1932];
assign g[3979] = b[10] & g[1932];
assign g[2957] = a[10] & g[1933];
assign g[3980] = b[10] & g[1933];
assign g[2958] = a[10] & g[1934];
assign g[3981] = b[10] & g[1934];
assign g[2959] = a[10] & g[1935];
assign g[3982] = b[10] & g[1935];
assign g[2960] = a[10] & g[1936];
assign g[3983] = b[10] & g[1936];
assign g[2961] = a[10] & g[1937];
assign g[3984] = b[10] & g[1937];
assign g[2962] = a[10] & g[1938];
assign g[3985] = b[10] & g[1938];
assign g[2963] = a[10] & g[1939];
assign g[3986] = b[10] & g[1939];
assign g[2964] = a[10] & g[1940];
assign g[3987] = b[10] & g[1940];
assign g[2965] = a[10] & g[1941];
assign g[3988] = b[10] & g[1941];
assign g[2966] = a[10] & g[1942];
assign g[3989] = b[10] & g[1942];
assign g[2967] = a[10] & g[1943];
assign g[3990] = b[10] & g[1943];
assign g[2968] = a[10] & g[1944];
assign g[3991] = b[10] & g[1944];
assign g[2969] = a[10] & g[1945];
assign g[3992] = b[10] & g[1945];
assign g[2970] = a[10] & g[1946];
assign g[3993] = b[10] & g[1946];
assign g[2971] = a[10] & g[1947];
assign g[3994] = b[10] & g[1947];
assign g[2972] = a[10] & g[1948];
assign g[3995] = b[10] & g[1948];
assign g[2973] = a[10] & g[1949];
assign g[3996] = b[10] & g[1949];
assign g[2974] = a[10] & g[1950];
assign g[3997] = b[10] & g[1950];
assign g[2975] = a[10] & g[1951];
assign g[3998] = b[10] & g[1951];
assign g[2976] = a[10] & g[1952];
assign g[3999] = b[10] & g[1952];
assign g[2977] = a[10] & g[1953];
assign g[4000] = b[10] & g[1953];
assign g[2978] = a[10] & g[1954];
assign g[4001] = b[10] & g[1954];
assign g[2979] = a[10] & g[1955];
assign g[4002] = b[10] & g[1955];
assign g[2980] = a[10] & g[1956];
assign g[4003] = b[10] & g[1956];
assign g[2981] = a[10] & g[1957];
assign g[4004] = b[10] & g[1957];
assign g[2982] = a[10] & g[1958];
assign g[4005] = b[10] & g[1958];
assign g[2983] = a[10] & g[1959];
assign g[4006] = b[10] & g[1959];
assign g[2984] = a[10] & g[1960];
assign g[4007] = b[10] & g[1960];
assign g[2985] = a[10] & g[1961];
assign g[4008] = b[10] & g[1961];
assign g[2986] = a[10] & g[1962];
assign g[4009] = b[10] & g[1962];
assign g[2987] = a[10] & g[1963];
assign g[4010] = b[10] & g[1963];
assign g[2988] = a[10] & g[1964];
assign g[4011] = b[10] & g[1964];
assign g[2989] = a[10] & g[1965];
assign g[4012] = b[10] & g[1965];
assign g[2990] = a[10] & g[1966];
assign g[4013] = b[10] & g[1966];
assign g[2991] = a[10] & g[1967];
assign g[4014] = b[10] & g[1967];
assign g[2992] = a[10] & g[1968];
assign g[4015] = b[10] & g[1968];
assign g[2993] = a[10] & g[1969];
assign g[4016] = b[10] & g[1969];
assign g[2994] = a[10] & g[1970];
assign g[4017] = b[10] & g[1970];
assign g[2995] = a[10] & g[1971];
assign g[4018] = b[10] & g[1971];
assign g[2996] = a[10] & g[1972];
assign g[4019] = b[10] & g[1972];
assign g[2997] = a[10] & g[1973];
assign g[4020] = b[10] & g[1973];
assign g[2998] = a[10] & g[1974];
assign g[4021] = b[10] & g[1974];
assign g[2999] = a[10] & g[1975];
assign g[4022] = b[10] & g[1975];
assign g[3000] = a[10] & g[1976];
assign g[4023] = b[10] & g[1976];
assign g[3001] = a[10] & g[1977];
assign g[4024] = b[10] & g[1977];
assign g[3002] = a[10] & g[1978];
assign g[4025] = b[10] & g[1978];
assign g[3003] = a[10] & g[1979];
assign g[4026] = b[10] & g[1979];
assign g[3004] = a[10] & g[1980];
assign g[4027] = b[10] & g[1980];
assign g[3005] = a[10] & g[1981];
assign g[4028] = b[10] & g[1981];
assign g[3006] = a[10] & g[1982];
assign g[4029] = b[10] & g[1982];
assign g[3007] = a[10] & g[1983];
assign g[4030] = b[10] & g[1983];
assign g[3008] = a[10] & g[1984];
assign g[4031] = b[10] & g[1984];
assign g[3009] = a[10] & g[1985];
assign g[4032] = b[10] & g[1985];
assign g[3010] = a[10] & g[1986];
assign g[4033] = b[10] & g[1986];
assign g[3011] = a[10] & g[1987];
assign g[4034] = b[10] & g[1987];
assign g[3012] = a[10] & g[1988];
assign g[4035] = b[10] & g[1988];
assign g[3013] = a[10] & g[1989];
assign g[4036] = b[10] & g[1989];
assign g[3014] = a[10] & g[1990];
assign g[4037] = b[10] & g[1990];
assign g[3015] = a[10] & g[1991];
assign g[4038] = b[10] & g[1991];
assign g[3016] = a[10] & g[1992];
assign g[4039] = b[10] & g[1992];
assign g[3017] = a[10] & g[1993];
assign g[4040] = b[10] & g[1993];
assign g[3018] = a[10] & g[1994];
assign g[4041] = b[10] & g[1994];
assign g[3019] = a[10] & g[1995];
assign g[4042] = b[10] & g[1995];
assign g[3020] = a[10] & g[1996];
assign g[4043] = b[10] & g[1996];
assign g[3021] = a[10] & g[1997];
assign g[4044] = b[10] & g[1997];
assign g[3022] = a[10] & g[1998];
assign g[4045] = b[10] & g[1998];
assign g[3023] = a[10] & g[1999];
assign g[4046] = b[10] & g[1999];
assign g[3024] = a[10] & g[2000];
assign g[4047] = b[10] & g[2000];
assign g[3025] = a[10] & g[2001];
assign g[4048] = b[10] & g[2001];
assign g[3026] = a[10] & g[2002];
assign g[4049] = b[10] & g[2002];
assign g[3027] = a[10] & g[2003];
assign g[4050] = b[10] & g[2003];
assign g[3028] = a[10] & g[2004];
assign g[4051] = b[10] & g[2004];
assign g[3029] = a[10] & g[2005];
assign g[4052] = b[10] & g[2005];
assign g[3030] = a[10] & g[2006];
assign g[4053] = b[10] & g[2006];
assign g[3031] = a[10] & g[2007];
assign g[4054] = b[10] & g[2007];
assign g[3032] = a[10] & g[2008];
assign g[4055] = b[10] & g[2008];
assign g[3033] = a[10] & g[2009];
assign g[4056] = b[10] & g[2009];
assign g[3034] = a[10] & g[2010];
assign g[4057] = b[10] & g[2010];
assign g[3035] = a[10] & g[2011];
assign g[4058] = b[10] & g[2011];
assign g[3036] = a[10] & g[2012];
assign g[4059] = b[10] & g[2012];
assign g[3037] = a[10] & g[2013];
assign g[4060] = b[10] & g[2013];
assign g[3038] = a[10] & g[2014];
assign g[4061] = b[10] & g[2014];
assign g[3039] = a[10] & g[2015];
assign g[4062] = b[10] & g[2015];
assign g[3040] = a[10] & g[2016];
assign g[4063] = b[10] & g[2016];
assign g[3041] = a[10] & g[2017];
assign g[4064] = b[10] & g[2017];
assign g[3042] = a[10] & g[2018];
assign g[4065] = b[10] & g[2018];
assign g[3043] = a[10] & g[2019];
assign g[4066] = b[10] & g[2019];
assign g[3044] = a[10] & g[2020];
assign g[4067] = b[10] & g[2020];
assign g[3045] = a[10] & g[2021];
assign g[4068] = b[10] & g[2021];
assign g[3046] = a[10] & g[2022];
assign g[4069] = b[10] & g[2022];
assign g[3047] = a[10] & g[2023];
assign g[4070] = b[10] & g[2023];
assign g[3048] = a[10] & g[2024];
assign g[4071] = b[10] & g[2024];
assign g[3049] = a[10] & g[2025];
assign g[4072] = b[10] & g[2025];
assign g[3050] = a[10] & g[2026];
assign g[4073] = b[10] & g[2026];
assign g[3051] = a[10] & g[2027];
assign g[4074] = b[10] & g[2027];
assign g[3052] = a[10] & g[2028];
assign g[4075] = b[10] & g[2028];
assign g[3053] = a[10] & g[2029];
assign g[4076] = b[10] & g[2029];
assign g[3054] = a[10] & g[2030];
assign g[4077] = b[10] & g[2030];
assign g[3055] = a[10] & g[2031];
assign g[4078] = b[10] & g[2031];
assign g[3056] = a[10] & g[2032];
assign g[4079] = b[10] & g[2032];
assign g[3057] = a[10] & g[2033];
assign g[4080] = b[10] & g[2033];
assign g[3058] = a[10] & g[2034];
assign g[4081] = b[10] & g[2034];
assign g[3059] = a[10] & g[2035];
assign g[4082] = b[10] & g[2035];
//Assigning outputs for input bit 12
assign g[4083] = a[11] & b[11];
assign g[4084] = a[11] & g[2036];
assign g[6131] = b[11] & g[2036];
assign g[4085] = a[11] & g[2037];
assign g[6132] = b[11] & g[2037];
assign g[4086] = a[11] & g[2038];
assign g[6133] = b[11] & g[2038];
assign g[4087] = a[11] & g[2039];
assign g[6134] = b[11] & g[2039];
assign g[4088] = a[11] & g[2040];
assign g[6135] = b[11] & g[2040];
assign g[4089] = a[11] & g[2041];
assign g[6136] = b[11] & g[2041];
assign g[4090] = a[11] & g[2042];
assign g[6137] = b[11] & g[2042];
assign g[4091] = a[11] & g[2043];
assign g[6138] = b[11] & g[2043];
assign g[4092] = a[11] & g[2044];
assign g[6139] = b[11] & g[2044];
assign g[4093] = a[11] & g[2045];
assign g[6140] = b[11] & g[2045];
assign g[4094] = a[11] & g[2046];
assign g[6141] = b[11] & g[2046];
assign g[4095] = a[11] & g[2047];
assign g[6142] = b[11] & g[2047];
assign g[4096] = a[11] & g[2048];
assign g[6143] = b[11] & g[2048];
assign g[4097] = a[11] & g[2049];
assign g[6144] = b[11] & g[2049];
assign g[4098] = a[11] & g[2050];
assign g[6145] = b[11] & g[2050];
assign g[4099] = a[11] & g[2051];
assign g[6146] = b[11] & g[2051];
assign g[4100] = a[11] & g[2052];
assign g[6147] = b[11] & g[2052];
assign g[4101] = a[11] & g[2053];
assign g[6148] = b[11] & g[2053];
assign g[4102] = a[11] & g[2054];
assign g[6149] = b[11] & g[2054];
assign g[4103] = a[11] & g[2055];
assign g[6150] = b[11] & g[2055];
assign g[4104] = a[11] & g[2056];
assign g[6151] = b[11] & g[2056];
assign g[4105] = a[11] & g[2057];
assign g[6152] = b[11] & g[2057];
assign g[4106] = a[11] & g[2058];
assign g[6153] = b[11] & g[2058];
assign g[4107] = a[11] & g[2059];
assign g[6154] = b[11] & g[2059];
assign g[4108] = a[11] & g[2060];
assign g[6155] = b[11] & g[2060];
assign g[4109] = a[11] & g[2061];
assign g[6156] = b[11] & g[2061];
assign g[4110] = a[11] & g[2062];
assign g[6157] = b[11] & g[2062];
assign g[4111] = a[11] & g[2063];
assign g[6158] = b[11] & g[2063];
assign g[4112] = a[11] & g[2064];
assign g[6159] = b[11] & g[2064];
assign g[4113] = a[11] & g[2065];
assign g[6160] = b[11] & g[2065];
assign g[4114] = a[11] & g[2066];
assign g[6161] = b[11] & g[2066];
assign g[4115] = a[11] & g[2067];
assign g[6162] = b[11] & g[2067];
assign g[4116] = a[11] & g[2068];
assign g[6163] = b[11] & g[2068];
assign g[4117] = a[11] & g[2069];
assign g[6164] = b[11] & g[2069];
assign g[4118] = a[11] & g[2070];
assign g[6165] = b[11] & g[2070];
assign g[4119] = a[11] & g[2071];
assign g[6166] = b[11] & g[2071];
assign g[4120] = a[11] & g[2072];
assign g[6167] = b[11] & g[2072];
assign g[4121] = a[11] & g[2073];
assign g[6168] = b[11] & g[2073];
assign g[4122] = a[11] & g[2074];
assign g[6169] = b[11] & g[2074];
assign g[4123] = a[11] & g[2075];
assign g[6170] = b[11] & g[2075];
assign g[4124] = a[11] & g[2076];
assign g[6171] = b[11] & g[2076];
assign g[4125] = a[11] & g[2077];
assign g[6172] = b[11] & g[2077];
assign g[4126] = a[11] & g[2078];
assign g[6173] = b[11] & g[2078];
assign g[4127] = a[11] & g[2079];
assign g[6174] = b[11] & g[2079];
assign g[4128] = a[11] & g[2080];
assign g[6175] = b[11] & g[2080];
assign g[4129] = a[11] & g[2081];
assign g[6176] = b[11] & g[2081];
assign g[4130] = a[11] & g[2082];
assign g[6177] = b[11] & g[2082];
assign g[4131] = a[11] & g[2083];
assign g[6178] = b[11] & g[2083];
assign g[4132] = a[11] & g[2084];
assign g[6179] = b[11] & g[2084];
assign g[4133] = a[11] & g[2085];
assign g[6180] = b[11] & g[2085];
assign g[4134] = a[11] & g[2086];
assign g[6181] = b[11] & g[2086];
assign g[4135] = a[11] & g[2087];
assign g[6182] = b[11] & g[2087];
assign g[4136] = a[11] & g[2088];
assign g[6183] = b[11] & g[2088];
assign g[4137] = a[11] & g[2089];
assign g[6184] = b[11] & g[2089];
assign g[4138] = a[11] & g[2090];
assign g[6185] = b[11] & g[2090];
assign g[4139] = a[11] & g[2091];
assign g[6186] = b[11] & g[2091];
assign g[4140] = a[11] & g[2092];
assign g[6187] = b[11] & g[2092];
assign g[4141] = a[11] & g[2093];
assign g[6188] = b[11] & g[2093];
assign g[4142] = a[11] & g[2094];
assign g[6189] = b[11] & g[2094];
assign g[4143] = a[11] & g[2095];
assign g[6190] = b[11] & g[2095];
assign g[4144] = a[11] & g[2096];
assign g[6191] = b[11] & g[2096];
assign g[4145] = a[11] & g[2097];
assign g[6192] = b[11] & g[2097];
assign g[4146] = a[11] & g[2098];
assign g[6193] = b[11] & g[2098];
assign g[4147] = a[11] & g[2099];
assign g[6194] = b[11] & g[2099];
assign g[4148] = a[11] & g[2100];
assign g[6195] = b[11] & g[2100];
assign g[4149] = a[11] & g[2101];
assign g[6196] = b[11] & g[2101];
assign g[4150] = a[11] & g[2102];
assign g[6197] = b[11] & g[2102];
assign g[4151] = a[11] & g[2103];
assign g[6198] = b[11] & g[2103];
assign g[4152] = a[11] & g[2104];
assign g[6199] = b[11] & g[2104];
assign g[4153] = a[11] & g[2105];
assign g[6200] = b[11] & g[2105];
assign g[4154] = a[11] & g[2106];
assign g[6201] = b[11] & g[2106];
assign g[4155] = a[11] & g[2107];
assign g[6202] = b[11] & g[2107];
assign g[4156] = a[11] & g[2108];
assign g[6203] = b[11] & g[2108];
assign g[4157] = a[11] & g[2109];
assign g[6204] = b[11] & g[2109];
assign g[4158] = a[11] & g[2110];
assign g[6205] = b[11] & g[2110];
assign g[4159] = a[11] & g[2111];
assign g[6206] = b[11] & g[2111];
assign g[4160] = a[11] & g[2112];
assign g[6207] = b[11] & g[2112];
assign g[4161] = a[11] & g[2113];
assign g[6208] = b[11] & g[2113];
assign g[4162] = a[11] & g[2114];
assign g[6209] = b[11] & g[2114];
assign g[4163] = a[11] & g[2115];
assign g[6210] = b[11] & g[2115];
assign g[4164] = a[11] & g[2116];
assign g[6211] = b[11] & g[2116];
assign g[4165] = a[11] & g[2117];
assign g[6212] = b[11] & g[2117];
assign g[4166] = a[11] & g[2118];
assign g[6213] = b[11] & g[2118];
assign g[4167] = a[11] & g[2119];
assign g[6214] = b[11] & g[2119];
assign g[4168] = a[11] & g[2120];
assign g[6215] = b[11] & g[2120];
assign g[4169] = a[11] & g[2121];
assign g[6216] = b[11] & g[2121];
assign g[4170] = a[11] & g[2122];
assign g[6217] = b[11] & g[2122];
assign g[4171] = a[11] & g[2123];
assign g[6218] = b[11] & g[2123];
assign g[4172] = a[11] & g[2124];
assign g[6219] = b[11] & g[2124];
assign g[4173] = a[11] & g[2125];
assign g[6220] = b[11] & g[2125];
assign g[4174] = a[11] & g[2126];
assign g[6221] = b[11] & g[2126];
assign g[4175] = a[11] & g[2127];
assign g[6222] = b[11] & g[2127];
assign g[4176] = a[11] & g[2128];
assign g[6223] = b[11] & g[2128];
assign g[4177] = a[11] & g[2129];
assign g[6224] = b[11] & g[2129];
assign g[4178] = a[11] & g[2130];
assign g[6225] = b[11] & g[2130];
assign g[4179] = a[11] & g[2131];
assign g[6226] = b[11] & g[2131];
assign g[4180] = a[11] & g[2132];
assign g[6227] = b[11] & g[2132];
assign g[4181] = a[11] & g[2133];
assign g[6228] = b[11] & g[2133];
assign g[4182] = a[11] & g[2134];
assign g[6229] = b[11] & g[2134];
assign g[4183] = a[11] & g[2135];
assign g[6230] = b[11] & g[2135];
assign g[4184] = a[11] & g[2136];
assign g[6231] = b[11] & g[2136];
assign g[4185] = a[11] & g[2137];
assign g[6232] = b[11] & g[2137];
assign g[4186] = a[11] & g[2138];
assign g[6233] = b[11] & g[2138];
assign g[4187] = a[11] & g[2139];
assign g[6234] = b[11] & g[2139];
assign g[4188] = a[11] & g[2140];
assign g[6235] = b[11] & g[2140];
assign g[4189] = a[11] & g[2141];
assign g[6236] = b[11] & g[2141];
assign g[4190] = a[11] & g[2142];
assign g[6237] = b[11] & g[2142];
assign g[4191] = a[11] & g[2143];
assign g[6238] = b[11] & g[2143];
assign g[4192] = a[11] & g[2144];
assign g[6239] = b[11] & g[2144];
assign g[4193] = a[11] & g[2145];
assign g[6240] = b[11] & g[2145];
assign g[4194] = a[11] & g[2146];
assign g[6241] = b[11] & g[2146];
assign g[4195] = a[11] & g[2147];
assign g[6242] = b[11] & g[2147];
assign g[4196] = a[11] & g[2148];
assign g[6243] = b[11] & g[2148];
assign g[4197] = a[11] & g[2149];
assign g[6244] = b[11] & g[2149];
assign g[4198] = a[11] & g[2150];
assign g[6245] = b[11] & g[2150];
assign g[4199] = a[11] & g[2151];
assign g[6246] = b[11] & g[2151];
assign g[4200] = a[11] & g[2152];
assign g[6247] = b[11] & g[2152];
assign g[4201] = a[11] & g[2153];
assign g[6248] = b[11] & g[2153];
assign g[4202] = a[11] & g[2154];
assign g[6249] = b[11] & g[2154];
assign g[4203] = a[11] & g[2155];
assign g[6250] = b[11] & g[2155];
assign g[4204] = a[11] & g[2156];
assign g[6251] = b[11] & g[2156];
assign g[4205] = a[11] & g[2157];
assign g[6252] = b[11] & g[2157];
assign g[4206] = a[11] & g[2158];
assign g[6253] = b[11] & g[2158];
assign g[4207] = a[11] & g[2159];
assign g[6254] = b[11] & g[2159];
assign g[4208] = a[11] & g[2160];
assign g[6255] = b[11] & g[2160];
assign g[4209] = a[11] & g[2161];
assign g[6256] = b[11] & g[2161];
assign g[4210] = a[11] & g[2162];
assign g[6257] = b[11] & g[2162];
assign g[4211] = a[11] & g[2163];
assign g[6258] = b[11] & g[2163];
assign g[4212] = a[11] & g[2164];
assign g[6259] = b[11] & g[2164];
assign g[4213] = a[11] & g[2165];
assign g[6260] = b[11] & g[2165];
assign g[4214] = a[11] & g[2166];
assign g[6261] = b[11] & g[2166];
assign g[4215] = a[11] & g[2167];
assign g[6262] = b[11] & g[2167];
assign g[4216] = a[11] & g[2168];
assign g[6263] = b[11] & g[2168];
assign g[4217] = a[11] & g[2169];
assign g[6264] = b[11] & g[2169];
assign g[4218] = a[11] & g[2170];
assign g[6265] = b[11] & g[2170];
assign g[4219] = a[11] & g[2171];
assign g[6266] = b[11] & g[2171];
assign g[4220] = a[11] & g[2172];
assign g[6267] = b[11] & g[2172];
assign g[4221] = a[11] & g[2173];
assign g[6268] = b[11] & g[2173];
assign g[4222] = a[11] & g[2174];
assign g[6269] = b[11] & g[2174];
assign g[4223] = a[11] & g[2175];
assign g[6270] = b[11] & g[2175];
assign g[4224] = a[11] & g[2176];
assign g[6271] = b[11] & g[2176];
assign g[4225] = a[11] & g[2177];
assign g[6272] = b[11] & g[2177];
assign g[4226] = a[11] & g[2178];
assign g[6273] = b[11] & g[2178];
assign g[4227] = a[11] & g[2179];
assign g[6274] = b[11] & g[2179];
assign g[4228] = a[11] & g[2180];
assign g[6275] = b[11] & g[2180];
assign g[4229] = a[11] & g[2181];
assign g[6276] = b[11] & g[2181];
assign g[4230] = a[11] & g[2182];
assign g[6277] = b[11] & g[2182];
assign g[4231] = a[11] & g[2183];
assign g[6278] = b[11] & g[2183];
assign g[4232] = a[11] & g[2184];
assign g[6279] = b[11] & g[2184];
assign g[4233] = a[11] & g[2185];
assign g[6280] = b[11] & g[2185];
assign g[4234] = a[11] & g[2186];
assign g[6281] = b[11] & g[2186];
assign g[4235] = a[11] & g[2187];
assign g[6282] = b[11] & g[2187];
assign g[4236] = a[11] & g[2188];
assign g[6283] = b[11] & g[2188];
assign g[4237] = a[11] & g[2189];
assign g[6284] = b[11] & g[2189];
assign g[4238] = a[11] & g[2190];
assign g[6285] = b[11] & g[2190];
assign g[4239] = a[11] & g[2191];
assign g[6286] = b[11] & g[2191];
assign g[4240] = a[11] & g[2192];
assign g[6287] = b[11] & g[2192];
assign g[4241] = a[11] & g[2193];
assign g[6288] = b[11] & g[2193];
assign g[4242] = a[11] & g[2194];
assign g[6289] = b[11] & g[2194];
assign g[4243] = a[11] & g[2195];
assign g[6290] = b[11] & g[2195];
assign g[4244] = a[11] & g[2196];
assign g[6291] = b[11] & g[2196];
assign g[4245] = a[11] & g[2197];
assign g[6292] = b[11] & g[2197];
assign g[4246] = a[11] & g[2198];
assign g[6293] = b[11] & g[2198];
assign g[4247] = a[11] & g[2199];
assign g[6294] = b[11] & g[2199];
assign g[4248] = a[11] & g[2200];
assign g[6295] = b[11] & g[2200];
assign g[4249] = a[11] & g[2201];
assign g[6296] = b[11] & g[2201];
assign g[4250] = a[11] & g[2202];
assign g[6297] = b[11] & g[2202];
assign g[4251] = a[11] & g[2203];
assign g[6298] = b[11] & g[2203];
assign g[4252] = a[11] & g[2204];
assign g[6299] = b[11] & g[2204];
assign g[4253] = a[11] & g[2205];
assign g[6300] = b[11] & g[2205];
assign g[4254] = a[11] & g[2206];
assign g[6301] = b[11] & g[2206];
assign g[4255] = a[11] & g[2207];
assign g[6302] = b[11] & g[2207];
assign g[4256] = a[11] & g[2208];
assign g[6303] = b[11] & g[2208];
assign g[4257] = a[11] & g[2209];
assign g[6304] = b[11] & g[2209];
assign g[4258] = a[11] & g[2210];
assign g[6305] = b[11] & g[2210];
assign g[4259] = a[11] & g[2211];
assign g[6306] = b[11] & g[2211];
assign g[4260] = a[11] & g[2212];
assign g[6307] = b[11] & g[2212];
assign g[4261] = a[11] & g[2213];
assign g[6308] = b[11] & g[2213];
assign g[4262] = a[11] & g[2214];
assign g[6309] = b[11] & g[2214];
assign g[4263] = a[11] & g[2215];
assign g[6310] = b[11] & g[2215];
assign g[4264] = a[11] & g[2216];
assign g[6311] = b[11] & g[2216];
assign g[4265] = a[11] & g[2217];
assign g[6312] = b[11] & g[2217];
assign g[4266] = a[11] & g[2218];
assign g[6313] = b[11] & g[2218];
assign g[4267] = a[11] & g[2219];
assign g[6314] = b[11] & g[2219];
assign g[4268] = a[11] & g[2220];
assign g[6315] = b[11] & g[2220];
assign g[4269] = a[11] & g[2221];
assign g[6316] = b[11] & g[2221];
assign g[4270] = a[11] & g[2222];
assign g[6317] = b[11] & g[2222];
assign g[4271] = a[11] & g[2223];
assign g[6318] = b[11] & g[2223];
assign g[4272] = a[11] & g[2224];
assign g[6319] = b[11] & g[2224];
assign g[4273] = a[11] & g[2225];
assign g[6320] = b[11] & g[2225];
assign g[4274] = a[11] & g[2226];
assign g[6321] = b[11] & g[2226];
assign g[4275] = a[11] & g[2227];
assign g[6322] = b[11] & g[2227];
assign g[4276] = a[11] & g[2228];
assign g[6323] = b[11] & g[2228];
assign g[4277] = a[11] & g[2229];
assign g[6324] = b[11] & g[2229];
assign g[4278] = a[11] & g[2230];
assign g[6325] = b[11] & g[2230];
assign g[4279] = a[11] & g[2231];
assign g[6326] = b[11] & g[2231];
assign g[4280] = a[11] & g[2232];
assign g[6327] = b[11] & g[2232];
assign g[4281] = a[11] & g[2233];
assign g[6328] = b[11] & g[2233];
assign g[4282] = a[11] & g[2234];
assign g[6329] = b[11] & g[2234];
assign g[4283] = a[11] & g[2235];
assign g[6330] = b[11] & g[2235];
assign g[4284] = a[11] & g[2236];
assign g[6331] = b[11] & g[2236];
assign g[4285] = a[11] & g[2237];
assign g[6332] = b[11] & g[2237];
assign g[4286] = a[11] & g[2238];
assign g[6333] = b[11] & g[2238];
assign g[4287] = a[11] & g[2239];
assign g[6334] = b[11] & g[2239];
assign g[4288] = a[11] & g[2240];
assign g[6335] = b[11] & g[2240];
assign g[4289] = a[11] & g[2241];
assign g[6336] = b[11] & g[2241];
assign g[4290] = a[11] & g[2242];
assign g[6337] = b[11] & g[2242];
assign g[4291] = a[11] & g[2243];
assign g[6338] = b[11] & g[2243];
assign g[4292] = a[11] & g[2244];
assign g[6339] = b[11] & g[2244];
assign g[4293] = a[11] & g[2245];
assign g[6340] = b[11] & g[2245];
assign g[4294] = a[11] & g[2246];
assign g[6341] = b[11] & g[2246];
assign g[4295] = a[11] & g[2247];
assign g[6342] = b[11] & g[2247];
assign g[4296] = a[11] & g[2248];
assign g[6343] = b[11] & g[2248];
assign g[4297] = a[11] & g[2249];
assign g[6344] = b[11] & g[2249];
assign g[4298] = a[11] & g[2250];
assign g[6345] = b[11] & g[2250];
assign g[4299] = a[11] & g[2251];
assign g[6346] = b[11] & g[2251];
assign g[4300] = a[11] & g[2252];
assign g[6347] = b[11] & g[2252];
assign g[4301] = a[11] & g[2253];
assign g[6348] = b[11] & g[2253];
assign g[4302] = a[11] & g[2254];
assign g[6349] = b[11] & g[2254];
assign g[4303] = a[11] & g[2255];
assign g[6350] = b[11] & g[2255];
assign g[4304] = a[11] & g[2256];
assign g[6351] = b[11] & g[2256];
assign g[4305] = a[11] & g[2257];
assign g[6352] = b[11] & g[2257];
assign g[4306] = a[11] & g[2258];
assign g[6353] = b[11] & g[2258];
assign g[4307] = a[11] & g[2259];
assign g[6354] = b[11] & g[2259];
assign g[4308] = a[11] & g[2260];
assign g[6355] = b[11] & g[2260];
assign g[4309] = a[11] & g[2261];
assign g[6356] = b[11] & g[2261];
assign g[4310] = a[11] & g[2262];
assign g[6357] = b[11] & g[2262];
assign g[4311] = a[11] & g[2263];
assign g[6358] = b[11] & g[2263];
assign g[4312] = a[11] & g[2264];
assign g[6359] = b[11] & g[2264];
assign g[4313] = a[11] & g[2265];
assign g[6360] = b[11] & g[2265];
assign g[4314] = a[11] & g[2266];
assign g[6361] = b[11] & g[2266];
assign g[4315] = a[11] & g[2267];
assign g[6362] = b[11] & g[2267];
assign g[4316] = a[11] & g[2268];
assign g[6363] = b[11] & g[2268];
assign g[4317] = a[11] & g[2269];
assign g[6364] = b[11] & g[2269];
assign g[4318] = a[11] & g[2270];
assign g[6365] = b[11] & g[2270];
assign g[4319] = a[11] & g[2271];
assign g[6366] = b[11] & g[2271];
assign g[4320] = a[11] & g[2272];
assign g[6367] = b[11] & g[2272];
assign g[4321] = a[11] & g[2273];
assign g[6368] = b[11] & g[2273];
assign g[4322] = a[11] & g[2274];
assign g[6369] = b[11] & g[2274];
assign g[4323] = a[11] & g[2275];
assign g[6370] = b[11] & g[2275];
assign g[4324] = a[11] & g[2276];
assign g[6371] = b[11] & g[2276];
assign g[4325] = a[11] & g[2277];
assign g[6372] = b[11] & g[2277];
assign g[4326] = a[11] & g[2278];
assign g[6373] = b[11] & g[2278];
assign g[4327] = a[11] & g[2279];
assign g[6374] = b[11] & g[2279];
assign g[4328] = a[11] & g[2280];
assign g[6375] = b[11] & g[2280];
assign g[4329] = a[11] & g[2281];
assign g[6376] = b[11] & g[2281];
assign g[4330] = a[11] & g[2282];
assign g[6377] = b[11] & g[2282];
assign g[4331] = a[11] & g[2283];
assign g[6378] = b[11] & g[2283];
assign g[4332] = a[11] & g[2284];
assign g[6379] = b[11] & g[2284];
assign g[4333] = a[11] & g[2285];
assign g[6380] = b[11] & g[2285];
assign g[4334] = a[11] & g[2286];
assign g[6381] = b[11] & g[2286];
assign g[4335] = a[11] & g[2287];
assign g[6382] = b[11] & g[2287];
assign g[4336] = a[11] & g[2288];
assign g[6383] = b[11] & g[2288];
assign g[4337] = a[11] & g[2289];
assign g[6384] = b[11] & g[2289];
assign g[4338] = a[11] & g[2290];
assign g[6385] = b[11] & g[2290];
assign g[4339] = a[11] & g[2291];
assign g[6386] = b[11] & g[2291];
assign g[4340] = a[11] & g[2292];
assign g[6387] = b[11] & g[2292];
assign g[4341] = a[11] & g[2293];
assign g[6388] = b[11] & g[2293];
assign g[4342] = a[11] & g[2294];
assign g[6389] = b[11] & g[2294];
assign g[4343] = a[11] & g[2295];
assign g[6390] = b[11] & g[2295];
assign g[4344] = a[11] & g[2296];
assign g[6391] = b[11] & g[2296];
assign g[4345] = a[11] & g[2297];
assign g[6392] = b[11] & g[2297];
assign g[4346] = a[11] & g[2298];
assign g[6393] = b[11] & g[2298];
assign g[4347] = a[11] & g[2299];
assign g[6394] = b[11] & g[2299];
assign g[4348] = a[11] & g[2300];
assign g[6395] = b[11] & g[2300];
assign g[4349] = a[11] & g[2301];
assign g[6396] = b[11] & g[2301];
assign g[4350] = a[11] & g[2302];
assign g[6397] = b[11] & g[2302];
assign g[4351] = a[11] & g[2303];
assign g[6398] = b[11] & g[2303];
assign g[4352] = a[11] & g[2304];
assign g[6399] = b[11] & g[2304];
assign g[4353] = a[11] & g[2305];
assign g[6400] = b[11] & g[2305];
assign g[4354] = a[11] & g[2306];
assign g[6401] = b[11] & g[2306];
assign g[4355] = a[11] & g[2307];
assign g[6402] = b[11] & g[2307];
assign g[4356] = a[11] & g[2308];
assign g[6403] = b[11] & g[2308];
assign g[4357] = a[11] & g[2309];
assign g[6404] = b[11] & g[2309];
assign g[4358] = a[11] & g[2310];
assign g[6405] = b[11] & g[2310];
assign g[4359] = a[11] & g[2311];
assign g[6406] = b[11] & g[2311];
assign g[4360] = a[11] & g[2312];
assign g[6407] = b[11] & g[2312];
assign g[4361] = a[11] & g[2313];
assign g[6408] = b[11] & g[2313];
assign g[4362] = a[11] & g[2314];
assign g[6409] = b[11] & g[2314];
assign g[4363] = a[11] & g[2315];
assign g[6410] = b[11] & g[2315];
assign g[4364] = a[11] & g[2316];
assign g[6411] = b[11] & g[2316];
assign g[4365] = a[11] & g[2317];
assign g[6412] = b[11] & g[2317];
assign g[4366] = a[11] & g[2318];
assign g[6413] = b[11] & g[2318];
assign g[4367] = a[11] & g[2319];
assign g[6414] = b[11] & g[2319];
assign g[4368] = a[11] & g[2320];
assign g[6415] = b[11] & g[2320];
assign g[4369] = a[11] & g[2321];
assign g[6416] = b[11] & g[2321];
assign g[4370] = a[11] & g[2322];
assign g[6417] = b[11] & g[2322];
assign g[4371] = a[11] & g[2323];
assign g[6418] = b[11] & g[2323];
assign g[4372] = a[11] & g[2324];
assign g[6419] = b[11] & g[2324];
assign g[4373] = a[11] & g[2325];
assign g[6420] = b[11] & g[2325];
assign g[4374] = a[11] & g[2326];
assign g[6421] = b[11] & g[2326];
assign g[4375] = a[11] & g[2327];
assign g[6422] = b[11] & g[2327];
assign g[4376] = a[11] & g[2328];
assign g[6423] = b[11] & g[2328];
assign g[4377] = a[11] & g[2329];
assign g[6424] = b[11] & g[2329];
assign g[4378] = a[11] & g[2330];
assign g[6425] = b[11] & g[2330];
assign g[4379] = a[11] & g[2331];
assign g[6426] = b[11] & g[2331];
assign g[4380] = a[11] & g[2332];
assign g[6427] = b[11] & g[2332];
assign g[4381] = a[11] & g[2333];
assign g[6428] = b[11] & g[2333];
assign g[4382] = a[11] & g[2334];
assign g[6429] = b[11] & g[2334];
assign g[4383] = a[11] & g[2335];
assign g[6430] = b[11] & g[2335];
assign g[4384] = a[11] & g[2336];
assign g[6431] = b[11] & g[2336];
assign g[4385] = a[11] & g[2337];
assign g[6432] = b[11] & g[2337];
assign g[4386] = a[11] & g[2338];
assign g[6433] = b[11] & g[2338];
assign g[4387] = a[11] & g[2339];
assign g[6434] = b[11] & g[2339];
assign g[4388] = a[11] & g[2340];
assign g[6435] = b[11] & g[2340];
assign g[4389] = a[11] & g[2341];
assign g[6436] = b[11] & g[2341];
assign g[4390] = a[11] & g[2342];
assign g[6437] = b[11] & g[2342];
assign g[4391] = a[11] & g[2343];
assign g[6438] = b[11] & g[2343];
assign g[4392] = a[11] & g[2344];
assign g[6439] = b[11] & g[2344];
assign g[4393] = a[11] & g[2345];
assign g[6440] = b[11] & g[2345];
assign g[4394] = a[11] & g[2346];
assign g[6441] = b[11] & g[2346];
assign g[4395] = a[11] & g[2347];
assign g[6442] = b[11] & g[2347];
assign g[4396] = a[11] & g[2348];
assign g[6443] = b[11] & g[2348];
assign g[4397] = a[11] & g[2349];
assign g[6444] = b[11] & g[2349];
assign g[4398] = a[11] & g[2350];
assign g[6445] = b[11] & g[2350];
assign g[4399] = a[11] & g[2351];
assign g[6446] = b[11] & g[2351];
assign g[4400] = a[11] & g[2352];
assign g[6447] = b[11] & g[2352];
assign g[4401] = a[11] & g[2353];
assign g[6448] = b[11] & g[2353];
assign g[4402] = a[11] & g[2354];
assign g[6449] = b[11] & g[2354];
assign g[4403] = a[11] & g[2355];
assign g[6450] = b[11] & g[2355];
assign g[4404] = a[11] & g[2356];
assign g[6451] = b[11] & g[2356];
assign g[4405] = a[11] & g[2357];
assign g[6452] = b[11] & g[2357];
assign g[4406] = a[11] & g[2358];
assign g[6453] = b[11] & g[2358];
assign g[4407] = a[11] & g[2359];
assign g[6454] = b[11] & g[2359];
assign g[4408] = a[11] & g[2360];
assign g[6455] = b[11] & g[2360];
assign g[4409] = a[11] & g[2361];
assign g[6456] = b[11] & g[2361];
assign g[4410] = a[11] & g[2362];
assign g[6457] = b[11] & g[2362];
assign g[4411] = a[11] & g[2363];
assign g[6458] = b[11] & g[2363];
assign g[4412] = a[11] & g[2364];
assign g[6459] = b[11] & g[2364];
assign g[4413] = a[11] & g[2365];
assign g[6460] = b[11] & g[2365];
assign g[4414] = a[11] & g[2366];
assign g[6461] = b[11] & g[2366];
assign g[4415] = a[11] & g[2367];
assign g[6462] = b[11] & g[2367];
assign g[4416] = a[11] & g[2368];
assign g[6463] = b[11] & g[2368];
assign g[4417] = a[11] & g[2369];
assign g[6464] = b[11] & g[2369];
assign g[4418] = a[11] & g[2370];
assign g[6465] = b[11] & g[2370];
assign g[4419] = a[11] & g[2371];
assign g[6466] = b[11] & g[2371];
assign g[4420] = a[11] & g[2372];
assign g[6467] = b[11] & g[2372];
assign g[4421] = a[11] & g[2373];
assign g[6468] = b[11] & g[2373];
assign g[4422] = a[11] & g[2374];
assign g[6469] = b[11] & g[2374];
assign g[4423] = a[11] & g[2375];
assign g[6470] = b[11] & g[2375];
assign g[4424] = a[11] & g[2376];
assign g[6471] = b[11] & g[2376];
assign g[4425] = a[11] & g[2377];
assign g[6472] = b[11] & g[2377];
assign g[4426] = a[11] & g[2378];
assign g[6473] = b[11] & g[2378];
assign g[4427] = a[11] & g[2379];
assign g[6474] = b[11] & g[2379];
assign g[4428] = a[11] & g[2380];
assign g[6475] = b[11] & g[2380];
assign g[4429] = a[11] & g[2381];
assign g[6476] = b[11] & g[2381];
assign g[4430] = a[11] & g[2382];
assign g[6477] = b[11] & g[2382];
assign g[4431] = a[11] & g[2383];
assign g[6478] = b[11] & g[2383];
assign g[4432] = a[11] & g[2384];
assign g[6479] = b[11] & g[2384];
assign g[4433] = a[11] & g[2385];
assign g[6480] = b[11] & g[2385];
assign g[4434] = a[11] & g[2386];
assign g[6481] = b[11] & g[2386];
assign g[4435] = a[11] & g[2387];
assign g[6482] = b[11] & g[2387];
assign g[4436] = a[11] & g[2388];
assign g[6483] = b[11] & g[2388];
assign g[4437] = a[11] & g[2389];
assign g[6484] = b[11] & g[2389];
assign g[4438] = a[11] & g[2390];
assign g[6485] = b[11] & g[2390];
assign g[4439] = a[11] & g[2391];
assign g[6486] = b[11] & g[2391];
assign g[4440] = a[11] & g[2392];
assign g[6487] = b[11] & g[2392];
assign g[4441] = a[11] & g[2393];
assign g[6488] = b[11] & g[2393];
assign g[4442] = a[11] & g[2394];
assign g[6489] = b[11] & g[2394];
assign g[4443] = a[11] & g[2395];
assign g[6490] = b[11] & g[2395];
assign g[4444] = a[11] & g[2396];
assign g[6491] = b[11] & g[2396];
assign g[4445] = a[11] & g[2397];
assign g[6492] = b[11] & g[2397];
assign g[4446] = a[11] & g[2398];
assign g[6493] = b[11] & g[2398];
assign g[4447] = a[11] & g[2399];
assign g[6494] = b[11] & g[2399];
assign g[4448] = a[11] & g[2400];
assign g[6495] = b[11] & g[2400];
assign g[4449] = a[11] & g[2401];
assign g[6496] = b[11] & g[2401];
assign g[4450] = a[11] & g[2402];
assign g[6497] = b[11] & g[2402];
assign g[4451] = a[11] & g[2403];
assign g[6498] = b[11] & g[2403];
assign g[4452] = a[11] & g[2404];
assign g[6499] = b[11] & g[2404];
assign g[4453] = a[11] & g[2405];
assign g[6500] = b[11] & g[2405];
assign g[4454] = a[11] & g[2406];
assign g[6501] = b[11] & g[2406];
assign g[4455] = a[11] & g[2407];
assign g[6502] = b[11] & g[2407];
assign g[4456] = a[11] & g[2408];
assign g[6503] = b[11] & g[2408];
assign g[4457] = a[11] & g[2409];
assign g[6504] = b[11] & g[2409];
assign g[4458] = a[11] & g[2410];
assign g[6505] = b[11] & g[2410];
assign g[4459] = a[11] & g[2411];
assign g[6506] = b[11] & g[2411];
assign g[4460] = a[11] & g[2412];
assign g[6507] = b[11] & g[2412];
assign g[4461] = a[11] & g[2413];
assign g[6508] = b[11] & g[2413];
assign g[4462] = a[11] & g[2414];
assign g[6509] = b[11] & g[2414];
assign g[4463] = a[11] & g[2415];
assign g[6510] = b[11] & g[2415];
assign g[4464] = a[11] & g[2416];
assign g[6511] = b[11] & g[2416];
assign g[4465] = a[11] & g[2417];
assign g[6512] = b[11] & g[2417];
assign g[4466] = a[11] & g[2418];
assign g[6513] = b[11] & g[2418];
assign g[4467] = a[11] & g[2419];
assign g[6514] = b[11] & g[2419];
assign g[4468] = a[11] & g[2420];
assign g[6515] = b[11] & g[2420];
assign g[4469] = a[11] & g[2421];
assign g[6516] = b[11] & g[2421];
assign g[4470] = a[11] & g[2422];
assign g[6517] = b[11] & g[2422];
assign g[4471] = a[11] & g[2423];
assign g[6518] = b[11] & g[2423];
assign g[4472] = a[11] & g[2424];
assign g[6519] = b[11] & g[2424];
assign g[4473] = a[11] & g[2425];
assign g[6520] = b[11] & g[2425];
assign g[4474] = a[11] & g[2426];
assign g[6521] = b[11] & g[2426];
assign g[4475] = a[11] & g[2427];
assign g[6522] = b[11] & g[2427];
assign g[4476] = a[11] & g[2428];
assign g[6523] = b[11] & g[2428];
assign g[4477] = a[11] & g[2429];
assign g[6524] = b[11] & g[2429];
assign g[4478] = a[11] & g[2430];
assign g[6525] = b[11] & g[2430];
assign g[4479] = a[11] & g[2431];
assign g[6526] = b[11] & g[2431];
assign g[4480] = a[11] & g[2432];
assign g[6527] = b[11] & g[2432];
assign g[4481] = a[11] & g[2433];
assign g[6528] = b[11] & g[2433];
assign g[4482] = a[11] & g[2434];
assign g[6529] = b[11] & g[2434];
assign g[4483] = a[11] & g[2435];
assign g[6530] = b[11] & g[2435];
assign g[4484] = a[11] & g[2436];
assign g[6531] = b[11] & g[2436];
assign g[4485] = a[11] & g[2437];
assign g[6532] = b[11] & g[2437];
assign g[4486] = a[11] & g[2438];
assign g[6533] = b[11] & g[2438];
assign g[4487] = a[11] & g[2439];
assign g[6534] = b[11] & g[2439];
assign g[4488] = a[11] & g[2440];
assign g[6535] = b[11] & g[2440];
assign g[4489] = a[11] & g[2441];
assign g[6536] = b[11] & g[2441];
assign g[4490] = a[11] & g[2442];
assign g[6537] = b[11] & g[2442];
assign g[4491] = a[11] & g[2443];
assign g[6538] = b[11] & g[2443];
assign g[4492] = a[11] & g[2444];
assign g[6539] = b[11] & g[2444];
assign g[4493] = a[11] & g[2445];
assign g[6540] = b[11] & g[2445];
assign g[4494] = a[11] & g[2446];
assign g[6541] = b[11] & g[2446];
assign g[4495] = a[11] & g[2447];
assign g[6542] = b[11] & g[2447];
assign g[4496] = a[11] & g[2448];
assign g[6543] = b[11] & g[2448];
assign g[4497] = a[11] & g[2449];
assign g[6544] = b[11] & g[2449];
assign g[4498] = a[11] & g[2450];
assign g[6545] = b[11] & g[2450];
assign g[4499] = a[11] & g[2451];
assign g[6546] = b[11] & g[2451];
assign g[4500] = a[11] & g[2452];
assign g[6547] = b[11] & g[2452];
assign g[4501] = a[11] & g[2453];
assign g[6548] = b[11] & g[2453];
assign g[4502] = a[11] & g[2454];
assign g[6549] = b[11] & g[2454];
assign g[4503] = a[11] & g[2455];
assign g[6550] = b[11] & g[2455];
assign g[4504] = a[11] & g[2456];
assign g[6551] = b[11] & g[2456];
assign g[4505] = a[11] & g[2457];
assign g[6552] = b[11] & g[2457];
assign g[4506] = a[11] & g[2458];
assign g[6553] = b[11] & g[2458];
assign g[4507] = a[11] & g[2459];
assign g[6554] = b[11] & g[2459];
assign g[4508] = a[11] & g[2460];
assign g[6555] = b[11] & g[2460];
assign g[4509] = a[11] & g[2461];
assign g[6556] = b[11] & g[2461];
assign g[4510] = a[11] & g[2462];
assign g[6557] = b[11] & g[2462];
assign g[4511] = a[11] & g[2463];
assign g[6558] = b[11] & g[2463];
assign g[4512] = a[11] & g[2464];
assign g[6559] = b[11] & g[2464];
assign g[4513] = a[11] & g[2465];
assign g[6560] = b[11] & g[2465];
assign g[4514] = a[11] & g[2466];
assign g[6561] = b[11] & g[2466];
assign g[4515] = a[11] & g[2467];
assign g[6562] = b[11] & g[2467];
assign g[4516] = a[11] & g[2468];
assign g[6563] = b[11] & g[2468];
assign g[4517] = a[11] & g[2469];
assign g[6564] = b[11] & g[2469];
assign g[4518] = a[11] & g[2470];
assign g[6565] = b[11] & g[2470];
assign g[4519] = a[11] & g[2471];
assign g[6566] = b[11] & g[2471];
assign g[4520] = a[11] & g[2472];
assign g[6567] = b[11] & g[2472];
assign g[4521] = a[11] & g[2473];
assign g[6568] = b[11] & g[2473];
assign g[4522] = a[11] & g[2474];
assign g[6569] = b[11] & g[2474];
assign g[4523] = a[11] & g[2475];
assign g[6570] = b[11] & g[2475];
assign g[4524] = a[11] & g[2476];
assign g[6571] = b[11] & g[2476];
assign g[4525] = a[11] & g[2477];
assign g[6572] = b[11] & g[2477];
assign g[4526] = a[11] & g[2478];
assign g[6573] = b[11] & g[2478];
assign g[4527] = a[11] & g[2479];
assign g[6574] = b[11] & g[2479];
assign g[4528] = a[11] & g[2480];
assign g[6575] = b[11] & g[2480];
assign g[4529] = a[11] & g[2481];
assign g[6576] = b[11] & g[2481];
assign g[4530] = a[11] & g[2482];
assign g[6577] = b[11] & g[2482];
assign g[4531] = a[11] & g[2483];
assign g[6578] = b[11] & g[2483];
assign g[4532] = a[11] & g[2484];
assign g[6579] = b[11] & g[2484];
assign g[4533] = a[11] & g[2485];
assign g[6580] = b[11] & g[2485];
assign g[4534] = a[11] & g[2486];
assign g[6581] = b[11] & g[2486];
assign g[4535] = a[11] & g[2487];
assign g[6582] = b[11] & g[2487];
assign g[4536] = a[11] & g[2488];
assign g[6583] = b[11] & g[2488];
assign g[4537] = a[11] & g[2489];
assign g[6584] = b[11] & g[2489];
assign g[4538] = a[11] & g[2490];
assign g[6585] = b[11] & g[2490];
assign g[4539] = a[11] & g[2491];
assign g[6586] = b[11] & g[2491];
assign g[4540] = a[11] & g[2492];
assign g[6587] = b[11] & g[2492];
assign g[4541] = a[11] & g[2493];
assign g[6588] = b[11] & g[2493];
assign g[4542] = a[11] & g[2494];
assign g[6589] = b[11] & g[2494];
assign g[4543] = a[11] & g[2495];
assign g[6590] = b[11] & g[2495];
assign g[4544] = a[11] & g[2496];
assign g[6591] = b[11] & g[2496];
assign g[4545] = a[11] & g[2497];
assign g[6592] = b[11] & g[2497];
assign g[4546] = a[11] & g[2498];
assign g[6593] = b[11] & g[2498];
assign g[4547] = a[11] & g[2499];
assign g[6594] = b[11] & g[2499];
assign g[4548] = a[11] & g[2500];
assign g[6595] = b[11] & g[2500];
assign g[4549] = a[11] & g[2501];
assign g[6596] = b[11] & g[2501];
assign g[4550] = a[11] & g[2502];
assign g[6597] = b[11] & g[2502];
assign g[4551] = a[11] & g[2503];
assign g[6598] = b[11] & g[2503];
assign g[4552] = a[11] & g[2504];
assign g[6599] = b[11] & g[2504];
assign g[4553] = a[11] & g[2505];
assign g[6600] = b[11] & g[2505];
assign g[4554] = a[11] & g[2506];
assign g[6601] = b[11] & g[2506];
assign g[4555] = a[11] & g[2507];
assign g[6602] = b[11] & g[2507];
assign g[4556] = a[11] & g[2508];
assign g[6603] = b[11] & g[2508];
assign g[4557] = a[11] & g[2509];
assign g[6604] = b[11] & g[2509];
assign g[4558] = a[11] & g[2510];
assign g[6605] = b[11] & g[2510];
assign g[4559] = a[11] & g[2511];
assign g[6606] = b[11] & g[2511];
assign g[4560] = a[11] & g[2512];
assign g[6607] = b[11] & g[2512];
assign g[4561] = a[11] & g[2513];
assign g[6608] = b[11] & g[2513];
assign g[4562] = a[11] & g[2514];
assign g[6609] = b[11] & g[2514];
assign g[4563] = a[11] & g[2515];
assign g[6610] = b[11] & g[2515];
assign g[4564] = a[11] & g[2516];
assign g[6611] = b[11] & g[2516];
assign g[4565] = a[11] & g[2517];
assign g[6612] = b[11] & g[2517];
assign g[4566] = a[11] & g[2518];
assign g[6613] = b[11] & g[2518];
assign g[4567] = a[11] & g[2519];
assign g[6614] = b[11] & g[2519];
assign g[4568] = a[11] & g[2520];
assign g[6615] = b[11] & g[2520];
assign g[4569] = a[11] & g[2521];
assign g[6616] = b[11] & g[2521];
assign g[4570] = a[11] & g[2522];
assign g[6617] = b[11] & g[2522];
assign g[4571] = a[11] & g[2523];
assign g[6618] = b[11] & g[2523];
assign g[4572] = a[11] & g[2524];
assign g[6619] = b[11] & g[2524];
assign g[4573] = a[11] & g[2525];
assign g[6620] = b[11] & g[2525];
assign g[4574] = a[11] & g[2526];
assign g[6621] = b[11] & g[2526];
assign g[4575] = a[11] & g[2527];
assign g[6622] = b[11] & g[2527];
assign g[4576] = a[11] & g[2528];
assign g[6623] = b[11] & g[2528];
assign g[4577] = a[11] & g[2529];
assign g[6624] = b[11] & g[2529];
assign g[4578] = a[11] & g[2530];
assign g[6625] = b[11] & g[2530];
assign g[4579] = a[11] & g[2531];
assign g[6626] = b[11] & g[2531];
assign g[4580] = a[11] & g[2532];
assign g[6627] = b[11] & g[2532];
assign g[4581] = a[11] & g[2533];
assign g[6628] = b[11] & g[2533];
assign g[4582] = a[11] & g[2534];
assign g[6629] = b[11] & g[2534];
assign g[4583] = a[11] & g[2535];
assign g[6630] = b[11] & g[2535];
assign g[4584] = a[11] & g[2536];
assign g[6631] = b[11] & g[2536];
assign g[4585] = a[11] & g[2537];
assign g[6632] = b[11] & g[2537];
assign g[4586] = a[11] & g[2538];
assign g[6633] = b[11] & g[2538];
assign g[4587] = a[11] & g[2539];
assign g[6634] = b[11] & g[2539];
assign g[4588] = a[11] & g[2540];
assign g[6635] = b[11] & g[2540];
assign g[4589] = a[11] & g[2541];
assign g[6636] = b[11] & g[2541];
assign g[4590] = a[11] & g[2542];
assign g[6637] = b[11] & g[2542];
assign g[4591] = a[11] & g[2543];
assign g[6638] = b[11] & g[2543];
assign g[4592] = a[11] & g[2544];
assign g[6639] = b[11] & g[2544];
assign g[4593] = a[11] & g[2545];
assign g[6640] = b[11] & g[2545];
assign g[4594] = a[11] & g[2546];
assign g[6641] = b[11] & g[2546];
assign g[4595] = a[11] & g[2547];
assign g[6642] = b[11] & g[2547];
assign g[4596] = a[11] & g[2548];
assign g[6643] = b[11] & g[2548];
assign g[4597] = a[11] & g[2549];
assign g[6644] = b[11] & g[2549];
assign g[4598] = a[11] & g[2550];
assign g[6645] = b[11] & g[2550];
assign g[4599] = a[11] & g[2551];
assign g[6646] = b[11] & g[2551];
assign g[4600] = a[11] & g[2552];
assign g[6647] = b[11] & g[2552];
assign g[4601] = a[11] & g[2553];
assign g[6648] = b[11] & g[2553];
assign g[4602] = a[11] & g[2554];
assign g[6649] = b[11] & g[2554];
assign g[4603] = a[11] & g[2555];
assign g[6650] = b[11] & g[2555];
assign g[4604] = a[11] & g[2556];
assign g[6651] = b[11] & g[2556];
assign g[4605] = a[11] & g[2557];
assign g[6652] = b[11] & g[2557];
assign g[4606] = a[11] & g[2558];
assign g[6653] = b[11] & g[2558];
assign g[4607] = a[11] & g[2559];
assign g[6654] = b[11] & g[2559];
assign g[4608] = a[11] & g[2560];
assign g[6655] = b[11] & g[2560];
assign g[4609] = a[11] & g[2561];
assign g[6656] = b[11] & g[2561];
assign g[4610] = a[11] & g[2562];
assign g[6657] = b[11] & g[2562];
assign g[4611] = a[11] & g[2563];
assign g[6658] = b[11] & g[2563];
assign g[4612] = a[11] & g[2564];
assign g[6659] = b[11] & g[2564];
assign g[4613] = a[11] & g[2565];
assign g[6660] = b[11] & g[2565];
assign g[4614] = a[11] & g[2566];
assign g[6661] = b[11] & g[2566];
assign g[4615] = a[11] & g[2567];
assign g[6662] = b[11] & g[2567];
assign g[4616] = a[11] & g[2568];
assign g[6663] = b[11] & g[2568];
assign g[4617] = a[11] & g[2569];
assign g[6664] = b[11] & g[2569];
assign g[4618] = a[11] & g[2570];
assign g[6665] = b[11] & g[2570];
assign g[4619] = a[11] & g[2571];
assign g[6666] = b[11] & g[2571];
assign g[4620] = a[11] & g[2572];
assign g[6667] = b[11] & g[2572];
assign g[4621] = a[11] & g[2573];
assign g[6668] = b[11] & g[2573];
assign g[4622] = a[11] & g[2574];
assign g[6669] = b[11] & g[2574];
assign g[4623] = a[11] & g[2575];
assign g[6670] = b[11] & g[2575];
assign g[4624] = a[11] & g[2576];
assign g[6671] = b[11] & g[2576];
assign g[4625] = a[11] & g[2577];
assign g[6672] = b[11] & g[2577];
assign g[4626] = a[11] & g[2578];
assign g[6673] = b[11] & g[2578];
assign g[4627] = a[11] & g[2579];
assign g[6674] = b[11] & g[2579];
assign g[4628] = a[11] & g[2580];
assign g[6675] = b[11] & g[2580];
assign g[4629] = a[11] & g[2581];
assign g[6676] = b[11] & g[2581];
assign g[4630] = a[11] & g[2582];
assign g[6677] = b[11] & g[2582];
assign g[4631] = a[11] & g[2583];
assign g[6678] = b[11] & g[2583];
assign g[4632] = a[11] & g[2584];
assign g[6679] = b[11] & g[2584];
assign g[4633] = a[11] & g[2585];
assign g[6680] = b[11] & g[2585];
assign g[4634] = a[11] & g[2586];
assign g[6681] = b[11] & g[2586];
assign g[4635] = a[11] & g[2587];
assign g[6682] = b[11] & g[2587];
assign g[4636] = a[11] & g[2588];
assign g[6683] = b[11] & g[2588];
assign g[4637] = a[11] & g[2589];
assign g[6684] = b[11] & g[2589];
assign g[4638] = a[11] & g[2590];
assign g[6685] = b[11] & g[2590];
assign g[4639] = a[11] & g[2591];
assign g[6686] = b[11] & g[2591];
assign g[4640] = a[11] & g[2592];
assign g[6687] = b[11] & g[2592];
assign g[4641] = a[11] & g[2593];
assign g[6688] = b[11] & g[2593];
assign g[4642] = a[11] & g[2594];
assign g[6689] = b[11] & g[2594];
assign g[4643] = a[11] & g[2595];
assign g[6690] = b[11] & g[2595];
assign g[4644] = a[11] & g[2596];
assign g[6691] = b[11] & g[2596];
assign g[4645] = a[11] & g[2597];
assign g[6692] = b[11] & g[2597];
assign g[4646] = a[11] & g[2598];
assign g[6693] = b[11] & g[2598];
assign g[4647] = a[11] & g[2599];
assign g[6694] = b[11] & g[2599];
assign g[4648] = a[11] & g[2600];
assign g[6695] = b[11] & g[2600];
assign g[4649] = a[11] & g[2601];
assign g[6696] = b[11] & g[2601];
assign g[4650] = a[11] & g[2602];
assign g[6697] = b[11] & g[2602];
assign g[4651] = a[11] & g[2603];
assign g[6698] = b[11] & g[2603];
assign g[4652] = a[11] & g[2604];
assign g[6699] = b[11] & g[2604];
assign g[4653] = a[11] & g[2605];
assign g[6700] = b[11] & g[2605];
assign g[4654] = a[11] & g[2606];
assign g[6701] = b[11] & g[2606];
assign g[4655] = a[11] & g[2607];
assign g[6702] = b[11] & g[2607];
assign g[4656] = a[11] & g[2608];
assign g[6703] = b[11] & g[2608];
assign g[4657] = a[11] & g[2609];
assign g[6704] = b[11] & g[2609];
assign g[4658] = a[11] & g[2610];
assign g[6705] = b[11] & g[2610];
assign g[4659] = a[11] & g[2611];
assign g[6706] = b[11] & g[2611];
assign g[4660] = a[11] & g[2612];
assign g[6707] = b[11] & g[2612];
assign g[4661] = a[11] & g[2613];
assign g[6708] = b[11] & g[2613];
assign g[4662] = a[11] & g[2614];
assign g[6709] = b[11] & g[2614];
assign g[4663] = a[11] & g[2615];
assign g[6710] = b[11] & g[2615];
assign g[4664] = a[11] & g[2616];
assign g[6711] = b[11] & g[2616];
assign g[4665] = a[11] & g[2617];
assign g[6712] = b[11] & g[2617];
assign g[4666] = a[11] & g[2618];
assign g[6713] = b[11] & g[2618];
assign g[4667] = a[11] & g[2619];
assign g[6714] = b[11] & g[2619];
assign g[4668] = a[11] & g[2620];
assign g[6715] = b[11] & g[2620];
assign g[4669] = a[11] & g[2621];
assign g[6716] = b[11] & g[2621];
assign g[4670] = a[11] & g[2622];
assign g[6717] = b[11] & g[2622];
assign g[4671] = a[11] & g[2623];
assign g[6718] = b[11] & g[2623];
assign g[4672] = a[11] & g[2624];
assign g[6719] = b[11] & g[2624];
assign g[4673] = a[11] & g[2625];
assign g[6720] = b[11] & g[2625];
assign g[4674] = a[11] & g[2626];
assign g[6721] = b[11] & g[2626];
assign g[4675] = a[11] & g[2627];
assign g[6722] = b[11] & g[2627];
assign g[4676] = a[11] & g[2628];
assign g[6723] = b[11] & g[2628];
assign g[4677] = a[11] & g[2629];
assign g[6724] = b[11] & g[2629];
assign g[4678] = a[11] & g[2630];
assign g[6725] = b[11] & g[2630];
assign g[4679] = a[11] & g[2631];
assign g[6726] = b[11] & g[2631];
assign g[4680] = a[11] & g[2632];
assign g[6727] = b[11] & g[2632];
assign g[4681] = a[11] & g[2633];
assign g[6728] = b[11] & g[2633];
assign g[4682] = a[11] & g[2634];
assign g[6729] = b[11] & g[2634];
assign g[4683] = a[11] & g[2635];
assign g[6730] = b[11] & g[2635];
assign g[4684] = a[11] & g[2636];
assign g[6731] = b[11] & g[2636];
assign g[4685] = a[11] & g[2637];
assign g[6732] = b[11] & g[2637];
assign g[4686] = a[11] & g[2638];
assign g[6733] = b[11] & g[2638];
assign g[4687] = a[11] & g[2639];
assign g[6734] = b[11] & g[2639];
assign g[4688] = a[11] & g[2640];
assign g[6735] = b[11] & g[2640];
assign g[4689] = a[11] & g[2641];
assign g[6736] = b[11] & g[2641];
assign g[4690] = a[11] & g[2642];
assign g[6737] = b[11] & g[2642];
assign g[4691] = a[11] & g[2643];
assign g[6738] = b[11] & g[2643];
assign g[4692] = a[11] & g[2644];
assign g[6739] = b[11] & g[2644];
assign g[4693] = a[11] & g[2645];
assign g[6740] = b[11] & g[2645];
assign g[4694] = a[11] & g[2646];
assign g[6741] = b[11] & g[2646];
assign g[4695] = a[11] & g[2647];
assign g[6742] = b[11] & g[2647];
assign g[4696] = a[11] & g[2648];
assign g[6743] = b[11] & g[2648];
assign g[4697] = a[11] & g[2649];
assign g[6744] = b[11] & g[2649];
assign g[4698] = a[11] & g[2650];
assign g[6745] = b[11] & g[2650];
assign g[4699] = a[11] & g[2651];
assign g[6746] = b[11] & g[2651];
assign g[4700] = a[11] & g[2652];
assign g[6747] = b[11] & g[2652];
assign g[4701] = a[11] & g[2653];
assign g[6748] = b[11] & g[2653];
assign g[4702] = a[11] & g[2654];
assign g[6749] = b[11] & g[2654];
assign g[4703] = a[11] & g[2655];
assign g[6750] = b[11] & g[2655];
assign g[4704] = a[11] & g[2656];
assign g[6751] = b[11] & g[2656];
assign g[4705] = a[11] & g[2657];
assign g[6752] = b[11] & g[2657];
assign g[4706] = a[11] & g[2658];
assign g[6753] = b[11] & g[2658];
assign g[4707] = a[11] & g[2659];
assign g[6754] = b[11] & g[2659];
assign g[4708] = a[11] & g[2660];
assign g[6755] = b[11] & g[2660];
assign g[4709] = a[11] & g[2661];
assign g[6756] = b[11] & g[2661];
assign g[4710] = a[11] & g[2662];
assign g[6757] = b[11] & g[2662];
assign g[4711] = a[11] & g[2663];
assign g[6758] = b[11] & g[2663];
assign g[4712] = a[11] & g[2664];
assign g[6759] = b[11] & g[2664];
assign g[4713] = a[11] & g[2665];
assign g[6760] = b[11] & g[2665];
assign g[4714] = a[11] & g[2666];
assign g[6761] = b[11] & g[2666];
assign g[4715] = a[11] & g[2667];
assign g[6762] = b[11] & g[2667];
assign g[4716] = a[11] & g[2668];
assign g[6763] = b[11] & g[2668];
assign g[4717] = a[11] & g[2669];
assign g[6764] = b[11] & g[2669];
assign g[4718] = a[11] & g[2670];
assign g[6765] = b[11] & g[2670];
assign g[4719] = a[11] & g[2671];
assign g[6766] = b[11] & g[2671];
assign g[4720] = a[11] & g[2672];
assign g[6767] = b[11] & g[2672];
assign g[4721] = a[11] & g[2673];
assign g[6768] = b[11] & g[2673];
assign g[4722] = a[11] & g[2674];
assign g[6769] = b[11] & g[2674];
assign g[4723] = a[11] & g[2675];
assign g[6770] = b[11] & g[2675];
assign g[4724] = a[11] & g[2676];
assign g[6771] = b[11] & g[2676];
assign g[4725] = a[11] & g[2677];
assign g[6772] = b[11] & g[2677];
assign g[4726] = a[11] & g[2678];
assign g[6773] = b[11] & g[2678];
assign g[4727] = a[11] & g[2679];
assign g[6774] = b[11] & g[2679];
assign g[4728] = a[11] & g[2680];
assign g[6775] = b[11] & g[2680];
assign g[4729] = a[11] & g[2681];
assign g[6776] = b[11] & g[2681];
assign g[4730] = a[11] & g[2682];
assign g[6777] = b[11] & g[2682];
assign g[4731] = a[11] & g[2683];
assign g[6778] = b[11] & g[2683];
assign g[4732] = a[11] & g[2684];
assign g[6779] = b[11] & g[2684];
assign g[4733] = a[11] & g[2685];
assign g[6780] = b[11] & g[2685];
assign g[4734] = a[11] & g[2686];
assign g[6781] = b[11] & g[2686];
assign g[4735] = a[11] & g[2687];
assign g[6782] = b[11] & g[2687];
assign g[4736] = a[11] & g[2688];
assign g[6783] = b[11] & g[2688];
assign g[4737] = a[11] & g[2689];
assign g[6784] = b[11] & g[2689];
assign g[4738] = a[11] & g[2690];
assign g[6785] = b[11] & g[2690];
assign g[4739] = a[11] & g[2691];
assign g[6786] = b[11] & g[2691];
assign g[4740] = a[11] & g[2692];
assign g[6787] = b[11] & g[2692];
assign g[4741] = a[11] & g[2693];
assign g[6788] = b[11] & g[2693];
assign g[4742] = a[11] & g[2694];
assign g[6789] = b[11] & g[2694];
assign g[4743] = a[11] & g[2695];
assign g[6790] = b[11] & g[2695];
assign g[4744] = a[11] & g[2696];
assign g[6791] = b[11] & g[2696];
assign g[4745] = a[11] & g[2697];
assign g[6792] = b[11] & g[2697];
assign g[4746] = a[11] & g[2698];
assign g[6793] = b[11] & g[2698];
assign g[4747] = a[11] & g[2699];
assign g[6794] = b[11] & g[2699];
assign g[4748] = a[11] & g[2700];
assign g[6795] = b[11] & g[2700];
assign g[4749] = a[11] & g[2701];
assign g[6796] = b[11] & g[2701];
assign g[4750] = a[11] & g[2702];
assign g[6797] = b[11] & g[2702];
assign g[4751] = a[11] & g[2703];
assign g[6798] = b[11] & g[2703];
assign g[4752] = a[11] & g[2704];
assign g[6799] = b[11] & g[2704];
assign g[4753] = a[11] & g[2705];
assign g[6800] = b[11] & g[2705];
assign g[4754] = a[11] & g[2706];
assign g[6801] = b[11] & g[2706];
assign g[4755] = a[11] & g[2707];
assign g[6802] = b[11] & g[2707];
assign g[4756] = a[11] & g[2708];
assign g[6803] = b[11] & g[2708];
assign g[4757] = a[11] & g[2709];
assign g[6804] = b[11] & g[2709];
assign g[4758] = a[11] & g[2710];
assign g[6805] = b[11] & g[2710];
assign g[4759] = a[11] & g[2711];
assign g[6806] = b[11] & g[2711];
assign g[4760] = a[11] & g[2712];
assign g[6807] = b[11] & g[2712];
assign g[4761] = a[11] & g[2713];
assign g[6808] = b[11] & g[2713];
assign g[4762] = a[11] & g[2714];
assign g[6809] = b[11] & g[2714];
assign g[4763] = a[11] & g[2715];
assign g[6810] = b[11] & g[2715];
assign g[4764] = a[11] & g[2716];
assign g[6811] = b[11] & g[2716];
assign g[4765] = a[11] & g[2717];
assign g[6812] = b[11] & g[2717];
assign g[4766] = a[11] & g[2718];
assign g[6813] = b[11] & g[2718];
assign g[4767] = a[11] & g[2719];
assign g[6814] = b[11] & g[2719];
assign g[4768] = a[11] & g[2720];
assign g[6815] = b[11] & g[2720];
assign g[4769] = a[11] & g[2721];
assign g[6816] = b[11] & g[2721];
assign g[4770] = a[11] & g[2722];
assign g[6817] = b[11] & g[2722];
assign g[4771] = a[11] & g[2723];
assign g[6818] = b[11] & g[2723];
assign g[4772] = a[11] & g[2724];
assign g[6819] = b[11] & g[2724];
assign g[4773] = a[11] & g[2725];
assign g[6820] = b[11] & g[2725];
assign g[4774] = a[11] & g[2726];
assign g[6821] = b[11] & g[2726];
assign g[4775] = a[11] & g[2727];
assign g[6822] = b[11] & g[2727];
assign g[4776] = a[11] & g[2728];
assign g[6823] = b[11] & g[2728];
assign g[4777] = a[11] & g[2729];
assign g[6824] = b[11] & g[2729];
assign g[4778] = a[11] & g[2730];
assign g[6825] = b[11] & g[2730];
assign g[4779] = a[11] & g[2731];
assign g[6826] = b[11] & g[2731];
assign g[4780] = a[11] & g[2732];
assign g[6827] = b[11] & g[2732];
assign g[4781] = a[11] & g[2733];
assign g[6828] = b[11] & g[2733];
assign g[4782] = a[11] & g[2734];
assign g[6829] = b[11] & g[2734];
assign g[4783] = a[11] & g[2735];
assign g[6830] = b[11] & g[2735];
assign g[4784] = a[11] & g[2736];
assign g[6831] = b[11] & g[2736];
assign g[4785] = a[11] & g[2737];
assign g[6832] = b[11] & g[2737];
assign g[4786] = a[11] & g[2738];
assign g[6833] = b[11] & g[2738];
assign g[4787] = a[11] & g[2739];
assign g[6834] = b[11] & g[2739];
assign g[4788] = a[11] & g[2740];
assign g[6835] = b[11] & g[2740];
assign g[4789] = a[11] & g[2741];
assign g[6836] = b[11] & g[2741];
assign g[4790] = a[11] & g[2742];
assign g[6837] = b[11] & g[2742];
assign g[4791] = a[11] & g[2743];
assign g[6838] = b[11] & g[2743];
assign g[4792] = a[11] & g[2744];
assign g[6839] = b[11] & g[2744];
assign g[4793] = a[11] & g[2745];
assign g[6840] = b[11] & g[2745];
assign g[4794] = a[11] & g[2746];
assign g[6841] = b[11] & g[2746];
assign g[4795] = a[11] & g[2747];
assign g[6842] = b[11] & g[2747];
assign g[4796] = a[11] & g[2748];
assign g[6843] = b[11] & g[2748];
assign g[4797] = a[11] & g[2749];
assign g[6844] = b[11] & g[2749];
assign g[4798] = a[11] & g[2750];
assign g[6845] = b[11] & g[2750];
assign g[4799] = a[11] & g[2751];
assign g[6846] = b[11] & g[2751];
assign g[4800] = a[11] & g[2752];
assign g[6847] = b[11] & g[2752];
assign g[4801] = a[11] & g[2753];
assign g[6848] = b[11] & g[2753];
assign g[4802] = a[11] & g[2754];
assign g[6849] = b[11] & g[2754];
assign g[4803] = a[11] & g[2755];
assign g[6850] = b[11] & g[2755];
assign g[4804] = a[11] & g[2756];
assign g[6851] = b[11] & g[2756];
assign g[4805] = a[11] & g[2757];
assign g[6852] = b[11] & g[2757];
assign g[4806] = a[11] & g[2758];
assign g[6853] = b[11] & g[2758];
assign g[4807] = a[11] & g[2759];
assign g[6854] = b[11] & g[2759];
assign g[4808] = a[11] & g[2760];
assign g[6855] = b[11] & g[2760];
assign g[4809] = a[11] & g[2761];
assign g[6856] = b[11] & g[2761];
assign g[4810] = a[11] & g[2762];
assign g[6857] = b[11] & g[2762];
assign g[4811] = a[11] & g[2763];
assign g[6858] = b[11] & g[2763];
assign g[4812] = a[11] & g[2764];
assign g[6859] = b[11] & g[2764];
assign g[4813] = a[11] & g[2765];
assign g[6860] = b[11] & g[2765];
assign g[4814] = a[11] & g[2766];
assign g[6861] = b[11] & g[2766];
assign g[4815] = a[11] & g[2767];
assign g[6862] = b[11] & g[2767];
assign g[4816] = a[11] & g[2768];
assign g[6863] = b[11] & g[2768];
assign g[4817] = a[11] & g[2769];
assign g[6864] = b[11] & g[2769];
assign g[4818] = a[11] & g[2770];
assign g[6865] = b[11] & g[2770];
assign g[4819] = a[11] & g[2771];
assign g[6866] = b[11] & g[2771];
assign g[4820] = a[11] & g[2772];
assign g[6867] = b[11] & g[2772];
assign g[4821] = a[11] & g[2773];
assign g[6868] = b[11] & g[2773];
assign g[4822] = a[11] & g[2774];
assign g[6869] = b[11] & g[2774];
assign g[4823] = a[11] & g[2775];
assign g[6870] = b[11] & g[2775];
assign g[4824] = a[11] & g[2776];
assign g[6871] = b[11] & g[2776];
assign g[4825] = a[11] & g[2777];
assign g[6872] = b[11] & g[2777];
assign g[4826] = a[11] & g[2778];
assign g[6873] = b[11] & g[2778];
assign g[4827] = a[11] & g[2779];
assign g[6874] = b[11] & g[2779];
assign g[4828] = a[11] & g[2780];
assign g[6875] = b[11] & g[2780];
assign g[4829] = a[11] & g[2781];
assign g[6876] = b[11] & g[2781];
assign g[4830] = a[11] & g[2782];
assign g[6877] = b[11] & g[2782];
assign g[4831] = a[11] & g[2783];
assign g[6878] = b[11] & g[2783];
assign g[4832] = a[11] & g[2784];
assign g[6879] = b[11] & g[2784];
assign g[4833] = a[11] & g[2785];
assign g[6880] = b[11] & g[2785];
assign g[4834] = a[11] & g[2786];
assign g[6881] = b[11] & g[2786];
assign g[4835] = a[11] & g[2787];
assign g[6882] = b[11] & g[2787];
assign g[4836] = a[11] & g[2788];
assign g[6883] = b[11] & g[2788];
assign g[4837] = a[11] & g[2789];
assign g[6884] = b[11] & g[2789];
assign g[4838] = a[11] & g[2790];
assign g[6885] = b[11] & g[2790];
assign g[4839] = a[11] & g[2791];
assign g[6886] = b[11] & g[2791];
assign g[4840] = a[11] & g[2792];
assign g[6887] = b[11] & g[2792];
assign g[4841] = a[11] & g[2793];
assign g[6888] = b[11] & g[2793];
assign g[4842] = a[11] & g[2794];
assign g[6889] = b[11] & g[2794];
assign g[4843] = a[11] & g[2795];
assign g[6890] = b[11] & g[2795];
assign g[4844] = a[11] & g[2796];
assign g[6891] = b[11] & g[2796];
assign g[4845] = a[11] & g[2797];
assign g[6892] = b[11] & g[2797];
assign g[4846] = a[11] & g[2798];
assign g[6893] = b[11] & g[2798];
assign g[4847] = a[11] & g[2799];
assign g[6894] = b[11] & g[2799];
assign g[4848] = a[11] & g[2800];
assign g[6895] = b[11] & g[2800];
assign g[4849] = a[11] & g[2801];
assign g[6896] = b[11] & g[2801];
assign g[4850] = a[11] & g[2802];
assign g[6897] = b[11] & g[2802];
assign g[4851] = a[11] & g[2803];
assign g[6898] = b[11] & g[2803];
assign g[4852] = a[11] & g[2804];
assign g[6899] = b[11] & g[2804];
assign g[4853] = a[11] & g[2805];
assign g[6900] = b[11] & g[2805];
assign g[4854] = a[11] & g[2806];
assign g[6901] = b[11] & g[2806];
assign g[4855] = a[11] & g[2807];
assign g[6902] = b[11] & g[2807];
assign g[4856] = a[11] & g[2808];
assign g[6903] = b[11] & g[2808];
assign g[4857] = a[11] & g[2809];
assign g[6904] = b[11] & g[2809];
assign g[4858] = a[11] & g[2810];
assign g[6905] = b[11] & g[2810];
assign g[4859] = a[11] & g[2811];
assign g[6906] = b[11] & g[2811];
assign g[4860] = a[11] & g[2812];
assign g[6907] = b[11] & g[2812];
assign g[4861] = a[11] & g[2813];
assign g[6908] = b[11] & g[2813];
assign g[4862] = a[11] & g[2814];
assign g[6909] = b[11] & g[2814];
assign g[4863] = a[11] & g[2815];
assign g[6910] = b[11] & g[2815];
assign g[4864] = a[11] & g[2816];
assign g[6911] = b[11] & g[2816];
assign g[4865] = a[11] & g[2817];
assign g[6912] = b[11] & g[2817];
assign g[4866] = a[11] & g[2818];
assign g[6913] = b[11] & g[2818];
assign g[4867] = a[11] & g[2819];
assign g[6914] = b[11] & g[2819];
assign g[4868] = a[11] & g[2820];
assign g[6915] = b[11] & g[2820];
assign g[4869] = a[11] & g[2821];
assign g[6916] = b[11] & g[2821];
assign g[4870] = a[11] & g[2822];
assign g[6917] = b[11] & g[2822];
assign g[4871] = a[11] & g[2823];
assign g[6918] = b[11] & g[2823];
assign g[4872] = a[11] & g[2824];
assign g[6919] = b[11] & g[2824];
assign g[4873] = a[11] & g[2825];
assign g[6920] = b[11] & g[2825];
assign g[4874] = a[11] & g[2826];
assign g[6921] = b[11] & g[2826];
assign g[4875] = a[11] & g[2827];
assign g[6922] = b[11] & g[2827];
assign g[4876] = a[11] & g[2828];
assign g[6923] = b[11] & g[2828];
assign g[4877] = a[11] & g[2829];
assign g[6924] = b[11] & g[2829];
assign g[4878] = a[11] & g[2830];
assign g[6925] = b[11] & g[2830];
assign g[4879] = a[11] & g[2831];
assign g[6926] = b[11] & g[2831];
assign g[4880] = a[11] & g[2832];
assign g[6927] = b[11] & g[2832];
assign g[4881] = a[11] & g[2833];
assign g[6928] = b[11] & g[2833];
assign g[4882] = a[11] & g[2834];
assign g[6929] = b[11] & g[2834];
assign g[4883] = a[11] & g[2835];
assign g[6930] = b[11] & g[2835];
assign g[4884] = a[11] & g[2836];
assign g[6931] = b[11] & g[2836];
assign g[4885] = a[11] & g[2837];
assign g[6932] = b[11] & g[2837];
assign g[4886] = a[11] & g[2838];
assign g[6933] = b[11] & g[2838];
assign g[4887] = a[11] & g[2839];
assign g[6934] = b[11] & g[2839];
assign g[4888] = a[11] & g[2840];
assign g[6935] = b[11] & g[2840];
assign g[4889] = a[11] & g[2841];
assign g[6936] = b[11] & g[2841];
assign g[4890] = a[11] & g[2842];
assign g[6937] = b[11] & g[2842];
assign g[4891] = a[11] & g[2843];
assign g[6938] = b[11] & g[2843];
assign g[4892] = a[11] & g[2844];
assign g[6939] = b[11] & g[2844];
assign g[4893] = a[11] & g[2845];
assign g[6940] = b[11] & g[2845];
assign g[4894] = a[11] & g[2846];
assign g[6941] = b[11] & g[2846];
assign g[4895] = a[11] & g[2847];
assign g[6942] = b[11] & g[2847];
assign g[4896] = a[11] & g[2848];
assign g[6943] = b[11] & g[2848];
assign g[4897] = a[11] & g[2849];
assign g[6944] = b[11] & g[2849];
assign g[4898] = a[11] & g[2850];
assign g[6945] = b[11] & g[2850];
assign g[4899] = a[11] & g[2851];
assign g[6946] = b[11] & g[2851];
assign g[4900] = a[11] & g[2852];
assign g[6947] = b[11] & g[2852];
assign g[4901] = a[11] & g[2853];
assign g[6948] = b[11] & g[2853];
assign g[4902] = a[11] & g[2854];
assign g[6949] = b[11] & g[2854];
assign g[4903] = a[11] & g[2855];
assign g[6950] = b[11] & g[2855];
assign g[4904] = a[11] & g[2856];
assign g[6951] = b[11] & g[2856];
assign g[4905] = a[11] & g[2857];
assign g[6952] = b[11] & g[2857];
assign g[4906] = a[11] & g[2858];
assign g[6953] = b[11] & g[2858];
assign g[4907] = a[11] & g[2859];
assign g[6954] = b[11] & g[2859];
assign g[4908] = a[11] & g[2860];
assign g[6955] = b[11] & g[2860];
assign g[4909] = a[11] & g[2861];
assign g[6956] = b[11] & g[2861];
assign g[4910] = a[11] & g[2862];
assign g[6957] = b[11] & g[2862];
assign g[4911] = a[11] & g[2863];
assign g[6958] = b[11] & g[2863];
assign g[4912] = a[11] & g[2864];
assign g[6959] = b[11] & g[2864];
assign g[4913] = a[11] & g[2865];
assign g[6960] = b[11] & g[2865];
assign g[4914] = a[11] & g[2866];
assign g[6961] = b[11] & g[2866];
assign g[4915] = a[11] & g[2867];
assign g[6962] = b[11] & g[2867];
assign g[4916] = a[11] & g[2868];
assign g[6963] = b[11] & g[2868];
assign g[4917] = a[11] & g[2869];
assign g[6964] = b[11] & g[2869];
assign g[4918] = a[11] & g[2870];
assign g[6965] = b[11] & g[2870];
assign g[4919] = a[11] & g[2871];
assign g[6966] = b[11] & g[2871];
assign g[4920] = a[11] & g[2872];
assign g[6967] = b[11] & g[2872];
assign g[4921] = a[11] & g[2873];
assign g[6968] = b[11] & g[2873];
assign g[4922] = a[11] & g[2874];
assign g[6969] = b[11] & g[2874];
assign g[4923] = a[11] & g[2875];
assign g[6970] = b[11] & g[2875];
assign g[4924] = a[11] & g[2876];
assign g[6971] = b[11] & g[2876];
assign g[4925] = a[11] & g[2877];
assign g[6972] = b[11] & g[2877];
assign g[4926] = a[11] & g[2878];
assign g[6973] = b[11] & g[2878];
assign g[4927] = a[11] & g[2879];
assign g[6974] = b[11] & g[2879];
assign g[4928] = a[11] & g[2880];
assign g[6975] = b[11] & g[2880];
assign g[4929] = a[11] & g[2881];
assign g[6976] = b[11] & g[2881];
assign g[4930] = a[11] & g[2882];
assign g[6977] = b[11] & g[2882];
assign g[4931] = a[11] & g[2883];
assign g[6978] = b[11] & g[2883];
assign g[4932] = a[11] & g[2884];
assign g[6979] = b[11] & g[2884];
assign g[4933] = a[11] & g[2885];
assign g[6980] = b[11] & g[2885];
assign g[4934] = a[11] & g[2886];
assign g[6981] = b[11] & g[2886];
assign g[4935] = a[11] & g[2887];
assign g[6982] = b[11] & g[2887];
assign g[4936] = a[11] & g[2888];
assign g[6983] = b[11] & g[2888];
assign g[4937] = a[11] & g[2889];
assign g[6984] = b[11] & g[2889];
assign g[4938] = a[11] & g[2890];
assign g[6985] = b[11] & g[2890];
assign g[4939] = a[11] & g[2891];
assign g[6986] = b[11] & g[2891];
assign g[4940] = a[11] & g[2892];
assign g[6987] = b[11] & g[2892];
assign g[4941] = a[11] & g[2893];
assign g[6988] = b[11] & g[2893];
assign g[4942] = a[11] & g[2894];
assign g[6989] = b[11] & g[2894];
assign g[4943] = a[11] & g[2895];
assign g[6990] = b[11] & g[2895];
assign g[4944] = a[11] & g[2896];
assign g[6991] = b[11] & g[2896];
assign g[4945] = a[11] & g[2897];
assign g[6992] = b[11] & g[2897];
assign g[4946] = a[11] & g[2898];
assign g[6993] = b[11] & g[2898];
assign g[4947] = a[11] & g[2899];
assign g[6994] = b[11] & g[2899];
assign g[4948] = a[11] & g[2900];
assign g[6995] = b[11] & g[2900];
assign g[4949] = a[11] & g[2901];
assign g[6996] = b[11] & g[2901];
assign g[4950] = a[11] & g[2902];
assign g[6997] = b[11] & g[2902];
assign g[4951] = a[11] & g[2903];
assign g[6998] = b[11] & g[2903];
assign g[4952] = a[11] & g[2904];
assign g[6999] = b[11] & g[2904];
assign g[4953] = a[11] & g[2905];
assign g[7000] = b[11] & g[2905];
assign g[4954] = a[11] & g[2906];
assign g[7001] = b[11] & g[2906];
assign g[4955] = a[11] & g[2907];
assign g[7002] = b[11] & g[2907];
assign g[4956] = a[11] & g[2908];
assign g[7003] = b[11] & g[2908];
assign g[4957] = a[11] & g[2909];
assign g[7004] = b[11] & g[2909];
assign g[4958] = a[11] & g[2910];
assign g[7005] = b[11] & g[2910];
assign g[4959] = a[11] & g[2911];
assign g[7006] = b[11] & g[2911];
assign g[4960] = a[11] & g[2912];
assign g[7007] = b[11] & g[2912];
assign g[4961] = a[11] & g[2913];
assign g[7008] = b[11] & g[2913];
assign g[4962] = a[11] & g[2914];
assign g[7009] = b[11] & g[2914];
assign g[4963] = a[11] & g[2915];
assign g[7010] = b[11] & g[2915];
assign g[4964] = a[11] & g[2916];
assign g[7011] = b[11] & g[2916];
assign g[4965] = a[11] & g[2917];
assign g[7012] = b[11] & g[2917];
assign g[4966] = a[11] & g[2918];
assign g[7013] = b[11] & g[2918];
assign g[4967] = a[11] & g[2919];
assign g[7014] = b[11] & g[2919];
assign g[4968] = a[11] & g[2920];
assign g[7015] = b[11] & g[2920];
assign g[4969] = a[11] & g[2921];
assign g[7016] = b[11] & g[2921];
assign g[4970] = a[11] & g[2922];
assign g[7017] = b[11] & g[2922];
assign g[4971] = a[11] & g[2923];
assign g[7018] = b[11] & g[2923];
assign g[4972] = a[11] & g[2924];
assign g[7019] = b[11] & g[2924];
assign g[4973] = a[11] & g[2925];
assign g[7020] = b[11] & g[2925];
assign g[4974] = a[11] & g[2926];
assign g[7021] = b[11] & g[2926];
assign g[4975] = a[11] & g[2927];
assign g[7022] = b[11] & g[2927];
assign g[4976] = a[11] & g[2928];
assign g[7023] = b[11] & g[2928];
assign g[4977] = a[11] & g[2929];
assign g[7024] = b[11] & g[2929];
assign g[4978] = a[11] & g[2930];
assign g[7025] = b[11] & g[2930];
assign g[4979] = a[11] & g[2931];
assign g[7026] = b[11] & g[2931];
assign g[4980] = a[11] & g[2932];
assign g[7027] = b[11] & g[2932];
assign g[4981] = a[11] & g[2933];
assign g[7028] = b[11] & g[2933];
assign g[4982] = a[11] & g[2934];
assign g[7029] = b[11] & g[2934];
assign g[4983] = a[11] & g[2935];
assign g[7030] = b[11] & g[2935];
assign g[4984] = a[11] & g[2936];
assign g[7031] = b[11] & g[2936];
assign g[4985] = a[11] & g[2937];
assign g[7032] = b[11] & g[2937];
assign g[4986] = a[11] & g[2938];
assign g[7033] = b[11] & g[2938];
assign g[4987] = a[11] & g[2939];
assign g[7034] = b[11] & g[2939];
assign g[4988] = a[11] & g[2940];
assign g[7035] = b[11] & g[2940];
assign g[4989] = a[11] & g[2941];
assign g[7036] = b[11] & g[2941];
assign g[4990] = a[11] & g[2942];
assign g[7037] = b[11] & g[2942];
assign g[4991] = a[11] & g[2943];
assign g[7038] = b[11] & g[2943];
assign g[4992] = a[11] & g[2944];
assign g[7039] = b[11] & g[2944];
assign g[4993] = a[11] & g[2945];
assign g[7040] = b[11] & g[2945];
assign g[4994] = a[11] & g[2946];
assign g[7041] = b[11] & g[2946];
assign g[4995] = a[11] & g[2947];
assign g[7042] = b[11] & g[2947];
assign g[4996] = a[11] & g[2948];
assign g[7043] = b[11] & g[2948];
assign g[4997] = a[11] & g[2949];
assign g[7044] = b[11] & g[2949];
assign g[4998] = a[11] & g[2950];
assign g[7045] = b[11] & g[2950];
assign g[4999] = a[11] & g[2951];
assign g[7046] = b[11] & g[2951];
assign g[5000] = a[11] & g[2952];
assign g[7047] = b[11] & g[2952];
assign g[5001] = a[11] & g[2953];
assign g[7048] = b[11] & g[2953];
assign g[5002] = a[11] & g[2954];
assign g[7049] = b[11] & g[2954];
assign g[5003] = a[11] & g[2955];
assign g[7050] = b[11] & g[2955];
assign g[5004] = a[11] & g[2956];
assign g[7051] = b[11] & g[2956];
assign g[5005] = a[11] & g[2957];
assign g[7052] = b[11] & g[2957];
assign g[5006] = a[11] & g[2958];
assign g[7053] = b[11] & g[2958];
assign g[5007] = a[11] & g[2959];
assign g[7054] = b[11] & g[2959];
assign g[5008] = a[11] & g[2960];
assign g[7055] = b[11] & g[2960];
assign g[5009] = a[11] & g[2961];
assign g[7056] = b[11] & g[2961];
assign g[5010] = a[11] & g[2962];
assign g[7057] = b[11] & g[2962];
assign g[5011] = a[11] & g[2963];
assign g[7058] = b[11] & g[2963];
assign g[5012] = a[11] & g[2964];
assign g[7059] = b[11] & g[2964];
assign g[5013] = a[11] & g[2965];
assign g[7060] = b[11] & g[2965];
assign g[5014] = a[11] & g[2966];
assign g[7061] = b[11] & g[2966];
assign g[5015] = a[11] & g[2967];
assign g[7062] = b[11] & g[2967];
assign g[5016] = a[11] & g[2968];
assign g[7063] = b[11] & g[2968];
assign g[5017] = a[11] & g[2969];
assign g[7064] = b[11] & g[2969];
assign g[5018] = a[11] & g[2970];
assign g[7065] = b[11] & g[2970];
assign g[5019] = a[11] & g[2971];
assign g[7066] = b[11] & g[2971];
assign g[5020] = a[11] & g[2972];
assign g[7067] = b[11] & g[2972];
assign g[5021] = a[11] & g[2973];
assign g[7068] = b[11] & g[2973];
assign g[5022] = a[11] & g[2974];
assign g[7069] = b[11] & g[2974];
assign g[5023] = a[11] & g[2975];
assign g[7070] = b[11] & g[2975];
assign g[5024] = a[11] & g[2976];
assign g[7071] = b[11] & g[2976];
assign g[5025] = a[11] & g[2977];
assign g[7072] = b[11] & g[2977];
assign g[5026] = a[11] & g[2978];
assign g[7073] = b[11] & g[2978];
assign g[5027] = a[11] & g[2979];
assign g[7074] = b[11] & g[2979];
assign g[5028] = a[11] & g[2980];
assign g[7075] = b[11] & g[2980];
assign g[5029] = a[11] & g[2981];
assign g[7076] = b[11] & g[2981];
assign g[5030] = a[11] & g[2982];
assign g[7077] = b[11] & g[2982];
assign g[5031] = a[11] & g[2983];
assign g[7078] = b[11] & g[2983];
assign g[5032] = a[11] & g[2984];
assign g[7079] = b[11] & g[2984];
assign g[5033] = a[11] & g[2985];
assign g[7080] = b[11] & g[2985];
assign g[5034] = a[11] & g[2986];
assign g[7081] = b[11] & g[2986];
assign g[5035] = a[11] & g[2987];
assign g[7082] = b[11] & g[2987];
assign g[5036] = a[11] & g[2988];
assign g[7083] = b[11] & g[2988];
assign g[5037] = a[11] & g[2989];
assign g[7084] = b[11] & g[2989];
assign g[5038] = a[11] & g[2990];
assign g[7085] = b[11] & g[2990];
assign g[5039] = a[11] & g[2991];
assign g[7086] = b[11] & g[2991];
assign g[5040] = a[11] & g[2992];
assign g[7087] = b[11] & g[2992];
assign g[5041] = a[11] & g[2993];
assign g[7088] = b[11] & g[2993];
assign g[5042] = a[11] & g[2994];
assign g[7089] = b[11] & g[2994];
assign g[5043] = a[11] & g[2995];
assign g[7090] = b[11] & g[2995];
assign g[5044] = a[11] & g[2996];
assign g[7091] = b[11] & g[2996];
assign g[5045] = a[11] & g[2997];
assign g[7092] = b[11] & g[2997];
assign g[5046] = a[11] & g[2998];
assign g[7093] = b[11] & g[2998];
assign g[5047] = a[11] & g[2999];
assign g[7094] = b[11] & g[2999];
assign g[5048] = a[11] & g[3000];
assign g[7095] = b[11] & g[3000];
assign g[5049] = a[11] & g[3001];
assign g[7096] = b[11] & g[3001];
assign g[5050] = a[11] & g[3002];
assign g[7097] = b[11] & g[3002];
assign g[5051] = a[11] & g[3003];
assign g[7098] = b[11] & g[3003];
assign g[5052] = a[11] & g[3004];
assign g[7099] = b[11] & g[3004];
assign g[5053] = a[11] & g[3005];
assign g[7100] = b[11] & g[3005];
assign g[5054] = a[11] & g[3006];
assign g[7101] = b[11] & g[3006];
assign g[5055] = a[11] & g[3007];
assign g[7102] = b[11] & g[3007];
assign g[5056] = a[11] & g[3008];
assign g[7103] = b[11] & g[3008];
assign g[5057] = a[11] & g[3009];
assign g[7104] = b[11] & g[3009];
assign g[5058] = a[11] & g[3010];
assign g[7105] = b[11] & g[3010];
assign g[5059] = a[11] & g[3011];
assign g[7106] = b[11] & g[3011];
assign g[5060] = a[11] & g[3012];
assign g[7107] = b[11] & g[3012];
assign g[5061] = a[11] & g[3013];
assign g[7108] = b[11] & g[3013];
assign g[5062] = a[11] & g[3014];
assign g[7109] = b[11] & g[3014];
assign g[5063] = a[11] & g[3015];
assign g[7110] = b[11] & g[3015];
assign g[5064] = a[11] & g[3016];
assign g[7111] = b[11] & g[3016];
assign g[5065] = a[11] & g[3017];
assign g[7112] = b[11] & g[3017];
assign g[5066] = a[11] & g[3018];
assign g[7113] = b[11] & g[3018];
assign g[5067] = a[11] & g[3019];
assign g[7114] = b[11] & g[3019];
assign g[5068] = a[11] & g[3020];
assign g[7115] = b[11] & g[3020];
assign g[5069] = a[11] & g[3021];
assign g[7116] = b[11] & g[3021];
assign g[5070] = a[11] & g[3022];
assign g[7117] = b[11] & g[3022];
assign g[5071] = a[11] & g[3023];
assign g[7118] = b[11] & g[3023];
assign g[5072] = a[11] & g[3024];
assign g[7119] = b[11] & g[3024];
assign g[5073] = a[11] & g[3025];
assign g[7120] = b[11] & g[3025];
assign g[5074] = a[11] & g[3026];
assign g[7121] = b[11] & g[3026];
assign g[5075] = a[11] & g[3027];
assign g[7122] = b[11] & g[3027];
assign g[5076] = a[11] & g[3028];
assign g[7123] = b[11] & g[3028];
assign g[5077] = a[11] & g[3029];
assign g[7124] = b[11] & g[3029];
assign g[5078] = a[11] & g[3030];
assign g[7125] = b[11] & g[3030];
assign g[5079] = a[11] & g[3031];
assign g[7126] = b[11] & g[3031];
assign g[5080] = a[11] & g[3032];
assign g[7127] = b[11] & g[3032];
assign g[5081] = a[11] & g[3033];
assign g[7128] = b[11] & g[3033];
assign g[5082] = a[11] & g[3034];
assign g[7129] = b[11] & g[3034];
assign g[5083] = a[11] & g[3035];
assign g[7130] = b[11] & g[3035];
assign g[5084] = a[11] & g[3036];
assign g[7131] = b[11] & g[3036];
assign g[5085] = a[11] & g[3037];
assign g[7132] = b[11] & g[3037];
assign g[5086] = a[11] & g[3038];
assign g[7133] = b[11] & g[3038];
assign g[5087] = a[11] & g[3039];
assign g[7134] = b[11] & g[3039];
assign g[5088] = a[11] & g[3040];
assign g[7135] = b[11] & g[3040];
assign g[5089] = a[11] & g[3041];
assign g[7136] = b[11] & g[3041];
assign g[5090] = a[11] & g[3042];
assign g[7137] = b[11] & g[3042];
assign g[5091] = a[11] & g[3043];
assign g[7138] = b[11] & g[3043];
assign g[5092] = a[11] & g[3044];
assign g[7139] = b[11] & g[3044];
assign g[5093] = a[11] & g[3045];
assign g[7140] = b[11] & g[3045];
assign g[5094] = a[11] & g[3046];
assign g[7141] = b[11] & g[3046];
assign g[5095] = a[11] & g[3047];
assign g[7142] = b[11] & g[3047];
assign g[5096] = a[11] & g[3048];
assign g[7143] = b[11] & g[3048];
assign g[5097] = a[11] & g[3049];
assign g[7144] = b[11] & g[3049];
assign g[5098] = a[11] & g[3050];
assign g[7145] = b[11] & g[3050];
assign g[5099] = a[11] & g[3051];
assign g[7146] = b[11] & g[3051];
assign g[5100] = a[11] & g[3052];
assign g[7147] = b[11] & g[3052];
assign g[5101] = a[11] & g[3053];
assign g[7148] = b[11] & g[3053];
assign g[5102] = a[11] & g[3054];
assign g[7149] = b[11] & g[3054];
assign g[5103] = a[11] & g[3055];
assign g[7150] = b[11] & g[3055];
assign g[5104] = a[11] & g[3056];
assign g[7151] = b[11] & g[3056];
assign g[5105] = a[11] & g[3057];
assign g[7152] = b[11] & g[3057];
assign g[5106] = a[11] & g[3058];
assign g[7153] = b[11] & g[3058];
assign g[5107] = a[11] & g[3059];
assign g[7154] = b[11] & g[3059];
assign g[5108] = a[11] & g[3060];
assign g[7155] = b[11] & g[3060];
assign g[5109] = a[11] & g[3061];
assign g[7156] = b[11] & g[3061];
assign g[5110] = a[11] & g[3062];
assign g[7157] = b[11] & g[3062];
assign g[5111] = a[11] & g[3063];
assign g[7158] = b[11] & g[3063];
assign g[5112] = a[11] & g[3064];
assign g[7159] = b[11] & g[3064];
assign g[5113] = a[11] & g[3065];
assign g[7160] = b[11] & g[3065];
assign g[5114] = a[11] & g[3066];
assign g[7161] = b[11] & g[3066];
assign g[5115] = a[11] & g[3067];
assign g[7162] = b[11] & g[3067];
assign g[5116] = a[11] & g[3068];
assign g[7163] = b[11] & g[3068];
assign g[5117] = a[11] & g[3069];
assign g[7164] = b[11] & g[3069];
assign g[5118] = a[11] & g[3070];
assign g[7165] = b[11] & g[3070];
assign g[5119] = a[11] & g[3071];
assign g[7166] = b[11] & g[3071];
assign g[5120] = a[11] & g[3072];
assign g[7167] = b[11] & g[3072];
assign g[5121] = a[11] & g[3073];
assign g[7168] = b[11] & g[3073];
assign g[5122] = a[11] & g[3074];
assign g[7169] = b[11] & g[3074];
assign g[5123] = a[11] & g[3075];
assign g[7170] = b[11] & g[3075];
assign g[5124] = a[11] & g[3076];
assign g[7171] = b[11] & g[3076];
assign g[5125] = a[11] & g[3077];
assign g[7172] = b[11] & g[3077];
assign g[5126] = a[11] & g[3078];
assign g[7173] = b[11] & g[3078];
assign g[5127] = a[11] & g[3079];
assign g[7174] = b[11] & g[3079];
assign g[5128] = a[11] & g[3080];
assign g[7175] = b[11] & g[3080];
assign g[5129] = a[11] & g[3081];
assign g[7176] = b[11] & g[3081];
assign g[5130] = a[11] & g[3082];
assign g[7177] = b[11] & g[3082];
assign g[5131] = a[11] & g[3083];
assign g[7178] = b[11] & g[3083];
assign g[5132] = a[11] & g[3084];
assign g[7179] = b[11] & g[3084];
assign g[5133] = a[11] & g[3085];
assign g[7180] = b[11] & g[3085];
assign g[5134] = a[11] & g[3086];
assign g[7181] = b[11] & g[3086];
assign g[5135] = a[11] & g[3087];
assign g[7182] = b[11] & g[3087];
assign g[5136] = a[11] & g[3088];
assign g[7183] = b[11] & g[3088];
assign g[5137] = a[11] & g[3089];
assign g[7184] = b[11] & g[3089];
assign g[5138] = a[11] & g[3090];
assign g[7185] = b[11] & g[3090];
assign g[5139] = a[11] & g[3091];
assign g[7186] = b[11] & g[3091];
assign g[5140] = a[11] & g[3092];
assign g[7187] = b[11] & g[3092];
assign g[5141] = a[11] & g[3093];
assign g[7188] = b[11] & g[3093];
assign g[5142] = a[11] & g[3094];
assign g[7189] = b[11] & g[3094];
assign g[5143] = a[11] & g[3095];
assign g[7190] = b[11] & g[3095];
assign g[5144] = a[11] & g[3096];
assign g[7191] = b[11] & g[3096];
assign g[5145] = a[11] & g[3097];
assign g[7192] = b[11] & g[3097];
assign g[5146] = a[11] & g[3098];
assign g[7193] = b[11] & g[3098];
assign g[5147] = a[11] & g[3099];
assign g[7194] = b[11] & g[3099];
assign g[5148] = a[11] & g[3100];
assign g[7195] = b[11] & g[3100];
assign g[5149] = a[11] & g[3101];
assign g[7196] = b[11] & g[3101];
assign g[5150] = a[11] & g[3102];
assign g[7197] = b[11] & g[3102];
assign g[5151] = a[11] & g[3103];
assign g[7198] = b[11] & g[3103];
assign g[5152] = a[11] & g[3104];
assign g[7199] = b[11] & g[3104];
assign g[5153] = a[11] & g[3105];
assign g[7200] = b[11] & g[3105];
assign g[5154] = a[11] & g[3106];
assign g[7201] = b[11] & g[3106];
assign g[5155] = a[11] & g[3107];
assign g[7202] = b[11] & g[3107];
assign g[5156] = a[11] & g[3108];
assign g[7203] = b[11] & g[3108];
assign g[5157] = a[11] & g[3109];
assign g[7204] = b[11] & g[3109];
assign g[5158] = a[11] & g[3110];
assign g[7205] = b[11] & g[3110];
assign g[5159] = a[11] & g[3111];
assign g[7206] = b[11] & g[3111];
assign g[5160] = a[11] & g[3112];
assign g[7207] = b[11] & g[3112];
assign g[5161] = a[11] & g[3113];
assign g[7208] = b[11] & g[3113];
assign g[5162] = a[11] & g[3114];
assign g[7209] = b[11] & g[3114];
assign g[5163] = a[11] & g[3115];
assign g[7210] = b[11] & g[3115];
assign g[5164] = a[11] & g[3116];
assign g[7211] = b[11] & g[3116];
assign g[5165] = a[11] & g[3117];
assign g[7212] = b[11] & g[3117];
assign g[5166] = a[11] & g[3118];
assign g[7213] = b[11] & g[3118];
assign g[5167] = a[11] & g[3119];
assign g[7214] = b[11] & g[3119];
assign g[5168] = a[11] & g[3120];
assign g[7215] = b[11] & g[3120];
assign g[5169] = a[11] & g[3121];
assign g[7216] = b[11] & g[3121];
assign g[5170] = a[11] & g[3122];
assign g[7217] = b[11] & g[3122];
assign g[5171] = a[11] & g[3123];
assign g[7218] = b[11] & g[3123];
assign g[5172] = a[11] & g[3124];
assign g[7219] = b[11] & g[3124];
assign g[5173] = a[11] & g[3125];
assign g[7220] = b[11] & g[3125];
assign g[5174] = a[11] & g[3126];
assign g[7221] = b[11] & g[3126];
assign g[5175] = a[11] & g[3127];
assign g[7222] = b[11] & g[3127];
assign g[5176] = a[11] & g[3128];
assign g[7223] = b[11] & g[3128];
assign g[5177] = a[11] & g[3129];
assign g[7224] = b[11] & g[3129];
assign g[5178] = a[11] & g[3130];
assign g[7225] = b[11] & g[3130];
assign g[5179] = a[11] & g[3131];
assign g[7226] = b[11] & g[3131];
assign g[5180] = a[11] & g[3132];
assign g[7227] = b[11] & g[3132];
assign g[5181] = a[11] & g[3133];
assign g[7228] = b[11] & g[3133];
assign g[5182] = a[11] & g[3134];
assign g[7229] = b[11] & g[3134];
assign g[5183] = a[11] & g[3135];
assign g[7230] = b[11] & g[3135];
assign g[5184] = a[11] & g[3136];
assign g[7231] = b[11] & g[3136];
assign g[5185] = a[11] & g[3137];
assign g[7232] = b[11] & g[3137];
assign g[5186] = a[11] & g[3138];
assign g[7233] = b[11] & g[3138];
assign g[5187] = a[11] & g[3139];
assign g[7234] = b[11] & g[3139];
assign g[5188] = a[11] & g[3140];
assign g[7235] = b[11] & g[3140];
assign g[5189] = a[11] & g[3141];
assign g[7236] = b[11] & g[3141];
assign g[5190] = a[11] & g[3142];
assign g[7237] = b[11] & g[3142];
assign g[5191] = a[11] & g[3143];
assign g[7238] = b[11] & g[3143];
assign g[5192] = a[11] & g[3144];
assign g[7239] = b[11] & g[3144];
assign g[5193] = a[11] & g[3145];
assign g[7240] = b[11] & g[3145];
assign g[5194] = a[11] & g[3146];
assign g[7241] = b[11] & g[3146];
assign g[5195] = a[11] & g[3147];
assign g[7242] = b[11] & g[3147];
assign g[5196] = a[11] & g[3148];
assign g[7243] = b[11] & g[3148];
assign g[5197] = a[11] & g[3149];
assign g[7244] = b[11] & g[3149];
assign g[5198] = a[11] & g[3150];
assign g[7245] = b[11] & g[3150];
assign g[5199] = a[11] & g[3151];
assign g[7246] = b[11] & g[3151];
assign g[5200] = a[11] & g[3152];
assign g[7247] = b[11] & g[3152];
assign g[5201] = a[11] & g[3153];
assign g[7248] = b[11] & g[3153];
assign g[5202] = a[11] & g[3154];
assign g[7249] = b[11] & g[3154];
assign g[5203] = a[11] & g[3155];
assign g[7250] = b[11] & g[3155];
assign g[5204] = a[11] & g[3156];
assign g[7251] = b[11] & g[3156];
assign g[5205] = a[11] & g[3157];
assign g[7252] = b[11] & g[3157];
assign g[5206] = a[11] & g[3158];
assign g[7253] = b[11] & g[3158];
assign g[5207] = a[11] & g[3159];
assign g[7254] = b[11] & g[3159];
assign g[5208] = a[11] & g[3160];
assign g[7255] = b[11] & g[3160];
assign g[5209] = a[11] & g[3161];
assign g[7256] = b[11] & g[3161];
assign g[5210] = a[11] & g[3162];
assign g[7257] = b[11] & g[3162];
assign g[5211] = a[11] & g[3163];
assign g[7258] = b[11] & g[3163];
assign g[5212] = a[11] & g[3164];
assign g[7259] = b[11] & g[3164];
assign g[5213] = a[11] & g[3165];
assign g[7260] = b[11] & g[3165];
assign g[5214] = a[11] & g[3166];
assign g[7261] = b[11] & g[3166];
assign g[5215] = a[11] & g[3167];
assign g[7262] = b[11] & g[3167];
assign g[5216] = a[11] & g[3168];
assign g[7263] = b[11] & g[3168];
assign g[5217] = a[11] & g[3169];
assign g[7264] = b[11] & g[3169];
assign g[5218] = a[11] & g[3170];
assign g[7265] = b[11] & g[3170];
assign g[5219] = a[11] & g[3171];
assign g[7266] = b[11] & g[3171];
assign g[5220] = a[11] & g[3172];
assign g[7267] = b[11] & g[3172];
assign g[5221] = a[11] & g[3173];
assign g[7268] = b[11] & g[3173];
assign g[5222] = a[11] & g[3174];
assign g[7269] = b[11] & g[3174];
assign g[5223] = a[11] & g[3175];
assign g[7270] = b[11] & g[3175];
assign g[5224] = a[11] & g[3176];
assign g[7271] = b[11] & g[3176];
assign g[5225] = a[11] & g[3177];
assign g[7272] = b[11] & g[3177];
assign g[5226] = a[11] & g[3178];
assign g[7273] = b[11] & g[3178];
assign g[5227] = a[11] & g[3179];
assign g[7274] = b[11] & g[3179];
assign g[5228] = a[11] & g[3180];
assign g[7275] = b[11] & g[3180];
assign g[5229] = a[11] & g[3181];
assign g[7276] = b[11] & g[3181];
assign g[5230] = a[11] & g[3182];
assign g[7277] = b[11] & g[3182];
assign g[5231] = a[11] & g[3183];
assign g[7278] = b[11] & g[3183];
assign g[5232] = a[11] & g[3184];
assign g[7279] = b[11] & g[3184];
assign g[5233] = a[11] & g[3185];
assign g[7280] = b[11] & g[3185];
assign g[5234] = a[11] & g[3186];
assign g[7281] = b[11] & g[3186];
assign g[5235] = a[11] & g[3187];
assign g[7282] = b[11] & g[3187];
assign g[5236] = a[11] & g[3188];
assign g[7283] = b[11] & g[3188];
assign g[5237] = a[11] & g[3189];
assign g[7284] = b[11] & g[3189];
assign g[5238] = a[11] & g[3190];
assign g[7285] = b[11] & g[3190];
assign g[5239] = a[11] & g[3191];
assign g[7286] = b[11] & g[3191];
assign g[5240] = a[11] & g[3192];
assign g[7287] = b[11] & g[3192];
assign g[5241] = a[11] & g[3193];
assign g[7288] = b[11] & g[3193];
assign g[5242] = a[11] & g[3194];
assign g[7289] = b[11] & g[3194];
assign g[5243] = a[11] & g[3195];
assign g[7290] = b[11] & g[3195];
assign g[5244] = a[11] & g[3196];
assign g[7291] = b[11] & g[3196];
assign g[5245] = a[11] & g[3197];
assign g[7292] = b[11] & g[3197];
assign g[5246] = a[11] & g[3198];
assign g[7293] = b[11] & g[3198];
assign g[5247] = a[11] & g[3199];
assign g[7294] = b[11] & g[3199];
assign g[5248] = a[11] & g[3200];
assign g[7295] = b[11] & g[3200];
assign g[5249] = a[11] & g[3201];
assign g[7296] = b[11] & g[3201];
assign g[5250] = a[11] & g[3202];
assign g[7297] = b[11] & g[3202];
assign g[5251] = a[11] & g[3203];
assign g[7298] = b[11] & g[3203];
assign g[5252] = a[11] & g[3204];
assign g[7299] = b[11] & g[3204];
assign g[5253] = a[11] & g[3205];
assign g[7300] = b[11] & g[3205];
assign g[5254] = a[11] & g[3206];
assign g[7301] = b[11] & g[3206];
assign g[5255] = a[11] & g[3207];
assign g[7302] = b[11] & g[3207];
assign g[5256] = a[11] & g[3208];
assign g[7303] = b[11] & g[3208];
assign g[5257] = a[11] & g[3209];
assign g[7304] = b[11] & g[3209];
assign g[5258] = a[11] & g[3210];
assign g[7305] = b[11] & g[3210];
assign g[5259] = a[11] & g[3211];
assign g[7306] = b[11] & g[3211];
assign g[5260] = a[11] & g[3212];
assign g[7307] = b[11] & g[3212];
assign g[5261] = a[11] & g[3213];
assign g[7308] = b[11] & g[3213];
assign g[5262] = a[11] & g[3214];
assign g[7309] = b[11] & g[3214];
assign g[5263] = a[11] & g[3215];
assign g[7310] = b[11] & g[3215];
assign g[5264] = a[11] & g[3216];
assign g[7311] = b[11] & g[3216];
assign g[5265] = a[11] & g[3217];
assign g[7312] = b[11] & g[3217];
assign g[5266] = a[11] & g[3218];
assign g[7313] = b[11] & g[3218];
assign g[5267] = a[11] & g[3219];
assign g[7314] = b[11] & g[3219];
assign g[5268] = a[11] & g[3220];
assign g[7315] = b[11] & g[3220];
assign g[5269] = a[11] & g[3221];
assign g[7316] = b[11] & g[3221];
assign g[5270] = a[11] & g[3222];
assign g[7317] = b[11] & g[3222];
assign g[5271] = a[11] & g[3223];
assign g[7318] = b[11] & g[3223];
assign g[5272] = a[11] & g[3224];
assign g[7319] = b[11] & g[3224];
assign g[5273] = a[11] & g[3225];
assign g[7320] = b[11] & g[3225];
assign g[5274] = a[11] & g[3226];
assign g[7321] = b[11] & g[3226];
assign g[5275] = a[11] & g[3227];
assign g[7322] = b[11] & g[3227];
assign g[5276] = a[11] & g[3228];
assign g[7323] = b[11] & g[3228];
assign g[5277] = a[11] & g[3229];
assign g[7324] = b[11] & g[3229];
assign g[5278] = a[11] & g[3230];
assign g[7325] = b[11] & g[3230];
assign g[5279] = a[11] & g[3231];
assign g[7326] = b[11] & g[3231];
assign g[5280] = a[11] & g[3232];
assign g[7327] = b[11] & g[3232];
assign g[5281] = a[11] & g[3233];
assign g[7328] = b[11] & g[3233];
assign g[5282] = a[11] & g[3234];
assign g[7329] = b[11] & g[3234];
assign g[5283] = a[11] & g[3235];
assign g[7330] = b[11] & g[3235];
assign g[5284] = a[11] & g[3236];
assign g[7331] = b[11] & g[3236];
assign g[5285] = a[11] & g[3237];
assign g[7332] = b[11] & g[3237];
assign g[5286] = a[11] & g[3238];
assign g[7333] = b[11] & g[3238];
assign g[5287] = a[11] & g[3239];
assign g[7334] = b[11] & g[3239];
assign g[5288] = a[11] & g[3240];
assign g[7335] = b[11] & g[3240];
assign g[5289] = a[11] & g[3241];
assign g[7336] = b[11] & g[3241];
assign g[5290] = a[11] & g[3242];
assign g[7337] = b[11] & g[3242];
assign g[5291] = a[11] & g[3243];
assign g[7338] = b[11] & g[3243];
assign g[5292] = a[11] & g[3244];
assign g[7339] = b[11] & g[3244];
assign g[5293] = a[11] & g[3245];
assign g[7340] = b[11] & g[3245];
assign g[5294] = a[11] & g[3246];
assign g[7341] = b[11] & g[3246];
assign g[5295] = a[11] & g[3247];
assign g[7342] = b[11] & g[3247];
assign g[5296] = a[11] & g[3248];
assign g[7343] = b[11] & g[3248];
assign g[5297] = a[11] & g[3249];
assign g[7344] = b[11] & g[3249];
assign g[5298] = a[11] & g[3250];
assign g[7345] = b[11] & g[3250];
assign g[5299] = a[11] & g[3251];
assign g[7346] = b[11] & g[3251];
assign g[5300] = a[11] & g[3252];
assign g[7347] = b[11] & g[3252];
assign g[5301] = a[11] & g[3253];
assign g[7348] = b[11] & g[3253];
assign g[5302] = a[11] & g[3254];
assign g[7349] = b[11] & g[3254];
assign g[5303] = a[11] & g[3255];
assign g[7350] = b[11] & g[3255];
assign g[5304] = a[11] & g[3256];
assign g[7351] = b[11] & g[3256];
assign g[5305] = a[11] & g[3257];
assign g[7352] = b[11] & g[3257];
assign g[5306] = a[11] & g[3258];
assign g[7353] = b[11] & g[3258];
assign g[5307] = a[11] & g[3259];
assign g[7354] = b[11] & g[3259];
assign g[5308] = a[11] & g[3260];
assign g[7355] = b[11] & g[3260];
assign g[5309] = a[11] & g[3261];
assign g[7356] = b[11] & g[3261];
assign g[5310] = a[11] & g[3262];
assign g[7357] = b[11] & g[3262];
assign g[5311] = a[11] & g[3263];
assign g[7358] = b[11] & g[3263];
assign g[5312] = a[11] & g[3264];
assign g[7359] = b[11] & g[3264];
assign g[5313] = a[11] & g[3265];
assign g[7360] = b[11] & g[3265];
assign g[5314] = a[11] & g[3266];
assign g[7361] = b[11] & g[3266];
assign g[5315] = a[11] & g[3267];
assign g[7362] = b[11] & g[3267];
assign g[5316] = a[11] & g[3268];
assign g[7363] = b[11] & g[3268];
assign g[5317] = a[11] & g[3269];
assign g[7364] = b[11] & g[3269];
assign g[5318] = a[11] & g[3270];
assign g[7365] = b[11] & g[3270];
assign g[5319] = a[11] & g[3271];
assign g[7366] = b[11] & g[3271];
assign g[5320] = a[11] & g[3272];
assign g[7367] = b[11] & g[3272];
assign g[5321] = a[11] & g[3273];
assign g[7368] = b[11] & g[3273];
assign g[5322] = a[11] & g[3274];
assign g[7369] = b[11] & g[3274];
assign g[5323] = a[11] & g[3275];
assign g[7370] = b[11] & g[3275];
assign g[5324] = a[11] & g[3276];
assign g[7371] = b[11] & g[3276];
assign g[5325] = a[11] & g[3277];
assign g[7372] = b[11] & g[3277];
assign g[5326] = a[11] & g[3278];
assign g[7373] = b[11] & g[3278];
assign g[5327] = a[11] & g[3279];
assign g[7374] = b[11] & g[3279];
assign g[5328] = a[11] & g[3280];
assign g[7375] = b[11] & g[3280];
assign g[5329] = a[11] & g[3281];
assign g[7376] = b[11] & g[3281];
assign g[5330] = a[11] & g[3282];
assign g[7377] = b[11] & g[3282];
assign g[5331] = a[11] & g[3283];
assign g[7378] = b[11] & g[3283];
assign g[5332] = a[11] & g[3284];
assign g[7379] = b[11] & g[3284];
assign g[5333] = a[11] & g[3285];
assign g[7380] = b[11] & g[3285];
assign g[5334] = a[11] & g[3286];
assign g[7381] = b[11] & g[3286];
assign g[5335] = a[11] & g[3287];
assign g[7382] = b[11] & g[3287];
assign g[5336] = a[11] & g[3288];
assign g[7383] = b[11] & g[3288];
assign g[5337] = a[11] & g[3289];
assign g[7384] = b[11] & g[3289];
assign g[5338] = a[11] & g[3290];
assign g[7385] = b[11] & g[3290];
assign g[5339] = a[11] & g[3291];
assign g[7386] = b[11] & g[3291];
assign g[5340] = a[11] & g[3292];
assign g[7387] = b[11] & g[3292];
assign g[5341] = a[11] & g[3293];
assign g[7388] = b[11] & g[3293];
assign g[5342] = a[11] & g[3294];
assign g[7389] = b[11] & g[3294];
assign g[5343] = a[11] & g[3295];
assign g[7390] = b[11] & g[3295];
assign g[5344] = a[11] & g[3296];
assign g[7391] = b[11] & g[3296];
assign g[5345] = a[11] & g[3297];
assign g[7392] = b[11] & g[3297];
assign g[5346] = a[11] & g[3298];
assign g[7393] = b[11] & g[3298];
assign g[5347] = a[11] & g[3299];
assign g[7394] = b[11] & g[3299];
assign g[5348] = a[11] & g[3300];
assign g[7395] = b[11] & g[3300];
assign g[5349] = a[11] & g[3301];
assign g[7396] = b[11] & g[3301];
assign g[5350] = a[11] & g[3302];
assign g[7397] = b[11] & g[3302];
assign g[5351] = a[11] & g[3303];
assign g[7398] = b[11] & g[3303];
assign g[5352] = a[11] & g[3304];
assign g[7399] = b[11] & g[3304];
assign g[5353] = a[11] & g[3305];
assign g[7400] = b[11] & g[3305];
assign g[5354] = a[11] & g[3306];
assign g[7401] = b[11] & g[3306];
assign g[5355] = a[11] & g[3307];
assign g[7402] = b[11] & g[3307];
assign g[5356] = a[11] & g[3308];
assign g[7403] = b[11] & g[3308];
assign g[5357] = a[11] & g[3309];
assign g[7404] = b[11] & g[3309];
assign g[5358] = a[11] & g[3310];
assign g[7405] = b[11] & g[3310];
assign g[5359] = a[11] & g[3311];
assign g[7406] = b[11] & g[3311];
assign g[5360] = a[11] & g[3312];
assign g[7407] = b[11] & g[3312];
assign g[5361] = a[11] & g[3313];
assign g[7408] = b[11] & g[3313];
assign g[5362] = a[11] & g[3314];
assign g[7409] = b[11] & g[3314];
assign g[5363] = a[11] & g[3315];
assign g[7410] = b[11] & g[3315];
assign g[5364] = a[11] & g[3316];
assign g[7411] = b[11] & g[3316];
assign g[5365] = a[11] & g[3317];
assign g[7412] = b[11] & g[3317];
assign g[5366] = a[11] & g[3318];
assign g[7413] = b[11] & g[3318];
assign g[5367] = a[11] & g[3319];
assign g[7414] = b[11] & g[3319];
assign g[5368] = a[11] & g[3320];
assign g[7415] = b[11] & g[3320];
assign g[5369] = a[11] & g[3321];
assign g[7416] = b[11] & g[3321];
assign g[5370] = a[11] & g[3322];
assign g[7417] = b[11] & g[3322];
assign g[5371] = a[11] & g[3323];
assign g[7418] = b[11] & g[3323];
assign g[5372] = a[11] & g[3324];
assign g[7419] = b[11] & g[3324];
assign g[5373] = a[11] & g[3325];
assign g[7420] = b[11] & g[3325];
assign g[5374] = a[11] & g[3326];
assign g[7421] = b[11] & g[3326];
assign g[5375] = a[11] & g[3327];
assign g[7422] = b[11] & g[3327];
assign g[5376] = a[11] & g[3328];
assign g[7423] = b[11] & g[3328];
assign g[5377] = a[11] & g[3329];
assign g[7424] = b[11] & g[3329];
assign g[5378] = a[11] & g[3330];
assign g[7425] = b[11] & g[3330];
assign g[5379] = a[11] & g[3331];
assign g[7426] = b[11] & g[3331];
assign g[5380] = a[11] & g[3332];
assign g[7427] = b[11] & g[3332];
assign g[5381] = a[11] & g[3333];
assign g[7428] = b[11] & g[3333];
assign g[5382] = a[11] & g[3334];
assign g[7429] = b[11] & g[3334];
assign g[5383] = a[11] & g[3335];
assign g[7430] = b[11] & g[3335];
assign g[5384] = a[11] & g[3336];
assign g[7431] = b[11] & g[3336];
assign g[5385] = a[11] & g[3337];
assign g[7432] = b[11] & g[3337];
assign g[5386] = a[11] & g[3338];
assign g[7433] = b[11] & g[3338];
assign g[5387] = a[11] & g[3339];
assign g[7434] = b[11] & g[3339];
assign g[5388] = a[11] & g[3340];
assign g[7435] = b[11] & g[3340];
assign g[5389] = a[11] & g[3341];
assign g[7436] = b[11] & g[3341];
assign g[5390] = a[11] & g[3342];
assign g[7437] = b[11] & g[3342];
assign g[5391] = a[11] & g[3343];
assign g[7438] = b[11] & g[3343];
assign g[5392] = a[11] & g[3344];
assign g[7439] = b[11] & g[3344];
assign g[5393] = a[11] & g[3345];
assign g[7440] = b[11] & g[3345];
assign g[5394] = a[11] & g[3346];
assign g[7441] = b[11] & g[3346];
assign g[5395] = a[11] & g[3347];
assign g[7442] = b[11] & g[3347];
assign g[5396] = a[11] & g[3348];
assign g[7443] = b[11] & g[3348];
assign g[5397] = a[11] & g[3349];
assign g[7444] = b[11] & g[3349];
assign g[5398] = a[11] & g[3350];
assign g[7445] = b[11] & g[3350];
assign g[5399] = a[11] & g[3351];
assign g[7446] = b[11] & g[3351];
assign g[5400] = a[11] & g[3352];
assign g[7447] = b[11] & g[3352];
assign g[5401] = a[11] & g[3353];
assign g[7448] = b[11] & g[3353];
assign g[5402] = a[11] & g[3354];
assign g[7449] = b[11] & g[3354];
assign g[5403] = a[11] & g[3355];
assign g[7450] = b[11] & g[3355];
assign g[5404] = a[11] & g[3356];
assign g[7451] = b[11] & g[3356];
assign g[5405] = a[11] & g[3357];
assign g[7452] = b[11] & g[3357];
assign g[5406] = a[11] & g[3358];
assign g[7453] = b[11] & g[3358];
assign g[5407] = a[11] & g[3359];
assign g[7454] = b[11] & g[3359];
assign g[5408] = a[11] & g[3360];
assign g[7455] = b[11] & g[3360];
assign g[5409] = a[11] & g[3361];
assign g[7456] = b[11] & g[3361];
assign g[5410] = a[11] & g[3362];
assign g[7457] = b[11] & g[3362];
assign g[5411] = a[11] & g[3363];
assign g[7458] = b[11] & g[3363];
assign g[5412] = a[11] & g[3364];
assign g[7459] = b[11] & g[3364];
assign g[5413] = a[11] & g[3365];
assign g[7460] = b[11] & g[3365];
assign g[5414] = a[11] & g[3366];
assign g[7461] = b[11] & g[3366];
assign g[5415] = a[11] & g[3367];
assign g[7462] = b[11] & g[3367];
assign g[5416] = a[11] & g[3368];
assign g[7463] = b[11] & g[3368];
assign g[5417] = a[11] & g[3369];
assign g[7464] = b[11] & g[3369];
assign g[5418] = a[11] & g[3370];
assign g[7465] = b[11] & g[3370];
assign g[5419] = a[11] & g[3371];
assign g[7466] = b[11] & g[3371];
assign g[5420] = a[11] & g[3372];
assign g[7467] = b[11] & g[3372];
assign g[5421] = a[11] & g[3373];
assign g[7468] = b[11] & g[3373];
assign g[5422] = a[11] & g[3374];
assign g[7469] = b[11] & g[3374];
assign g[5423] = a[11] & g[3375];
assign g[7470] = b[11] & g[3375];
assign g[5424] = a[11] & g[3376];
assign g[7471] = b[11] & g[3376];
assign g[5425] = a[11] & g[3377];
assign g[7472] = b[11] & g[3377];
assign g[5426] = a[11] & g[3378];
assign g[7473] = b[11] & g[3378];
assign g[5427] = a[11] & g[3379];
assign g[7474] = b[11] & g[3379];
assign g[5428] = a[11] & g[3380];
assign g[7475] = b[11] & g[3380];
assign g[5429] = a[11] & g[3381];
assign g[7476] = b[11] & g[3381];
assign g[5430] = a[11] & g[3382];
assign g[7477] = b[11] & g[3382];
assign g[5431] = a[11] & g[3383];
assign g[7478] = b[11] & g[3383];
assign g[5432] = a[11] & g[3384];
assign g[7479] = b[11] & g[3384];
assign g[5433] = a[11] & g[3385];
assign g[7480] = b[11] & g[3385];
assign g[5434] = a[11] & g[3386];
assign g[7481] = b[11] & g[3386];
assign g[5435] = a[11] & g[3387];
assign g[7482] = b[11] & g[3387];
assign g[5436] = a[11] & g[3388];
assign g[7483] = b[11] & g[3388];
assign g[5437] = a[11] & g[3389];
assign g[7484] = b[11] & g[3389];
assign g[5438] = a[11] & g[3390];
assign g[7485] = b[11] & g[3390];
assign g[5439] = a[11] & g[3391];
assign g[7486] = b[11] & g[3391];
assign g[5440] = a[11] & g[3392];
assign g[7487] = b[11] & g[3392];
assign g[5441] = a[11] & g[3393];
assign g[7488] = b[11] & g[3393];
assign g[5442] = a[11] & g[3394];
assign g[7489] = b[11] & g[3394];
assign g[5443] = a[11] & g[3395];
assign g[7490] = b[11] & g[3395];
assign g[5444] = a[11] & g[3396];
assign g[7491] = b[11] & g[3396];
assign g[5445] = a[11] & g[3397];
assign g[7492] = b[11] & g[3397];
assign g[5446] = a[11] & g[3398];
assign g[7493] = b[11] & g[3398];
assign g[5447] = a[11] & g[3399];
assign g[7494] = b[11] & g[3399];
assign g[5448] = a[11] & g[3400];
assign g[7495] = b[11] & g[3400];
assign g[5449] = a[11] & g[3401];
assign g[7496] = b[11] & g[3401];
assign g[5450] = a[11] & g[3402];
assign g[7497] = b[11] & g[3402];
assign g[5451] = a[11] & g[3403];
assign g[7498] = b[11] & g[3403];
assign g[5452] = a[11] & g[3404];
assign g[7499] = b[11] & g[3404];
assign g[5453] = a[11] & g[3405];
assign g[7500] = b[11] & g[3405];
assign g[5454] = a[11] & g[3406];
assign g[7501] = b[11] & g[3406];
assign g[5455] = a[11] & g[3407];
assign g[7502] = b[11] & g[3407];
assign g[5456] = a[11] & g[3408];
assign g[7503] = b[11] & g[3408];
assign g[5457] = a[11] & g[3409];
assign g[7504] = b[11] & g[3409];
assign g[5458] = a[11] & g[3410];
assign g[7505] = b[11] & g[3410];
assign g[5459] = a[11] & g[3411];
assign g[7506] = b[11] & g[3411];
assign g[5460] = a[11] & g[3412];
assign g[7507] = b[11] & g[3412];
assign g[5461] = a[11] & g[3413];
assign g[7508] = b[11] & g[3413];
assign g[5462] = a[11] & g[3414];
assign g[7509] = b[11] & g[3414];
assign g[5463] = a[11] & g[3415];
assign g[7510] = b[11] & g[3415];
assign g[5464] = a[11] & g[3416];
assign g[7511] = b[11] & g[3416];
assign g[5465] = a[11] & g[3417];
assign g[7512] = b[11] & g[3417];
assign g[5466] = a[11] & g[3418];
assign g[7513] = b[11] & g[3418];
assign g[5467] = a[11] & g[3419];
assign g[7514] = b[11] & g[3419];
assign g[5468] = a[11] & g[3420];
assign g[7515] = b[11] & g[3420];
assign g[5469] = a[11] & g[3421];
assign g[7516] = b[11] & g[3421];
assign g[5470] = a[11] & g[3422];
assign g[7517] = b[11] & g[3422];
assign g[5471] = a[11] & g[3423];
assign g[7518] = b[11] & g[3423];
assign g[5472] = a[11] & g[3424];
assign g[7519] = b[11] & g[3424];
assign g[5473] = a[11] & g[3425];
assign g[7520] = b[11] & g[3425];
assign g[5474] = a[11] & g[3426];
assign g[7521] = b[11] & g[3426];
assign g[5475] = a[11] & g[3427];
assign g[7522] = b[11] & g[3427];
assign g[5476] = a[11] & g[3428];
assign g[7523] = b[11] & g[3428];
assign g[5477] = a[11] & g[3429];
assign g[7524] = b[11] & g[3429];
assign g[5478] = a[11] & g[3430];
assign g[7525] = b[11] & g[3430];
assign g[5479] = a[11] & g[3431];
assign g[7526] = b[11] & g[3431];
assign g[5480] = a[11] & g[3432];
assign g[7527] = b[11] & g[3432];
assign g[5481] = a[11] & g[3433];
assign g[7528] = b[11] & g[3433];
assign g[5482] = a[11] & g[3434];
assign g[7529] = b[11] & g[3434];
assign g[5483] = a[11] & g[3435];
assign g[7530] = b[11] & g[3435];
assign g[5484] = a[11] & g[3436];
assign g[7531] = b[11] & g[3436];
assign g[5485] = a[11] & g[3437];
assign g[7532] = b[11] & g[3437];
assign g[5486] = a[11] & g[3438];
assign g[7533] = b[11] & g[3438];
assign g[5487] = a[11] & g[3439];
assign g[7534] = b[11] & g[3439];
assign g[5488] = a[11] & g[3440];
assign g[7535] = b[11] & g[3440];
assign g[5489] = a[11] & g[3441];
assign g[7536] = b[11] & g[3441];
assign g[5490] = a[11] & g[3442];
assign g[7537] = b[11] & g[3442];
assign g[5491] = a[11] & g[3443];
assign g[7538] = b[11] & g[3443];
assign g[5492] = a[11] & g[3444];
assign g[7539] = b[11] & g[3444];
assign g[5493] = a[11] & g[3445];
assign g[7540] = b[11] & g[3445];
assign g[5494] = a[11] & g[3446];
assign g[7541] = b[11] & g[3446];
assign g[5495] = a[11] & g[3447];
assign g[7542] = b[11] & g[3447];
assign g[5496] = a[11] & g[3448];
assign g[7543] = b[11] & g[3448];
assign g[5497] = a[11] & g[3449];
assign g[7544] = b[11] & g[3449];
assign g[5498] = a[11] & g[3450];
assign g[7545] = b[11] & g[3450];
assign g[5499] = a[11] & g[3451];
assign g[7546] = b[11] & g[3451];
assign g[5500] = a[11] & g[3452];
assign g[7547] = b[11] & g[3452];
assign g[5501] = a[11] & g[3453];
assign g[7548] = b[11] & g[3453];
assign g[5502] = a[11] & g[3454];
assign g[7549] = b[11] & g[3454];
assign g[5503] = a[11] & g[3455];
assign g[7550] = b[11] & g[3455];
assign g[5504] = a[11] & g[3456];
assign g[7551] = b[11] & g[3456];
assign g[5505] = a[11] & g[3457];
assign g[7552] = b[11] & g[3457];
assign g[5506] = a[11] & g[3458];
assign g[7553] = b[11] & g[3458];
assign g[5507] = a[11] & g[3459];
assign g[7554] = b[11] & g[3459];
assign g[5508] = a[11] & g[3460];
assign g[7555] = b[11] & g[3460];
assign g[5509] = a[11] & g[3461];
assign g[7556] = b[11] & g[3461];
assign g[5510] = a[11] & g[3462];
assign g[7557] = b[11] & g[3462];
assign g[5511] = a[11] & g[3463];
assign g[7558] = b[11] & g[3463];
assign g[5512] = a[11] & g[3464];
assign g[7559] = b[11] & g[3464];
assign g[5513] = a[11] & g[3465];
assign g[7560] = b[11] & g[3465];
assign g[5514] = a[11] & g[3466];
assign g[7561] = b[11] & g[3466];
assign g[5515] = a[11] & g[3467];
assign g[7562] = b[11] & g[3467];
assign g[5516] = a[11] & g[3468];
assign g[7563] = b[11] & g[3468];
assign g[5517] = a[11] & g[3469];
assign g[7564] = b[11] & g[3469];
assign g[5518] = a[11] & g[3470];
assign g[7565] = b[11] & g[3470];
assign g[5519] = a[11] & g[3471];
assign g[7566] = b[11] & g[3471];
assign g[5520] = a[11] & g[3472];
assign g[7567] = b[11] & g[3472];
assign g[5521] = a[11] & g[3473];
assign g[7568] = b[11] & g[3473];
assign g[5522] = a[11] & g[3474];
assign g[7569] = b[11] & g[3474];
assign g[5523] = a[11] & g[3475];
assign g[7570] = b[11] & g[3475];
assign g[5524] = a[11] & g[3476];
assign g[7571] = b[11] & g[3476];
assign g[5525] = a[11] & g[3477];
assign g[7572] = b[11] & g[3477];
assign g[5526] = a[11] & g[3478];
assign g[7573] = b[11] & g[3478];
assign g[5527] = a[11] & g[3479];
assign g[7574] = b[11] & g[3479];
assign g[5528] = a[11] & g[3480];
assign g[7575] = b[11] & g[3480];
assign g[5529] = a[11] & g[3481];
assign g[7576] = b[11] & g[3481];
assign g[5530] = a[11] & g[3482];
assign g[7577] = b[11] & g[3482];
assign g[5531] = a[11] & g[3483];
assign g[7578] = b[11] & g[3483];
assign g[5532] = a[11] & g[3484];
assign g[7579] = b[11] & g[3484];
assign g[5533] = a[11] & g[3485];
assign g[7580] = b[11] & g[3485];
assign g[5534] = a[11] & g[3486];
assign g[7581] = b[11] & g[3486];
assign g[5535] = a[11] & g[3487];
assign g[7582] = b[11] & g[3487];
assign g[5536] = a[11] & g[3488];
assign g[7583] = b[11] & g[3488];
assign g[5537] = a[11] & g[3489];
assign g[7584] = b[11] & g[3489];
assign g[5538] = a[11] & g[3490];
assign g[7585] = b[11] & g[3490];
assign g[5539] = a[11] & g[3491];
assign g[7586] = b[11] & g[3491];
assign g[5540] = a[11] & g[3492];
assign g[7587] = b[11] & g[3492];
assign g[5541] = a[11] & g[3493];
assign g[7588] = b[11] & g[3493];
assign g[5542] = a[11] & g[3494];
assign g[7589] = b[11] & g[3494];
assign g[5543] = a[11] & g[3495];
assign g[7590] = b[11] & g[3495];
assign g[5544] = a[11] & g[3496];
assign g[7591] = b[11] & g[3496];
assign g[5545] = a[11] & g[3497];
assign g[7592] = b[11] & g[3497];
assign g[5546] = a[11] & g[3498];
assign g[7593] = b[11] & g[3498];
assign g[5547] = a[11] & g[3499];
assign g[7594] = b[11] & g[3499];
assign g[5548] = a[11] & g[3500];
assign g[7595] = b[11] & g[3500];
assign g[5549] = a[11] & g[3501];
assign g[7596] = b[11] & g[3501];
assign g[5550] = a[11] & g[3502];
assign g[7597] = b[11] & g[3502];
assign g[5551] = a[11] & g[3503];
assign g[7598] = b[11] & g[3503];
assign g[5552] = a[11] & g[3504];
assign g[7599] = b[11] & g[3504];
assign g[5553] = a[11] & g[3505];
assign g[7600] = b[11] & g[3505];
assign g[5554] = a[11] & g[3506];
assign g[7601] = b[11] & g[3506];
assign g[5555] = a[11] & g[3507];
assign g[7602] = b[11] & g[3507];
assign g[5556] = a[11] & g[3508];
assign g[7603] = b[11] & g[3508];
assign g[5557] = a[11] & g[3509];
assign g[7604] = b[11] & g[3509];
assign g[5558] = a[11] & g[3510];
assign g[7605] = b[11] & g[3510];
assign g[5559] = a[11] & g[3511];
assign g[7606] = b[11] & g[3511];
assign g[5560] = a[11] & g[3512];
assign g[7607] = b[11] & g[3512];
assign g[5561] = a[11] & g[3513];
assign g[7608] = b[11] & g[3513];
assign g[5562] = a[11] & g[3514];
assign g[7609] = b[11] & g[3514];
assign g[5563] = a[11] & g[3515];
assign g[7610] = b[11] & g[3515];
assign g[5564] = a[11] & g[3516];
assign g[7611] = b[11] & g[3516];
assign g[5565] = a[11] & g[3517];
assign g[7612] = b[11] & g[3517];
assign g[5566] = a[11] & g[3518];
assign g[7613] = b[11] & g[3518];
assign g[5567] = a[11] & g[3519];
assign g[7614] = b[11] & g[3519];
assign g[5568] = a[11] & g[3520];
assign g[7615] = b[11] & g[3520];
assign g[5569] = a[11] & g[3521];
assign g[7616] = b[11] & g[3521];
assign g[5570] = a[11] & g[3522];
assign g[7617] = b[11] & g[3522];
assign g[5571] = a[11] & g[3523];
assign g[7618] = b[11] & g[3523];
assign g[5572] = a[11] & g[3524];
assign g[7619] = b[11] & g[3524];
assign g[5573] = a[11] & g[3525];
assign g[7620] = b[11] & g[3525];
assign g[5574] = a[11] & g[3526];
assign g[7621] = b[11] & g[3526];
assign g[5575] = a[11] & g[3527];
assign g[7622] = b[11] & g[3527];
assign g[5576] = a[11] & g[3528];
assign g[7623] = b[11] & g[3528];
assign g[5577] = a[11] & g[3529];
assign g[7624] = b[11] & g[3529];
assign g[5578] = a[11] & g[3530];
assign g[7625] = b[11] & g[3530];
assign g[5579] = a[11] & g[3531];
assign g[7626] = b[11] & g[3531];
assign g[5580] = a[11] & g[3532];
assign g[7627] = b[11] & g[3532];
assign g[5581] = a[11] & g[3533];
assign g[7628] = b[11] & g[3533];
assign g[5582] = a[11] & g[3534];
assign g[7629] = b[11] & g[3534];
assign g[5583] = a[11] & g[3535];
assign g[7630] = b[11] & g[3535];
assign g[5584] = a[11] & g[3536];
assign g[7631] = b[11] & g[3536];
assign g[5585] = a[11] & g[3537];
assign g[7632] = b[11] & g[3537];
assign g[5586] = a[11] & g[3538];
assign g[7633] = b[11] & g[3538];
assign g[5587] = a[11] & g[3539];
assign g[7634] = b[11] & g[3539];
assign g[5588] = a[11] & g[3540];
assign g[7635] = b[11] & g[3540];
assign g[5589] = a[11] & g[3541];
assign g[7636] = b[11] & g[3541];
assign g[5590] = a[11] & g[3542];
assign g[7637] = b[11] & g[3542];
assign g[5591] = a[11] & g[3543];
assign g[7638] = b[11] & g[3543];
assign g[5592] = a[11] & g[3544];
assign g[7639] = b[11] & g[3544];
assign g[5593] = a[11] & g[3545];
assign g[7640] = b[11] & g[3545];
assign g[5594] = a[11] & g[3546];
assign g[7641] = b[11] & g[3546];
assign g[5595] = a[11] & g[3547];
assign g[7642] = b[11] & g[3547];
assign g[5596] = a[11] & g[3548];
assign g[7643] = b[11] & g[3548];
assign g[5597] = a[11] & g[3549];
assign g[7644] = b[11] & g[3549];
assign g[5598] = a[11] & g[3550];
assign g[7645] = b[11] & g[3550];
assign g[5599] = a[11] & g[3551];
assign g[7646] = b[11] & g[3551];
assign g[5600] = a[11] & g[3552];
assign g[7647] = b[11] & g[3552];
assign g[5601] = a[11] & g[3553];
assign g[7648] = b[11] & g[3553];
assign g[5602] = a[11] & g[3554];
assign g[7649] = b[11] & g[3554];
assign g[5603] = a[11] & g[3555];
assign g[7650] = b[11] & g[3555];
assign g[5604] = a[11] & g[3556];
assign g[7651] = b[11] & g[3556];
assign g[5605] = a[11] & g[3557];
assign g[7652] = b[11] & g[3557];
assign g[5606] = a[11] & g[3558];
assign g[7653] = b[11] & g[3558];
assign g[5607] = a[11] & g[3559];
assign g[7654] = b[11] & g[3559];
assign g[5608] = a[11] & g[3560];
assign g[7655] = b[11] & g[3560];
assign g[5609] = a[11] & g[3561];
assign g[7656] = b[11] & g[3561];
assign g[5610] = a[11] & g[3562];
assign g[7657] = b[11] & g[3562];
assign g[5611] = a[11] & g[3563];
assign g[7658] = b[11] & g[3563];
assign g[5612] = a[11] & g[3564];
assign g[7659] = b[11] & g[3564];
assign g[5613] = a[11] & g[3565];
assign g[7660] = b[11] & g[3565];
assign g[5614] = a[11] & g[3566];
assign g[7661] = b[11] & g[3566];
assign g[5615] = a[11] & g[3567];
assign g[7662] = b[11] & g[3567];
assign g[5616] = a[11] & g[3568];
assign g[7663] = b[11] & g[3568];
assign g[5617] = a[11] & g[3569];
assign g[7664] = b[11] & g[3569];
assign g[5618] = a[11] & g[3570];
assign g[7665] = b[11] & g[3570];
assign g[5619] = a[11] & g[3571];
assign g[7666] = b[11] & g[3571];
assign g[5620] = a[11] & g[3572];
assign g[7667] = b[11] & g[3572];
assign g[5621] = a[11] & g[3573];
assign g[7668] = b[11] & g[3573];
assign g[5622] = a[11] & g[3574];
assign g[7669] = b[11] & g[3574];
assign g[5623] = a[11] & g[3575];
assign g[7670] = b[11] & g[3575];
assign g[5624] = a[11] & g[3576];
assign g[7671] = b[11] & g[3576];
assign g[5625] = a[11] & g[3577];
assign g[7672] = b[11] & g[3577];
assign g[5626] = a[11] & g[3578];
assign g[7673] = b[11] & g[3578];
assign g[5627] = a[11] & g[3579];
assign g[7674] = b[11] & g[3579];
assign g[5628] = a[11] & g[3580];
assign g[7675] = b[11] & g[3580];
assign g[5629] = a[11] & g[3581];
assign g[7676] = b[11] & g[3581];
assign g[5630] = a[11] & g[3582];
assign g[7677] = b[11] & g[3582];
assign g[5631] = a[11] & g[3583];
assign g[7678] = b[11] & g[3583];
assign g[5632] = a[11] & g[3584];
assign g[7679] = b[11] & g[3584];
assign g[5633] = a[11] & g[3585];
assign g[7680] = b[11] & g[3585];
assign g[5634] = a[11] & g[3586];
assign g[7681] = b[11] & g[3586];
assign g[5635] = a[11] & g[3587];
assign g[7682] = b[11] & g[3587];
assign g[5636] = a[11] & g[3588];
assign g[7683] = b[11] & g[3588];
assign g[5637] = a[11] & g[3589];
assign g[7684] = b[11] & g[3589];
assign g[5638] = a[11] & g[3590];
assign g[7685] = b[11] & g[3590];
assign g[5639] = a[11] & g[3591];
assign g[7686] = b[11] & g[3591];
assign g[5640] = a[11] & g[3592];
assign g[7687] = b[11] & g[3592];
assign g[5641] = a[11] & g[3593];
assign g[7688] = b[11] & g[3593];
assign g[5642] = a[11] & g[3594];
assign g[7689] = b[11] & g[3594];
assign g[5643] = a[11] & g[3595];
assign g[7690] = b[11] & g[3595];
assign g[5644] = a[11] & g[3596];
assign g[7691] = b[11] & g[3596];
assign g[5645] = a[11] & g[3597];
assign g[7692] = b[11] & g[3597];
assign g[5646] = a[11] & g[3598];
assign g[7693] = b[11] & g[3598];
assign g[5647] = a[11] & g[3599];
assign g[7694] = b[11] & g[3599];
assign g[5648] = a[11] & g[3600];
assign g[7695] = b[11] & g[3600];
assign g[5649] = a[11] & g[3601];
assign g[7696] = b[11] & g[3601];
assign g[5650] = a[11] & g[3602];
assign g[7697] = b[11] & g[3602];
assign g[5651] = a[11] & g[3603];
assign g[7698] = b[11] & g[3603];
assign g[5652] = a[11] & g[3604];
assign g[7699] = b[11] & g[3604];
assign g[5653] = a[11] & g[3605];
assign g[7700] = b[11] & g[3605];
assign g[5654] = a[11] & g[3606];
assign g[7701] = b[11] & g[3606];
assign g[5655] = a[11] & g[3607];
assign g[7702] = b[11] & g[3607];
assign g[5656] = a[11] & g[3608];
assign g[7703] = b[11] & g[3608];
assign g[5657] = a[11] & g[3609];
assign g[7704] = b[11] & g[3609];
assign g[5658] = a[11] & g[3610];
assign g[7705] = b[11] & g[3610];
assign g[5659] = a[11] & g[3611];
assign g[7706] = b[11] & g[3611];
assign g[5660] = a[11] & g[3612];
assign g[7707] = b[11] & g[3612];
assign g[5661] = a[11] & g[3613];
assign g[7708] = b[11] & g[3613];
assign g[5662] = a[11] & g[3614];
assign g[7709] = b[11] & g[3614];
assign g[5663] = a[11] & g[3615];
assign g[7710] = b[11] & g[3615];
assign g[5664] = a[11] & g[3616];
assign g[7711] = b[11] & g[3616];
assign g[5665] = a[11] & g[3617];
assign g[7712] = b[11] & g[3617];
assign g[5666] = a[11] & g[3618];
assign g[7713] = b[11] & g[3618];
assign g[5667] = a[11] & g[3619];
assign g[7714] = b[11] & g[3619];
assign g[5668] = a[11] & g[3620];
assign g[7715] = b[11] & g[3620];
assign g[5669] = a[11] & g[3621];
assign g[7716] = b[11] & g[3621];
assign g[5670] = a[11] & g[3622];
assign g[7717] = b[11] & g[3622];
assign g[5671] = a[11] & g[3623];
assign g[7718] = b[11] & g[3623];
assign g[5672] = a[11] & g[3624];
assign g[7719] = b[11] & g[3624];
assign g[5673] = a[11] & g[3625];
assign g[7720] = b[11] & g[3625];
assign g[5674] = a[11] & g[3626];
assign g[7721] = b[11] & g[3626];
assign g[5675] = a[11] & g[3627];
assign g[7722] = b[11] & g[3627];
assign g[5676] = a[11] & g[3628];
assign g[7723] = b[11] & g[3628];
assign g[5677] = a[11] & g[3629];
assign g[7724] = b[11] & g[3629];
assign g[5678] = a[11] & g[3630];
assign g[7725] = b[11] & g[3630];
assign g[5679] = a[11] & g[3631];
assign g[7726] = b[11] & g[3631];
assign g[5680] = a[11] & g[3632];
assign g[7727] = b[11] & g[3632];
assign g[5681] = a[11] & g[3633];
assign g[7728] = b[11] & g[3633];
assign g[5682] = a[11] & g[3634];
assign g[7729] = b[11] & g[3634];
assign g[5683] = a[11] & g[3635];
assign g[7730] = b[11] & g[3635];
assign g[5684] = a[11] & g[3636];
assign g[7731] = b[11] & g[3636];
assign g[5685] = a[11] & g[3637];
assign g[7732] = b[11] & g[3637];
assign g[5686] = a[11] & g[3638];
assign g[7733] = b[11] & g[3638];
assign g[5687] = a[11] & g[3639];
assign g[7734] = b[11] & g[3639];
assign g[5688] = a[11] & g[3640];
assign g[7735] = b[11] & g[3640];
assign g[5689] = a[11] & g[3641];
assign g[7736] = b[11] & g[3641];
assign g[5690] = a[11] & g[3642];
assign g[7737] = b[11] & g[3642];
assign g[5691] = a[11] & g[3643];
assign g[7738] = b[11] & g[3643];
assign g[5692] = a[11] & g[3644];
assign g[7739] = b[11] & g[3644];
assign g[5693] = a[11] & g[3645];
assign g[7740] = b[11] & g[3645];
assign g[5694] = a[11] & g[3646];
assign g[7741] = b[11] & g[3646];
assign g[5695] = a[11] & g[3647];
assign g[7742] = b[11] & g[3647];
assign g[5696] = a[11] & g[3648];
assign g[7743] = b[11] & g[3648];
assign g[5697] = a[11] & g[3649];
assign g[7744] = b[11] & g[3649];
assign g[5698] = a[11] & g[3650];
assign g[7745] = b[11] & g[3650];
assign g[5699] = a[11] & g[3651];
assign g[7746] = b[11] & g[3651];
assign g[5700] = a[11] & g[3652];
assign g[7747] = b[11] & g[3652];
assign g[5701] = a[11] & g[3653];
assign g[7748] = b[11] & g[3653];
assign g[5702] = a[11] & g[3654];
assign g[7749] = b[11] & g[3654];
assign g[5703] = a[11] & g[3655];
assign g[7750] = b[11] & g[3655];
assign g[5704] = a[11] & g[3656];
assign g[7751] = b[11] & g[3656];
assign g[5705] = a[11] & g[3657];
assign g[7752] = b[11] & g[3657];
assign g[5706] = a[11] & g[3658];
assign g[7753] = b[11] & g[3658];
assign g[5707] = a[11] & g[3659];
assign g[7754] = b[11] & g[3659];
assign g[5708] = a[11] & g[3660];
assign g[7755] = b[11] & g[3660];
assign g[5709] = a[11] & g[3661];
assign g[7756] = b[11] & g[3661];
assign g[5710] = a[11] & g[3662];
assign g[7757] = b[11] & g[3662];
assign g[5711] = a[11] & g[3663];
assign g[7758] = b[11] & g[3663];
assign g[5712] = a[11] & g[3664];
assign g[7759] = b[11] & g[3664];
assign g[5713] = a[11] & g[3665];
assign g[7760] = b[11] & g[3665];
assign g[5714] = a[11] & g[3666];
assign g[7761] = b[11] & g[3666];
assign g[5715] = a[11] & g[3667];
assign g[7762] = b[11] & g[3667];
assign g[5716] = a[11] & g[3668];
assign g[7763] = b[11] & g[3668];
assign g[5717] = a[11] & g[3669];
assign g[7764] = b[11] & g[3669];
assign g[5718] = a[11] & g[3670];
assign g[7765] = b[11] & g[3670];
assign g[5719] = a[11] & g[3671];
assign g[7766] = b[11] & g[3671];
assign g[5720] = a[11] & g[3672];
assign g[7767] = b[11] & g[3672];
assign g[5721] = a[11] & g[3673];
assign g[7768] = b[11] & g[3673];
assign g[5722] = a[11] & g[3674];
assign g[7769] = b[11] & g[3674];
assign g[5723] = a[11] & g[3675];
assign g[7770] = b[11] & g[3675];
assign g[5724] = a[11] & g[3676];
assign g[7771] = b[11] & g[3676];
assign g[5725] = a[11] & g[3677];
assign g[7772] = b[11] & g[3677];
assign g[5726] = a[11] & g[3678];
assign g[7773] = b[11] & g[3678];
assign g[5727] = a[11] & g[3679];
assign g[7774] = b[11] & g[3679];
assign g[5728] = a[11] & g[3680];
assign g[7775] = b[11] & g[3680];
assign g[5729] = a[11] & g[3681];
assign g[7776] = b[11] & g[3681];
assign g[5730] = a[11] & g[3682];
assign g[7777] = b[11] & g[3682];
assign g[5731] = a[11] & g[3683];
assign g[7778] = b[11] & g[3683];
assign g[5732] = a[11] & g[3684];
assign g[7779] = b[11] & g[3684];
assign g[5733] = a[11] & g[3685];
assign g[7780] = b[11] & g[3685];
assign g[5734] = a[11] & g[3686];
assign g[7781] = b[11] & g[3686];
assign g[5735] = a[11] & g[3687];
assign g[7782] = b[11] & g[3687];
assign g[5736] = a[11] & g[3688];
assign g[7783] = b[11] & g[3688];
assign g[5737] = a[11] & g[3689];
assign g[7784] = b[11] & g[3689];
assign g[5738] = a[11] & g[3690];
assign g[7785] = b[11] & g[3690];
assign g[5739] = a[11] & g[3691];
assign g[7786] = b[11] & g[3691];
assign g[5740] = a[11] & g[3692];
assign g[7787] = b[11] & g[3692];
assign g[5741] = a[11] & g[3693];
assign g[7788] = b[11] & g[3693];
assign g[5742] = a[11] & g[3694];
assign g[7789] = b[11] & g[3694];
assign g[5743] = a[11] & g[3695];
assign g[7790] = b[11] & g[3695];
assign g[5744] = a[11] & g[3696];
assign g[7791] = b[11] & g[3696];
assign g[5745] = a[11] & g[3697];
assign g[7792] = b[11] & g[3697];
assign g[5746] = a[11] & g[3698];
assign g[7793] = b[11] & g[3698];
assign g[5747] = a[11] & g[3699];
assign g[7794] = b[11] & g[3699];
assign g[5748] = a[11] & g[3700];
assign g[7795] = b[11] & g[3700];
assign g[5749] = a[11] & g[3701];
assign g[7796] = b[11] & g[3701];
assign g[5750] = a[11] & g[3702];
assign g[7797] = b[11] & g[3702];
assign g[5751] = a[11] & g[3703];
assign g[7798] = b[11] & g[3703];
assign g[5752] = a[11] & g[3704];
assign g[7799] = b[11] & g[3704];
assign g[5753] = a[11] & g[3705];
assign g[7800] = b[11] & g[3705];
assign g[5754] = a[11] & g[3706];
assign g[7801] = b[11] & g[3706];
assign g[5755] = a[11] & g[3707];
assign g[7802] = b[11] & g[3707];
assign g[5756] = a[11] & g[3708];
assign g[7803] = b[11] & g[3708];
assign g[5757] = a[11] & g[3709];
assign g[7804] = b[11] & g[3709];
assign g[5758] = a[11] & g[3710];
assign g[7805] = b[11] & g[3710];
assign g[5759] = a[11] & g[3711];
assign g[7806] = b[11] & g[3711];
assign g[5760] = a[11] & g[3712];
assign g[7807] = b[11] & g[3712];
assign g[5761] = a[11] & g[3713];
assign g[7808] = b[11] & g[3713];
assign g[5762] = a[11] & g[3714];
assign g[7809] = b[11] & g[3714];
assign g[5763] = a[11] & g[3715];
assign g[7810] = b[11] & g[3715];
assign g[5764] = a[11] & g[3716];
assign g[7811] = b[11] & g[3716];
assign g[5765] = a[11] & g[3717];
assign g[7812] = b[11] & g[3717];
assign g[5766] = a[11] & g[3718];
assign g[7813] = b[11] & g[3718];
assign g[5767] = a[11] & g[3719];
assign g[7814] = b[11] & g[3719];
assign g[5768] = a[11] & g[3720];
assign g[7815] = b[11] & g[3720];
assign g[5769] = a[11] & g[3721];
assign g[7816] = b[11] & g[3721];
assign g[5770] = a[11] & g[3722];
assign g[7817] = b[11] & g[3722];
assign g[5771] = a[11] & g[3723];
assign g[7818] = b[11] & g[3723];
assign g[5772] = a[11] & g[3724];
assign g[7819] = b[11] & g[3724];
assign g[5773] = a[11] & g[3725];
assign g[7820] = b[11] & g[3725];
assign g[5774] = a[11] & g[3726];
assign g[7821] = b[11] & g[3726];
assign g[5775] = a[11] & g[3727];
assign g[7822] = b[11] & g[3727];
assign g[5776] = a[11] & g[3728];
assign g[7823] = b[11] & g[3728];
assign g[5777] = a[11] & g[3729];
assign g[7824] = b[11] & g[3729];
assign g[5778] = a[11] & g[3730];
assign g[7825] = b[11] & g[3730];
assign g[5779] = a[11] & g[3731];
assign g[7826] = b[11] & g[3731];
assign g[5780] = a[11] & g[3732];
assign g[7827] = b[11] & g[3732];
assign g[5781] = a[11] & g[3733];
assign g[7828] = b[11] & g[3733];
assign g[5782] = a[11] & g[3734];
assign g[7829] = b[11] & g[3734];
assign g[5783] = a[11] & g[3735];
assign g[7830] = b[11] & g[3735];
assign g[5784] = a[11] & g[3736];
assign g[7831] = b[11] & g[3736];
assign g[5785] = a[11] & g[3737];
assign g[7832] = b[11] & g[3737];
assign g[5786] = a[11] & g[3738];
assign g[7833] = b[11] & g[3738];
assign g[5787] = a[11] & g[3739];
assign g[7834] = b[11] & g[3739];
assign g[5788] = a[11] & g[3740];
assign g[7835] = b[11] & g[3740];
assign g[5789] = a[11] & g[3741];
assign g[7836] = b[11] & g[3741];
assign g[5790] = a[11] & g[3742];
assign g[7837] = b[11] & g[3742];
assign g[5791] = a[11] & g[3743];
assign g[7838] = b[11] & g[3743];
assign g[5792] = a[11] & g[3744];
assign g[7839] = b[11] & g[3744];
assign g[5793] = a[11] & g[3745];
assign g[7840] = b[11] & g[3745];
assign g[5794] = a[11] & g[3746];
assign g[7841] = b[11] & g[3746];
assign g[5795] = a[11] & g[3747];
assign g[7842] = b[11] & g[3747];
assign g[5796] = a[11] & g[3748];
assign g[7843] = b[11] & g[3748];
assign g[5797] = a[11] & g[3749];
assign g[7844] = b[11] & g[3749];
assign g[5798] = a[11] & g[3750];
assign g[7845] = b[11] & g[3750];
assign g[5799] = a[11] & g[3751];
assign g[7846] = b[11] & g[3751];
assign g[5800] = a[11] & g[3752];
assign g[7847] = b[11] & g[3752];
assign g[5801] = a[11] & g[3753];
assign g[7848] = b[11] & g[3753];
assign g[5802] = a[11] & g[3754];
assign g[7849] = b[11] & g[3754];
assign g[5803] = a[11] & g[3755];
assign g[7850] = b[11] & g[3755];
assign g[5804] = a[11] & g[3756];
assign g[7851] = b[11] & g[3756];
assign g[5805] = a[11] & g[3757];
assign g[7852] = b[11] & g[3757];
assign g[5806] = a[11] & g[3758];
assign g[7853] = b[11] & g[3758];
assign g[5807] = a[11] & g[3759];
assign g[7854] = b[11] & g[3759];
assign g[5808] = a[11] & g[3760];
assign g[7855] = b[11] & g[3760];
assign g[5809] = a[11] & g[3761];
assign g[7856] = b[11] & g[3761];
assign g[5810] = a[11] & g[3762];
assign g[7857] = b[11] & g[3762];
assign g[5811] = a[11] & g[3763];
assign g[7858] = b[11] & g[3763];
assign g[5812] = a[11] & g[3764];
assign g[7859] = b[11] & g[3764];
assign g[5813] = a[11] & g[3765];
assign g[7860] = b[11] & g[3765];
assign g[5814] = a[11] & g[3766];
assign g[7861] = b[11] & g[3766];
assign g[5815] = a[11] & g[3767];
assign g[7862] = b[11] & g[3767];
assign g[5816] = a[11] & g[3768];
assign g[7863] = b[11] & g[3768];
assign g[5817] = a[11] & g[3769];
assign g[7864] = b[11] & g[3769];
assign g[5818] = a[11] & g[3770];
assign g[7865] = b[11] & g[3770];
assign g[5819] = a[11] & g[3771];
assign g[7866] = b[11] & g[3771];
assign g[5820] = a[11] & g[3772];
assign g[7867] = b[11] & g[3772];
assign g[5821] = a[11] & g[3773];
assign g[7868] = b[11] & g[3773];
assign g[5822] = a[11] & g[3774];
assign g[7869] = b[11] & g[3774];
assign g[5823] = a[11] & g[3775];
assign g[7870] = b[11] & g[3775];
assign g[5824] = a[11] & g[3776];
assign g[7871] = b[11] & g[3776];
assign g[5825] = a[11] & g[3777];
assign g[7872] = b[11] & g[3777];
assign g[5826] = a[11] & g[3778];
assign g[7873] = b[11] & g[3778];
assign g[5827] = a[11] & g[3779];
assign g[7874] = b[11] & g[3779];
assign g[5828] = a[11] & g[3780];
assign g[7875] = b[11] & g[3780];
assign g[5829] = a[11] & g[3781];
assign g[7876] = b[11] & g[3781];
assign g[5830] = a[11] & g[3782];
assign g[7877] = b[11] & g[3782];
assign g[5831] = a[11] & g[3783];
assign g[7878] = b[11] & g[3783];
assign g[5832] = a[11] & g[3784];
assign g[7879] = b[11] & g[3784];
assign g[5833] = a[11] & g[3785];
assign g[7880] = b[11] & g[3785];
assign g[5834] = a[11] & g[3786];
assign g[7881] = b[11] & g[3786];
assign g[5835] = a[11] & g[3787];
assign g[7882] = b[11] & g[3787];
assign g[5836] = a[11] & g[3788];
assign g[7883] = b[11] & g[3788];
assign g[5837] = a[11] & g[3789];
assign g[7884] = b[11] & g[3789];
assign g[5838] = a[11] & g[3790];
assign g[7885] = b[11] & g[3790];
assign g[5839] = a[11] & g[3791];
assign g[7886] = b[11] & g[3791];
assign g[5840] = a[11] & g[3792];
assign g[7887] = b[11] & g[3792];
assign g[5841] = a[11] & g[3793];
assign g[7888] = b[11] & g[3793];
assign g[5842] = a[11] & g[3794];
assign g[7889] = b[11] & g[3794];
assign g[5843] = a[11] & g[3795];
assign g[7890] = b[11] & g[3795];
assign g[5844] = a[11] & g[3796];
assign g[7891] = b[11] & g[3796];
assign g[5845] = a[11] & g[3797];
assign g[7892] = b[11] & g[3797];
assign g[5846] = a[11] & g[3798];
assign g[7893] = b[11] & g[3798];
assign g[5847] = a[11] & g[3799];
assign g[7894] = b[11] & g[3799];
assign g[5848] = a[11] & g[3800];
assign g[7895] = b[11] & g[3800];
assign g[5849] = a[11] & g[3801];
assign g[7896] = b[11] & g[3801];
assign g[5850] = a[11] & g[3802];
assign g[7897] = b[11] & g[3802];
assign g[5851] = a[11] & g[3803];
assign g[7898] = b[11] & g[3803];
assign g[5852] = a[11] & g[3804];
assign g[7899] = b[11] & g[3804];
assign g[5853] = a[11] & g[3805];
assign g[7900] = b[11] & g[3805];
assign g[5854] = a[11] & g[3806];
assign g[7901] = b[11] & g[3806];
assign g[5855] = a[11] & g[3807];
assign g[7902] = b[11] & g[3807];
assign g[5856] = a[11] & g[3808];
assign g[7903] = b[11] & g[3808];
assign g[5857] = a[11] & g[3809];
assign g[7904] = b[11] & g[3809];
assign g[5858] = a[11] & g[3810];
assign g[7905] = b[11] & g[3810];
assign g[5859] = a[11] & g[3811];
assign g[7906] = b[11] & g[3811];
assign g[5860] = a[11] & g[3812];
assign g[7907] = b[11] & g[3812];
assign g[5861] = a[11] & g[3813];
assign g[7908] = b[11] & g[3813];
assign g[5862] = a[11] & g[3814];
assign g[7909] = b[11] & g[3814];
assign g[5863] = a[11] & g[3815];
assign g[7910] = b[11] & g[3815];
assign g[5864] = a[11] & g[3816];
assign g[7911] = b[11] & g[3816];
assign g[5865] = a[11] & g[3817];
assign g[7912] = b[11] & g[3817];
assign g[5866] = a[11] & g[3818];
assign g[7913] = b[11] & g[3818];
assign g[5867] = a[11] & g[3819];
assign g[7914] = b[11] & g[3819];
assign g[5868] = a[11] & g[3820];
assign g[7915] = b[11] & g[3820];
assign g[5869] = a[11] & g[3821];
assign g[7916] = b[11] & g[3821];
assign g[5870] = a[11] & g[3822];
assign g[7917] = b[11] & g[3822];
assign g[5871] = a[11] & g[3823];
assign g[7918] = b[11] & g[3823];
assign g[5872] = a[11] & g[3824];
assign g[7919] = b[11] & g[3824];
assign g[5873] = a[11] & g[3825];
assign g[7920] = b[11] & g[3825];
assign g[5874] = a[11] & g[3826];
assign g[7921] = b[11] & g[3826];
assign g[5875] = a[11] & g[3827];
assign g[7922] = b[11] & g[3827];
assign g[5876] = a[11] & g[3828];
assign g[7923] = b[11] & g[3828];
assign g[5877] = a[11] & g[3829];
assign g[7924] = b[11] & g[3829];
assign g[5878] = a[11] & g[3830];
assign g[7925] = b[11] & g[3830];
assign g[5879] = a[11] & g[3831];
assign g[7926] = b[11] & g[3831];
assign g[5880] = a[11] & g[3832];
assign g[7927] = b[11] & g[3832];
assign g[5881] = a[11] & g[3833];
assign g[7928] = b[11] & g[3833];
assign g[5882] = a[11] & g[3834];
assign g[7929] = b[11] & g[3834];
assign g[5883] = a[11] & g[3835];
assign g[7930] = b[11] & g[3835];
assign g[5884] = a[11] & g[3836];
assign g[7931] = b[11] & g[3836];
assign g[5885] = a[11] & g[3837];
assign g[7932] = b[11] & g[3837];
assign g[5886] = a[11] & g[3838];
assign g[7933] = b[11] & g[3838];
assign g[5887] = a[11] & g[3839];
assign g[7934] = b[11] & g[3839];
assign g[5888] = a[11] & g[3840];
assign g[7935] = b[11] & g[3840];
assign g[5889] = a[11] & g[3841];
assign g[7936] = b[11] & g[3841];
assign g[5890] = a[11] & g[3842];
assign g[7937] = b[11] & g[3842];
assign g[5891] = a[11] & g[3843];
assign g[7938] = b[11] & g[3843];
assign g[5892] = a[11] & g[3844];
assign g[7939] = b[11] & g[3844];
assign g[5893] = a[11] & g[3845];
assign g[7940] = b[11] & g[3845];
assign g[5894] = a[11] & g[3846];
assign g[7941] = b[11] & g[3846];
assign g[5895] = a[11] & g[3847];
assign g[7942] = b[11] & g[3847];
assign g[5896] = a[11] & g[3848];
assign g[7943] = b[11] & g[3848];
assign g[5897] = a[11] & g[3849];
assign g[7944] = b[11] & g[3849];
assign g[5898] = a[11] & g[3850];
assign g[7945] = b[11] & g[3850];
assign g[5899] = a[11] & g[3851];
assign g[7946] = b[11] & g[3851];
assign g[5900] = a[11] & g[3852];
assign g[7947] = b[11] & g[3852];
assign g[5901] = a[11] & g[3853];
assign g[7948] = b[11] & g[3853];
assign g[5902] = a[11] & g[3854];
assign g[7949] = b[11] & g[3854];
assign g[5903] = a[11] & g[3855];
assign g[7950] = b[11] & g[3855];
assign g[5904] = a[11] & g[3856];
assign g[7951] = b[11] & g[3856];
assign g[5905] = a[11] & g[3857];
assign g[7952] = b[11] & g[3857];
assign g[5906] = a[11] & g[3858];
assign g[7953] = b[11] & g[3858];
assign g[5907] = a[11] & g[3859];
assign g[7954] = b[11] & g[3859];
assign g[5908] = a[11] & g[3860];
assign g[7955] = b[11] & g[3860];
assign g[5909] = a[11] & g[3861];
assign g[7956] = b[11] & g[3861];
assign g[5910] = a[11] & g[3862];
assign g[7957] = b[11] & g[3862];
assign g[5911] = a[11] & g[3863];
assign g[7958] = b[11] & g[3863];
assign g[5912] = a[11] & g[3864];
assign g[7959] = b[11] & g[3864];
assign g[5913] = a[11] & g[3865];
assign g[7960] = b[11] & g[3865];
assign g[5914] = a[11] & g[3866];
assign g[7961] = b[11] & g[3866];
assign g[5915] = a[11] & g[3867];
assign g[7962] = b[11] & g[3867];
assign g[5916] = a[11] & g[3868];
assign g[7963] = b[11] & g[3868];
assign g[5917] = a[11] & g[3869];
assign g[7964] = b[11] & g[3869];
assign g[5918] = a[11] & g[3870];
assign g[7965] = b[11] & g[3870];
assign g[5919] = a[11] & g[3871];
assign g[7966] = b[11] & g[3871];
assign g[5920] = a[11] & g[3872];
assign g[7967] = b[11] & g[3872];
assign g[5921] = a[11] & g[3873];
assign g[7968] = b[11] & g[3873];
assign g[5922] = a[11] & g[3874];
assign g[7969] = b[11] & g[3874];
assign g[5923] = a[11] & g[3875];
assign g[7970] = b[11] & g[3875];
assign g[5924] = a[11] & g[3876];
assign g[7971] = b[11] & g[3876];
assign g[5925] = a[11] & g[3877];
assign g[7972] = b[11] & g[3877];
assign g[5926] = a[11] & g[3878];
assign g[7973] = b[11] & g[3878];
assign g[5927] = a[11] & g[3879];
assign g[7974] = b[11] & g[3879];
assign g[5928] = a[11] & g[3880];
assign g[7975] = b[11] & g[3880];
assign g[5929] = a[11] & g[3881];
assign g[7976] = b[11] & g[3881];
assign g[5930] = a[11] & g[3882];
assign g[7977] = b[11] & g[3882];
assign g[5931] = a[11] & g[3883];
assign g[7978] = b[11] & g[3883];
assign g[5932] = a[11] & g[3884];
assign g[7979] = b[11] & g[3884];
assign g[5933] = a[11] & g[3885];
assign g[7980] = b[11] & g[3885];
assign g[5934] = a[11] & g[3886];
assign g[7981] = b[11] & g[3886];
assign g[5935] = a[11] & g[3887];
assign g[7982] = b[11] & g[3887];
assign g[5936] = a[11] & g[3888];
assign g[7983] = b[11] & g[3888];
assign g[5937] = a[11] & g[3889];
assign g[7984] = b[11] & g[3889];
assign g[5938] = a[11] & g[3890];
assign g[7985] = b[11] & g[3890];
assign g[5939] = a[11] & g[3891];
assign g[7986] = b[11] & g[3891];
assign g[5940] = a[11] & g[3892];
assign g[7987] = b[11] & g[3892];
assign g[5941] = a[11] & g[3893];
assign g[7988] = b[11] & g[3893];
assign g[5942] = a[11] & g[3894];
assign g[7989] = b[11] & g[3894];
assign g[5943] = a[11] & g[3895];
assign g[7990] = b[11] & g[3895];
assign g[5944] = a[11] & g[3896];
assign g[7991] = b[11] & g[3896];
assign g[5945] = a[11] & g[3897];
assign g[7992] = b[11] & g[3897];
assign g[5946] = a[11] & g[3898];
assign g[7993] = b[11] & g[3898];
assign g[5947] = a[11] & g[3899];
assign g[7994] = b[11] & g[3899];
assign g[5948] = a[11] & g[3900];
assign g[7995] = b[11] & g[3900];
assign g[5949] = a[11] & g[3901];
assign g[7996] = b[11] & g[3901];
assign g[5950] = a[11] & g[3902];
assign g[7997] = b[11] & g[3902];
assign g[5951] = a[11] & g[3903];
assign g[7998] = b[11] & g[3903];
assign g[5952] = a[11] & g[3904];
assign g[7999] = b[11] & g[3904];
assign g[5953] = a[11] & g[3905];
assign g[8000] = b[11] & g[3905];
assign g[5954] = a[11] & g[3906];
assign g[8001] = b[11] & g[3906];
assign g[5955] = a[11] & g[3907];
assign g[8002] = b[11] & g[3907];
assign g[5956] = a[11] & g[3908];
assign g[8003] = b[11] & g[3908];
assign g[5957] = a[11] & g[3909];
assign g[8004] = b[11] & g[3909];
assign g[5958] = a[11] & g[3910];
assign g[8005] = b[11] & g[3910];
assign g[5959] = a[11] & g[3911];
assign g[8006] = b[11] & g[3911];
assign g[5960] = a[11] & g[3912];
assign g[8007] = b[11] & g[3912];
assign g[5961] = a[11] & g[3913];
assign g[8008] = b[11] & g[3913];
assign g[5962] = a[11] & g[3914];
assign g[8009] = b[11] & g[3914];
assign g[5963] = a[11] & g[3915];
assign g[8010] = b[11] & g[3915];
assign g[5964] = a[11] & g[3916];
assign g[8011] = b[11] & g[3916];
assign g[5965] = a[11] & g[3917];
assign g[8012] = b[11] & g[3917];
assign g[5966] = a[11] & g[3918];
assign g[8013] = b[11] & g[3918];
assign g[5967] = a[11] & g[3919];
assign g[8014] = b[11] & g[3919];
assign g[5968] = a[11] & g[3920];
assign g[8015] = b[11] & g[3920];
assign g[5969] = a[11] & g[3921];
assign g[8016] = b[11] & g[3921];
assign g[5970] = a[11] & g[3922];
assign g[8017] = b[11] & g[3922];
assign g[5971] = a[11] & g[3923];
assign g[8018] = b[11] & g[3923];
assign g[5972] = a[11] & g[3924];
assign g[8019] = b[11] & g[3924];
assign g[5973] = a[11] & g[3925];
assign g[8020] = b[11] & g[3925];
assign g[5974] = a[11] & g[3926];
assign g[8021] = b[11] & g[3926];
assign g[5975] = a[11] & g[3927];
assign g[8022] = b[11] & g[3927];
assign g[5976] = a[11] & g[3928];
assign g[8023] = b[11] & g[3928];
assign g[5977] = a[11] & g[3929];
assign g[8024] = b[11] & g[3929];
assign g[5978] = a[11] & g[3930];
assign g[8025] = b[11] & g[3930];
assign g[5979] = a[11] & g[3931];
assign g[8026] = b[11] & g[3931];
assign g[5980] = a[11] & g[3932];
assign g[8027] = b[11] & g[3932];
assign g[5981] = a[11] & g[3933];
assign g[8028] = b[11] & g[3933];
assign g[5982] = a[11] & g[3934];
assign g[8029] = b[11] & g[3934];
assign g[5983] = a[11] & g[3935];
assign g[8030] = b[11] & g[3935];
assign g[5984] = a[11] & g[3936];
assign g[8031] = b[11] & g[3936];
assign g[5985] = a[11] & g[3937];
assign g[8032] = b[11] & g[3937];
assign g[5986] = a[11] & g[3938];
assign g[8033] = b[11] & g[3938];
assign g[5987] = a[11] & g[3939];
assign g[8034] = b[11] & g[3939];
assign g[5988] = a[11] & g[3940];
assign g[8035] = b[11] & g[3940];
assign g[5989] = a[11] & g[3941];
assign g[8036] = b[11] & g[3941];
assign g[5990] = a[11] & g[3942];
assign g[8037] = b[11] & g[3942];
assign g[5991] = a[11] & g[3943];
assign g[8038] = b[11] & g[3943];
assign g[5992] = a[11] & g[3944];
assign g[8039] = b[11] & g[3944];
assign g[5993] = a[11] & g[3945];
assign g[8040] = b[11] & g[3945];
assign g[5994] = a[11] & g[3946];
assign g[8041] = b[11] & g[3946];
assign g[5995] = a[11] & g[3947];
assign g[8042] = b[11] & g[3947];
assign g[5996] = a[11] & g[3948];
assign g[8043] = b[11] & g[3948];
assign g[5997] = a[11] & g[3949];
assign g[8044] = b[11] & g[3949];
assign g[5998] = a[11] & g[3950];
assign g[8045] = b[11] & g[3950];
assign g[5999] = a[11] & g[3951];
assign g[8046] = b[11] & g[3951];
assign g[6000] = a[11] & g[3952];
assign g[8047] = b[11] & g[3952];
assign g[6001] = a[11] & g[3953];
assign g[8048] = b[11] & g[3953];
assign g[6002] = a[11] & g[3954];
assign g[8049] = b[11] & g[3954];
assign g[6003] = a[11] & g[3955];
assign g[8050] = b[11] & g[3955];
assign g[6004] = a[11] & g[3956];
assign g[8051] = b[11] & g[3956];
assign g[6005] = a[11] & g[3957];
assign g[8052] = b[11] & g[3957];
assign g[6006] = a[11] & g[3958];
assign g[8053] = b[11] & g[3958];
assign g[6007] = a[11] & g[3959];
assign g[8054] = b[11] & g[3959];
assign g[6008] = a[11] & g[3960];
assign g[8055] = b[11] & g[3960];
assign g[6009] = a[11] & g[3961];
assign g[8056] = b[11] & g[3961];
assign g[6010] = a[11] & g[3962];
assign g[8057] = b[11] & g[3962];
assign g[6011] = a[11] & g[3963];
assign g[8058] = b[11] & g[3963];
assign g[6012] = a[11] & g[3964];
assign g[8059] = b[11] & g[3964];
assign g[6013] = a[11] & g[3965];
assign g[8060] = b[11] & g[3965];
assign g[6014] = a[11] & g[3966];
assign g[8061] = b[11] & g[3966];
assign g[6015] = a[11] & g[3967];
assign g[8062] = b[11] & g[3967];
assign g[6016] = a[11] & g[3968];
assign g[8063] = b[11] & g[3968];
assign g[6017] = a[11] & g[3969];
assign g[8064] = b[11] & g[3969];
assign g[6018] = a[11] & g[3970];
assign g[8065] = b[11] & g[3970];
assign g[6019] = a[11] & g[3971];
assign g[8066] = b[11] & g[3971];
assign g[6020] = a[11] & g[3972];
assign g[8067] = b[11] & g[3972];
assign g[6021] = a[11] & g[3973];
assign g[8068] = b[11] & g[3973];
assign g[6022] = a[11] & g[3974];
assign g[8069] = b[11] & g[3974];
assign g[6023] = a[11] & g[3975];
assign g[8070] = b[11] & g[3975];
assign g[6024] = a[11] & g[3976];
assign g[8071] = b[11] & g[3976];
assign g[6025] = a[11] & g[3977];
assign g[8072] = b[11] & g[3977];
assign g[6026] = a[11] & g[3978];
assign g[8073] = b[11] & g[3978];
assign g[6027] = a[11] & g[3979];
assign g[8074] = b[11] & g[3979];
assign g[6028] = a[11] & g[3980];
assign g[8075] = b[11] & g[3980];
assign g[6029] = a[11] & g[3981];
assign g[8076] = b[11] & g[3981];
assign g[6030] = a[11] & g[3982];
assign g[8077] = b[11] & g[3982];
assign g[6031] = a[11] & g[3983];
assign g[8078] = b[11] & g[3983];
assign g[6032] = a[11] & g[3984];
assign g[8079] = b[11] & g[3984];
assign g[6033] = a[11] & g[3985];
assign g[8080] = b[11] & g[3985];
assign g[6034] = a[11] & g[3986];
assign g[8081] = b[11] & g[3986];
assign g[6035] = a[11] & g[3987];
assign g[8082] = b[11] & g[3987];
assign g[6036] = a[11] & g[3988];
assign g[8083] = b[11] & g[3988];
assign g[6037] = a[11] & g[3989];
assign g[8084] = b[11] & g[3989];
assign g[6038] = a[11] & g[3990];
assign g[8085] = b[11] & g[3990];
assign g[6039] = a[11] & g[3991];
assign g[8086] = b[11] & g[3991];
assign g[6040] = a[11] & g[3992];
assign g[8087] = b[11] & g[3992];
assign g[6041] = a[11] & g[3993];
assign g[8088] = b[11] & g[3993];
assign g[6042] = a[11] & g[3994];
assign g[8089] = b[11] & g[3994];
assign g[6043] = a[11] & g[3995];
assign g[8090] = b[11] & g[3995];
assign g[6044] = a[11] & g[3996];
assign g[8091] = b[11] & g[3996];
assign g[6045] = a[11] & g[3997];
assign g[8092] = b[11] & g[3997];
assign g[6046] = a[11] & g[3998];
assign g[8093] = b[11] & g[3998];
assign g[6047] = a[11] & g[3999];
assign g[8094] = b[11] & g[3999];
assign g[6048] = a[11] & g[4000];
assign g[8095] = b[11] & g[4000];
assign g[6049] = a[11] & g[4001];
assign g[8096] = b[11] & g[4001];
assign g[6050] = a[11] & g[4002];
assign g[8097] = b[11] & g[4002];
assign g[6051] = a[11] & g[4003];
assign g[8098] = b[11] & g[4003];
assign g[6052] = a[11] & g[4004];
assign g[8099] = b[11] & g[4004];
assign g[6053] = a[11] & g[4005];
assign g[8100] = b[11] & g[4005];
assign g[6054] = a[11] & g[4006];
assign g[8101] = b[11] & g[4006];
assign g[6055] = a[11] & g[4007];
assign g[8102] = b[11] & g[4007];
assign g[6056] = a[11] & g[4008];
assign g[8103] = b[11] & g[4008];
assign g[6057] = a[11] & g[4009];
assign g[8104] = b[11] & g[4009];
assign g[6058] = a[11] & g[4010];
assign g[8105] = b[11] & g[4010];
assign g[6059] = a[11] & g[4011];
assign g[8106] = b[11] & g[4011];
assign g[6060] = a[11] & g[4012];
assign g[8107] = b[11] & g[4012];
assign g[6061] = a[11] & g[4013];
assign g[8108] = b[11] & g[4013];
assign g[6062] = a[11] & g[4014];
assign g[8109] = b[11] & g[4014];
assign g[6063] = a[11] & g[4015];
assign g[8110] = b[11] & g[4015];
assign g[6064] = a[11] & g[4016];
assign g[8111] = b[11] & g[4016];
assign g[6065] = a[11] & g[4017];
assign g[8112] = b[11] & g[4017];
assign g[6066] = a[11] & g[4018];
assign g[8113] = b[11] & g[4018];
assign g[6067] = a[11] & g[4019];
assign g[8114] = b[11] & g[4019];
assign g[6068] = a[11] & g[4020];
assign g[8115] = b[11] & g[4020];
assign g[6069] = a[11] & g[4021];
assign g[8116] = b[11] & g[4021];
assign g[6070] = a[11] & g[4022];
assign g[8117] = b[11] & g[4022];
assign g[6071] = a[11] & g[4023];
assign g[8118] = b[11] & g[4023];
assign g[6072] = a[11] & g[4024];
assign g[8119] = b[11] & g[4024];
assign g[6073] = a[11] & g[4025];
assign g[8120] = b[11] & g[4025];
assign g[6074] = a[11] & g[4026];
assign g[8121] = b[11] & g[4026];
assign g[6075] = a[11] & g[4027];
assign g[8122] = b[11] & g[4027];
assign g[6076] = a[11] & g[4028];
assign g[8123] = b[11] & g[4028];
assign g[6077] = a[11] & g[4029];
assign g[8124] = b[11] & g[4029];
assign g[6078] = a[11] & g[4030];
assign g[8125] = b[11] & g[4030];
assign g[6079] = a[11] & g[4031];
assign g[8126] = b[11] & g[4031];
assign g[6080] = a[11] & g[4032];
assign g[8127] = b[11] & g[4032];
assign g[6081] = a[11] & g[4033];
assign g[8128] = b[11] & g[4033];
assign g[6082] = a[11] & g[4034];
assign g[8129] = b[11] & g[4034];
assign g[6083] = a[11] & g[4035];
assign g[8130] = b[11] & g[4035];
assign g[6084] = a[11] & g[4036];
assign g[8131] = b[11] & g[4036];
assign g[6085] = a[11] & g[4037];
assign g[8132] = b[11] & g[4037];
assign g[6086] = a[11] & g[4038];
assign g[8133] = b[11] & g[4038];
assign g[6087] = a[11] & g[4039];
assign g[8134] = b[11] & g[4039];
assign g[6088] = a[11] & g[4040];
assign g[8135] = b[11] & g[4040];
assign g[6089] = a[11] & g[4041];
assign g[8136] = b[11] & g[4041];
assign g[6090] = a[11] & g[4042];
assign g[8137] = b[11] & g[4042];
assign g[6091] = a[11] & g[4043];
assign g[8138] = b[11] & g[4043];
assign g[6092] = a[11] & g[4044];
assign g[8139] = b[11] & g[4044];
assign g[6093] = a[11] & g[4045];
assign g[8140] = b[11] & g[4045];
assign g[6094] = a[11] & g[4046];
assign g[8141] = b[11] & g[4046];
assign g[6095] = a[11] & g[4047];
assign g[8142] = b[11] & g[4047];
assign g[6096] = a[11] & g[4048];
assign g[8143] = b[11] & g[4048];
assign g[6097] = a[11] & g[4049];
assign g[8144] = b[11] & g[4049];
assign g[6098] = a[11] & g[4050];
assign g[8145] = b[11] & g[4050];
assign g[6099] = a[11] & g[4051];
assign g[8146] = b[11] & g[4051];
assign g[6100] = a[11] & g[4052];
assign g[8147] = b[11] & g[4052];
assign g[6101] = a[11] & g[4053];
assign g[8148] = b[11] & g[4053];
assign g[6102] = a[11] & g[4054];
assign g[8149] = b[11] & g[4054];
assign g[6103] = a[11] & g[4055];
assign g[8150] = b[11] & g[4055];
assign g[6104] = a[11] & g[4056];
assign g[8151] = b[11] & g[4056];
assign g[6105] = a[11] & g[4057];
assign g[8152] = b[11] & g[4057];
assign g[6106] = a[11] & g[4058];
assign g[8153] = b[11] & g[4058];
assign g[6107] = a[11] & g[4059];
assign g[8154] = b[11] & g[4059];
assign g[6108] = a[11] & g[4060];
assign g[8155] = b[11] & g[4060];
assign g[6109] = a[11] & g[4061];
assign g[8156] = b[11] & g[4061];
assign g[6110] = a[11] & g[4062];
assign g[8157] = b[11] & g[4062];
assign g[6111] = a[11] & g[4063];
assign g[8158] = b[11] & g[4063];
assign g[6112] = a[11] & g[4064];
assign g[8159] = b[11] & g[4064];
assign g[6113] = a[11] & g[4065];
assign g[8160] = b[11] & g[4065];
assign g[6114] = a[11] & g[4066];
assign g[8161] = b[11] & g[4066];
assign g[6115] = a[11] & g[4067];
assign g[8162] = b[11] & g[4067];
assign g[6116] = a[11] & g[4068];
assign g[8163] = b[11] & g[4068];
assign g[6117] = a[11] & g[4069];
assign g[8164] = b[11] & g[4069];
assign g[6118] = a[11] & g[4070];
assign g[8165] = b[11] & g[4070];
assign g[6119] = a[11] & g[4071];
assign g[8166] = b[11] & g[4071];
assign g[6120] = a[11] & g[4072];
assign g[8167] = b[11] & g[4072];
assign g[6121] = a[11] & g[4073];
assign g[8168] = b[11] & g[4073];
assign g[6122] = a[11] & g[4074];
assign g[8169] = b[11] & g[4074];
assign g[6123] = a[11] & g[4075];
assign g[8170] = b[11] & g[4075];
assign g[6124] = a[11] & g[4076];
assign g[8171] = b[11] & g[4076];
assign g[6125] = a[11] & g[4077];
assign g[8172] = b[11] & g[4077];
assign g[6126] = a[11] & g[4078];
assign g[8173] = b[11] & g[4078];
assign g[6127] = a[11] & g[4079];
assign g[8174] = b[11] & g[4079];
assign g[6128] = a[11] & g[4080];
assign g[8175] = b[11] & g[4080];
assign g[6129] = a[11] & g[4081];
assign g[8176] = b[11] & g[4081];
assign g[6130] = a[11] & g[4082];
assign g[8177] = b[11] & g[4082];
//Assigning outputs for input bit 13
assign g[8178] = a[12] & b[12];
assign g[8179] = a[12] & g[4083];
assign g[12274] = b[12] & g[4083];
assign g[8180] = a[12] & g[4084];
assign g[12275] = b[12] & g[4084];
assign g[8181] = a[12] & g[4085];
assign g[12276] = b[12] & g[4085];
assign g[8182] = a[12] & g[4086];
assign g[12277] = b[12] & g[4086];
assign g[8183] = a[12] & g[4087];
assign g[12278] = b[12] & g[4087];
assign g[8184] = a[12] & g[4088];
assign g[12279] = b[12] & g[4088];
assign g[8185] = a[12] & g[4089];
assign g[12280] = b[12] & g[4089];
assign g[8186] = a[12] & g[4090];
assign g[12281] = b[12] & g[4090];
assign g[8187] = a[12] & g[4091];
assign g[12282] = b[12] & g[4091];
assign g[8188] = a[12] & g[4092];
assign g[12283] = b[12] & g[4092];
assign g[8189] = a[12] & g[4093];
assign g[12284] = b[12] & g[4093];
assign g[8190] = a[12] & g[4094];
assign g[12285] = b[12] & g[4094];
assign g[8191] = a[12] & g[4095];
assign g[12286] = b[12] & g[4095];
assign g[8192] = a[12] & g[4096];
assign g[12287] = b[12] & g[4096];
assign g[8193] = a[12] & g[4097];
assign g[12288] = b[12] & g[4097];
assign g[8194] = a[12] & g[4098];
assign g[12289] = b[12] & g[4098];
assign g[8195] = a[12] & g[4099];
assign g[12290] = b[12] & g[4099];
assign g[8196] = a[12] & g[4100];
assign g[12291] = b[12] & g[4100];
assign g[8197] = a[12] & g[4101];
assign g[12292] = b[12] & g[4101];
assign g[8198] = a[12] & g[4102];
assign g[12293] = b[12] & g[4102];
assign g[8199] = a[12] & g[4103];
assign g[12294] = b[12] & g[4103];
assign g[8200] = a[12] & g[4104];
assign g[12295] = b[12] & g[4104];
assign g[8201] = a[12] & g[4105];
assign g[12296] = b[12] & g[4105];
assign g[8202] = a[12] & g[4106];
assign g[12297] = b[12] & g[4106];
assign g[8203] = a[12] & g[4107];
assign g[12298] = b[12] & g[4107];
assign g[8204] = a[12] & g[4108];
assign g[12299] = b[12] & g[4108];
assign g[8205] = a[12] & g[4109];
assign g[12300] = b[12] & g[4109];
assign g[8206] = a[12] & g[4110];
assign g[12301] = b[12] & g[4110];
assign g[8207] = a[12] & g[4111];
assign g[12302] = b[12] & g[4111];
assign g[8208] = a[12] & g[4112];
assign g[12303] = b[12] & g[4112];
assign g[8209] = a[12] & g[4113];
assign g[12304] = b[12] & g[4113];
assign g[8210] = a[12] & g[4114];
assign g[12305] = b[12] & g[4114];
assign g[8211] = a[12] & g[4115];
assign g[12306] = b[12] & g[4115];
assign g[8212] = a[12] & g[4116];
assign g[12307] = b[12] & g[4116];
assign g[8213] = a[12] & g[4117];
assign g[12308] = b[12] & g[4117];
assign g[8214] = a[12] & g[4118];
assign g[12309] = b[12] & g[4118];
assign g[8215] = a[12] & g[4119];
assign g[12310] = b[12] & g[4119];
assign g[8216] = a[12] & g[4120];
assign g[12311] = b[12] & g[4120];
assign g[8217] = a[12] & g[4121];
assign g[12312] = b[12] & g[4121];
assign g[8218] = a[12] & g[4122];
assign g[12313] = b[12] & g[4122];
assign g[8219] = a[12] & g[4123];
assign g[12314] = b[12] & g[4123];
assign g[8220] = a[12] & g[4124];
assign g[12315] = b[12] & g[4124];
assign g[8221] = a[12] & g[4125];
assign g[12316] = b[12] & g[4125];
assign g[8222] = a[12] & g[4126];
assign g[12317] = b[12] & g[4126];
assign g[8223] = a[12] & g[4127];
assign g[12318] = b[12] & g[4127];
assign g[8224] = a[12] & g[4128];
assign g[12319] = b[12] & g[4128];
assign g[8225] = a[12] & g[4129];
assign g[12320] = b[12] & g[4129];
assign g[8226] = a[12] & g[4130];
assign g[12321] = b[12] & g[4130];
assign g[8227] = a[12] & g[4131];
assign g[12322] = b[12] & g[4131];
assign g[8228] = a[12] & g[4132];
assign g[12323] = b[12] & g[4132];
assign g[8229] = a[12] & g[4133];
assign g[12324] = b[12] & g[4133];
assign g[8230] = a[12] & g[4134];
assign g[12325] = b[12] & g[4134];
assign g[8231] = a[12] & g[4135];
assign g[12326] = b[12] & g[4135];
assign g[8232] = a[12] & g[4136];
assign g[12327] = b[12] & g[4136];
assign g[8233] = a[12] & g[4137];
assign g[12328] = b[12] & g[4137];
assign g[8234] = a[12] & g[4138];
assign g[12329] = b[12] & g[4138];
assign g[8235] = a[12] & g[4139];
assign g[12330] = b[12] & g[4139];
assign g[8236] = a[12] & g[4140];
assign g[12331] = b[12] & g[4140];
assign g[8237] = a[12] & g[4141];
assign g[12332] = b[12] & g[4141];
assign g[8238] = a[12] & g[4142];
assign g[12333] = b[12] & g[4142];
assign g[8239] = a[12] & g[4143];
assign g[12334] = b[12] & g[4143];
assign g[8240] = a[12] & g[4144];
assign g[12335] = b[12] & g[4144];
assign g[8241] = a[12] & g[4145];
assign g[12336] = b[12] & g[4145];
assign g[8242] = a[12] & g[4146];
assign g[12337] = b[12] & g[4146];
assign g[8243] = a[12] & g[4147];
assign g[12338] = b[12] & g[4147];
assign g[8244] = a[12] & g[4148];
assign g[12339] = b[12] & g[4148];
assign g[8245] = a[12] & g[4149];
assign g[12340] = b[12] & g[4149];
assign g[8246] = a[12] & g[4150];
assign g[12341] = b[12] & g[4150];
assign g[8247] = a[12] & g[4151];
assign g[12342] = b[12] & g[4151];
assign g[8248] = a[12] & g[4152];
assign g[12343] = b[12] & g[4152];
assign g[8249] = a[12] & g[4153];
assign g[12344] = b[12] & g[4153];
assign g[8250] = a[12] & g[4154];
assign g[12345] = b[12] & g[4154];
assign g[8251] = a[12] & g[4155];
assign g[12346] = b[12] & g[4155];
assign g[8252] = a[12] & g[4156];
assign g[12347] = b[12] & g[4156];
assign g[8253] = a[12] & g[4157];
assign g[12348] = b[12] & g[4157];
assign g[8254] = a[12] & g[4158];
assign g[12349] = b[12] & g[4158];
assign g[8255] = a[12] & g[4159];
assign g[12350] = b[12] & g[4159];
assign g[8256] = a[12] & g[4160];
assign g[12351] = b[12] & g[4160];
assign g[8257] = a[12] & g[4161];
assign g[12352] = b[12] & g[4161];
assign g[8258] = a[12] & g[4162];
assign g[12353] = b[12] & g[4162];
assign g[8259] = a[12] & g[4163];
assign g[12354] = b[12] & g[4163];
assign g[8260] = a[12] & g[4164];
assign g[12355] = b[12] & g[4164];
assign g[8261] = a[12] & g[4165];
assign g[12356] = b[12] & g[4165];
assign g[8262] = a[12] & g[4166];
assign g[12357] = b[12] & g[4166];
assign g[8263] = a[12] & g[4167];
assign g[12358] = b[12] & g[4167];
assign g[8264] = a[12] & g[4168];
assign g[12359] = b[12] & g[4168];
assign g[8265] = a[12] & g[4169];
assign g[12360] = b[12] & g[4169];
assign g[8266] = a[12] & g[4170];
assign g[12361] = b[12] & g[4170];
assign g[8267] = a[12] & g[4171];
assign g[12362] = b[12] & g[4171];
assign g[8268] = a[12] & g[4172];
assign g[12363] = b[12] & g[4172];
assign g[8269] = a[12] & g[4173];
assign g[12364] = b[12] & g[4173];
assign g[8270] = a[12] & g[4174];
assign g[12365] = b[12] & g[4174];
assign g[8271] = a[12] & g[4175];
assign g[12366] = b[12] & g[4175];
assign g[8272] = a[12] & g[4176];
assign g[12367] = b[12] & g[4176];
assign g[8273] = a[12] & g[4177];
assign g[12368] = b[12] & g[4177];
assign g[8274] = a[12] & g[4178];
assign g[12369] = b[12] & g[4178];
assign g[8275] = a[12] & g[4179];
assign g[12370] = b[12] & g[4179];
assign g[8276] = a[12] & g[4180];
assign g[12371] = b[12] & g[4180];
assign g[8277] = a[12] & g[4181];
assign g[12372] = b[12] & g[4181];
assign g[8278] = a[12] & g[4182];
assign g[12373] = b[12] & g[4182];
assign g[8279] = a[12] & g[4183];
assign g[12374] = b[12] & g[4183];
assign g[8280] = a[12] & g[4184];
assign g[12375] = b[12] & g[4184];
assign g[8281] = a[12] & g[4185];
assign g[12376] = b[12] & g[4185];
assign g[8282] = a[12] & g[4186];
assign g[12377] = b[12] & g[4186];
assign g[8283] = a[12] & g[4187];
assign g[12378] = b[12] & g[4187];
assign g[8284] = a[12] & g[4188];
assign g[12379] = b[12] & g[4188];
assign g[8285] = a[12] & g[4189];
assign g[12380] = b[12] & g[4189];
assign g[8286] = a[12] & g[4190];
assign g[12381] = b[12] & g[4190];
assign g[8287] = a[12] & g[4191];
assign g[12382] = b[12] & g[4191];
assign g[8288] = a[12] & g[4192];
assign g[12383] = b[12] & g[4192];
assign g[8289] = a[12] & g[4193];
assign g[12384] = b[12] & g[4193];
assign g[8290] = a[12] & g[4194];
assign g[12385] = b[12] & g[4194];
assign g[8291] = a[12] & g[4195];
assign g[12386] = b[12] & g[4195];
assign g[8292] = a[12] & g[4196];
assign g[12387] = b[12] & g[4196];
assign g[8293] = a[12] & g[4197];
assign g[12388] = b[12] & g[4197];
assign g[8294] = a[12] & g[4198];
assign g[12389] = b[12] & g[4198];
assign g[8295] = a[12] & g[4199];
assign g[12390] = b[12] & g[4199];
assign g[8296] = a[12] & g[4200];
assign g[12391] = b[12] & g[4200];
assign g[8297] = a[12] & g[4201];
assign g[12392] = b[12] & g[4201];
assign g[8298] = a[12] & g[4202];
assign g[12393] = b[12] & g[4202];
assign g[8299] = a[12] & g[4203];
assign g[12394] = b[12] & g[4203];
assign g[8300] = a[12] & g[4204];
assign g[12395] = b[12] & g[4204];
assign g[8301] = a[12] & g[4205];
assign g[12396] = b[12] & g[4205];
assign g[8302] = a[12] & g[4206];
assign g[12397] = b[12] & g[4206];
assign g[8303] = a[12] & g[4207];
assign g[12398] = b[12] & g[4207];
assign g[8304] = a[12] & g[4208];
assign g[12399] = b[12] & g[4208];
assign g[8305] = a[12] & g[4209];
assign g[12400] = b[12] & g[4209];
assign g[8306] = a[12] & g[4210];
assign g[12401] = b[12] & g[4210];
assign g[8307] = a[12] & g[4211];
assign g[12402] = b[12] & g[4211];
assign g[8308] = a[12] & g[4212];
assign g[12403] = b[12] & g[4212];
assign g[8309] = a[12] & g[4213];
assign g[12404] = b[12] & g[4213];
assign g[8310] = a[12] & g[4214];
assign g[12405] = b[12] & g[4214];
assign g[8311] = a[12] & g[4215];
assign g[12406] = b[12] & g[4215];
assign g[8312] = a[12] & g[4216];
assign g[12407] = b[12] & g[4216];
assign g[8313] = a[12] & g[4217];
assign g[12408] = b[12] & g[4217];
assign g[8314] = a[12] & g[4218];
assign g[12409] = b[12] & g[4218];
assign g[8315] = a[12] & g[4219];
assign g[12410] = b[12] & g[4219];
assign g[8316] = a[12] & g[4220];
assign g[12411] = b[12] & g[4220];
assign g[8317] = a[12] & g[4221];
assign g[12412] = b[12] & g[4221];
assign g[8318] = a[12] & g[4222];
assign g[12413] = b[12] & g[4222];
assign g[8319] = a[12] & g[4223];
assign g[12414] = b[12] & g[4223];
assign g[8320] = a[12] & g[4224];
assign g[12415] = b[12] & g[4224];
assign g[8321] = a[12] & g[4225];
assign g[12416] = b[12] & g[4225];
assign g[8322] = a[12] & g[4226];
assign g[12417] = b[12] & g[4226];
assign g[8323] = a[12] & g[4227];
assign g[12418] = b[12] & g[4227];
assign g[8324] = a[12] & g[4228];
assign g[12419] = b[12] & g[4228];
assign g[8325] = a[12] & g[4229];
assign g[12420] = b[12] & g[4229];
assign g[8326] = a[12] & g[4230];
assign g[12421] = b[12] & g[4230];
assign g[8327] = a[12] & g[4231];
assign g[12422] = b[12] & g[4231];
assign g[8328] = a[12] & g[4232];
assign g[12423] = b[12] & g[4232];
assign g[8329] = a[12] & g[4233];
assign g[12424] = b[12] & g[4233];
assign g[8330] = a[12] & g[4234];
assign g[12425] = b[12] & g[4234];
assign g[8331] = a[12] & g[4235];
assign g[12426] = b[12] & g[4235];
assign g[8332] = a[12] & g[4236];
assign g[12427] = b[12] & g[4236];
assign g[8333] = a[12] & g[4237];
assign g[12428] = b[12] & g[4237];
assign g[8334] = a[12] & g[4238];
assign g[12429] = b[12] & g[4238];
assign g[8335] = a[12] & g[4239];
assign g[12430] = b[12] & g[4239];
assign g[8336] = a[12] & g[4240];
assign g[12431] = b[12] & g[4240];
assign g[8337] = a[12] & g[4241];
assign g[12432] = b[12] & g[4241];
assign g[8338] = a[12] & g[4242];
assign g[12433] = b[12] & g[4242];
assign g[8339] = a[12] & g[4243];
assign g[12434] = b[12] & g[4243];
assign g[8340] = a[12] & g[4244];
assign g[12435] = b[12] & g[4244];
assign g[8341] = a[12] & g[4245];
assign g[12436] = b[12] & g[4245];
assign g[8342] = a[12] & g[4246];
assign g[12437] = b[12] & g[4246];
assign g[8343] = a[12] & g[4247];
assign g[12438] = b[12] & g[4247];
assign g[8344] = a[12] & g[4248];
assign g[12439] = b[12] & g[4248];
assign g[8345] = a[12] & g[4249];
assign g[12440] = b[12] & g[4249];
assign g[8346] = a[12] & g[4250];
assign g[12441] = b[12] & g[4250];
assign g[8347] = a[12] & g[4251];
assign g[12442] = b[12] & g[4251];
assign g[8348] = a[12] & g[4252];
assign g[12443] = b[12] & g[4252];
assign g[8349] = a[12] & g[4253];
assign g[12444] = b[12] & g[4253];
assign g[8350] = a[12] & g[4254];
assign g[12445] = b[12] & g[4254];
assign g[8351] = a[12] & g[4255];
assign g[12446] = b[12] & g[4255];
assign g[8352] = a[12] & g[4256];
assign g[12447] = b[12] & g[4256];
assign g[8353] = a[12] & g[4257];
assign g[12448] = b[12] & g[4257];
assign g[8354] = a[12] & g[4258];
assign g[12449] = b[12] & g[4258];
assign g[8355] = a[12] & g[4259];
assign g[12450] = b[12] & g[4259];
assign g[8356] = a[12] & g[4260];
assign g[12451] = b[12] & g[4260];
assign g[8357] = a[12] & g[4261];
assign g[12452] = b[12] & g[4261];
assign g[8358] = a[12] & g[4262];
assign g[12453] = b[12] & g[4262];
assign g[8359] = a[12] & g[4263];
assign g[12454] = b[12] & g[4263];
assign g[8360] = a[12] & g[4264];
assign g[12455] = b[12] & g[4264];
assign g[8361] = a[12] & g[4265];
assign g[12456] = b[12] & g[4265];
assign g[8362] = a[12] & g[4266];
assign g[12457] = b[12] & g[4266];
assign g[8363] = a[12] & g[4267];
assign g[12458] = b[12] & g[4267];
assign g[8364] = a[12] & g[4268];
assign g[12459] = b[12] & g[4268];
assign g[8365] = a[12] & g[4269];
assign g[12460] = b[12] & g[4269];
assign g[8366] = a[12] & g[4270];
assign g[12461] = b[12] & g[4270];
assign g[8367] = a[12] & g[4271];
assign g[12462] = b[12] & g[4271];
assign g[8368] = a[12] & g[4272];
assign g[12463] = b[12] & g[4272];
assign g[8369] = a[12] & g[4273];
assign g[12464] = b[12] & g[4273];
assign g[8370] = a[12] & g[4274];
assign g[12465] = b[12] & g[4274];
assign g[8371] = a[12] & g[4275];
assign g[12466] = b[12] & g[4275];
assign g[8372] = a[12] & g[4276];
assign g[12467] = b[12] & g[4276];
assign g[8373] = a[12] & g[4277];
assign g[12468] = b[12] & g[4277];
assign g[8374] = a[12] & g[4278];
assign g[12469] = b[12] & g[4278];
assign g[8375] = a[12] & g[4279];
assign g[12470] = b[12] & g[4279];
assign g[8376] = a[12] & g[4280];
assign g[12471] = b[12] & g[4280];
assign g[8377] = a[12] & g[4281];
assign g[12472] = b[12] & g[4281];
assign g[8378] = a[12] & g[4282];
assign g[12473] = b[12] & g[4282];
assign g[8379] = a[12] & g[4283];
assign g[12474] = b[12] & g[4283];
assign g[8380] = a[12] & g[4284];
assign g[12475] = b[12] & g[4284];
assign g[8381] = a[12] & g[4285];
assign g[12476] = b[12] & g[4285];
assign g[8382] = a[12] & g[4286];
assign g[12477] = b[12] & g[4286];
assign g[8383] = a[12] & g[4287];
assign g[12478] = b[12] & g[4287];
assign g[8384] = a[12] & g[4288];
assign g[12479] = b[12] & g[4288];
assign g[8385] = a[12] & g[4289];
assign g[12480] = b[12] & g[4289];
assign g[8386] = a[12] & g[4290];
assign g[12481] = b[12] & g[4290];
assign g[8387] = a[12] & g[4291];
assign g[12482] = b[12] & g[4291];
assign g[8388] = a[12] & g[4292];
assign g[12483] = b[12] & g[4292];
assign g[8389] = a[12] & g[4293];
assign g[12484] = b[12] & g[4293];
assign g[8390] = a[12] & g[4294];
assign g[12485] = b[12] & g[4294];
assign g[8391] = a[12] & g[4295];
assign g[12486] = b[12] & g[4295];
assign g[8392] = a[12] & g[4296];
assign g[12487] = b[12] & g[4296];
assign g[8393] = a[12] & g[4297];
assign g[12488] = b[12] & g[4297];
assign g[8394] = a[12] & g[4298];
assign g[12489] = b[12] & g[4298];
assign g[8395] = a[12] & g[4299];
assign g[12490] = b[12] & g[4299];
assign g[8396] = a[12] & g[4300];
assign g[12491] = b[12] & g[4300];
assign g[8397] = a[12] & g[4301];
assign g[12492] = b[12] & g[4301];
assign g[8398] = a[12] & g[4302];
assign g[12493] = b[12] & g[4302];
assign g[8399] = a[12] & g[4303];
assign g[12494] = b[12] & g[4303];
assign g[8400] = a[12] & g[4304];
assign g[12495] = b[12] & g[4304];
assign g[8401] = a[12] & g[4305];
assign g[12496] = b[12] & g[4305];
assign g[8402] = a[12] & g[4306];
assign g[12497] = b[12] & g[4306];
assign g[8403] = a[12] & g[4307];
assign g[12498] = b[12] & g[4307];
assign g[8404] = a[12] & g[4308];
assign g[12499] = b[12] & g[4308];
assign g[8405] = a[12] & g[4309];
assign g[12500] = b[12] & g[4309];
assign g[8406] = a[12] & g[4310];
assign g[12501] = b[12] & g[4310];
assign g[8407] = a[12] & g[4311];
assign g[12502] = b[12] & g[4311];
assign g[8408] = a[12] & g[4312];
assign g[12503] = b[12] & g[4312];
assign g[8409] = a[12] & g[4313];
assign g[12504] = b[12] & g[4313];
assign g[8410] = a[12] & g[4314];
assign g[12505] = b[12] & g[4314];
assign g[8411] = a[12] & g[4315];
assign g[12506] = b[12] & g[4315];
assign g[8412] = a[12] & g[4316];
assign g[12507] = b[12] & g[4316];
assign g[8413] = a[12] & g[4317];
assign g[12508] = b[12] & g[4317];
assign g[8414] = a[12] & g[4318];
assign g[12509] = b[12] & g[4318];
assign g[8415] = a[12] & g[4319];
assign g[12510] = b[12] & g[4319];
assign g[8416] = a[12] & g[4320];
assign g[12511] = b[12] & g[4320];
assign g[8417] = a[12] & g[4321];
assign g[12512] = b[12] & g[4321];
assign g[8418] = a[12] & g[4322];
assign g[12513] = b[12] & g[4322];
assign g[8419] = a[12] & g[4323];
assign g[12514] = b[12] & g[4323];
assign g[8420] = a[12] & g[4324];
assign g[12515] = b[12] & g[4324];
assign g[8421] = a[12] & g[4325];
assign g[12516] = b[12] & g[4325];
assign g[8422] = a[12] & g[4326];
assign g[12517] = b[12] & g[4326];
assign g[8423] = a[12] & g[4327];
assign g[12518] = b[12] & g[4327];
assign g[8424] = a[12] & g[4328];
assign g[12519] = b[12] & g[4328];
assign g[8425] = a[12] & g[4329];
assign g[12520] = b[12] & g[4329];
assign g[8426] = a[12] & g[4330];
assign g[12521] = b[12] & g[4330];
assign g[8427] = a[12] & g[4331];
assign g[12522] = b[12] & g[4331];
assign g[8428] = a[12] & g[4332];
assign g[12523] = b[12] & g[4332];
assign g[8429] = a[12] & g[4333];
assign g[12524] = b[12] & g[4333];
assign g[8430] = a[12] & g[4334];
assign g[12525] = b[12] & g[4334];
assign g[8431] = a[12] & g[4335];
assign g[12526] = b[12] & g[4335];
assign g[8432] = a[12] & g[4336];
assign g[12527] = b[12] & g[4336];
assign g[8433] = a[12] & g[4337];
assign g[12528] = b[12] & g[4337];
assign g[8434] = a[12] & g[4338];
assign g[12529] = b[12] & g[4338];
assign g[8435] = a[12] & g[4339];
assign g[12530] = b[12] & g[4339];
assign g[8436] = a[12] & g[4340];
assign g[12531] = b[12] & g[4340];
assign g[8437] = a[12] & g[4341];
assign g[12532] = b[12] & g[4341];
assign g[8438] = a[12] & g[4342];
assign g[12533] = b[12] & g[4342];
assign g[8439] = a[12] & g[4343];
assign g[12534] = b[12] & g[4343];
assign g[8440] = a[12] & g[4344];
assign g[12535] = b[12] & g[4344];
assign g[8441] = a[12] & g[4345];
assign g[12536] = b[12] & g[4345];
assign g[8442] = a[12] & g[4346];
assign g[12537] = b[12] & g[4346];
assign g[8443] = a[12] & g[4347];
assign g[12538] = b[12] & g[4347];
assign g[8444] = a[12] & g[4348];
assign g[12539] = b[12] & g[4348];
assign g[8445] = a[12] & g[4349];
assign g[12540] = b[12] & g[4349];
assign g[8446] = a[12] & g[4350];
assign g[12541] = b[12] & g[4350];
assign g[8447] = a[12] & g[4351];
assign g[12542] = b[12] & g[4351];
assign g[8448] = a[12] & g[4352];
assign g[12543] = b[12] & g[4352];
assign g[8449] = a[12] & g[4353];
assign g[12544] = b[12] & g[4353];
assign g[8450] = a[12] & g[4354];
assign g[12545] = b[12] & g[4354];
assign g[8451] = a[12] & g[4355];
assign g[12546] = b[12] & g[4355];
assign g[8452] = a[12] & g[4356];
assign g[12547] = b[12] & g[4356];
assign g[8453] = a[12] & g[4357];
assign g[12548] = b[12] & g[4357];
assign g[8454] = a[12] & g[4358];
assign g[12549] = b[12] & g[4358];
assign g[8455] = a[12] & g[4359];
assign g[12550] = b[12] & g[4359];
assign g[8456] = a[12] & g[4360];
assign g[12551] = b[12] & g[4360];
assign g[8457] = a[12] & g[4361];
assign g[12552] = b[12] & g[4361];
assign g[8458] = a[12] & g[4362];
assign g[12553] = b[12] & g[4362];
assign g[8459] = a[12] & g[4363];
assign g[12554] = b[12] & g[4363];
assign g[8460] = a[12] & g[4364];
assign g[12555] = b[12] & g[4364];
assign g[8461] = a[12] & g[4365];
assign g[12556] = b[12] & g[4365];
assign g[8462] = a[12] & g[4366];
assign g[12557] = b[12] & g[4366];
assign g[8463] = a[12] & g[4367];
assign g[12558] = b[12] & g[4367];
assign g[8464] = a[12] & g[4368];
assign g[12559] = b[12] & g[4368];
assign g[8465] = a[12] & g[4369];
assign g[12560] = b[12] & g[4369];
assign g[8466] = a[12] & g[4370];
assign g[12561] = b[12] & g[4370];
assign g[8467] = a[12] & g[4371];
assign g[12562] = b[12] & g[4371];
assign g[8468] = a[12] & g[4372];
assign g[12563] = b[12] & g[4372];
assign g[8469] = a[12] & g[4373];
assign g[12564] = b[12] & g[4373];
assign g[8470] = a[12] & g[4374];
assign g[12565] = b[12] & g[4374];
assign g[8471] = a[12] & g[4375];
assign g[12566] = b[12] & g[4375];
assign g[8472] = a[12] & g[4376];
assign g[12567] = b[12] & g[4376];
assign g[8473] = a[12] & g[4377];
assign g[12568] = b[12] & g[4377];
assign g[8474] = a[12] & g[4378];
assign g[12569] = b[12] & g[4378];
assign g[8475] = a[12] & g[4379];
assign g[12570] = b[12] & g[4379];
assign g[8476] = a[12] & g[4380];
assign g[12571] = b[12] & g[4380];
assign g[8477] = a[12] & g[4381];
assign g[12572] = b[12] & g[4381];
assign g[8478] = a[12] & g[4382];
assign g[12573] = b[12] & g[4382];
assign g[8479] = a[12] & g[4383];
assign g[12574] = b[12] & g[4383];
assign g[8480] = a[12] & g[4384];
assign g[12575] = b[12] & g[4384];
assign g[8481] = a[12] & g[4385];
assign g[12576] = b[12] & g[4385];
assign g[8482] = a[12] & g[4386];
assign g[12577] = b[12] & g[4386];
assign g[8483] = a[12] & g[4387];
assign g[12578] = b[12] & g[4387];
assign g[8484] = a[12] & g[4388];
assign g[12579] = b[12] & g[4388];
assign g[8485] = a[12] & g[4389];
assign g[12580] = b[12] & g[4389];
assign g[8486] = a[12] & g[4390];
assign g[12581] = b[12] & g[4390];
assign g[8487] = a[12] & g[4391];
assign g[12582] = b[12] & g[4391];
assign g[8488] = a[12] & g[4392];
assign g[12583] = b[12] & g[4392];
assign g[8489] = a[12] & g[4393];
assign g[12584] = b[12] & g[4393];
assign g[8490] = a[12] & g[4394];
assign g[12585] = b[12] & g[4394];
assign g[8491] = a[12] & g[4395];
assign g[12586] = b[12] & g[4395];
assign g[8492] = a[12] & g[4396];
assign g[12587] = b[12] & g[4396];
assign g[8493] = a[12] & g[4397];
assign g[12588] = b[12] & g[4397];
assign g[8494] = a[12] & g[4398];
assign g[12589] = b[12] & g[4398];
assign g[8495] = a[12] & g[4399];
assign g[12590] = b[12] & g[4399];
assign g[8496] = a[12] & g[4400];
assign g[12591] = b[12] & g[4400];
assign g[8497] = a[12] & g[4401];
assign g[12592] = b[12] & g[4401];
assign g[8498] = a[12] & g[4402];
assign g[12593] = b[12] & g[4402];
assign g[8499] = a[12] & g[4403];
assign g[12594] = b[12] & g[4403];
assign g[8500] = a[12] & g[4404];
assign g[12595] = b[12] & g[4404];
assign g[8501] = a[12] & g[4405];
assign g[12596] = b[12] & g[4405];
assign g[8502] = a[12] & g[4406];
assign g[12597] = b[12] & g[4406];
assign g[8503] = a[12] & g[4407];
assign g[12598] = b[12] & g[4407];
assign g[8504] = a[12] & g[4408];
assign g[12599] = b[12] & g[4408];
assign g[8505] = a[12] & g[4409];
assign g[12600] = b[12] & g[4409];
assign g[8506] = a[12] & g[4410];
assign g[12601] = b[12] & g[4410];
assign g[8507] = a[12] & g[4411];
assign g[12602] = b[12] & g[4411];
assign g[8508] = a[12] & g[4412];
assign g[12603] = b[12] & g[4412];
assign g[8509] = a[12] & g[4413];
assign g[12604] = b[12] & g[4413];
assign g[8510] = a[12] & g[4414];
assign g[12605] = b[12] & g[4414];
assign g[8511] = a[12] & g[4415];
assign g[12606] = b[12] & g[4415];
assign g[8512] = a[12] & g[4416];
assign g[12607] = b[12] & g[4416];
assign g[8513] = a[12] & g[4417];
assign g[12608] = b[12] & g[4417];
assign g[8514] = a[12] & g[4418];
assign g[12609] = b[12] & g[4418];
assign g[8515] = a[12] & g[4419];
assign g[12610] = b[12] & g[4419];
assign g[8516] = a[12] & g[4420];
assign g[12611] = b[12] & g[4420];
assign g[8517] = a[12] & g[4421];
assign g[12612] = b[12] & g[4421];
assign g[8518] = a[12] & g[4422];
assign g[12613] = b[12] & g[4422];
assign g[8519] = a[12] & g[4423];
assign g[12614] = b[12] & g[4423];
assign g[8520] = a[12] & g[4424];
assign g[12615] = b[12] & g[4424];
assign g[8521] = a[12] & g[4425];
assign g[12616] = b[12] & g[4425];
assign g[8522] = a[12] & g[4426];
assign g[12617] = b[12] & g[4426];
assign g[8523] = a[12] & g[4427];
assign g[12618] = b[12] & g[4427];
assign g[8524] = a[12] & g[4428];
assign g[12619] = b[12] & g[4428];
assign g[8525] = a[12] & g[4429];
assign g[12620] = b[12] & g[4429];
assign g[8526] = a[12] & g[4430];
assign g[12621] = b[12] & g[4430];
assign g[8527] = a[12] & g[4431];
assign g[12622] = b[12] & g[4431];
assign g[8528] = a[12] & g[4432];
assign g[12623] = b[12] & g[4432];
assign g[8529] = a[12] & g[4433];
assign g[12624] = b[12] & g[4433];
assign g[8530] = a[12] & g[4434];
assign g[12625] = b[12] & g[4434];
assign g[8531] = a[12] & g[4435];
assign g[12626] = b[12] & g[4435];
assign g[8532] = a[12] & g[4436];
assign g[12627] = b[12] & g[4436];
assign g[8533] = a[12] & g[4437];
assign g[12628] = b[12] & g[4437];
assign g[8534] = a[12] & g[4438];
assign g[12629] = b[12] & g[4438];
assign g[8535] = a[12] & g[4439];
assign g[12630] = b[12] & g[4439];
assign g[8536] = a[12] & g[4440];
assign g[12631] = b[12] & g[4440];
assign g[8537] = a[12] & g[4441];
assign g[12632] = b[12] & g[4441];
assign g[8538] = a[12] & g[4442];
assign g[12633] = b[12] & g[4442];
assign g[8539] = a[12] & g[4443];
assign g[12634] = b[12] & g[4443];
assign g[8540] = a[12] & g[4444];
assign g[12635] = b[12] & g[4444];
assign g[8541] = a[12] & g[4445];
assign g[12636] = b[12] & g[4445];
assign g[8542] = a[12] & g[4446];
assign g[12637] = b[12] & g[4446];
assign g[8543] = a[12] & g[4447];
assign g[12638] = b[12] & g[4447];
assign g[8544] = a[12] & g[4448];
assign g[12639] = b[12] & g[4448];
assign g[8545] = a[12] & g[4449];
assign g[12640] = b[12] & g[4449];
assign g[8546] = a[12] & g[4450];
assign g[12641] = b[12] & g[4450];
assign g[8547] = a[12] & g[4451];
assign g[12642] = b[12] & g[4451];
assign g[8548] = a[12] & g[4452];
assign g[12643] = b[12] & g[4452];
assign g[8549] = a[12] & g[4453];
assign g[12644] = b[12] & g[4453];
assign g[8550] = a[12] & g[4454];
assign g[12645] = b[12] & g[4454];
assign g[8551] = a[12] & g[4455];
assign g[12646] = b[12] & g[4455];
assign g[8552] = a[12] & g[4456];
assign g[12647] = b[12] & g[4456];
assign g[8553] = a[12] & g[4457];
assign g[12648] = b[12] & g[4457];
assign g[8554] = a[12] & g[4458];
assign g[12649] = b[12] & g[4458];
assign g[8555] = a[12] & g[4459];
assign g[12650] = b[12] & g[4459];
assign g[8556] = a[12] & g[4460];
assign g[12651] = b[12] & g[4460];
assign g[8557] = a[12] & g[4461];
assign g[12652] = b[12] & g[4461];
assign g[8558] = a[12] & g[4462];
assign g[12653] = b[12] & g[4462];
assign g[8559] = a[12] & g[4463];
assign g[12654] = b[12] & g[4463];
assign g[8560] = a[12] & g[4464];
assign g[12655] = b[12] & g[4464];
assign g[8561] = a[12] & g[4465];
assign g[12656] = b[12] & g[4465];
assign g[8562] = a[12] & g[4466];
assign g[12657] = b[12] & g[4466];
assign g[8563] = a[12] & g[4467];
assign g[12658] = b[12] & g[4467];
assign g[8564] = a[12] & g[4468];
assign g[12659] = b[12] & g[4468];
assign g[8565] = a[12] & g[4469];
assign g[12660] = b[12] & g[4469];
assign g[8566] = a[12] & g[4470];
assign g[12661] = b[12] & g[4470];
assign g[8567] = a[12] & g[4471];
assign g[12662] = b[12] & g[4471];
assign g[8568] = a[12] & g[4472];
assign g[12663] = b[12] & g[4472];
assign g[8569] = a[12] & g[4473];
assign g[12664] = b[12] & g[4473];
assign g[8570] = a[12] & g[4474];
assign g[12665] = b[12] & g[4474];
assign g[8571] = a[12] & g[4475];
assign g[12666] = b[12] & g[4475];
assign g[8572] = a[12] & g[4476];
assign g[12667] = b[12] & g[4476];
assign g[8573] = a[12] & g[4477];
assign g[12668] = b[12] & g[4477];
assign g[8574] = a[12] & g[4478];
assign g[12669] = b[12] & g[4478];
assign g[8575] = a[12] & g[4479];
assign g[12670] = b[12] & g[4479];
assign g[8576] = a[12] & g[4480];
assign g[12671] = b[12] & g[4480];
assign g[8577] = a[12] & g[4481];
assign g[12672] = b[12] & g[4481];
assign g[8578] = a[12] & g[4482];
assign g[12673] = b[12] & g[4482];
assign g[8579] = a[12] & g[4483];
assign g[12674] = b[12] & g[4483];
assign g[8580] = a[12] & g[4484];
assign g[12675] = b[12] & g[4484];
assign g[8581] = a[12] & g[4485];
assign g[12676] = b[12] & g[4485];
assign g[8582] = a[12] & g[4486];
assign g[12677] = b[12] & g[4486];
assign g[8583] = a[12] & g[4487];
assign g[12678] = b[12] & g[4487];
assign g[8584] = a[12] & g[4488];
assign g[12679] = b[12] & g[4488];
assign g[8585] = a[12] & g[4489];
assign g[12680] = b[12] & g[4489];
assign g[8586] = a[12] & g[4490];
assign g[12681] = b[12] & g[4490];
assign g[8587] = a[12] & g[4491];
assign g[12682] = b[12] & g[4491];
assign g[8588] = a[12] & g[4492];
assign g[12683] = b[12] & g[4492];
assign g[8589] = a[12] & g[4493];
assign g[12684] = b[12] & g[4493];
assign g[8590] = a[12] & g[4494];
assign g[12685] = b[12] & g[4494];
assign g[8591] = a[12] & g[4495];
assign g[12686] = b[12] & g[4495];
assign g[8592] = a[12] & g[4496];
assign g[12687] = b[12] & g[4496];
assign g[8593] = a[12] & g[4497];
assign g[12688] = b[12] & g[4497];
assign g[8594] = a[12] & g[4498];
assign g[12689] = b[12] & g[4498];
assign g[8595] = a[12] & g[4499];
assign g[12690] = b[12] & g[4499];
assign g[8596] = a[12] & g[4500];
assign g[12691] = b[12] & g[4500];
assign g[8597] = a[12] & g[4501];
assign g[12692] = b[12] & g[4501];
assign g[8598] = a[12] & g[4502];
assign g[12693] = b[12] & g[4502];
assign g[8599] = a[12] & g[4503];
assign g[12694] = b[12] & g[4503];
assign g[8600] = a[12] & g[4504];
assign g[12695] = b[12] & g[4504];
assign g[8601] = a[12] & g[4505];
assign g[12696] = b[12] & g[4505];
assign g[8602] = a[12] & g[4506];
assign g[12697] = b[12] & g[4506];
assign g[8603] = a[12] & g[4507];
assign g[12698] = b[12] & g[4507];
assign g[8604] = a[12] & g[4508];
assign g[12699] = b[12] & g[4508];
assign g[8605] = a[12] & g[4509];
assign g[12700] = b[12] & g[4509];
assign g[8606] = a[12] & g[4510];
assign g[12701] = b[12] & g[4510];
assign g[8607] = a[12] & g[4511];
assign g[12702] = b[12] & g[4511];
assign g[8608] = a[12] & g[4512];
assign g[12703] = b[12] & g[4512];
assign g[8609] = a[12] & g[4513];
assign g[12704] = b[12] & g[4513];
assign g[8610] = a[12] & g[4514];
assign g[12705] = b[12] & g[4514];
assign g[8611] = a[12] & g[4515];
assign g[12706] = b[12] & g[4515];
assign g[8612] = a[12] & g[4516];
assign g[12707] = b[12] & g[4516];
assign g[8613] = a[12] & g[4517];
assign g[12708] = b[12] & g[4517];
assign g[8614] = a[12] & g[4518];
assign g[12709] = b[12] & g[4518];
assign g[8615] = a[12] & g[4519];
assign g[12710] = b[12] & g[4519];
assign g[8616] = a[12] & g[4520];
assign g[12711] = b[12] & g[4520];
assign g[8617] = a[12] & g[4521];
assign g[12712] = b[12] & g[4521];
assign g[8618] = a[12] & g[4522];
assign g[12713] = b[12] & g[4522];
assign g[8619] = a[12] & g[4523];
assign g[12714] = b[12] & g[4523];
assign g[8620] = a[12] & g[4524];
assign g[12715] = b[12] & g[4524];
assign g[8621] = a[12] & g[4525];
assign g[12716] = b[12] & g[4525];
assign g[8622] = a[12] & g[4526];
assign g[12717] = b[12] & g[4526];
assign g[8623] = a[12] & g[4527];
assign g[12718] = b[12] & g[4527];
assign g[8624] = a[12] & g[4528];
assign g[12719] = b[12] & g[4528];
assign g[8625] = a[12] & g[4529];
assign g[12720] = b[12] & g[4529];
assign g[8626] = a[12] & g[4530];
assign g[12721] = b[12] & g[4530];
assign g[8627] = a[12] & g[4531];
assign g[12722] = b[12] & g[4531];
assign g[8628] = a[12] & g[4532];
assign g[12723] = b[12] & g[4532];
assign g[8629] = a[12] & g[4533];
assign g[12724] = b[12] & g[4533];
assign g[8630] = a[12] & g[4534];
assign g[12725] = b[12] & g[4534];
assign g[8631] = a[12] & g[4535];
assign g[12726] = b[12] & g[4535];
assign g[8632] = a[12] & g[4536];
assign g[12727] = b[12] & g[4536];
assign g[8633] = a[12] & g[4537];
assign g[12728] = b[12] & g[4537];
assign g[8634] = a[12] & g[4538];
assign g[12729] = b[12] & g[4538];
assign g[8635] = a[12] & g[4539];
assign g[12730] = b[12] & g[4539];
assign g[8636] = a[12] & g[4540];
assign g[12731] = b[12] & g[4540];
assign g[8637] = a[12] & g[4541];
assign g[12732] = b[12] & g[4541];
assign g[8638] = a[12] & g[4542];
assign g[12733] = b[12] & g[4542];
assign g[8639] = a[12] & g[4543];
assign g[12734] = b[12] & g[4543];
assign g[8640] = a[12] & g[4544];
assign g[12735] = b[12] & g[4544];
assign g[8641] = a[12] & g[4545];
assign g[12736] = b[12] & g[4545];
assign g[8642] = a[12] & g[4546];
assign g[12737] = b[12] & g[4546];
assign g[8643] = a[12] & g[4547];
assign g[12738] = b[12] & g[4547];
assign g[8644] = a[12] & g[4548];
assign g[12739] = b[12] & g[4548];
assign g[8645] = a[12] & g[4549];
assign g[12740] = b[12] & g[4549];
assign g[8646] = a[12] & g[4550];
assign g[12741] = b[12] & g[4550];
assign g[8647] = a[12] & g[4551];
assign g[12742] = b[12] & g[4551];
assign g[8648] = a[12] & g[4552];
assign g[12743] = b[12] & g[4552];
assign g[8649] = a[12] & g[4553];
assign g[12744] = b[12] & g[4553];
assign g[8650] = a[12] & g[4554];
assign g[12745] = b[12] & g[4554];
assign g[8651] = a[12] & g[4555];
assign g[12746] = b[12] & g[4555];
assign g[8652] = a[12] & g[4556];
assign g[12747] = b[12] & g[4556];
assign g[8653] = a[12] & g[4557];
assign g[12748] = b[12] & g[4557];
assign g[8654] = a[12] & g[4558];
assign g[12749] = b[12] & g[4558];
assign g[8655] = a[12] & g[4559];
assign g[12750] = b[12] & g[4559];
assign g[8656] = a[12] & g[4560];
assign g[12751] = b[12] & g[4560];
assign g[8657] = a[12] & g[4561];
assign g[12752] = b[12] & g[4561];
assign g[8658] = a[12] & g[4562];
assign g[12753] = b[12] & g[4562];
assign g[8659] = a[12] & g[4563];
assign g[12754] = b[12] & g[4563];
assign g[8660] = a[12] & g[4564];
assign g[12755] = b[12] & g[4564];
assign g[8661] = a[12] & g[4565];
assign g[12756] = b[12] & g[4565];
assign g[8662] = a[12] & g[4566];
assign g[12757] = b[12] & g[4566];
assign g[8663] = a[12] & g[4567];
assign g[12758] = b[12] & g[4567];
assign g[8664] = a[12] & g[4568];
assign g[12759] = b[12] & g[4568];
assign g[8665] = a[12] & g[4569];
assign g[12760] = b[12] & g[4569];
assign g[8666] = a[12] & g[4570];
assign g[12761] = b[12] & g[4570];
assign g[8667] = a[12] & g[4571];
assign g[12762] = b[12] & g[4571];
assign g[8668] = a[12] & g[4572];
assign g[12763] = b[12] & g[4572];
assign g[8669] = a[12] & g[4573];
assign g[12764] = b[12] & g[4573];
assign g[8670] = a[12] & g[4574];
assign g[12765] = b[12] & g[4574];
assign g[8671] = a[12] & g[4575];
assign g[12766] = b[12] & g[4575];
assign g[8672] = a[12] & g[4576];
assign g[12767] = b[12] & g[4576];
assign g[8673] = a[12] & g[4577];
assign g[12768] = b[12] & g[4577];
assign g[8674] = a[12] & g[4578];
assign g[12769] = b[12] & g[4578];
assign g[8675] = a[12] & g[4579];
assign g[12770] = b[12] & g[4579];
assign g[8676] = a[12] & g[4580];
assign g[12771] = b[12] & g[4580];
assign g[8677] = a[12] & g[4581];
assign g[12772] = b[12] & g[4581];
assign g[8678] = a[12] & g[4582];
assign g[12773] = b[12] & g[4582];
assign g[8679] = a[12] & g[4583];
assign g[12774] = b[12] & g[4583];
assign g[8680] = a[12] & g[4584];
assign g[12775] = b[12] & g[4584];
assign g[8681] = a[12] & g[4585];
assign g[12776] = b[12] & g[4585];
assign g[8682] = a[12] & g[4586];
assign g[12777] = b[12] & g[4586];
assign g[8683] = a[12] & g[4587];
assign g[12778] = b[12] & g[4587];
assign g[8684] = a[12] & g[4588];
assign g[12779] = b[12] & g[4588];
assign g[8685] = a[12] & g[4589];
assign g[12780] = b[12] & g[4589];
assign g[8686] = a[12] & g[4590];
assign g[12781] = b[12] & g[4590];
assign g[8687] = a[12] & g[4591];
assign g[12782] = b[12] & g[4591];
assign g[8688] = a[12] & g[4592];
assign g[12783] = b[12] & g[4592];
assign g[8689] = a[12] & g[4593];
assign g[12784] = b[12] & g[4593];
assign g[8690] = a[12] & g[4594];
assign g[12785] = b[12] & g[4594];
assign g[8691] = a[12] & g[4595];
assign g[12786] = b[12] & g[4595];
assign g[8692] = a[12] & g[4596];
assign g[12787] = b[12] & g[4596];
assign g[8693] = a[12] & g[4597];
assign g[12788] = b[12] & g[4597];
assign g[8694] = a[12] & g[4598];
assign g[12789] = b[12] & g[4598];
assign g[8695] = a[12] & g[4599];
assign g[12790] = b[12] & g[4599];
assign g[8696] = a[12] & g[4600];
assign g[12791] = b[12] & g[4600];
assign g[8697] = a[12] & g[4601];
assign g[12792] = b[12] & g[4601];
assign g[8698] = a[12] & g[4602];
assign g[12793] = b[12] & g[4602];
assign g[8699] = a[12] & g[4603];
assign g[12794] = b[12] & g[4603];
assign g[8700] = a[12] & g[4604];
assign g[12795] = b[12] & g[4604];
assign g[8701] = a[12] & g[4605];
assign g[12796] = b[12] & g[4605];
assign g[8702] = a[12] & g[4606];
assign g[12797] = b[12] & g[4606];
assign g[8703] = a[12] & g[4607];
assign g[12798] = b[12] & g[4607];
assign g[8704] = a[12] & g[4608];
assign g[12799] = b[12] & g[4608];
assign g[8705] = a[12] & g[4609];
assign g[12800] = b[12] & g[4609];
assign g[8706] = a[12] & g[4610];
assign g[12801] = b[12] & g[4610];
assign g[8707] = a[12] & g[4611];
assign g[12802] = b[12] & g[4611];
assign g[8708] = a[12] & g[4612];
assign g[12803] = b[12] & g[4612];
assign g[8709] = a[12] & g[4613];
assign g[12804] = b[12] & g[4613];
assign g[8710] = a[12] & g[4614];
assign g[12805] = b[12] & g[4614];
assign g[8711] = a[12] & g[4615];
assign g[12806] = b[12] & g[4615];
assign g[8712] = a[12] & g[4616];
assign g[12807] = b[12] & g[4616];
assign g[8713] = a[12] & g[4617];
assign g[12808] = b[12] & g[4617];
assign g[8714] = a[12] & g[4618];
assign g[12809] = b[12] & g[4618];
assign g[8715] = a[12] & g[4619];
assign g[12810] = b[12] & g[4619];
assign g[8716] = a[12] & g[4620];
assign g[12811] = b[12] & g[4620];
assign g[8717] = a[12] & g[4621];
assign g[12812] = b[12] & g[4621];
assign g[8718] = a[12] & g[4622];
assign g[12813] = b[12] & g[4622];
assign g[8719] = a[12] & g[4623];
assign g[12814] = b[12] & g[4623];
assign g[8720] = a[12] & g[4624];
assign g[12815] = b[12] & g[4624];
assign g[8721] = a[12] & g[4625];
assign g[12816] = b[12] & g[4625];
assign g[8722] = a[12] & g[4626];
assign g[12817] = b[12] & g[4626];
assign g[8723] = a[12] & g[4627];
assign g[12818] = b[12] & g[4627];
assign g[8724] = a[12] & g[4628];
assign g[12819] = b[12] & g[4628];
assign g[8725] = a[12] & g[4629];
assign g[12820] = b[12] & g[4629];
assign g[8726] = a[12] & g[4630];
assign g[12821] = b[12] & g[4630];
assign g[8727] = a[12] & g[4631];
assign g[12822] = b[12] & g[4631];
assign g[8728] = a[12] & g[4632];
assign g[12823] = b[12] & g[4632];
assign g[8729] = a[12] & g[4633];
assign g[12824] = b[12] & g[4633];
assign g[8730] = a[12] & g[4634];
assign g[12825] = b[12] & g[4634];
assign g[8731] = a[12] & g[4635];
assign g[12826] = b[12] & g[4635];
assign g[8732] = a[12] & g[4636];
assign g[12827] = b[12] & g[4636];
assign g[8733] = a[12] & g[4637];
assign g[12828] = b[12] & g[4637];
assign g[8734] = a[12] & g[4638];
assign g[12829] = b[12] & g[4638];
assign g[8735] = a[12] & g[4639];
assign g[12830] = b[12] & g[4639];
assign g[8736] = a[12] & g[4640];
assign g[12831] = b[12] & g[4640];
assign g[8737] = a[12] & g[4641];
assign g[12832] = b[12] & g[4641];
assign g[8738] = a[12] & g[4642];
assign g[12833] = b[12] & g[4642];
assign g[8739] = a[12] & g[4643];
assign g[12834] = b[12] & g[4643];
assign g[8740] = a[12] & g[4644];
assign g[12835] = b[12] & g[4644];
assign g[8741] = a[12] & g[4645];
assign g[12836] = b[12] & g[4645];
assign g[8742] = a[12] & g[4646];
assign g[12837] = b[12] & g[4646];
assign g[8743] = a[12] & g[4647];
assign g[12838] = b[12] & g[4647];
assign g[8744] = a[12] & g[4648];
assign g[12839] = b[12] & g[4648];
assign g[8745] = a[12] & g[4649];
assign g[12840] = b[12] & g[4649];
assign g[8746] = a[12] & g[4650];
assign g[12841] = b[12] & g[4650];
assign g[8747] = a[12] & g[4651];
assign g[12842] = b[12] & g[4651];
assign g[8748] = a[12] & g[4652];
assign g[12843] = b[12] & g[4652];
assign g[8749] = a[12] & g[4653];
assign g[12844] = b[12] & g[4653];
assign g[8750] = a[12] & g[4654];
assign g[12845] = b[12] & g[4654];
assign g[8751] = a[12] & g[4655];
assign g[12846] = b[12] & g[4655];
assign g[8752] = a[12] & g[4656];
assign g[12847] = b[12] & g[4656];
assign g[8753] = a[12] & g[4657];
assign g[12848] = b[12] & g[4657];
assign g[8754] = a[12] & g[4658];
assign g[12849] = b[12] & g[4658];
assign g[8755] = a[12] & g[4659];
assign g[12850] = b[12] & g[4659];
assign g[8756] = a[12] & g[4660];
assign g[12851] = b[12] & g[4660];
assign g[8757] = a[12] & g[4661];
assign g[12852] = b[12] & g[4661];
assign g[8758] = a[12] & g[4662];
assign g[12853] = b[12] & g[4662];
assign g[8759] = a[12] & g[4663];
assign g[12854] = b[12] & g[4663];
assign g[8760] = a[12] & g[4664];
assign g[12855] = b[12] & g[4664];
assign g[8761] = a[12] & g[4665];
assign g[12856] = b[12] & g[4665];
assign g[8762] = a[12] & g[4666];
assign g[12857] = b[12] & g[4666];
assign g[8763] = a[12] & g[4667];
assign g[12858] = b[12] & g[4667];
assign g[8764] = a[12] & g[4668];
assign g[12859] = b[12] & g[4668];
assign g[8765] = a[12] & g[4669];
assign g[12860] = b[12] & g[4669];
assign g[8766] = a[12] & g[4670];
assign g[12861] = b[12] & g[4670];
assign g[8767] = a[12] & g[4671];
assign g[12862] = b[12] & g[4671];
assign g[8768] = a[12] & g[4672];
assign g[12863] = b[12] & g[4672];
assign g[8769] = a[12] & g[4673];
assign g[12864] = b[12] & g[4673];
assign g[8770] = a[12] & g[4674];
assign g[12865] = b[12] & g[4674];
assign g[8771] = a[12] & g[4675];
assign g[12866] = b[12] & g[4675];
assign g[8772] = a[12] & g[4676];
assign g[12867] = b[12] & g[4676];
assign g[8773] = a[12] & g[4677];
assign g[12868] = b[12] & g[4677];
assign g[8774] = a[12] & g[4678];
assign g[12869] = b[12] & g[4678];
assign g[8775] = a[12] & g[4679];
assign g[12870] = b[12] & g[4679];
assign g[8776] = a[12] & g[4680];
assign g[12871] = b[12] & g[4680];
assign g[8777] = a[12] & g[4681];
assign g[12872] = b[12] & g[4681];
assign g[8778] = a[12] & g[4682];
assign g[12873] = b[12] & g[4682];
assign g[8779] = a[12] & g[4683];
assign g[12874] = b[12] & g[4683];
assign g[8780] = a[12] & g[4684];
assign g[12875] = b[12] & g[4684];
assign g[8781] = a[12] & g[4685];
assign g[12876] = b[12] & g[4685];
assign g[8782] = a[12] & g[4686];
assign g[12877] = b[12] & g[4686];
assign g[8783] = a[12] & g[4687];
assign g[12878] = b[12] & g[4687];
assign g[8784] = a[12] & g[4688];
assign g[12879] = b[12] & g[4688];
assign g[8785] = a[12] & g[4689];
assign g[12880] = b[12] & g[4689];
assign g[8786] = a[12] & g[4690];
assign g[12881] = b[12] & g[4690];
assign g[8787] = a[12] & g[4691];
assign g[12882] = b[12] & g[4691];
assign g[8788] = a[12] & g[4692];
assign g[12883] = b[12] & g[4692];
assign g[8789] = a[12] & g[4693];
assign g[12884] = b[12] & g[4693];
assign g[8790] = a[12] & g[4694];
assign g[12885] = b[12] & g[4694];
assign g[8791] = a[12] & g[4695];
assign g[12886] = b[12] & g[4695];
assign g[8792] = a[12] & g[4696];
assign g[12887] = b[12] & g[4696];
assign g[8793] = a[12] & g[4697];
assign g[12888] = b[12] & g[4697];
assign g[8794] = a[12] & g[4698];
assign g[12889] = b[12] & g[4698];
assign g[8795] = a[12] & g[4699];
assign g[12890] = b[12] & g[4699];
assign g[8796] = a[12] & g[4700];
assign g[12891] = b[12] & g[4700];
assign g[8797] = a[12] & g[4701];
assign g[12892] = b[12] & g[4701];
assign g[8798] = a[12] & g[4702];
assign g[12893] = b[12] & g[4702];
assign g[8799] = a[12] & g[4703];
assign g[12894] = b[12] & g[4703];
assign g[8800] = a[12] & g[4704];
assign g[12895] = b[12] & g[4704];
assign g[8801] = a[12] & g[4705];
assign g[12896] = b[12] & g[4705];
assign g[8802] = a[12] & g[4706];
assign g[12897] = b[12] & g[4706];
assign g[8803] = a[12] & g[4707];
assign g[12898] = b[12] & g[4707];
assign g[8804] = a[12] & g[4708];
assign g[12899] = b[12] & g[4708];
assign g[8805] = a[12] & g[4709];
assign g[12900] = b[12] & g[4709];
assign g[8806] = a[12] & g[4710];
assign g[12901] = b[12] & g[4710];
assign g[8807] = a[12] & g[4711];
assign g[12902] = b[12] & g[4711];
assign g[8808] = a[12] & g[4712];
assign g[12903] = b[12] & g[4712];
assign g[8809] = a[12] & g[4713];
assign g[12904] = b[12] & g[4713];
assign g[8810] = a[12] & g[4714];
assign g[12905] = b[12] & g[4714];
assign g[8811] = a[12] & g[4715];
assign g[12906] = b[12] & g[4715];
assign g[8812] = a[12] & g[4716];
assign g[12907] = b[12] & g[4716];
assign g[8813] = a[12] & g[4717];
assign g[12908] = b[12] & g[4717];
assign g[8814] = a[12] & g[4718];
assign g[12909] = b[12] & g[4718];
assign g[8815] = a[12] & g[4719];
assign g[12910] = b[12] & g[4719];
assign g[8816] = a[12] & g[4720];
assign g[12911] = b[12] & g[4720];
assign g[8817] = a[12] & g[4721];
assign g[12912] = b[12] & g[4721];
assign g[8818] = a[12] & g[4722];
assign g[12913] = b[12] & g[4722];
assign g[8819] = a[12] & g[4723];
assign g[12914] = b[12] & g[4723];
assign g[8820] = a[12] & g[4724];
assign g[12915] = b[12] & g[4724];
assign g[8821] = a[12] & g[4725];
assign g[12916] = b[12] & g[4725];
assign g[8822] = a[12] & g[4726];
assign g[12917] = b[12] & g[4726];
assign g[8823] = a[12] & g[4727];
assign g[12918] = b[12] & g[4727];
assign g[8824] = a[12] & g[4728];
assign g[12919] = b[12] & g[4728];
assign g[8825] = a[12] & g[4729];
assign g[12920] = b[12] & g[4729];
assign g[8826] = a[12] & g[4730];
assign g[12921] = b[12] & g[4730];
assign g[8827] = a[12] & g[4731];
assign g[12922] = b[12] & g[4731];
assign g[8828] = a[12] & g[4732];
assign g[12923] = b[12] & g[4732];
assign g[8829] = a[12] & g[4733];
assign g[12924] = b[12] & g[4733];
assign g[8830] = a[12] & g[4734];
assign g[12925] = b[12] & g[4734];
assign g[8831] = a[12] & g[4735];
assign g[12926] = b[12] & g[4735];
assign g[8832] = a[12] & g[4736];
assign g[12927] = b[12] & g[4736];
assign g[8833] = a[12] & g[4737];
assign g[12928] = b[12] & g[4737];
assign g[8834] = a[12] & g[4738];
assign g[12929] = b[12] & g[4738];
assign g[8835] = a[12] & g[4739];
assign g[12930] = b[12] & g[4739];
assign g[8836] = a[12] & g[4740];
assign g[12931] = b[12] & g[4740];
assign g[8837] = a[12] & g[4741];
assign g[12932] = b[12] & g[4741];
assign g[8838] = a[12] & g[4742];
assign g[12933] = b[12] & g[4742];
assign g[8839] = a[12] & g[4743];
assign g[12934] = b[12] & g[4743];
assign g[8840] = a[12] & g[4744];
assign g[12935] = b[12] & g[4744];
assign g[8841] = a[12] & g[4745];
assign g[12936] = b[12] & g[4745];
assign g[8842] = a[12] & g[4746];
assign g[12937] = b[12] & g[4746];
assign g[8843] = a[12] & g[4747];
assign g[12938] = b[12] & g[4747];
assign g[8844] = a[12] & g[4748];
assign g[12939] = b[12] & g[4748];
assign g[8845] = a[12] & g[4749];
assign g[12940] = b[12] & g[4749];
assign g[8846] = a[12] & g[4750];
assign g[12941] = b[12] & g[4750];
assign g[8847] = a[12] & g[4751];
assign g[12942] = b[12] & g[4751];
assign g[8848] = a[12] & g[4752];
assign g[12943] = b[12] & g[4752];
assign g[8849] = a[12] & g[4753];
assign g[12944] = b[12] & g[4753];
assign g[8850] = a[12] & g[4754];
assign g[12945] = b[12] & g[4754];
assign g[8851] = a[12] & g[4755];
assign g[12946] = b[12] & g[4755];
assign g[8852] = a[12] & g[4756];
assign g[12947] = b[12] & g[4756];
assign g[8853] = a[12] & g[4757];
assign g[12948] = b[12] & g[4757];
assign g[8854] = a[12] & g[4758];
assign g[12949] = b[12] & g[4758];
assign g[8855] = a[12] & g[4759];
assign g[12950] = b[12] & g[4759];
assign g[8856] = a[12] & g[4760];
assign g[12951] = b[12] & g[4760];
assign g[8857] = a[12] & g[4761];
assign g[12952] = b[12] & g[4761];
assign g[8858] = a[12] & g[4762];
assign g[12953] = b[12] & g[4762];
assign g[8859] = a[12] & g[4763];
assign g[12954] = b[12] & g[4763];
assign g[8860] = a[12] & g[4764];
assign g[12955] = b[12] & g[4764];
assign g[8861] = a[12] & g[4765];
assign g[12956] = b[12] & g[4765];
assign g[8862] = a[12] & g[4766];
assign g[12957] = b[12] & g[4766];
assign g[8863] = a[12] & g[4767];
assign g[12958] = b[12] & g[4767];
assign g[8864] = a[12] & g[4768];
assign g[12959] = b[12] & g[4768];
assign g[8865] = a[12] & g[4769];
assign g[12960] = b[12] & g[4769];
assign g[8866] = a[12] & g[4770];
assign g[12961] = b[12] & g[4770];
assign g[8867] = a[12] & g[4771];
assign g[12962] = b[12] & g[4771];
assign g[8868] = a[12] & g[4772];
assign g[12963] = b[12] & g[4772];
assign g[8869] = a[12] & g[4773];
assign g[12964] = b[12] & g[4773];
assign g[8870] = a[12] & g[4774];
assign g[12965] = b[12] & g[4774];
assign g[8871] = a[12] & g[4775];
assign g[12966] = b[12] & g[4775];
assign g[8872] = a[12] & g[4776];
assign g[12967] = b[12] & g[4776];
assign g[8873] = a[12] & g[4777];
assign g[12968] = b[12] & g[4777];
assign g[8874] = a[12] & g[4778];
assign g[12969] = b[12] & g[4778];
assign g[8875] = a[12] & g[4779];
assign g[12970] = b[12] & g[4779];
assign g[8876] = a[12] & g[4780];
assign g[12971] = b[12] & g[4780];
assign g[8877] = a[12] & g[4781];
assign g[12972] = b[12] & g[4781];
assign g[8878] = a[12] & g[4782];
assign g[12973] = b[12] & g[4782];
assign g[8879] = a[12] & g[4783];
assign g[12974] = b[12] & g[4783];
assign g[8880] = a[12] & g[4784];
assign g[12975] = b[12] & g[4784];
assign g[8881] = a[12] & g[4785];
assign g[12976] = b[12] & g[4785];
assign g[8882] = a[12] & g[4786];
assign g[12977] = b[12] & g[4786];
assign g[8883] = a[12] & g[4787];
assign g[12978] = b[12] & g[4787];
assign g[8884] = a[12] & g[4788];
assign g[12979] = b[12] & g[4788];
assign g[8885] = a[12] & g[4789];
assign g[12980] = b[12] & g[4789];
assign g[8886] = a[12] & g[4790];
assign g[12981] = b[12] & g[4790];
assign g[8887] = a[12] & g[4791];
assign g[12982] = b[12] & g[4791];
assign g[8888] = a[12] & g[4792];
assign g[12983] = b[12] & g[4792];
assign g[8889] = a[12] & g[4793];
assign g[12984] = b[12] & g[4793];
assign g[8890] = a[12] & g[4794];
assign g[12985] = b[12] & g[4794];
assign g[8891] = a[12] & g[4795];
assign g[12986] = b[12] & g[4795];
assign g[8892] = a[12] & g[4796];
assign g[12987] = b[12] & g[4796];
assign g[8893] = a[12] & g[4797];
assign g[12988] = b[12] & g[4797];
assign g[8894] = a[12] & g[4798];
assign g[12989] = b[12] & g[4798];
assign g[8895] = a[12] & g[4799];
assign g[12990] = b[12] & g[4799];
assign g[8896] = a[12] & g[4800];
assign g[12991] = b[12] & g[4800];
assign g[8897] = a[12] & g[4801];
assign g[12992] = b[12] & g[4801];
assign g[8898] = a[12] & g[4802];
assign g[12993] = b[12] & g[4802];
assign g[8899] = a[12] & g[4803];
assign g[12994] = b[12] & g[4803];
assign g[8900] = a[12] & g[4804];
assign g[12995] = b[12] & g[4804];
assign g[8901] = a[12] & g[4805];
assign g[12996] = b[12] & g[4805];
assign g[8902] = a[12] & g[4806];
assign g[12997] = b[12] & g[4806];
assign g[8903] = a[12] & g[4807];
assign g[12998] = b[12] & g[4807];
assign g[8904] = a[12] & g[4808];
assign g[12999] = b[12] & g[4808];
assign g[8905] = a[12] & g[4809];
assign g[13000] = b[12] & g[4809];
assign g[8906] = a[12] & g[4810];
assign g[13001] = b[12] & g[4810];
assign g[8907] = a[12] & g[4811];
assign g[13002] = b[12] & g[4811];
assign g[8908] = a[12] & g[4812];
assign g[13003] = b[12] & g[4812];
assign g[8909] = a[12] & g[4813];
assign g[13004] = b[12] & g[4813];
assign g[8910] = a[12] & g[4814];
assign g[13005] = b[12] & g[4814];
assign g[8911] = a[12] & g[4815];
assign g[13006] = b[12] & g[4815];
assign g[8912] = a[12] & g[4816];
assign g[13007] = b[12] & g[4816];
assign g[8913] = a[12] & g[4817];
assign g[13008] = b[12] & g[4817];
assign g[8914] = a[12] & g[4818];
assign g[13009] = b[12] & g[4818];
assign g[8915] = a[12] & g[4819];
assign g[13010] = b[12] & g[4819];
assign g[8916] = a[12] & g[4820];
assign g[13011] = b[12] & g[4820];
assign g[8917] = a[12] & g[4821];
assign g[13012] = b[12] & g[4821];
assign g[8918] = a[12] & g[4822];
assign g[13013] = b[12] & g[4822];
assign g[8919] = a[12] & g[4823];
assign g[13014] = b[12] & g[4823];
assign g[8920] = a[12] & g[4824];
assign g[13015] = b[12] & g[4824];
assign g[8921] = a[12] & g[4825];
assign g[13016] = b[12] & g[4825];
assign g[8922] = a[12] & g[4826];
assign g[13017] = b[12] & g[4826];
assign g[8923] = a[12] & g[4827];
assign g[13018] = b[12] & g[4827];
assign g[8924] = a[12] & g[4828];
assign g[13019] = b[12] & g[4828];
assign g[8925] = a[12] & g[4829];
assign g[13020] = b[12] & g[4829];
assign g[8926] = a[12] & g[4830];
assign g[13021] = b[12] & g[4830];
assign g[8927] = a[12] & g[4831];
assign g[13022] = b[12] & g[4831];
assign g[8928] = a[12] & g[4832];
assign g[13023] = b[12] & g[4832];
assign g[8929] = a[12] & g[4833];
assign g[13024] = b[12] & g[4833];
assign g[8930] = a[12] & g[4834];
assign g[13025] = b[12] & g[4834];
assign g[8931] = a[12] & g[4835];
assign g[13026] = b[12] & g[4835];
assign g[8932] = a[12] & g[4836];
assign g[13027] = b[12] & g[4836];
assign g[8933] = a[12] & g[4837];
assign g[13028] = b[12] & g[4837];
assign g[8934] = a[12] & g[4838];
assign g[13029] = b[12] & g[4838];
assign g[8935] = a[12] & g[4839];
assign g[13030] = b[12] & g[4839];
assign g[8936] = a[12] & g[4840];
assign g[13031] = b[12] & g[4840];
assign g[8937] = a[12] & g[4841];
assign g[13032] = b[12] & g[4841];
assign g[8938] = a[12] & g[4842];
assign g[13033] = b[12] & g[4842];
assign g[8939] = a[12] & g[4843];
assign g[13034] = b[12] & g[4843];
assign g[8940] = a[12] & g[4844];
assign g[13035] = b[12] & g[4844];
assign g[8941] = a[12] & g[4845];
assign g[13036] = b[12] & g[4845];
assign g[8942] = a[12] & g[4846];
assign g[13037] = b[12] & g[4846];
assign g[8943] = a[12] & g[4847];
assign g[13038] = b[12] & g[4847];
assign g[8944] = a[12] & g[4848];
assign g[13039] = b[12] & g[4848];
assign g[8945] = a[12] & g[4849];
assign g[13040] = b[12] & g[4849];
assign g[8946] = a[12] & g[4850];
assign g[13041] = b[12] & g[4850];
assign g[8947] = a[12] & g[4851];
assign g[13042] = b[12] & g[4851];
assign g[8948] = a[12] & g[4852];
assign g[13043] = b[12] & g[4852];
assign g[8949] = a[12] & g[4853];
assign g[13044] = b[12] & g[4853];
assign g[8950] = a[12] & g[4854];
assign g[13045] = b[12] & g[4854];
assign g[8951] = a[12] & g[4855];
assign g[13046] = b[12] & g[4855];
assign g[8952] = a[12] & g[4856];
assign g[13047] = b[12] & g[4856];
assign g[8953] = a[12] & g[4857];
assign g[13048] = b[12] & g[4857];
assign g[8954] = a[12] & g[4858];
assign g[13049] = b[12] & g[4858];
assign g[8955] = a[12] & g[4859];
assign g[13050] = b[12] & g[4859];
assign g[8956] = a[12] & g[4860];
assign g[13051] = b[12] & g[4860];
assign g[8957] = a[12] & g[4861];
assign g[13052] = b[12] & g[4861];
assign g[8958] = a[12] & g[4862];
assign g[13053] = b[12] & g[4862];
assign g[8959] = a[12] & g[4863];
assign g[13054] = b[12] & g[4863];
assign g[8960] = a[12] & g[4864];
assign g[13055] = b[12] & g[4864];
assign g[8961] = a[12] & g[4865];
assign g[13056] = b[12] & g[4865];
assign g[8962] = a[12] & g[4866];
assign g[13057] = b[12] & g[4866];
assign g[8963] = a[12] & g[4867];
assign g[13058] = b[12] & g[4867];
assign g[8964] = a[12] & g[4868];
assign g[13059] = b[12] & g[4868];
assign g[8965] = a[12] & g[4869];
assign g[13060] = b[12] & g[4869];
assign g[8966] = a[12] & g[4870];
assign g[13061] = b[12] & g[4870];
assign g[8967] = a[12] & g[4871];
assign g[13062] = b[12] & g[4871];
assign g[8968] = a[12] & g[4872];
assign g[13063] = b[12] & g[4872];
assign g[8969] = a[12] & g[4873];
assign g[13064] = b[12] & g[4873];
assign g[8970] = a[12] & g[4874];
assign g[13065] = b[12] & g[4874];
assign g[8971] = a[12] & g[4875];
assign g[13066] = b[12] & g[4875];
assign g[8972] = a[12] & g[4876];
assign g[13067] = b[12] & g[4876];
assign g[8973] = a[12] & g[4877];
assign g[13068] = b[12] & g[4877];
assign g[8974] = a[12] & g[4878];
assign g[13069] = b[12] & g[4878];
assign g[8975] = a[12] & g[4879];
assign g[13070] = b[12] & g[4879];
assign g[8976] = a[12] & g[4880];
assign g[13071] = b[12] & g[4880];
assign g[8977] = a[12] & g[4881];
assign g[13072] = b[12] & g[4881];
assign g[8978] = a[12] & g[4882];
assign g[13073] = b[12] & g[4882];
assign g[8979] = a[12] & g[4883];
assign g[13074] = b[12] & g[4883];
assign g[8980] = a[12] & g[4884];
assign g[13075] = b[12] & g[4884];
assign g[8981] = a[12] & g[4885];
assign g[13076] = b[12] & g[4885];
assign g[8982] = a[12] & g[4886];
assign g[13077] = b[12] & g[4886];
assign g[8983] = a[12] & g[4887];
assign g[13078] = b[12] & g[4887];
assign g[8984] = a[12] & g[4888];
assign g[13079] = b[12] & g[4888];
assign g[8985] = a[12] & g[4889];
assign g[13080] = b[12] & g[4889];
assign g[8986] = a[12] & g[4890];
assign g[13081] = b[12] & g[4890];
assign g[8987] = a[12] & g[4891];
assign g[13082] = b[12] & g[4891];
assign g[8988] = a[12] & g[4892];
assign g[13083] = b[12] & g[4892];
assign g[8989] = a[12] & g[4893];
assign g[13084] = b[12] & g[4893];
assign g[8990] = a[12] & g[4894];
assign g[13085] = b[12] & g[4894];
assign g[8991] = a[12] & g[4895];
assign g[13086] = b[12] & g[4895];
assign g[8992] = a[12] & g[4896];
assign g[13087] = b[12] & g[4896];
assign g[8993] = a[12] & g[4897];
assign g[13088] = b[12] & g[4897];
assign g[8994] = a[12] & g[4898];
assign g[13089] = b[12] & g[4898];
assign g[8995] = a[12] & g[4899];
assign g[13090] = b[12] & g[4899];
assign g[8996] = a[12] & g[4900];
assign g[13091] = b[12] & g[4900];
assign g[8997] = a[12] & g[4901];
assign g[13092] = b[12] & g[4901];
assign g[8998] = a[12] & g[4902];
assign g[13093] = b[12] & g[4902];
assign g[8999] = a[12] & g[4903];
assign g[13094] = b[12] & g[4903];
assign g[9000] = a[12] & g[4904];
assign g[13095] = b[12] & g[4904];
assign g[9001] = a[12] & g[4905];
assign g[13096] = b[12] & g[4905];
assign g[9002] = a[12] & g[4906];
assign g[13097] = b[12] & g[4906];
assign g[9003] = a[12] & g[4907];
assign g[13098] = b[12] & g[4907];
assign g[9004] = a[12] & g[4908];
assign g[13099] = b[12] & g[4908];
assign g[9005] = a[12] & g[4909];
assign g[13100] = b[12] & g[4909];
assign g[9006] = a[12] & g[4910];
assign g[13101] = b[12] & g[4910];
assign g[9007] = a[12] & g[4911];
assign g[13102] = b[12] & g[4911];
assign g[9008] = a[12] & g[4912];
assign g[13103] = b[12] & g[4912];
assign g[9009] = a[12] & g[4913];
assign g[13104] = b[12] & g[4913];
assign g[9010] = a[12] & g[4914];
assign g[13105] = b[12] & g[4914];
assign g[9011] = a[12] & g[4915];
assign g[13106] = b[12] & g[4915];
assign g[9012] = a[12] & g[4916];
assign g[13107] = b[12] & g[4916];
assign g[9013] = a[12] & g[4917];
assign g[13108] = b[12] & g[4917];
assign g[9014] = a[12] & g[4918];
assign g[13109] = b[12] & g[4918];
assign g[9015] = a[12] & g[4919];
assign g[13110] = b[12] & g[4919];
assign g[9016] = a[12] & g[4920];
assign g[13111] = b[12] & g[4920];
assign g[9017] = a[12] & g[4921];
assign g[13112] = b[12] & g[4921];
assign g[9018] = a[12] & g[4922];
assign g[13113] = b[12] & g[4922];
assign g[9019] = a[12] & g[4923];
assign g[13114] = b[12] & g[4923];
assign g[9020] = a[12] & g[4924];
assign g[13115] = b[12] & g[4924];
assign g[9021] = a[12] & g[4925];
assign g[13116] = b[12] & g[4925];
assign g[9022] = a[12] & g[4926];
assign g[13117] = b[12] & g[4926];
assign g[9023] = a[12] & g[4927];
assign g[13118] = b[12] & g[4927];
assign g[9024] = a[12] & g[4928];
assign g[13119] = b[12] & g[4928];
assign g[9025] = a[12] & g[4929];
assign g[13120] = b[12] & g[4929];
assign g[9026] = a[12] & g[4930];
assign g[13121] = b[12] & g[4930];
assign g[9027] = a[12] & g[4931];
assign g[13122] = b[12] & g[4931];
assign g[9028] = a[12] & g[4932];
assign g[13123] = b[12] & g[4932];
assign g[9029] = a[12] & g[4933];
assign g[13124] = b[12] & g[4933];
assign g[9030] = a[12] & g[4934];
assign g[13125] = b[12] & g[4934];
assign g[9031] = a[12] & g[4935];
assign g[13126] = b[12] & g[4935];
assign g[9032] = a[12] & g[4936];
assign g[13127] = b[12] & g[4936];
assign g[9033] = a[12] & g[4937];
assign g[13128] = b[12] & g[4937];
assign g[9034] = a[12] & g[4938];
assign g[13129] = b[12] & g[4938];
assign g[9035] = a[12] & g[4939];
assign g[13130] = b[12] & g[4939];
assign g[9036] = a[12] & g[4940];
assign g[13131] = b[12] & g[4940];
assign g[9037] = a[12] & g[4941];
assign g[13132] = b[12] & g[4941];
assign g[9038] = a[12] & g[4942];
assign g[13133] = b[12] & g[4942];
assign g[9039] = a[12] & g[4943];
assign g[13134] = b[12] & g[4943];
assign g[9040] = a[12] & g[4944];
assign g[13135] = b[12] & g[4944];
assign g[9041] = a[12] & g[4945];
assign g[13136] = b[12] & g[4945];
assign g[9042] = a[12] & g[4946];
assign g[13137] = b[12] & g[4946];
assign g[9043] = a[12] & g[4947];
assign g[13138] = b[12] & g[4947];
assign g[9044] = a[12] & g[4948];
assign g[13139] = b[12] & g[4948];
assign g[9045] = a[12] & g[4949];
assign g[13140] = b[12] & g[4949];
assign g[9046] = a[12] & g[4950];
assign g[13141] = b[12] & g[4950];
assign g[9047] = a[12] & g[4951];
assign g[13142] = b[12] & g[4951];
assign g[9048] = a[12] & g[4952];
assign g[13143] = b[12] & g[4952];
assign g[9049] = a[12] & g[4953];
assign g[13144] = b[12] & g[4953];
assign g[9050] = a[12] & g[4954];
assign g[13145] = b[12] & g[4954];
assign g[9051] = a[12] & g[4955];
assign g[13146] = b[12] & g[4955];
assign g[9052] = a[12] & g[4956];
assign g[13147] = b[12] & g[4956];
assign g[9053] = a[12] & g[4957];
assign g[13148] = b[12] & g[4957];
assign g[9054] = a[12] & g[4958];
assign g[13149] = b[12] & g[4958];
assign g[9055] = a[12] & g[4959];
assign g[13150] = b[12] & g[4959];
assign g[9056] = a[12] & g[4960];
assign g[13151] = b[12] & g[4960];
assign g[9057] = a[12] & g[4961];
assign g[13152] = b[12] & g[4961];
assign g[9058] = a[12] & g[4962];
assign g[13153] = b[12] & g[4962];
assign g[9059] = a[12] & g[4963];
assign g[13154] = b[12] & g[4963];
assign g[9060] = a[12] & g[4964];
assign g[13155] = b[12] & g[4964];
assign g[9061] = a[12] & g[4965];
assign g[13156] = b[12] & g[4965];
assign g[9062] = a[12] & g[4966];
assign g[13157] = b[12] & g[4966];
assign g[9063] = a[12] & g[4967];
assign g[13158] = b[12] & g[4967];
assign g[9064] = a[12] & g[4968];
assign g[13159] = b[12] & g[4968];
assign g[9065] = a[12] & g[4969];
assign g[13160] = b[12] & g[4969];
assign g[9066] = a[12] & g[4970];
assign g[13161] = b[12] & g[4970];
assign g[9067] = a[12] & g[4971];
assign g[13162] = b[12] & g[4971];
assign g[9068] = a[12] & g[4972];
assign g[13163] = b[12] & g[4972];
assign g[9069] = a[12] & g[4973];
assign g[13164] = b[12] & g[4973];
assign g[9070] = a[12] & g[4974];
assign g[13165] = b[12] & g[4974];
assign g[9071] = a[12] & g[4975];
assign g[13166] = b[12] & g[4975];
assign g[9072] = a[12] & g[4976];
assign g[13167] = b[12] & g[4976];
assign g[9073] = a[12] & g[4977];
assign g[13168] = b[12] & g[4977];
assign g[9074] = a[12] & g[4978];
assign g[13169] = b[12] & g[4978];
assign g[9075] = a[12] & g[4979];
assign g[13170] = b[12] & g[4979];
assign g[9076] = a[12] & g[4980];
assign g[13171] = b[12] & g[4980];
assign g[9077] = a[12] & g[4981];
assign g[13172] = b[12] & g[4981];
assign g[9078] = a[12] & g[4982];
assign g[13173] = b[12] & g[4982];
assign g[9079] = a[12] & g[4983];
assign g[13174] = b[12] & g[4983];
assign g[9080] = a[12] & g[4984];
assign g[13175] = b[12] & g[4984];
assign g[9081] = a[12] & g[4985];
assign g[13176] = b[12] & g[4985];
assign g[9082] = a[12] & g[4986];
assign g[13177] = b[12] & g[4986];
assign g[9083] = a[12] & g[4987];
assign g[13178] = b[12] & g[4987];
assign g[9084] = a[12] & g[4988];
assign g[13179] = b[12] & g[4988];
assign g[9085] = a[12] & g[4989];
assign g[13180] = b[12] & g[4989];
assign g[9086] = a[12] & g[4990];
assign g[13181] = b[12] & g[4990];
assign g[9087] = a[12] & g[4991];
assign g[13182] = b[12] & g[4991];
assign g[9088] = a[12] & g[4992];
assign g[13183] = b[12] & g[4992];
assign g[9089] = a[12] & g[4993];
assign g[13184] = b[12] & g[4993];
assign g[9090] = a[12] & g[4994];
assign g[13185] = b[12] & g[4994];
assign g[9091] = a[12] & g[4995];
assign g[13186] = b[12] & g[4995];
assign g[9092] = a[12] & g[4996];
assign g[13187] = b[12] & g[4996];
assign g[9093] = a[12] & g[4997];
assign g[13188] = b[12] & g[4997];
assign g[9094] = a[12] & g[4998];
assign g[13189] = b[12] & g[4998];
assign g[9095] = a[12] & g[4999];
assign g[13190] = b[12] & g[4999];
assign g[9096] = a[12] & g[5000];
assign g[13191] = b[12] & g[5000];
assign g[9097] = a[12] & g[5001];
assign g[13192] = b[12] & g[5001];
assign g[9098] = a[12] & g[5002];
assign g[13193] = b[12] & g[5002];
assign g[9099] = a[12] & g[5003];
assign g[13194] = b[12] & g[5003];
assign g[9100] = a[12] & g[5004];
assign g[13195] = b[12] & g[5004];
assign g[9101] = a[12] & g[5005];
assign g[13196] = b[12] & g[5005];
assign g[9102] = a[12] & g[5006];
assign g[13197] = b[12] & g[5006];
assign g[9103] = a[12] & g[5007];
assign g[13198] = b[12] & g[5007];
assign g[9104] = a[12] & g[5008];
assign g[13199] = b[12] & g[5008];
assign g[9105] = a[12] & g[5009];
assign g[13200] = b[12] & g[5009];
assign g[9106] = a[12] & g[5010];
assign g[13201] = b[12] & g[5010];
assign g[9107] = a[12] & g[5011];
assign g[13202] = b[12] & g[5011];
assign g[9108] = a[12] & g[5012];
assign g[13203] = b[12] & g[5012];
assign g[9109] = a[12] & g[5013];
assign g[13204] = b[12] & g[5013];
assign g[9110] = a[12] & g[5014];
assign g[13205] = b[12] & g[5014];
assign g[9111] = a[12] & g[5015];
assign g[13206] = b[12] & g[5015];
assign g[9112] = a[12] & g[5016];
assign g[13207] = b[12] & g[5016];
assign g[9113] = a[12] & g[5017];
assign g[13208] = b[12] & g[5017];
assign g[9114] = a[12] & g[5018];
assign g[13209] = b[12] & g[5018];
assign g[9115] = a[12] & g[5019];
assign g[13210] = b[12] & g[5019];
assign g[9116] = a[12] & g[5020];
assign g[13211] = b[12] & g[5020];
assign g[9117] = a[12] & g[5021];
assign g[13212] = b[12] & g[5021];
assign g[9118] = a[12] & g[5022];
assign g[13213] = b[12] & g[5022];
assign g[9119] = a[12] & g[5023];
assign g[13214] = b[12] & g[5023];
assign g[9120] = a[12] & g[5024];
assign g[13215] = b[12] & g[5024];
assign g[9121] = a[12] & g[5025];
assign g[13216] = b[12] & g[5025];
assign g[9122] = a[12] & g[5026];
assign g[13217] = b[12] & g[5026];
assign g[9123] = a[12] & g[5027];
assign g[13218] = b[12] & g[5027];
assign g[9124] = a[12] & g[5028];
assign g[13219] = b[12] & g[5028];
assign g[9125] = a[12] & g[5029];
assign g[13220] = b[12] & g[5029];
assign g[9126] = a[12] & g[5030];
assign g[13221] = b[12] & g[5030];
assign g[9127] = a[12] & g[5031];
assign g[13222] = b[12] & g[5031];
assign g[9128] = a[12] & g[5032];
assign g[13223] = b[12] & g[5032];
assign g[9129] = a[12] & g[5033];
assign g[13224] = b[12] & g[5033];
assign g[9130] = a[12] & g[5034];
assign g[13225] = b[12] & g[5034];
assign g[9131] = a[12] & g[5035];
assign g[13226] = b[12] & g[5035];
assign g[9132] = a[12] & g[5036];
assign g[13227] = b[12] & g[5036];
assign g[9133] = a[12] & g[5037];
assign g[13228] = b[12] & g[5037];
assign g[9134] = a[12] & g[5038];
assign g[13229] = b[12] & g[5038];
assign g[9135] = a[12] & g[5039];
assign g[13230] = b[12] & g[5039];
assign g[9136] = a[12] & g[5040];
assign g[13231] = b[12] & g[5040];
assign g[9137] = a[12] & g[5041];
assign g[13232] = b[12] & g[5041];
assign g[9138] = a[12] & g[5042];
assign g[13233] = b[12] & g[5042];
assign g[9139] = a[12] & g[5043];
assign g[13234] = b[12] & g[5043];
assign g[9140] = a[12] & g[5044];
assign g[13235] = b[12] & g[5044];
assign g[9141] = a[12] & g[5045];
assign g[13236] = b[12] & g[5045];
assign g[9142] = a[12] & g[5046];
assign g[13237] = b[12] & g[5046];
assign g[9143] = a[12] & g[5047];
assign g[13238] = b[12] & g[5047];
assign g[9144] = a[12] & g[5048];
assign g[13239] = b[12] & g[5048];
assign g[9145] = a[12] & g[5049];
assign g[13240] = b[12] & g[5049];
assign g[9146] = a[12] & g[5050];
assign g[13241] = b[12] & g[5050];
assign g[9147] = a[12] & g[5051];
assign g[13242] = b[12] & g[5051];
assign g[9148] = a[12] & g[5052];
assign g[13243] = b[12] & g[5052];
assign g[9149] = a[12] & g[5053];
assign g[13244] = b[12] & g[5053];
assign g[9150] = a[12] & g[5054];
assign g[13245] = b[12] & g[5054];
assign g[9151] = a[12] & g[5055];
assign g[13246] = b[12] & g[5055];
assign g[9152] = a[12] & g[5056];
assign g[13247] = b[12] & g[5056];
assign g[9153] = a[12] & g[5057];
assign g[13248] = b[12] & g[5057];
assign g[9154] = a[12] & g[5058];
assign g[13249] = b[12] & g[5058];
assign g[9155] = a[12] & g[5059];
assign g[13250] = b[12] & g[5059];
assign g[9156] = a[12] & g[5060];
assign g[13251] = b[12] & g[5060];
assign g[9157] = a[12] & g[5061];
assign g[13252] = b[12] & g[5061];
assign g[9158] = a[12] & g[5062];
assign g[13253] = b[12] & g[5062];
assign g[9159] = a[12] & g[5063];
assign g[13254] = b[12] & g[5063];
assign g[9160] = a[12] & g[5064];
assign g[13255] = b[12] & g[5064];
assign g[9161] = a[12] & g[5065];
assign g[13256] = b[12] & g[5065];
assign g[9162] = a[12] & g[5066];
assign g[13257] = b[12] & g[5066];
assign g[9163] = a[12] & g[5067];
assign g[13258] = b[12] & g[5067];
assign g[9164] = a[12] & g[5068];
assign g[13259] = b[12] & g[5068];
assign g[9165] = a[12] & g[5069];
assign g[13260] = b[12] & g[5069];
assign g[9166] = a[12] & g[5070];
assign g[13261] = b[12] & g[5070];
assign g[9167] = a[12] & g[5071];
assign g[13262] = b[12] & g[5071];
assign g[9168] = a[12] & g[5072];
assign g[13263] = b[12] & g[5072];
assign g[9169] = a[12] & g[5073];
assign g[13264] = b[12] & g[5073];
assign g[9170] = a[12] & g[5074];
assign g[13265] = b[12] & g[5074];
assign g[9171] = a[12] & g[5075];
assign g[13266] = b[12] & g[5075];
assign g[9172] = a[12] & g[5076];
assign g[13267] = b[12] & g[5076];
assign g[9173] = a[12] & g[5077];
assign g[13268] = b[12] & g[5077];
assign g[9174] = a[12] & g[5078];
assign g[13269] = b[12] & g[5078];
assign g[9175] = a[12] & g[5079];
assign g[13270] = b[12] & g[5079];
assign g[9176] = a[12] & g[5080];
assign g[13271] = b[12] & g[5080];
assign g[9177] = a[12] & g[5081];
assign g[13272] = b[12] & g[5081];
assign g[9178] = a[12] & g[5082];
assign g[13273] = b[12] & g[5082];
assign g[9179] = a[12] & g[5083];
assign g[13274] = b[12] & g[5083];
assign g[9180] = a[12] & g[5084];
assign g[13275] = b[12] & g[5084];
assign g[9181] = a[12] & g[5085];
assign g[13276] = b[12] & g[5085];
assign g[9182] = a[12] & g[5086];
assign g[13277] = b[12] & g[5086];
assign g[9183] = a[12] & g[5087];
assign g[13278] = b[12] & g[5087];
assign g[9184] = a[12] & g[5088];
assign g[13279] = b[12] & g[5088];
assign g[9185] = a[12] & g[5089];
assign g[13280] = b[12] & g[5089];
assign g[9186] = a[12] & g[5090];
assign g[13281] = b[12] & g[5090];
assign g[9187] = a[12] & g[5091];
assign g[13282] = b[12] & g[5091];
assign g[9188] = a[12] & g[5092];
assign g[13283] = b[12] & g[5092];
assign g[9189] = a[12] & g[5093];
assign g[13284] = b[12] & g[5093];
assign g[9190] = a[12] & g[5094];
assign g[13285] = b[12] & g[5094];
assign g[9191] = a[12] & g[5095];
assign g[13286] = b[12] & g[5095];
assign g[9192] = a[12] & g[5096];
assign g[13287] = b[12] & g[5096];
assign g[9193] = a[12] & g[5097];
assign g[13288] = b[12] & g[5097];
assign g[9194] = a[12] & g[5098];
assign g[13289] = b[12] & g[5098];
assign g[9195] = a[12] & g[5099];
assign g[13290] = b[12] & g[5099];
assign g[9196] = a[12] & g[5100];
assign g[13291] = b[12] & g[5100];
assign g[9197] = a[12] & g[5101];
assign g[13292] = b[12] & g[5101];
assign g[9198] = a[12] & g[5102];
assign g[13293] = b[12] & g[5102];
assign g[9199] = a[12] & g[5103];
assign g[13294] = b[12] & g[5103];
assign g[9200] = a[12] & g[5104];
assign g[13295] = b[12] & g[5104];
assign g[9201] = a[12] & g[5105];
assign g[13296] = b[12] & g[5105];
assign g[9202] = a[12] & g[5106];
assign g[13297] = b[12] & g[5106];
assign g[9203] = a[12] & g[5107];
assign g[13298] = b[12] & g[5107];
assign g[9204] = a[12] & g[5108];
assign g[13299] = b[12] & g[5108];
assign g[9205] = a[12] & g[5109];
assign g[13300] = b[12] & g[5109];
assign g[9206] = a[12] & g[5110];
assign g[13301] = b[12] & g[5110];
assign g[9207] = a[12] & g[5111];
assign g[13302] = b[12] & g[5111];
assign g[9208] = a[12] & g[5112];
assign g[13303] = b[12] & g[5112];
assign g[9209] = a[12] & g[5113];
assign g[13304] = b[12] & g[5113];
assign g[9210] = a[12] & g[5114];
assign g[13305] = b[12] & g[5114];
assign g[9211] = a[12] & g[5115];
assign g[13306] = b[12] & g[5115];
assign g[9212] = a[12] & g[5116];
assign g[13307] = b[12] & g[5116];
assign g[9213] = a[12] & g[5117];
assign g[13308] = b[12] & g[5117];
assign g[9214] = a[12] & g[5118];
assign g[13309] = b[12] & g[5118];
assign g[9215] = a[12] & g[5119];
assign g[13310] = b[12] & g[5119];
assign g[9216] = a[12] & g[5120];
assign g[13311] = b[12] & g[5120];
assign g[9217] = a[12] & g[5121];
assign g[13312] = b[12] & g[5121];
assign g[9218] = a[12] & g[5122];
assign g[13313] = b[12] & g[5122];
assign g[9219] = a[12] & g[5123];
assign g[13314] = b[12] & g[5123];
assign g[9220] = a[12] & g[5124];
assign g[13315] = b[12] & g[5124];
assign g[9221] = a[12] & g[5125];
assign g[13316] = b[12] & g[5125];
assign g[9222] = a[12] & g[5126];
assign g[13317] = b[12] & g[5126];
assign g[9223] = a[12] & g[5127];
assign g[13318] = b[12] & g[5127];
assign g[9224] = a[12] & g[5128];
assign g[13319] = b[12] & g[5128];
assign g[9225] = a[12] & g[5129];
assign g[13320] = b[12] & g[5129];
assign g[9226] = a[12] & g[5130];
assign g[13321] = b[12] & g[5130];
assign g[9227] = a[12] & g[5131];
assign g[13322] = b[12] & g[5131];
assign g[9228] = a[12] & g[5132];
assign g[13323] = b[12] & g[5132];
assign g[9229] = a[12] & g[5133];
assign g[13324] = b[12] & g[5133];
assign g[9230] = a[12] & g[5134];
assign g[13325] = b[12] & g[5134];
assign g[9231] = a[12] & g[5135];
assign g[13326] = b[12] & g[5135];
assign g[9232] = a[12] & g[5136];
assign g[13327] = b[12] & g[5136];
assign g[9233] = a[12] & g[5137];
assign g[13328] = b[12] & g[5137];
assign g[9234] = a[12] & g[5138];
assign g[13329] = b[12] & g[5138];
assign g[9235] = a[12] & g[5139];
assign g[13330] = b[12] & g[5139];
assign g[9236] = a[12] & g[5140];
assign g[13331] = b[12] & g[5140];
assign g[9237] = a[12] & g[5141];
assign g[13332] = b[12] & g[5141];
assign g[9238] = a[12] & g[5142];
assign g[13333] = b[12] & g[5142];
assign g[9239] = a[12] & g[5143];
assign g[13334] = b[12] & g[5143];
assign g[9240] = a[12] & g[5144];
assign g[13335] = b[12] & g[5144];
assign g[9241] = a[12] & g[5145];
assign g[13336] = b[12] & g[5145];
assign g[9242] = a[12] & g[5146];
assign g[13337] = b[12] & g[5146];
assign g[9243] = a[12] & g[5147];
assign g[13338] = b[12] & g[5147];
assign g[9244] = a[12] & g[5148];
assign g[13339] = b[12] & g[5148];
assign g[9245] = a[12] & g[5149];
assign g[13340] = b[12] & g[5149];
assign g[9246] = a[12] & g[5150];
assign g[13341] = b[12] & g[5150];
assign g[9247] = a[12] & g[5151];
assign g[13342] = b[12] & g[5151];
assign g[9248] = a[12] & g[5152];
assign g[13343] = b[12] & g[5152];
assign g[9249] = a[12] & g[5153];
assign g[13344] = b[12] & g[5153];
assign g[9250] = a[12] & g[5154];
assign g[13345] = b[12] & g[5154];
assign g[9251] = a[12] & g[5155];
assign g[13346] = b[12] & g[5155];
assign g[9252] = a[12] & g[5156];
assign g[13347] = b[12] & g[5156];
assign g[9253] = a[12] & g[5157];
assign g[13348] = b[12] & g[5157];
assign g[9254] = a[12] & g[5158];
assign g[13349] = b[12] & g[5158];
assign g[9255] = a[12] & g[5159];
assign g[13350] = b[12] & g[5159];
assign g[9256] = a[12] & g[5160];
assign g[13351] = b[12] & g[5160];
assign g[9257] = a[12] & g[5161];
assign g[13352] = b[12] & g[5161];
assign g[9258] = a[12] & g[5162];
assign g[13353] = b[12] & g[5162];
assign g[9259] = a[12] & g[5163];
assign g[13354] = b[12] & g[5163];
assign g[9260] = a[12] & g[5164];
assign g[13355] = b[12] & g[5164];
assign g[9261] = a[12] & g[5165];
assign g[13356] = b[12] & g[5165];
assign g[9262] = a[12] & g[5166];
assign g[13357] = b[12] & g[5166];
assign g[9263] = a[12] & g[5167];
assign g[13358] = b[12] & g[5167];
assign g[9264] = a[12] & g[5168];
assign g[13359] = b[12] & g[5168];
assign g[9265] = a[12] & g[5169];
assign g[13360] = b[12] & g[5169];
assign g[9266] = a[12] & g[5170];
assign g[13361] = b[12] & g[5170];
assign g[9267] = a[12] & g[5171];
assign g[13362] = b[12] & g[5171];
assign g[9268] = a[12] & g[5172];
assign g[13363] = b[12] & g[5172];
assign g[9269] = a[12] & g[5173];
assign g[13364] = b[12] & g[5173];
assign g[9270] = a[12] & g[5174];
assign g[13365] = b[12] & g[5174];
assign g[9271] = a[12] & g[5175];
assign g[13366] = b[12] & g[5175];
assign g[9272] = a[12] & g[5176];
assign g[13367] = b[12] & g[5176];
assign g[9273] = a[12] & g[5177];
assign g[13368] = b[12] & g[5177];
assign g[9274] = a[12] & g[5178];
assign g[13369] = b[12] & g[5178];
assign g[9275] = a[12] & g[5179];
assign g[13370] = b[12] & g[5179];
assign g[9276] = a[12] & g[5180];
assign g[13371] = b[12] & g[5180];
assign g[9277] = a[12] & g[5181];
assign g[13372] = b[12] & g[5181];
assign g[9278] = a[12] & g[5182];
assign g[13373] = b[12] & g[5182];
assign g[9279] = a[12] & g[5183];
assign g[13374] = b[12] & g[5183];
assign g[9280] = a[12] & g[5184];
assign g[13375] = b[12] & g[5184];
assign g[9281] = a[12] & g[5185];
assign g[13376] = b[12] & g[5185];
assign g[9282] = a[12] & g[5186];
assign g[13377] = b[12] & g[5186];
assign g[9283] = a[12] & g[5187];
assign g[13378] = b[12] & g[5187];
assign g[9284] = a[12] & g[5188];
assign g[13379] = b[12] & g[5188];
assign g[9285] = a[12] & g[5189];
assign g[13380] = b[12] & g[5189];
assign g[9286] = a[12] & g[5190];
assign g[13381] = b[12] & g[5190];
assign g[9287] = a[12] & g[5191];
assign g[13382] = b[12] & g[5191];
assign g[9288] = a[12] & g[5192];
assign g[13383] = b[12] & g[5192];
assign g[9289] = a[12] & g[5193];
assign g[13384] = b[12] & g[5193];
assign g[9290] = a[12] & g[5194];
assign g[13385] = b[12] & g[5194];
assign g[9291] = a[12] & g[5195];
assign g[13386] = b[12] & g[5195];
assign g[9292] = a[12] & g[5196];
assign g[13387] = b[12] & g[5196];
assign g[9293] = a[12] & g[5197];
assign g[13388] = b[12] & g[5197];
assign g[9294] = a[12] & g[5198];
assign g[13389] = b[12] & g[5198];
assign g[9295] = a[12] & g[5199];
assign g[13390] = b[12] & g[5199];
assign g[9296] = a[12] & g[5200];
assign g[13391] = b[12] & g[5200];
assign g[9297] = a[12] & g[5201];
assign g[13392] = b[12] & g[5201];
assign g[9298] = a[12] & g[5202];
assign g[13393] = b[12] & g[5202];
assign g[9299] = a[12] & g[5203];
assign g[13394] = b[12] & g[5203];
assign g[9300] = a[12] & g[5204];
assign g[13395] = b[12] & g[5204];
assign g[9301] = a[12] & g[5205];
assign g[13396] = b[12] & g[5205];
assign g[9302] = a[12] & g[5206];
assign g[13397] = b[12] & g[5206];
assign g[9303] = a[12] & g[5207];
assign g[13398] = b[12] & g[5207];
assign g[9304] = a[12] & g[5208];
assign g[13399] = b[12] & g[5208];
assign g[9305] = a[12] & g[5209];
assign g[13400] = b[12] & g[5209];
assign g[9306] = a[12] & g[5210];
assign g[13401] = b[12] & g[5210];
assign g[9307] = a[12] & g[5211];
assign g[13402] = b[12] & g[5211];
assign g[9308] = a[12] & g[5212];
assign g[13403] = b[12] & g[5212];
assign g[9309] = a[12] & g[5213];
assign g[13404] = b[12] & g[5213];
assign g[9310] = a[12] & g[5214];
assign g[13405] = b[12] & g[5214];
assign g[9311] = a[12] & g[5215];
assign g[13406] = b[12] & g[5215];
assign g[9312] = a[12] & g[5216];
assign g[13407] = b[12] & g[5216];
assign g[9313] = a[12] & g[5217];
assign g[13408] = b[12] & g[5217];
assign g[9314] = a[12] & g[5218];
assign g[13409] = b[12] & g[5218];
assign g[9315] = a[12] & g[5219];
assign g[13410] = b[12] & g[5219];
assign g[9316] = a[12] & g[5220];
assign g[13411] = b[12] & g[5220];
assign g[9317] = a[12] & g[5221];
assign g[13412] = b[12] & g[5221];
assign g[9318] = a[12] & g[5222];
assign g[13413] = b[12] & g[5222];
assign g[9319] = a[12] & g[5223];
assign g[13414] = b[12] & g[5223];
assign g[9320] = a[12] & g[5224];
assign g[13415] = b[12] & g[5224];
assign g[9321] = a[12] & g[5225];
assign g[13416] = b[12] & g[5225];
assign g[9322] = a[12] & g[5226];
assign g[13417] = b[12] & g[5226];
assign g[9323] = a[12] & g[5227];
assign g[13418] = b[12] & g[5227];
assign g[9324] = a[12] & g[5228];
assign g[13419] = b[12] & g[5228];
assign g[9325] = a[12] & g[5229];
assign g[13420] = b[12] & g[5229];
assign g[9326] = a[12] & g[5230];
assign g[13421] = b[12] & g[5230];
assign g[9327] = a[12] & g[5231];
assign g[13422] = b[12] & g[5231];
assign g[9328] = a[12] & g[5232];
assign g[13423] = b[12] & g[5232];
assign g[9329] = a[12] & g[5233];
assign g[13424] = b[12] & g[5233];
assign g[9330] = a[12] & g[5234];
assign g[13425] = b[12] & g[5234];
assign g[9331] = a[12] & g[5235];
assign g[13426] = b[12] & g[5235];
assign g[9332] = a[12] & g[5236];
assign g[13427] = b[12] & g[5236];
assign g[9333] = a[12] & g[5237];
assign g[13428] = b[12] & g[5237];
assign g[9334] = a[12] & g[5238];
assign g[13429] = b[12] & g[5238];
assign g[9335] = a[12] & g[5239];
assign g[13430] = b[12] & g[5239];
assign g[9336] = a[12] & g[5240];
assign g[13431] = b[12] & g[5240];
assign g[9337] = a[12] & g[5241];
assign g[13432] = b[12] & g[5241];
assign g[9338] = a[12] & g[5242];
assign g[13433] = b[12] & g[5242];
assign g[9339] = a[12] & g[5243];
assign g[13434] = b[12] & g[5243];
assign g[9340] = a[12] & g[5244];
assign g[13435] = b[12] & g[5244];
assign g[9341] = a[12] & g[5245];
assign g[13436] = b[12] & g[5245];
assign g[9342] = a[12] & g[5246];
assign g[13437] = b[12] & g[5246];
assign g[9343] = a[12] & g[5247];
assign g[13438] = b[12] & g[5247];
assign g[9344] = a[12] & g[5248];
assign g[13439] = b[12] & g[5248];
assign g[9345] = a[12] & g[5249];
assign g[13440] = b[12] & g[5249];
assign g[9346] = a[12] & g[5250];
assign g[13441] = b[12] & g[5250];
assign g[9347] = a[12] & g[5251];
assign g[13442] = b[12] & g[5251];
assign g[9348] = a[12] & g[5252];
assign g[13443] = b[12] & g[5252];
assign g[9349] = a[12] & g[5253];
assign g[13444] = b[12] & g[5253];
assign g[9350] = a[12] & g[5254];
assign g[13445] = b[12] & g[5254];
assign g[9351] = a[12] & g[5255];
assign g[13446] = b[12] & g[5255];
assign g[9352] = a[12] & g[5256];
assign g[13447] = b[12] & g[5256];
assign g[9353] = a[12] & g[5257];
assign g[13448] = b[12] & g[5257];
assign g[9354] = a[12] & g[5258];
assign g[13449] = b[12] & g[5258];
assign g[9355] = a[12] & g[5259];
assign g[13450] = b[12] & g[5259];
assign g[9356] = a[12] & g[5260];
assign g[13451] = b[12] & g[5260];
assign g[9357] = a[12] & g[5261];
assign g[13452] = b[12] & g[5261];
assign g[9358] = a[12] & g[5262];
assign g[13453] = b[12] & g[5262];
assign g[9359] = a[12] & g[5263];
assign g[13454] = b[12] & g[5263];
assign g[9360] = a[12] & g[5264];
assign g[13455] = b[12] & g[5264];
assign g[9361] = a[12] & g[5265];
assign g[13456] = b[12] & g[5265];
assign g[9362] = a[12] & g[5266];
assign g[13457] = b[12] & g[5266];
assign g[9363] = a[12] & g[5267];
assign g[13458] = b[12] & g[5267];
assign g[9364] = a[12] & g[5268];
assign g[13459] = b[12] & g[5268];
assign g[9365] = a[12] & g[5269];
assign g[13460] = b[12] & g[5269];
assign g[9366] = a[12] & g[5270];
assign g[13461] = b[12] & g[5270];
assign g[9367] = a[12] & g[5271];
assign g[13462] = b[12] & g[5271];
assign g[9368] = a[12] & g[5272];
assign g[13463] = b[12] & g[5272];
assign g[9369] = a[12] & g[5273];
assign g[13464] = b[12] & g[5273];
assign g[9370] = a[12] & g[5274];
assign g[13465] = b[12] & g[5274];
assign g[9371] = a[12] & g[5275];
assign g[13466] = b[12] & g[5275];
assign g[9372] = a[12] & g[5276];
assign g[13467] = b[12] & g[5276];
assign g[9373] = a[12] & g[5277];
assign g[13468] = b[12] & g[5277];
assign g[9374] = a[12] & g[5278];
assign g[13469] = b[12] & g[5278];
assign g[9375] = a[12] & g[5279];
assign g[13470] = b[12] & g[5279];
assign g[9376] = a[12] & g[5280];
assign g[13471] = b[12] & g[5280];
assign g[9377] = a[12] & g[5281];
assign g[13472] = b[12] & g[5281];
assign g[9378] = a[12] & g[5282];
assign g[13473] = b[12] & g[5282];
assign g[9379] = a[12] & g[5283];
assign g[13474] = b[12] & g[5283];
assign g[9380] = a[12] & g[5284];
assign g[13475] = b[12] & g[5284];
assign g[9381] = a[12] & g[5285];
assign g[13476] = b[12] & g[5285];
assign g[9382] = a[12] & g[5286];
assign g[13477] = b[12] & g[5286];
assign g[9383] = a[12] & g[5287];
assign g[13478] = b[12] & g[5287];
assign g[9384] = a[12] & g[5288];
assign g[13479] = b[12] & g[5288];
assign g[9385] = a[12] & g[5289];
assign g[13480] = b[12] & g[5289];
assign g[9386] = a[12] & g[5290];
assign g[13481] = b[12] & g[5290];
assign g[9387] = a[12] & g[5291];
assign g[13482] = b[12] & g[5291];
assign g[9388] = a[12] & g[5292];
assign g[13483] = b[12] & g[5292];
assign g[9389] = a[12] & g[5293];
assign g[13484] = b[12] & g[5293];
assign g[9390] = a[12] & g[5294];
assign g[13485] = b[12] & g[5294];
assign g[9391] = a[12] & g[5295];
assign g[13486] = b[12] & g[5295];
assign g[9392] = a[12] & g[5296];
assign g[13487] = b[12] & g[5296];
assign g[9393] = a[12] & g[5297];
assign g[13488] = b[12] & g[5297];
assign g[9394] = a[12] & g[5298];
assign g[13489] = b[12] & g[5298];
assign g[9395] = a[12] & g[5299];
assign g[13490] = b[12] & g[5299];
assign g[9396] = a[12] & g[5300];
assign g[13491] = b[12] & g[5300];
assign g[9397] = a[12] & g[5301];
assign g[13492] = b[12] & g[5301];
assign g[9398] = a[12] & g[5302];
assign g[13493] = b[12] & g[5302];
assign g[9399] = a[12] & g[5303];
assign g[13494] = b[12] & g[5303];
assign g[9400] = a[12] & g[5304];
assign g[13495] = b[12] & g[5304];
assign g[9401] = a[12] & g[5305];
assign g[13496] = b[12] & g[5305];
assign g[9402] = a[12] & g[5306];
assign g[13497] = b[12] & g[5306];
assign g[9403] = a[12] & g[5307];
assign g[13498] = b[12] & g[5307];
assign g[9404] = a[12] & g[5308];
assign g[13499] = b[12] & g[5308];
assign g[9405] = a[12] & g[5309];
assign g[13500] = b[12] & g[5309];
assign g[9406] = a[12] & g[5310];
assign g[13501] = b[12] & g[5310];
assign g[9407] = a[12] & g[5311];
assign g[13502] = b[12] & g[5311];
assign g[9408] = a[12] & g[5312];
assign g[13503] = b[12] & g[5312];
assign g[9409] = a[12] & g[5313];
assign g[13504] = b[12] & g[5313];
assign g[9410] = a[12] & g[5314];
assign g[13505] = b[12] & g[5314];
assign g[9411] = a[12] & g[5315];
assign g[13506] = b[12] & g[5315];
assign g[9412] = a[12] & g[5316];
assign g[13507] = b[12] & g[5316];
assign g[9413] = a[12] & g[5317];
assign g[13508] = b[12] & g[5317];
assign g[9414] = a[12] & g[5318];
assign g[13509] = b[12] & g[5318];
assign g[9415] = a[12] & g[5319];
assign g[13510] = b[12] & g[5319];
assign g[9416] = a[12] & g[5320];
assign g[13511] = b[12] & g[5320];
assign g[9417] = a[12] & g[5321];
assign g[13512] = b[12] & g[5321];
assign g[9418] = a[12] & g[5322];
assign g[13513] = b[12] & g[5322];
assign g[9419] = a[12] & g[5323];
assign g[13514] = b[12] & g[5323];
assign g[9420] = a[12] & g[5324];
assign g[13515] = b[12] & g[5324];
assign g[9421] = a[12] & g[5325];
assign g[13516] = b[12] & g[5325];
assign g[9422] = a[12] & g[5326];
assign g[13517] = b[12] & g[5326];
assign g[9423] = a[12] & g[5327];
assign g[13518] = b[12] & g[5327];
assign g[9424] = a[12] & g[5328];
assign g[13519] = b[12] & g[5328];
assign g[9425] = a[12] & g[5329];
assign g[13520] = b[12] & g[5329];
assign g[9426] = a[12] & g[5330];
assign g[13521] = b[12] & g[5330];
assign g[9427] = a[12] & g[5331];
assign g[13522] = b[12] & g[5331];
assign g[9428] = a[12] & g[5332];
assign g[13523] = b[12] & g[5332];
assign g[9429] = a[12] & g[5333];
assign g[13524] = b[12] & g[5333];
assign g[9430] = a[12] & g[5334];
assign g[13525] = b[12] & g[5334];
assign g[9431] = a[12] & g[5335];
assign g[13526] = b[12] & g[5335];
assign g[9432] = a[12] & g[5336];
assign g[13527] = b[12] & g[5336];
assign g[9433] = a[12] & g[5337];
assign g[13528] = b[12] & g[5337];
assign g[9434] = a[12] & g[5338];
assign g[13529] = b[12] & g[5338];
assign g[9435] = a[12] & g[5339];
assign g[13530] = b[12] & g[5339];
assign g[9436] = a[12] & g[5340];
assign g[13531] = b[12] & g[5340];
assign g[9437] = a[12] & g[5341];
assign g[13532] = b[12] & g[5341];
assign g[9438] = a[12] & g[5342];
assign g[13533] = b[12] & g[5342];
assign g[9439] = a[12] & g[5343];
assign g[13534] = b[12] & g[5343];
assign g[9440] = a[12] & g[5344];
assign g[13535] = b[12] & g[5344];
assign g[9441] = a[12] & g[5345];
assign g[13536] = b[12] & g[5345];
assign g[9442] = a[12] & g[5346];
assign g[13537] = b[12] & g[5346];
assign g[9443] = a[12] & g[5347];
assign g[13538] = b[12] & g[5347];
assign g[9444] = a[12] & g[5348];
assign g[13539] = b[12] & g[5348];
assign g[9445] = a[12] & g[5349];
assign g[13540] = b[12] & g[5349];
assign g[9446] = a[12] & g[5350];
assign g[13541] = b[12] & g[5350];
assign g[9447] = a[12] & g[5351];
assign g[13542] = b[12] & g[5351];
assign g[9448] = a[12] & g[5352];
assign g[13543] = b[12] & g[5352];
assign g[9449] = a[12] & g[5353];
assign g[13544] = b[12] & g[5353];
assign g[9450] = a[12] & g[5354];
assign g[13545] = b[12] & g[5354];
assign g[9451] = a[12] & g[5355];
assign g[13546] = b[12] & g[5355];
assign g[9452] = a[12] & g[5356];
assign g[13547] = b[12] & g[5356];
assign g[9453] = a[12] & g[5357];
assign g[13548] = b[12] & g[5357];
assign g[9454] = a[12] & g[5358];
assign g[13549] = b[12] & g[5358];
assign g[9455] = a[12] & g[5359];
assign g[13550] = b[12] & g[5359];
assign g[9456] = a[12] & g[5360];
assign g[13551] = b[12] & g[5360];
assign g[9457] = a[12] & g[5361];
assign g[13552] = b[12] & g[5361];
assign g[9458] = a[12] & g[5362];
assign g[13553] = b[12] & g[5362];
assign g[9459] = a[12] & g[5363];
assign g[13554] = b[12] & g[5363];
assign g[9460] = a[12] & g[5364];
assign g[13555] = b[12] & g[5364];
assign g[9461] = a[12] & g[5365];
assign g[13556] = b[12] & g[5365];
assign g[9462] = a[12] & g[5366];
assign g[13557] = b[12] & g[5366];
assign g[9463] = a[12] & g[5367];
assign g[13558] = b[12] & g[5367];
assign g[9464] = a[12] & g[5368];
assign g[13559] = b[12] & g[5368];
assign g[9465] = a[12] & g[5369];
assign g[13560] = b[12] & g[5369];
assign g[9466] = a[12] & g[5370];
assign g[13561] = b[12] & g[5370];
assign g[9467] = a[12] & g[5371];
assign g[13562] = b[12] & g[5371];
assign g[9468] = a[12] & g[5372];
assign g[13563] = b[12] & g[5372];
assign g[9469] = a[12] & g[5373];
assign g[13564] = b[12] & g[5373];
assign g[9470] = a[12] & g[5374];
assign g[13565] = b[12] & g[5374];
assign g[9471] = a[12] & g[5375];
assign g[13566] = b[12] & g[5375];
assign g[9472] = a[12] & g[5376];
assign g[13567] = b[12] & g[5376];
assign g[9473] = a[12] & g[5377];
assign g[13568] = b[12] & g[5377];
assign g[9474] = a[12] & g[5378];
assign g[13569] = b[12] & g[5378];
assign g[9475] = a[12] & g[5379];
assign g[13570] = b[12] & g[5379];
assign g[9476] = a[12] & g[5380];
assign g[13571] = b[12] & g[5380];
assign g[9477] = a[12] & g[5381];
assign g[13572] = b[12] & g[5381];
assign g[9478] = a[12] & g[5382];
assign g[13573] = b[12] & g[5382];
assign g[9479] = a[12] & g[5383];
assign g[13574] = b[12] & g[5383];
assign g[9480] = a[12] & g[5384];
assign g[13575] = b[12] & g[5384];
assign g[9481] = a[12] & g[5385];
assign g[13576] = b[12] & g[5385];
assign g[9482] = a[12] & g[5386];
assign g[13577] = b[12] & g[5386];
assign g[9483] = a[12] & g[5387];
assign g[13578] = b[12] & g[5387];
assign g[9484] = a[12] & g[5388];
assign g[13579] = b[12] & g[5388];
assign g[9485] = a[12] & g[5389];
assign g[13580] = b[12] & g[5389];
assign g[9486] = a[12] & g[5390];
assign g[13581] = b[12] & g[5390];
assign g[9487] = a[12] & g[5391];
assign g[13582] = b[12] & g[5391];
assign g[9488] = a[12] & g[5392];
assign g[13583] = b[12] & g[5392];
assign g[9489] = a[12] & g[5393];
assign g[13584] = b[12] & g[5393];
assign g[9490] = a[12] & g[5394];
assign g[13585] = b[12] & g[5394];
assign g[9491] = a[12] & g[5395];
assign g[13586] = b[12] & g[5395];
assign g[9492] = a[12] & g[5396];
assign g[13587] = b[12] & g[5396];
assign g[9493] = a[12] & g[5397];
assign g[13588] = b[12] & g[5397];
assign g[9494] = a[12] & g[5398];
assign g[13589] = b[12] & g[5398];
assign g[9495] = a[12] & g[5399];
assign g[13590] = b[12] & g[5399];
assign g[9496] = a[12] & g[5400];
assign g[13591] = b[12] & g[5400];
assign g[9497] = a[12] & g[5401];
assign g[13592] = b[12] & g[5401];
assign g[9498] = a[12] & g[5402];
assign g[13593] = b[12] & g[5402];
assign g[9499] = a[12] & g[5403];
assign g[13594] = b[12] & g[5403];
assign g[9500] = a[12] & g[5404];
assign g[13595] = b[12] & g[5404];
assign g[9501] = a[12] & g[5405];
assign g[13596] = b[12] & g[5405];
assign g[9502] = a[12] & g[5406];
assign g[13597] = b[12] & g[5406];
assign g[9503] = a[12] & g[5407];
assign g[13598] = b[12] & g[5407];
assign g[9504] = a[12] & g[5408];
assign g[13599] = b[12] & g[5408];
assign g[9505] = a[12] & g[5409];
assign g[13600] = b[12] & g[5409];
assign g[9506] = a[12] & g[5410];
assign g[13601] = b[12] & g[5410];
assign g[9507] = a[12] & g[5411];
assign g[13602] = b[12] & g[5411];
assign g[9508] = a[12] & g[5412];
assign g[13603] = b[12] & g[5412];
assign g[9509] = a[12] & g[5413];
assign g[13604] = b[12] & g[5413];
assign g[9510] = a[12] & g[5414];
assign g[13605] = b[12] & g[5414];
assign g[9511] = a[12] & g[5415];
assign g[13606] = b[12] & g[5415];
assign g[9512] = a[12] & g[5416];
assign g[13607] = b[12] & g[5416];
assign g[9513] = a[12] & g[5417];
assign g[13608] = b[12] & g[5417];
assign g[9514] = a[12] & g[5418];
assign g[13609] = b[12] & g[5418];
assign g[9515] = a[12] & g[5419];
assign g[13610] = b[12] & g[5419];
assign g[9516] = a[12] & g[5420];
assign g[13611] = b[12] & g[5420];
assign g[9517] = a[12] & g[5421];
assign g[13612] = b[12] & g[5421];
assign g[9518] = a[12] & g[5422];
assign g[13613] = b[12] & g[5422];
assign g[9519] = a[12] & g[5423];
assign g[13614] = b[12] & g[5423];
assign g[9520] = a[12] & g[5424];
assign g[13615] = b[12] & g[5424];
assign g[9521] = a[12] & g[5425];
assign g[13616] = b[12] & g[5425];
assign g[9522] = a[12] & g[5426];
assign g[13617] = b[12] & g[5426];
assign g[9523] = a[12] & g[5427];
assign g[13618] = b[12] & g[5427];
assign g[9524] = a[12] & g[5428];
assign g[13619] = b[12] & g[5428];
assign g[9525] = a[12] & g[5429];
assign g[13620] = b[12] & g[5429];
assign g[9526] = a[12] & g[5430];
assign g[13621] = b[12] & g[5430];
assign g[9527] = a[12] & g[5431];
assign g[13622] = b[12] & g[5431];
assign g[9528] = a[12] & g[5432];
assign g[13623] = b[12] & g[5432];
assign g[9529] = a[12] & g[5433];
assign g[13624] = b[12] & g[5433];
assign g[9530] = a[12] & g[5434];
assign g[13625] = b[12] & g[5434];
assign g[9531] = a[12] & g[5435];
assign g[13626] = b[12] & g[5435];
assign g[9532] = a[12] & g[5436];
assign g[13627] = b[12] & g[5436];
assign g[9533] = a[12] & g[5437];
assign g[13628] = b[12] & g[5437];
assign g[9534] = a[12] & g[5438];
assign g[13629] = b[12] & g[5438];
assign g[9535] = a[12] & g[5439];
assign g[13630] = b[12] & g[5439];
assign g[9536] = a[12] & g[5440];
assign g[13631] = b[12] & g[5440];
assign g[9537] = a[12] & g[5441];
assign g[13632] = b[12] & g[5441];
assign g[9538] = a[12] & g[5442];
assign g[13633] = b[12] & g[5442];
assign g[9539] = a[12] & g[5443];
assign g[13634] = b[12] & g[5443];
assign g[9540] = a[12] & g[5444];
assign g[13635] = b[12] & g[5444];
assign g[9541] = a[12] & g[5445];
assign g[13636] = b[12] & g[5445];
assign g[9542] = a[12] & g[5446];
assign g[13637] = b[12] & g[5446];
assign g[9543] = a[12] & g[5447];
assign g[13638] = b[12] & g[5447];
assign g[9544] = a[12] & g[5448];
assign g[13639] = b[12] & g[5448];
assign g[9545] = a[12] & g[5449];
assign g[13640] = b[12] & g[5449];
assign g[9546] = a[12] & g[5450];
assign g[13641] = b[12] & g[5450];
assign g[9547] = a[12] & g[5451];
assign g[13642] = b[12] & g[5451];
assign g[9548] = a[12] & g[5452];
assign g[13643] = b[12] & g[5452];
assign g[9549] = a[12] & g[5453];
assign g[13644] = b[12] & g[5453];
assign g[9550] = a[12] & g[5454];
assign g[13645] = b[12] & g[5454];
assign g[9551] = a[12] & g[5455];
assign g[13646] = b[12] & g[5455];
assign g[9552] = a[12] & g[5456];
assign g[13647] = b[12] & g[5456];
assign g[9553] = a[12] & g[5457];
assign g[13648] = b[12] & g[5457];
assign g[9554] = a[12] & g[5458];
assign g[13649] = b[12] & g[5458];
assign g[9555] = a[12] & g[5459];
assign g[13650] = b[12] & g[5459];
assign g[9556] = a[12] & g[5460];
assign g[13651] = b[12] & g[5460];
assign g[9557] = a[12] & g[5461];
assign g[13652] = b[12] & g[5461];
assign g[9558] = a[12] & g[5462];
assign g[13653] = b[12] & g[5462];
assign g[9559] = a[12] & g[5463];
assign g[13654] = b[12] & g[5463];
assign g[9560] = a[12] & g[5464];
assign g[13655] = b[12] & g[5464];
assign g[9561] = a[12] & g[5465];
assign g[13656] = b[12] & g[5465];
assign g[9562] = a[12] & g[5466];
assign g[13657] = b[12] & g[5466];
assign g[9563] = a[12] & g[5467];
assign g[13658] = b[12] & g[5467];
assign g[9564] = a[12] & g[5468];
assign g[13659] = b[12] & g[5468];
assign g[9565] = a[12] & g[5469];
assign g[13660] = b[12] & g[5469];
assign g[9566] = a[12] & g[5470];
assign g[13661] = b[12] & g[5470];
assign g[9567] = a[12] & g[5471];
assign g[13662] = b[12] & g[5471];
assign g[9568] = a[12] & g[5472];
assign g[13663] = b[12] & g[5472];
assign g[9569] = a[12] & g[5473];
assign g[13664] = b[12] & g[5473];
assign g[9570] = a[12] & g[5474];
assign g[13665] = b[12] & g[5474];
assign g[9571] = a[12] & g[5475];
assign g[13666] = b[12] & g[5475];
assign g[9572] = a[12] & g[5476];
assign g[13667] = b[12] & g[5476];
assign g[9573] = a[12] & g[5477];
assign g[13668] = b[12] & g[5477];
assign g[9574] = a[12] & g[5478];
assign g[13669] = b[12] & g[5478];
assign g[9575] = a[12] & g[5479];
assign g[13670] = b[12] & g[5479];
assign g[9576] = a[12] & g[5480];
assign g[13671] = b[12] & g[5480];
assign g[9577] = a[12] & g[5481];
assign g[13672] = b[12] & g[5481];
assign g[9578] = a[12] & g[5482];
assign g[13673] = b[12] & g[5482];
assign g[9579] = a[12] & g[5483];
assign g[13674] = b[12] & g[5483];
assign g[9580] = a[12] & g[5484];
assign g[13675] = b[12] & g[5484];
assign g[9581] = a[12] & g[5485];
assign g[13676] = b[12] & g[5485];
assign g[9582] = a[12] & g[5486];
assign g[13677] = b[12] & g[5486];
assign g[9583] = a[12] & g[5487];
assign g[13678] = b[12] & g[5487];
assign g[9584] = a[12] & g[5488];
assign g[13679] = b[12] & g[5488];
assign g[9585] = a[12] & g[5489];
assign g[13680] = b[12] & g[5489];
assign g[9586] = a[12] & g[5490];
assign g[13681] = b[12] & g[5490];
assign g[9587] = a[12] & g[5491];
assign g[13682] = b[12] & g[5491];
assign g[9588] = a[12] & g[5492];
assign g[13683] = b[12] & g[5492];
assign g[9589] = a[12] & g[5493];
assign g[13684] = b[12] & g[5493];
assign g[9590] = a[12] & g[5494];
assign g[13685] = b[12] & g[5494];
assign g[9591] = a[12] & g[5495];
assign g[13686] = b[12] & g[5495];
assign g[9592] = a[12] & g[5496];
assign g[13687] = b[12] & g[5496];
assign g[9593] = a[12] & g[5497];
assign g[13688] = b[12] & g[5497];
assign g[9594] = a[12] & g[5498];
assign g[13689] = b[12] & g[5498];
assign g[9595] = a[12] & g[5499];
assign g[13690] = b[12] & g[5499];
assign g[9596] = a[12] & g[5500];
assign g[13691] = b[12] & g[5500];
assign g[9597] = a[12] & g[5501];
assign g[13692] = b[12] & g[5501];
assign g[9598] = a[12] & g[5502];
assign g[13693] = b[12] & g[5502];
assign g[9599] = a[12] & g[5503];
assign g[13694] = b[12] & g[5503];
assign g[9600] = a[12] & g[5504];
assign g[13695] = b[12] & g[5504];
assign g[9601] = a[12] & g[5505];
assign g[13696] = b[12] & g[5505];
assign g[9602] = a[12] & g[5506];
assign g[13697] = b[12] & g[5506];
assign g[9603] = a[12] & g[5507];
assign g[13698] = b[12] & g[5507];
assign g[9604] = a[12] & g[5508];
assign g[13699] = b[12] & g[5508];
assign g[9605] = a[12] & g[5509];
assign g[13700] = b[12] & g[5509];
assign g[9606] = a[12] & g[5510];
assign g[13701] = b[12] & g[5510];
assign g[9607] = a[12] & g[5511];
assign g[13702] = b[12] & g[5511];
assign g[9608] = a[12] & g[5512];
assign g[13703] = b[12] & g[5512];
assign g[9609] = a[12] & g[5513];
assign g[13704] = b[12] & g[5513];
assign g[9610] = a[12] & g[5514];
assign g[13705] = b[12] & g[5514];
assign g[9611] = a[12] & g[5515];
assign g[13706] = b[12] & g[5515];
assign g[9612] = a[12] & g[5516];
assign g[13707] = b[12] & g[5516];
assign g[9613] = a[12] & g[5517];
assign g[13708] = b[12] & g[5517];
assign g[9614] = a[12] & g[5518];
assign g[13709] = b[12] & g[5518];
assign g[9615] = a[12] & g[5519];
assign g[13710] = b[12] & g[5519];
assign g[9616] = a[12] & g[5520];
assign g[13711] = b[12] & g[5520];
assign g[9617] = a[12] & g[5521];
assign g[13712] = b[12] & g[5521];
assign g[9618] = a[12] & g[5522];
assign g[13713] = b[12] & g[5522];
assign g[9619] = a[12] & g[5523];
assign g[13714] = b[12] & g[5523];
assign g[9620] = a[12] & g[5524];
assign g[13715] = b[12] & g[5524];
assign g[9621] = a[12] & g[5525];
assign g[13716] = b[12] & g[5525];
assign g[9622] = a[12] & g[5526];
assign g[13717] = b[12] & g[5526];
assign g[9623] = a[12] & g[5527];
assign g[13718] = b[12] & g[5527];
assign g[9624] = a[12] & g[5528];
assign g[13719] = b[12] & g[5528];
assign g[9625] = a[12] & g[5529];
assign g[13720] = b[12] & g[5529];
assign g[9626] = a[12] & g[5530];
assign g[13721] = b[12] & g[5530];
assign g[9627] = a[12] & g[5531];
assign g[13722] = b[12] & g[5531];
assign g[9628] = a[12] & g[5532];
assign g[13723] = b[12] & g[5532];
assign g[9629] = a[12] & g[5533];
assign g[13724] = b[12] & g[5533];
assign g[9630] = a[12] & g[5534];
assign g[13725] = b[12] & g[5534];
assign g[9631] = a[12] & g[5535];
assign g[13726] = b[12] & g[5535];
assign g[9632] = a[12] & g[5536];
assign g[13727] = b[12] & g[5536];
assign g[9633] = a[12] & g[5537];
assign g[13728] = b[12] & g[5537];
assign g[9634] = a[12] & g[5538];
assign g[13729] = b[12] & g[5538];
assign g[9635] = a[12] & g[5539];
assign g[13730] = b[12] & g[5539];
assign g[9636] = a[12] & g[5540];
assign g[13731] = b[12] & g[5540];
assign g[9637] = a[12] & g[5541];
assign g[13732] = b[12] & g[5541];
assign g[9638] = a[12] & g[5542];
assign g[13733] = b[12] & g[5542];
assign g[9639] = a[12] & g[5543];
assign g[13734] = b[12] & g[5543];
assign g[9640] = a[12] & g[5544];
assign g[13735] = b[12] & g[5544];
assign g[9641] = a[12] & g[5545];
assign g[13736] = b[12] & g[5545];
assign g[9642] = a[12] & g[5546];
assign g[13737] = b[12] & g[5546];
assign g[9643] = a[12] & g[5547];
assign g[13738] = b[12] & g[5547];
assign g[9644] = a[12] & g[5548];
assign g[13739] = b[12] & g[5548];
assign g[9645] = a[12] & g[5549];
assign g[13740] = b[12] & g[5549];
assign g[9646] = a[12] & g[5550];
assign g[13741] = b[12] & g[5550];
assign g[9647] = a[12] & g[5551];
assign g[13742] = b[12] & g[5551];
assign g[9648] = a[12] & g[5552];
assign g[13743] = b[12] & g[5552];
assign g[9649] = a[12] & g[5553];
assign g[13744] = b[12] & g[5553];
assign g[9650] = a[12] & g[5554];
assign g[13745] = b[12] & g[5554];
assign g[9651] = a[12] & g[5555];
assign g[13746] = b[12] & g[5555];
assign g[9652] = a[12] & g[5556];
assign g[13747] = b[12] & g[5556];
assign g[9653] = a[12] & g[5557];
assign g[13748] = b[12] & g[5557];
assign g[9654] = a[12] & g[5558];
assign g[13749] = b[12] & g[5558];
assign g[9655] = a[12] & g[5559];
assign g[13750] = b[12] & g[5559];
assign g[9656] = a[12] & g[5560];
assign g[13751] = b[12] & g[5560];
assign g[9657] = a[12] & g[5561];
assign g[13752] = b[12] & g[5561];
assign g[9658] = a[12] & g[5562];
assign g[13753] = b[12] & g[5562];
assign g[9659] = a[12] & g[5563];
assign g[13754] = b[12] & g[5563];
assign g[9660] = a[12] & g[5564];
assign g[13755] = b[12] & g[5564];
assign g[9661] = a[12] & g[5565];
assign g[13756] = b[12] & g[5565];
assign g[9662] = a[12] & g[5566];
assign g[13757] = b[12] & g[5566];
assign g[9663] = a[12] & g[5567];
assign g[13758] = b[12] & g[5567];
assign g[9664] = a[12] & g[5568];
assign g[13759] = b[12] & g[5568];
assign g[9665] = a[12] & g[5569];
assign g[13760] = b[12] & g[5569];
assign g[9666] = a[12] & g[5570];
assign g[13761] = b[12] & g[5570];
assign g[9667] = a[12] & g[5571];
assign g[13762] = b[12] & g[5571];
assign g[9668] = a[12] & g[5572];
assign g[13763] = b[12] & g[5572];
assign g[9669] = a[12] & g[5573];
assign g[13764] = b[12] & g[5573];
assign g[9670] = a[12] & g[5574];
assign g[13765] = b[12] & g[5574];
assign g[9671] = a[12] & g[5575];
assign g[13766] = b[12] & g[5575];
assign g[9672] = a[12] & g[5576];
assign g[13767] = b[12] & g[5576];
assign g[9673] = a[12] & g[5577];
assign g[13768] = b[12] & g[5577];
assign g[9674] = a[12] & g[5578];
assign g[13769] = b[12] & g[5578];
assign g[9675] = a[12] & g[5579];
assign g[13770] = b[12] & g[5579];
assign g[9676] = a[12] & g[5580];
assign g[13771] = b[12] & g[5580];
assign g[9677] = a[12] & g[5581];
assign g[13772] = b[12] & g[5581];
assign g[9678] = a[12] & g[5582];
assign g[13773] = b[12] & g[5582];
assign g[9679] = a[12] & g[5583];
assign g[13774] = b[12] & g[5583];
assign g[9680] = a[12] & g[5584];
assign g[13775] = b[12] & g[5584];
assign g[9681] = a[12] & g[5585];
assign g[13776] = b[12] & g[5585];
assign g[9682] = a[12] & g[5586];
assign g[13777] = b[12] & g[5586];
assign g[9683] = a[12] & g[5587];
assign g[13778] = b[12] & g[5587];
assign g[9684] = a[12] & g[5588];
assign g[13779] = b[12] & g[5588];
assign g[9685] = a[12] & g[5589];
assign g[13780] = b[12] & g[5589];
assign g[9686] = a[12] & g[5590];
assign g[13781] = b[12] & g[5590];
assign g[9687] = a[12] & g[5591];
assign g[13782] = b[12] & g[5591];
assign g[9688] = a[12] & g[5592];
assign g[13783] = b[12] & g[5592];
assign g[9689] = a[12] & g[5593];
assign g[13784] = b[12] & g[5593];
assign g[9690] = a[12] & g[5594];
assign g[13785] = b[12] & g[5594];
assign g[9691] = a[12] & g[5595];
assign g[13786] = b[12] & g[5595];
assign g[9692] = a[12] & g[5596];
assign g[13787] = b[12] & g[5596];
assign g[9693] = a[12] & g[5597];
assign g[13788] = b[12] & g[5597];
assign g[9694] = a[12] & g[5598];
assign g[13789] = b[12] & g[5598];
assign g[9695] = a[12] & g[5599];
assign g[13790] = b[12] & g[5599];
assign g[9696] = a[12] & g[5600];
assign g[13791] = b[12] & g[5600];
assign g[9697] = a[12] & g[5601];
assign g[13792] = b[12] & g[5601];
assign g[9698] = a[12] & g[5602];
assign g[13793] = b[12] & g[5602];
assign g[9699] = a[12] & g[5603];
assign g[13794] = b[12] & g[5603];
assign g[9700] = a[12] & g[5604];
assign g[13795] = b[12] & g[5604];
assign g[9701] = a[12] & g[5605];
assign g[13796] = b[12] & g[5605];
assign g[9702] = a[12] & g[5606];
assign g[13797] = b[12] & g[5606];
assign g[9703] = a[12] & g[5607];
assign g[13798] = b[12] & g[5607];
assign g[9704] = a[12] & g[5608];
assign g[13799] = b[12] & g[5608];
assign g[9705] = a[12] & g[5609];
assign g[13800] = b[12] & g[5609];
assign g[9706] = a[12] & g[5610];
assign g[13801] = b[12] & g[5610];
assign g[9707] = a[12] & g[5611];
assign g[13802] = b[12] & g[5611];
assign g[9708] = a[12] & g[5612];
assign g[13803] = b[12] & g[5612];
assign g[9709] = a[12] & g[5613];
assign g[13804] = b[12] & g[5613];
assign g[9710] = a[12] & g[5614];
assign g[13805] = b[12] & g[5614];
assign g[9711] = a[12] & g[5615];
assign g[13806] = b[12] & g[5615];
assign g[9712] = a[12] & g[5616];
assign g[13807] = b[12] & g[5616];
assign g[9713] = a[12] & g[5617];
assign g[13808] = b[12] & g[5617];
assign g[9714] = a[12] & g[5618];
assign g[13809] = b[12] & g[5618];
assign g[9715] = a[12] & g[5619];
assign g[13810] = b[12] & g[5619];
assign g[9716] = a[12] & g[5620];
assign g[13811] = b[12] & g[5620];
assign g[9717] = a[12] & g[5621];
assign g[13812] = b[12] & g[5621];
assign g[9718] = a[12] & g[5622];
assign g[13813] = b[12] & g[5622];
assign g[9719] = a[12] & g[5623];
assign g[13814] = b[12] & g[5623];
assign g[9720] = a[12] & g[5624];
assign g[13815] = b[12] & g[5624];
assign g[9721] = a[12] & g[5625];
assign g[13816] = b[12] & g[5625];
assign g[9722] = a[12] & g[5626];
assign g[13817] = b[12] & g[5626];
assign g[9723] = a[12] & g[5627];
assign g[13818] = b[12] & g[5627];
assign g[9724] = a[12] & g[5628];
assign g[13819] = b[12] & g[5628];
assign g[9725] = a[12] & g[5629];
assign g[13820] = b[12] & g[5629];
assign g[9726] = a[12] & g[5630];
assign g[13821] = b[12] & g[5630];
assign g[9727] = a[12] & g[5631];
assign g[13822] = b[12] & g[5631];
assign g[9728] = a[12] & g[5632];
assign g[13823] = b[12] & g[5632];
assign g[9729] = a[12] & g[5633];
assign g[13824] = b[12] & g[5633];
assign g[9730] = a[12] & g[5634];
assign g[13825] = b[12] & g[5634];
assign g[9731] = a[12] & g[5635];
assign g[13826] = b[12] & g[5635];
assign g[9732] = a[12] & g[5636];
assign g[13827] = b[12] & g[5636];
assign g[9733] = a[12] & g[5637];
assign g[13828] = b[12] & g[5637];
assign g[9734] = a[12] & g[5638];
assign g[13829] = b[12] & g[5638];
assign g[9735] = a[12] & g[5639];
assign g[13830] = b[12] & g[5639];
assign g[9736] = a[12] & g[5640];
assign g[13831] = b[12] & g[5640];
assign g[9737] = a[12] & g[5641];
assign g[13832] = b[12] & g[5641];
assign g[9738] = a[12] & g[5642];
assign g[13833] = b[12] & g[5642];
assign g[9739] = a[12] & g[5643];
assign g[13834] = b[12] & g[5643];
assign g[9740] = a[12] & g[5644];
assign g[13835] = b[12] & g[5644];
assign g[9741] = a[12] & g[5645];
assign g[13836] = b[12] & g[5645];
assign g[9742] = a[12] & g[5646];
assign g[13837] = b[12] & g[5646];
assign g[9743] = a[12] & g[5647];
assign g[13838] = b[12] & g[5647];
assign g[9744] = a[12] & g[5648];
assign g[13839] = b[12] & g[5648];
assign g[9745] = a[12] & g[5649];
assign g[13840] = b[12] & g[5649];
assign g[9746] = a[12] & g[5650];
assign g[13841] = b[12] & g[5650];
assign g[9747] = a[12] & g[5651];
assign g[13842] = b[12] & g[5651];
assign g[9748] = a[12] & g[5652];
assign g[13843] = b[12] & g[5652];
assign g[9749] = a[12] & g[5653];
assign g[13844] = b[12] & g[5653];
assign g[9750] = a[12] & g[5654];
assign g[13845] = b[12] & g[5654];
assign g[9751] = a[12] & g[5655];
assign g[13846] = b[12] & g[5655];
assign g[9752] = a[12] & g[5656];
assign g[13847] = b[12] & g[5656];
assign g[9753] = a[12] & g[5657];
assign g[13848] = b[12] & g[5657];
assign g[9754] = a[12] & g[5658];
assign g[13849] = b[12] & g[5658];
assign g[9755] = a[12] & g[5659];
assign g[13850] = b[12] & g[5659];
assign g[9756] = a[12] & g[5660];
assign g[13851] = b[12] & g[5660];
assign g[9757] = a[12] & g[5661];
assign g[13852] = b[12] & g[5661];
assign g[9758] = a[12] & g[5662];
assign g[13853] = b[12] & g[5662];
assign g[9759] = a[12] & g[5663];
assign g[13854] = b[12] & g[5663];
assign g[9760] = a[12] & g[5664];
assign g[13855] = b[12] & g[5664];
assign g[9761] = a[12] & g[5665];
assign g[13856] = b[12] & g[5665];
assign g[9762] = a[12] & g[5666];
assign g[13857] = b[12] & g[5666];
assign g[9763] = a[12] & g[5667];
assign g[13858] = b[12] & g[5667];
assign g[9764] = a[12] & g[5668];
assign g[13859] = b[12] & g[5668];
assign g[9765] = a[12] & g[5669];
assign g[13860] = b[12] & g[5669];
assign g[9766] = a[12] & g[5670];
assign g[13861] = b[12] & g[5670];
assign g[9767] = a[12] & g[5671];
assign g[13862] = b[12] & g[5671];
assign g[9768] = a[12] & g[5672];
assign g[13863] = b[12] & g[5672];
assign g[9769] = a[12] & g[5673];
assign g[13864] = b[12] & g[5673];
assign g[9770] = a[12] & g[5674];
assign g[13865] = b[12] & g[5674];
assign g[9771] = a[12] & g[5675];
assign g[13866] = b[12] & g[5675];
assign g[9772] = a[12] & g[5676];
assign g[13867] = b[12] & g[5676];
assign g[9773] = a[12] & g[5677];
assign g[13868] = b[12] & g[5677];
assign g[9774] = a[12] & g[5678];
assign g[13869] = b[12] & g[5678];
assign g[9775] = a[12] & g[5679];
assign g[13870] = b[12] & g[5679];
assign g[9776] = a[12] & g[5680];
assign g[13871] = b[12] & g[5680];
assign g[9777] = a[12] & g[5681];
assign g[13872] = b[12] & g[5681];
assign g[9778] = a[12] & g[5682];
assign g[13873] = b[12] & g[5682];
assign g[9779] = a[12] & g[5683];
assign g[13874] = b[12] & g[5683];
assign g[9780] = a[12] & g[5684];
assign g[13875] = b[12] & g[5684];
assign g[9781] = a[12] & g[5685];
assign g[13876] = b[12] & g[5685];
assign g[9782] = a[12] & g[5686];
assign g[13877] = b[12] & g[5686];
assign g[9783] = a[12] & g[5687];
assign g[13878] = b[12] & g[5687];
assign g[9784] = a[12] & g[5688];
assign g[13879] = b[12] & g[5688];
assign g[9785] = a[12] & g[5689];
assign g[13880] = b[12] & g[5689];
assign g[9786] = a[12] & g[5690];
assign g[13881] = b[12] & g[5690];
assign g[9787] = a[12] & g[5691];
assign g[13882] = b[12] & g[5691];
assign g[9788] = a[12] & g[5692];
assign g[13883] = b[12] & g[5692];
assign g[9789] = a[12] & g[5693];
assign g[13884] = b[12] & g[5693];
assign g[9790] = a[12] & g[5694];
assign g[13885] = b[12] & g[5694];
assign g[9791] = a[12] & g[5695];
assign g[13886] = b[12] & g[5695];
assign g[9792] = a[12] & g[5696];
assign g[13887] = b[12] & g[5696];
assign g[9793] = a[12] & g[5697];
assign g[13888] = b[12] & g[5697];
assign g[9794] = a[12] & g[5698];
assign g[13889] = b[12] & g[5698];
assign g[9795] = a[12] & g[5699];
assign g[13890] = b[12] & g[5699];
assign g[9796] = a[12] & g[5700];
assign g[13891] = b[12] & g[5700];
assign g[9797] = a[12] & g[5701];
assign g[13892] = b[12] & g[5701];
assign g[9798] = a[12] & g[5702];
assign g[13893] = b[12] & g[5702];
assign g[9799] = a[12] & g[5703];
assign g[13894] = b[12] & g[5703];
assign g[9800] = a[12] & g[5704];
assign g[13895] = b[12] & g[5704];
assign g[9801] = a[12] & g[5705];
assign g[13896] = b[12] & g[5705];
assign g[9802] = a[12] & g[5706];
assign g[13897] = b[12] & g[5706];
assign g[9803] = a[12] & g[5707];
assign g[13898] = b[12] & g[5707];
assign g[9804] = a[12] & g[5708];
assign g[13899] = b[12] & g[5708];
assign g[9805] = a[12] & g[5709];
assign g[13900] = b[12] & g[5709];
assign g[9806] = a[12] & g[5710];
assign g[13901] = b[12] & g[5710];
assign g[9807] = a[12] & g[5711];
assign g[13902] = b[12] & g[5711];
assign g[9808] = a[12] & g[5712];
assign g[13903] = b[12] & g[5712];
assign g[9809] = a[12] & g[5713];
assign g[13904] = b[12] & g[5713];
assign g[9810] = a[12] & g[5714];
assign g[13905] = b[12] & g[5714];
assign g[9811] = a[12] & g[5715];
assign g[13906] = b[12] & g[5715];
assign g[9812] = a[12] & g[5716];
assign g[13907] = b[12] & g[5716];
assign g[9813] = a[12] & g[5717];
assign g[13908] = b[12] & g[5717];
assign g[9814] = a[12] & g[5718];
assign g[13909] = b[12] & g[5718];
assign g[9815] = a[12] & g[5719];
assign g[13910] = b[12] & g[5719];
assign g[9816] = a[12] & g[5720];
assign g[13911] = b[12] & g[5720];
assign g[9817] = a[12] & g[5721];
assign g[13912] = b[12] & g[5721];
assign g[9818] = a[12] & g[5722];
assign g[13913] = b[12] & g[5722];
assign g[9819] = a[12] & g[5723];
assign g[13914] = b[12] & g[5723];
assign g[9820] = a[12] & g[5724];
assign g[13915] = b[12] & g[5724];
assign g[9821] = a[12] & g[5725];
assign g[13916] = b[12] & g[5725];
assign g[9822] = a[12] & g[5726];
assign g[13917] = b[12] & g[5726];
assign g[9823] = a[12] & g[5727];
assign g[13918] = b[12] & g[5727];
assign g[9824] = a[12] & g[5728];
assign g[13919] = b[12] & g[5728];
assign g[9825] = a[12] & g[5729];
assign g[13920] = b[12] & g[5729];
assign g[9826] = a[12] & g[5730];
assign g[13921] = b[12] & g[5730];
assign g[9827] = a[12] & g[5731];
assign g[13922] = b[12] & g[5731];
assign g[9828] = a[12] & g[5732];
assign g[13923] = b[12] & g[5732];
assign g[9829] = a[12] & g[5733];
assign g[13924] = b[12] & g[5733];
assign g[9830] = a[12] & g[5734];
assign g[13925] = b[12] & g[5734];
assign g[9831] = a[12] & g[5735];
assign g[13926] = b[12] & g[5735];
assign g[9832] = a[12] & g[5736];
assign g[13927] = b[12] & g[5736];
assign g[9833] = a[12] & g[5737];
assign g[13928] = b[12] & g[5737];
assign g[9834] = a[12] & g[5738];
assign g[13929] = b[12] & g[5738];
assign g[9835] = a[12] & g[5739];
assign g[13930] = b[12] & g[5739];
assign g[9836] = a[12] & g[5740];
assign g[13931] = b[12] & g[5740];
assign g[9837] = a[12] & g[5741];
assign g[13932] = b[12] & g[5741];
assign g[9838] = a[12] & g[5742];
assign g[13933] = b[12] & g[5742];
assign g[9839] = a[12] & g[5743];
assign g[13934] = b[12] & g[5743];
assign g[9840] = a[12] & g[5744];
assign g[13935] = b[12] & g[5744];
assign g[9841] = a[12] & g[5745];
assign g[13936] = b[12] & g[5745];
assign g[9842] = a[12] & g[5746];
assign g[13937] = b[12] & g[5746];
assign g[9843] = a[12] & g[5747];
assign g[13938] = b[12] & g[5747];
assign g[9844] = a[12] & g[5748];
assign g[13939] = b[12] & g[5748];
assign g[9845] = a[12] & g[5749];
assign g[13940] = b[12] & g[5749];
assign g[9846] = a[12] & g[5750];
assign g[13941] = b[12] & g[5750];
assign g[9847] = a[12] & g[5751];
assign g[13942] = b[12] & g[5751];
assign g[9848] = a[12] & g[5752];
assign g[13943] = b[12] & g[5752];
assign g[9849] = a[12] & g[5753];
assign g[13944] = b[12] & g[5753];
assign g[9850] = a[12] & g[5754];
assign g[13945] = b[12] & g[5754];
assign g[9851] = a[12] & g[5755];
assign g[13946] = b[12] & g[5755];
assign g[9852] = a[12] & g[5756];
assign g[13947] = b[12] & g[5756];
assign g[9853] = a[12] & g[5757];
assign g[13948] = b[12] & g[5757];
assign g[9854] = a[12] & g[5758];
assign g[13949] = b[12] & g[5758];
assign g[9855] = a[12] & g[5759];
assign g[13950] = b[12] & g[5759];
assign g[9856] = a[12] & g[5760];
assign g[13951] = b[12] & g[5760];
assign g[9857] = a[12] & g[5761];
assign g[13952] = b[12] & g[5761];
assign g[9858] = a[12] & g[5762];
assign g[13953] = b[12] & g[5762];
assign g[9859] = a[12] & g[5763];
assign g[13954] = b[12] & g[5763];
assign g[9860] = a[12] & g[5764];
assign g[13955] = b[12] & g[5764];
assign g[9861] = a[12] & g[5765];
assign g[13956] = b[12] & g[5765];
assign g[9862] = a[12] & g[5766];
assign g[13957] = b[12] & g[5766];
assign g[9863] = a[12] & g[5767];
assign g[13958] = b[12] & g[5767];
assign g[9864] = a[12] & g[5768];
assign g[13959] = b[12] & g[5768];
assign g[9865] = a[12] & g[5769];
assign g[13960] = b[12] & g[5769];
assign g[9866] = a[12] & g[5770];
assign g[13961] = b[12] & g[5770];
assign g[9867] = a[12] & g[5771];
assign g[13962] = b[12] & g[5771];
assign g[9868] = a[12] & g[5772];
assign g[13963] = b[12] & g[5772];
assign g[9869] = a[12] & g[5773];
assign g[13964] = b[12] & g[5773];
assign g[9870] = a[12] & g[5774];
assign g[13965] = b[12] & g[5774];
assign g[9871] = a[12] & g[5775];
assign g[13966] = b[12] & g[5775];
assign g[9872] = a[12] & g[5776];
assign g[13967] = b[12] & g[5776];
assign g[9873] = a[12] & g[5777];
assign g[13968] = b[12] & g[5777];
assign g[9874] = a[12] & g[5778];
assign g[13969] = b[12] & g[5778];
assign g[9875] = a[12] & g[5779];
assign g[13970] = b[12] & g[5779];
assign g[9876] = a[12] & g[5780];
assign g[13971] = b[12] & g[5780];
assign g[9877] = a[12] & g[5781];
assign g[13972] = b[12] & g[5781];
assign g[9878] = a[12] & g[5782];
assign g[13973] = b[12] & g[5782];
assign g[9879] = a[12] & g[5783];
assign g[13974] = b[12] & g[5783];
assign g[9880] = a[12] & g[5784];
assign g[13975] = b[12] & g[5784];
assign g[9881] = a[12] & g[5785];
assign g[13976] = b[12] & g[5785];
assign g[9882] = a[12] & g[5786];
assign g[13977] = b[12] & g[5786];
assign g[9883] = a[12] & g[5787];
assign g[13978] = b[12] & g[5787];
assign g[9884] = a[12] & g[5788];
assign g[13979] = b[12] & g[5788];
assign g[9885] = a[12] & g[5789];
assign g[13980] = b[12] & g[5789];
assign g[9886] = a[12] & g[5790];
assign g[13981] = b[12] & g[5790];
assign g[9887] = a[12] & g[5791];
assign g[13982] = b[12] & g[5791];
assign g[9888] = a[12] & g[5792];
assign g[13983] = b[12] & g[5792];
assign g[9889] = a[12] & g[5793];
assign g[13984] = b[12] & g[5793];
assign g[9890] = a[12] & g[5794];
assign g[13985] = b[12] & g[5794];
assign g[9891] = a[12] & g[5795];
assign g[13986] = b[12] & g[5795];
assign g[9892] = a[12] & g[5796];
assign g[13987] = b[12] & g[5796];
assign g[9893] = a[12] & g[5797];
assign g[13988] = b[12] & g[5797];
assign g[9894] = a[12] & g[5798];
assign g[13989] = b[12] & g[5798];
assign g[9895] = a[12] & g[5799];
assign g[13990] = b[12] & g[5799];
assign g[9896] = a[12] & g[5800];
assign g[13991] = b[12] & g[5800];
assign g[9897] = a[12] & g[5801];
assign g[13992] = b[12] & g[5801];
assign g[9898] = a[12] & g[5802];
assign g[13993] = b[12] & g[5802];
assign g[9899] = a[12] & g[5803];
assign g[13994] = b[12] & g[5803];
assign g[9900] = a[12] & g[5804];
assign g[13995] = b[12] & g[5804];
assign g[9901] = a[12] & g[5805];
assign g[13996] = b[12] & g[5805];
assign g[9902] = a[12] & g[5806];
assign g[13997] = b[12] & g[5806];
assign g[9903] = a[12] & g[5807];
assign g[13998] = b[12] & g[5807];
assign g[9904] = a[12] & g[5808];
assign g[13999] = b[12] & g[5808];
assign g[9905] = a[12] & g[5809];
assign g[14000] = b[12] & g[5809];
assign g[9906] = a[12] & g[5810];
assign g[14001] = b[12] & g[5810];
assign g[9907] = a[12] & g[5811];
assign g[14002] = b[12] & g[5811];
assign g[9908] = a[12] & g[5812];
assign g[14003] = b[12] & g[5812];
assign g[9909] = a[12] & g[5813];
assign g[14004] = b[12] & g[5813];
assign g[9910] = a[12] & g[5814];
assign g[14005] = b[12] & g[5814];
assign g[9911] = a[12] & g[5815];
assign g[14006] = b[12] & g[5815];
assign g[9912] = a[12] & g[5816];
assign g[14007] = b[12] & g[5816];
assign g[9913] = a[12] & g[5817];
assign g[14008] = b[12] & g[5817];
assign g[9914] = a[12] & g[5818];
assign g[14009] = b[12] & g[5818];
assign g[9915] = a[12] & g[5819];
assign g[14010] = b[12] & g[5819];
assign g[9916] = a[12] & g[5820];
assign g[14011] = b[12] & g[5820];
assign g[9917] = a[12] & g[5821];
assign g[14012] = b[12] & g[5821];
assign g[9918] = a[12] & g[5822];
assign g[14013] = b[12] & g[5822];
assign g[9919] = a[12] & g[5823];
assign g[14014] = b[12] & g[5823];
assign g[9920] = a[12] & g[5824];
assign g[14015] = b[12] & g[5824];
assign g[9921] = a[12] & g[5825];
assign g[14016] = b[12] & g[5825];
assign g[9922] = a[12] & g[5826];
assign g[14017] = b[12] & g[5826];
assign g[9923] = a[12] & g[5827];
assign g[14018] = b[12] & g[5827];
assign g[9924] = a[12] & g[5828];
assign g[14019] = b[12] & g[5828];
assign g[9925] = a[12] & g[5829];
assign g[14020] = b[12] & g[5829];
assign g[9926] = a[12] & g[5830];
assign g[14021] = b[12] & g[5830];
assign g[9927] = a[12] & g[5831];
assign g[14022] = b[12] & g[5831];
assign g[9928] = a[12] & g[5832];
assign g[14023] = b[12] & g[5832];
assign g[9929] = a[12] & g[5833];
assign g[14024] = b[12] & g[5833];
assign g[9930] = a[12] & g[5834];
assign g[14025] = b[12] & g[5834];
assign g[9931] = a[12] & g[5835];
assign g[14026] = b[12] & g[5835];
assign g[9932] = a[12] & g[5836];
assign g[14027] = b[12] & g[5836];
assign g[9933] = a[12] & g[5837];
assign g[14028] = b[12] & g[5837];
assign g[9934] = a[12] & g[5838];
assign g[14029] = b[12] & g[5838];
assign g[9935] = a[12] & g[5839];
assign g[14030] = b[12] & g[5839];
assign g[9936] = a[12] & g[5840];
assign g[14031] = b[12] & g[5840];
assign g[9937] = a[12] & g[5841];
assign g[14032] = b[12] & g[5841];
assign g[9938] = a[12] & g[5842];
assign g[14033] = b[12] & g[5842];
assign g[9939] = a[12] & g[5843];
assign g[14034] = b[12] & g[5843];
assign g[9940] = a[12] & g[5844];
assign g[14035] = b[12] & g[5844];
assign g[9941] = a[12] & g[5845];
assign g[14036] = b[12] & g[5845];
assign g[9942] = a[12] & g[5846];
assign g[14037] = b[12] & g[5846];
assign g[9943] = a[12] & g[5847];
assign g[14038] = b[12] & g[5847];
assign g[9944] = a[12] & g[5848];
assign g[14039] = b[12] & g[5848];
assign g[9945] = a[12] & g[5849];
assign g[14040] = b[12] & g[5849];
assign g[9946] = a[12] & g[5850];
assign g[14041] = b[12] & g[5850];
assign g[9947] = a[12] & g[5851];
assign g[14042] = b[12] & g[5851];
assign g[9948] = a[12] & g[5852];
assign g[14043] = b[12] & g[5852];
assign g[9949] = a[12] & g[5853];
assign g[14044] = b[12] & g[5853];
assign g[9950] = a[12] & g[5854];
assign g[14045] = b[12] & g[5854];
assign g[9951] = a[12] & g[5855];
assign g[14046] = b[12] & g[5855];
assign g[9952] = a[12] & g[5856];
assign g[14047] = b[12] & g[5856];
assign g[9953] = a[12] & g[5857];
assign g[14048] = b[12] & g[5857];
assign g[9954] = a[12] & g[5858];
assign g[14049] = b[12] & g[5858];
assign g[9955] = a[12] & g[5859];
assign g[14050] = b[12] & g[5859];
assign g[9956] = a[12] & g[5860];
assign g[14051] = b[12] & g[5860];
assign g[9957] = a[12] & g[5861];
assign g[14052] = b[12] & g[5861];
assign g[9958] = a[12] & g[5862];
assign g[14053] = b[12] & g[5862];
assign g[9959] = a[12] & g[5863];
assign g[14054] = b[12] & g[5863];
assign g[9960] = a[12] & g[5864];
assign g[14055] = b[12] & g[5864];
assign g[9961] = a[12] & g[5865];
assign g[14056] = b[12] & g[5865];
assign g[9962] = a[12] & g[5866];
assign g[14057] = b[12] & g[5866];
assign g[9963] = a[12] & g[5867];
assign g[14058] = b[12] & g[5867];
assign g[9964] = a[12] & g[5868];
assign g[14059] = b[12] & g[5868];
assign g[9965] = a[12] & g[5869];
assign g[14060] = b[12] & g[5869];
assign g[9966] = a[12] & g[5870];
assign g[14061] = b[12] & g[5870];
assign g[9967] = a[12] & g[5871];
assign g[14062] = b[12] & g[5871];
assign g[9968] = a[12] & g[5872];
assign g[14063] = b[12] & g[5872];
assign g[9969] = a[12] & g[5873];
assign g[14064] = b[12] & g[5873];
assign g[9970] = a[12] & g[5874];
assign g[14065] = b[12] & g[5874];
assign g[9971] = a[12] & g[5875];
assign g[14066] = b[12] & g[5875];
assign g[9972] = a[12] & g[5876];
assign g[14067] = b[12] & g[5876];
assign g[9973] = a[12] & g[5877];
assign g[14068] = b[12] & g[5877];
assign g[9974] = a[12] & g[5878];
assign g[14069] = b[12] & g[5878];
assign g[9975] = a[12] & g[5879];
assign g[14070] = b[12] & g[5879];
assign g[9976] = a[12] & g[5880];
assign g[14071] = b[12] & g[5880];
assign g[9977] = a[12] & g[5881];
assign g[14072] = b[12] & g[5881];
assign g[9978] = a[12] & g[5882];
assign g[14073] = b[12] & g[5882];
assign g[9979] = a[12] & g[5883];
assign g[14074] = b[12] & g[5883];
assign g[9980] = a[12] & g[5884];
assign g[14075] = b[12] & g[5884];
assign g[9981] = a[12] & g[5885];
assign g[14076] = b[12] & g[5885];
assign g[9982] = a[12] & g[5886];
assign g[14077] = b[12] & g[5886];
assign g[9983] = a[12] & g[5887];
assign g[14078] = b[12] & g[5887];
assign g[9984] = a[12] & g[5888];
assign g[14079] = b[12] & g[5888];
assign g[9985] = a[12] & g[5889];
assign g[14080] = b[12] & g[5889];
assign g[9986] = a[12] & g[5890];
assign g[14081] = b[12] & g[5890];
assign g[9987] = a[12] & g[5891];
assign g[14082] = b[12] & g[5891];
assign g[9988] = a[12] & g[5892];
assign g[14083] = b[12] & g[5892];
assign g[9989] = a[12] & g[5893];
assign g[14084] = b[12] & g[5893];
assign g[9990] = a[12] & g[5894];
assign g[14085] = b[12] & g[5894];
assign g[9991] = a[12] & g[5895];
assign g[14086] = b[12] & g[5895];
assign g[9992] = a[12] & g[5896];
assign g[14087] = b[12] & g[5896];
assign g[9993] = a[12] & g[5897];
assign g[14088] = b[12] & g[5897];
assign g[9994] = a[12] & g[5898];
assign g[14089] = b[12] & g[5898];
assign g[9995] = a[12] & g[5899];
assign g[14090] = b[12] & g[5899];
assign g[9996] = a[12] & g[5900];
assign g[14091] = b[12] & g[5900];
assign g[9997] = a[12] & g[5901];
assign g[14092] = b[12] & g[5901];
assign g[9998] = a[12] & g[5902];
assign g[14093] = b[12] & g[5902];
assign g[9999] = a[12] & g[5903];
assign g[14094] = b[12] & g[5903];
assign g[10000] = a[12] & g[5904];
assign g[14095] = b[12] & g[5904];
assign g[10001] = a[12] & g[5905];
assign g[14096] = b[12] & g[5905];
assign g[10002] = a[12] & g[5906];
assign g[14097] = b[12] & g[5906];
assign g[10003] = a[12] & g[5907];
assign g[14098] = b[12] & g[5907];
assign g[10004] = a[12] & g[5908];
assign g[14099] = b[12] & g[5908];
assign g[10005] = a[12] & g[5909];
assign g[14100] = b[12] & g[5909];
assign g[10006] = a[12] & g[5910];
assign g[14101] = b[12] & g[5910];
assign g[10007] = a[12] & g[5911];
assign g[14102] = b[12] & g[5911];
assign g[10008] = a[12] & g[5912];
assign g[14103] = b[12] & g[5912];
assign g[10009] = a[12] & g[5913];
assign g[14104] = b[12] & g[5913];
assign g[10010] = a[12] & g[5914];
assign g[14105] = b[12] & g[5914];
assign g[10011] = a[12] & g[5915];
assign g[14106] = b[12] & g[5915];
assign g[10012] = a[12] & g[5916];
assign g[14107] = b[12] & g[5916];
assign g[10013] = a[12] & g[5917];
assign g[14108] = b[12] & g[5917];
assign g[10014] = a[12] & g[5918];
assign g[14109] = b[12] & g[5918];
assign g[10015] = a[12] & g[5919];
assign g[14110] = b[12] & g[5919];
assign g[10016] = a[12] & g[5920];
assign g[14111] = b[12] & g[5920];
assign g[10017] = a[12] & g[5921];
assign g[14112] = b[12] & g[5921];
assign g[10018] = a[12] & g[5922];
assign g[14113] = b[12] & g[5922];
assign g[10019] = a[12] & g[5923];
assign g[14114] = b[12] & g[5923];
assign g[10020] = a[12] & g[5924];
assign g[14115] = b[12] & g[5924];
assign g[10021] = a[12] & g[5925];
assign g[14116] = b[12] & g[5925];
assign g[10022] = a[12] & g[5926];
assign g[14117] = b[12] & g[5926];
assign g[10023] = a[12] & g[5927];
assign g[14118] = b[12] & g[5927];
assign g[10024] = a[12] & g[5928];
assign g[14119] = b[12] & g[5928];
assign g[10025] = a[12] & g[5929];
assign g[14120] = b[12] & g[5929];
assign g[10026] = a[12] & g[5930];
assign g[14121] = b[12] & g[5930];
assign g[10027] = a[12] & g[5931];
assign g[14122] = b[12] & g[5931];
assign g[10028] = a[12] & g[5932];
assign g[14123] = b[12] & g[5932];
assign g[10029] = a[12] & g[5933];
assign g[14124] = b[12] & g[5933];
assign g[10030] = a[12] & g[5934];
assign g[14125] = b[12] & g[5934];
assign g[10031] = a[12] & g[5935];
assign g[14126] = b[12] & g[5935];
assign g[10032] = a[12] & g[5936];
assign g[14127] = b[12] & g[5936];
assign g[10033] = a[12] & g[5937];
assign g[14128] = b[12] & g[5937];
assign g[10034] = a[12] & g[5938];
assign g[14129] = b[12] & g[5938];
assign g[10035] = a[12] & g[5939];
assign g[14130] = b[12] & g[5939];
assign g[10036] = a[12] & g[5940];
assign g[14131] = b[12] & g[5940];
assign g[10037] = a[12] & g[5941];
assign g[14132] = b[12] & g[5941];
assign g[10038] = a[12] & g[5942];
assign g[14133] = b[12] & g[5942];
assign g[10039] = a[12] & g[5943];
assign g[14134] = b[12] & g[5943];
assign g[10040] = a[12] & g[5944];
assign g[14135] = b[12] & g[5944];
assign g[10041] = a[12] & g[5945];
assign g[14136] = b[12] & g[5945];
assign g[10042] = a[12] & g[5946];
assign g[14137] = b[12] & g[5946];
assign g[10043] = a[12] & g[5947];
assign g[14138] = b[12] & g[5947];
assign g[10044] = a[12] & g[5948];
assign g[14139] = b[12] & g[5948];
assign g[10045] = a[12] & g[5949];
assign g[14140] = b[12] & g[5949];
assign g[10046] = a[12] & g[5950];
assign g[14141] = b[12] & g[5950];
assign g[10047] = a[12] & g[5951];
assign g[14142] = b[12] & g[5951];
assign g[10048] = a[12] & g[5952];
assign g[14143] = b[12] & g[5952];
assign g[10049] = a[12] & g[5953];
assign g[14144] = b[12] & g[5953];
assign g[10050] = a[12] & g[5954];
assign g[14145] = b[12] & g[5954];
assign g[10051] = a[12] & g[5955];
assign g[14146] = b[12] & g[5955];
assign g[10052] = a[12] & g[5956];
assign g[14147] = b[12] & g[5956];
assign g[10053] = a[12] & g[5957];
assign g[14148] = b[12] & g[5957];
assign g[10054] = a[12] & g[5958];
assign g[14149] = b[12] & g[5958];
assign g[10055] = a[12] & g[5959];
assign g[14150] = b[12] & g[5959];
assign g[10056] = a[12] & g[5960];
assign g[14151] = b[12] & g[5960];
assign g[10057] = a[12] & g[5961];
assign g[14152] = b[12] & g[5961];
assign g[10058] = a[12] & g[5962];
assign g[14153] = b[12] & g[5962];
assign g[10059] = a[12] & g[5963];
assign g[14154] = b[12] & g[5963];
assign g[10060] = a[12] & g[5964];
assign g[14155] = b[12] & g[5964];
assign g[10061] = a[12] & g[5965];
assign g[14156] = b[12] & g[5965];
assign g[10062] = a[12] & g[5966];
assign g[14157] = b[12] & g[5966];
assign g[10063] = a[12] & g[5967];
assign g[14158] = b[12] & g[5967];
assign g[10064] = a[12] & g[5968];
assign g[14159] = b[12] & g[5968];
assign g[10065] = a[12] & g[5969];
assign g[14160] = b[12] & g[5969];
assign g[10066] = a[12] & g[5970];
assign g[14161] = b[12] & g[5970];
assign g[10067] = a[12] & g[5971];
assign g[14162] = b[12] & g[5971];
assign g[10068] = a[12] & g[5972];
assign g[14163] = b[12] & g[5972];
assign g[10069] = a[12] & g[5973];
assign g[14164] = b[12] & g[5973];
assign g[10070] = a[12] & g[5974];
assign g[14165] = b[12] & g[5974];
assign g[10071] = a[12] & g[5975];
assign g[14166] = b[12] & g[5975];
assign g[10072] = a[12] & g[5976];
assign g[14167] = b[12] & g[5976];
assign g[10073] = a[12] & g[5977];
assign g[14168] = b[12] & g[5977];
assign g[10074] = a[12] & g[5978];
assign g[14169] = b[12] & g[5978];
assign g[10075] = a[12] & g[5979];
assign g[14170] = b[12] & g[5979];
assign g[10076] = a[12] & g[5980];
assign g[14171] = b[12] & g[5980];
assign g[10077] = a[12] & g[5981];
assign g[14172] = b[12] & g[5981];
assign g[10078] = a[12] & g[5982];
assign g[14173] = b[12] & g[5982];
assign g[10079] = a[12] & g[5983];
assign g[14174] = b[12] & g[5983];
assign g[10080] = a[12] & g[5984];
assign g[14175] = b[12] & g[5984];
assign g[10081] = a[12] & g[5985];
assign g[14176] = b[12] & g[5985];
assign g[10082] = a[12] & g[5986];
assign g[14177] = b[12] & g[5986];
assign g[10083] = a[12] & g[5987];
assign g[14178] = b[12] & g[5987];
assign g[10084] = a[12] & g[5988];
assign g[14179] = b[12] & g[5988];
assign g[10085] = a[12] & g[5989];
assign g[14180] = b[12] & g[5989];
assign g[10086] = a[12] & g[5990];
assign g[14181] = b[12] & g[5990];
assign g[10087] = a[12] & g[5991];
assign g[14182] = b[12] & g[5991];
assign g[10088] = a[12] & g[5992];
assign g[14183] = b[12] & g[5992];
assign g[10089] = a[12] & g[5993];
assign g[14184] = b[12] & g[5993];
assign g[10090] = a[12] & g[5994];
assign g[14185] = b[12] & g[5994];
assign g[10091] = a[12] & g[5995];
assign g[14186] = b[12] & g[5995];
assign g[10092] = a[12] & g[5996];
assign g[14187] = b[12] & g[5996];
assign g[10093] = a[12] & g[5997];
assign g[14188] = b[12] & g[5997];
assign g[10094] = a[12] & g[5998];
assign g[14189] = b[12] & g[5998];
assign g[10095] = a[12] & g[5999];
assign g[14190] = b[12] & g[5999];
assign g[10096] = a[12] & g[6000];
assign g[14191] = b[12] & g[6000];
assign g[10097] = a[12] & g[6001];
assign g[14192] = b[12] & g[6001];
assign g[10098] = a[12] & g[6002];
assign g[14193] = b[12] & g[6002];
assign g[10099] = a[12] & g[6003];
assign g[14194] = b[12] & g[6003];
assign g[10100] = a[12] & g[6004];
assign g[14195] = b[12] & g[6004];
assign g[10101] = a[12] & g[6005];
assign g[14196] = b[12] & g[6005];
assign g[10102] = a[12] & g[6006];
assign g[14197] = b[12] & g[6006];
assign g[10103] = a[12] & g[6007];
assign g[14198] = b[12] & g[6007];
assign g[10104] = a[12] & g[6008];
assign g[14199] = b[12] & g[6008];
assign g[10105] = a[12] & g[6009];
assign g[14200] = b[12] & g[6009];
assign g[10106] = a[12] & g[6010];
assign g[14201] = b[12] & g[6010];
assign g[10107] = a[12] & g[6011];
assign g[14202] = b[12] & g[6011];
assign g[10108] = a[12] & g[6012];
assign g[14203] = b[12] & g[6012];
assign g[10109] = a[12] & g[6013];
assign g[14204] = b[12] & g[6013];
assign g[10110] = a[12] & g[6014];
assign g[14205] = b[12] & g[6014];
assign g[10111] = a[12] & g[6015];
assign g[14206] = b[12] & g[6015];
assign g[10112] = a[12] & g[6016];
assign g[14207] = b[12] & g[6016];
assign g[10113] = a[12] & g[6017];
assign g[14208] = b[12] & g[6017];
assign g[10114] = a[12] & g[6018];
assign g[14209] = b[12] & g[6018];
assign g[10115] = a[12] & g[6019];
assign g[14210] = b[12] & g[6019];
assign g[10116] = a[12] & g[6020];
assign g[14211] = b[12] & g[6020];
assign g[10117] = a[12] & g[6021];
assign g[14212] = b[12] & g[6021];
assign g[10118] = a[12] & g[6022];
assign g[14213] = b[12] & g[6022];
assign g[10119] = a[12] & g[6023];
assign g[14214] = b[12] & g[6023];
assign g[10120] = a[12] & g[6024];
assign g[14215] = b[12] & g[6024];
assign g[10121] = a[12] & g[6025];
assign g[14216] = b[12] & g[6025];
assign g[10122] = a[12] & g[6026];
assign g[14217] = b[12] & g[6026];
assign g[10123] = a[12] & g[6027];
assign g[14218] = b[12] & g[6027];
assign g[10124] = a[12] & g[6028];
assign g[14219] = b[12] & g[6028];
assign g[10125] = a[12] & g[6029];
assign g[14220] = b[12] & g[6029];
assign g[10126] = a[12] & g[6030];
assign g[14221] = b[12] & g[6030];
assign g[10127] = a[12] & g[6031];
assign g[14222] = b[12] & g[6031];
assign g[10128] = a[12] & g[6032];
assign g[14223] = b[12] & g[6032];
assign g[10129] = a[12] & g[6033];
assign g[14224] = b[12] & g[6033];
assign g[10130] = a[12] & g[6034];
assign g[14225] = b[12] & g[6034];
assign g[10131] = a[12] & g[6035];
assign g[14226] = b[12] & g[6035];
assign g[10132] = a[12] & g[6036];
assign g[14227] = b[12] & g[6036];
assign g[10133] = a[12] & g[6037];
assign g[14228] = b[12] & g[6037];
assign g[10134] = a[12] & g[6038];
assign g[14229] = b[12] & g[6038];
assign g[10135] = a[12] & g[6039];
assign g[14230] = b[12] & g[6039];
assign g[10136] = a[12] & g[6040];
assign g[14231] = b[12] & g[6040];
assign g[10137] = a[12] & g[6041];
assign g[14232] = b[12] & g[6041];
assign g[10138] = a[12] & g[6042];
assign g[14233] = b[12] & g[6042];
assign g[10139] = a[12] & g[6043];
assign g[14234] = b[12] & g[6043];
assign g[10140] = a[12] & g[6044];
assign g[14235] = b[12] & g[6044];
assign g[10141] = a[12] & g[6045];
assign g[14236] = b[12] & g[6045];
assign g[10142] = a[12] & g[6046];
assign g[14237] = b[12] & g[6046];
assign g[10143] = a[12] & g[6047];
assign g[14238] = b[12] & g[6047];
assign g[10144] = a[12] & g[6048];
assign g[14239] = b[12] & g[6048];
assign g[10145] = a[12] & g[6049];
assign g[14240] = b[12] & g[6049];
assign g[10146] = a[12] & g[6050];
assign g[14241] = b[12] & g[6050];
assign g[10147] = a[12] & g[6051];
assign g[14242] = b[12] & g[6051];
assign g[10148] = a[12] & g[6052];
assign g[14243] = b[12] & g[6052];
assign g[10149] = a[12] & g[6053];
assign g[14244] = b[12] & g[6053];
assign g[10150] = a[12] & g[6054];
assign g[14245] = b[12] & g[6054];
assign g[10151] = a[12] & g[6055];
assign g[14246] = b[12] & g[6055];
assign g[10152] = a[12] & g[6056];
assign g[14247] = b[12] & g[6056];
assign g[10153] = a[12] & g[6057];
assign g[14248] = b[12] & g[6057];
assign g[10154] = a[12] & g[6058];
assign g[14249] = b[12] & g[6058];
assign g[10155] = a[12] & g[6059];
assign g[14250] = b[12] & g[6059];
assign g[10156] = a[12] & g[6060];
assign g[14251] = b[12] & g[6060];
assign g[10157] = a[12] & g[6061];
assign g[14252] = b[12] & g[6061];
assign g[10158] = a[12] & g[6062];
assign g[14253] = b[12] & g[6062];
assign g[10159] = a[12] & g[6063];
assign g[14254] = b[12] & g[6063];
assign g[10160] = a[12] & g[6064];
assign g[14255] = b[12] & g[6064];
assign g[10161] = a[12] & g[6065];
assign g[14256] = b[12] & g[6065];
assign g[10162] = a[12] & g[6066];
assign g[14257] = b[12] & g[6066];
assign g[10163] = a[12] & g[6067];
assign g[14258] = b[12] & g[6067];
assign g[10164] = a[12] & g[6068];
assign g[14259] = b[12] & g[6068];
assign g[10165] = a[12] & g[6069];
assign g[14260] = b[12] & g[6069];
assign g[10166] = a[12] & g[6070];
assign g[14261] = b[12] & g[6070];
assign g[10167] = a[12] & g[6071];
assign g[14262] = b[12] & g[6071];
assign g[10168] = a[12] & g[6072];
assign g[14263] = b[12] & g[6072];
assign g[10169] = a[12] & g[6073];
assign g[14264] = b[12] & g[6073];
assign g[10170] = a[12] & g[6074];
assign g[14265] = b[12] & g[6074];
assign g[10171] = a[12] & g[6075];
assign g[14266] = b[12] & g[6075];
assign g[10172] = a[12] & g[6076];
assign g[14267] = b[12] & g[6076];
assign g[10173] = a[12] & g[6077];
assign g[14268] = b[12] & g[6077];
assign g[10174] = a[12] & g[6078];
assign g[14269] = b[12] & g[6078];
assign g[10175] = a[12] & g[6079];
assign g[14270] = b[12] & g[6079];
assign g[10176] = a[12] & g[6080];
assign g[14271] = b[12] & g[6080];
assign g[10177] = a[12] & g[6081];
assign g[14272] = b[12] & g[6081];
assign g[10178] = a[12] & g[6082];
assign g[14273] = b[12] & g[6082];
assign g[10179] = a[12] & g[6083];
assign g[14274] = b[12] & g[6083];
assign g[10180] = a[12] & g[6084];
assign g[14275] = b[12] & g[6084];
assign g[10181] = a[12] & g[6085];
assign g[14276] = b[12] & g[6085];
assign g[10182] = a[12] & g[6086];
assign g[14277] = b[12] & g[6086];
assign g[10183] = a[12] & g[6087];
assign g[14278] = b[12] & g[6087];
assign g[10184] = a[12] & g[6088];
assign g[14279] = b[12] & g[6088];
assign g[10185] = a[12] & g[6089];
assign g[14280] = b[12] & g[6089];
assign g[10186] = a[12] & g[6090];
assign g[14281] = b[12] & g[6090];
assign g[10187] = a[12] & g[6091];
assign g[14282] = b[12] & g[6091];
assign g[10188] = a[12] & g[6092];
assign g[14283] = b[12] & g[6092];
assign g[10189] = a[12] & g[6093];
assign g[14284] = b[12] & g[6093];
assign g[10190] = a[12] & g[6094];
assign g[14285] = b[12] & g[6094];
assign g[10191] = a[12] & g[6095];
assign g[14286] = b[12] & g[6095];
assign g[10192] = a[12] & g[6096];
assign g[14287] = b[12] & g[6096];
assign g[10193] = a[12] & g[6097];
assign g[14288] = b[12] & g[6097];
assign g[10194] = a[12] & g[6098];
assign g[14289] = b[12] & g[6098];
assign g[10195] = a[12] & g[6099];
assign g[14290] = b[12] & g[6099];
assign g[10196] = a[12] & g[6100];
assign g[14291] = b[12] & g[6100];
assign g[10197] = a[12] & g[6101];
assign g[14292] = b[12] & g[6101];
assign g[10198] = a[12] & g[6102];
assign g[14293] = b[12] & g[6102];
assign g[10199] = a[12] & g[6103];
assign g[14294] = b[12] & g[6103];
assign g[10200] = a[12] & g[6104];
assign g[14295] = b[12] & g[6104];
assign g[10201] = a[12] & g[6105];
assign g[14296] = b[12] & g[6105];
assign g[10202] = a[12] & g[6106];
assign g[14297] = b[12] & g[6106];
assign g[10203] = a[12] & g[6107];
assign g[14298] = b[12] & g[6107];
assign g[10204] = a[12] & g[6108];
assign g[14299] = b[12] & g[6108];
assign g[10205] = a[12] & g[6109];
assign g[14300] = b[12] & g[6109];
assign g[10206] = a[12] & g[6110];
assign g[14301] = b[12] & g[6110];
assign g[10207] = a[12] & g[6111];
assign g[14302] = b[12] & g[6111];
assign g[10208] = a[12] & g[6112];
assign g[14303] = b[12] & g[6112];
assign g[10209] = a[12] & g[6113];
assign g[14304] = b[12] & g[6113];
assign g[10210] = a[12] & g[6114];
assign g[14305] = b[12] & g[6114];
assign g[10211] = a[12] & g[6115];
assign g[14306] = b[12] & g[6115];
assign g[10212] = a[12] & g[6116];
assign g[14307] = b[12] & g[6116];
assign g[10213] = a[12] & g[6117];
assign g[14308] = b[12] & g[6117];
assign g[10214] = a[12] & g[6118];
assign g[14309] = b[12] & g[6118];
assign g[10215] = a[12] & g[6119];
assign g[14310] = b[12] & g[6119];
assign g[10216] = a[12] & g[6120];
assign g[14311] = b[12] & g[6120];
assign g[10217] = a[12] & g[6121];
assign g[14312] = b[12] & g[6121];
assign g[10218] = a[12] & g[6122];
assign g[14313] = b[12] & g[6122];
assign g[10219] = a[12] & g[6123];
assign g[14314] = b[12] & g[6123];
assign g[10220] = a[12] & g[6124];
assign g[14315] = b[12] & g[6124];
assign g[10221] = a[12] & g[6125];
assign g[14316] = b[12] & g[6125];
assign g[10222] = a[12] & g[6126];
assign g[14317] = b[12] & g[6126];
assign g[10223] = a[12] & g[6127];
assign g[14318] = b[12] & g[6127];
assign g[10224] = a[12] & g[6128];
assign g[14319] = b[12] & g[6128];
assign g[10225] = a[12] & g[6129];
assign g[14320] = b[12] & g[6129];
assign g[10226] = a[12] & g[6130];
assign g[14321] = b[12] & g[6130];
assign g[10227] = a[12] & g[6131];
assign g[14322] = b[12] & g[6131];
assign g[10228] = a[12] & g[6132];
assign g[14323] = b[12] & g[6132];
assign g[10229] = a[12] & g[6133];
assign g[14324] = b[12] & g[6133];
assign g[10230] = a[12] & g[6134];
assign g[14325] = b[12] & g[6134];
assign g[10231] = a[12] & g[6135];
assign g[14326] = b[12] & g[6135];
assign g[10232] = a[12] & g[6136];
assign g[14327] = b[12] & g[6136];
assign g[10233] = a[12] & g[6137];
assign g[14328] = b[12] & g[6137];
assign g[10234] = a[12] & g[6138];
assign g[14329] = b[12] & g[6138];
assign g[10235] = a[12] & g[6139];
assign g[14330] = b[12] & g[6139];
assign g[10236] = a[12] & g[6140];
assign g[14331] = b[12] & g[6140];
assign g[10237] = a[12] & g[6141];
assign g[14332] = b[12] & g[6141];
assign g[10238] = a[12] & g[6142];
assign g[14333] = b[12] & g[6142];
assign g[10239] = a[12] & g[6143];
assign g[14334] = b[12] & g[6143];
assign g[10240] = a[12] & g[6144];
assign g[14335] = b[12] & g[6144];
assign g[10241] = a[12] & g[6145];
assign g[14336] = b[12] & g[6145];
assign g[10242] = a[12] & g[6146];
assign g[14337] = b[12] & g[6146];
assign g[10243] = a[12] & g[6147];
assign g[14338] = b[12] & g[6147];
assign g[10244] = a[12] & g[6148];
assign g[14339] = b[12] & g[6148];
assign g[10245] = a[12] & g[6149];
assign g[14340] = b[12] & g[6149];
assign g[10246] = a[12] & g[6150];
assign g[14341] = b[12] & g[6150];
assign g[10247] = a[12] & g[6151];
assign g[14342] = b[12] & g[6151];
assign g[10248] = a[12] & g[6152];
assign g[14343] = b[12] & g[6152];
assign g[10249] = a[12] & g[6153];
assign g[14344] = b[12] & g[6153];
assign g[10250] = a[12] & g[6154];
assign g[14345] = b[12] & g[6154];
assign g[10251] = a[12] & g[6155];
assign g[14346] = b[12] & g[6155];
assign g[10252] = a[12] & g[6156];
assign g[14347] = b[12] & g[6156];
assign g[10253] = a[12] & g[6157];
assign g[14348] = b[12] & g[6157];
assign g[10254] = a[12] & g[6158];
assign g[14349] = b[12] & g[6158];
assign g[10255] = a[12] & g[6159];
assign g[14350] = b[12] & g[6159];
assign g[10256] = a[12] & g[6160];
assign g[14351] = b[12] & g[6160];
assign g[10257] = a[12] & g[6161];
assign g[14352] = b[12] & g[6161];
assign g[10258] = a[12] & g[6162];
assign g[14353] = b[12] & g[6162];
assign g[10259] = a[12] & g[6163];
assign g[14354] = b[12] & g[6163];
assign g[10260] = a[12] & g[6164];
assign g[14355] = b[12] & g[6164];
assign g[10261] = a[12] & g[6165];
assign g[14356] = b[12] & g[6165];
assign g[10262] = a[12] & g[6166];
assign g[14357] = b[12] & g[6166];
assign g[10263] = a[12] & g[6167];
assign g[14358] = b[12] & g[6167];
assign g[10264] = a[12] & g[6168];
assign g[14359] = b[12] & g[6168];
assign g[10265] = a[12] & g[6169];
assign g[14360] = b[12] & g[6169];
assign g[10266] = a[12] & g[6170];
assign g[14361] = b[12] & g[6170];
assign g[10267] = a[12] & g[6171];
assign g[14362] = b[12] & g[6171];
assign g[10268] = a[12] & g[6172];
assign g[14363] = b[12] & g[6172];
assign g[10269] = a[12] & g[6173];
assign g[14364] = b[12] & g[6173];
assign g[10270] = a[12] & g[6174];
assign g[14365] = b[12] & g[6174];
assign g[10271] = a[12] & g[6175];
assign g[14366] = b[12] & g[6175];
assign g[10272] = a[12] & g[6176];
assign g[14367] = b[12] & g[6176];
assign g[10273] = a[12] & g[6177];
assign g[14368] = b[12] & g[6177];
assign g[10274] = a[12] & g[6178];
assign g[14369] = b[12] & g[6178];
assign g[10275] = a[12] & g[6179];
assign g[14370] = b[12] & g[6179];
assign g[10276] = a[12] & g[6180];
assign g[14371] = b[12] & g[6180];
assign g[10277] = a[12] & g[6181];
assign g[14372] = b[12] & g[6181];
assign g[10278] = a[12] & g[6182];
assign g[14373] = b[12] & g[6182];
assign g[10279] = a[12] & g[6183];
assign g[14374] = b[12] & g[6183];
assign g[10280] = a[12] & g[6184];
assign g[14375] = b[12] & g[6184];
assign g[10281] = a[12] & g[6185];
assign g[14376] = b[12] & g[6185];
assign g[10282] = a[12] & g[6186];
assign g[14377] = b[12] & g[6186];
assign g[10283] = a[12] & g[6187];
assign g[14378] = b[12] & g[6187];
assign g[10284] = a[12] & g[6188];
assign g[14379] = b[12] & g[6188];
assign g[10285] = a[12] & g[6189];
assign g[14380] = b[12] & g[6189];
assign g[10286] = a[12] & g[6190];
assign g[14381] = b[12] & g[6190];
assign g[10287] = a[12] & g[6191];
assign g[14382] = b[12] & g[6191];
assign g[10288] = a[12] & g[6192];
assign g[14383] = b[12] & g[6192];
assign g[10289] = a[12] & g[6193];
assign g[14384] = b[12] & g[6193];
assign g[10290] = a[12] & g[6194];
assign g[14385] = b[12] & g[6194];
assign g[10291] = a[12] & g[6195];
assign g[14386] = b[12] & g[6195];
assign g[10292] = a[12] & g[6196];
assign g[14387] = b[12] & g[6196];
assign g[10293] = a[12] & g[6197];
assign g[14388] = b[12] & g[6197];
assign g[10294] = a[12] & g[6198];
assign g[14389] = b[12] & g[6198];
assign g[10295] = a[12] & g[6199];
assign g[14390] = b[12] & g[6199];
assign g[10296] = a[12] & g[6200];
assign g[14391] = b[12] & g[6200];
assign g[10297] = a[12] & g[6201];
assign g[14392] = b[12] & g[6201];
assign g[10298] = a[12] & g[6202];
assign g[14393] = b[12] & g[6202];
assign g[10299] = a[12] & g[6203];
assign g[14394] = b[12] & g[6203];
assign g[10300] = a[12] & g[6204];
assign g[14395] = b[12] & g[6204];
assign g[10301] = a[12] & g[6205];
assign g[14396] = b[12] & g[6205];
assign g[10302] = a[12] & g[6206];
assign g[14397] = b[12] & g[6206];
assign g[10303] = a[12] & g[6207];
assign g[14398] = b[12] & g[6207];
assign g[10304] = a[12] & g[6208];
assign g[14399] = b[12] & g[6208];
assign g[10305] = a[12] & g[6209];
assign g[14400] = b[12] & g[6209];
assign g[10306] = a[12] & g[6210];
assign g[14401] = b[12] & g[6210];
assign g[10307] = a[12] & g[6211];
assign g[14402] = b[12] & g[6211];
assign g[10308] = a[12] & g[6212];
assign g[14403] = b[12] & g[6212];
assign g[10309] = a[12] & g[6213];
assign g[14404] = b[12] & g[6213];
assign g[10310] = a[12] & g[6214];
assign g[14405] = b[12] & g[6214];
assign g[10311] = a[12] & g[6215];
assign g[14406] = b[12] & g[6215];
assign g[10312] = a[12] & g[6216];
assign g[14407] = b[12] & g[6216];
assign g[10313] = a[12] & g[6217];
assign g[14408] = b[12] & g[6217];
assign g[10314] = a[12] & g[6218];
assign g[14409] = b[12] & g[6218];
assign g[10315] = a[12] & g[6219];
assign g[14410] = b[12] & g[6219];
assign g[10316] = a[12] & g[6220];
assign g[14411] = b[12] & g[6220];
assign g[10317] = a[12] & g[6221];
assign g[14412] = b[12] & g[6221];
assign g[10318] = a[12] & g[6222];
assign g[14413] = b[12] & g[6222];
assign g[10319] = a[12] & g[6223];
assign g[14414] = b[12] & g[6223];
assign g[10320] = a[12] & g[6224];
assign g[14415] = b[12] & g[6224];
assign g[10321] = a[12] & g[6225];
assign g[14416] = b[12] & g[6225];
assign g[10322] = a[12] & g[6226];
assign g[14417] = b[12] & g[6226];
assign g[10323] = a[12] & g[6227];
assign g[14418] = b[12] & g[6227];
assign g[10324] = a[12] & g[6228];
assign g[14419] = b[12] & g[6228];
assign g[10325] = a[12] & g[6229];
assign g[14420] = b[12] & g[6229];
assign g[10326] = a[12] & g[6230];
assign g[14421] = b[12] & g[6230];
assign g[10327] = a[12] & g[6231];
assign g[14422] = b[12] & g[6231];
assign g[10328] = a[12] & g[6232];
assign g[14423] = b[12] & g[6232];
assign g[10329] = a[12] & g[6233];
assign g[14424] = b[12] & g[6233];
assign g[10330] = a[12] & g[6234];
assign g[14425] = b[12] & g[6234];
assign g[10331] = a[12] & g[6235];
assign g[14426] = b[12] & g[6235];
assign g[10332] = a[12] & g[6236];
assign g[14427] = b[12] & g[6236];
assign g[10333] = a[12] & g[6237];
assign g[14428] = b[12] & g[6237];
assign g[10334] = a[12] & g[6238];
assign g[14429] = b[12] & g[6238];
assign g[10335] = a[12] & g[6239];
assign g[14430] = b[12] & g[6239];
assign g[10336] = a[12] & g[6240];
assign g[14431] = b[12] & g[6240];
assign g[10337] = a[12] & g[6241];
assign g[14432] = b[12] & g[6241];
assign g[10338] = a[12] & g[6242];
assign g[14433] = b[12] & g[6242];
assign g[10339] = a[12] & g[6243];
assign g[14434] = b[12] & g[6243];
assign g[10340] = a[12] & g[6244];
assign g[14435] = b[12] & g[6244];
assign g[10341] = a[12] & g[6245];
assign g[14436] = b[12] & g[6245];
assign g[10342] = a[12] & g[6246];
assign g[14437] = b[12] & g[6246];
assign g[10343] = a[12] & g[6247];
assign g[14438] = b[12] & g[6247];
assign g[10344] = a[12] & g[6248];
assign g[14439] = b[12] & g[6248];
assign g[10345] = a[12] & g[6249];
assign g[14440] = b[12] & g[6249];
assign g[10346] = a[12] & g[6250];
assign g[14441] = b[12] & g[6250];
assign g[10347] = a[12] & g[6251];
assign g[14442] = b[12] & g[6251];
assign g[10348] = a[12] & g[6252];
assign g[14443] = b[12] & g[6252];
assign g[10349] = a[12] & g[6253];
assign g[14444] = b[12] & g[6253];
assign g[10350] = a[12] & g[6254];
assign g[14445] = b[12] & g[6254];
assign g[10351] = a[12] & g[6255];
assign g[14446] = b[12] & g[6255];
assign g[10352] = a[12] & g[6256];
assign g[14447] = b[12] & g[6256];
assign g[10353] = a[12] & g[6257];
assign g[14448] = b[12] & g[6257];
assign g[10354] = a[12] & g[6258];
assign g[14449] = b[12] & g[6258];
assign g[10355] = a[12] & g[6259];
assign g[14450] = b[12] & g[6259];
assign g[10356] = a[12] & g[6260];
assign g[14451] = b[12] & g[6260];
assign g[10357] = a[12] & g[6261];
assign g[14452] = b[12] & g[6261];
assign g[10358] = a[12] & g[6262];
assign g[14453] = b[12] & g[6262];
assign g[10359] = a[12] & g[6263];
assign g[14454] = b[12] & g[6263];
assign g[10360] = a[12] & g[6264];
assign g[14455] = b[12] & g[6264];
assign g[10361] = a[12] & g[6265];
assign g[14456] = b[12] & g[6265];
assign g[10362] = a[12] & g[6266];
assign g[14457] = b[12] & g[6266];
assign g[10363] = a[12] & g[6267];
assign g[14458] = b[12] & g[6267];
assign g[10364] = a[12] & g[6268];
assign g[14459] = b[12] & g[6268];
assign g[10365] = a[12] & g[6269];
assign g[14460] = b[12] & g[6269];
assign g[10366] = a[12] & g[6270];
assign g[14461] = b[12] & g[6270];
assign g[10367] = a[12] & g[6271];
assign g[14462] = b[12] & g[6271];
assign g[10368] = a[12] & g[6272];
assign g[14463] = b[12] & g[6272];
assign g[10369] = a[12] & g[6273];
assign g[14464] = b[12] & g[6273];
assign g[10370] = a[12] & g[6274];
assign g[14465] = b[12] & g[6274];
assign g[10371] = a[12] & g[6275];
assign g[14466] = b[12] & g[6275];
assign g[10372] = a[12] & g[6276];
assign g[14467] = b[12] & g[6276];
assign g[10373] = a[12] & g[6277];
assign g[14468] = b[12] & g[6277];
assign g[10374] = a[12] & g[6278];
assign g[14469] = b[12] & g[6278];
assign g[10375] = a[12] & g[6279];
assign g[14470] = b[12] & g[6279];
assign g[10376] = a[12] & g[6280];
assign g[14471] = b[12] & g[6280];
assign g[10377] = a[12] & g[6281];
assign g[14472] = b[12] & g[6281];
assign g[10378] = a[12] & g[6282];
assign g[14473] = b[12] & g[6282];
assign g[10379] = a[12] & g[6283];
assign g[14474] = b[12] & g[6283];
assign g[10380] = a[12] & g[6284];
assign g[14475] = b[12] & g[6284];
assign g[10381] = a[12] & g[6285];
assign g[14476] = b[12] & g[6285];
assign g[10382] = a[12] & g[6286];
assign g[14477] = b[12] & g[6286];
assign g[10383] = a[12] & g[6287];
assign g[14478] = b[12] & g[6287];
assign g[10384] = a[12] & g[6288];
assign g[14479] = b[12] & g[6288];
assign g[10385] = a[12] & g[6289];
assign g[14480] = b[12] & g[6289];
assign g[10386] = a[12] & g[6290];
assign g[14481] = b[12] & g[6290];
assign g[10387] = a[12] & g[6291];
assign g[14482] = b[12] & g[6291];
assign g[10388] = a[12] & g[6292];
assign g[14483] = b[12] & g[6292];
assign g[10389] = a[12] & g[6293];
assign g[14484] = b[12] & g[6293];
assign g[10390] = a[12] & g[6294];
assign g[14485] = b[12] & g[6294];
assign g[10391] = a[12] & g[6295];
assign g[14486] = b[12] & g[6295];
assign g[10392] = a[12] & g[6296];
assign g[14487] = b[12] & g[6296];
assign g[10393] = a[12] & g[6297];
assign g[14488] = b[12] & g[6297];
assign g[10394] = a[12] & g[6298];
assign g[14489] = b[12] & g[6298];
assign g[10395] = a[12] & g[6299];
assign g[14490] = b[12] & g[6299];
assign g[10396] = a[12] & g[6300];
assign g[14491] = b[12] & g[6300];
assign g[10397] = a[12] & g[6301];
assign g[14492] = b[12] & g[6301];
assign g[10398] = a[12] & g[6302];
assign g[14493] = b[12] & g[6302];
assign g[10399] = a[12] & g[6303];
assign g[14494] = b[12] & g[6303];
assign g[10400] = a[12] & g[6304];
assign g[14495] = b[12] & g[6304];
assign g[10401] = a[12] & g[6305];
assign g[14496] = b[12] & g[6305];
assign g[10402] = a[12] & g[6306];
assign g[14497] = b[12] & g[6306];
assign g[10403] = a[12] & g[6307];
assign g[14498] = b[12] & g[6307];
assign g[10404] = a[12] & g[6308];
assign g[14499] = b[12] & g[6308];
assign g[10405] = a[12] & g[6309];
assign g[14500] = b[12] & g[6309];
assign g[10406] = a[12] & g[6310];
assign g[14501] = b[12] & g[6310];
assign g[10407] = a[12] & g[6311];
assign g[14502] = b[12] & g[6311];
assign g[10408] = a[12] & g[6312];
assign g[14503] = b[12] & g[6312];
assign g[10409] = a[12] & g[6313];
assign g[14504] = b[12] & g[6313];
assign g[10410] = a[12] & g[6314];
assign g[14505] = b[12] & g[6314];
assign g[10411] = a[12] & g[6315];
assign g[14506] = b[12] & g[6315];
assign g[10412] = a[12] & g[6316];
assign g[14507] = b[12] & g[6316];
assign g[10413] = a[12] & g[6317];
assign g[14508] = b[12] & g[6317];
assign g[10414] = a[12] & g[6318];
assign g[14509] = b[12] & g[6318];
assign g[10415] = a[12] & g[6319];
assign g[14510] = b[12] & g[6319];
assign g[10416] = a[12] & g[6320];
assign g[14511] = b[12] & g[6320];
assign g[10417] = a[12] & g[6321];
assign g[14512] = b[12] & g[6321];
assign g[10418] = a[12] & g[6322];
assign g[14513] = b[12] & g[6322];
assign g[10419] = a[12] & g[6323];
assign g[14514] = b[12] & g[6323];
assign g[10420] = a[12] & g[6324];
assign g[14515] = b[12] & g[6324];
assign g[10421] = a[12] & g[6325];
assign g[14516] = b[12] & g[6325];
assign g[10422] = a[12] & g[6326];
assign g[14517] = b[12] & g[6326];
assign g[10423] = a[12] & g[6327];
assign g[14518] = b[12] & g[6327];
assign g[10424] = a[12] & g[6328];
assign g[14519] = b[12] & g[6328];
assign g[10425] = a[12] & g[6329];
assign g[14520] = b[12] & g[6329];
assign g[10426] = a[12] & g[6330];
assign g[14521] = b[12] & g[6330];
assign g[10427] = a[12] & g[6331];
assign g[14522] = b[12] & g[6331];
assign g[10428] = a[12] & g[6332];
assign g[14523] = b[12] & g[6332];
assign g[10429] = a[12] & g[6333];
assign g[14524] = b[12] & g[6333];
assign g[10430] = a[12] & g[6334];
assign g[14525] = b[12] & g[6334];
assign g[10431] = a[12] & g[6335];
assign g[14526] = b[12] & g[6335];
assign g[10432] = a[12] & g[6336];
assign g[14527] = b[12] & g[6336];
assign g[10433] = a[12] & g[6337];
assign g[14528] = b[12] & g[6337];
assign g[10434] = a[12] & g[6338];
assign g[14529] = b[12] & g[6338];
assign g[10435] = a[12] & g[6339];
assign g[14530] = b[12] & g[6339];
assign g[10436] = a[12] & g[6340];
assign g[14531] = b[12] & g[6340];
assign g[10437] = a[12] & g[6341];
assign g[14532] = b[12] & g[6341];
assign g[10438] = a[12] & g[6342];
assign g[14533] = b[12] & g[6342];
assign g[10439] = a[12] & g[6343];
assign g[14534] = b[12] & g[6343];
assign g[10440] = a[12] & g[6344];
assign g[14535] = b[12] & g[6344];
assign g[10441] = a[12] & g[6345];
assign g[14536] = b[12] & g[6345];
assign g[10442] = a[12] & g[6346];
assign g[14537] = b[12] & g[6346];
assign g[10443] = a[12] & g[6347];
assign g[14538] = b[12] & g[6347];
assign g[10444] = a[12] & g[6348];
assign g[14539] = b[12] & g[6348];
assign g[10445] = a[12] & g[6349];
assign g[14540] = b[12] & g[6349];
assign g[10446] = a[12] & g[6350];
assign g[14541] = b[12] & g[6350];
assign g[10447] = a[12] & g[6351];
assign g[14542] = b[12] & g[6351];
assign g[10448] = a[12] & g[6352];
assign g[14543] = b[12] & g[6352];
assign g[10449] = a[12] & g[6353];
assign g[14544] = b[12] & g[6353];
assign g[10450] = a[12] & g[6354];
assign g[14545] = b[12] & g[6354];
assign g[10451] = a[12] & g[6355];
assign g[14546] = b[12] & g[6355];
assign g[10452] = a[12] & g[6356];
assign g[14547] = b[12] & g[6356];
assign g[10453] = a[12] & g[6357];
assign g[14548] = b[12] & g[6357];
assign g[10454] = a[12] & g[6358];
assign g[14549] = b[12] & g[6358];
assign g[10455] = a[12] & g[6359];
assign g[14550] = b[12] & g[6359];
assign g[10456] = a[12] & g[6360];
assign g[14551] = b[12] & g[6360];
assign g[10457] = a[12] & g[6361];
assign g[14552] = b[12] & g[6361];
assign g[10458] = a[12] & g[6362];
assign g[14553] = b[12] & g[6362];
assign g[10459] = a[12] & g[6363];
assign g[14554] = b[12] & g[6363];
assign g[10460] = a[12] & g[6364];
assign g[14555] = b[12] & g[6364];
assign g[10461] = a[12] & g[6365];
assign g[14556] = b[12] & g[6365];
assign g[10462] = a[12] & g[6366];
assign g[14557] = b[12] & g[6366];
assign g[10463] = a[12] & g[6367];
assign g[14558] = b[12] & g[6367];
assign g[10464] = a[12] & g[6368];
assign g[14559] = b[12] & g[6368];
assign g[10465] = a[12] & g[6369];
assign g[14560] = b[12] & g[6369];
assign g[10466] = a[12] & g[6370];
assign g[14561] = b[12] & g[6370];
assign g[10467] = a[12] & g[6371];
assign g[14562] = b[12] & g[6371];
assign g[10468] = a[12] & g[6372];
assign g[14563] = b[12] & g[6372];
assign g[10469] = a[12] & g[6373];
assign g[14564] = b[12] & g[6373];
assign g[10470] = a[12] & g[6374];
assign g[14565] = b[12] & g[6374];
assign g[10471] = a[12] & g[6375];
assign g[14566] = b[12] & g[6375];
assign g[10472] = a[12] & g[6376];
assign g[14567] = b[12] & g[6376];
assign g[10473] = a[12] & g[6377];
assign g[14568] = b[12] & g[6377];
assign g[10474] = a[12] & g[6378];
assign g[14569] = b[12] & g[6378];
assign g[10475] = a[12] & g[6379];
assign g[14570] = b[12] & g[6379];
assign g[10476] = a[12] & g[6380];
assign g[14571] = b[12] & g[6380];
assign g[10477] = a[12] & g[6381];
assign g[14572] = b[12] & g[6381];
assign g[10478] = a[12] & g[6382];
assign g[14573] = b[12] & g[6382];
assign g[10479] = a[12] & g[6383];
assign g[14574] = b[12] & g[6383];
assign g[10480] = a[12] & g[6384];
assign g[14575] = b[12] & g[6384];
assign g[10481] = a[12] & g[6385];
assign g[14576] = b[12] & g[6385];
assign g[10482] = a[12] & g[6386];
assign g[14577] = b[12] & g[6386];
assign g[10483] = a[12] & g[6387];
assign g[14578] = b[12] & g[6387];
assign g[10484] = a[12] & g[6388];
assign g[14579] = b[12] & g[6388];
assign g[10485] = a[12] & g[6389];
assign g[14580] = b[12] & g[6389];
assign g[10486] = a[12] & g[6390];
assign g[14581] = b[12] & g[6390];
assign g[10487] = a[12] & g[6391];
assign g[14582] = b[12] & g[6391];
assign g[10488] = a[12] & g[6392];
assign g[14583] = b[12] & g[6392];
assign g[10489] = a[12] & g[6393];
assign g[14584] = b[12] & g[6393];
assign g[10490] = a[12] & g[6394];
assign g[14585] = b[12] & g[6394];
assign g[10491] = a[12] & g[6395];
assign g[14586] = b[12] & g[6395];
assign g[10492] = a[12] & g[6396];
assign g[14587] = b[12] & g[6396];
assign g[10493] = a[12] & g[6397];
assign g[14588] = b[12] & g[6397];
assign g[10494] = a[12] & g[6398];
assign g[14589] = b[12] & g[6398];
assign g[10495] = a[12] & g[6399];
assign g[14590] = b[12] & g[6399];
assign g[10496] = a[12] & g[6400];
assign g[14591] = b[12] & g[6400];
assign g[10497] = a[12] & g[6401];
assign g[14592] = b[12] & g[6401];
assign g[10498] = a[12] & g[6402];
assign g[14593] = b[12] & g[6402];
assign g[10499] = a[12] & g[6403];
assign g[14594] = b[12] & g[6403];
assign g[10500] = a[12] & g[6404];
assign g[14595] = b[12] & g[6404];
assign g[10501] = a[12] & g[6405];
assign g[14596] = b[12] & g[6405];
assign g[10502] = a[12] & g[6406];
assign g[14597] = b[12] & g[6406];
assign g[10503] = a[12] & g[6407];
assign g[14598] = b[12] & g[6407];
assign g[10504] = a[12] & g[6408];
assign g[14599] = b[12] & g[6408];
assign g[10505] = a[12] & g[6409];
assign g[14600] = b[12] & g[6409];
assign g[10506] = a[12] & g[6410];
assign g[14601] = b[12] & g[6410];
assign g[10507] = a[12] & g[6411];
assign g[14602] = b[12] & g[6411];
assign g[10508] = a[12] & g[6412];
assign g[14603] = b[12] & g[6412];
assign g[10509] = a[12] & g[6413];
assign g[14604] = b[12] & g[6413];
assign g[10510] = a[12] & g[6414];
assign g[14605] = b[12] & g[6414];
assign g[10511] = a[12] & g[6415];
assign g[14606] = b[12] & g[6415];
assign g[10512] = a[12] & g[6416];
assign g[14607] = b[12] & g[6416];
assign g[10513] = a[12] & g[6417];
assign g[14608] = b[12] & g[6417];
assign g[10514] = a[12] & g[6418];
assign g[14609] = b[12] & g[6418];
assign g[10515] = a[12] & g[6419];
assign g[14610] = b[12] & g[6419];
assign g[10516] = a[12] & g[6420];
assign g[14611] = b[12] & g[6420];
assign g[10517] = a[12] & g[6421];
assign g[14612] = b[12] & g[6421];
assign g[10518] = a[12] & g[6422];
assign g[14613] = b[12] & g[6422];
assign g[10519] = a[12] & g[6423];
assign g[14614] = b[12] & g[6423];
assign g[10520] = a[12] & g[6424];
assign g[14615] = b[12] & g[6424];
assign g[10521] = a[12] & g[6425];
assign g[14616] = b[12] & g[6425];
assign g[10522] = a[12] & g[6426];
assign g[14617] = b[12] & g[6426];
assign g[10523] = a[12] & g[6427];
assign g[14618] = b[12] & g[6427];
assign g[10524] = a[12] & g[6428];
assign g[14619] = b[12] & g[6428];
assign g[10525] = a[12] & g[6429];
assign g[14620] = b[12] & g[6429];
assign g[10526] = a[12] & g[6430];
assign g[14621] = b[12] & g[6430];
assign g[10527] = a[12] & g[6431];
assign g[14622] = b[12] & g[6431];
assign g[10528] = a[12] & g[6432];
assign g[14623] = b[12] & g[6432];
assign g[10529] = a[12] & g[6433];
assign g[14624] = b[12] & g[6433];
assign g[10530] = a[12] & g[6434];
assign g[14625] = b[12] & g[6434];
assign g[10531] = a[12] & g[6435];
assign g[14626] = b[12] & g[6435];
assign g[10532] = a[12] & g[6436];
assign g[14627] = b[12] & g[6436];
assign g[10533] = a[12] & g[6437];
assign g[14628] = b[12] & g[6437];
assign g[10534] = a[12] & g[6438];
assign g[14629] = b[12] & g[6438];
assign g[10535] = a[12] & g[6439];
assign g[14630] = b[12] & g[6439];
assign g[10536] = a[12] & g[6440];
assign g[14631] = b[12] & g[6440];
assign g[10537] = a[12] & g[6441];
assign g[14632] = b[12] & g[6441];
assign g[10538] = a[12] & g[6442];
assign g[14633] = b[12] & g[6442];
assign g[10539] = a[12] & g[6443];
assign g[14634] = b[12] & g[6443];
assign g[10540] = a[12] & g[6444];
assign g[14635] = b[12] & g[6444];
assign g[10541] = a[12] & g[6445];
assign g[14636] = b[12] & g[6445];
assign g[10542] = a[12] & g[6446];
assign g[14637] = b[12] & g[6446];
assign g[10543] = a[12] & g[6447];
assign g[14638] = b[12] & g[6447];
assign g[10544] = a[12] & g[6448];
assign g[14639] = b[12] & g[6448];
assign g[10545] = a[12] & g[6449];
assign g[14640] = b[12] & g[6449];
assign g[10546] = a[12] & g[6450];
assign g[14641] = b[12] & g[6450];
assign g[10547] = a[12] & g[6451];
assign g[14642] = b[12] & g[6451];
assign g[10548] = a[12] & g[6452];
assign g[14643] = b[12] & g[6452];
assign g[10549] = a[12] & g[6453];
assign g[14644] = b[12] & g[6453];
assign g[10550] = a[12] & g[6454];
assign g[14645] = b[12] & g[6454];
assign g[10551] = a[12] & g[6455];
assign g[14646] = b[12] & g[6455];
assign g[10552] = a[12] & g[6456];
assign g[14647] = b[12] & g[6456];
assign g[10553] = a[12] & g[6457];
assign g[14648] = b[12] & g[6457];
assign g[10554] = a[12] & g[6458];
assign g[14649] = b[12] & g[6458];
assign g[10555] = a[12] & g[6459];
assign g[14650] = b[12] & g[6459];
assign g[10556] = a[12] & g[6460];
assign g[14651] = b[12] & g[6460];
assign g[10557] = a[12] & g[6461];
assign g[14652] = b[12] & g[6461];
assign g[10558] = a[12] & g[6462];
assign g[14653] = b[12] & g[6462];
assign g[10559] = a[12] & g[6463];
assign g[14654] = b[12] & g[6463];
assign g[10560] = a[12] & g[6464];
assign g[14655] = b[12] & g[6464];
assign g[10561] = a[12] & g[6465];
assign g[14656] = b[12] & g[6465];
assign g[10562] = a[12] & g[6466];
assign g[14657] = b[12] & g[6466];
assign g[10563] = a[12] & g[6467];
assign g[14658] = b[12] & g[6467];
assign g[10564] = a[12] & g[6468];
assign g[14659] = b[12] & g[6468];
assign g[10565] = a[12] & g[6469];
assign g[14660] = b[12] & g[6469];
assign g[10566] = a[12] & g[6470];
assign g[14661] = b[12] & g[6470];
assign g[10567] = a[12] & g[6471];
assign g[14662] = b[12] & g[6471];
assign g[10568] = a[12] & g[6472];
assign g[14663] = b[12] & g[6472];
assign g[10569] = a[12] & g[6473];
assign g[14664] = b[12] & g[6473];
assign g[10570] = a[12] & g[6474];
assign g[14665] = b[12] & g[6474];
assign g[10571] = a[12] & g[6475];
assign g[14666] = b[12] & g[6475];
assign g[10572] = a[12] & g[6476];
assign g[14667] = b[12] & g[6476];
assign g[10573] = a[12] & g[6477];
assign g[14668] = b[12] & g[6477];
assign g[10574] = a[12] & g[6478];
assign g[14669] = b[12] & g[6478];
assign g[10575] = a[12] & g[6479];
assign g[14670] = b[12] & g[6479];
assign g[10576] = a[12] & g[6480];
assign g[14671] = b[12] & g[6480];
assign g[10577] = a[12] & g[6481];
assign g[14672] = b[12] & g[6481];
assign g[10578] = a[12] & g[6482];
assign g[14673] = b[12] & g[6482];
assign g[10579] = a[12] & g[6483];
assign g[14674] = b[12] & g[6483];
assign g[10580] = a[12] & g[6484];
assign g[14675] = b[12] & g[6484];
assign g[10581] = a[12] & g[6485];
assign g[14676] = b[12] & g[6485];
assign g[10582] = a[12] & g[6486];
assign g[14677] = b[12] & g[6486];
assign g[10583] = a[12] & g[6487];
assign g[14678] = b[12] & g[6487];
assign g[10584] = a[12] & g[6488];
assign g[14679] = b[12] & g[6488];
assign g[10585] = a[12] & g[6489];
assign g[14680] = b[12] & g[6489];
assign g[10586] = a[12] & g[6490];
assign g[14681] = b[12] & g[6490];
assign g[10587] = a[12] & g[6491];
assign g[14682] = b[12] & g[6491];
assign g[10588] = a[12] & g[6492];
assign g[14683] = b[12] & g[6492];
assign g[10589] = a[12] & g[6493];
assign g[14684] = b[12] & g[6493];
assign g[10590] = a[12] & g[6494];
assign g[14685] = b[12] & g[6494];
assign g[10591] = a[12] & g[6495];
assign g[14686] = b[12] & g[6495];
assign g[10592] = a[12] & g[6496];
assign g[14687] = b[12] & g[6496];
assign g[10593] = a[12] & g[6497];
assign g[14688] = b[12] & g[6497];
assign g[10594] = a[12] & g[6498];
assign g[14689] = b[12] & g[6498];
assign g[10595] = a[12] & g[6499];
assign g[14690] = b[12] & g[6499];
assign g[10596] = a[12] & g[6500];
assign g[14691] = b[12] & g[6500];
assign g[10597] = a[12] & g[6501];
assign g[14692] = b[12] & g[6501];
assign g[10598] = a[12] & g[6502];
assign g[14693] = b[12] & g[6502];
assign g[10599] = a[12] & g[6503];
assign g[14694] = b[12] & g[6503];
assign g[10600] = a[12] & g[6504];
assign g[14695] = b[12] & g[6504];
assign g[10601] = a[12] & g[6505];
assign g[14696] = b[12] & g[6505];
assign g[10602] = a[12] & g[6506];
assign g[14697] = b[12] & g[6506];
assign g[10603] = a[12] & g[6507];
assign g[14698] = b[12] & g[6507];
assign g[10604] = a[12] & g[6508];
assign g[14699] = b[12] & g[6508];
assign g[10605] = a[12] & g[6509];
assign g[14700] = b[12] & g[6509];
assign g[10606] = a[12] & g[6510];
assign g[14701] = b[12] & g[6510];
assign g[10607] = a[12] & g[6511];
assign g[14702] = b[12] & g[6511];
assign g[10608] = a[12] & g[6512];
assign g[14703] = b[12] & g[6512];
assign g[10609] = a[12] & g[6513];
assign g[14704] = b[12] & g[6513];
assign g[10610] = a[12] & g[6514];
assign g[14705] = b[12] & g[6514];
assign g[10611] = a[12] & g[6515];
assign g[14706] = b[12] & g[6515];
assign g[10612] = a[12] & g[6516];
assign g[14707] = b[12] & g[6516];
assign g[10613] = a[12] & g[6517];
assign g[14708] = b[12] & g[6517];
assign g[10614] = a[12] & g[6518];
assign g[14709] = b[12] & g[6518];
assign g[10615] = a[12] & g[6519];
assign g[14710] = b[12] & g[6519];
assign g[10616] = a[12] & g[6520];
assign g[14711] = b[12] & g[6520];
assign g[10617] = a[12] & g[6521];
assign g[14712] = b[12] & g[6521];
assign g[10618] = a[12] & g[6522];
assign g[14713] = b[12] & g[6522];
assign g[10619] = a[12] & g[6523];
assign g[14714] = b[12] & g[6523];
assign g[10620] = a[12] & g[6524];
assign g[14715] = b[12] & g[6524];
assign g[10621] = a[12] & g[6525];
assign g[14716] = b[12] & g[6525];
assign g[10622] = a[12] & g[6526];
assign g[14717] = b[12] & g[6526];
assign g[10623] = a[12] & g[6527];
assign g[14718] = b[12] & g[6527];
assign g[10624] = a[12] & g[6528];
assign g[14719] = b[12] & g[6528];
assign g[10625] = a[12] & g[6529];
assign g[14720] = b[12] & g[6529];
assign g[10626] = a[12] & g[6530];
assign g[14721] = b[12] & g[6530];
assign g[10627] = a[12] & g[6531];
assign g[14722] = b[12] & g[6531];
assign g[10628] = a[12] & g[6532];
assign g[14723] = b[12] & g[6532];
assign g[10629] = a[12] & g[6533];
assign g[14724] = b[12] & g[6533];
assign g[10630] = a[12] & g[6534];
assign g[14725] = b[12] & g[6534];
assign g[10631] = a[12] & g[6535];
assign g[14726] = b[12] & g[6535];
assign g[10632] = a[12] & g[6536];
assign g[14727] = b[12] & g[6536];
assign g[10633] = a[12] & g[6537];
assign g[14728] = b[12] & g[6537];
assign g[10634] = a[12] & g[6538];
assign g[14729] = b[12] & g[6538];
assign g[10635] = a[12] & g[6539];
assign g[14730] = b[12] & g[6539];
assign g[10636] = a[12] & g[6540];
assign g[14731] = b[12] & g[6540];
assign g[10637] = a[12] & g[6541];
assign g[14732] = b[12] & g[6541];
assign g[10638] = a[12] & g[6542];
assign g[14733] = b[12] & g[6542];
assign g[10639] = a[12] & g[6543];
assign g[14734] = b[12] & g[6543];
assign g[10640] = a[12] & g[6544];
assign g[14735] = b[12] & g[6544];
assign g[10641] = a[12] & g[6545];
assign g[14736] = b[12] & g[6545];
assign g[10642] = a[12] & g[6546];
assign g[14737] = b[12] & g[6546];
assign g[10643] = a[12] & g[6547];
assign g[14738] = b[12] & g[6547];
assign g[10644] = a[12] & g[6548];
assign g[14739] = b[12] & g[6548];
assign g[10645] = a[12] & g[6549];
assign g[14740] = b[12] & g[6549];
assign g[10646] = a[12] & g[6550];
assign g[14741] = b[12] & g[6550];
assign g[10647] = a[12] & g[6551];
assign g[14742] = b[12] & g[6551];
assign g[10648] = a[12] & g[6552];
assign g[14743] = b[12] & g[6552];
assign g[10649] = a[12] & g[6553];
assign g[14744] = b[12] & g[6553];
assign g[10650] = a[12] & g[6554];
assign g[14745] = b[12] & g[6554];
assign g[10651] = a[12] & g[6555];
assign g[14746] = b[12] & g[6555];
assign g[10652] = a[12] & g[6556];
assign g[14747] = b[12] & g[6556];
assign g[10653] = a[12] & g[6557];
assign g[14748] = b[12] & g[6557];
assign g[10654] = a[12] & g[6558];
assign g[14749] = b[12] & g[6558];
assign g[10655] = a[12] & g[6559];
assign g[14750] = b[12] & g[6559];
assign g[10656] = a[12] & g[6560];
assign g[14751] = b[12] & g[6560];
assign g[10657] = a[12] & g[6561];
assign g[14752] = b[12] & g[6561];
assign g[10658] = a[12] & g[6562];
assign g[14753] = b[12] & g[6562];
assign g[10659] = a[12] & g[6563];
assign g[14754] = b[12] & g[6563];
assign g[10660] = a[12] & g[6564];
assign g[14755] = b[12] & g[6564];
assign g[10661] = a[12] & g[6565];
assign g[14756] = b[12] & g[6565];
assign g[10662] = a[12] & g[6566];
assign g[14757] = b[12] & g[6566];
assign g[10663] = a[12] & g[6567];
assign g[14758] = b[12] & g[6567];
assign g[10664] = a[12] & g[6568];
assign g[14759] = b[12] & g[6568];
assign g[10665] = a[12] & g[6569];
assign g[14760] = b[12] & g[6569];
assign g[10666] = a[12] & g[6570];
assign g[14761] = b[12] & g[6570];
assign g[10667] = a[12] & g[6571];
assign g[14762] = b[12] & g[6571];
assign g[10668] = a[12] & g[6572];
assign g[14763] = b[12] & g[6572];
assign g[10669] = a[12] & g[6573];
assign g[14764] = b[12] & g[6573];
assign g[10670] = a[12] & g[6574];
assign g[14765] = b[12] & g[6574];
assign g[10671] = a[12] & g[6575];
assign g[14766] = b[12] & g[6575];
assign g[10672] = a[12] & g[6576];
assign g[14767] = b[12] & g[6576];
assign g[10673] = a[12] & g[6577];
assign g[14768] = b[12] & g[6577];
assign g[10674] = a[12] & g[6578];
assign g[14769] = b[12] & g[6578];
assign g[10675] = a[12] & g[6579];
assign g[14770] = b[12] & g[6579];
assign g[10676] = a[12] & g[6580];
assign g[14771] = b[12] & g[6580];
assign g[10677] = a[12] & g[6581];
assign g[14772] = b[12] & g[6581];
assign g[10678] = a[12] & g[6582];
assign g[14773] = b[12] & g[6582];
assign g[10679] = a[12] & g[6583];
assign g[14774] = b[12] & g[6583];
assign g[10680] = a[12] & g[6584];
assign g[14775] = b[12] & g[6584];
assign g[10681] = a[12] & g[6585];
assign g[14776] = b[12] & g[6585];
assign g[10682] = a[12] & g[6586];
assign g[14777] = b[12] & g[6586];
assign g[10683] = a[12] & g[6587];
assign g[14778] = b[12] & g[6587];
assign g[10684] = a[12] & g[6588];
assign g[14779] = b[12] & g[6588];
assign g[10685] = a[12] & g[6589];
assign g[14780] = b[12] & g[6589];
assign g[10686] = a[12] & g[6590];
assign g[14781] = b[12] & g[6590];
assign g[10687] = a[12] & g[6591];
assign g[14782] = b[12] & g[6591];
assign g[10688] = a[12] & g[6592];
assign g[14783] = b[12] & g[6592];
assign g[10689] = a[12] & g[6593];
assign g[14784] = b[12] & g[6593];
assign g[10690] = a[12] & g[6594];
assign g[14785] = b[12] & g[6594];
assign g[10691] = a[12] & g[6595];
assign g[14786] = b[12] & g[6595];
assign g[10692] = a[12] & g[6596];
assign g[14787] = b[12] & g[6596];
assign g[10693] = a[12] & g[6597];
assign g[14788] = b[12] & g[6597];
assign g[10694] = a[12] & g[6598];
assign g[14789] = b[12] & g[6598];
assign g[10695] = a[12] & g[6599];
assign g[14790] = b[12] & g[6599];
assign g[10696] = a[12] & g[6600];
assign g[14791] = b[12] & g[6600];
assign g[10697] = a[12] & g[6601];
assign g[14792] = b[12] & g[6601];
assign g[10698] = a[12] & g[6602];
assign g[14793] = b[12] & g[6602];
assign g[10699] = a[12] & g[6603];
assign g[14794] = b[12] & g[6603];
assign g[10700] = a[12] & g[6604];
assign g[14795] = b[12] & g[6604];
assign g[10701] = a[12] & g[6605];
assign g[14796] = b[12] & g[6605];
assign g[10702] = a[12] & g[6606];
assign g[14797] = b[12] & g[6606];
assign g[10703] = a[12] & g[6607];
assign g[14798] = b[12] & g[6607];
assign g[10704] = a[12] & g[6608];
assign g[14799] = b[12] & g[6608];
assign g[10705] = a[12] & g[6609];
assign g[14800] = b[12] & g[6609];
assign g[10706] = a[12] & g[6610];
assign g[14801] = b[12] & g[6610];
assign g[10707] = a[12] & g[6611];
assign g[14802] = b[12] & g[6611];
assign g[10708] = a[12] & g[6612];
assign g[14803] = b[12] & g[6612];
assign g[10709] = a[12] & g[6613];
assign g[14804] = b[12] & g[6613];
assign g[10710] = a[12] & g[6614];
assign g[14805] = b[12] & g[6614];
assign g[10711] = a[12] & g[6615];
assign g[14806] = b[12] & g[6615];
assign g[10712] = a[12] & g[6616];
assign g[14807] = b[12] & g[6616];
assign g[10713] = a[12] & g[6617];
assign g[14808] = b[12] & g[6617];
assign g[10714] = a[12] & g[6618];
assign g[14809] = b[12] & g[6618];
assign g[10715] = a[12] & g[6619];
assign g[14810] = b[12] & g[6619];
assign g[10716] = a[12] & g[6620];
assign g[14811] = b[12] & g[6620];
assign g[10717] = a[12] & g[6621];
assign g[14812] = b[12] & g[6621];
assign g[10718] = a[12] & g[6622];
assign g[14813] = b[12] & g[6622];
assign g[10719] = a[12] & g[6623];
assign g[14814] = b[12] & g[6623];
assign g[10720] = a[12] & g[6624];
assign g[14815] = b[12] & g[6624];
assign g[10721] = a[12] & g[6625];
assign g[14816] = b[12] & g[6625];
assign g[10722] = a[12] & g[6626];
assign g[14817] = b[12] & g[6626];
assign g[10723] = a[12] & g[6627];
assign g[14818] = b[12] & g[6627];
assign g[10724] = a[12] & g[6628];
assign g[14819] = b[12] & g[6628];
assign g[10725] = a[12] & g[6629];
assign g[14820] = b[12] & g[6629];
assign g[10726] = a[12] & g[6630];
assign g[14821] = b[12] & g[6630];
assign g[10727] = a[12] & g[6631];
assign g[14822] = b[12] & g[6631];
assign g[10728] = a[12] & g[6632];
assign g[14823] = b[12] & g[6632];
assign g[10729] = a[12] & g[6633];
assign g[14824] = b[12] & g[6633];
assign g[10730] = a[12] & g[6634];
assign g[14825] = b[12] & g[6634];
assign g[10731] = a[12] & g[6635];
assign g[14826] = b[12] & g[6635];
assign g[10732] = a[12] & g[6636];
assign g[14827] = b[12] & g[6636];
assign g[10733] = a[12] & g[6637];
assign g[14828] = b[12] & g[6637];
assign g[10734] = a[12] & g[6638];
assign g[14829] = b[12] & g[6638];
assign g[10735] = a[12] & g[6639];
assign g[14830] = b[12] & g[6639];
assign g[10736] = a[12] & g[6640];
assign g[14831] = b[12] & g[6640];
assign g[10737] = a[12] & g[6641];
assign g[14832] = b[12] & g[6641];
assign g[10738] = a[12] & g[6642];
assign g[14833] = b[12] & g[6642];
assign g[10739] = a[12] & g[6643];
assign g[14834] = b[12] & g[6643];
assign g[10740] = a[12] & g[6644];
assign g[14835] = b[12] & g[6644];
assign g[10741] = a[12] & g[6645];
assign g[14836] = b[12] & g[6645];
assign g[10742] = a[12] & g[6646];
assign g[14837] = b[12] & g[6646];
assign g[10743] = a[12] & g[6647];
assign g[14838] = b[12] & g[6647];
assign g[10744] = a[12] & g[6648];
assign g[14839] = b[12] & g[6648];
assign g[10745] = a[12] & g[6649];
assign g[14840] = b[12] & g[6649];
assign g[10746] = a[12] & g[6650];
assign g[14841] = b[12] & g[6650];
assign g[10747] = a[12] & g[6651];
assign g[14842] = b[12] & g[6651];
assign g[10748] = a[12] & g[6652];
assign g[14843] = b[12] & g[6652];
assign g[10749] = a[12] & g[6653];
assign g[14844] = b[12] & g[6653];
assign g[10750] = a[12] & g[6654];
assign g[14845] = b[12] & g[6654];
assign g[10751] = a[12] & g[6655];
assign g[14846] = b[12] & g[6655];
assign g[10752] = a[12] & g[6656];
assign g[14847] = b[12] & g[6656];
assign g[10753] = a[12] & g[6657];
assign g[14848] = b[12] & g[6657];
assign g[10754] = a[12] & g[6658];
assign g[14849] = b[12] & g[6658];
assign g[10755] = a[12] & g[6659];
assign g[14850] = b[12] & g[6659];
assign g[10756] = a[12] & g[6660];
assign g[14851] = b[12] & g[6660];
assign g[10757] = a[12] & g[6661];
assign g[14852] = b[12] & g[6661];
assign g[10758] = a[12] & g[6662];
assign g[14853] = b[12] & g[6662];
assign g[10759] = a[12] & g[6663];
assign g[14854] = b[12] & g[6663];
assign g[10760] = a[12] & g[6664];
assign g[14855] = b[12] & g[6664];
assign g[10761] = a[12] & g[6665];
assign g[14856] = b[12] & g[6665];
assign g[10762] = a[12] & g[6666];
assign g[14857] = b[12] & g[6666];
assign g[10763] = a[12] & g[6667];
assign g[14858] = b[12] & g[6667];
assign g[10764] = a[12] & g[6668];
assign g[14859] = b[12] & g[6668];
assign g[10765] = a[12] & g[6669];
assign g[14860] = b[12] & g[6669];
assign g[10766] = a[12] & g[6670];
assign g[14861] = b[12] & g[6670];
assign g[10767] = a[12] & g[6671];
assign g[14862] = b[12] & g[6671];
assign g[10768] = a[12] & g[6672];
assign g[14863] = b[12] & g[6672];
assign g[10769] = a[12] & g[6673];
assign g[14864] = b[12] & g[6673];
assign g[10770] = a[12] & g[6674];
assign g[14865] = b[12] & g[6674];
assign g[10771] = a[12] & g[6675];
assign g[14866] = b[12] & g[6675];
assign g[10772] = a[12] & g[6676];
assign g[14867] = b[12] & g[6676];
assign g[10773] = a[12] & g[6677];
assign g[14868] = b[12] & g[6677];
assign g[10774] = a[12] & g[6678];
assign g[14869] = b[12] & g[6678];
assign g[10775] = a[12] & g[6679];
assign g[14870] = b[12] & g[6679];
assign g[10776] = a[12] & g[6680];
assign g[14871] = b[12] & g[6680];
assign g[10777] = a[12] & g[6681];
assign g[14872] = b[12] & g[6681];
assign g[10778] = a[12] & g[6682];
assign g[14873] = b[12] & g[6682];
assign g[10779] = a[12] & g[6683];
assign g[14874] = b[12] & g[6683];
assign g[10780] = a[12] & g[6684];
assign g[14875] = b[12] & g[6684];
assign g[10781] = a[12] & g[6685];
assign g[14876] = b[12] & g[6685];
assign g[10782] = a[12] & g[6686];
assign g[14877] = b[12] & g[6686];
assign g[10783] = a[12] & g[6687];
assign g[14878] = b[12] & g[6687];
assign g[10784] = a[12] & g[6688];
assign g[14879] = b[12] & g[6688];
assign g[10785] = a[12] & g[6689];
assign g[14880] = b[12] & g[6689];
assign g[10786] = a[12] & g[6690];
assign g[14881] = b[12] & g[6690];
assign g[10787] = a[12] & g[6691];
assign g[14882] = b[12] & g[6691];
assign g[10788] = a[12] & g[6692];
assign g[14883] = b[12] & g[6692];
assign g[10789] = a[12] & g[6693];
assign g[14884] = b[12] & g[6693];
assign g[10790] = a[12] & g[6694];
assign g[14885] = b[12] & g[6694];
assign g[10791] = a[12] & g[6695];
assign g[14886] = b[12] & g[6695];
assign g[10792] = a[12] & g[6696];
assign g[14887] = b[12] & g[6696];
assign g[10793] = a[12] & g[6697];
assign g[14888] = b[12] & g[6697];
assign g[10794] = a[12] & g[6698];
assign g[14889] = b[12] & g[6698];
assign g[10795] = a[12] & g[6699];
assign g[14890] = b[12] & g[6699];
assign g[10796] = a[12] & g[6700];
assign g[14891] = b[12] & g[6700];
assign g[10797] = a[12] & g[6701];
assign g[14892] = b[12] & g[6701];
assign g[10798] = a[12] & g[6702];
assign g[14893] = b[12] & g[6702];
assign g[10799] = a[12] & g[6703];
assign g[14894] = b[12] & g[6703];
assign g[10800] = a[12] & g[6704];
assign g[14895] = b[12] & g[6704];
assign g[10801] = a[12] & g[6705];
assign g[14896] = b[12] & g[6705];
assign g[10802] = a[12] & g[6706];
assign g[14897] = b[12] & g[6706];
assign g[10803] = a[12] & g[6707];
assign g[14898] = b[12] & g[6707];
assign g[10804] = a[12] & g[6708];
assign g[14899] = b[12] & g[6708];
assign g[10805] = a[12] & g[6709];
assign g[14900] = b[12] & g[6709];
assign g[10806] = a[12] & g[6710];
assign g[14901] = b[12] & g[6710];
assign g[10807] = a[12] & g[6711];
assign g[14902] = b[12] & g[6711];
assign g[10808] = a[12] & g[6712];
assign g[14903] = b[12] & g[6712];
assign g[10809] = a[12] & g[6713];
assign g[14904] = b[12] & g[6713];
assign g[10810] = a[12] & g[6714];
assign g[14905] = b[12] & g[6714];
assign g[10811] = a[12] & g[6715];
assign g[14906] = b[12] & g[6715];
assign g[10812] = a[12] & g[6716];
assign g[14907] = b[12] & g[6716];
assign g[10813] = a[12] & g[6717];
assign g[14908] = b[12] & g[6717];
assign g[10814] = a[12] & g[6718];
assign g[14909] = b[12] & g[6718];
assign g[10815] = a[12] & g[6719];
assign g[14910] = b[12] & g[6719];
assign g[10816] = a[12] & g[6720];
assign g[14911] = b[12] & g[6720];
assign g[10817] = a[12] & g[6721];
assign g[14912] = b[12] & g[6721];
assign g[10818] = a[12] & g[6722];
assign g[14913] = b[12] & g[6722];
assign g[10819] = a[12] & g[6723];
assign g[14914] = b[12] & g[6723];
assign g[10820] = a[12] & g[6724];
assign g[14915] = b[12] & g[6724];
assign g[10821] = a[12] & g[6725];
assign g[14916] = b[12] & g[6725];
assign g[10822] = a[12] & g[6726];
assign g[14917] = b[12] & g[6726];
assign g[10823] = a[12] & g[6727];
assign g[14918] = b[12] & g[6727];
assign g[10824] = a[12] & g[6728];
assign g[14919] = b[12] & g[6728];
assign g[10825] = a[12] & g[6729];
assign g[14920] = b[12] & g[6729];
assign g[10826] = a[12] & g[6730];
assign g[14921] = b[12] & g[6730];
assign g[10827] = a[12] & g[6731];
assign g[14922] = b[12] & g[6731];
assign g[10828] = a[12] & g[6732];
assign g[14923] = b[12] & g[6732];
assign g[10829] = a[12] & g[6733];
assign g[14924] = b[12] & g[6733];
assign g[10830] = a[12] & g[6734];
assign g[14925] = b[12] & g[6734];
assign g[10831] = a[12] & g[6735];
assign g[14926] = b[12] & g[6735];
assign g[10832] = a[12] & g[6736];
assign g[14927] = b[12] & g[6736];
assign g[10833] = a[12] & g[6737];
assign g[14928] = b[12] & g[6737];
assign g[10834] = a[12] & g[6738];
assign g[14929] = b[12] & g[6738];
assign g[10835] = a[12] & g[6739];
assign g[14930] = b[12] & g[6739];
assign g[10836] = a[12] & g[6740];
assign g[14931] = b[12] & g[6740];
assign g[10837] = a[12] & g[6741];
assign g[14932] = b[12] & g[6741];
assign g[10838] = a[12] & g[6742];
assign g[14933] = b[12] & g[6742];
assign g[10839] = a[12] & g[6743];
assign g[14934] = b[12] & g[6743];
assign g[10840] = a[12] & g[6744];
assign g[14935] = b[12] & g[6744];
assign g[10841] = a[12] & g[6745];
assign g[14936] = b[12] & g[6745];
assign g[10842] = a[12] & g[6746];
assign g[14937] = b[12] & g[6746];
assign g[10843] = a[12] & g[6747];
assign g[14938] = b[12] & g[6747];
assign g[10844] = a[12] & g[6748];
assign g[14939] = b[12] & g[6748];
assign g[10845] = a[12] & g[6749];
assign g[14940] = b[12] & g[6749];
assign g[10846] = a[12] & g[6750];
assign g[14941] = b[12] & g[6750];
assign g[10847] = a[12] & g[6751];
assign g[14942] = b[12] & g[6751];
assign g[10848] = a[12] & g[6752];
assign g[14943] = b[12] & g[6752];
assign g[10849] = a[12] & g[6753];
assign g[14944] = b[12] & g[6753];
assign g[10850] = a[12] & g[6754];
assign g[14945] = b[12] & g[6754];
assign g[10851] = a[12] & g[6755];
assign g[14946] = b[12] & g[6755];
assign g[10852] = a[12] & g[6756];
assign g[14947] = b[12] & g[6756];
assign g[10853] = a[12] & g[6757];
assign g[14948] = b[12] & g[6757];
assign g[10854] = a[12] & g[6758];
assign g[14949] = b[12] & g[6758];
assign g[10855] = a[12] & g[6759];
assign g[14950] = b[12] & g[6759];
assign g[10856] = a[12] & g[6760];
assign g[14951] = b[12] & g[6760];
assign g[10857] = a[12] & g[6761];
assign g[14952] = b[12] & g[6761];
assign g[10858] = a[12] & g[6762];
assign g[14953] = b[12] & g[6762];
assign g[10859] = a[12] & g[6763];
assign g[14954] = b[12] & g[6763];
assign g[10860] = a[12] & g[6764];
assign g[14955] = b[12] & g[6764];
assign g[10861] = a[12] & g[6765];
assign g[14956] = b[12] & g[6765];
assign g[10862] = a[12] & g[6766];
assign g[14957] = b[12] & g[6766];
assign g[10863] = a[12] & g[6767];
assign g[14958] = b[12] & g[6767];
assign g[10864] = a[12] & g[6768];
assign g[14959] = b[12] & g[6768];
assign g[10865] = a[12] & g[6769];
assign g[14960] = b[12] & g[6769];
assign g[10866] = a[12] & g[6770];
assign g[14961] = b[12] & g[6770];
assign g[10867] = a[12] & g[6771];
assign g[14962] = b[12] & g[6771];
assign g[10868] = a[12] & g[6772];
assign g[14963] = b[12] & g[6772];
assign g[10869] = a[12] & g[6773];
assign g[14964] = b[12] & g[6773];
assign g[10870] = a[12] & g[6774];
assign g[14965] = b[12] & g[6774];
assign g[10871] = a[12] & g[6775];
assign g[14966] = b[12] & g[6775];
assign g[10872] = a[12] & g[6776];
assign g[14967] = b[12] & g[6776];
assign g[10873] = a[12] & g[6777];
assign g[14968] = b[12] & g[6777];
assign g[10874] = a[12] & g[6778];
assign g[14969] = b[12] & g[6778];
assign g[10875] = a[12] & g[6779];
assign g[14970] = b[12] & g[6779];
assign g[10876] = a[12] & g[6780];
assign g[14971] = b[12] & g[6780];
assign g[10877] = a[12] & g[6781];
assign g[14972] = b[12] & g[6781];
assign g[10878] = a[12] & g[6782];
assign g[14973] = b[12] & g[6782];
assign g[10879] = a[12] & g[6783];
assign g[14974] = b[12] & g[6783];
assign g[10880] = a[12] & g[6784];
assign g[14975] = b[12] & g[6784];
assign g[10881] = a[12] & g[6785];
assign g[14976] = b[12] & g[6785];
assign g[10882] = a[12] & g[6786];
assign g[14977] = b[12] & g[6786];
assign g[10883] = a[12] & g[6787];
assign g[14978] = b[12] & g[6787];
assign g[10884] = a[12] & g[6788];
assign g[14979] = b[12] & g[6788];
assign g[10885] = a[12] & g[6789];
assign g[14980] = b[12] & g[6789];
assign g[10886] = a[12] & g[6790];
assign g[14981] = b[12] & g[6790];
assign g[10887] = a[12] & g[6791];
assign g[14982] = b[12] & g[6791];
assign g[10888] = a[12] & g[6792];
assign g[14983] = b[12] & g[6792];
assign g[10889] = a[12] & g[6793];
assign g[14984] = b[12] & g[6793];
assign g[10890] = a[12] & g[6794];
assign g[14985] = b[12] & g[6794];
assign g[10891] = a[12] & g[6795];
assign g[14986] = b[12] & g[6795];
assign g[10892] = a[12] & g[6796];
assign g[14987] = b[12] & g[6796];
assign g[10893] = a[12] & g[6797];
assign g[14988] = b[12] & g[6797];
assign g[10894] = a[12] & g[6798];
assign g[14989] = b[12] & g[6798];
assign g[10895] = a[12] & g[6799];
assign g[14990] = b[12] & g[6799];
assign g[10896] = a[12] & g[6800];
assign g[14991] = b[12] & g[6800];
assign g[10897] = a[12] & g[6801];
assign g[14992] = b[12] & g[6801];
assign g[10898] = a[12] & g[6802];
assign g[14993] = b[12] & g[6802];
assign g[10899] = a[12] & g[6803];
assign g[14994] = b[12] & g[6803];
assign g[10900] = a[12] & g[6804];
assign g[14995] = b[12] & g[6804];
assign g[10901] = a[12] & g[6805];
assign g[14996] = b[12] & g[6805];
assign g[10902] = a[12] & g[6806];
assign g[14997] = b[12] & g[6806];
assign g[10903] = a[12] & g[6807];
assign g[14998] = b[12] & g[6807];
assign g[10904] = a[12] & g[6808];
assign g[14999] = b[12] & g[6808];
assign g[10905] = a[12] & g[6809];
assign g[15000] = b[12] & g[6809];
assign g[10906] = a[12] & g[6810];
assign g[15001] = b[12] & g[6810];
assign g[10907] = a[12] & g[6811];
assign g[15002] = b[12] & g[6811];
assign g[10908] = a[12] & g[6812];
assign g[15003] = b[12] & g[6812];
assign g[10909] = a[12] & g[6813];
assign g[15004] = b[12] & g[6813];
assign g[10910] = a[12] & g[6814];
assign g[15005] = b[12] & g[6814];
assign g[10911] = a[12] & g[6815];
assign g[15006] = b[12] & g[6815];
assign g[10912] = a[12] & g[6816];
assign g[15007] = b[12] & g[6816];
assign g[10913] = a[12] & g[6817];
assign g[15008] = b[12] & g[6817];
assign g[10914] = a[12] & g[6818];
assign g[15009] = b[12] & g[6818];
assign g[10915] = a[12] & g[6819];
assign g[15010] = b[12] & g[6819];
assign g[10916] = a[12] & g[6820];
assign g[15011] = b[12] & g[6820];
assign g[10917] = a[12] & g[6821];
assign g[15012] = b[12] & g[6821];
assign g[10918] = a[12] & g[6822];
assign g[15013] = b[12] & g[6822];
assign g[10919] = a[12] & g[6823];
assign g[15014] = b[12] & g[6823];
assign g[10920] = a[12] & g[6824];
assign g[15015] = b[12] & g[6824];
assign g[10921] = a[12] & g[6825];
assign g[15016] = b[12] & g[6825];
assign g[10922] = a[12] & g[6826];
assign g[15017] = b[12] & g[6826];
assign g[10923] = a[12] & g[6827];
assign g[15018] = b[12] & g[6827];
assign g[10924] = a[12] & g[6828];
assign g[15019] = b[12] & g[6828];
assign g[10925] = a[12] & g[6829];
assign g[15020] = b[12] & g[6829];
assign g[10926] = a[12] & g[6830];
assign g[15021] = b[12] & g[6830];
assign g[10927] = a[12] & g[6831];
assign g[15022] = b[12] & g[6831];
assign g[10928] = a[12] & g[6832];
assign g[15023] = b[12] & g[6832];
assign g[10929] = a[12] & g[6833];
assign g[15024] = b[12] & g[6833];
assign g[10930] = a[12] & g[6834];
assign g[15025] = b[12] & g[6834];
assign g[10931] = a[12] & g[6835];
assign g[15026] = b[12] & g[6835];
assign g[10932] = a[12] & g[6836];
assign g[15027] = b[12] & g[6836];
assign g[10933] = a[12] & g[6837];
assign g[15028] = b[12] & g[6837];
assign g[10934] = a[12] & g[6838];
assign g[15029] = b[12] & g[6838];
assign g[10935] = a[12] & g[6839];
assign g[15030] = b[12] & g[6839];
assign g[10936] = a[12] & g[6840];
assign g[15031] = b[12] & g[6840];
assign g[10937] = a[12] & g[6841];
assign g[15032] = b[12] & g[6841];
assign g[10938] = a[12] & g[6842];
assign g[15033] = b[12] & g[6842];
assign g[10939] = a[12] & g[6843];
assign g[15034] = b[12] & g[6843];
assign g[10940] = a[12] & g[6844];
assign g[15035] = b[12] & g[6844];
assign g[10941] = a[12] & g[6845];
assign g[15036] = b[12] & g[6845];
assign g[10942] = a[12] & g[6846];
assign g[15037] = b[12] & g[6846];
assign g[10943] = a[12] & g[6847];
assign g[15038] = b[12] & g[6847];
assign g[10944] = a[12] & g[6848];
assign g[15039] = b[12] & g[6848];
assign g[10945] = a[12] & g[6849];
assign g[15040] = b[12] & g[6849];
assign g[10946] = a[12] & g[6850];
assign g[15041] = b[12] & g[6850];
assign g[10947] = a[12] & g[6851];
assign g[15042] = b[12] & g[6851];
assign g[10948] = a[12] & g[6852];
assign g[15043] = b[12] & g[6852];
assign g[10949] = a[12] & g[6853];
assign g[15044] = b[12] & g[6853];
assign g[10950] = a[12] & g[6854];
assign g[15045] = b[12] & g[6854];
assign g[10951] = a[12] & g[6855];
assign g[15046] = b[12] & g[6855];
assign g[10952] = a[12] & g[6856];
assign g[15047] = b[12] & g[6856];
assign g[10953] = a[12] & g[6857];
assign g[15048] = b[12] & g[6857];
assign g[10954] = a[12] & g[6858];
assign g[15049] = b[12] & g[6858];
assign g[10955] = a[12] & g[6859];
assign g[15050] = b[12] & g[6859];
assign g[10956] = a[12] & g[6860];
assign g[15051] = b[12] & g[6860];
assign g[10957] = a[12] & g[6861];
assign g[15052] = b[12] & g[6861];
assign g[10958] = a[12] & g[6862];
assign g[15053] = b[12] & g[6862];
assign g[10959] = a[12] & g[6863];
assign g[15054] = b[12] & g[6863];
assign g[10960] = a[12] & g[6864];
assign g[15055] = b[12] & g[6864];
assign g[10961] = a[12] & g[6865];
assign g[15056] = b[12] & g[6865];
assign g[10962] = a[12] & g[6866];
assign g[15057] = b[12] & g[6866];
assign g[10963] = a[12] & g[6867];
assign g[15058] = b[12] & g[6867];
assign g[10964] = a[12] & g[6868];
assign g[15059] = b[12] & g[6868];
assign g[10965] = a[12] & g[6869];
assign g[15060] = b[12] & g[6869];
assign g[10966] = a[12] & g[6870];
assign g[15061] = b[12] & g[6870];
assign g[10967] = a[12] & g[6871];
assign g[15062] = b[12] & g[6871];
assign g[10968] = a[12] & g[6872];
assign g[15063] = b[12] & g[6872];
assign g[10969] = a[12] & g[6873];
assign g[15064] = b[12] & g[6873];
assign g[10970] = a[12] & g[6874];
assign g[15065] = b[12] & g[6874];
assign g[10971] = a[12] & g[6875];
assign g[15066] = b[12] & g[6875];
assign g[10972] = a[12] & g[6876];
assign g[15067] = b[12] & g[6876];
assign g[10973] = a[12] & g[6877];
assign g[15068] = b[12] & g[6877];
assign g[10974] = a[12] & g[6878];
assign g[15069] = b[12] & g[6878];
assign g[10975] = a[12] & g[6879];
assign g[15070] = b[12] & g[6879];
assign g[10976] = a[12] & g[6880];
assign g[15071] = b[12] & g[6880];
assign g[10977] = a[12] & g[6881];
assign g[15072] = b[12] & g[6881];
assign g[10978] = a[12] & g[6882];
assign g[15073] = b[12] & g[6882];
assign g[10979] = a[12] & g[6883];
assign g[15074] = b[12] & g[6883];
assign g[10980] = a[12] & g[6884];
assign g[15075] = b[12] & g[6884];
assign g[10981] = a[12] & g[6885];
assign g[15076] = b[12] & g[6885];
assign g[10982] = a[12] & g[6886];
assign g[15077] = b[12] & g[6886];
assign g[10983] = a[12] & g[6887];
assign g[15078] = b[12] & g[6887];
assign g[10984] = a[12] & g[6888];
assign g[15079] = b[12] & g[6888];
assign g[10985] = a[12] & g[6889];
assign g[15080] = b[12] & g[6889];
assign g[10986] = a[12] & g[6890];
assign g[15081] = b[12] & g[6890];
assign g[10987] = a[12] & g[6891];
assign g[15082] = b[12] & g[6891];
assign g[10988] = a[12] & g[6892];
assign g[15083] = b[12] & g[6892];
assign g[10989] = a[12] & g[6893];
assign g[15084] = b[12] & g[6893];
assign g[10990] = a[12] & g[6894];
assign g[15085] = b[12] & g[6894];
assign g[10991] = a[12] & g[6895];
assign g[15086] = b[12] & g[6895];
assign g[10992] = a[12] & g[6896];
assign g[15087] = b[12] & g[6896];
assign g[10993] = a[12] & g[6897];
assign g[15088] = b[12] & g[6897];
assign g[10994] = a[12] & g[6898];
assign g[15089] = b[12] & g[6898];
assign g[10995] = a[12] & g[6899];
assign g[15090] = b[12] & g[6899];
assign g[10996] = a[12] & g[6900];
assign g[15091] = b[12] & g[6900];
assign g[10997] = a[12] & g[6901];
assign g[15092] = b[12] & g[6901];
assign g[10998] = a[12] & g[6902];
assign g[15093] = b[12] & g[6902];
assign g[10999] = a[12] & g[6903];
assign g[15094] = b[12] & g[6903];
assign g[11000] = a[12] & g[6904];
assign g[15095] = b[12] & g[6904];
assign g[11001] = a[12] & g[6905];
assign g[15096] = b[12] & g[6905];
assign g[11002] = a[12] & g[6906];
assign g[15097] = b[12] & g[6906];
assign g[11003] = a[12] & g[6907];
assign g[15098] = b[12] & g[6907];
assign g[11004] = a[12] & g[6908];
assign g[15099] = b[12] & g[6908];
assign g[11005] = a[12] & g[6909];
assign g[15100] = b[12] & g[6909];
assign g[11006] = a[12] & g[6910];
assign g[15101] = b[12] & g[6910];
assign g[11007] = a[12] & g[6911];
assign g[15102] = b[12] & g[6911];
assign g[11008] = a[12] & g[6912];
assign g[15103] = b[12] & g[6912];
assign g[11009] = a[12] & g[6913];
assign g[15104] = b[12] & g[6913];
assign g[11010] = a[12] & g[6914];
assign g[15105] = b[12] & g[6914];
assign g[11011] = a[12] & g[6915];
assign g[15106] = b[12] & g[6915];
assign g[11012] = a[12] & g[6916];
assign g[15107] = b[12] & g[6916];
assign g[11013] = a[12] & g[6917];
assign g[15108] = b[12] & g[6917];
assign g[11014] = a[12] & g[6918];
assign g[15109] = b[12] & g[6918];
assign g[11015] = a[12] & g[6919];
assign g[15110] = b[12] & g[6919];
assign g[11016] = a[12] & g[6920];
assign g[15111] = b[12] & g[6920];
assign g[11017] = a[12] & g[6921];
assign g[15112] = b[12] & g[6921];
assign g[11018] = a[12] & g[6922];
assign g[15113] = b[12] & g[6922];
assign g[11019] = a[12] & g[6923];
assign g[15114] = b[12] & g[6923];
assign g[11020] = a[12] & g[6924];
assign g[15115] = b[12] & g[6924];
assign g[11021] = a[12] & g[6925];
assign g[15116] = b[12] & g[6925];
assign g[11022] = a[12] & g[6926];
assign g[15117] = b[12] & g[6926];
assign g[11023] = a[12] & g[6927];
assign g[15118] = b[12] & g[6927];
assign g[11024] = a[12] & g[6928];
assign g[15119] = b[12] & g[6928];
assign g[11025] = a[12] & g[6929];
assign g[15120] = b[12] & g[6929];
assign g[11026] = a[12] & g[6930];
assign g[15121] = b[12] & g[6930];
assign g[11027] = a[12] & g[6931];
assign g[15122] = b[12] & g[6931];
assign g[11028] = a[12] & g[6932];
assign g[15123] = b[12] & g[6932];
assign g[11029] = a[12] & g[6933];
assign g[15124] = b[12] & g[6933];
assign g[11030] = a[12] & g[6934];
assign g[15125] = b[12] & g[6934];
assign g[11031] = a[12] & g[6935];
assign g[15126] = b[12] & g[6935];
assign g[11032] = a[12] & g[6936];
assign g[15127] = b[12] & g[6936];
assign g[11033] = a[12] & g[6937];
assign g[15128] = b[12] & g[6937];
assign g[11034] = a[12] & g[6938];
assign g[15129] = b[12] & g[6938];
assign g[11035] = a[12] & g[6939];
assign g[15130] = b[12] & g[6939];
assign g[11036] = a[12] & g[6940];
assign g[15131] = b[12] & g[6940];
assign g[11037] = a[12] & g[6941];
assign g[15132] = b[12] & g[6941];
assign g[11038] = a[12] & g[6942];
assign g[15133] = b[12] & g[6942];
assign g[11039] = a[12] & g[6943];
assign g[15134] = b[12] & g[6943];
assign g[11040] = a[12] & g[6944];
assign g[15135] = b[12] & g[6944];
assign g[11041] = a[12] & g[6945];
assign g[15136] = b[12] & g[6945];
assign g[11042] = a[12] & g[6946];
assign g[15137] = b[12] & g[6946];
assign g[11043] = a[12] & g[6947];
assign g[15138] = b[12] & g[6947];
assign g[11044] = a[12] & g[6948];
assign g[15139] = b[12] & g[6948];
assign g[11045] = a[12] & g[6949];
assign g[15140] = b[12] & g[6949];
assign g[11046] = a[12] & g[6950];
assign g[15141] = b[12] & g[6950];
assign g[11047] = a[12] & g[6951];
assign g[15142] = b[12] & g[6951];
assign g[11048] = a[12] & g[6952];
assign g[15143] = b[12] & g[6952];
assign g[11049] = a[12] & g[6953];
assign g[15144] = b[12] & g[6953];
assign g[11050] = a[12] & g[6954];
assign g[15145] = b[12] & g[6954];
assign g[11051] = a[12] & g[6955];
assign g[15146] = b[12] & g[6955];
assign g[11052] = a[12] & g[6956];
assign g[15147] = b[12] & g[6956];
assign g[11053] = a[12] & g[6957];
assign g[15148] = b[12] & g[6957];
assign g[11054] = a[12] & g[6958];
assign g[15149] = b[12] & g[6958];
assign g[11055] = a[12] & g[6959];
assign g[15150] = b[12] & g[6959];
assign g[11056] = a[12] & g[6960];
assign g[15151] = b[12] & g[6960];
assign g[11057] = a[12] & g[6961];
assign g[15152] = b[12] & g[6961];
assign g[11058] = a[12] & g[6962];
assign g[15153] = b[12] & g[6962];
assign g[11059] = a[12] & g[6963];
assign g[15154] = b[12] & g[6963];
assign g[11060] = a[12] & g[6964];
assign g[15155] = b[12] & g[6964];
assign g[11061] = a[12] & g[6965];
assign g[15156] = b[12] & g[6965];
assign g[11062] = a[12] & g[6966];
assign g[15157] = b[12] & g[6966];
assign g[11063] = a[12] & g[6967];
assign g[15158] = b[12] & g[6967];
assign g[11064] = a[12] & g[6968];
assign g[15159] = b[12] & g[6968];
assign g[11065] = a[12] & g[6969];
assign g[15160] = b[12] & g[6969];
assign g[11066] = a[12] & g[6970];
assign g[15161] = b[12] & g[6970];
assign g[11067] = a[12] & g[6971];
assign g[15162] = b[12] & g[6971];
assign g[11068] = a[12] & g[6972];
assign g[15163] = b[12] & g[6972];
assign g[11069] = a[12] & g[6973];
assign g[15164] = b[12] & g[6973];
assign g[11070] = a[12] & g[6974];
assign g[15165] = b[12] & g[6974];
assign g[11071] = a[12] & g[6975];
assign g[15166] = b[12] & g[6975];
assign g[11072] = a[12] & g[6976];
assign g[15167] = b[12] & g[6976];
assign g[11073] = a[12] & g[6977];
assign g[15168] = b[12] & g[6977];
assign g[11074] = a[12] & g[6978];
assign g[15169] = b[12] & g[6978];
assign g[11075] = a[12] & g[6979];
assign g[15170] = b[12] & g[6979];
assign g[11076] = a[12] & g[6980];
assign g[15171] = b[12] & g[6980];
assign g[11077] = a[12] & g[6981];
assign g[15172] = b[12] & g[6981];
assign g[11078] = a[12] & g[6982];
assign g[15173] = b[12] & g[6982];
assign g[11079] = a[12] & g[6983];
assign g[15174] = b[12] & g[6983];
assign g[11080] = a[12] & g[6984];
assign g[15175] = b[12] & g[6984];
assign g[11081] = a[12] & g[6985];
assign g[15176] = b[12] & g[6985];
assign g[11082] = a[12] & g[6986];
assign g[15177] = b[12] & g[6986];
assign g[11083] = a[12] & g[6987];
assign g[15178] = b[12] & g[6987];
assign g[11084] = a[12] & g[6988];
assign g[15179] = b[12] & g[6988];
assign g[11085] = a[12] & g[6989];
assign g[15180] = b[12] & g[6989];
assign g[11086] = a[12] & g[6990];
assign g[15181] = b[12] & g[6990];
assign g[11087] = a[12] & g[6991];
assign g[15182] = b[12] & g[6991];
assign g[11088] = a[12] & g[6992];
assign g[15183] = b[12] & g[6992];
assign g[11089] = a[12] & g[6993];
assign g[15184] = b[12] & g[6993];
assign g[11090] = a[12] & g[6994];
assign g[15185] = b[12] & g[6994];
assign g[11091] = a[12] & g[6995];
assign g[15186] = b[12] & g[6995];
assign g[11092] = a[12] & g[6996];
assign g[15187] = b[12] & g[6996];
assign g[11093] = a[12] & g[6997];
assign g[15188] = b[12] & g[6997];
assign g[11094] = a[12] & g[6998];
assign g[15189] = b[12] & g[6998];
assign g[11095] = a[12] & g[6999];
assign g[15190] = b[12] & g[6999];
assign g[11096] = a[12] & g[7000];
assign g[15191] = b[12] & g[7000];
assign g[11097] = a[12] & g[7001];
assign g[15192] = b[12] & g[7001];
assign g[11098] = a[12] & g[7002];
assign g[15193] = b[12] & g[7002];
assign g[11099] = a[12] & g[7003];
assign g[15194] = b[12] & g[7003];
assign g[11100] = a[12] & g[7004];
assign g[15195] = b[12] & g[7004];
assign g[11101] = a[12] & g[7005];
assign g[15196] = b[12] & g[7005];
assign g[11102] = a[12] & g[7006];
assign g[15197] = b[12] & g[7006];
assign g[11103] = a[12] & g[7007];
assign g[15198] = b[12] & g[7007];
assign g[11104] = a[12] & g[7008];
assign g[15199] = b[12] & g[7008];
assign g[11105] = a[12] & g[7009];
assign g[15200] = b[12] & g[7009];
assign g[11106] = a[12] & g[7010];
assign g[15201] = b[12] & g[7010];
assign g[11107] = a[12] & g[7011];
assign g[15202] = b[12] & g[7011];
assign g[11108] = a[12] & g[7012];
assign g[15203] = b[12] & g[7012];
assign g[11109] = a[12] & g[7013];
assign g[15204] = b[12] & g[7013];
assign g[11110] = a[12] & g[7014];
assign g[15205] = b[12] & g[7014];
assign g[11111] = a[12] & g[7015];
assign g[15206] = b[12] & g[7015];
assign g[11112] = a[12] & g[7016];
assign g[15207] = b[12] & g[7016];
assign g[11113] = a[12] & g[7017];
assign g[15208] = b[12] & g[7017];
assign g[11114] = a[12] & g[7018];
assign g[15209] = b[12] & g[7018];
assign g[11115] = a[12] & g[7019];
assign g[15210] = b[12] & g[7019];
assign g[11116] = a[12] & g[7020];
assign g[15211] = b[12] & g[7020];
assign g[11117] = a[12] & g[7021];
assign g[15212] = b[12] & g[7021];
assign g[11118] = a[12] & g[7022];
assign g[15213] = b[12] & g[7022];
assign g[11119] = a[12] & g[7023];
assign g[15214] = b[12] & g[7023];
assign g[11120] = a[12] & g[7024];
assign g[15215] = b[12] & g[7024];
assign g[11121] = a[12] & g[7025];
assign g[15216] = b[12] & g[7025];
assign g[11122] = a[12] & g[7026];
assign g[15217] = b[12] & g[7026];
assign g[11123] = a[12] & g[7027];
assign g[15218] = b[12] & g[7027];
assign g[11124] = a[12] & g[7028];
assign g[15219] = b[12] & g[7028];
assign g[11125] = a[12] & g[7029];
assign g[15220] = b[12] & g[7029];
assign g[11126] = a[12] & g[7030];
assign g[15221] = b[12] & g[7030];
assign g[11127] = a[12] & g[7031];
assign g[15222] = b[12] & g[7031];
assign g[11128] = a[12] & g[7032];
assign g[15223] = b[12] & g[7032];
assign g[11129] = a[12] & g[7033];
assign g[15224] = b[12] & g[7033];
assign g[11130] = a[12] & g[7034];
assign g[15225] = b[12] & g[7034];
assign g[11131] = a[12] & g[7035];
assign g[15226] = b[12] & g[7035];
assign g[11132] = a[12] & g[7036];
assign g[15227] = b[12] & g[7036];
assign g[11133] = a[12] & g[7037];
assign g[15228] = b[12] & g[7037];
assign g[11134] = a[12] & g[7038];
assign g[15229] = b[12] & g[7038];
assign g[11135] = a[12] & g[7039];
assign g[15230] = b[12] & g[7039];
assign g[11136] = a[12] & g[7040];
assign g[15231] = b[12] & g[7040];
assign g[11137] = a[12] & g[7041];
assign g[15232] = b[12] & g[7041];
assign g[11138] = a[12] & g[7042];
assign g[15233] = b[12] & g[7042];
assign g[11139] = a[12] & g[7043];
assign g[15234] = b[12] & g[7043];
assign g[11140] = a[12] & g[7044];
assign g[15235] = b[12] & g[7044];
assign g[11141] = a[12] & g[7045];
assign g[15236] = b[12] & g[7045];
assign g[11142] = a[12] & g[7046];
assign g[15237] = b[12] & g[7046];
assign g[11143] = a[12] & g[7047];
assign g[15238] = b[12] & g[7047];
assign g[11144] = a[12] & g[7048];
assign g[15239] = b[12] & g[7048];
assign g[11145] = a[12] & g[7049];
assign g[15240] = b[12] & g[7049];
assign g[11146] = a[12] & g[7050];
assign g[15241] = b[12] & g[7050];
assign g[11147] = a[12] & g[7051];
assign g[15242] = b[12] & g[7051];
assign g[11148] = a[12] & g[7052];
assign g[15243] = b[12] & g[7052];
assign g[11149] = a[12] & g[7053];
assign g[15244] = b[12] & g[7053];
assign g[11150] = a[12] & g[7054];
assign g[15245] = b[12] & g[7054];
assign g[11151] = a[12] & g[7055];
assign g[15246] = b[12] & g[7055];
assign g[11152] = a[12] & g[7056];
assign g[15247] = b[12] & g[7056];
assign g[11153] = a[12] & g[7057];
assign g[15248] = b[12] & g[7057];
assign g[11154] = a[12] & g[7058];
assign g[15249] = b[12] & g[7058];
assign g[11155] = a[12] & g[7059];
assign g[15250] = b[12] & g[7059];
assign g[11156] = a[12] & g[7060];
assign g[15251] = b[12] & g[7060];
assign g[11157] = a[12] & g[7061];
assign g[15252] = b[12] & g[7061];
assign g[11158] = a[12] & g[7062];
assign g[15253] = b[12] & g[7062];
assign g[11159] = a[12] & g[7063];
assign g[15254] = b[12] & g[7063];
assign g[11160] = a[12] & g[7064];
assign g[15255] = b[12] & g[7064];
assign g[11161] = a[12] & g[7065];
assign g[15256] = b[12] & g[7065];
assign g[11162] = a[12] & g[7066];
assign g[15257] = b[12] & g[7066];
assign g[11163] = a[12] & g[7067];
assign g[15258] = b[12] & g[7067];
assign g[11164] = a[12] & g[7068];
assign g[15259] = b[12] & g[7068];
assign g[11165] = a[12] & g[7069];
assign g[15260] = b[12] & g[7069];
assign g[11166] = a[12] & g[7070];
assign g[15261] = b[12] & g[7070];
assign g[11167] = a[12] & g[7071];
assign g[15262] = b[12] & g[7071];
assign g[11168] = a[12] & g[7072];
assign g[15263] = b[12] & g[7072];
assign g[11169] = a[12] & g[7073];
assign g[15264] = b[12] & g[7073];
assign g[11170] = a[12] & g[7074];
assign g[15265] = b[12] & g[7074];
assign g[11171] = a[12] & g[7075];
assign g[15266] = b[12] & g[7075];
assign g[11172] = a[12] & g[7076];
assign g[15267] = b[12] & g[7076];
assign g[11173] = a[12] & g[7077];
assign g[15268] = b[12] & g[7077];
assign g[11174] = a[12] & g[7078];
assign g[15269] = b[12] & g[7078];
assign g[11175] = a[12] & g[7079];
assign g[15270] = b[12] & g[7079];
assign g[11176] = a[12] & g[7080];
assign g[15271] = b[12] & g[7080];
assign g[11177] = a[12] & g[7081];
assign g[15272] = b[12] & g[7081];
assign g[11178] = a[12] & g[7082];
assign g[15273] = b[12] & g[7082];
assign g[11179] = a[12] & g[7083];
assign g[15274] = b[12] & g[7083];
assign g[11180] = a[12] & g[7084];
assign g[15275] = b[12] & g[7084];
assign g[11181] = a[12] & g[7085];
assign g[15276] = b[12] & g[7085];
assign g[11182] = a[12] & g[7086];
assign g[15277] = b[12] & g[7086];
assign g[11183] = a[12] & g[7087];
assign g[15278] = b[12] & g[7087];
assign g[11184] = a[12] & g[7088];
assign g[15279] = b[12] & g[7088];
assign g[11185] = a[12] & g[7089];
assign g[15280] = b[12] & g[7089];
assign g[11186] = a[12] & g[7090];
assign g[15281] = b[12] & g[7090];
assign g[11187] = a[12] & g[7091];
assign g[15282] = b[12] & g[7091];
assign g[11188] = a[12] & g[7092];
assign g[15283] = b[12] & g[7092];
assign g[11189] = a[12] & g[7093];
assign g[15284] = b[12] & g[7093];
assign g[11190] = a[12] & g[7094];
assign g[15285] = b[12] & g[7094];
assign g[11191] = a[12] & g[7095];
assign g[15286] = b[12] & g[7095];
assign g[11192] = a[12] & g[7096];
assign g[15287] = b[12] & g[7096];
assign g[11193] = a[12] & g[7097];
assign g[15288] = b[12] & g[7097];
assign g[11194] = a[12] & g[7098];
assign g[15289] = b[12] & g[7098];
assign g[11195] = a[12] & g[7099];
assign g[15290] = b[12] & g[7099];
assign g[11196] = a[12] & g[7100];
assign g[15291] = b[12] & g[7100];
assign g[11197] = a[12] & g[7101];
assign g[15292] = b[12] & g[7101];
assign g[11198] = a[12] & g[7102];
assign g[15293] = b[12] & g[7102];
assign g[11199] = a[12] & g[7103];
assign g[15294] = b[12] & g[7103];
assign g[11200] = a[12] & g[7104];
assign g[15295] = b[12] & g[7104];
assign g[11201] = a[12] & g[7105];
assign g[15296] = b[12] & g[7105];
assign g[11202] = a[12] & g[7106];
assign g[15297] = b[12] & g[7106];
assign g[11203] = a[12] & g[7107];
assign g[15298] = b[12] & g[7107];
assign g[11204] = a[12] & g[7108];
assign g[15299] = b[12] & g[7108];
assign g[11205] = a[12] & g[7109];
assign g[15300] = b[12] & g[7109];
assign g[11206] = a[12] & g[7110];
assign g[15301] = b[12] & g[7110];
assign g[11207] = a[12] & g[7111];
assign g[15302] = b[12] & g[7111];
assign g[11208] = a[12] & g[7112];
assign g[15303] = b[12] & g[7112];
assign g[11209] = a[12] & g[7113];
assign g[15304] = b[12] & g[7113];
assign g[11210] = a[12] & g[7114];
assign g[15305] = b[12] & g[7114];
assign g[11211] = a[12] & g[7115];
assign g[15306] = b[12] & g[7115];
assign g[11212] = a[12] & g[7116];
assign g[15307] = b[12] & g[7116];
assign g[11213] = a[12] & g[7117];
assign g[15308] = b[12] & g[7117];
assign g[11214] = a[12] & g[7118];
assign g[15309] = b[12] & g[7118];
assign g[11215] = a[12] & g[7119];
assign g[15310] = b[12] & g[7119];
assign g[11216] = a[12] & g[7120];
assign g[15311] = b[12] & g[7120];
assign g[11217] = a[12] & g[7121];
assign g[15312] = b[12] & g[7121];
assign g[11218] = a[12] & g[7122];
assign g[15313] = b[12] & g[7122];
assign g[11219] = a[12] & g[7123];
assign g[15314] = b[12] & g[7123];
assign g[11220] = a[12] & g[7124];
assign g[15315] = b[12] & g[7124];
assign g[11221] = a[12] & g[7125];
assign g[15316] = b[12] & g[7125];
assign g[11222] = a[12] & g[7126];
assign g[15317] = b[12] & g[7126];
assign g[11223] = a[12] & g[7127];
assign g[15318] = b[12] & g[7127];
assign g[11224] = a[12] & g[7128];
assign g[15319] = b[12] & g[7128];
assign g[11225] = a[12] & g[7129];
assign g[15320] = b[12] & g[7129];
assign g[11226] = a[12] & g[7130];
assign g[15321] = b[12] & g[7130];
assign g[11227] = a[12] & g[7131];
assign g[15322] = b[12] & g[7131];
assign g[11228] = a[12] & g[7132];
assign g[15323] = b[12] & g[7132];
assign g[11229] = a[12] & g[7133];
assign g[15324] = b[12] & g[7133];
assign g[11230] = a[12] & g[7134];
assign g[15325] = b[12] & g[7134];
assign g[11231] = a[12] & g[7135];
assign g[15326] = b[12] & g[7135];
assign g[11232] = a[12] & g[7136];
assign g[15327] = b[12] & g[7136];
assign g[11233] = a[12] & g[7137];
assign g[15328] = b[12] & g[7137];
assign g[11234] = a[12] & g[7138];
assign g[15329] = b[12] & g[7138];
assign g[11235] = a[12] & g[7139];
assign g[15330] = b[12] & g[7139];
assign g[11236] = a[12] & g[7140];
assign g[15331] = b[12] & g[7140];
assign g[11237] = a[12] & g[7141];
assign g[15332] = b[12] & g[7141];
assign g[11238] = a[12] & g[7142];
assign g[15333] = b[12] & g[7142];
assign g[11239] = a[12] & g[7143];
assign g[15334] = b[12] & g[7143];
assign g[11240] = a[12] & g[7144];
assign g[15335] = b[12] & g[7144];
assign g[11241] = a[12] & g[7145];
assign g[15336] = b[12] & g[7145];
assign g[11242] = a[12] & g[7146];
assign g[15337] = b[12] & g[7146];
assign g[11243] = a[12] & g[7147];
assign g[15338] = b[12] & g[7147];
assign g[11244] = a[12] & g[7148];
assign g[15339] = b[12] & g[7148];
assign g[11245] = a[12] & g[7149];
assign g[15340] = b[12] & g[7149];
assign g[11246] = a[12] & g[7150];
assign g[15341] = b[12] & g[7150];
assign g[11247] = a[12] & g[7151];
assign g[15342] = b[12] & g[7151];
assign g[11248] = a[12] & g[7152];
assign g[15343] = b[12] & g[7152];
assign g[11249] = a[12] & g[7153];
assign g[15344] = b[12] & g[7153];
assign g[11250] = a[12] & g[7154];
assign g[15345] = b[12] & g[7154];
assign g[11251] = a[12] & g[7155];
assign g[15346] = b[12] & g[7155];
assign g[11252] = a[12] & g[7156];
assign g[15347] = b[12] & g[7156];
assign g[11253] = a[12] & g[7157];
assign g[15348] = b[12] & g[7157];
assign g[11254] = a[12] & g[7158];
assign g[15349] = b[12] & g[7158];
assign g[11255] = a[12] & g[7159];
assign g[15350] = b[12] & g[7159];
assign g[11256] = a[12] & g[7160];
assign g[15351] = b[12] & g[7160];
assign g[11257] = a[12] & g[7161];
assign g[15352] = b[12] & g[7161];
assign g[11258] = a[12] & g[7162];
assign g[15353] = b[12] & g[7162];
assign g[11259] = a[12] & g[7163];
assign g[15354] = b[12] & g[7163];
assign g[11260] = a[12] & g[7164];
assign g[15355] = b[12] & g[7164];
assign g[11261] = a[12] & g[7165];
assign g[15356] = b[12] & g[7165];
assign g[11262] = a[12] & g[7166];
assign g[15357] = b[12] & g[7166];
assign g[11263] = a[12] & g[7167];
assign g[15358] = b[12] & g[7167];
assign g[11264] = a[12] & g[7168];
assign g[15359] = b[12] & g[7168];
assign g[11265] = a[12] & g[7169];
assign g[15360] = b[12] & g[7169];
assign g[11266] = a[12] & g[7170];
assign g[15361] = b[12] & g[7170];
assign g[11267] = a[12] & g[7171];
assign g[15362] = b[12] & g[7171];
assign g[11268] = a[12] & g[7172];
assign g[15363] = b[12] & g[7172];
assign g[11269] = a[12] & g[7173];
assign g[15364] = b[12] & g[7173];
assign g[11270] = a[12] & g[7174];
assign g[15365] = b[12] & g[7174];
assign g[11271] = a[12] & g[7175];
assign g[15366] = b[12] & g[7175];
assign g[11272] = a[12] & g[7176];
assign g[15367] = b[12] & g[7176];
assign g[11273] = a[12] & g[7177];
assign g[15368] = b[12] & g[7177];
assign g[11274] = a[12] & g[7178];
assign g[15369] = b[12] & g[7178];
assign g[11275] = a[12] & g[7179];
assign g[15370] = b[12] & g[7179];
assign g[11276] = a[12] & g[7180];
assign g[15371] = b[12] & g[7180];
assign g[11277] = a[12] & g[7181];
assign g[15372] = b[12] & g[7181];
assign g[11278] = a[12] & g[7182];
assign g[15373] = b[12] & g[7182];
assign g[11279] = a[12] & g[7183];
assign g[15374] = b[12] & g[7183];
assign g[11280] = a[12] & g[7184];
assign g[15375] = b[12] & g[7184];
assign g[11281] = a[12] & g[7185];
assign g[15376] = b[12] & g[7185];
assign g[11282] = a[12] & g[7186];
assign g[15377] = b[12] & g[7186];
assign g[11283] = a[12] & g[7187];
assign g[15378] = b[12] & g[7187];
assign g[11284] = a[12] & g[7188];
assign g[15379] = b[12] & g[7188];
assign g[11285] = a[12] & g[7189];
assign g[15380] = b[12] & g[7189];
assign g[11286] = a[12] & g[7190];
assign g[15381] = b[12] & g[7190];
assign g[11287] = a[12] & g[7191];
assign g[15382] = b[12] & g[7191];
assign g[11288] = a[12] & g[7192];
assign g[15383] = b[12] & g[7192];
assign g[11289] = a[12] & g[7193];
assign g[15384] = b[12] & g[7193];
assign g[11290] = a[12] & g[7194];
assign g[15385] = b[12] & g[7194];
assign g[11291] = a[12] & g[7195];
assign g[15386] = b[12] & g[7195];
assign g[11292] = a[12] & g[7196];
assign g[15387] = b[12] & g[7196];
assign g[11293] = a[12] & g[7197];
assign g[15388] = b[12] & g[7197];
assign g[11294] = a[12] & g[7198];
assign g[15389] = b[12] & g[7198];
assign g[11295] = a[12] & g[7199];
assign g[15390] = b[12] & g[7199];
assign g[11296] = a[12] & g[7200];
assign g[15391] = b[12] & g[7200];
assign g[11297] = a[12] & g[7201];
assign g[15392] = b[12] & g[7201];
assign g[11298] = a[12] & g[7202];
assign g[15393] = b[12] & g[7202];
assign g[11299] = a[12] & g[7203];
assign g[15394] = b[12] & g[7203];
assign g[11300] = a[12] & g[7204];
assign g[15395] = b[12] & g[7204];
assign g[11301] = a[12] & g[7205];
assign g[15396] = b[12] & g[7205];
assign g[11302] = a[12] & g[7206];
assign g[15397] = b[12] & g[7206];
assign g[11303] = a[12] & g[7207];
assign g[15398] = b[12] & g[7207];
assign g[11304] = a[12] & g[7208];
assign g[15399] = b[12] & g[7208];
assign g[11305] = a[12] & g[7209];
assign g[15400] = b[12] & g[7209];
assign g[11306] = a[12] & g[7210];
assign g[15401] = b[12] & g[7210];
assign g[11307] = a[12] & g[7211];
assign g[15402] = b[12] & g[7211];
assign g[11308] = a[12] & g[7212];
assign g[15403] = b[12] & g[7212];
assign g[11309] = a[12] & g[7213];
assign g[15404] = b[12] & g[7213];
assign g[11310] = a[12] & g[7214];
assign g[15405] = b[12] & g[7214];
assign g[11311] = a[12] & g[7215];
assign g[15406] = b[12] & g[7215];
assign g[11312] = a[12] & g[7216];
assign g[15407] = b[12] & g[7216];
assign g[11313] = a[12] & g[7217];
assign g[15408] = b[12] & g[7217];
assign g[11314] = a[12] & g[7218];
assign g[15409] = b[12] & g[7218];
assign g[11315] = a[12] & g[7219];
assign g[15410] = b[12] & g[7219];
assign g[11316] = a[12] & g[7220];
assign g[15411] = b[12] & g[7220];
assign g[11317] = a[12] & g[7221];
assign g[15412] = b[12] & g[7221];
assign g[11318] = a[12] & g[7222];
assign g[15413] = b[12] & g[7222];
assign g[11319] = a[12] & g[7223];
assign g[15414] = b[12] & g[7223];
assign g[11320] = a[12] & g[7224];
assign g[15415] = b[12] & g[7224];
assign g[11321] = a[12] & g[7225];
assign g[15416] = b[12] & g[7225];
assign g[11322] = a[12] & g[7226];
assign g[15417] = b[12] & g[7226];
assign g[11323] = a[12] & g[7227];
assign g[15418] = b[12] & g[7227];
assign g[11324] = a[12] & g[7228];
assign g[15419] = b[12] & g[7228];
assign g[11325] = a[12] & g[7229];
assign g[15420] = b[12] & g[7229];
assign g[11326] = a[12] & g[7230];
assign g[15421] = b[12] & g[7230];
assign g[11327] = a[12] & g[7231];
assign g[15422] = b[12] & g[7231];
assign g[11328] = a[12] & g[7232];
assign g[15423] = b[12] & g[7232];
assign g[11329] = a[12] & g[7233];
assign g[15424] = b[12] & g[7233];
assign g[11330] = a[12] & g[7234];
assign g[15425] = b[12] & g[7234];
assign g[11331] = a[12] & g[7235];
assign g[15426] = b[12] & g[7235];
assign g[11332] = a[12] & g[7236];
assign g[15427] = b[12] & g[7236];
assign g[11333] = a[12] & g[7237];
assign g[15428] = b[12] & g[7237];
assign g[11334] = a[12] & g[7238];
assign g[15429] = b[12] & g[7238];
assign g[11335] = a[12] & g[7239];
assign g[15430] = b[12] & g[7239];
assign g[11336] = a[12] & g[7240];
assign g[15431] = b[12] & g[7240];
assign g[11337] = a[12] & g[7241];
assign g[15432] = b[12] & g[7241];
assign g[11338] = a[12] & g[7242];
assign g[15433] = b[12] & g[7242];
assign g[11339] = a[12] & g[7243];
assign g[15434] = b[12] & g[7243];
assign g[11340] = a[12] & g[7244];
assign g[15435] = b[12] & g[7244];
assign g[11341] = a[12] & g[7245];
assign g[15436] = b[12] & g[7245];
assign g[11342] = a[12] & g[7246];
assign g[15437] = b[12] & g[7246];
assign g[11343] = a[12] & g[7247];
assign g[15438] = b[12] & g[7247];
assign g[11344] = a[12] & g[7248];
assign g[15439] = b[12] & g[7248];
assign g[11345] = a[12] & g[7249];
assign g[15440] = b[12] & g[7249];
assign g[11346] = a[12] & g[7250];
assign g[15441] = b[12] & g[7250];
assign g[11347] = a[12] & g[7251];
assign g[15442] = b[12] & g[7251];
assign g[11348] = a[12] & g[7252];
assign g[15443] = b[12] & g[7252];
assign g[11349] = a[12] & g[7253];
assign g[15444] = b[12] & g[7253];
assign g[11350] = a[12] & g[7254];
assign g[15445] = b[12] & g[7254];
assign g[11351] = a[12] & g[7255];
assign g[15446] = b[12] & g[7255];
assign g[11352] = a[12] & g[7256];
assign g[15447] = b[12] & g[7256];
assign g[11353] = a[12] & g[7257];
assign g[15448] = b[12] & g[7257];
assign g[11354] = a[12] & g[7258];
assign g[15449] = b[12] & g[7258];
assign g[11355] = a[12] & g[7259];
assign g[15450] = b[12] & g[7259];
assign g[11356] = a[12] & g[7260];
assign g[15451] = b[12] & g[7260];
assign g[11357] = a[12] & g[7261];
assign g[15452] = b[12] & g[7261];
assign g[11358] = a[12] & g[7262];
assign g[15453] = b[12] & g[7262];
assign g[11359] = a[12] & g[7263];
assign g[15454] = b[12] & g[7263];
assign g[11360] = a[12] & g[7264];
assign g[15455] = b[12] & g[7264];
assign g[11361] = a[12] & g[7265];
assign g[15456] = b[12] & g[7265];
assign g[11362] = a[12] & g[7266];
assign g[15457] = b[12] & g[7266];
assign g[11363] = a[12] & g[7267];
assign g[15458] = b[12] & g[7267];
assign g[11364] = a[12] & g[7268];
assign g[15459] = b[12] & g[7268];
assign g[11365] = a[12] & g[7269];
assign g[15460] = b[12] & g[7269];
assign g[11366] = a[12] & g[7270];
assign g[15461] = b[12] & g[7270];
assign g[11367] = a[12] & g[7271];
assign g[15462] = b[12] & g[7271];
assign g[11368] = a[12] & g[7272];
assign g[15463] = b[12] & g[7272];
assign g[11369] = a[12] & g[7273];
assign g[15464] = b[12] & g[7273];
assign g[11370] = a[12] & g[7274];
assign g[15465] = b[12] & g[7274];
assign g[11371] = a[12] & g[7275];
assign g[15466] = b[12] & g[7275];
assign g[11372] = a[12] & g[7276];
assign g[15467] = b[12] & g[7276];
assign g[11373] = a[12] & g[7277];
assign g[15468] = b[12] & g[7277];
assign g[11374] = a[12] & g[7278];
assign g[15469] = b[12] & g[7278];
assign g[11375] = a[12] & g[7279];
assign g[15470] = b[12] & g[7279];
assign g[11376] = a[12] & g[7280];
assign g[15471] = b[12] & g[7280];
assign g[11377] = a[12] & g[7281];
assign g[15472] = b[12] & g[7281];
assign g[11378] = a[12] & g[7282];
assign g[15473] = b[12] & g[7282];
assign g[11379] = a[12] & g[7283];
assign g[15474] = b[12] & g[7283];
assign g[11380] = a[12] & g[7284];
assign g[15475] = b[12] & g[7284];
assign g[11381] = a[12] & g[7285];
assign g[15476] = b[12] & g[7285];
assign g[11382] = a[12] & g[7286];
assign g[15477] = b[12] & g[7286];
assign g[11383] = a[12] & g[7287];
assign g[15478] = b[12] & g[7287];
assign g[11384] = a[12] & g[7288];
assign g[15479] = b[12] & g[7288];
assign g[11385] = a[12] & g[7289];
assign g[15480] = b[12] & g[7289];
assign g[11386] = a[12] & g[7290];
assign g[15481] = b[12] & g[7290];
assign g[11387] = a[12] & g[7291];
assign g[15482] = b[12] & g[7291];
assign g[11388] = a[12] & g[7292];
assign g[15483] = b[12] & g[7292];
assign g[11389] = a[12] & g[7293];
assign g[15484] = b[12] & g[7293];
assign g[11390] = a[12] & g[7294];
assign g[15485] = b[12] & g[7294];
assign g[11391] = a[12] & g[7295];
assign g[15486] = b[12] & g[7295];
assign g[11392] = a[12] & g[7296];
assign g[15487] = b[12] & g[7296];
assign g[11393] = a[12] & g[7297];
assign g[15488] = b[12] & g[7297];
assign g[11394] = a[12] & g[7298];
assign g[15489] = b[12] & g[7298];
assign g[11395] = a[12] & g[7299];
assign g[15490] = b[12] & g[7299];
assign g[11396] = a[12] & g[7300];
assign g[15491] = b[12] & g[7300];
assign g[11397] = a[12] & g[7301];
assign g[15492] = b[12] & g[7301];
assign g[11398] = a[12] & g[7302];
assign g[15493] = b[12] & g[7302];
assign g[11399] = a[12] & g[7303];
assign g[15494] = b[12] & g[7303];
assign g[11400] = a[12] & g[7304];
assign g[15495] = b[12] & g[7304];
assign g[11401] = a[12] & g[7305];
assign g[15496] = b[12] & g[7305];
assign g[11402] = a[12] & g[7306];
assign g[15497] = b[12] & g[7306];
assign g[11403] = a[12] & g[7307];
assign g[15498] = b[12] & g[7307];
assign g[11404] = a[12] & g[7308];
assign g[15499] = b[12] & g[7308];
assign g[11405] = a[12] & g[7309];
assign g[15500] = b[12] & g[7309];
assign g[11406] = a[12] & g[7310];
assign g[15501] = b[12] & g[7310];
assign g[11407] = a[12] & g[7311];
assign g[15502] = b[12] & g[7311];
assign g[11408] = a[12] & g[7312];
assign g[15503] = b[12] & g[7312];
assign g[11409] = a[12] & g[7313];
assign g[15504] = b[12] & g[7313];
assign g[11410] = a[12] & g[7314];
assign g[15505] = b[12] & g[7314];
assign g[11411] = a[12] & g[7315];
assign g[15506] = b[12] & g[7315];
assign g[11412] = a[12] & g[7316];
assign g[15507] = b[12] & g[7316];
assign g[11413] = a[12] & g[7317];
assign g[15508] = b[12] & g[7317];
assign g[11414] = a[12] & g[7318];
assign g[15509] = b[12] & g[7318];
assign g[11415] = a[12] & g[7319];
assign g[15510] = b[12] & g[7319];
assign g[11416] = a[12] & g[7320];
assign g[15511] = b[12] & g[7320];
assign g[11417] = a[12] & g[7321];
assign g[15512] = b[12] & g[7321];
assign g[11418] = a[12] & g[7322];
assign g[15513] = b[12] & g[7322];
assign g[11419] = a[12] & g[7323];
assign g[15514] = b[12] & g[7323];
assign g[11420] = a[12] & g[7324];
assign g[15515] = b[12] & g[7324];
assign g[11421] = a[12] & g[7325];
assign g[15516] = b[12] & g[7325];
assign g[11422] = a[12] & g[7326];
assign g[15517] = b[12] & g[7326];
assign g[11423] = a[12] & g[7327];
assign g[15518] = b[12] & g[7327];
assign g[11424] = a[12] & g[7328];
assign g[15519] = b[12] & g[7328];
assign g[11425] = a[12] & g[7329];
assign g[15520] = b[12] & g[7329];
assign g[11426] = a[12] & g[7330];
assign g[15521] = b[12] & g[7330];
assign g[11427] = a[12] & g[7331];
assign g[15522] = b[12] & g[7331];
assign g[11428] = a[12] & g[7332];
assign g[15523] = b[12] & g[7332];
assign g[11429] = a[12] & g[7333];
assign g[15524] = b[12] & g[7333];
assign g[11430] = a[12] & g[7334];
assign g[15525] = b[12] & g[7334];
assign g[11431] = a[12] & g[7335];
assign g[15526] = b[12] & g[7335];
assign g[11432] = a[12] & g[7336];
assign g[15527] = b[12] & g[7336];
assign g[11433] = a[12] & g[7337];
assign g[15528] = b[12] & g[7337];
assign g[11434] = a[12] & g[7338];
assign g[15529] = b[12] & g[7338];
assign g[11435] = a[12] & g[7339];
assign g[15530] = b[12] & g[7339];
assign g[11436] = a[12] & g[7340];
assign g[15531] = b[12] & g[7340];
assign g[11437] = a[12] & g[7341];
assign g[15532] = b[12] & g[7341];
assign g[11438] = a[12] & g[7342];
assign g[15533] = b[12] & g[7342];
assign g[11439] = a[12] & g[7343];
assign g[15534] = b[12] & g[7343];
assign g[11440] = a[12] & g[7344];
assign g[15535] = b[12] & g[7344];
assign g[11441] = a[12] & g[7345];
assign g[15536] = b[12] & g[7345];
assign g[11442] = a[12] & g[7346];
assign g[15537] = b[12] & g[7346];
assign g[11443] = a[12] & g[7347];
assign g[15538] = b[12] & g[7347];
assign g[11444] = a[12] & g[7348];
assign g[15539] = b[12] & g[7348];
assign g[11445] = a[12] & g[7349];
assign g[15540] = b[12] & g[7349];
assign g[11446] = a[12] & g[7350];
assign g[15541] = b[12] & g[7350];
assign g[11447] = a[12] & g[7351];
assign g[15542] = b[12] & g[7351];
assign g[11448] = a[12] & g[7352];
assign g[15543] = b[12] & g[7352];
assign g[11449] = a[12] & g[7353];
assign g[15544] = b[12] & g[7353];
assign g[11450] = a[12] & g[7354];
assign g[15545] = b[12] & g[7354];
assign g[11451] = a[12] & g[7355];
assign g[15546] = b[12] & g[7355];
assign g[11452] = a[12] & g[7356];
assign g[15547] = b[12] & g[7356];
assign g[11453] = a[12] & g[7357];
assign g[15548] = b[12] & g[7357];
assign g[11454] = a[12] & g[7358];
assign g[15549] = b[12] & g[7358];
assign g[11455] = a[12] & g[7359];
assign g[15550] = b[12] & g[7359];
assign g[11456] = a[12] & g[7360];
assign g[15551] = b[12] & g[7360];
assign g[11457] = a[12] & g[7361];
assign g[15552] = b[12] & g[7361];
assign g[11458] = a[12] & g[7362];
assign g[15553] = b[12] & g[7362];
assign g[11459] = a[12] & g[7363];
assign g[15554] = b[12] & g[7363];
assign g[11460] = a[12] & g[7364];
assign g[15555] = b[12] & g[7364];
assign g[11461] = a[12] & g[7365];
assign g[15556] = b[12] & g[7365];
assign g[11462] = a[12] & g[7366];
assign g[15557] = b[12] & g[7366];
assign g[11463] = a[12] & g[7367];
assign g[15558] = b[12] & g[7367];
assign g[11464] = a[12] & g[7368];
assign g[15559] = b[12] & g[7368];
assign g[11465] = a[12] & g[7369];
assign g[15560] = b[12] & g[7369];
assign g[11466] = a[12] & g[7370];
assign g[15561] = b[12] & g[7370];
assign g[11467] = a[12] & g[7371];
assign g[15562] = b[12] & g[7371];
assign g[11468] = a[12] & g[7372];
assign g[15563] = b[12] & g[7372];
assign g[11469] = a[12] & g[7373];
assign g[15564] = b[12] & g[7373];
assign g[11470] = a[12] & g[7374];
assign g[15565] = b[12] & g[7374];
assign g[11471] = a[12] & g[7375];
assign g[15566] = b[12] & g[7375];
assign g[11472] = a[12] & g[7376];
assign g[15567] = b[12] & g[7376];
assign g[11473] = a[12] & g[7377];
assign g[15568] = b[12] & g[7377];
assign g[11474] = a[12] & g[7378];
assign g[15569] = b[12] & g[7378];
assign g[11475] = a[12] & g[7379];
assign g[15570] = b[12] & g[7379];
assign g[11476] = a[12] & g[7380];
assign g[15571] = b[12] & g[7380];
assign g[11477] = a[12] & g[7381];
assign g[15572] = b[12] & g[7381];
assign g[11478] = a[12] & g[7382];
assign g[15573] = b[12] & g[7382];
assign g[11479] = a[12] & g[7383];
assign g[15574] = b[12] & g[7383];
assign g[11480] = a[12] & g[7384];
assign g[15575] = b[12] & g[7384];
assign g[11481] = a[12] & g[7385];
assign g[15576] = b[12] & g[7385];
assign g[11482] = a[12] & g[7386];
assign g[15577] = b[12] & g[7386];
assign g[11483] = a[12] & g[7387];
assign g[15578] = b[12] & g[7387];
assign g[11484] = a[12] & g[7388];
assign g[15579] = b[12] & g[7388];
assign g[11485] = a[12] & g[7389];
assign g[15580] = b[12] & g[7389];
assign g[11486] = a[12] & g[7390];
assign g[15581] = b[12] & g[7390];
assign g[11487] = a[12] & g[7391];
assign g[15582] = b[12] & g[7391];
assign g[11488] = a[12] & g[7392];
assign g[15583] = b[12] & g[7392];
assign g[11489] = a[12] & g[7393];
assign g[15584] = b[12] & g[7393];
assign g[11490] = a[12] & g[7394];
assign g[15585] = b[12] & g[7394];
assign g[11491] = a[12] & g[7395];
assign g[15586] = b[12] & g[7395];
assign g[11492] = a[12] & g[7396];
assign g[15587] = b[12] & g[7396];
assign g[11493] = a[12] & g[7397];
assign g[15588] = b[12] & g[7397];
assign g[11494] = a[12] & g[7398];
assign g[15589] = b[12] & g[7398];
assign g[11495] = a[12] & g[7399];
assign g[15590] = b[12] & g[7399];
assign g[11496] = a[12] & g[7400];
assign g[15591] = b[12] & g[7400];
assign g[11497] = a[12] & g[7401];
assign g[15592] = b[12] & g[7401];
assign g[11498] = a[12] & g[7402];
assign g[15593] = b[12] & g[7402];
assign g[11499] = a[12] & g[7403];
assign g[15594] = b[12] & g[7403];
assign g[11500] = a[12] & g[7404];
assign g[15595] = b[12] & g[7404];
assign g[11501] = a[12] & g[7405];
assign g[15596] = b[12] & g[7405];
assign g[11502] = a[12] & g[7406];
assign g[15597] = b[12] & g[7406];
assign g[11503] = a[12] & g[7407];
assign g[15598] = b[12] & g[7407];
assign g[11504] = a[12] & g[7408];
assign g[15599] = b[12] & g[7408];
assign g[11505] = a[12] & g[7409];
assign g[15600] = b[12] & g[7409];
assign g[11506] = a[12] & g[7410];
assign g[15601] = b[12] & g[7410];
assign g[11507] = a[12] & g[7411];
assign g[15602] = b[12] & g[7411];
assign g[11508] = a[12] & g[7412];
assign g[15603] = b[12] & g[7412];
assign g[11509] = a[12] & g[7413];
assign g[15604] = b[12] & g[7413];
assign g[11510] = a[12] & g[7414];
assign g[15605] = b[12] & g[7414];
assign g[11511] = a[12] & g[7415];
assign g[15606] = b[12] & g[7415];
assign g[11512] = a[12] & g[7416];
assign g[15607] = b[12] & g[7416];
assign g[11513] = a[12] & g[7417];
assign g[15608] = b[12] & g[7417];
assign g[11514] = a[12] & g[7418];
assign g[15609] = b[12] & g[7418];
assign g[11515] = a[12] & g[7419];
assign g[15610] = b[12] & g[7419];
assign g[11516] = a[12] & g[7420];
assign g[15611] = b[12] & g[7420];
assign g[11517] = a[12] & g[7421];
assign g[15612] = b[12] & g[7421];
assign g[11518] = a[12] & g[7422];
assign g[15613] = b[12] & g[7422];
assign g[11519] = a[12] & g[7423];
assign g[15614] = b[12] & g[7423];
assign g[11520] = a[12] & g[7424];
assign g[15615] = b[12] & g[7424];
assign g[11521] = a[12] & g[7425];
assign g[15616] = b[12] & g[7425];
assign g[11522] = a[12] & g[7426];
assign g[15617] = b[12] & g[7426];
assign g[11523] = a[12] & g[7427];
assign g[15618] = b[12] & g[7427];
assign g[11524] = a[12] & g[7428];
assign g[15619] = b[12] & g[7428];
assign g[11525] = a[12] & g[7429];
assign g[15620] = b[12] & g[7429];
assign g[11526] = a[12] & g[7430];
assign g[15621] = b[12] & g[7430];
assign g[11527] = a[12] & g[7431];
assign g[15622] = b[12] & g[7431];
assign g[11528] = a[12] & g[7432];
assign g[15623] = b[12] & g[7432];
assign g[11529] = a[12] & g[7433];
assign g[15624] = b[12] & g[7433];
assign g[11530] = a[12] & g[7434];
assign g[15625] = b[12] & g[7434];
assign g[11531] = a[12] & g[7435];
assign g[15626] = b[12] & g[7435];
assign g[11532] = a[12] & g[7436];
assign g[15627] = b[12] & g[7436];
assign g[11533] = a[12] & g[7437];
assign g[15628] = b[12] & g[7437];
assign g[11534] = a[12] & g[7438];
assign g[15629] = b[12] & g[7438];
assign g[11535] = a[12] & g[7439];
assign g[15630] = b[12] & g[7439];
assign g[11536] = a[12] & g[7440];
assign g[15631] = b[12] & g[7440];
assign g[11537] = a[12] & g[7441];
assign g[15632] = b[12] & g[7441];
assign g[11538] = a[12] & g[7442];
assign g[15633] = b[12] & g[7442];
assign g[11539] = a[12] & g[7443];
assign g[15634] = b[12] & g[7443];
assign g[11540] = a[12] & g[7444];
assign g[15635] = b[12] & g[7444];
assign g[11541] = a[12] & g[7445];
assign g[15636] = b[12] & g[7445];
assign g[11542] = a[12] & g[7446];
assign g[15637] = b[12] & g[7446];
assign g[11543] = a[12] & g[7447];
assign g[15638] = b[12] & g[7447];
assign g[11544] = a[12] & g[7448];
assign g[15639] = b[12] & g[7448];
assign g[11545] = a[12] & g[7449];
assign g[15640] = b[12] & g[7449];
assign g[11546] = a[12] & g[7450];
assign g[15641] = b[12] & g[7450];
assign g[11547] = a[12] & g[7451];
assign g[15642] = b[12] & g[7451];
assign g[11548] = a[12] & g[7452];
assign g[15643] = b[12] & g[7452];
assign g[11549] = a[12] & g[7453];
assign g[15644] = b[12] & g[7453];
assign g[11550] = a[12] & g[7454];
assign g[15645] = b[12] & g[7454];
assign g[11551] = a[12] & g[7455];
assign g[15646] = b[12] & g[7455];
assign g[11552] = a[12] & g[7456];
assign g[15647] = b[12] & g[7456];
assign g[11553] = a[12] & g[7457];
assign g[15648] = b[12] & g[7457];
assign g[11554] = a[12] & g[7458];
assign g[15649] = b[12] & g[7458];
assign g[11555] = a[12] & g[7459];
assign g[15650] = b[12] & g[7459];
assign g[11556] = a[12] & g[7460];
assign g[15651] = b[12] & g[7460];
assign g[11557] = a[12] & g[7461];
assign g[15652] = b[12] & g[7461];
assign g[11558] = a[12] & g[7462];
assign g[15653] = b[12] & g[7462];
assign g[11559] = a[12] & g[7463];
assign g[15654] = b[12] & g[7463];
assign g[11560] = a[12] & g[7464];
assign g[15655] = b[12] & g[7464];
assign g[11561] = a[12] & g[7465];
assign g[15656] = b[12] & g[7465];
assign g[11562] = a[12] & g[7466];
assign g[15657] = b[12] & g[7466];
assign g[11563] = a[12] & g[7467];
assign g[15658] = b[12] & g[7467];
assign g[11564] = a[12] & g[7468];
assign g[15659] = b[12] & g[7468];
assign g[11565] = a[12] & g[7469];
assign g[15660] = b[12] & g[7469];
assign g[11566] = a[12] & g[7470];
assign g[15661] = b[12] & g[7470];
assign g[11567] = a[12] & g[7471];
assign g[15662] = b[12] & g[7471];
assign g[11568] = a[12] & g[7472];
assign g[15663] = b[12] & g[7472];
assign g[11569] = a[12] & g[7473];
assign g[15664] = b[12] & g[7473];
assign g[11570] = a[12] & g[7474];
assign g[15665] = b[12] & g[7474];
assign g[11571] = a[12] & g[7475];
assign g[15666] = b[12] & g[7475];
assign g[11572] = a[12] & g[7476];
assign g[15667] = b[12] & g[7476];
assign g[11573] = a[12] & g[7477];
assign g[15668] = b[12] & g[7477];
assign g[11574] = a[12] & g[7478];
assign g[15669] = b[12] & g[7478];
assign g[11575] = a[12] & g[7479];
assign g[15670] = b[12] & g[7479];
assign g[11576] = a[12] & g[7480];
assign g[15671] = b[12] & g[7480];
assign g[11577] = a[12] & g[7481];
assign g[15672] = b[12] & g[7481];
assign g[11578] = a[12] & g[7482];
assign g[15673] = b[12] & g[7482];
assign g[11579] = a[12] & g[7483];
assign g[15674] = b[12] & g[7483];
assign g[11580] = a[12] & g[7484];
assign g[15675] = b[12] & g[7484];
assign g[11581] = a[12] & g[7485];
assign g[15676] = b[12] & g[7485];
assign g[11582] = a[12] & g[7486];
assign g[15677] = b[12] & g[7486];
assign g[11583] = a[12] & g[7487];
assign g[15678] = b[12] & g[7487];
assign g[11584] = a[12] & g[7488];
assign g[15679] = b[12] & g[7488];
assign g[11585] = a[12] & g[7489];
assign g[15680] = b[12] & g[7489];
assign g[11586] = a[12] & g[7490];
assign g[15681] = b[12] & g[7490];
assign g[11587] = a[12] & g[7491];
assign g[15682] = b[12] & g[7491];
assign g[11588] = a[12] & g[7492];
assign g[15683] = b[12] & g[7492];
assign g[11589] = a[12] & g[7493];
assign g[15684] = b[12] & g[7493];
assign g[11590] = a[12] & g[7494];
assign g[15685] = b[12] & g[7494];
assign g[11591] = a[12] & g[7495];
assign g[15686] = b[12] & g[7495];
assign g[11592] = a[12] & g[7496];
assign g[15687] = b[12] & g[7496];
assign g[11593] = a[12] & g[7497];
assign g[15688] = b[12] & g[7497];
assign g[11594] = a[12] & g[7498];
assign g[15689] = b[12] & g[7498];
assign g[11595] = a[12] & g[7499];
assign g[15690] = b[12] & g[7499];
assign g[11596] = a[12] & g[7500];
assign g[15691] = b[12] & g[7500];
assign g[11597] = a[12] & g[7501];
assign g[15692] = b[12] & g[7501];
assign g[11598] = a[12] & g[7502];
assign g[15693] = b[12] & g[7502];
assign g[11599] = a[12] & g[7503];
assign g[15694] = b[12] & g[7503];
assign g[11600] = a[12] & g[7504];
assign g[15695] = b[12] & g[7504];
assign g[11601] = a[12] & g[7505];
assign g[15696] = b[12] & g[7505];
assign g[11602] = a[12] & g[7506];
assign g[15697] = b[12] & g[7506];
assign g[11603] = a[12] & g[7507];
assign g[15698] = b[12] & g[7507];
assign g[11604] = a[12] & g[7508];
assign g[15699] = b[12] & g[7508];
assign g[11605] = a[12] & g[7509];
assign g[15700] = b[12] & g[7509];
assign g[11606] = a[12] & g[7510];
assign g[15701] = b[12] & g[7510];
assign g[11607] = a[12] & g[7511];
assign g[15702] = b[12] & g[7511];
assign g[11608] = a[12] & g[7512];
assign g[15703] = b[12] & g[7512];
assign g[11609] = a[12] & g[7513];
assign g[15704] = b[12] & g[7513];
assign g[11610] = a[12] & g[7514];
assign g[15705] = b[12] & g[7514];
assign g[11611] = a[12] & g[7515];
assign g[15706] = b[12] & g[7515];
assign g[11612] = a[12] & g[7516];
assign g[15707] = b[12] & g[7516];
assign g[11613] = a[12] & g[7517];
assign g[15708] = b[12] & g[7517];
assign g[11614] = a[12] & g[7518];
assign g[15709] = b[12] & g[7518];
assign g[11615] = a[12] & g[7519];
assign g[15710] = b[12] & g[7519];
assign g[11616] = a[12] & g[7520];
assign g[15711] = b[12] & g[7520];
assign g[11617] = a[12] & g[7521];
assign g[15712] = b[12] & g[7521];
assign g[11618] = a[12] & g[7522];
assign g[15713] = b[12] & g[7522];
assign g[11619] = a[12] & g[7523];
assign g[15714] = b[12] & g[7523];
assign g[11620] = a[12] & g[7524];
assign g[15715] = b[12] & g[7524];
assign g[11621] = a[12] & g[7525];
assign g[15716] = b[12] & g[7525];
assign g[11622] = a[12] & g[7526];
assign g[15717] = b[12] & g[7526];
assign g[11623] = a[12] & g[7527];
assign g[15718] = b[12] & g[7527];
assign g[11624] = a[12] & g[7528];
assign g[15719] = b[12] & g[7528];
assign g[11625] = a[12] & g[7529];
assign g[15720] = b[12] & g[7529];
assign g[11626] = a[12] & g[7530];
assign g[15721] = b[12] & g[7530];
assign g[11627] = a[12] & g[7531];
assign g[15722] = b[12] & g[7531];
assign g[11628] = a[12] & g[7532];
assign g[15723] = b[12] & g[7532];
assign g[11629] = a[12] & g[7533];
assign g[15724] = b[12] & g[7533];
assign g[11630] = a[12] & g[7534];
assign g[15725] = b[12] & g[7534];
assign g[11631] = a[12] & g[7535];
assign g[15726] = b[12] & g[7535];
assign g[11632] = a[12] & g[7536];
assign g[15727] = b[12] & g[7536];
assign g[11633] = a[12] & g[7537];
assign g[15728] = b[12] & g[7537];
assign g[11634] = a[12] & g[7538];
assign g[15729] = b[12] & g[7538];
assign g[11635] = a[12] & g[7539];
assign g[15730] = b[12] & g[7539];
assign g[11636] = a[12] & g[7540];
assign g[15731] = b[12] & g[7540];
assign g[11637] = a[12] & g[7541];
assign g[15732] = b[12] & g[7541];
assign g[11638] = a[12] & g[7542];
assign g[15733] = b[12] & g[7542];
assign g[11639] = a[12] & g[7543];
assign g[15734] = b[12] & g[7543];
assign g[11640] = a[12] & g[7544];
assign g[15735] = b[12] & g[7544];
assign g[11641] = a[12] & g[7545];
assign g[15736] = b[12] & g[7545];
assign g[11642] = a[12] & g[7546];
assign g[15737] = b[12] & g[7546];
assign g[11643] = a[12] & g[7547];
assign g[15738] = b[12] & g[7547];
assign g[11644] = a[12] & g[7548];
assign g[15739] = b[12] & g[7548];
assign g[11645] = a[12] & g[7549];
assign g[15740] = b[12] & g[7549];
assign g[11646] = a[12] & g[7550];
assign g[15741] = b[12] & g[7550];
assign g[11647] = a[12] & g[7551];
assign g[15742] = b[12] & g[7551];
assign g[11648] = a[12] & g[7552];
assign g[15743] = b[12] & g[7552];
assign g[11649] = a[12] & g[7553];
assign g[15744] = b[12] & g[7553];
assign g[11650] = a[12] & g[7554];
assign g[15745] = b[12] & g[7554];
assign g[11651] = a[12] & g[7555];
assign g[15746] = b[12] & g[7555];
assign g[11652] = a[12] & g[7556];
assign g[15747] = b[12] & g[7556];
assign g[11653] = a[12] & g[7557];
assign g[15748] = b[12] & g[7557];
assign g[11654] = a[12] & g[7558];
assign g[15749] = b[12] & g[7558];
assign g[11655] = a[12] & g[7559];
assign g[15750] = b[12] & g[7559];
assign g[11656] = a[12] & g[7560];
assign g[15751] = b[12] & g[7560];
assign g[11657] = a[12] & g[7561];
assign g[15752] = b[12] & g[7561];
assign g[11658] = a[12] & g[7562];
assign g[15753] = b[12] & g[7562];
assign g[11659] = a[12] & g[7563];
assign g[15754] = b[12] & g[7563];
assign g[11660] = a[12] & g[7564];
assign g[15755] = b[12] & g[7564];
assign g[11661] = a[12] & g[7565];
assign g[15756] = b[12] & g[7565];
assign g[11662] = a[12] & g[7566];
assign g[15757] = b[12] & g[7566];
assign g[11663] = a[12] & g[7567];
assign g[15758] = b[12] & g[7567];
assign g[11664] = a[12] & g[7568];
assign g[15759] = b[12] & g[7568];
assign g[11665] = a[12] & g[7569];
assign g[15760] = b[12] & g[7569];
assign g[11666] = a[12] & g[7570];
assign g[15761] = b[12] & g[7570];
assign g[11667] = a[12] & g[7571];
assign g[15762] = b[12] & g[7571];
assign g[11668] = a[12] & g[7572];
assign g[15763] = b[12] & g[7572];
assign g[11669] = a[12] & g[7573];
assign g[15764] = b[12] & g[7573];
assign g[11670] = a[12] & g[7574];
assign g[15765] = b[12] & g[7574];
assign g[11671] = a[12] & g[7575];
assign g[15766] = b[12] & g[7575];
assign g[11672] = a[12] & g[7576];
assign g[15767] = b[12] & g[7576];
assign g[11673] = a[12] & g[7577];
assign g[15768] = b[12] & g[7577];
assign g[11674] = a[12] & g[7578];
assign g[15769] = b[12] & g[7578];
assign g[11675] = a[12] & g[7579];
assign g[15770] = b[12] & g[7579];
assign g[11676] = a[12] & g[7580];
assign g[15771] = b[12] & g[7580];
assign g[11677] = a[12] & g[7581];
assign g[15772] = b[12] & g[7581];
assign g[11678] = a[12] & g[7582];
assign g[15773] = b[12] & g[7582];
assign g[11679] = a[12] & g[7583];
assign g[15774] = b[12] & g[7583];
assign g[11680] = a[12] & g[7584];
assign g[15775] = b[12] & g[7584];
assign g[11681] = a[12] & g[7585];
assign g[15776] = b[12] & g[7585];
assign g[11682] = a[12] & g[7586];
assign g[15777] = b[12] & g[7586];
assign g[11683] = a[12] & g[7587];
assign g[15778] = b[12] & g[7587];
assign g[11684] = a[12] & g[7588];
assign g[15779] = b[12] & g[7588];
assign g[11685] = a[12] & g[7589];
assign g[15780] = b[12] & g[7589];
assign g[11686] = a[12] & g[7590];
assign g[15781] = b[12] & g[7590];
assign g[11687] = a[12] & g[7591];
assign g[15782] = b[12] & g[7591];
assign g[11688] = a[12] & g[7592];
assign g[15783] = b[12] & g[7592];
assign g[11689] = a[12] & g[7593];
assign g[15784] = b[12] & g[7593];
assign g[11690] = a[12] & g[7594];
assign g[15785] = b[12] & g[7594];
assign g[11691] = a[12] & g[7595];
assign g[15786] = b[12] & g[7595];
assign g[11692] = a[12] & g[7596];
assign g[15787] = b[12] & g[7596];
assign g[11693] = a[12] & g[7597];
assign g[15788] = b[12] & g[7597];
assign g[11694] = a[12] & g[7598];
assign g[15789] = b[12] & g[7598];
assign g[11695] = a[12] & g[7599];
assign g[15790] = b[12] & g[7599];
assign g[11696] = a[12] & g[7600];
assign g[15791] = b[12] & g[7600];
assign g[11697] = a[12] & g[7601];
assign g[15792] = b[12] & g[7601];
assign g[11698] = a[12] & g[7602];
assign g[15793] = b[12] & g[7602];
assign g[11699] = a[12] & g[7603];
assign g[15794] = b[12] & g[7603];
assign g[11700] = a[12] & g[7604];
assign g[15795] = b[12] & g[7604];
assign g[11701] = a[12] & g[7605];
assign g[15796] = b[12] & g[7605];
assign g[11702] = a[12] & g[7606];
assign g[15797] = b[12] & g[7606];
assign g[11703] = a[12] & g[7607];
assign g[15798] = b[12] & g[7607];
assign g[11704] = a[12] & g[7608];
assign g[15799] = b[12] & g[7608];
assign g[11705] = a[12] & g[7609];
assign g[15800] = b[12] & g[7609];
assign g[11706] = a[12] & g[7610];
assign g[15801] = b[12] & g[7610];
assign g[11707] = a[12] & g[7611];
assign g[15802] = b[12] & g[7611];
assign g[11708] = a[12] & g[7612];
assign g[15803] = b[12] & g[7612];
assign g[11709] = a[12] & g[7613];
assign g[15804] = b[12] & g[7613];
assign g[11710] = a[12] & g[7614];
assign g[15805] = b[12] & g[7614];
assign g[11711] = a[12] & g[7615];
assign g[15806] = b[12] & g[7615];
assign g[11712] = a[12] & g[7616];
assign g[15807] = b[12] & g[7616];
assign g[11713] = a[12] & g[7617];
assign g[15808] = b[12] & g[7617];
assign g[11714] = a[12] & g[7618];
assign g[15809] = b[12] & g[7618];
assign g[11715] = a[12] & g[7619];
assign g[15810] = b[12] & g[7619];
assign g[11716] = a[12] & g[7620];
assign g[15811] = b[12] & g[7620];
assign g[11717] = a[12] & g[7621];
assign g[15812] = b[12] & g[7621];
assign g[11718] = a[12] & g[7622];
assign g[15813] = b[12] & g[7622];
assign g[11719] = a[12] & g[7623];
assign g[15814] = b[12] & g[7623];
assign g[11720] = a[12] & g[7624];
assign g[15815] = b[12] & g[7624];
assign g[11721] = a[12] & g[7625];
assign g[15816] = b[12] & g[7625];
assign g[11722] = a[12] & g[7626];
assign g[15817] = b[12] & g[7626];
assign g[11723] = a[12] & g[7627];
assign g[15818] = b[12] & g[7627];
assign g[11724] = a[12] & g[7628];
assign g[15819] = b[12] & g[7628];
assign g[11725] = a[12] & g[7629];
assign g[15820] = b[12] & g[7629];
assign g[11726] = a[12] & g[7630];
assign g[15821] = b[12] & g[7630];
assign g[11727] = a[12] & g[7631];
assign g[15822] = b[12] & g[7631];
assign g[11728] = a[12] & g[7632];
assign g[15823] = b[12] & g[7632];
assign g[11729] = a[12] & g[7633];
assign g[15824] = b[12] & g[7633];
assign g[11730] = a[12] & g[7634];
assign g[15825] = b[12] & g[7634];
assign g[11731] = a[12] & g[7635];
assign g[15826] = b[12] & g[7635];
assign g[11732] = a[12] & g[7636];
assign g[15827] = b[12] & g[7636];
assign g[11733] = a[12] & g[7637];
assign g[15828] = b[12] & g[7637];
assign g[11734] = a[12] & g[7638];
assign g[15829] = b[12] & g[7638];
assign g[11735] = a[12] & g[7639];
assign g[15830] = b[12] & g[7639];
assign g[11736] = a[12] & g[7640];
assign g[15831] = b[12] & g[7640];
assign g[11737] = a[12] & g[7641];
assign g[15832] = b[12] & g[7641];
assign g[11738] = a[12] & g[7642];
assign g[15833] = b[12] & g[7642];
assign g[11739] = a[12] & g[7643];
assign g[15834] = b[12] & g[7643];
assign g[11740] = a[12] & g[7644];
assign g[15835] = b[12] & g[7644];
assign g[11741] = a[12] & g[7645];
assign g[15836] = b[12] & g[7645];
assign g[11742] = a[12] & g[7646];
assign g[15837] = b[12] & g[7646];
assign g[11743] = a[12] & g[7647];
assign g[15838] = b[12] & g[7647];
assign g[11744] = a[12] & g[7648];
assign g[15839] = b[12] & g[7648];
assign g[11745] = a[12] & g[7649];
assign g[15840] = b[12] & g[7649];
assign g[11746] = a[12] & g[7650];
assign g[15841] = b[12] & g[7650];
assign g[11747] = a[12] & g[7651];
assign g[15842] = b[12] & g[7651];
assign g[11748] = a[12] & g[7652];
assign g[15843] = b[12] & g[7652];
assign g[11749] = a[12] & g[7653];
assign g[15844] = b[12] & g[7653];
assign g[11750] = a[12] & g[7654];
assign g[15845] = b[12] & g[7654];
assign g[11751] = a[12] & g[7655];
assign g[15846] = b[12] & g[7655];
assign g[11752] = a[12] & g[7656];
assign g[15847] = b[12] & g[7656];
assign g[11753] = a[12] & g[7657];
assign g[15848] = b[12] & g[7657];
assign g[11754] = a[12] & g[7658];
assign g[15849] = b[12] & g[7658];
assign g[11755] = a[12] & g[7659];
assign g[15850] = b[12] & g[7659];
assign g[11756] = a[12] & g[7660];
assign g[15851] = b[12] & g[7660];
assign g[11757] = a[12] & g[7661];
assign g[15852] = b[12] & g[7661];
assign g[11758] = a[12] & g[7662];
assign g[15853] = b[12] & g[7662];
assign g[11759] = a[12] & g[7663];
assign g[15854] = b[12] & g[7663];
assign g[11760] = a[12] & g[7664];
assign g[15855] = b[12] & g[7664];
assign g[11761] = a[12] & g[7665];
assign g[15856] = b[12] & g[7665];
assign g[11762] = a[12] & g[7666];
assign g[15857] = b[12] & g[7666];
assign g[11763] = a[12] & g[7667];
assign g[15858] = b[12] & g[7667];
assign g[11764] = a[12] & g[7668];
assign g[15859] = b[12] & g[7668];
assign g[11765] = a[12] & g[7669];
assign g[15860] = b[12] & g[7669];
assign g[11766] = a[12] & g[7670];
assign g[15861] = b[12] & g[7670];
assign g[11767] = a[12] & g[7671];
assign g[15862] = b[12] & g[7671];
assign g[11768] = a[12] & g[7672];
assign g[15863] = b[12] & g[7672];
assign g[11769] = a[12] & g[7673];
assign g[15864] = b[12] & g[7673];
assign g[11770] = a[12] & g[7674];
assign g[15865] = b[12] & g[7674];
assign g[11771] = a[12] & g[7675];
assign g[15866] = b[12] & g[7675];
assign g[11772] = a[12] & g[7676];
assign g[15867] = b[12] & g[7676];
assign g[11773] = a[12] & g[7677];
assign g[15868] = b[12] & g[7677];
assign g[11774] = a[12] & g[7678];
assign g[15869] = b[12] & g[7678];
assign g[11775] = a[12] & g[7679];
assign g[15870] = b[12] & g[7679];
assign g[11776] = a[12] & g[7680];
assign g[15871] = b[12] & g[7680];
assign g[11777] = a[12] & g[7681];
assign g[15872] = b[12] & g[7681];
assign g[11778] = a[12] & g[7682];
assign g[15873] = b[12] & g[7682];
assign g[11779] = a[12] & g[7683];
assign g[15874] = b[12] & g[7683];
assign g[11780] = a[12] & g[7684];
assign g[15875] = b[12] & g[7684];
assign g[11781] = a[12] & g[7685];
assign g[15876] = b[12] & g[7685];
assign g[11782] = a[12] & g[7686];
assign g[15877] = b[12] & g[7686];
assign g[11783] = a[12] & g[7687];
assign g[15878] = b[12] & g[7687];
assign g[11784] = a[12] & g[7688];
assign g[15879] = b[12] & g[7688];
assign g[11785] = a[12] & g[7689];
assign g[15880] = b[12] & g[7689];
assign g[11786] = a[12] & g[7690];
assign g[15881] = b[12] & g[7690];
assign g[11787] = a[12] & g[7691];
assign g[15882] = b[12] & g[7691];
assign g[11788] = a[12] & g[7692];
assign g[15883] = b[12] & g[7692];
assign g[11789] = a[12] & g[7693];
assign g[15884] = b[12] & g[7693];
assign g[11790] = a[12] & g[7694];
assign g[15885] = b[12] & g[7694];
assign g[11791] = a[12] & g[7695];
assign g[15886] = b[12] & g[7695];
assign g[11792] = a[12] & g[7696];
assign g[15887] = b[12] & g[7696];
assign g[11793] = a[12] & g[7697];
assign g[15888] = b[12] & g[7697];
assign g[11794] = a[12] & g[7698];
assign g[15889] = b[12] & g[7698];
assign g[11795] = a[12] & g[7699];
assign g[15890] = b[12] & g[7699];
assign g[11796] = a[12] & g[7700];
assign g[15891] = b[12] & g[7700];
assign g[11797] = a[12] & g[7701];
assign g[15892] = b[12] & g[7701];
assign g[11798] = a[12] & g[7702];
assign g[15893] = b[12] & g[7702];
assign g[11799] = a[12] & g[7703];
assign g[15894] = b[12] & g[7703];
assign g[11800] = a[12] & g[7704];
assign g[15895] = b[12] & g[7704];
assign g[11801] = a[12] & g[7705];
assign g[15896] = b[12] & g[7705];
assign g[11802] = a[12] & g[7706];
assign g[15897] = b[12] & g[7706];
assign g[11803] = a[12] & g[7707];
assign g[15898] = b[12] & g[7707];
assign g[11804] = a[12] & g[7708];
assign g[15899] = b[12] & g[7708];
assign g[11805] = a[12] & g[7709];
assign g[15900] = b[12] & g[7709];
assign g[11806] = a[12] & g[7710];
assign g[15901] = b[12] & g[7710];
assign g[11807] = a[12] & g[7711];
assign g[15902] = b[12] & g[7711];
assign g[11808] = a[12] & g[7712];
assign g[15903] = b[12] & g[7712];
assign g[11809] = a[12] & g[7713];
assign g[15904] = b[12] & g[7713];
assign g[11810] = a[12] & g[7714];
assign g[15905] = b[12] & g[7714];
assign g[11811] = a[12] & g[7715];
assign g[15906] = b[12] & g[7715];
assign g[11812] = a[12] & g[7716];
assign g[15907] = b[12] & g[7716];
assign g[11813] = a[12] & g[7717];
assign g[15908] = b[12] & g[7717];
assign g[11814] = a[12] & g[7718];
assign g[15909] = b[12] & g[7718];
assign g[11815] = a[12] & g[7719];
assign g[15910] = b[12] & g[7719];
assign g[11816] = a[12] & g[7720];
assign g[15911] = b[12] & g[7720];
assign g[11817] = a[12] & g[7721];
assign g[15912] = b[12] & g[7721];
assign g[11818] = a[12] & g[7722];
assign g[15913] = b[12] & g[7722];
assign g[11819] = a[12] & g[7723];
assign g[15914] = b[12] & g[7723];
assign g[11820] = a[12] & g[7724];
assign g[15915] = b[12] & g[7724];
assign g[11821] = a[12] & g[7725];
assign g[15916] = b[12] & g[7725];
assign g[11822] = a[12] & g[7726];
assign g[15917] = b[12] & g[7726];
assign g[11823] = a[12] & g[7727];
assign g[15918] = b[12] & g[7727];
assign g[11824] = a[12] & g[7728];
assign g[15919] = b[12] & g[7728];
assign g[11825] = a[12] & g[7729];
assign g[15920] = b[12] & g[7729];
assign g[11826] = a[12] & g[7730];
assign g[15921] = b[12] & g[7730];
assign g[11827] = a[12] & g[7731];
assign g[15922] = b[12] & g[7731];
assign g[11828] = a[12] & g[7732];
assign g[15923] = b[12] & g[7732];
assign g[11829] = a[12] & g[7733];
assign g[15924] = b[12] & g[7733];
assign g[11830] = a[12] & g[7734];
assign g[15925] = b[12] & g[7734];
assign g[11831] = a[12] & g[7735];
assign g[15926] = b[12] & g[7735];
assign g[11832] = a[12] & g[7736];
assign g[15927] = b[12] & g[7736];
assign g[11833] = a[12] & g[7737];
assign g[15928] = b[12] & g[7737];
assign g[11834] = a[12] & g[7738];
assign g[15929] = b[12] & g[7738];
assign g[11835] = a[12] & g[7739];
assign g[15930] = b[12] & g[7739];
assign g[11836] = a[12] & g[7740];
assign g[15931] = b[12] & g[7740];
assign g[11837] = a[12] & g[7741];
assign g[15932] = b[12] & g[7741];
assign g[11838] = a[12] & g[7742];
assign g[15933] = b[12] & g[7742];
assign g[11839] = a[12] & g[7743];
assign g[15934] = b[12] & g[7743];
assign g[11840] = a[12] & g[7744];
assign g[15935] = b[12] & g[7744];
assign g[11841] = a[12] & g[7745];
assign g[15936] = b[12] & g[7745];
assign g[11842] = a[12] & g[7746];
assign g[15937] = b[12] & g[7746];
assign g[11843] = a[12] & g[7747];
assign g[15938] = b[12] & g[7747];
assign g[11844] = a[12] & g[7748];
assign g[15939] = b[12] & g[7748];
assign g[11845] = a[12] & g[7749];
assign g[15940] = b[12] & g[7749];
assign g[11846] = a[12] & g[7750];
assign g[15941] = b[12] & g[7750];
assign g[11847] = a[12] & g[7751];
assign g[15942] = b[12] & g[7751];
assign g[11848] = a[12] & g[7752];
assign g[15943] = b[12] & g[7752];
assign g[11849] = a[12] & g[7753];
assign g[15944] = b[12] & g[7753];
assign g[11850] = a[12] & g[7754];
assign g[15945] = b[12] & g[7754];
assign g[11851] = a[12] & g[7755];
assign g[15946] = b[12] & g[7755];
assign g[11852] = a[12] & g[7756];
assign g[15947] = b[12] & g[7756];
assign g[11853] = a[12] & g[7757];
assign g[15948] = b[12] & g[7757];
assign g[11854] = a[12] & g[7758];
assign g[15949] = b[12] & g[7758];
assign g[11855] = a[12] & g[7759];
assign g[15950] = b[12] & g[7759];
assign g[11856] = a[12] & g[7760];
assign g[15951] = b[12] & g[7760];
assign g[11857] = a[12] & g[7761];
assign g[15952] = b[12] & g[7761];
assign g[11858] = a[12] & g[7762];
assign g[15953] = b[12] & g[7762];
assign g[11859] = a[12] & g[7763];
assign g[15954] = b[12] & g[7763];
assign g[11860] = a[12] & g[7764];
assign g[15955] = b[12] & g[7764];
assign g[11861] = a[12] & g[7765];
assign g[15956] = b[12] & g[7765];
assign g[11862] = a[12] & g[7766];
assign g[15957] = b[12] & g[7766];
assign g[11863] = a[12] & g[7767];
assign g[15958] = b[12] & g[7767];
assign g[11864] = a[12] & g[7768];
assign g[15959] = b[12] & g[7768];
assign g[11865] = a[12] & g[7769];
assign g[15960] = b[12] & g[7769];
assign g[11866] = a[12] & g[7770];
assign g[15961] = b[12] & g[7770];
assign g[11867] = a[12] & g[7771];
assign g[15962] = b[12] & g[7771];
assign g[11868] = a[12] & g[7772];
assign g[15963] = b[12] & g[7772];
assign g[11869] = a[12] & g[7773];
assign g[15964] = b[12] & g[7773];
assign g[11870] = a[12] & g[7774];
assign g[15965] = b[12] & g[7774];
assign g[11871] = a[12] & g[7775];
assign g[15966] = b[12] & g[7775];
assign g[11872] = a[12] & g[7776];
assign g[15967] = b[12] & g[7776];
assign g[11873] = a[12] & g[7777];
assign g[15968] = b[12] & g[7777];
assign g[11874] = a[12] & g[7778];
assign g[15969] = b[12] & g[7778];
assign g[11875] = a[12] & g[7779];
assign g[15970] = b[12] & g[7779];
assign g[11876] = a[12] & g[7780];
assign g[15971] = b[12] & g[7780];
assign g[11877] = a[12] & g[7781];
assign g[15972] = b[12] & g[7781];
assign g[11878] = a[12] & g[7782];
assign g[15973] = b[12] & g[7782];
assign g[11879] = a[12] & g[7783];
assign g[15974] = b[12] & g[7783];
assign g[11880] = a[12] & g[7784];
assign g[15975] = b[12] & g[7784];
assign g[11881] = a[12] & g[7785];
assign g[15976] = b[12] & g[7785];
assign g[11882] = a[12] & g[7786];
assign g[15977] = b[12] & g[7786];
assign g[11883] = a[12] & g[7787];
assign g[15978] = b[12] & g[7787];
assign g[11884] = a[12] & g[7788];
assign g[15979] = b[12] & g[7788];
assign g[11885] = a[12] & g[7789];
assign g[15980] = b[12] & g[7789];
assign g[11886] = a[12] & g[7790];
assign g[15981] = b[12] & g[7790];
assign g[11887] = a[12] & g[7791];
assign g[15982] = b[12] & g[7791];
assign g[11888] = a[12] & g[7792];
assign g[15983] = b[12] & g[7792];
assign g[11889] = a[12] & g[7793];
assign g[15984] = b[12] & g[7793];
assign g[11890] = a[12] & g[7794];
assign g[15985] = b[12] & g[7794];
assign g[11891] = a[12] & g[7795];
assign g[15986] = b[12] & g[7795];
assign g[11892] = a[12] & g[7796];
assign g[15987] = b[12] & g[7796];
assign g[11893] = a[12] & g[7797];
assign g[15988] = b[12] & g[7797];
assign g[11894] = a[12] & g[7798];
assign g[15989] = b[12] & g[7798];
assign g[11895] = a[12] & g[7799];
assign g[15990] = b[12] & g[7799];
assign g[11896] = a[12] & g[7800];
assign g[15991] = b[12] & g[7800];
assign g[11897] = a[12] & g[7801];
assign g[15992] = b[12] & g[7801];
assign g[11898] = a[12] & g[7802];
assign g[15993] = b[12] & g[7802];
assign g[11899] = a[12] & g[7803];
assign g[15994] = b[12] & g[7803];
assign g[11900] = a[12] & g[7804];
assign g[15995] = b[12] & g[7804];
assign g[11901] = a[12] & g[7805];
assign g[15996] = b[12] & g[7805];
assign g[11902] = a[12] & g[7806];
assign g[15997] = b[12] & g[7806];
assign g[11903] = a[12] & g[7807];
assign g[15998] = b[12] & g[7807];
assign g[11904] = a[12] & g[7808];
assign g[15999] = b[12] & g[7808];
assign g[11905] = a[12] & g[7809];
assign g[16000] = b[12] & g[7809];
assign g[11906] = a[12] & g[7810];
assign g[16001] = b[12] & g[7810];
assign g[11907] = a[12] & g[7811];
assign g[16002] = b[12] & g[7811];
assign g[11908] = a[12] & g[7812];
assign g[16003] = b[12] & g[7812];
assign g[11909] = a[12] & g[7813];
assign g[16004] = b[12] & g[7813];
assign g[11910] = a[12] & g[7814];
assign g[16005] = b[12] & g[7814];
assign g[11911] = a[12] & g[7815];
assign g[16006] = b[12] & g[7815];
assign g[11912] = a[12] & g[7816];
assign g[16007] = b[12] & g[7816];
assign g[11913] = a[12] & g[7817];
assign g[16008] = b[12] & g[7817];
assign g[11914] = a[12] & g[7818];
assign g[16009] = b[12] & g[7818];
assign g[11915] = a[12] & g[7819];
assign g[16010] = b[12] & g[7819];
assign g[11916] = a[12] & g[7820];
assign g[16011] = b[12] & g[7820];
assign g[11917] = a[12] & g[7821];
assign g[16012] = b[12] & g[7821];
assign g[11918] = a[12] & g[7822];
assign g[16013] = b[12] & g[7822];
assign g[11919] = a[12] & g[7823];
assign g[16014] = b[12] & g[7823];
assign g[11920] = a[12] & g[7824];
assign g[16015] = b[12] & g[7824];
assign g[11921] = a[12] & g[7825];
assign g[16016] = b[12] & g[7825];
assign g[11922] = a[12] & g[7826];
assign g[16017] = b[12] & g[7826];
assign g[11923] = a[12] & g[7827];
assign g[16018] = b[12] & g[7827];
assign g[11924] = a[12] & g[7828];
assign g[16019] = b[12] & g[7828];
assign g[11925] = a[12] & g[7829];
assign g[16020] = b[12] & g[7829];
assign g[11926] = a[12] & g[7830];
assign g[16021] = b[12] & g[7830];
assign g[11927] = a[12] & g[7831];
assign g[16022] = b[12] & g[7831];
assign g[11928] = a[12] & g[7832];
assign g[16023] = b[12] & g[7832];
assign g[11929] = a[12] & g[7833];
assign g[16024] = b[12] & g[7833];
assign g[11930] = a[12] & g[7834];
assign g[16025] = b[12] & g[7834];
assign g[11931] = a[12] & g[7835];
assign g[16026] = b[12] & g[7835];
assign g[11932] = a[12] & g[7836];
assign g[16027] = b[12] & g[7836];
assign g[11933] = a[12] & g[7837];
assign g[16028] = b[12] & g[7837];
assign g[11934] = a[12] & g[7838];
assign g[16029] = b[12] & g[7838];
assign g[11935] = a[12] & g[7839];
assign g[16030] = b[12] & g[7839];
assign g[11936] = a[12] & g[7840];
assign g[16031] = b[12] & g[7840];
assign g[11937] = a[12] & g[7841];
assign g[16032] = b[12] & g[7841];
assign g[11938] = a[12] & g[7842];
assign g[16033] = b[12] & g[7842];
assign g[11939] = a[12] & g[7843];
assign g[16034] = b[12] & g[7843];
assign g[11940] = a[12] & g[7844];
assign g[16035] = b[12] & g[7844];
assign g[11941] = a[12] & g[7845];
assign g[16036] = b[12] & g[7845];
assign g[11942] = a[12] & g[7846];
assign g[16037] = b[12] & g[7846];
assign g[11943] = a[12] & g[7847];
assign g[16038] = b[12] & g[7847];
assign g[11944] = a[12] & g[7848];
assign g[16039] = b[12] & g[7848];
assign g[11945] = a[12] & g[7849];
assign g[16040] = b[12] & g[7849];
assign g[11946] = a[12] & g[7850];
assign g[16041] = b[12] & g[7850];
assign g[11947] = a[12] & g[7851];
assign g[16042] = b[12] & g[7851];
assign g[11948] = a[12] & g[7852];
assign g[16043] = b[12] & g[7852];
assign g[11949] = a[12] & g[7853];
assign g[16044] = b[12] & g[7853];
assign g[11950] = a[12] & g[7854];
assign g[16045] = b[12] & g[7854];
assign g[11951] = a[12] & g[7855];
assign g[16046] = b[12] & g[7855];
assign g[11952] = a[12] & g[7856];
assign g[16047] = b[12] & g[7856];
assign g[11953] = a[12] & g[7857];
assign g[16048] = b[12] & g[7857];
assign g[11954] = a[12] & g[7858];
assign g[16049] = b[12] & g[7858];
assign g[11955] = a[12] & g[7859];
assign g[16050] = b[12] & g[7859];
assign g[11956] = a[12] & g[7860];
assign g[16051] = b[12] & g[7860];
assign g[11957] = a[12] & g[7861];
assign g[16052] = b[12] & g[7861];
assign g[11958] = a[12] & g[7862];
assign g[16053] = b[12] & g[7862];
assign g[11959] = a[12] & g[7863];
assign g[16054] = b[12] & g[7863];
assign g[11960] = a[12] & g[7864];
assign g[16055] = b[12] & g[7864];
assign g[11961] = a[12] & g[7865];
assign g[16056] = b[12] & g[7865];
assign g[11962] = a[12] & g[7866];
assign g[16057] = b[12] & g[7866];
assign g[11963] = a[12] & g[7867];
assign g[16058] = b[12] & g[7867];
assign g[11964] = a[12] & g[7868];
assign g[16059] = b[12] & g[7868];
assign g[11965] = a[12] & g[7869];
assign g[16060] = b[12] & g[7869];
assign g[11966] = a[12] & g[7870];
assign g[16061] = b[12] & g[7870];
assign g[11967] = a[12] & g[7871];
assign g[16062] = b[12] & g[7871];
assign g[11968] = a[12] & g[7872];
assign g[16063] = b[12] & g[7872];
assign g[11969] = a[12] & g[7873];
assign g[16064] = b[12] & g[7873];
assign g[11970] = a[12] & g[7874];
assign g[16065] = b[12] & g[7874];
assign g[11971] = a[12] & g[7875];
assign g[16066] = b[12] & g[7875];
assign g[11972] = a[12] & g[7876];
assign g[16067] = b[12] & g[7876];
assign g[11973] = a[12] & g[7877];
assign g[16068] = b[12] & g[7877];
assign g[11974] = a[12] & g[7878];
assign g[16069] = b[12] & g[7878];
assign g[11975] = a[12] & g[7879];
assign g[16070] = b[12] & g[7879];
assign g[11976] = a[12] & g[7880];
assign g[16071] = b[12] & g[7880];
assign g[11977] = a[12] & g[7881];
assign g[16072] = b[12] & g[7881];
assign g[11978] = a[12] & g[7882];
assign g[16073] = b[12] & g[7882];
assign g[11979] = a[12] & g[7883];
assign g[16074] = b[12] & g[7883];
assign g[11980] = a[12] & g[7884];
assign g[16075] = b[12] & g[7884];
assign g[11981] = a[12] & g[7885];
assign g[16076] = b[12] & g[7885];
assign g[11982] = a[12] & g[7886];
assign g[16077] = b[12] & g[7886];
assign g[11983] = a[12] & g[7887];
assign g[16078] = b[12] & g[7887];
assign g[11984] = a[12] & g[7888];
assign g[16079] = b[12] & g[7888];
assign g[11985] = a[12] & g[7889];
assign g[16080] = b[12] & g[7889];
assign g[11986] = a[12] & g[7890];
assign g[16081] = b[12] & g[7890];
assign g[11987] = a[12] & g[7891];
assign g[16082] = b[12] & g[7891];
assign g[11988] = a[12] & g[7892];
assign g[16083] = b[12] & g[7892];
assign g[11989] = a[12] & g[7893];
assign g[16084] = b[12] & g[7893];
assign g[11990] = a[12] & g[7894];
assign g[16085] = b[12] & g[7894];
assign g[11991] = a[12] & g[7895];
assign g[16086] = b[12] & g[7895];
assign g[11992] = a[12] & g[7896];
assign g[16087] = b[12] & g[7896];
assign g[11993] = a[12] & g[7897];
assign g[16088] = b[12] & g[7897];
assign g[11994] = a[12] & g[7898];
assign g[16089] = b[12] & g[7898];
assign g[11995] = a[12] & g[7899];
assign g[16090] = b[12] & g[7899];
assign g[11996] = a[12] & g[7900];
assign g[16091] = b[12] & g[7900];
assign g[11997] = a[12] & g[7901];
assign g[16092] = b[12] & g[7901];
assign g[11998] = a[12] & g[7902];
assign g[16093] = b[12] & g[7902];
assign g[11999] = a[12] & g[7903];
assign g[16094] = b[12] & g[7903];
assign g[12000] = a[12] & g[7904];
assign g[16095] = b[12] & g[7904];
assign g[12001] = a[12] & g[7905];
assign g[16096] = b[12] & g[7905];
assign g[12002] = a[12] & g[7906];
assign g[16097] = b[12] & g[7906];
assign g[12003] = a[12] & g[7907];
assign g[16098] = b[12] & g[7907];
assign g[12004] = a[12] & g[7908];
assign g[16099] = b[12] & g[7908];
assign g[12005] = a[12] & g[7909];
assign g[16100] = b[12] & g[7909];
assign g[12006] = a[12] & g[7910];
assign g[16101] = b[12] & g[7910];
assign g[12007] = a[12] & g[7911];
assign g[16102] = b[12] & g[7911];
assign g[12008] = a[12] & g[7912];
assign g[16103] = b[12] & g[7912];
assign g[12009] = a[12] & g[7913];
assign g[16104] = b[12] & g[7913];
assign g[12010] = a[12] & g[7914];
assign g[16105] = b[12] & g[7914];
assign g[12011] = a[12] & g[7915];
assign g[16106] = b[12] & g[7915];
assign g[12012] = a[12] & g[7916];
assign g[16107] = b[12] & g[7916];
assign g[12013] = a[12] & g[7917];
assign g[16108] = b[12] & g[7917];
assign g[12014] = a[12] & g[7918];
assign g[16109] = b[12] & g[7918];
assign g[12015] = a[12] & g[7919];
assign g[16110] = b[12] & g[7919];
assign g[12016] = a[12] & g[7920];
assign g[16111] = b[12] & g[7920];
assign g[12017] = a[12] & g[7921];
assign g[16112] = b[12] & g[7921];
assign g[12018] = a[12] & g[7922];
assign g[16113] = b[12] & g[7922];
assign g[12019] = a[12] & g[7923];
assign g[16114] = b[12] & g[7923];
assign g[12020] = a[12] & g[7924];
assign g[16115] = b[12] & g[7924];
assign g[12021] = a[12] & g[7925];
assign g[16116] = b[12] & g[7925];
assign g[12022] = a[12] & g[7926];
assign g[16117] = b[12] & g[7926];
assign g[12023] = a[12] & g[7927];
assign g[16118] = b[12] & g[7927];
assign g[12024] = a[12] & g[7928];
assign g[16119] = b[12] & g[7928];
assign g[12025] = a[12] & g[7929];
assign g[16120] = b[12] & g[7929];
assign g[12026] = a[12] & g[7930];
assign g[16121] = b[12] & g[7930];
assign g[12027] = a[12] & g[7931];
assign g[16122] = b[12] & g[7931];
assign g[12028] = a[12] & g[7932];
assign g[16123] = b[12] & g[7932];
assign g[12029] = a[12] & g[7933];
assign g[16124] = b[12] & g[7933];
assign g[12030] = a[12] & g[7934];
assign g[16125] = b[12] & g[7934];
assign g[12031] = a[12] & g[7935];
assign g[16126] = b[12] & g[7935];
assign g[12032] = a[12] & g[7936];
assign g[16127] = b[12] & g[7936];
assign g[12033] = a[12] & g[7937];
assign g[16128] = b[12] & g[7937];
assign g[12034] = a[12] & g[7938];
assign g[16129] = b[12] & g[7938];
assign g[12035] = a[12] & g[7939];
assign g[16130] = b[12] & g[7939];
assign g[12036] = a[12] & g[7940];
assign g[16131] = b[12] & g[7940];
assign g[12037] = a[12] & g[7941];
assign g[16132] = b[12] & g[7941];
assign g[12038] = a[12] & g[7942];
assign g[16133] = b[12] & g[7942];
assign g[12039] = a[12] & g[7943];
assign g[16134] = b[12] & g[7943];
assign g[12040] = a[12] & g[7944];
assign g[16135] = b[12] & g[7944];
assign g[12041] = a[12] & g[7945];
assign g[16136] = b[12] & g[7945];
assign g[12042] = a[12] & g[7946];
assign g[16137] = b[12] & g[7946];
assign g[12043] = a[12] & g[7947];
assign g[16138] = b[12] & g[7947];
assign g[12044] = a[12] & g[7948];
assign g[16139] = b[12] & g[7948];
assign g[12045] = a[12] & g[7949];
assign g[16140] = b[12] & g[7949];
assign g[12046] = a[12] & g[7950];
assign g[16141] = b[12] & g[7950];
assign g[12047] = a[12] & g[7951];
assign g[16142] = b[12] & g[7951];
assign g[12048] = a[12] & g[7952];
assign g[16143] = b[12] & g[7952];
assign g[12049] = a[12] & g[7953];
assign g[16144] = b[12] & g[7953];
assign g[12050] = a[12] & g[7954];
assign g[16145] = b[12] & g[7954];
assign g[12051] = a[12] & g[7955];
assign g[16146] = b[12] & g[7955];
assign g[12052] = a[12] & g[7956];
assign g[16147] = b[12] & g[7956];
assign g[12053] = a[12] & g[7957];
assign g[16148] = b[12] & g[7957];
assign g[12054] = a[12] & g[7958];
assign g[16149] = b[12] & g[7958];
assign g[12055] = a[12] & g[7959];
assign g[16150] = b[12] & g[7959];
assign g[12056] = a[12] & g[7960];
assign g[16151] = b[12] & g[7960];
assign g[12057] = a[12] & g[7961];
assign g[16152] = b[12] & g[7961];
assign g[12058] = a[12] & g[7962];
assign g[16153] = b[12] & g[7962];
assign g[12059] = a[12] & g[7963];
assign g[16154] = b[12] & g[7963];
assign g[12060] = a[12] & g[7964];
assign g[16155] = b[12] & g[7964];
assign g[12061] = a[12] & g[7965];
assign g[16156] = b[12] & g[7965];
assign g[12062] = a[12] & g[7966];
assign g[16157] = b[12] & g[7966];
assign g[12063] = a[12] & g[7967];
assign g[16158] = b[12] & g[7967];
assign g[12064] = a[12] & g[7968];
assign g[16159] = b[12] & g[7968];
assign g[12065] = a[12] & g[7969];
assign g[16160] = b[12] & g[7969];
assign g[12066] = a[12] & g[7970];
assign g[16161] = b[12] & g[7970];
assign g[12067] = a[12] & g[7971];
assign g[16162] = b[12] & g[7971];
assign g[12068] = a[12] & g[7972];
assign g[16163] = b[12] & g[7972];
assign g[12069] = a[12] & g[7973];
assign g[16164] = b[12] & g[7973];
assign g[12070] = a[12] & g[7974];
assign g[16165] = b[12] & g[7974];
assign g[12071] = a[12] & g[7975];
assign g[16166] = b[12] & g[7975];
assign g[12072] = a[12] & g[7976];
assign g[16167] = b[12] & g[7976];
assign g[12073] = a[12] & g[7977];
assign g[16168] = b[12] & g[7977];
assign g[12074] = a[12] & g[7978];
assign g[16169] = b[12] & g[7978];
assign g[12075] = a[12] & g[7979];
assign g[16170] = b[12] & g[7979];
assign g[12076] = a[12] & g[7980];
assign g[16171] = b[12] & g[7980];
assign g[12077] = a[12] & g[7981];
assign g[16172] = b[12] & g[7981];
assign g[12078] = a[12] & g[7982];
assign g[16173] = b[12] & g[7982];
assign g[12079] = a[12] & g[7983];
assign g[16174] = b[12] & g[7983];
assign g[12080] = a[12] & g[7984];
assign g[16175] = b[12] & g[7984];
assign g[12081] = a[12] & g[7985];
assign g[16176] = b[12] & g[7985];
assign g[12082] = a[12] & g[7986];
assign g[16177] = b[12] & g[7986];
assign g[12083] = a[12] & g[7987];
assign g[16178] = b[12] & g[7987];
assign g[12084] = a[12] & g[7988];
assign g[16179] = b[12] & g[7988];
assign g[12085] = a[12] & g[7989];
assign g[16180] = b[12] & g[7989];
assign g[12086] = a[12] & g[7990];
assign g[16181] = b[12] & g[7990];
assign g[12087] = a[12] & g[7991];
assign g[16182] = b[12] & g[7991];
assign g[12088] = a[12] & g[7992];
assign g[16183] = b[12] & g[7992];
assign g[12089] = a[12] & g[7993];
assign g[16184] = b[12] & g[7993];
assign g[12090] = a[12] & g[7994];
assign g[16185] = b[12] & g[7994];
assign g[12091] = a[12] & g[7995];
assign g[16186] = b[12] & g[7995];
assign g[12092] = a[12] & g[7996];
assign g[16187] = b[12] & g[7996];
assign g[12093] = a[12] & g[7997];
assign g[16188] = b[12] & g[7997];
assign g[12094] = a[12] & g[7998];
assign g[16189] = b[12] & g[7998];
assign g[12095] = a[12] & g[7999];
assign g[16190] = b[12] & g[7999];
assign g[12096] = a[12] & g[8000];
assign g[16191] = b[12] & g[8000];
assign g[12097] = a[12] & g[8001];
assign g[16192] = b[12] & g[8001];
assign g[12098] = a[12] & g[8002];
assign g[16193] = b[12] & g[8002];
assign g[12099] = a[12] & g[8003];
assign g[16194] = b[12] & g[8003];
assign g[12100] = a[12] & g[8004];
assign g[16195] = b[12] & g[8004];
assign g[12101] = a[12] & g[8005];
assign g[16196] = b[12] & g[8005];
assign g[12102] = a[12] & g[8006];
assign g[16197] = b[12] & g[8006];
assign g[12103] = a[12] & g[8007];
assign g[16198] = b[12] & g[8007];
assign g[12104] = a[12] & g[8008];
assign g[16199] = b[12] & g[8008];
assign g[12105] = a[12] & g[8009];
assign g[16200] = b[12] & g[8009];
assign g[12106] = a[12] & g[8010];
assign g[16201] = b[12] & g[8010];
assign g[12107] = a[12] & g[8011];
assign g[16202] = b[12] & g[8011];
assign g[12108] = a[12] & g[8012];
assign g[16203] = b[12] & g[8012];
assign g[12109] = a[12] & g[8013];
assign g[16204] = b[12] & g[8013];
assign g[12110] = a[12] & g[8014];
assign g[16205] = b[12] & g[8014];
assign g[12111] = a[12] & g[8015];
assign g[16206] = b[12] & g[8015];
assign g[12112] = a[12] & g[8016];
assign g[16207] = b[12] & g[8016];
assign g[12113] = a[12] & g[8017];
assign g[16208] = b[12] & g[8017];
assign g[12114] = a[12] & g[8018];
assign g[16209] = b[12] & g[8018];
assign g[12115] = a[12] & g[8019];
assign g[16210] = b[12] & g[8019];
assign g[12116] = a[12] & g[8020];
assign g[16211] = b[12] & g[8020];
assign g[12117] = a[12] & g[8021];
assign g[16212] = b[12] & g[8021];
assign g[12118] = a[12] & g[8022];
assign g[16213] = b[12] & g[8022];
assign g[12119] = a[12] & g[8023];
assign g[16214] = b[12] & g[8023];
assign g[12120] = a[12] & g[8024];
assign g[16215] = b[12] & g[8024];
assign g[12121] = a[12] & g[8025];
assign g[16216] = b[12] & g[8025];
assign g[12122] = a[12] & g[8026];
assign g[16217] = b[12] & g[8026];
assign g[12123] = a[12] & g[8027];
assign g[16218] = b[12] & g[8027];
assign g[12124] = a[12] & g[8028];
assign g[16219] = b[12] & g[8028];
assign g[12125] = a[12] & g[8029];
assign g[16220] = b[12] & g[8029];
assign g[12126] = a[12] & g[8030];
assign g[16221] = b[12] & g[8030];
assign g[12127] = a[12] & g[8031];
assign g[16222] = b[12] & g[8031];
assign g[12128] = a[12] & g[8032];
assign g[16223] = b[12] & g[8032];
assign g[12129] = a[12] & g[8033];
assign g[16224] = b[12] & g[8033];
assign g[12130] = a[12] & g[8034];
assign g[16225] = b[12] & g[8034];
assign g[12131] = a[12] & g[8035];
assign g[16226] = b[12] & g[8035];
assign g[12132] = a[12] & g[8036];
assign g[16227] = b[12] & g[8036];
assign g[12133] = a[12] & g[8037];
assign g[16228] = b[12] & g[8037];
assign g[12134] = a[12] & g[8038];
assign g[16229] = b[12] & g[8038];
assign g[12135] = a[12] & g[8039];
assign g[16230] = b[12] & g[8039];
assign g[12136] = a[12] & g[8040];
assign g[16231] = b[12] & g[8040];
assign g[12137] = a[12] & g[8041];
assign g[16232] = b[12] & g[8041];
assign g[12138] = a[12] & g[8042];
assign g[16233] = b[12] & g[8042];
assign g[12139] = a[12] & g[8043];
assign g[16234] = b[12] & g[8043];
assign g[12140] = a[12] & g[8044];
assign g[16235] = b[12] & g[8044];
assign g[12141] = a[12] & g[8045];
assign g[16236] = b[12] & g[8045];
assign g[12142] = a[12] & g[8046];
assign g[16237] = b[12] & g[8046];
assign g[12143] = a[12] & g[8047];
assign g[16238] = b[12] & g[8047];
assign g[12144] = a[12] & g[8048];
assign g[16239] = b[12] & g[8048];
assign g[12145] = a[12] & g[8049];
assign g[16240] = b[12] & g[8049];
assign g[12146] = a[12] & g[8050];
assign g[16241] = b[12] & g[8050];
assign g[12147] = a[12] & g[8051];
assign g[16242] = b[12] & g[8051];
assign g[12148] = a[12] & g[8052];
assign g[16243] = b[12] & g[8052];
assign g[12149] = a[12] & g[8053];
assign g[16244] = b[12] & g[8053];
assign g[12150] = a[12] & g[8054];
assign g[16245] = b[12] & g[8054];
assign g[12151] = a[12] & g[8055];
assign g[16246] = b[12] & g[8055];
assign g[12152] = a[12] & g[8056];
assign g[16247] = b[12] & g[8056];
assign g[12153] = a[12] & g[8057];
assign g[16248] = b[12] & g[8057];
assign g[12154] = a[12] & g[8058];
assign g[16249] = b[12] & g[8058];
assign g[12155] = a[12] & g[8059];
assign g[16250] = b[12] & g[8059];
assign g[12156] = a[12] & g[8060];
assign g[16251] = b[12] & g[8060];
assign g[12157] = a[12] & g[8061];
assign g[16252] = b[12] & g[8061];
assign g[12158] = a[12] & g[8062];
assign g[16253] = b[12] & g[8062];
assign g[12159] = a[12] & g[8063];
assign g[16254] = b[12] & g[8063];
assign g[12160] = a[12] & g[8064];
assign g[16255] = b[12] & g[8064];
assign g[12161] = a[12] & g[8065];
assign g[16256] = b[12] & g[8065];
assign g[12162] = a[12] & g[8066];
assign g[16257] = b[12] & g[8066];
assign g[12163] = a[12] & g[8067];
assign g[16258] = b[12] & g[8067];
assign g[12164] = a[12] & g[8068];
assign g[16259] = b[12] & g[8068];
assign g[12165] = a[12] & g[8069];
assign g[16260] = b[12] & g[8069];
assign g[12166] = a[12] & g[8070];
assign g[16261] = b[12] & g[8070];
assign g[12167] = a[12] & g[8071];
assign g[16262] = b[12] & g[8071];
assign g[12168] = a[12] & g[8072];
assign g[16263] = b[12] & g[8072];
assign g[12169] = a[12] & g[8073];
assign g[16264] = b[12] & g[8073];
assign g[12170] = a[12] & g[8074];
assign g[16265] = b[12] & g[8074];
assign g[12171] = a[12] & g[8075];
assign g[16266] = b[12] & g[8075];
assign g[12172] = a[12] & g[8076];
assign g[16267] = b[12] & g[8076];
assign g[12173] = a[12] & g[8077];
assign g[16268] = b[12] & g[8077];
assign g[12174] = a[12] & g[8078];
assign g[16269] = b[12] & g[8078];
assign g[12175] = a[12] & g[8079];
assign g[16270] = b[12] & g[8079];
assign g[12176] = a[12] & g[8080];
assign g[16271] = b[12] & g[8080];
assign g[12177] = a[12] & g[8081];
assign g[16272] = b[12] & g[8081];
assign g[12178] = a[12] & g[8082];
assign g[16273] = b[12] & g[8082];
assign g[12179] = a[12] & g[8083];
assign g[16274] = b[12] & g[8083];
assign g[12180] = a[12] & g[8084];
assign g[16275] = b[12] & g[8084];
assign g[12181] = a[12] & g[8085];
assign g[16276] = b[12] & g[8085];
assign g[12182] = a[12] & g[8086];
assign g[16277] = b[12] & g[8086];
assign g[12183] = a[12] & g[8087];
assign g[16278] = b[12] & g[8087];
assign g[12184] = a[12] & g[8088];
assign g[16279] = b[12] & g[8088];
assign g[12185] = a[12] & g[8089];
assign g[16280] = b[12] & g[8089];
assign g[12186] = a[12] & g[8090];
assign g[16281] = b[12] & g[8090];
assign g[12187] = a[12] & g[8091];
assign g[16282] = b[12] & g[8091];
assign g[12188] = a[12] & g[8092];
assign g[16283] = b[12] & g[8092];
assign g[12189] = a[12] & g[8093];
assign g[16284] = b[12] & g[8093];
assign g[12190] = a[12] & g[8094];
assign g[16285] = b[12] & g[8094];
assign g[12191] = a[12] & g[8095];
assign g[16286] = b[12] & g[8095];
assign g[12192] = a[12] & g[8096];
assign g[16287] = b[12] & g[8096];
assign g[12193] = a[12] & g[8097];
assign g[16288] = b[12] & g[8097];
assign g[12194] = a[12] & g[8098];
assign g[16289] = b[12] & g[8098];
assign g[12195] = a[12] & g[8099];
assign g[16290] = b[12] & g[8099];
assign g[12196] = a[12] & g[8100];
assign g[16291] = b[12] & g[8100];
assign g[12197] = a[12] & g[8101];
assign g[16292] = b[12] & g[8101];
assign g[12198] = a[12] & g[8102];
assign g[16293] = b[12] & g[8102];
assign g[12199] = a[12] & g[8103];
assign g[16294] = b[12] & g[8103];
assign g[12200] = a[12] & g[8104];
assign g[16295] = b[12] & g[8104];
assign g[12201] = a[12] & g[8105];
assign g[16296] = b[12] & g[8105];
assign g[12202] = a[12] & g[8106];
assign g[16297] = b[12] & g[8106];
assign g[12203] = a[12] & g[8107];
assign g[16298] = b[12] & g[8107];
assign g[12204] = a[12] & g[8108];
assign g[16299] = b[12] & g[8108];
assign g[12205] = a[12] & g[8109];
assign g[16300] = b[12] & g[8109];
assign g[12206] = a[12] & g[8110];
assign g[16301] = b[12] & g[8110];
assign g[12207] = a[12] & g[8111];
assign g[16302] = b[12] & g[8111];
assign g[12208] = a[12] & g[8112];
assign g[16303] = b[12] & g[8112];
assign g[12209] = a[12] & g[8113];
assign g[16304] = b[12] & g[8113];
assign g[12210] = a[12] & g[8114];
assign g[16305] = b[12] & g[8114];
assign g[12211] = a[12] & g[8115];
assign g[16306] = b[12] & g[8115];
assign g[12212] = a[12] & g[8116];
assign g[16307] = b[12] & g[8116];
assign g[12213] = a[12] & g[8117];
assign g[16308] = b[12] & g[8117];
assign g[12214] = a[12] & g[8118];
assign g[16309] = b[12] & g[8118];
assign g[12215] = a[12] & g[8119];
assign g[16310] = b[12] & g[8119];
assign g[12216] = a[12] & g[8120];
assign g[16311] = b[12] & g[8120];
assign g[12217] = a[12] & g[8121];
assign g[16312] = b[12] & g[8121];
assign g[12218] = a[12] & g[8122];
assign g[16313] = b[12] & g[8122];
assign g[12219] = a[12] & g[8123];
assign g[16314] = b[12] & g[8123];
assign g[12220] = a[12] & g[8124];
assign g[16315] = b[12] & g[8124];
assign g[12221] = a[12] & g[8125];
assign g[16316] = b[12] & g[8125];
assign g[12222] = a[12] & g[8126];
assign g[16317] = b[12] & g[8126];
assign g[12223] = a[12] & g[8127];
assign g[16318] = b[12] & g[8127];
assign g[12224] = a[12] & g[8128];
assign g[16319] = b[12] & g[8128];
assign g[12225] = a[12] & g[8129];
assign g[16320] = b[12] & g[8129];
assign g[12226] = a[12] & g[8130];
assign g[16321] = b[12] & g[8130];
assign g[12227] = a[12] & g[8131];
assign g[16322] = b[12] & g[8131];
assign g[12228] = a[12] & g[8132];
assign g[16323] = b[12] & g[8132];
assign g[12229] = a[12] & g[8133];
assign g[16324] = b[12] & g[8133];
assign g[12230] = a[12] & g[8134];
assign g[16325] = b[12] & g[8134];
assign g[12231] = a[12] & g[8135];
assign g[16326] = b[12] & g[8135];
assign g[12232] = a[12] & g[8136];
assign g[16327] = b[12] & g[8136];
assign g[12233] = a[12] & g[8137];
assign g[16328] = b[12] & g[8137];
assign g[12234] = a[12] & g[8138];
assign g[16329] = b[12] & g[8138];
assign g[12235] = a[12] & g[8139];
assign g[16330] = b[12] & g[8139];
assign g[12236] = a[12] & g[8140];
assign g[16331] = b[12] & g[8140];
assign g[12237] = a[12] & g[8141];
assign g[16332] = b[12] & g[8141];
assign g[12238] = a[12] & g[8142];
assign g[16333] = b[12] & g[8142];
assign g[12239] = a[12] & g[8143];
assign g[16334] = b[12] & g[8143];
assign g[12240] = a[12] & g[8144];
assign g[16335] = b[12] & g[8144];
assign g[12241] = a[12] & g[8145];
assign g[16336] = b[12] & g[8145];
assign g[12242] = a[12] & g[8146];
assign g[16337] = b[12] & g[8146];
assign g[12243] = a[12] & g[8147];
assign g[16338] = b[12] & g[8147];
assign g[12244] = a[12] & g[8148];
assign g[16339] = b[12] & g[8148];
assign g[12245] = a[12] & g[8149];
assign g[16340] = b[12] & g[8149];
assign g[12246] = a[12] & g[8150];
assign g[16341] = b[12] & g[8150];
assign g[12247] = a[12] & g[8151];
assign g[16342] = b[12] & g[8151];
assign g[12248] = a[12] & g[8152];
assign g[16343] = b[12] & g[8152];
assign g[12249] = a[12] & g[8153];
assign g[16344] = b[12] & g[8153];
assign g[12250] = a[12] & g[8154];
assign g[16345] = b[12] & g[8154];
assign g[12251] = a[12] & g[8155];
assign g[16346] = b[12] & g[8155];
assign g[12252] = a[12] & g[8156];
assign g[16347] = b[12] & g[8156];
assign g[12253] = a[12] & g[8157];
assign g[16348] = b[12] & g[8157];
assign g[12254] = a[12] & g[8158];
assign g[16349] = b[12] & g[8158];
assign g[12255] = a[12] & g[8159];
assign g[16350] = b[12] & g[8159];
assign g[12256] = a[12] & g[8160];
assign g[16351] = b[12] & g[8160];
assign g[12257] = a[12] & g[8161];
assign g[16352] = b[12] & g[8161];
assign g[12258] = a[12] & g[8162];
assign g[16353] = b[12] & g[8162];
assign g[12259] = a[12] & g[8163];
assign g[16354] = b[12] & g[8163];
assign g[12260] = a[12] & g[8164];
assign g[16355] = b[12] & g[8164];
assign g[12261] = a[12] & g[8165];
assign g[16356] = b[12] & g[8165];
assign g[12262] = a[12] & g[8166];
assign g[16357] = b[12] & g[8166];
assign g[12263] = a[12] & g[8167];
assign g[16358] = b[12] & g[8167];
assign g[12264] = a[12] & g[8168];
assign g[16359] = b[12] & g[8168];
assign g[12265] = a[12] & g[8169];
assign g[16360] = b[12] & g[8169];
assign g[12266] = a[12] & g[8170];
assign g[16361] = b[12] & g[8170];
assign g[12267] = a[12] & g[8171];
assign g[16362] = b[12] & g[8171];
assign g[12268] = a[12] & g[8172];
assign g[16363] = b[12] & g[8172];
assign g[12269] = a[12] & g[8173];
assign g[16364] = b[12] & g[8173];
assign g[12270] = a[12] & g[8174];
assign g[16365] = b[12] & g[8174];
assign g[12271] = a[12] & g[8175];
assign g[16366] = b[12] & g[8175];
assign g[12272] = a[12] & g[8176];
assign g[16367] = b[12] & g[8176];
assign g[12273] = a[12] & g[8177];
assign g[16368] = b[12] & g[8177];
//Assigning outputs for input bit 14
assign g[16369] = a[13] & b[13];
assign g[16370] = a[13] & g[8178];
assign g[24561] = b[13] & g[8178];
assign g[16371] = a[13] & g[8179];
assign g[24562] = b[13] & g[8179];
assign g[16372] = a[13] & g[8180];
assign g[24563] = b[13] & g[8180];
assign g[16373] = a[13] & g[8181];
assign g[24564] = b[13] & g[8181];
assign g[16374] = a[13] & g[8182];
assign g[24565] = b[13] & g[8182];
assign g[16375] = a[13] & g[8183];
assign g[24566] = b[13] & g[8183];
assign g[16376] = a[13] & g[8184];
assign g[24567] = b[13] & g[8184];
assign g[16377] = a[13] & g[8185];
assign g[24568] = b[13] & g[8185];
assign g[16378] = a[13] & g[8186];
assign g[24569] = b[13] & g[8186];
assign g[16379] = a[13] & g[8187];
assign g[24570] = b[13] & g[8187];
assign g[16380] = a[13] & g[8188];
assign g[24571] = b[13] & g[8188];
assign g[16381] = a[13] & g[8189];
assign g[24572] = b[13] & g[8189];
assign g[16382] = a[13] & g[8190];
assign g[24573] = b[13] & g[8190];
assign g[16383] = a[13] & g[8191];
assign g[24574] = b[13] & g[8191];
assign g[16384] = a[13] & g[8192];
assign g[24575] = b[13] & g[8192];
assign g[16385] = a[13] & g[8193];
assign g[24576] = b[13] & g[8193];
assign g[16386] = a[13] & g[8194];
assign g[24577] = b[13] & g[8194];
assign g[16387] = a[13] & g[8195];
assign g[24578] = b[13] & g[8195];
assign g[16388] = a[13] & g[8196];
assign g[24579] = b[13] & g[8196];
assign g[16389] = a[13] & g[8197];
assign g[24580] = b[13] & g[8197];
assign g[16390] = a[13] & g[8198];
assign g[24581] = b[13] & g[8198];
assign g[16391] = a[13] & g[8199];
assign g[24582] = b[13] & g[8199];
assign g[16392] = a[13] & g[8200];
assign g[24583] = b[13] & g[8200];
assign g[16393] = a[13] & g[8201];
assign g[24584] = b[13] & g[8201];
assign g[16394] = a[13] & g[8202];
assign g[24585] = b[13] & g[8202];
assign g[16395] = a[13] & g[8203];
assign g[24586] = b[13] & g[8203];
assign g[16396] = a[13] & g[8204];
assign g[24587] = b[13] & g[8204];
assign g[16397] = a[13] & g[8205];
assign g[24588] = b[13] & g[8205];
assign g[16398] = a[13] & g[8206];
assign g[24589] = b[13] & g[8206];
assign g[16399] = a[13] & g[8207];
assign g[24590] = b[13] & g[8207];
assign g[16400] = a[13] & g[8208];
assign g[24591] = b[13] & g[8208];
assign g[16401] = a[13] & g[8209];
assign g[24592] = b[13] & g[8209];
assign g[16402] = a[13] & g[8210];
assign g[24593] = b[13] & g[8210];
assign g[16403] = a[13] & g[8211];
assign g[24594] = b[13] & g[8211];
assign g[16404] = a[13] & g[8212];
assign g[24595] = b[13] & g[8212];
assign g[16405] = a[13] & g[8213];
assign g[24596] = b[13] & g[8213];
assign g[16406] = a[13] & g[8214];
assign g[24597] = b[13] & g[8214];
assign g[16407] = a[13] & g[8215];
assign g[24598] = b[13] & g[8215];
assign g[16408] = a[13] & g[8216];
assign g[24599] = b[13] & g[8216];
assign g[16409] = a[13] & g[8217];
assign g[24600] = b[13] & g[8217];
assign g[16410] = a[13] & g[8218];
assign g[24601] = b[13] & g[8218];
assign g[16411] = a[13] & g[8219];
assign g[24602] = b[13] & g[8219];
assign g[16412] = a[13] & g[8220];
assign g[24603] = b[13] & g[8220];
assign g[16413] = a[13] & g[8221];
assign g[24604] = b[13] & g[8221];
assign g[16414] = a[13] & g[8222];
assign g[24605] = b[13] & g[8222];
assign g[16415] = a[13] & g[8223];
assign g[24606] = b[13] & g[8223];
assign g[16416] = a[13] & g[8224];
assign g[24607] = b[13] & g[8224];
assign g[16417] = a[13] & g[8225];
assign g[24608] = b[13] & g[8225];
assign g[16418] = a[13] & g[8226];
assign g[24609] = b[13] & g[8226];
assign g[16419] = a[13] & g[8227];
assign g[24610] = b[13] & g[8227];
assign g[16420] = a[13] & g[8228];
assign g[24611] = b[13] & g[8228];
assign g[16421] = a[13] & g[8229];
assign g[24612] = b[13] & g[8229];
assign g[16422] = a[13] & g[8230];
assign g[24613] = b[13] & g[8230];
assign g[16423] = a[13] & g[8231];
assign g[24614] = b[13] & g[8231];
assign g[16424] = a[13] & g[8232];
assign g[24615] = b[13] & g[8232];
assign g[16425] = a[13] & g[8233];
assign g[24616] = b[13] & g[8233];
assign g[16426] = a[13] & g[8234];
assign g[24617] = b[13] & g[8234];
assign g[16427] = a[13] & g[8235];
assign g[24618] = b[13] & g[8235];
assign g[16428] = a[13] & g[8236];
assign g[24619] = b[13] & g[8236];
assign g[16429] = a[13] & g[8237];
assign g[24620] = b[13] & g[8237];
assign g[16430] = a[13] & g[8238];
assign g[24621] = b[13] & g[8238];
assign g[16431] = a[13] & g[8239];
assign g[24622] = b[13] & g[8239];
assign g[16432] = a[13] & g[8240];
assign g[24623] = b[13] & g[8240];
assign g[16433] = a[13] & g[8241];
assign g[24624] = b[13] & g[8241];
assign g[16434] = a[13] & g[8242];
assign g[24625] = b[13] & g[8242];
assign g[16435] = a[13] & g[8243];
assign g[24626] = b[13] & g[8243];
assign g[16436] = a[13] & g[8244];
assign g[24627] = b[13] & g[8244];
assign g[16437] = a[13] & g[8245];
assign g[24628] = b[13] & g[8245];
assign g[16438] = a[13] & g[8246];
assign g[24629] = b[13] & g[8246];
assign g[16439] = a[13] & g[8247];
assign g[24630] = b[13] & g[8247];
assign g[16440] = a[13] & g[8248];
assign g[24631] = b[13] & g[8248];
assign g[16441] = a[13] & g[8249];
assign g[24632] = b[13] & g[8249];
assign g[16442] = a[13] & g[8250];
assign g[24633] = b[13] & g[8250];
assign g[16443] = a[13] & g[8251];
assign g[24634] = b[13] & g[8251];
assign g[16444] = a[13] & g[8252];
assign g[24635] = b[13] & g[8252];
assign g[16445] = a[13] & g[8253];
assign g[24636] = b[13] & g[8253];
assign g[16446] = a[13] & g[8254];
assign g[24637] = b[13] & g[8254];
assign g[16447] = a[13] & g[8255];
assign g[24638] = b[13] & g[8255];
assign g[16448] = a[13] & g[8256];
assign g[24639] = b[13] & g[8256];
assign g[16449] = a[13] & g[8257];
assign g[24640] = b[13] & g[8257];
assign g[16450] = a[13] & g[8258];
assign g[24641] = b[13] & g[8258];
assign g[16451] = a[13] & g[8259];
assign g[24642] = b[13] & g[8259];
assign g[16452] = a[13] & g[8260];
assign g[24643] = b[13] & g[8260];
assign g[16453] = a[13] & g[8261];
assign g[24644] = b[13] & g[8261];
assign g[16454] = a[13] & g[8262];
assign g[24645] = b[13] & g[8262];
assign g[16455] = a[13] & g[8263];
assign g[24646] = b[13] & g[8263];
assign g[16456] = a[13] & g[8264];
assign g[24647] = b[13] & g[8264];
assign g[16457] = a[13] & g[8265];
assign g[24648] = b[13] & g[8265];
assign g[16458] = a[13] & g[8266];
assign g[24649] = b[13] & g[8266];
assign g[16459] = a[13] & g[8267];
assign g[24650] = b[13] & g[8267];
assign g[16460] = a[13] & g[8268];
assign g[24651] = b[13] & g[8268];
assign g[16461] = a[13] & g[8269];
assign g[24652] = b[13] & g[8269];
assign g[16462] = a[13] & g[8270];
assign g[24653] = b[13] & g[8270];
assign g[16463] = a[13] & g[8271];
assign g[24654] = b[13] & g[8271];
assign g[16464] = a[13] & g[8272];
assign g[24655] = b[13] & g[8272];
assign g[16465] = a[13] & g[8273];
assign g[24656] = b[13] & g[8273];
assign g[16466] = a[13] & g[8274];
assign g[24657] = b[13] & g[8274];
assign g[16467] = a[13] & g[8275];
assign g[24658] = b[13] & g[8275];
assign g[16468] = a[13] & g[8276];
assign g[24659] = b[13] & g[8276];
assign g[16469] = a[13] & g[8277];
assign g[24660] = b[13] & g[8277];
assign g[16470] = a[13] & g[8278];
assign g[24661] = b[13] & g[8278];
assign g[16471] = a[13] & g[8279];
assign g[24662] = b[13] & g[8279];
assign g[16472] = a[13] & g[8280];
assign g[24663] = b[13] & g[8280];
assign g[16473] = a[13] & g[8281];
assign g[24664] = b[13] & g[8281];
assign g[16474] = a[13] & g[8282];
assign g[24665] = b[13] & g[8282];
assign g[16475] = a[13] & g[8283];
assign g[24666] = b[13] & g[8283];
assign g[16476] = a[13] & g[8284];
assign g[24667] = b[13] & g[8284];
assign g[16477] = a[13] & g[8285];
assign g[24668] = b[13] & g[8285];
assign g[16478] = a[13] & g[8286];
assign g[24669] = b[13] & g[8286];
assign g[16479] = a[13] & g[8287];
assign g[24670] = b[13] & g[8287];
assign g[16480] = a[13] & g[8288];
assign g[24671] = b[13] & g[8288];
assign g[16481] = a[13] & g[8289];
assign g[24672] = b[13] & g[8289];
assign g[16482] = a[13] & g[8290];
assign g[24673] = b[13] & g[8290];
assign g[16483] = a[13] & g[8291];
assign g[24674] = b[13] & g[8291];
assign g[16484] = a[13] & g[8292];
assign g[24675] = b[13] & g[8292];
assign g[16485] = a[13] & g[8293];
assign g[24676] = b[13] & g[8293];
assign g[16486] = a[13] & g[8294];
assign g[24677] = b[13] & g[8294];
assign g[16487] = a[13] & g[8295];
assign g[24678] = b[13] & g[8295];
assign g[16488] = a[13] & g[8296];
assign g[24679] = b[13] & g[8296];
assign g[16489] = a[13] & g[8297];
assign g[24680] = b[13] & g[8297];
assign g[16490] = a[13] & g[8298];
assign g[24681] = b[13] & g[8298];
assign g[16491] = a[13] & g[8299];
assign g[24682] = b[13] & g[8299];
assign g[16492] = a[13] & g[8300];
assign g[24683] = b[13] & g[8300];
assign g[16493] = a[13] & g[8301];
assign g[24684] = b[13] & g[8301];
assign g[16494] = a[13] & g[8302];
assign g[24685] = b[13] & g[8302];
assign g[16495] = a[13] & g[8303];
assign g[24686] = b[13] & g[8303];
assign g[16496] = a[13] & g[8304];
assign g[24687] = b[13] & g[8304];
assign g[16497] = a[13] & g[8305];
assign g[24688] = b[13] & g[8305];
assign g[16498] = a[13] & g[8306];
assign g[24689] = b[13] & g[8306];
assign g[16499] = a[13] & g[8307];
assign g[24690] = b[13] & g[8307];
assign g[16500] = a[13] & g[8308];
assign g[24691] = b[13] & g[8308];
assign g[16501] = a[13] & g[8309];
assign g[24692] = b[13] & g[8309];
assign g[16502] = a[13] & g[8310];
assign g[24693] = b[13] & g[8310];
assign g[16503] = a[13] & g[8311];
assign g[24694] = b[13] & g[8311];
assign g[16504] = a[13] & g[8312];
assign g[24695] = b[13] & g[8312];
assign g[16505] = a[13] & g[8313];
assign g[24696] = b[13] & g[8313];
assign g[16506] = a[13] & g[8314];
assign g[24697] = b[13] & g[8314];
assign g[16507] = a[13] & g[8315];
assign g[24698] = b[13] & g[8315];
assign g[16508] = a[13] & g[8316];
assign g[24699] = b[13] & g[8316];
assign g[16509] = a[13] & g[8317];
assign g[24700] = b[13] & g[8317];
assign g[16510] = a[13] & g[8318];
assign g[24701] = b[13] & g[8318];
assign g[16511] = a[13] & g[8319];
assign g[24702] = b[13] & g[8319];
assign g[16512] = a[13] & g[8320];
assign g[24703] = b[13] & g[8320];
assign g[16513] = a[13] & g[8321];
assign g[24704] = b[13] & g[8321];
assign g[16514] = a[13] & g[8322];
assign g[24705] = b[13] & g[8322];
assign g[16515] = a[13] & g[8323];
assign g[24706] = b[13] & g[8323];
assign g[16516] = a[13] & g[8324];
assign g[24707] = b[13] & g[8324];
assign g[16517] = a[13] & g[8325];
assign g[24708] = b[13] & g[8325];
assign g[16518] = a[13] & g[8326];
assign g[24709] = b[13] & g[8326];
assign g[16519] = a[13] & g[8327];
assign g[24710] = b[13] & g[8327];
assign g[16520] = a[13] & g[8328];
assign g[24711] = b[13] & g[8328];
assign g[16521] = a[13] & g[8329];
assign g[24712] = b[13] & g[8329];
assign g[16522] = a[13] & g[8330];
assign g[24713] = b[13] & g[8330];
assign g[16523] = a[13] & g[8331];
assign g[24714] = b[13] & g[8331];
assign g[16524] = a[13] & g[8332];
assign g[24715] = b[13] & g[8332];
assign g[16525] = a[13] & g[8333];
assign g[24716] = b[13] & g[8333];
assign g[16526] = a[13] & g[8334];
assign g[24717] = b[13] & g[8334];
assign g[16527] = a[13] & g[8335];
assign g[24718] = b[13] & g[8335];
assign g[16528] = a[13] & g[8336];
assign g[24719] = b[13] & g[8336];
assign g[16529] = a[13] & g[8337];
assign g[24720] = b[13] & g[8337];
assign g[16530] = a[13] & g[8338];
assign g[24721] = b[13] & g[8338];
assign g[16531] = a[13] & g[8339];
assign g[24722] = b[13] & g[8339];
assign g[16532] = a[13] & g[8340];
assign g[24723] = b[13] & g[8340];
assign g[16533] = a[13] & g[8341];
assign g[24724] = b[13] & g[8341];
assign g[16534] = a[13] & g[8342];
assign g[24725] = b[13] & g[8342];
assign g[16535] = a[13] & g[8343];
assign g[24726] = b[13] & g[8343];
assign g[16536] = a[13] & g[8344];
assign g[24727] = b[13] & g[8344];
assign g[16537] = a[13] & g[8345];
assign g[24728] = b[13] & g[8345];
assign g[16538] = a[13] & g[8346];
assign g[24729] = b[13] & g[8346];
assign g[16539] = a[13] & g[8347];
assign g[24730] = b[13] & g[8347];
assign g[16540] = a[13] & g[8348];
assign g[24731] = b[13] & g[8348];
assign g[16541] = a[13] & g[8349];
assign g[24732] = b[13] & g[8349];
assign g[16542] = a[13] & g[8350];
assign g[24733] = b[13] & g[8350];
assign g[16543] = a[13] & g[8351];
assign g[24734] = b[13] & g[8351];
assign g[16544] = a[13] & g[8352];
assign g[24735] = b[13] & g[8352];
assign g[16545] = a[13] & g[8353];
assign g[24736] = b[13] & g[8353];
assign g[16546] = a[13] & g[8354];
assign g[24737] = b[13] & g[8354];
assign g[16547] = a[13] & g[8355];
assign g[24738] = b[13] & g[8355];
assign g[16548] = a[13] & g[8356];
assign g[24739] = b[13] & g[8356];
assign g[16549] = a[13] & g[8357];
assign g[24740] = b[13] & g[8357];
assign g[16550] = a[13] & g[8358];
assign g[24741] = b[13] & g[8358];
assign g[16551] = a[13] & g[8359];
assign g[24742] = b[13] & g[8359];
assign g[16552] = a[13] & g[8360];
assign g[24743] = b[13] & g[8360];
assign g[16553] = a[13] & g[8361];
assign g[24744] = b[13] & g[8361];
assign g[16554] = a[13] & g[8362];
assign g[24745] = b[13] & g[8362];
assign g[16555] = a[13] & g[8363];
assign g[24746] = b[13] & g[8363];
assign g[16556] = a[13] & g[8364];
assign g[24747] = b[13] & g[8364];
assign g[16557] = a[13] & g[8365];
assign g[24748] = b[13] & g[8365];
assign g[16558] = a[13] & g[8366];
assign g[24749] = b[13] & g[8366];
assign g[16559] = a[13] & g[8367];
assign g[24750] = b[13] & g[8367];
assign g[16560] = a[13] & g[8368];
assign g[24751] = b[13] & g[8368];
assign g[16561] = a[13] & g[8369];
assign g[24752] = b[13] & g[8369];
assign g[16562] = a[13] & g[8370];
assign g[24753] = b[13] & g[8370];
assign g[16563] = a[13] & g[8371];
assign g[24754] = b[13] & g[8371];
assign g[16564] = a[13] & g[8372];
assign g[24755] = b[13] & g[8372];
assign g[16565] = a[13] & g[8373];
assign g[24756] = b[13] & g[8373];
assign g[16566] = a[13] & g[8374];
assign g[24757] = b[13] & g[8374];
assign g[16567] = a[13] & g[8375];
assign g[24758] = b[13] & g[8375];
assign g[16568] = a[13] & g[8376];
assign g[24759] = b[13] & g[8376];
assign g[16569] = a[13] & g[8377];
assign g[24760] = b[13] & g[8377];
assign g[16570] = a[13] & g[8378];
assign g[24761] = b[13] & g[8378];
assign g[16571] = a[13] & g[8379];
assign g[24762] = b[13] & g[8379];
assign g[16572] = a[13] & g[8380];
assign g[24763] = b[13] & g[8380];
assign g[16573] = a[13] & g[8381];
assign g[24764] = b[13] & g[8381];
assign g[16574] = a[13] & g[8382];
assign g[24765] = b[13] & g[8382];
assign g[16575] = a[13] & g[8383];
assign g[24766] = b[13] & g[8383];
assign g[16576] = a[13] & g[8384];
assign g[24767] = b[13] & g[8384];
assign g[16577] = a[13] & g[8385];
assign g[24768] = b[13] & g[8385];
assign g[16578] = a[13] & g[8386];
assign g[24769] = b[13] & g[8386];
assign g[16579] = a[13] & g[8387];
assign g[24770] = b[13] & g[8387];
assign g[16580] = a[13] & g[8388];
assign g[24771] = b[13] & g[8388];
assign g[16581] = a[13] & g[8389];
assign g[24772] = b[13] & g[8389];
assign g[16582] = a[13] & g[8390];
assign g[24773] = b[13] & g[8390];
assign g[16583] = a[13] & g[8391];
assign g[24774] = b[13] & g[8391];
assign g[16584] = a[13] & g[8392];
assign g[24775] = b[13] & g[8392];
assign g[16585] = a[13] & g[8393];
assign g[24776] = b[13] & g[8393];
assign g[16586] = a[13] & g[8394];
assign g[24777] = b[13] & g[8394];
assign g[16587] = a[13] & g[8395];
assign g[24778] = b[13] & g[8395];
assign g[16588] = a[13] & g[8396];
assign g[24779] = b[13] & g[8396];
assign g[16589] = a[13] & g[8397];
assign g[24780] = b[13] & g[8397];
assign g[16590] = a[13] & g[8398];
assign g[24781] = b[13] & g[8398];
assign g[16591] = a[13] & g[8399];
assign g[24782] = b[13] & g[8399];
assign g[16592] = a[13] & g[8400];
assign g[24783] = b[13] & g[8400];
assign g[16593] = a[13] & g[8401];
assign g[24784] = b[13] & g[8401];
assign g[16594] = a[13] & g[8402];
assign g[24785] = b[13] & g[8402];
assign g[16595] = a[13] & g[8403];
assign g[24786] = b[13] & g[8403];
assign g[16596] = a[13] & g[8404];
assign g[24787] = b[13] & g[8404];
assign g[16597] = a[13] & g[8405];
assign g[24788] = b[13] & g[8405];
assign g[16598] = a[13] & g[8406];
assign g[24789] = b[13] & g[8406];
assign g[16599] = a[13] & g[8407];
assign g[24790] = b[13] & g[8407];
assign g[16600] = a[13] & g[8408];
assign g[24791] = b[13] & g[8408];
assign g[16601] = a[13] & g[8409];
assign g[24792] = b[13] & g[8409];
assign g[16602] = a[13] & g[8410];
assign g[24793] = b[13] & g[8410];
assign g[16603] = a[13] & g[8411];
assign g[24794] = b[13] & g[8411];
assign g[16604] = a[13] & g[8412];
assign g[24795] = b[13] & g[8412];
assign g[16605] = a[13] & g[8413];
assign g[24796] = b[13] & g[8413];
assign g[16606] = a[13] & g[8414];
assign g[24797] = b[13] & g[8414];
assign g[16607] = a[13] & g[8415];
assign g[24798] = b[13] & g[8415];
assign g[16608] = a[13] & g[8416];
assign g[24799] = b[13] & g[8416];
assign g[16609] = a[13] & g[8417];
assign g[24800] = b[13] & g[8417];
assign g[16610] = a[13] & g[8418];
assign g[24801] = b[13] & g[8418];
assign g[16611] = a[13] & g[8419];
assign g[24802] = b[13] & g[8419];
assign g[16612] = a[13] & g[8420];
assign g[24803] = b[13] & g[8420];
assign g[16613] = a[13] & g[8421];
assign g[24804] = b[13] & g[8421];
assign g[16614] = a[13] & g[8422];
assign g[24805] = b[13] & g[8422];
assign g[16615] = a[13] & g[8423];
assign g[24806] = b[13] & g[8423];
assign g[16616] = a[13] & g[8424];
assign g[24807] = b[13] & g[8424];
assign g[16617] = a[13] & g[8425];
assign g[24808] = b[13] & g[8425];
assign g[16618] = a[13] & g[8426];
assign g[24809] = b[13] & g[8426];
assign g[16619] = a[13] & g[8427];
assign g[24810] = b[13] & g[8427];
assign g[16620] = a[13] & g[8428];
assign g[24811] = b[13] & g[8428];
assign g[16621] = a[13] & g[8429];
assign g[24812] = b[13] & g[8429];
assign g[16622] = a[13] & g[8430];
assign g[24813] = b[13] & g[8430];
assign g[16623] = a[13] & g[8431];
assign g[24814] = b[13] & g[8431];
assign g[16624] = a[13] & g[8432];
assign g[24815] = b[13] & g[8432];
assign g[16625] = a[13] & g[8433];
assign g[24816] = b[13] & g[8433];
assign g[16626] = a[13] & g[8434];
assign g[24817] = b[13] & g[8434];
assign g[16627] = a[13] & g[8435];
assign g[24818] = b[13] & g[8435];
assign g[16628] = a[13] & g[8436];
assign g[24819] = b[13] & g[8436];
assign g[16629] = a[13] & g[8437];
assign g[24820] = b[13] & g[8437];
assign g[16630] = a[13] & g[8438];
assign g[24821] = b[13] & g[8438];
assign g[16631] = a[13] & g[8439];
assign g[24822] = b[13] & g[8439];
assign g[16632] = a[13] & g[8440];
assign g[24823] = b[13] & g[8440];
assign g[16633] = a[13] & g[8441];
assign g[24824] = b[13] & g[8441];
assign g[16634] = a[13] & g[8442];
assign g[24825] = b[13] & g[8442];
assign g[16635] = a[13] & g[8443];
assign g[24826] = b[13] & g[8443];
assign g[16636] = a[13] & g[8444];
assign g[24827] = b[13] & g[8444];
assign g[16637] = a[13] & g[8445];
assign g[24828] = b[13] & g[8445];
assign g[16638] = a[13] & g[8446];
assign g[24829] = b[13] & g[8446];
assign g[16639] = a[13] & g[8447];
assign g[24830] = b[13] & g[8447];
assign g[16640] = a[13] & g[8448];
assign g[24831] = b[13] & g[8448];
assign g[16641] = a[13] & g[8449];
assign g[24832] = b[13] & g[8449];
assign g[16642] = a[13] & g[8450];
assign g[24833] = b[13] & g[8450];
assign g[16643] = a[13] & g[8451];
assign g[24834] = b[13] & g[8451];
assign g[16644] = a[13] & g[8452];
assign g[24835] = b[13] & g[8452];
assign g[16645] = a[13] & g[8453];
assign g[24836] = b[13] & g[8453];
assign g[16646] = a[13] & g[8454];
assign g[24837] = b[13] & g[8454];
assign g[16647] = a[13] & g[8455];
assign g[24838] = b[13] & g[8455];
assign g[16648] = a[13] & g[8456];
assign g[24839] = b[13] & g[8456];
assign g[16649] = a[13] & g[8457];
assign g[24840] = b[13] & g[8457];
assign g[16650] = a[13] & g[8458];
assign g[24841] = b[13] & g[8458];
assign g[16651] = a[13] & g[8459];
assign g[24842] = b[13] & g[8459];
assign g[16652] = a[13] & g[8460];
assign g[24843] = b[13] & g[8460];
assign g[16653] = a[13] & g[8461];
assign g[24844] = b[13] & g[8461];
assign g[16654] = a[13] & g[8462];
assign g[24845] = b[13] & g[8462];
assign g[16655] = a[13] & g[8463];
assign g[24846] = b[13] & g[8463];
assign g[16656] = a[13] & g[8464];
assign g[24847] = b[13] & g[8464];
assign g[16657] = a[13] & g[8465];
assign g[24848] = b[13] & g[8465];
assign g[16658] = a[13] & g[8466];
assign g[24849] = b[13] & g[8466];
assign g[16659] = a[13] & g[8467];
assign g[24850] = b[13] & g[8467];
assign g[16660] = a[13] & g[8468];
assign g[24851] = b[13] & g[8468];
assign g[16661] = a[13] & g[8469];
assign g[24852] = b[13] & g[8469];
assign g[16662] = a[13] & g[8470];
assign g[24853] = b[13] & g[8470];
assign g[16663] = a[13] & g[8471];
assign g[24854] = b[13] & g[8471];
assign g[16664] = a[13] & g[8472];
assign g[24855] = b[13] & g[8472];
assign g[16665] = a[13] & g[8473];
assign g[24856] = b[13] & g[8473];
assign g[16666] = a[13] & g[8474];
assign g[24857] = b[13] & g[8474];
assign g[16667] = a[13] & g[8475];
assign g[24858] = b[13] & g[8475];
assign g[16668] = a[13] & g[8476];
assign g[24859] = b[13] & g[8476];
assign g[16669] = a[13] & g[8477];
assign g[24860] = b[13] & g[8477];
assign g[16670] = a[13] & g[8478];
assign g[24861] = b[13] & g[8478];
assign g[16671] = a[13] & g[8479];
assign g[24862] = b[13] & g[8479];
assign g[16672] = a[13] & g[8480];
assign g[24863] = b[13] & g[8480];
assign g[16673] = a[13] & g[8481];
assign g[24864] = b[13] & g[8481];
assign g[16674] = a[13] & g[8482];
assign g[24865] = b[13] & g[8482];
assign g[16675] = a[13] & g[8483];
assign g[24866] = b[13] & g[8483];
assign g[16676] = a[13] & g[8484];
assign g[24867] = b[13] & g[8484];
assign g[16677] = a[13] & g[8485];
assign g[24868] = b[13] & g[8485];
assign g[16678] = a[13] & g[8486];
assign g[24869] = b[13] & g[8486];
assign g[16679] = a[13] & g[8487];
assign g[24870] = b[13] & g[8487];
assign g[16680] = a[13] & g[8488];
assign g[24871] = b[13] & g[8488];
assign g[16681] = a[13] & g[8489];
assign g[24872] = b[13] & g[8489];
assign g[16682] = a[13] & g[8490];
assign g[24873] = b[13] & g[8490];
assign g[16683] = a[13] & g[8491];
assign g[24874] = b[13] & g[8491];
assign g[16684] = a[13] & g[8492];
assign g[24875] = b[13] & g[8492];
assign g[16685] = a[13] & g[8493];
assign g[24876] = b[13] & g[8493];
assign g[16686] = a[13] & g[8494];
assign g[24877] = b[13] & g[8494];
assign g[16687] = a[13] & g[8495];
assign g[24878] = b[13] & g[8495];
assign g[16688] = a[13] & g[8496];
assign g[24879] = b[13] & g[8496];
assign g[16689] = a[13] & g[8497];
assign g[24880] = b[13] & g[8497];
assign g[16690] = a[13] & g[8498];
assign g[24881] = b[13] & g[8498];
assign g[16691] = a[13] & g[8499];
assign g[24882] = b[13] & g[8499];
assign g[16692] = a[13] & g[8500];
assign g[24883] = b[13] & g[8500];
assign g[16693] = a[13] & g[8501];
assign g[24884] = b[13] & g[8501];
assign g[16694] = a[13] & g[8502];
assign g[24885] = b[13] & g[8502];
assign g[16695] = a[13] & g[8503];
assign g[24886] = b[13] & g[8503];
assign g[16696] = a[13] & g[8504];
assign g[24887] = b[13] & g[8504];
assign g[16697] = a[13] & g[8505];
assign g[24888] = b[13] & g[8505];
assign g[16698] = a[13] & g[8506];
assign g[24889] = b[13] & g[8506];
assign g[16699] = a[13] & g[8507];
assign g[24890] = b[13] & g[8507];
assign g[16700] = a[13] & g[8508];
assign g[24891] = b[13] & g[8508];
assign g[16701] = a[13] & g[8509];
assign g[24892] = b[13] & g[8509];
assign g[16702] = a[13] & g[8510];
assign g[24893] = b[13] & g[8510];
assign g[16703] = a[13] & g[8511];
assign g[24894] = b[13] & g[8511];
assign g[16704] = a[13] & g[8512];
assign g[24895] = b[13] & g[8512];
assign g[16705] = a[13] & g[8513];
assign g[24896] = b[13] & g[8513];
assign g[16706] = a[13] & g[8514];
assign g[24897] = b[13] & g[8514];
assign g[16707] = a[13] & g[8515];
assign g[24898] = b[13] & g[8515];
assign g[16708] = a[13] & g[8516];
assign g[24899] = b[13] & g[8516];
assign g[16709] = a[13] & g[8517];
assign g[24900] = b[13] & g[8517];
assign g[16710] = a[13] & g[8518];
assign g[24901] = b[13] & g[8518];
assign g[16711] = a[13] & g[8519];
assign g[24902] = b[13] & g[8519];
assign g[16712] = a[13] & g[8520];
assign g[24903] = b[13] & g[8520];
assign g[16713] = a[13] & g[8521];
assign g[24904] = b[13] & g[8521];
assign g[16714] = a[13] & g[8522];
assign g[24905] = b[13] & g[8522];
assign g[16715] = a[13] & g[8523];
assign g[24906] = b[13] & g[8523];
assign g[16716] = a[13] & g[8524];
assign g[24907] = b[13] & g[8524];
assign g[16717] = a[13] & g[8525];
assign g[24908] = b[13] & g[8525];
assign g[16718] = a[13] & g[8526];
assign g[24909] = b[13] & g[8526];
assign g[16719] = a[13] & g[8527];
assign g[24910] = b[13] & g[8527];
assign g[16720] = a[13] & g[8528];
assign g[24911] = b[13] & g[8528];
assign g[16721] = a[13] & g[8529];
assign g[24912] = b[13] & g[8529];
assign g[16722] = a[13] & g[8530];
assign g[24913] = b[13] & g[8530];
assign g[16723] = a[13] & g[8531];
assign g[24914] = b[13] & g[8531];
assign g[16724] = a[13] & g[8532];
assign g[24915] = b[13] & g[8532];
assign g[16725] = a[13] & g[8533];
assign g[24916] = b[13] & g[8533];
assign g[16726] = a[13] & g[8534];
assign g[24917] = b[13] & g[8534];
assign g[16727] = a[13] & g[8535];
assign g[24918] = b[13] & g[8535];
assign g[16728] = a[13] & g[8536];
assign g[24919] = b[13] & g[8536];
assign g[16729] = a[13] & g[8537];
assign g[24920] = b[13] & g[8537];
assign g[16730] = a[13] & g[8538];
assign g[24921] = b[13] & g[8538];
assign g[16731] = a[13] & g[8539];
assign g[24922] = b[13] & g[8539];
assign g[16732] = a[13] & g[8540];
assign g[24923] = b[13] & g[8540];
assign g[16733] = a[13] & g[8541];
assign g[24924] = b[13] & g[8541];
assign g[16734] = a[13] & g[8542];
assign g[24925] = b[13] & g[8542];
assign g[16735] = a[13] & g[8543];
assign g[24926] = b[13] & g[8543];
assign g[16736] = a[13] & g[8544];
assign g[24927] = b[13] & g[8544];
assign g[16737] = a[13] & g[8545];
assign g[24928] = b[13] & g[8545];
assign g[16738] = a[13] & g[8546];
assign g[24929] = b[13] & g[8546];
assign g[16739] = a[13] & g[8547];
assign g[24930] = b[13] & g[8547];
assign g[16740] = a[13] & g[8548];
assign g[24931] = b[13] & g[8548];
assign g[16741] = a[13] & g[8549];
assign g[24932] = b[13] & g[8549];
assign g[16742] = a[13] & g[8550];
assign g[24933] = b[13] & g[8550];
assign g[16743] = a[13] & g[8551];
assign g[24934] = b[13] & g[8551];
assign g[16744] = a[13] & g[8552];
assign g[24935] = b[13] & g[8552];
assign g[16745] = a[13] & g[8553];
assign g[24936] = b[13] & g[8553];
assign g[16746] = a[13] & g[8554];
assign g[24937] = b[13] & g[8554];
assign g[16747] = a[13] & g[8555];
assign g[24938] = b[13] & g[8555];
assign g[16748] = a[13] & g[8556];
assign g[24939] = b[13] & g[8556];
assign g[16749] = a[13] & g[8557];
assign g[24940] = b[13] & g[8557];
assign g[16750] = a[13] & g[8558];
assign g[24941] = b[13] & g[8558];
assign g[16751] = a[13] & g[8559];
assign g[24942] = b[13] & g[8559];
assign g[16752] = a[13] & g[8560];
assign g[24943] = b[13] & g[8560];
assign g[16753] = a[13] & g[8561];
assign g[24944] = b[13] & g[8561];
assign g[16754] = a[13] & g[8562];
assign g[24945] = b[13] & g[8562];
assign g[16755] = a[13] & g[8563];
assign g[24946] = b[13] & g[8563];
assign g[16756] = a[13] & g[8564];
assign g[24947] = b[13] & g[8564];
assign g[16757] = a[13] & g[8565];
assign g[24948] = b[13] & g[8565];
assign g[16758] = a[13] & g[8566];
assign g[24949] = b[13] & g[8566];
assign g[16759] = a[13] & g[8567];
assign g[24950] = b[13] & g[8567];
assign g[16760] = a[13] & g[8568];
assign g[24951] = b[13] & g[8568];
assign g[16761] = a[13] & g[8569];
assign g[24952] = b[13] & g[8569];
assign g[16762] = a[13] & g[8570];
assign g[24953] = b[13] & g[8570];
assign g[16763] = a[13] & g[8571];
assign g[24954] = b[13] & g[8571];
assign g[16764] = a[13] & g[8572];
assign g[24955] = b[13] & g[8572];
assign g[16765] = a[13] & g[8573];
assign g[24956] = b[13] & g[8573];
assign g[16766] = a[13] & g[8574];
assign g[24957] = b[13] & g[8574];
assign g[16767] = a[13] & g[8575];
assign g[24958] = b[13] & g[8575];
assign g[16768] = a[13] & g[8576];
assign g[24959] = b[13] & g[8576];
assign g[16769] = a[13] & g[8577];
assign g[24960] = b[13] & g[8577];
assign g[16770] = a[13] & g[8578];
assign g[24961] = b[13] & g[8578];
assign g[16771] = a[13] & g[8579];
assign g[24962] = b[13] & g[8579];
assign g[16772] = a[13] & g[8580];
assign g[24963] = b[13] & g[8580];
assign g[16773] = a[13] & g[8581];
assign g[24964] = b[13] & g[8581];
assign g[16774] = a[13] & g[8582];
assign g[24965] = b[13] & g[8582];
assign g[16775] = a[13] & g[8583];
assign g[24966] = b[13] & g[8583];
assign g[16776] = a[13] & g[8584];
assign g[24967] = b[13] & g[8584];
assign g[16777] = a[13] & g[8585];
assign g[24968] = b[13] & g[8585];
assign g[16778] = a[13] & g[8586];
assign g[24969] = b[13] & g[8586];
assign g[16779] = a[13] & g[8587];
assign g[24970] = b[13] & g[8587];
assign g[16780] = a[13] & g[8588];
assign g[24971] = b[13] & g[8588];
assign g[16781] = a[13] & g[8589];
assign g[24972] = b[13] & g[8589];
assign g[16782] = a[13] & g[8590];
assign g[24973] = b[13] & g[8590];
assign g[16783] = a[13] & g[8591];
assign g[24974] = b[13] & g[8591];
assign g[16784] = a[13] & g[8592];
assign g[24975] = b[13] & g[8592];
assign g[16785] = a[13] & g[8593];
assign g[24976] = b[13] & g[8593];
assign g[16786] = a[13] & g[8594];
assign g[24977] = b[13] & g[8594];
assign g[16787] = a[13] & g[8595];
assign g[24978] = b[13] & g[8595];
assign g[16788] = a[13] & g[8596];
assign g[24979] = b[13] & g[8596];
assign g[16789] = a[13] & g[8597];
assign g[24980] = b[13] & g[8597];
assign g[16790] = a[13] & g[8598];
assign g[24981] = b[13] & g[8598];
assign g[16791] = a[13] & g[8599];
assign g[24982] = b[13] & g[8599];
assign g[16792] = a[13] & g[8600];
assign g[24983] = b[13] & g[8600];
assign g[16793] = a[13] & g[8601];
assign g[24984] = b[13] & g[8601];
assign g[16794] = a[13] & g[8602];
assign g[24985] = b[13] & g[8602];
assign g[16795] = a[13] & g[8603];
assign g[24986] = b[13] & g[8603];
assign g[16796] = a[13] & g[8604];
assign g[24987] = b[13] & g[8604];
assign g[16797] = a[13] & g[8605];
assign g[24988] = b[13] & g[8605];
assign g[16798] = a[13] & g[8606];
assign g[24989] = b[13] & g[8606];
assign g[16799] = a[13] & g[8607];
assign g[24990] = b[13] & g[8607];
assign g[16800] = a[13] & g[8608];
assign g[24991] = b[13] & g[8608];
assign g[16801] = a[13] & g[8609];
assign g[24992] = b[13] & g[8609];
assign g[16802] = a[13] & g[8610];
assign g[24993] = b[13] & g[8610];
assign g[16803] = a[13] & g[8611];
assign g[24994] = b[13] & g[8611];
assign g[16804] = a[13] & g[8612];
assign g[24995] = b[13] & g[8612];
assign g[16805] = a[13] & g[8613];
assign g[24996] = b[13] & g[8613];
assign g[16806] = a[13] & g[8614];
assign g[24997] = b[13] & g[8614];
assign g[16807] = a[13] & g[8615];
assign g[24998] = b[13] & g[8615];
assign g[16808] = a[13] & g[8616];
assign g[24999] = b[13] & g[8616];
assign g[16809] = a[13] & g[8617];
assign g[25000] = b[13] & g[8617];
assign g[16810] = a[13] & g[8618];
assign g[25001] = b[13] & g[8618];
assign g[16811] = a[13] & g[8619];
assign g[25002] = b[13] & g[8619];
assign g[16812] = a[13] & g[8620];
assign g[25003] = b[13] & g[8620];
assign g[16813] = a[13] & g[8621];
assign g[25004] = b[13] & g[8621];
assign g[16814] = a[13] & g[8622];
assign g[25005] = b[13] & g[8622];
assign g[16815] = a[13] & g[8623];
assign g[25006] = b[13] & g[8623];
assign g[16816] = a[13] & g[8624];
assign g[25007] = b[13] & g[8624];
assign g[16817] = a[13] & g[8625];
assign g[25008] = b[13] & g[8625];
assign g[16818] = a[13] & g[8626];
assign g[25009] = b[13] & g[8626];
assign g[16819] = a[13] & g[8627];
assign g[25010] = b[13] & g[8627];
assign g[16820] = a[13] & g[8628];
assign g[25011] = b[13] & g[8628];
assign g[16821] = a[13] & g[8629];
assign g[25012] = b[13] & g[8629];
assign g[16822] = a[13] & g[8630];
assign g[25013] = b[13] & g[8630];
assign g[16823] = a[13] & g[8631];
assign g[25014] = b[13] & g[8631];
assign g[16824] = a[13] & g[8632];
assign g[25015] = b[13] & g[8632];
assign g[16825] = a[13] & g[8633];
assign g[25016] = b[13] & g[8633];
assign g[16826] = a[13] & g[8634];
assign g[25017] = b[13] & g[8634];
assign g[16827] = a[13] & g[8635];
assign g[25018] = b[13] & g[8635];
assign g[16828] = a[13] & g[8636];
assign g[25019] = b[13] & g[8636];
assign g[16829] = a[13] & g[8637];
assign g[25020] = b[13] & g[8637];
assign g[16830] = a[13] & g[8638];
assign g[25021] = b[13] & g[8638];
assign g[16831] = a[13] & g[8639];
assign g[25022] = b[13] & g[8639];
assign g[16832] = a[13] & g[8640];
assign g[25023] = b[13] & g[8640];
assign g[16833] = a[13] & g[8641];
assign g[25024] = b[13] & g[8641];
assign g[16834] = a[13] & g[8642];
assign g[25025] = b[13] & g[8642];
assign g[16835] = a[13] & g[8643];
assign g[25026] = b[13] & g[8643];
assign g[16836] = a[13] & g[8644];
assign g[25027] = b[13] & g[8644];
assign g[16837] = a[13] & g[8645];
assign g[25028] = b[13] & g[8645];
assign g[16838] = a[13] & g[8646];
assign g[25029] = b[13] & g[8646];
assign g[16839] = a[13] & g[8647];
assign g[25030] = b[13] & g[8647];
assign g[16840] = a[13] & g[8648];
assign g[25031] = b[13] & g[8648];
assign g[16841] = a[13] & g[8649];
assign g[25032] = b[13] & g[8649];
assign g[16842] = a[13] & g[8650];
assign g[25033] = b[13] & g[8650];
assign g[16843] = a[13] & g[8651];
assign g[25034] = b[13] & g[8651];
assign g[16844] = a[13] & g[8652];
assign g[25035] = b[13] & g[8652];
assign g[16845] = a[13] & g[8653];
assign g[25036] = b[13] & g[8653];
assign g[16846] = a[13] & g[8654];
assign g[25037] = b[13] & g[8654];
assign g[16847] = a[13] & g[8655];
assign g[25038] = b[13] & g[8655];
assign g[16848] = a[13] & g[8656];
assign g[25039] = b[13] & g[8656];
assign g[16849] = a[13] & g[8657];
assign g[25040] = b[13] & g[8657];
assign g[16850] = a[13] & g[8658];
assign g[25041] = b[13] & g[8658];
assign g[16851] = a[13] & g[8659];
assign g[25042] = b[13] & g[8659];
assign g[16852] = a[13] & g[8660];
assign g[25043] = b[13] & g[8660];
assign g[16853] = a[13] & g[8661];
assign g[25044] = b[13] & g[8661];
assign g[16854] = a[13] & g[8662];
assign g[25045] = b[13] & g[8662];
assign g[16855] = a[13] & g[8663];
assign g[25046] = b[13] & g[8663];
assign g[16856] = a[13] & g[8664];
assign g[25047] = b[13] & g[8664];
assign g[16857] = a[13] & g[8665];
assign g[25048] = b[13] & g[8665];
assign g[16858] = a[13] & g[8666];
assign g[25049] = b[13] & g[8666];
assign g[16859] = a[13] & g[8667];
assign g[25050] = b[13] & g[8667];
assign g[16860] = a[13] & g[8668];
assign g[25051] = b[13] & g[8668];
assign g[16861] = a[13] & g[8669];
assign g[25052] = b[13] & g[8669];
assign g[16862] = a[13] & g[8670];
assign g[25053] = b[13] & g[8670];
assign g[16863] = a[13] & g[8671];
assign g[25054] = b[13] & g[8671];
assign g[16864] = a[13] & g[8672];
assign g[25055] = b[13] & g[8672];
assign g[16865] = a[13] & g[8673];
assign g[25056] = b[13] & g[8673];
assign g[16866] = a[13] & g[8674];
assign g[25057] = b[13] & g[8674];
assign g[16867] = a[13] & g[8675];
assign g[25058] = b[13] & g[8675];
assign g[16868] = a[13] & g[8676];
assign g[25059] = b[13] & g[8676];
assign g[16869] = a[13] & g[8677];
assign g[25060] = b[13] & g[8677];
assign g[16870] = a[13] & g[8678];
assign g[25061] = b[13] & g[8678];
assign g[16871] = a[13] & g[8679];
assign g[25062] = b[13] & g[8679];
assign g[16872] = a[13] & g[8680];
assign g[25063] = b[13] & g[8680];
assign g[16873] = a[13] & g[8681];
assign g[25064] = b[13] & g[8681];
assign g[16874] = a[13] & g[8682];
assign g[25065] = b[13] & g[8682];
assign g[16875] = a[13] & g[8683];
assign g[25066] = b[13] & g[8683];
assign g[16876] = a[13] & g[8684];
assign g[25067] = b[13] & g[8684];
assign g[16877] = a[13] & g[8685];
assign g[25068] = b[13] & g[8685];
assign g[16878] = a[13] & g[8686];
assign g[25069] = b[13] & g[8686];
assign g[16879] = a[13] & g[8687];
assign g[25070] = b[13] & g[8687];
assign g[16880] = a[13] & g[8688];
assign g[25071] = b[13] & g[8688];
assign g[16881] = a[13] & g[8689];
assign g[25072] = b[13] & g[8689];
assign g[16882] = a[13] & g[8690];
assign g[25073] = b[13] & g[8690];
assign g[16883] = a[13] & g[8691];
assign g[25074] = b[13] & g[8691];
assign g[16884] = a[13] & g[8692];
assign g[25075] = b[13] & g[8692];
assign g[16885] = a[13] & g[8693];
assign g[25076] = b[13] & g[8693];
assign g[16886] = a[13] & g[8694];
assign g[25077] = b[13] & g[8694];
assign g[16887] = a[13] & g[8695];
assign g[25078] = b[13] & g[8695];
assign g[16888] = a[13] & g[8696];
assign g[25079] = b[13] & g[8696];
assign g[16889] = a[13] & g[8697];
assign g[25080] = b[13] & g[8697];
assign g[16890] = a[13] & g[8698];
assign g[25081] = b[13] & g[8698];
assign g[16891] = a[13] & g[8699];
assign g[25082] = b[13] & g[8699];
assign g[16892] = a[13] & g[8700];
assign g[25083] = b[13] & g[8700];
assign g[16893] = a[13] & g[8701];
assign g[25084] = b[13] & g[8701];
assign g[16894] = a[13] & g[8702];
assign g[25085] = b[13] & g[8702];
assign g[16895] = a[13] & g[8703];
assign g[25086] = b[13] & g[8703];
assign g[16896] = a[13] & g[8704];
assign g[25087] = b[13] & g[8704];
assign g[16897] = a[13] & g[8705];
assign g[25088] = b[13] & g[8705];
assign g[16898] = a[13] & g[8706];
assign g[25089] = b[13] & g[8706];
assign g[16899] = a[13] & g[8707];
assign g[25090] = b[13] & g[8707];
assign g[16900] = a[13] & g[8708];
assign g[25091] = b[13] & g[8708];
assign g[16901] = a[13] & g[8709];
assign g[25092] = b[13] & g[8709];
assign g[16902] = a[13] & g[8710];
assign g[25093] = b[13] & g[8710];
assign g[16903] = a[13] & g[8711];
assign g[25094] = b[13] & g[8711];
assign g[16904] = a[13] & g[8712];
assign g[25095] = b[13] & g[8712];
assign g[16905] = a[13] & g[8713];
assign g[25096] = b[13] & g[8713];
assign g[16906] = a[13] & g[8714];
assign g[25097] = b[13] & g[8714];
assign g[16907] = a[13] & g[8715];
assign g[25098] = b[13] & g[8715];
assign g[16908] = a[13] & g[8716];
assign g[25099] = b[13] & g[8716];
assign g[16909] = a[13] & g[8717];
assign g[25100] = b[13] & g[8717];
assign g[16910] = a[13] & g[8718];
assign g[25101] = b[13] & g[8718];
assign g[16911] = a[13] & g[8719];
assign g[25102] = b[13] & g[8719];
assign g[16912] = a[13] & g[8720];
assign g[25103] = b[13] & g[8720];
assign g[16913] = a[13] & g[8721];
assign g[25104] = b[13] & g[8721];
assign g[16914] = a[13] & g[8722];
assign g[25105] = b[13] & g[8722];
assign g[16915] = a[13] & g[8723];
assign g[25106] = b[13] & g[8723];
assign g[16916] = a[13] & g[8724];
assign g[25107] = b[13] & g[8724];
assign g[16917] = a[13] & g[8725];
assign g[25108] = b[13] & g[8725];
assign g[16918] = a[13] & g[8726];
assign g[25109] = b[13] & g[8726];
assign g[16919] = a[13] & g[8727];
assign g[25110] = b[13] & g[8727];
assign g[16920] = a[13] & g[8728];
assign g[25111] = b[13] & g[8728];
assign g[16921] = a[13] & g[8729];
assign g[25112] = b[13] & g[8729];
assign g[16922] = a[13] & g[8730];
assign g[25113] = b[13] & g[8730];
assign g[16923] = a[13] & g[8731];
assign g[25114] = b[13] & g[8731];
assign g[16924] = a[13] & g[8732];
assign g[25115] = b[13] & g[8732];
assign g[16925] = a[13] & g[8733];
assign g[25116] = b[13] & g[8733];
assign g[16926] = a[13] & g[8734];
assign g[25117] = b[13] & g[8734];
assign g[16927] = a[13] & g[8735];
assign g[25118] = b[13] & g[8735];
assign g[16928] = a[13] & g[8736];
assign g[25119] = b[13] & g[8736];
assign g[16929] = a[13] & g[8737];
assign g[25120] = b[13] & g[8737];
assign g[16930] = a[13] & g[8738];
assign g[25121] = b[13] & g[8738];
assign g[16931] = a[13] & g[8739];
assign g[25122] = b[13] & g[8739];
assign g[16932] = a[13] & g[8740];
assign g[25123] = b[13] & g[8740];
assign g[16933] = a[13] & g[8741];
assign g[25124] = b[13] & g[8741];
assign g[16934] = a[13] & g[8742];
assign g[25125] = b[13] & g[8742];
assign g[16935] = a[13] & g[8743];
assign g[25126] = b[13] & g[8743];
assign g[16936] = a[13] & g[8744];
assign g[25127] = b[13] & g[8744];
assign g[16937] = a[13] & g[8745];
assign g[25128] = b[13] & g[8745];
assign g[16938] = a[13] & g[8746];
assign g[25129] = b[13] & g[8746];
assign g[16939] = a[13] & g[8747];
assign g[25130] = b[13] & g[8747];
assign g[16940] = a[13] & g[8748];
assign g[25131] = b[13] & g[8748];
assign g[16941] = a[13] & g[8749];
assign g[25132] = b[13] & g[8749];
assign g[16942] = a[13] & g[8750];
assign g[25133] = b[13] & g[8750];
assign g[16943] = a[13] & g[8751];
assign g[25134] = b[13] & g[8751];
assign g[16944] = a[13] & g[8752];
assign g[25135] = b[13] & g[8752];
assign g[16945] = a[13] & g[8753];
assign g[25136] = b[13] & g[8753];
assign g[16946] = a[13] & g[8754];
assign g[25137] = b[13] & g[8754];
assign g[16947] = a[13] & g[8755];
assign g[25138] = b[13] & g[8755];
assign g[16948] = a[13] & g[8756];
assign g[25139] = b[13] & g[8756];
assign g[16949] = a[13] & g[8757];
assign g[25140] = b[13] & g[8757];
assign g[16950] = a[13] & g[8758];
assign g[25141] = b[13] & g[8758];
assign g[16951] = a[13] & g[8759];
assign g[25142] = b[13] & g[8759];
assign g[16952] = a[13] & g[8760];
assign g[25143] = b[13] & g[8760];
assign g[16953] = a[13] & g[8761];
assign g[25144] = b[13] & g[8761];
assign g[16954] = a[13] & g[8762];
assign g[25145] = b[13] & g[8762];
assign g[16955] = a[13] & g[8763];
assign g[25146] = b[13] & g[8763];
assign g[16956] = a[13] & g[8764];
assign g[25147] = b[13] & g[8764];
assign g[16957] = a[13] & g[8765];
assign g[25148] = b[13] & g[8765];
assign g[16958] = a[13] & g[8766];
assign g[25149] = b[13] & g[8766];
assign g[16959] = a[13] & g[8767];
assign g[25150] = b[13] & g[8767];
assign g[16960] = a[13] & g[8768];
assign g[25151] = b[13] & g[8768];
assign g[16961] = a[13] & g[8769];
assign g[25152] = b[13] & g[8769];
assign g[16962] = a[13] & g[8770];
assign g[25153] = b[13] & g[8770];
assign g[16963] = a[13] & g[8771];
assign g[25154] = b[13] & g[8771];
assign g[16964] = a[13] & g[8772];
assign g[25155] = b[13] & g[8772];
assign g[16965] = a[13] & g[8773];
assign g[25156] = b[13] & g[8773];
assign g[16966] = a[13] & g[8774];
assign g[25157] = b[13] & g[8774];
assign g[16967] = a[13] & g[8775];
assign g[25158] = b[13] & g[8775];
assign g[16968] = a[13] & g[8776];
assign g[25159] = b[13] & g[8776];
assign g[16969] = a[13] & g[8777];
assign g[25160] = b[13] & g[8777];
assign g[16970] = a[13] & g[8778];
assign g[25161] = b[13] & g[8778];
assign g[16971] = a[13] & g[8779];
assign g[25162] = b[13] & g[8779];
assign g[16972] = a[13] & g[8780];
assign g[25163] = b[13] & g[8780];
assign g[16973] = a[13] & g[8781];
assign g[25164] = b[13] & g[8781];
assign g[16974] = a[13] & g[8782];
assign g[25165] = b[13] & g[8782];
assign g[16975] = a[13] & g[8783];
assign g[25166] = b[13] & g[8783];
assign g[16976] = a[13] & g[8784];
assign g[25167] = b[13] & g[8784];
assign g[16977] = a[13] & g[8785];
assign g[25168] = b[13] & g[8785];
assign g[16978] = a[13] & g[8786];
assign g[25169] = b[13] & g[8786];
assign g[16979] = a[13] & g[8787];
assign g[25170] = b[13] & g[8787];
assign g[16980] = a[13] & g[8788];
assign g[25171] = b[13] & g[8788];
assign g[16981] = a[13] & g[8789];
assign g[25172] = b[13] & g[8789];
assign g[16982] = a[13] & g[8790];
assign g[25173] = b[13] & g[8790];
assign g[16983] = a[13] & g[8791];
assign g[25174] = b[13] & g[8791];
assign g[16984] = a[13] & g[8792];
assign g[25175] = b[13] & g[8792];
assign g[16985] = a[13] & g[8793];
assign g[25176] = b[13] & g[8793];
assign g[16986] = a[13] & g[8794];
assign g[25177] = b[13] & g[8794];
assign g[16987] = a[13] & g[8795];
assign g[25178] = b[13] & g[8795];
assign g[16988] = a[13] & g[8796];
assign g[25179] = b[13] & g[8796];
assign g[16989] = a[13] & g[8797];
assign g[25180] = b[13] & g[8797];
assign g[16990] = a[13] & g[8798];
assign g[25181] = b[13] & g[8798];
assign g[16991] = a[13] & g[8799];
assign g[25182] = b[13] & g[8799];
assign g[16992] = a[13] & g[8800];
assign g[25183] = b[13] & g[8800];
assign g[16993] = a[13] & g[8801];
assign g[25184] = b[13] & g[8801];
assign g[16994] = a[13] & g[8802];
assign g[25185] = b[13] & g[8802];
assign g[16995] = a[13] & g[8803];
assign g[25186] = b[13] & g[8803];
assign g[16996] = a[13] & g[8804];
assign g[25187] = b[13] & g[8804];
assign g[16997] = a[13] & g[8805];
assign g[25188] = b[13] & g[8805];
assign g[16998] = a[13] & g[8806];
assign g[25189] = b[13] & g[8806];
assign g[16999] = a[13] & g[8807];
assign g[25190] = b[13] & g[8807];
assign g[17000] = a[13] & g[8808];
assign g[25191] = b[13] & g[8808];
assign g[17001] = a[13] & g[8809];
assign g[25192] = b[13] & g[8809];
assign g[17002] = a[13] & g[8810];
assign g[25193] = b[13] & g[8810];
assign g[17003] = a[13] & g[8811];
assign g[25194] = b[13] & g[8811];
assign g[17004] = a[13] & g[8812];
assign g[25195] = b[13] & g[8812];
assign g[17005] = a[13] & g[8813];
assign g[25196] = b[13] & g[8813];
assign g[17006] = a[13] & g[8814];
assign g[25197] = b[13] & g[8814];
assign g[17007] = a[13] & g[8815];
assign g[25198] = b[13] & g[8815];
assign g[17008] = a[13] & g[8816];
assign g[25199] = b[13] & g[8816];
assign g[17009] = a[13] & g[8817];
assign g[25200] = b[13] & g[8817];
assign g[17010] = a[13] & g[8818];
assign g[25201] = b[13] & g[8818];
assign g[17011] = a[13] & g[8819];
assign g[25202] = b[13] & g[8819];
assign g[17012] = a[13] & g[8820];
assign g[25203] = b[13] & g[8820];
assign g[17013] = a[13] & g[8821];
assign g[25204] = b[13] & g[8821];
assign g[17014] = a[13] & g[8822];
assign g[25205] = b[13] & g[8822];
assign g[17015] = a[13] & g[8823];
assign g[25206] = b[13] & g[8823];
assign g[17016] = a[13] & g[8824];
assign g[25207] = b[13] & g[8824];
assign g[17017] = a[13] & g[8825];
assign g[25208] = b[13] & g[8825];
assign g[17018] = a[13] & g[8826];
assign g[25209] = b[13] & g[8826];
assign g[17019] = a[13] & g[8827];
assign g[25210] = b[13] & g[8827];
assign g[17020] = a[13] & g[8828];
assign g[25211] = b[13] & g[8828];
assign g[17021] = a[13] & g[8829];
assign g[25212] = b[13] & g[8829];
assign g[17022] = a[13] & g[8830];
assign g[25213] = b[13] & g[8830];
assign g[17023] = a[13] & g[8831];
assign g[25214] = b[13] & g[8831];
assign g[17024] = a[13] & g[8832];
assign g[25215] = b[13] & g[8832];
assign g[17025] = a[13] & g[8833];
assign g[25216] = b[13] & g[8833];
assign g[17026] = a[13] & g[8834];
assign g[25217] = b[13] & g[8834];
assign g[17027] = a[13] & g[8835];
assign g[25218] = b[13] & g[8835];
assign g[17028] = a[13] & g[8836];
assign g[25219] = b[13] & g[8836];
assign g[17029] = a[13] & g[8837];
assign g[25220] = b[13] & g[8837];
assign g[17030] = a[13] & g[8838];
assign g[25221] = b[13] & g[8838];
assign g[17031] = a[13] & g[8839];
assign g[25222] = b[13] & g[8839];
assign g[17032] = a[13] & g[8840];
assign g[25223] = b[13] & g[8840];
assign g[17033] = a[13] & g[8841];
assign g[25224] = b[13] & g[8841];
assign g[17034] = a[13] & g[8842];
assign g[25225] = b[13] & g[8842];
assign g[17035] = a[13] & g[8843];
assign g[25226] = b[13] & g[8843];
assign g[17036] = a[13] & g[8844];
assign g[25227] = b[13] & g[8844];
assign g[17037] = a[13] & g[8845];
assign g[25228] = b[13] & g[8845];
assign g[17038] = a[13] & g[8846];
assign g[25229] = b[13] & g[8846];
assign g[17039] = a[13] & g[8847];
assign g[25230] = b[13] & g[8847];
assign g[17040] = a[13] & g[8848];
assign g[25231] = b[13] & g[8848];
assign g[17041] = a[13] & g[8849];
assign g[25232] = b[13] & g[8849];
assign g[17042] = a[13] & g[8850];
assign g[25233] = b[13] & g[8850];
assign g[17043] = a[13] & g[8851];
assign g[25234] = b[13] & g[8851];
assign g[17044] = a[13] & g[8852];
assign g[25235] = b[13] & g[8852];
assign g[17045] = a[13] & g[8853];
assign g[25236] = b[13] & g[8853];
assign g[17046] = a[13] & g[8854];
assign g[25237] = b[13] & g[8854];
assign g[17047] = a[13] & g[8855];
assign g[25238] = b[13] & g[8855];
assign g[17048] = a[13] & g[8856];
assign g[25239] = b[13] & g[8856];
assign g[17049] = a[13] & g[8857];
assign g[25240] = b[13] & g[8857];
assign g[17050] = a[13] & g[8858];
assign g[25241] = b[13] & g[8858];
assign g[17051] = a[13] & g[8859];
assign g[25242] = b[13] & g[8859];
assign g[17052] = a[13] & g[8860];
assign g[25243] = b[13] & g[8860];
assign g[17053] = a[13] & g[8861];
assign g[25244] = b[13] & g[8861];
assign g[17054] = a[13] & g[8862];
assign g[25245] = b[13] & g[8862];
assign g[17055] = a[13] & g[8863];
assign g[25246] = b[13] & g[8863];
assign g[17056] = a[13] & g[8864];
assign g[25247] = b[13] & g[8864];
assign g[17057] = a[13] & g[8865];
assign g[25248] = b[13] & g[8865];
assign g[17058] = a[13] & g[8866];
assign g[25249] = b[13] & g[8866];
assign g[17059] = a[13] & g[8867];
assign g[25250] = b[13] & g[8867];
assign g[17060] = a[13] & g[8868];
assign g[25251] = b[13] & g[8868];
assign g[17061] = a[13] & g[8869];
assign g[25252] = b[13] & g[8869];
assign g[17062] = a[13] & g[8870];
assign g[25253] = b[13] & g[8870];
assign g[17063] = a[13] & g[8871];
assign g[25254] = b[13] & g[8871];
assign g[17064] = a[13] & g[8872];
assign g[25255] = b[13] & g[8872];
assign g[17065] = a[13] & g[8873];
assign g[25256] = b[13] & g[8873];
assign g[17066] = a[13] & g[8874];
assign g[25257] = b[13] & g[8874];
assign g[17067] = a[13] & g[8875];
assign g[25258] = b[13] & g[8875];
assign g[17068] = a[13] & g[8876];
assign g[25259] = b[13] & g[8876];
assign g[17069] = a[13] & g[8877];
assign g[25260] = b[13] & g[8877];
assign g[17070] = a[13] & g[8878];
assign g[25261] = b[13] & g[8878];
assign g[17071] = a[13] & g[8879];
assign g[25262] = b[13] & g[8879];
assign g[17072] = a[13] & g[8880];
assign g[25263] = b[13] & g[8880];
assign g[17073] = a[13] & g[8881];
assign g[25264] = b[13] & g[8881];
assign g[17074] = a[13] & g[8882];
assign g[25265] = b[13] & g[8882];
assign g[17075] = a[13] & g[8883];
assign g[25266] = b[13] & g[8883];
assign g[17076] = a[13] & g[8884];
assign g[25267] = b[13] & g[8884];
assign g[17077] = a[13] & g[8885];
assign g[25268] = b[13] & g[8885];
assign g[17078] = a[13] & g[8886];
assign g[25269] = b[13] & g[8886];
assign g[17079] = a[13] & g[8887];
assign g[25270] = b[13] & g[8887];
assign g[17080] = a[13] & g[8888];
assign g[25271] = b[13] & g[8888];
assign g[17081] = a[13] & g[8889];
assign g[25272] = b[13] & g[8889];
assign g[17082] = a[13] & g[8890];
assign g[25273] = b[13] & g[8890];
assign g[17083] = a[13] & g[8891];
assign g[25274] = b[13] & g[8891];
assign g[17084] = a[13] & g[8892];
assign g[25275] = b[13] & g[8892];
assign g[17085] = a[13] & g[8893];
assign g[25276] = b[13] & g[8893];
assign g[17086] = a[13] & g[8894];
assign g[25277] = b[13] & g[8894];
assign g[17087] = a[13] & g[8895];
assign g[25278] = b[13] & g[8895];
assign g[17088] = a[13] & g[8896];
assign g[25279] = b[13] & g[8896];
assign g[17089] = a[13] & g[8897];
assign g[25280] = b[13] & g[8897];
assign g[17090] = a[13] & g[8898];
assign g[25281] = b[13] & g[8898];
assign g[17091] = a[13] & g[8899];
assign g[25282] = b[13] & g[8899];
assign g[17092] = a[13] & g[8900];
assign g[25283] = b[13] & g[8900];
assign g[17093] = a[13] & g[8901];
assign g[25284] = b[13] & g[8901];
assign g[17094] = a[13] & g[8902];
assign g[25285] = b[13] & g[8902];
assign g[17095] = a[13] & g[8903];
assign g[25286] = b[13] & g[8903];
assign g[17096] = a[13] & g[8904];
assign g[25287] = b[13] & g[8904];
assign g[17097] = a[13] & g[8905];
assign g[25288] = b[13] & g[8905];
assign g[17098] = a[13] & g[8906];
assign g[25289] = b[13] & g[8906];
assign g[17099] = a[13] & g[8907];
assign g[25290] = b[13] & g[8907];
assign g[17100] = a[13] & g[8908];
assign g[25291] = b[13] & g[8908];
assign g[17101] = a[13] & g[8909];
assign g[25292] = b[13] & g[8909];
assign g[17102] = a[13] & g[8910];
assign g[25293] = b[13] & g[8910];
assign g[17103] = a[13] & g[8911];
assign g[25294] = b[13] & g[8911];
assign g[17104] = a[13] & g[8912];
assign g[25295] = b[13] & g[8912];
assign g[17105] = a[13] & g[8913];
assign g[25296] = b[13] & g[8913];
assign g[17106] = a[13] & g[8914];
assign g[25297] = b[13] & g[8914];
assign g[17107] = a[13] & g[8915];
assign g[25298] = b[13] & g[8915];
assign g[17108] = a[13] & g[8916];
assign g[25299] = b[13] & g[8916];
assign g[17109] = a[13] & g[8917];
assign g[25300] = b[13] & g[8917];
assign g[17110] = a[13] & g[8918];
assign g[25301] = b[13] & g[8918];
assign g[17111] = a[13] & g[8919];
assign g[25302] = b[13] & g[8919];
assign g[17112] = a[13] & g[8920];
assign g[25303] = b[13] & g[8920];
assign g[17113] = a[13] & g[8921];
assign g[25304] = b[13] & g[8921];
assign g[17114] = a[13] & g[8922];
assign g[25305] = b[13] & g[8922];
assign g[17115] = a[13] & g[8923];
assign g[25306] = b[13] & g[8923];
assign g[17116] = a[13] & g[8924];
assign g[25307] = b[13] & g[8924];
assign g[17117] = a[13] & g[8925];
assign g[25308] = b[13] & g[8925];
assign g[17118] = a[13] & g[8926];
assign g[25309] = b[13] & g[8926];
assign g[17119] = a[13] & g[8927];
assign g[25310] = b[13] & g[8927];
assign g[17120] = a[13] & g[8928];
assign g[25311] = b[13] & g[8928];
assign g[17121] = a[13] & g[8929];
assign g[25312] = b[13] & g[8929];
assign g[17122] = a[13] & g[8930];
assign g[25313] = b[13] & g[8930];
assign g[17123] = a[13] & g[8931];
assign g[25314] = b[13] & g[8931];
assign g[17124] = a[13] & g[8932];
assign g[25315] = b[13] & g[8932];
assign g[17125] = a[13] & g[8933];
assign g[25316] = b[13] & g[8933];
assign g[17126] = a[13] & g[8934];
assign g[25317] = b[13] & g[8934];
assign g[17127] = a[13] & g[8935];
assign g[25318] = b[13] & g[8935];
assign g[17128] = a[13] & g[8936];
assign g[25319] = b[13] & g[8936];
assign g[17129] = a[13] & g[8937];
assign g[25320] = b[13] & g[8937];
assign g[17130] = a[13] & g[8938];
assign g[25321] = b[13] & g[8938];
assign g[17131] = a[13] & g[8939];
assign g[25322] = b[13] & g[8939];
assign g[17132] = a[13] & g[8940];
assign g[25323] = b[13] & g[8940];
assign g[17133] = a[13] & g[8941];
assign g[25324] = b[13] & g[8941];
assign g[17134] = a[13] & g[8942];
assign g[25325] = b[13] & g[8942];
assign g[17135] = a[13] & g[8943];
assign g[25326] = b[13] & g[8943];
assign g[17136] = a[13] & g[8944];
assign g[25327] = b[13] & g[8944];
assign g[17137] = a[13] & g[8945];
assign g[25328] = b[13] & g[8945];
assign g[17138] = a[13] & g[8946];
assign g[25329] = b[13] & g[8946];
assign g[17139] = a[13] & g[8947];
assign g[25330] = b[13] & g[8947];
assign g[17140] = a[13] & g[8948];
assign g[25331] = b[13] & g[8948];
assign g[17141] = a[13] & g[8949];
assign g[25332] = b[13] & g[8949];
assign g[17142] = a[13] & g[8950];
assign g[25333] = b[13] & g[8950];
assign g[17143] = a[13] & g[8951];
assign g[25334] = b[13] & g[8951];
assign g[17144] = a[13] & g[8952];
assign g[25335] = b[13] & g[8952];
assign g[17145] = a[13] & g[8953];
assign g[25336] = b[13] & g[8953];
assign g[17146] = a[13] & g[8954];
assign g[25337] = b[13] & g[8954];
assign g[17147] = a[13] & g[8955];
assign g[25338] = b[13] & g[8955];
assign g[17148] = a[13] & g[8956];
assign g[25339] = b[13] & g[8956];
assign g[17149] = a[13] & g[8957];
assign g[25340] = b[13] & g[8957];
assign g[17150] = a[13] & g[8958];
assign g[25341] = b[13] & g[8958];
assign g[17151] = a[13] & g[8959];
assign g[25342] = b[13] & g[8959];
assign g[17152] = a[13] & g[8960];
assign g[25343] = b[13] & g[8960];
assign g[17153] = a[13] & g[8961];
assign g[25344] = b[13] & g[8961];
assign g[17154] = a[13] & g[8962];
assign g[25345] = b[13] & g[8962];
assign g[17155] = a[13] & g[8963];
assign g[25346] = b[13] & g[8963];
assign g[17156] = a[13] & g[8964];
assign g[25347] = b[13] & g[8964];
assign g[17157] = a[13] & g[8965];
assign g[25348] = b[13] & g[8965];
assign g[17158] = a[13] & g[8966];
assign g[25349] = b[13] & g[8966];
assign g[17159] = a[13] & g[8967];
assign g[25350] = b[13] & g[8967];
assign g[17160] = a[13] & g[8968];
assign g[25351] = b[13] & g[8968];
assign g[17161] = a[13] & g[8969];
assign g[25352] = b[13] & g[8969];
assign g[17162] = a[13] & g[8970];
assign g[25353] = b[13] & g[8970];
assign g[17163] = a[13] & g[8971];
assign g[25354] = b[13] & g[8971];
assign g[17164] = a[13] & g[8972];
assign g[25355] = b[13] & g[8972];
assign g[17165] = a[13] & g[8973];
assign g[25356] = b[13] & g[8973];
assign g[17166] = a[13] & g[8974];
assign g[25357] = b[13] & g[8974];
assign g[17167] = a[13] & g[8975];
assign g[25358] = b[13] & g[8975];
assign g[17168] = a[13] & g[8976];
assign g[25359] = b[13] & g[8976];
assign g[17169] = a[13] & g[8977];
assign g[25360] = b[13] & g[8977];
assign g[17170] = a[13] & g[8978];
assign g[25361] = b[13] & g[8978];
assign g[17171] = a[13] & g[8979];
assign g[25362] = b[13] & g[8979];
assign g[17172] = a[13] & g[8980];
assign g[25363] = b[13] & g[8980];
assign g[17173] = a[13] & g[8981];
assign g[25364] = b[13] & g[8981];
assign g[17174] = a[13] & g[8982];
assign g[25365] = b[13] & g[8982];
assign g[17175] = a[13] & g[8983];
assign g[25366] = b[13] & g[8983];
assign g[17176] = a[13] & g[8984];
assign g[25367] = b[13] & g[8984];
assign g[17177] = a[13] & g[8985];
assign g[25368] = b[13] & g[8985];
assign g[17178] = a[13] & g[8986];
assign g[25369] = b[13] & g[8986];
assign g[17179] = a[13] & g[8987];
assign g[25370] = b[13] & g[8987];
assign g[17180] = a[13] & g[8988];
assign g[25371] = b[13] & g[8988];
assign g[17181] = a[13] & g[8989];
assign g[25372] = b[13] & g[8989];
assign g[17182] = a[13] & g[8990];
assign g[25373] = b[13] & g[8990];
assign g[17183] = a[13] & g[8991];
assign g[25374] = b[13] & g[8991];
assign g[17184] = a[13] & g[8992];
assign g[25375] = b[13] & g[8992];
assign g[17185] = a[13] & g[8993];
assign g[25376] = b[13] & g[8993];
assign g[17186] = a[13] & g[8994];
assign g[25377] = b[13] & g[8994];
assign g[17187] = a[13] & g[8995];
assign g[25378] = b[13] & g[8995];
assign g[17188] = a[13] & g[8996];
assign g[25379] = b[13] & g[8996];
assign g[17189] = a[13] & g[8997];
assign g[25380] = b[13] & g[8997];
assign g[17190] = a[13] & g[8998];
assign g[25381] = b[13] & g[8998];
assign g[17191] = a[13] & g[8999];
assign g[25382] = b[13] & g[8999];
assign g[17192] = a[13] & g[9000];
assign g[25383] = b[13] & g[9000];
assign g[17193] = a[13] & g[9001];
assign g[25384] = b[13] & g[9001];
assign g[17194] = a[13] & g[9002];
assign g[25385] = b[13] & g[9002];
assign g[17195] = a[13] & g[9003];
assign g[25386] = b[13] & g[9003];
assign g[17196] = a[13] & g[9004];
assign g[25387] = b[13] & g[9004];
assign g[17197] = a[13] & g[9005];
assign g[25388] = b[13] & g[9005];
assign g[17198] = a[13] & g[9006];
assign g[25389] = b[13] & g[9006];
assign g[17199] = a[13] & g[9007];
assign g[25390] = b[13] & g[9007];
assign g[17200] = a[13] & g[9008];
assign g[25391] = b[13] & g[9008];
assign g[17201] = a[13] & g[9009];
assign g[25392] = b[13] & g[9009];
assign g[17202] = a[13] & g[9010];
assign g[25393] = b[13] & g[9010];
assign g[17203] = a[13] & g[9011];
assign g[25394] = b[13] & g[9011];
assign g[17204] = a[13] & g[9012];
assign g[25395] = b[13] & g[9012];
assign g[17205] = a[13] & g[9013];
assign g[25396] = b[13] & g[9013];
assign g[17206] = a[13] & g[9014];
assign g[25397] = b[13] & g[9014];
assign g[17207] = a[13] & g[9015];
assign g[25398] = b[13] & g[9015];
assign g[17208] = a[13] & g[9016];
assign g[25399] = b[13] & g[9016];
assign g[17209] = a[13] & g[9017];
assign g[25400] = b[13] & g[9017];
assign g[17210] = a[13] & g[9018];
assign g[25401] = b[13] & g[9018];
assign g[17211] = a[13] & g[9019];
assign g[25402] = b[13] & g[9019];
assign g[17212] = a[13] & g[9020];
assign g[25403] = b[13] & g[9020];
assign g[17213] = a[13] & g[9021];
assign g[25404] = b[13] & g[9021];
assign g[17214] = a[13] & g[9022];
assign g[25405] = b[13] & g[9022];
assign g[17215] = a[13] & g[9023];
assign g[25406] = b[13] & g[9023];
assign g[17216] = a[13] & g[9024];
assign g[25407] = b[13] & g[9024];
assign g[17217] = a[13] & g[9025];
assign g[25408] = b[13] & g[9025];
assign g[17218] = a[13] & g[9026];
assign g[25409] = b[13] & g[9026];
assign g[17219] = a[13] & g[9027];
assign g[25410] = b[13] & g[9027];
assign g[17220] = a[13] & g[9028];
assign g[25411] = b[13] & g[9028];
assign g[17221] = a[13] & g[9029];
assign g[25412] = b[13] & g[9029];
assign g[17222] = a[13] & g[9030];
assign g[25413] = b[13] & g[9030];
assign g[17223] = a[13] & g[9031];
assign g[25414] = b[13] & g[9031];
assign g[17224] = a[13] & g[9032];
assign g[25415] = b[13] & g[9032];
assign g[17225] = a[13] & g[9033];
assign g[25416] = b[13] & g[9033];
assign g[17226] = a[13] & g[9034];
assign g[25417] = b[13] & g[9034];
assign g[17227] = a[13] & g[9035];
assign g[25418] = b[13] & g[9035];
assign g[17228] = a[13] & g[9036];
assign g[25419] = b[13] & g[9036];
assign g[17229] = a[13] & g[9037];
assign g[25420] = b[13] & g[9037];
assign g[17230] = a[13] & g[9038];
assign g[25421] = b[13] & g[9038];
assign g[17231] = a[13] & g[9039];
assign g[25422] = b[13] & g[9039];
assign g[17232] = a[13] & g[9040];
assign g[25423] = b[13] & g[9040];
assign g[17233] = a[13] & g[9041];
assign g[25424] = b[13] & g[9041];
assign g[17234] = a[13] & g[9042];
assign g[25425] = b[13] & g[9042];
assign g[17235] = a[13] & g[9043];
assign g[25426] = b[13] & g[9043];
assign g[17236] = a[13] & g[9044];
assign g[25427] = b[13] & g[9044];
assign g[17237] = a[13] & g[9045];
assign g[25428] = b[13] & g[9045];
assign g[17238] = a[13] & g[9046];
assign g[25429] = b[13] & g[9046];
assign g[17239] = a[13] & g[9047];
assign g[25430] = b[13] & g[9047];
assign g[17240] = a[13] & g[9048];
assign g[25431] = b[13] & g[9048];
assign g[17241] = a[13] & g[9049];
assign g[25432] = b[13] & g[9049];
assign g[17242] = a[13] & g[9050];
assign g[25433] = b[13] & g[9050];
assign g[17243] = a[13] & g[9051];
assign g[25434] = b[13] & g[9051];
assign g[17244] = a[13] & g[9052];
assign g[25435] = b[13] & g[9052];
assign g[17245] = a[13] & g[9053];
assign g[25436] = b[13] & g[9053];
assign g[17246] = a[13] & g[9054];
assign g[25437] = b[13] & g[9054];
assign g[17247] = a[13] & g[9055];
assign g[25438] = b[13] & g[9055];
assign g[17248] = a[13] & g[9056];
assign g[25439] = b[13] & g[9056];
assign g[17249] = a[13] & g[9057];
assign g[25440] = b[13] & g[9057];
assign g[17250] = a[13] & g[9058];
assign g[25441] = b[13] & g[9058];
assign g[17251] = a[13] & g[9059];
assign g[25442] = b[13] & g[9059];
assign g[17252] = a[13] & g[9060];
assign g[25443] = b[13] & g[9060];
assign g[17253] = a[13] & g[9061];
assign g[25444] = b[13] & g[9061];
assign g[17254] = a[13] & g[9062];
assign g[25445] = b[13] & g[9062];
assign g[17255] = a[13] & g[9063];
assign g[25446] = b[13] & g[9063];
assign g[17256] = a[13] & g[9064];
assign g[25447] = b[13] & g[9064];
assign g[17257] = a[13] & g[9065];
assign g[25448] = b[13] & g[9065];
assign g[17258] = a[13] & g[9066];
assign g[25449] = b[13] & g[9066];
assign g[17259] = a[13] & g[9067];
assign g[25450] = b[13] & g[9067];
assign g[17260] = a[13] & g[9068];
assign g[25451] = b[13] & g[9068];
assign g[17261] = a[13] & g[9069];
assign g[25452] = b[13] & g[9069];
assign g[17262] = a[13] & g[9070];
assign g[25453] = b[13] & g[9070];
assign g[17263] = a[13] & g[9071];
assign g[25454] = b[13] & g[9071];
assign g[17264] = a[13] & g[9072];
assign g[25455] = b[13] & g[9072];
assign g[17265] = a[13] & g[9073];
assign g[25456] = b[13] & g[9073];
assign g[17266] = a[13] & g[9074];
assign g[25457] = b[13] & g[9074];
assign g[17267] = a[13] & g[9075];
assign g[25458] = b[13] & g[9075];
assign g[17268] = a[13] & g[9076];
assign g[25459] = b[13] & g[9076];
assign g[17269] = a[13] & g[9077];
assign g[25460] = b[13] & g[9077];
assign g[17270] = a[13] & g[9078];
assign g[25461] = b[13] & g[9078];
assign g[17271] = a[13] & g[9079];
assign g[25462] = b[13] & g[9079];
assign g[17272] = a[13] & g[9080];
assign g[25463] = b[13] & g[9080];
assign g[17273] = a[13] & g[9081];
assign g[25464] = b[13] & g[9081];
assign g[17274] = a[13] & g[9082];
assign g[25465] = b[13] & g[9082];
assign g[17275] = a[13] & g[9083];
assign g[25466] = b[13] & g[9083];
assign g[17276] = a[13] & g[9084];
assign g[25467] = b[13] & g[9084];
assign g[17277] = a[13] & g[9085];
assign g[25468] = b[13] & g[9085];
assign g[17278] = a[13] & g[9086];
assign g[25469] = b[13] & g[9086];
assign g[17279] = a[13] & g[9087];
assign g[25470] = b[13] & g[9087];
assign g[17280] = a[13] & g[9088];
assign g[25471] = b[13] & g[9088];
assign g[17281] = a[13] & g[9089];
assign g[25472] = b[13] & g[9089];
assign g[17282] = a[13] & g[9090];
assign g[25473] = b[13] & g[9090];
assign g[17283] = a[13] & g[9091];
assign g[25474] = b[13] & g[9091];
assign g[17284] = a[13] & g[9092];
assign g[25475] = b[13] & g[9092];
assign g[17285] = a[13] & g[9093];
assign g[25476] = b[13] & g[9093];
assign g[17286] = a[13] & g[9094];
assign g[25477] = b[13] & g[9094];
assign g[17287] = a[13] & g[9095];
assign g[25478] = b[13] & g[9095];
assign g[17288] = a[13] & g[9096];
assign g[25479] = b[13] & g[9096];
assign g[17289] = a[13] & g[9097];
assign g[25480] = b[13] & g[9097];
assign g[17290] = a[13] & g[9098];
assign g[25481] = b[13] & g[9098];
assign g[17291] = a[13] & g[9099];
assign g[25482] = b[13] & g[9099];
assign g[17292] = a[13] & g[9100];
assign g[25483] = b[13] & g[9100];
assign g[17293] = a[13] & g[9101];
assign g[25484] = b[13] & g[9101];
assign g[17294] = a[13] & g[9102];
assign g[25485] = b[13] & g[9102];
assign g[17295] = a[13] & g[9103];
assign g[25486] = b[13] & g[9103];
assign g[17296] = a[13] & g[9104];
assign g[25487] = b[13] & g[9104];
assign g[17297] = a[13] & g[9105];
assign g[25488] = b[13] & g[9105];
assign g[17298] = a[13] & g[9106];
assign g[25489] = b[13] & g[9106];
assign g[17299] = a[13] & g[9107];
assign g[25490] = b[13] & g[9107];
assign g[17300] = a[13] & g[9108];
assign g[25491] = b[13] & g[9108];
assign g[17301] = a[13] & g[9109];
assign g[25492] = b[13] & g[9109];
assign g[17302] = a[13] & g[9110];
assign g[25493] = b[13] & g[9110];
assign g[17303] = a[13] & g[9111];
assign g[25494] = b[13] & g[9111];
assign g[17304] = a[13] & g[9112];
assign g[25495] = b[13] & g[9112];
assign g[17305] = a[13] & g[9113];
assign g[25496] = b[13] & g[9113];
assign g[17306] = a[13] & g[9114];
assign g[25497] = b[13] & g[9114];
assign g[17307] = a[13] & g[9115];
assign g[25498] = b[13] & g[9115];
assign g[17308] = a[13] & g[9116];
assign g[25499] = b[13] & g[9116];
assign g[17309] = a[13] & g[9117];
assign g[25500] = b[13] & g[9117];
assign g[17310] = a[13] & g[9118];
assign g[25501] = b[13] & g[9118];
assign g[17311] = a[13] & g[9119];
assign g[25502] = b[13] & g[9119];
assign g[17312] = a[13] & g[9120];
assign g[25503] = b[13] & g[9120];
assign g[17313] = a[13] & g[9121];
assign g[25504] = b[13] & g[9121];
assign g[17314] = a[13] & g[9122];
assign g[25505] = b[13] & g[9122];
assign g[17315] = a[13] & g[9123];
assign g[25506] = b[13] & g[9123];
assign g[17316] = a[13] & g[9124];
assign g[25507] = b[13] & g[9124];
assign g[17317] = a[13] & g[9125];
assign g[25508] = b[13] & g[9125];
assign g[17318] = a[13] & g[9126];
assign g[25509] = b[13] & g[9126];
assign g[17319] = a[13] & g[9127];
assign g[25510] = b[13] & g[9127];
assign g[17320] = a[13] & g[9128];
assign g[25511] = b[13] & g[9128];
assign g[17321] = a[13] & g[9129];
assign g[25512] = b[13] & g[9129];
assign g[17322] = a[13] & g[9130];
assign g[25513] = b[13] & g[9130];
assign g[17323] = a[13] & g[9131];
assign g[25514] = b[13] & g[9131];
assign g[17324] = a[13] & g[9132];
assign g[25515] = b[13] & g[9132];
assign g[17325] = a[13] & g[9133];
assign g[25516] = b[13] & g[9133];
assign g[17326] = a[13] & g[9134];
assign g[25517] = b[13] & g[9134];
assign g[17327] = a[13] & g[9135];
assign g[25518] = b[13] & g[9135];
assign g[17328] = a[13] & g[9136];
assign g[25519] = b[13] & g[9136];
assign g[17329] = a[13] & g[9137];
assign g[25520] = b[13] & g[9137];
assign g[17330] = a[13] & g[9138];
assign g[25521] = b[13] & g[9138];
assign g[17331] = a[13] & g[9139];
assign g[25522] = b[13] & g[9139];
assign g[17332] = a[13] & g[9140];
assign g[25523] = b[13] & g[9140];
assign g[17333] = a[13] & g[9141];
assign g[25524] = b[13] & g[9141];
assign g[17334] = a[13] & g[9142];
assign g[25525] = b[13] & g[9142];
assign g[17335] = a[13] & g[9143];
assign g[25526] = b[13] & g[9143];
assign g[17336] = a[13] & g[9144];
assign g[25527] = b[13] & g[9144];
assign g[17337] = a[13] & g[9145];
assign g[25528] = b[13] & g[9145];
assign g[17338] = a[13] & g[9146];
assign g[25529] = b[13] & g[9146];
assign g[17339] = a[13] & g[9147];
assign g[25530] = b[13] & g[9147];
assign g[17340] = a[13] & g[9148];
assign g[25531] = b[13] & g[9148];
assign g[17341] = a[13] & g[9149];
assign g[25532] = b[13] & g[9149];
assign g[17342] = a[13] & g[9150];
assign g[25533] = b[13] & g[9150];
assign g[17343] = a[13] & g[9151];
assign g[25534] = b[13] & g[9151];
assign g[17344] = a[13] & g[9152];
assign g[25535] = b[13] & g[9152];
assign g[17345] = a[13] & g[9153];
assign g[25536] = b[13] & g[9153];
assign g[17346] = a[13] & g[9154];
assign g[25537] = b[13] & g[9154];
assign g[17347] = a[13] & g[9155];
assign g[25538] = b[13] & g[9155];
assign g[17348] = a[13] & g[9156];
assign g[25539] = b[13] & g[9156];
assign g[17349] = a[13] & g[9157];
assign g[25540] = b[13] & g[9157];
assign g[17350] = a[13] & g[9158];
assign g[25541] = b[13] & g[9158];
assign g[17351] = a[13] & g[9159];
assign g[25542] = b[13] & g[9159];
assign g[17352] = a[13] & g[9160];
assign g[25543] = b[13] & g[9160];
assign g[17353] = a[13] & g[9161];
assign g[25544] = b[13] & g[9161];
assign g[17354] = a[13] & g[9162];
assign g[25545] = b[13] & g[9162];
assign g[17355] = a[13] & g[9163];
assign g[25546] = b[13] & g[9163];
assign g[17356] = a[13] & g[9164];
assign g[25547] = b[13] & g[9164];
assign g[17357] = a[13] & g[9165];
assign g[25548] = b[13] & g[9165];
assign g[17358] = a[13] & g[9166];
assign g[25549] = b[13] & g[9166];
assign g[17359] = a[13] & g[9167];
assign g[25550] = b[13] & g[9167];
assign g[17360] = a[13] & g[9168];
assign g[25551] = b[13] & g[9168];
assign g[17361] = a[13] & g[9169];
assign g[25552] = b[13] & g[9169];
assign g[17362] = a[13] & g[9170];
assign g[25553] = b[13] & g[9170];
assign g[17363] = a[13] & g[9171];
assign g[25554] = b[13] & g[9171];
assign g[17364] = a[13] & g[9172];
assign g[25555] = b[13] & g[9172];
assign g[17365] = a[13] & g[9173];
assign g[25556] = b[13] & g[9173];
assign g[17366] = a[13] & g[9174];
assign g[25557] = b[13] & g[9174];
assign g[17367] = a[13] & g[9175];
assign g[25558] = b[13] & g[9175];
assign g[17368] = a[13] & g[9176];
assign g[25559] = b[13] & g[9176];
assign g[17369] = a[13] & g[9177];
assign g[25560] = b[13] & g[9177];
assign g[17370] = a[13] & g[9178];
assign g[25561] = b[13] & g[9178];
assign g[17371] = a[13] & g[9179];
assign g[25562] = b[13] & g[9179];
assign g[17372] = a[13] & g[9180];
assign g[25563] = b[13] & g[9180];
assign g[17373] = a[13] & g[9181];
assign g[25564] = b[13] & g[9181];
assign g[17374] = a[13] & g[9182];
assign g[25565] = b[13] & g[9182];
assign g[17375] = a[13] & g[9183];
assign g[25566] = b[13] & g[9183];
assign g[17376] = a[13] & g[9184];
assign g[25567] = b[13] & g[9184];
assign g[17377] = a[13] & g[9185];
assign g[25568] = b[13] & g[9185];
assign g[17378] = a[13] & g[9186];
assign g[25569] = b[13] & g[9186];
assign g[17379] = a[13] & g[9187];
assign g[25570] = b[13] & g[9187];
assign g[17380] = a[13] & g[9188];
assign g[25571] = b[13] & g[9188];
assign g[17381] = a[13] & g[9189];
assign g[25572] = b[13] & g[9189];
assign g[17382] = a[13] & g[9190];
assign g[25573] = b[13] & g[9190];
assign g[17383] = a[13] & g[9191];
assign g[25574] = b[13] & g[9191];
assign g[17384] = a[13] & g[9192];
assign g[25575] = b[13] & g[9192];
assign g[17385] = a[13] & g[9193];
assign g[25576] = b[13] & g[9193];
assign g[17386] = a[13] & g[9194];
assign g[25577] = b[13] & g[9194];
assign g[17387] = a[13] & g[9195];
assign g[25578] = b[13] & g[9195];
assign g[17388] = a[13] & g[9196];
assign g[25579] = b[13] & g[9196];
assign g[17389] = a[13] & g[9197];
assign g[25580] = b[13] & g[9197];
assign g[17390] = a[13] & g[9198];
assign g[25581] = b[13] & g[9198];
assign g[17391] = a[13] & g[9199];
assign g[25582] = b[13] & g[9199];
assign g[17392] = a[13] & g[9200];
assign g[25583] = b[13] & g[9200];
assign g[17393] = a[13] & g[9201];
assign g[25584] = b[13] & g[9201];
assign g[17394] = a[13] & g[9202];
assign g[25585] = b[13] & g[9202];
assign g[17395] = a[13] & g[9203];
assign g[25586] = b[13] & g[9203];
assign g[17396] = a[13] & g[9204];
assign g[25587] = b[13] & g[9204];
assign g[17397] = a[13] & g[9205];
assign g[25588] = b[13] & g[9205];
assign g[17398] = a[13] & g[9206];
assign g[25589] = b[13] & g[9206];
assign g[17399] = a[13] & g[9207];
assign g[25590] = b[13] & g[9207];
assign g[17400] = a[13] & g[9208];
assign g[25591] = b[13] & g[9208];
assign g[17401] = a[13] & g[9209];
assign g[25592] = b[13] & g[9209];
assign g[17402] = a[13] & g[9210];
assign g[25593] = b[13] & g[9210];
assign g[17403] = a[13] & g[9211];
assign g[25594] = b[13] & g[9211];
assign g[17404] = a[13] & g[9212];
assign g[25595] = b[13] & g[9212];
assign g[17405] = a[13] & g[9213];
assign g[25596] = b[13] & g[9213];
assign g[17406] = a[13] & g[9214];
assign g[25597] = b[13] & g[9214];
assign g[17407] = a[13] & g[9215];
assign g[25598] = b[13] & g[9215];
assign g[17408] = a[13] & g[9216];
assign g[25599] = b[13] & g[9216];
assign g[17409] = a[13] & g[9217];
assign g[25600] = b[13] & g[9217];
assign g[17410] = a[13] & g[9218];
assign g[25601] = b[13] & g[9218];
assign g[17411] = a[13] & g[9219];
assign g[25602] = b[13] & g[9219];
assign g[17412] = a[13] & g[9220];
assign g[25603] = b[13] & g[9220];
assign g[17413] = a[13] & g[9221];
assign g[25604] = b[13] & g[9221];
assign g[17414] = a[13] & g[9222];
assign g[25605] = b[13] & g[9222];
assign g[17415] = a[13] & g[9223];
assign g[25606] = b[13] & g[9223];
assign g[17416] = a[13] & g[9224];
assign g[25607] = b[13] & g[9224];
assign g[17417] = a[13] & g[9225];
assign g[25608] = b[13] & g[9225];
assign g[17418] = a[13] & g[9226];
assign g[25609] = b[13] & g[9226];
assign g[17419] = a[13] & g[9227];
assign g[25610] = b[13] & g[9227];
assign g[17420] = a[13] & g[9228];
assign g[25611] = b[13] & g[9228];
assign g[17421] = a[13] & g[9229];
assign g[25612] = b[13] & g[9229];
assign g[17422] = a[13] & g[9230];
assign g[25613] = b[13] & g[9230];
assign g[17423] = a[13] & g[9231];
assign g[25614] = b[13] & g[9231];
assign g[17424] = a[13] & g[9232];
assign g[25615] = b[13] & g[9232];
assign g[17425] = a[13] & g[9233];
assign g[25616] = b[13] & g[9233];
assign g[17426] = a[13] & g[9234];
assign g[25617] = b[13] & g[9234];
assign g[17427] = a[13] & g[9235];
assign g[25618] = b[13] & g[9235];
assign g[17428] = a[13] & g[9236];
assign g[25619] = b[13] & g[9236];
assign g[17429] = a[13] & g[9237];
assign g[25620] = b[13] & g[9237];
assign g[17430] = a[13] & g[9238];
assign g[25621] = b[13] & g[9238];
assign g[17431] = a[13] & g[9239];
assign g[25622] = b[13] & g[9239];
assign g[17432] = a[13] & g[9240];
assign g[25623] = b[13] & g[9240];
assign g[17433] = a[13] & g[9241];
assign g[25624] = b[13] & g[9241];
assign g[17434] = a[13] & g[9242];
assign g[25625] = b[13] & g[9242];
assign g[17435] = a[13] & g[9243];
assign g[25626] = b[13] & g[9243];
assign g[17436] = a[13] & g[9244];
assign g[25627] = b[13] & g[9244];
assign g[17437] = a[13] & g[9245];
assign g[25628] = b[13] & g[9245];
assign g[17438] = a[13] & g[9246];
assign g[25629] = b[13] & g[9246];
assign g[17439] = a[13] & g[9247];
assign g[25630] = b[13] & g[9247];
assign g[17440] = a[13] & g[9248];
assign g[25631] = b[13] & g[9248];
assign g[17441] = a[13] & g[9249];
assign g[25632] = b[13] & g[9249];
assign g[17442] = a[13] & g[9250];
assign g[25633] = b[13] & g[9250];
assign g[17443] = a[13] & g[9251];
assign g[25634] = b[13] & g[9251];
assign g[17444] = a[13] & g[9252];
assign g[25635] = b[13] & g[9252];
assign g[17445] = a[13] & g[9253];
assign g[25636] = b[13] & g[9253];
assign g[17446] = a[13] & g[9254];
assign g[25637] = b[13] & g[9254];
assign g[17447] = a[13] & g[9255];
assign g[25638] = b[13] & g[9255];
assign g[17448] = a[13] & g[9256];
assign g[25639] = b[13] & g[9256];
assign g[17449] = a[13] & g[9257];
assign g[25640] = b[13] & g[9257];
assign g[17450] = a[13] & g[9258];
assign g[25641] = b[13] & g[9258];
assign g[17451] = a[13] & g[9259];
assign g[25642] = b[13] & g[9259];
assign g[17452] = a[13] & g[9260];
assign g[25643] = b[13] & g[9260];
assign g[17453] = a[13] & g[9261];
assign g[25644] = b[13] & g[9261];
assign g[17454] = a[13] & g[9262];
assign g[25645] = b[13] & g[9262];
assign g[17455] = a[13] & g[9263];
assign g[25646] = b[13] & g[9263];
assign g[17456] = a[13] & g[9264];
assign g[25647] = b[13] & g[9264];
assign g[17457] = a[13] & g[9265];
assign g[25648] = b[13] & g[9265];
assign g[17458] = a[13] & g[9266];
assign g[25649] = b[13] & g[9266];
assign g[17459] = a[13] & g[9267];
assign g[25650] = b[13] & g[9267];
assign g[17460] = a[13] & g[9268];
assign g[25651] = b[13] & g[9268];
assign g[17461] = a[13] & g[9269];
assign g[25652] = b[13] & g[9269];
assign g[17462] = a[13] & g[9270];
assign g[25653] = b[13] & g[9270];
assign g[17463] = a[13] & g[9271];
assign g[25654] = b[13] & g[9271];
assign g[17464] = a[13] & g[9272];
assign g[25655] = b[13] & g[9272];
assign g[17465] = a[13] & g[9273];
assign g[25656] = b[13] & g[9273];
assign g[17466] = a[13] & g[9274];
assign g[25657] = b[13] & g[9274];
assign g[17467] = a[13] & g[9275];
assign g[25658] = b[13] & g[9275];
assign g[17468] = a[13] & g[9276];
assign g[25659] = b[13] & g[9276];
assign g[17469] = a[13] & g[9277];
assign g[25660] = b[13] & g[9277];
assign g[17470] = a[13] & g[9278];
assign g[25661] = b[13] & g[9278];
assign g[17471] = a[13] & g[9279];
assign g[25662] = b[13] & g[9279];
assign g[17472] = a[13] & g[9280];
assign g[25663] = b[13] & g[9280];
assign g[17473] = a[13] & g[9281];
assign g[25664] = b[13] & g[9281];
assign g[17474] = a[13] & g[9282];
assign g[25665] = b[13] & g[9282];
assign g[17475] = a[13] & g[9283];
assign g[25666] = b[13] & g[9283];
assign g[17476] = a[13] & g[9284];
assign g[25667] = b[13] & g[9284];
assign g[17477] = a[13] & g[9285];
assign g[25668] = b[13] & g[9285];
assign g[17478] = a[13] & g[9286];
assign g[25669] = b[13] & g[9286];
assign g[17479] = a[13] & g[9287];
assign g[25670] = b[13] & g[9287];
assign g[17480] = a[13] & g[9288];
assign g[25671] = b[13] & g[9288];
assign g[17481] = a[13] & g[9289];
assign g[25672] = b[13] & g[9289];
assign g[17482] = a[13] & g[9290];
assign g[25673] = b[13] & g[9290];
assign g[17483] = a[13] & g[9291];
assign g[25674] = b[13] & g[9291];
assign g[17484] = a[13] & g[9292];
assign g[25675] = b[13] & g[9292];
assign g[17485] = a[13] & g[9293];
assign g[25676] = b[13] & g[9293];
assign g[17486] = a[13] & g[9294];
assign g[25677] = b[13] & g[9294];
assign g[17487] = a[13] & g[9295];
assign g[25678] = b[13] & g[9295];
assign g[17488] = a[13] & g[9296];
assign g[25679] = b[13] & g[9296];
assign g[17489] = a[13] & g[9297];
assign g[25680] = b[13] & g[9297];
assign g[17490] = a[13] & g[9298];
assign g[25681] = b[13] & g[9298];
assign g[17491] = a[13] & g[9299];
assign g[25682] = b[13] & g[9299];
assign g[17492] = a[13] & g[9300];
assign g[25683] = b[13] & g[9300];
assign g[17493] = a[13] & g[9301];
assign g[25684] = b[13] & g[9301];
assign g[17494] = a[13] & g[9302];
assign g[25685] = b[13] & g[9302];
assign g[17495] = a[13] & g[9303];
assign g[25686] = b[13] & g[9303];
assign g[17496] = a[13] & g[9304];
assign g[25687] = b[13] & g[9304];
assign g[17497] = a[13] & g[9305];
assign g[25688] = b[13] & g[9305];
assign g[17498] = a[13] & g[9306];
assign g[25689] = b[13] & g[9306];
assign g[17499] = a[13] & g[9307];
assign g[25690] = b[13] & g[9307];
assign g[17500] = a[13] & g[9308];
assign g[25691] = b[13] & g[9308];
assign g[17501] = a[13] & g[9309];
assign g[25692] = b[13] & g[9309];
assign g[17502] = a[13] & g[9310];
assign g[25693] = b[13] & g[9310];
assign g[17503] = a[13] & g[9311];
assign g[25694] = b[13] & g[9311];
assign g[17504] = a[13] & g[9312];
assign g[25695] = b[13] & g[9312];
assign g[17505] = a[13] & g[9313];
assign g[25696] = b[13] & g[9313];
assign g[17506] = a[13] & g[9314];
assign g[25697] = b[13] & g[9314];
assign g[17507] = a[13] & g[9315];
assign g[25698] = b[13] & g[9315];
assign g[17508] = a[13] & g[9316];
assign g[25699] = b[13] & g[9316];
assign g[17509] = a[13] & g[9317];
assign g[25700] = b[13] & g[9317];
assign g[17510] = a[13] & g[9318];
assign g[25701] = b[13] & g[9318];
assign g[17511] = a[13] & g[9319];
assign g[25702] = b[13] & g[9319];
assign g[17512] = a[13] & g[9320];
assign g[25703] = b[13] & g[9320];
assign g[17513] = a[13] & g[9321];
assign g[25704] = b[13] & g[9321];
assign g[17514] = a[13] & g[9322];
assign g[25705] = b[13] & g[9322];
assign g[17515] = a[13] & g[9323];
assign g[25706] = b[13] & g[9323];
assign g[17516] = a[13] & g[9324];
assign g[25707] = b[13] & g[9324];
assign g[17517] = a[13] & g[9325];
assign g[25708] = b[13] & g[9325];
assign g[17518] = a[13] & g[9326];
assign g[25709] = b[13] & g[9326];
assign g[17519] = a[13] & g[9327];
assign g[25710] = b[13] & g[9327];
assign g[17520] = a[13] & g[9328];
assign g[25711] = b[13] & g[9328];
assign g[17521] = a[13] & g[9329];
assign g[25712] = b[13] & g[9329];
assign g[17522] = a[13] & g[9330];
assign g[25713] = b[13] & g[9330];
assign g[17523] = a[13] & g[9331];
assign g[25714] = b[13] & g[9331];
assign g[17524] = a[13] & g[9332];
assign g[25715] = b[13] & g[9332];
assign g[17525] = a[13] & g[9333];
assign g[25716] = b[13] & g[9333];
assign g[17526] = a[13] & g[9334];
assign g[25717] = b[13] & g[9334];
assign g[17527] = a[13] & g[9335];
assign g[25718] = b[13] & g[9335];
assign g[17528] = a[13] & g[9336];
assign g[25719] = b[13] & g[9336];
assign g[17529] = a[13] & g[9337];
assign g[25720] = b[13] & g[9337];
assign g[17530] = a[13] & g[9338];
assign g[25721] = b[13] & g[9338];
assign g[17531] = a[13] & g[9339];
assign g[25722] = b[13] & g[9339];
assign g[17532] = a[13] & g[9340];
assign g[25723] = b[13] & g[9340];
assign g[17533] = a[13] & g[9341];
assign g[25724] = b[13] & g[9341];
assign g[17534] = a[13] & g[9342];
assign g[25725] = b[13] & g[9342];
assign g[17535] = a[13] & g[9343];
assign g[25726] = b[13] & g[9343];
assign g[17536] = a[13] & g[9344];
assign g[25727] = b[13] & g[9344];
assign g[17537] = a[13] & g[9345];
assign g[25728] = b[13] & g[9345];
assign g[17538] = a[13] & g[9346];
assign g[25729] = b[13] & g[9346];
assign g[17539] = a[13] & g[9347];
assign g[25730] = b[13] & g[9347];
assign g[17540] = a[13] & g[9348];
assign g[25731] = b[13] & g[9348];
assign g[17541] = a[13] & g[9349];
assign g[25732] = b[13] & g[9349];
assign g[17542] = a[13] & g[9350];
assign g[25733] = b[13] & g[9350];
assign g[17543] = a[13] & g[9351];
assign g[25734] = b[13] & g[9351];
assign g[17544] = a[13] & g[9352];
assign g[25735] = b[13] & g[9352];
assign g[17545] = a[13] & g[9353];
assign g[25736] = b[13] & g[9353];
assign g[17546] = a[13] & g[9354];
assign g[25737] = b[13] & g[9354];
assign g[17547] = a[13] & g[9355];
assign g[25738] = b[13] & g[9355];
assign g[17548] = a[13] & g[9356];
assign g[25739] = b[13] & g[9356];
assign g[17549] = a[13] & g[9357];
assign g[25740] = b[13] & g[9357];
assign g[17550] = a[13] & g[9358];
assign g[25741] = b[13] & g[9358];
assign g[17551] = a[13] & g[9359];
assign g[25742] = b[13] & g[9359];
assign g[17552] = a[13] & g[9360];
assign g[25743] = b[13] & g[9360];
assign g[17553] = a[13] & g[9361];
assign g[25744] = b[13] & g[9361];
assign g[17554] = a[13] & g[9362];
assign g[25745] = b[13] & g[9362];
assign g[17555] = a[13] & g[9363];
assign g[25746] = b[13] & g[9363];
assign g[17556] = a[13] & g[9364];
assign g[25747] = b[13] & g[9364];
assign g[17557] = a[13] & g[9365];
assign g[25748] = b[13] & g[9365];
assign g[17558] = a[13] & g[9366];
assign g[25749] = b[13] & g[9366];
assign g[17559] = a[13] & g[9367];
assign g[25750] = b[13] & g[9367];
assign g[17560] = a[13] & g[9368];
assign g[25751] = b[13] & g[9368];
assign g[17561] = a[13] & g[9369];
assign g[25752] = b[13] & g[9369];
assign g[17562] = a[13] & g[9370];
assign g[25753] = b[13] & g[9370];
assign g[17563] = a[13] & g[9371];
assign g[25754] = b[13] & g[9371];
assign g[17564] = a[13] & g[9372];
assign g[25755] = b[13] & g[9372];
assign g[17565] = a[13] & g[9373];
assign g[25756] = b[13] & g[9373];
assign g[17566] = a[13] & g[9374];
assign g[25757] = b[13] & g[9374];
assign g[17567] = a[13] & g[9375];
assign g[25758] = b[13] & g[9375];
assign g[17568] = a[13] & g[9376];
assign g[25759] = b[13] & g[9376];
assign g[17569] = a[13] & g[9377];
assign g[25760] = b[13] & g[9377];
assign g[17570] = a[13] & g[9378];
assign g[25761] = b[13] & g[9378];
assign g[17571] = a[13] & g[9379];
assign g[25762] = b[13] & g[9379];
assign g[17572] = a[13] & g[9380];
assign g[25763] = b[13] & g[9380];
assign g[17573] = a[13] & g[9381];
assign g[25764] = b[13] & g[9381];
assign g[17574] = a[13] & g[9382];
assign g[25765] = b[13] & g[9382];
assign g[17575] = a[13] & g[9383];
assign g[25766] = b[13] & g[9383];
assign g[17576] = a[13] & g[9384];
assign g[25767] = b[13] & g[9384];
assign g[17577] = a[13] & g[9385];
assign g[25768] = b[13] & g[9385];
assign g[17578] = a[13] & g[9386];
assign g[25769] = b[13] & g[9386];
assign g[17579] = a[13] & g[9387];
assign g[25770] = b[13] & g[9387];
assign g[17580] = a[13] & g[9388];
assign g[25771] = b[13] & g[9388];
assign g[17581] = a[13] & g[9389];
assign g[25772] = b[13] & g[9389];
assign g[17582] = a[13] & g[9390];
assign g[25773] = b[13] & g[9390];
assign g[17583] = a[13] & g[9391];
assign g[25774] = b[13] & g[9391];
assign g[17584] = a[13] & g[9392];
assign g[25775] = b[13] & g[9392];
assign g[17585] = a[13] & g[9393];
assign g[25776] = b[13] & g[9393];
assign g[17586] = a[13] & g[9394];
assign g[25777] = b[13] & g[9394];
assign g[17587] = a[13] & g[9395];
assign g[25778] = b[13] & g[9395];
assign g[17588] = a[13] & g[9396];
assign g[25779] = b[13] & g[9396];
assign g[17589] = a[13] & g[9397];
assign g[25780] = b[13] & g[9397];
assign g[17590] = a[13] & g[9398];
assign g[25781] = b[13] & g[9398];
assign g[17591] = a[13] & g[9399];
assign g[25782] = b[13] & g[9399];
assign g[17592] = a[13] & g[9400];
assign g[25783] = b[13] & g[9400];
assign g[17593] = a[13] & g[9401];
assign g[25784] = b[13] & g[9401];
assign g[17594] = a[13] & g[9402];
assign g[25785] = b[13] & g[9402];
assign g[17595] = a[13] & g[9403];
assign g[25786] = b[13] & g[9403];
assign g[17596] = a[13] & g[9404];
assign g[25787] = b[13] & g[9404];
assign g[17597] = a[13] & g[9405];
assign g[25788] = b[13] & g[9405];
assign g[17598] = a[13] & g[9406];
assign g[25789] = b[13] & g[9406];
assign g[17599] = a[13] & g[9407];
assign g[25790] = b[13] & g[9407];
assign g[17600] = a[13] & g[9408];
assign g[25791] = b[13] & g[9408];
assign g[17601] = a[13] & g[9409];
assign g[25792] = b[13] & g[9409];
assign g[17602] = a[13] & g[9410];
assign g[25793] = b[13] & g[9410];
assign g[17603] = a[13] & g[9411];
assign g[25794] = b[13] & g[9411];
assign g[17604] = a[13] & g[9412];
assign g[25795] = b[13] & g[9412];
assign g[17605] = a[13] & g[9413];
assign g[25796] = b[13] & g[9413];
assign g[17606] = a[13] & g[9414];
assign g[25797] = b[13] & g[9414];
assign g[17607] = a[13] & g[9415];
assign g[25798] = b[13] & g[9415];
assign g[17608] = a[13] & g[9416];
assign g[25799] = b[13] & g[9416];
assign g[17609] = a[13] & g[9417];
assign g[25800] = b[13] & g[9417];
assign g[17610] = a[13] & g[9418];
assign g[25801] = b[13] & g[9418];
assign g[17611] = a[13] & g[9419];
assign g[25802] = b[13] & g[9419];
assign g[17612] = a[13] & g[9420];
assign g[25803] = b[13] & g[9420];
assign g[17613] = a[13] & g[9421];
assign g[25804] = b[13] & g[9421];
assign g[17614] = a[13] & g[9422];
assign g[25805] = b[13] & g[9422];
assign g[17615] = a[13] & g[9423];
assign g[25806] = b[13] & g[9423];
assign g[17616] = a[13] & g[9424];
assign g[25807] = b[13] & g[9424];
assign g[17617] = a[13] & g[9425];
assign g[25808] = b[13] & g[9425];
assign g[17618] = a[13] & g[9426];
assign g[25809] = b[13] & g[9426];
assign g[17619] = a[13] & g[9427];
assign g[25810] = b[13] & g[9427];
assign g[17620] = a[13] & g[9428];
assign g[25811] = b[13] & g[9428];
assign g[17621] = a[13] & g[9429];
assign g[25812] = b[13] & g[9429];
assign g[17622] = a[13] & g[9430];
assign g[25813] = b[13] & g[9430];
assign g[17623] = a[13] & g[9431];
assign g[25814] = b[13] & g[9431];
assign g[17624] = a[13] & g[9432];
assign g[25815] = b[13] & g[9432];
assign g[17625] = a[13] & g[9433];
assign g[25816] = b[13] & g[9433];
assign g[17626] = a[13] & g[9434];
assign g[25817] = b[13] & g[9434];
assign g[17627] = a[13] & g[9435];
assign g[25818] = b[13] & g[9435];
assign g[17628] = a[13] & g[9436];
assign g[25819] = b[13] & g[9436];
assign g[17629] = a[13] & g[9437];
assign g[25820] = b[13] & g[9437];
assign g[17630] = a[13] & g[9438];
assign g[25821] = b[13] & g[9438];
assign g[17631] = a[13] & g[9439];
assign g[25822] = b[13] & g[9439];
assign g[17632] = a[13] & g[9440];
assign g[25823] = b[13] & g[9440];
assign g[17633] = a[13] & g[9441];
assign g[25824] = b[13] & g[9441];
assign g[17634] = a[13] & g[9442];
assign g[25825] = b[13] & g[9442];
assign g[17635] = a[13] & g[9443];
assign g[25826] = b[13] & g[9443];
assign g[17636] = a[13] & g[9444];
assign g[25827] = b[13] & g[9444];
assign g[17637] = a[13] & g[9445];
assign g[25828] = b[13] & g[9445];
assign g[17638] = a[13] & g[9446];
assign g[25829] = b[13] & g[9446];
assign g[17639] = a[13] & g[9447];
assign g[25830] = b[13] & g[9447];
assign g[17640] = a[13] & g[9448];
assign g[25831] = b[13] & g[9448];
assign g[17641] = a[13] & g[9449];
assign g[25832] = b[13] & g[9449];
assign g[17642] = a[13] & g[9450];
assign g[25833] = b[13] & g[9450];
assign g[17643] = a[13] & g[9451];
assign g[25834] = b[13] & g[9451];
assign g[17644] = a[13] & g[9452];
assign g[25835] = b[13] & g[9452];
assign g[17645] = a[13] & g[9453];
assign g[25836] = b[13] & g[9453];
assign g[17646] = a[13] & g[9454];
assign g[25837] = b[13] & g[9454];
assign g[17647] = a[13] & g[9455];
assign g[25838] = b[13] & g[9455];
assign g[17648] = a[13] & g[9456];
assign g[25839] = b[13] & g[9456];
assign g[17649] = a[13] & g[9457];
assign g[25840] = b[13] & g[9457];
assign g[17650] = a[13] & g[9458];
assign g[25841] = b[13] & g[9458];
assign g[17651] = a[13] & g[9459];
assign g[25842] = b[13] & g[9459];
assign g[17652] = a[13] & g[9460];
assign g[25843] = b[13] & g[9460];
assign g[17653] = a[13] & g[9461];
assign g[25844] = b[13] & g[9461];
assign g[17654] = a[13] & g[9462];
assign g[25845] = b[13] & g[9462];
assign g[17655] = a[13] & g[9463];
assign g[25846] = b[13] & g[9463];
assign g[17656] = a[13] & g[9464];
assign g[25847] = b[13] & g[9464];
assign g[17657] = a[13] & g[9465];
assign g[25848] = b[13] & g[9465];
assign g[17658] = a[13] & g[9466];
assign g[25849] = b[13] & g[9466];
assign g[17659] = a[13] & g[9467];
assign g[25850] = b[13] & g[9467];
assign g[17660] = a[13] & g[9468];
assign g[25851] = b[13] & g[9468];
assign g[17661] = a[13] & g[9469];
assign g[25852] = b[13] & g[9469];
assign g[17662] = a[13] & g[9470];
assign g[25853] = b[13] & g[9470];
assign g[17663] = a[13] & g[9471];
assign g[25854] = b[13] & g[9471];
assign g[17664] = a[13] & g[9472];
assign g[25855] = b[13] & g[9472];
assign g[17665] = a[13] & g[9473];
assign g[25856] = b[13] & g[9473];
assign g[17666] = a[13] & g[9474];
assign g[25857] = b[13] & g[9474];
assign g[17667] = a[13] & g[9475];
assign g[25858] = b[13] & g[9475];
assign g[17668] = a[13] & g[9476];
assign g[25859] = b[13] & g[9476];
assign g[17669] = a[13] & g[9477];
assign g[25860] = b[13] & g[9477];
assign g[17670] = a[13] & g[9478];
assign g[25861] = b[13] & g[9478];
assign g[17671] = a[13] & g[9479];
assign g[25862] = b[13] & g[9479];
assign g[17672] = a[13] & g[9480];
assign g[25863] = b[13] & g[9480];
assign g[17673] = a[13] & g[9481];
assign g[25864] = b[13] & g[9481];
assign g[17674] = a[13] & g[9482];
assign g[25865] = b[13] & g[9482];
assign g[17675] = a[13] & g[9483];
assign g[25866] = b[13] & g[9483];
assign g[17676] = a[13] & g[9484];
assign g[25867] = b[13] & g[9484];
assign g[17677] = a[13] & g[9485];
assign g[25868] = b[13] & g[9485];
assign g[17678] = a[13] & g[9486];
assign g[25869] = b[13] & g[9486];
assign g[17679] = a[13] & g[9487];
assign g[25870] = b[13] & g[9487];
assign g[17680] = a[13] & g[9488];
assign g[25871] = b[13] & g[9488];
assign g[17681] = a[13] & g[9489];
assign g[25872] = b[13] & g[9489];
assign g[17682] = a[13] & g[9490];
assign g[25873] = b[13] & g[9490];
assign g[17683] = a[13] & g[9491];
assign g[25874] = b[13] & g[9491];
assign g[17684] = a[13] & g[9492];
assign g[25875] = b[13] & g[9492];
assign g[17685] = a[13] & g[9493];
assign g[25876] = b[13] & g[9493];
assign g[17686] = a[13] & g[9494];
assign g[25877] = b[13] & g[9494];
assign g[17687] = a[13] & g[9495];
assign g[25878] = b[13] & g[9495];
assign g[17688] = a[13] & g[9496];
assign g[25879] = b[13] & g[9496];
assign g[17689] = a[13] & g[9497];
assign g[25880] = b[13] & g[9497];
assign g[17690] = a[13] & g[9498];
assign g[25881] = b[13] & g[9498];
assign g[17691] = a[13] & g[9499];
assign g[25882] = b[13] & g[9499];
assign g[17692] = a[13] & g[9500];
assign g[25883] = b[13] & g[9500];
assign g[17693] = a[13] & g[9501];
assign g[25884] = b[13] & g[9501];
assign g[17694] = a[13] & g[9502];
assign g[25885] = b[13] & g[9502];
assign g[17695] = a[13] & g[9503];
assign g[25886] = b[13] & g[9503];
assign g[17696] = a[13] & g[9504];
assign g[25887] = b[13] & g[9504];
assign g[17697] = a[13] & g[9505];
assign g[25888] = b[13] & g[9505];
assign g[17698] = a[13] & g[9506];
assign g[25889] = b[13] & g[9506];
assign g[17699] = a[13] & g[9507];
assign g[25890] = b[13] & g[9507];
assign g[17700] = a[13] & g[9508];
assign g[25891] = b[13] & g[9508];
assign g[17701] = a[13] & g[9509];
assign g[25892] = b[13] & g[9509];
assign g[17702] = a[13] & g[9510];
assign g[25893] = b[13] & g[9510];
assign g[17703] = a[13] & g[9511];
assign g[25894] = b[13] & g[9511];
assign g[17704] = a[13] & g[9512];
assign g[25895] = b[13] & g[9512];
assign g[17705] = a[13] & g[9513];
assign g[25896] = b[13] & g[9513];
assign g[17706] = a[13] & g[9514];
assign g[25897] = b[13] & g[9514];
assign g[17707] = a[13] & g[9515];
assign g[25898] = b[13] & g[9515];
assign g[17708] = a[13] & g[9516];
assign g[25899] = b[13] & g[9516];
assign g[17709] = a[13] & g[9517];
assign g[25900] = b[13] & g[9517];
assign g[17710] = a[13] & g[9518];
assign g[25901] = b[13] & g[9518];
assign g[17711] = a[13] & g[9519];
assign g[25902] = b[13] & g[9519];
assign g[17712] = a[13] & g[9520];
assign g[25903] = b[13] & g[9520];
assign g[17713] = a[13] & g[9521];
assign g[25904] = b[13] & g[9521];
assign g[17714] = a[13] & g[9522];
assign g[25905] = b[13] & g[9522];
assign g[17715] = a[13] & g[9523];
assign g[25906] = b[13] & g[9523];
assign g[17716] = a[13] & g[9524];
assign g[25907] = b[13] & g[9524];
assign g[17717] = a[13] & g[9525];
assign g[25908] = b[13] & g[9525];
assign g[17718] = a[13] & g[9526];
assign g[25909] = b[13] & g[9526];
assign g[17719] = a[13] & g[9527];
assign g[25910] = b[13] & g[9527];
assign g[17720] = a[13] & g[9528];
assign g[25911] = b[13] & g[9528];
assign g[17721] = a[13] & g[9529];
assign g[25912] = b[13] & g[9529];
assign g[17722] = a[13] & g[9530];
assign g[25913] = b[13] & g[9530];
assign g[17723] = a[13] & g[9531];
assign g[25914] = b[13] & g[9531];
assign g[17724] = a[13] & g[9532];
assign g[25915] = b[13] & g[9532];
assign g[17725] = a[13] & g[9533];
assign g[25916] = b[13] & g[9533];
assign g[17726] = a[13] & g[9534];
assign g[25917] = b[13] & g[9534];
assign g[17727] = a[13] & g[9535];
assign g[25918] = b[13] & g[9535];
assign g[17728] = a[13] & g[9536];
assign g[25919] = b[13] & g[9536];
assign g[17729] = a[13] & g[9537];
assign g[25920] = b[13] & g[9537];
assign g[17730] = a[13] & g[9538];
assign g[25921] = b[13] & g[9538];
assign g[17731] = a[13] & g[9539];
assign g[25922] = b[13] & g[9539];
assign g[17732] = a[13] & g[9540];
assign g[25923] = b[13] & g[9540];
assign g[17733] = a[13] & g[9541];
assign g[25924] = b[13] & g[9541];
assign g[17734] = a[13] & g[9542];
assign g[25925] = b[13] & g[9542];
assign g[17735] = a[13] & g[9543];
assign g[25926] = b[13] & g[9543];
assign g[17736] = a[13] & g[9544];
assign g[25927] = b[13] & g[9544];
assign g[17737] = a[13] & g[9545];
assign g[25928] = b[13] & g[9545];
assign g[17738] = a[13] & g[9546];
assign g[25929] = b[13] & g[9546];
assign g[17739] = a[13] & g[9547];
assign g[25930] = b[13] & g[9547];
assign g[17740] = a[13] & g[9548];
assign g[25931] = b[13] & g[9548];
assign g[17741] = a[13] & g[9549];
assign g[25932] = b[13] & g[9549];
assign g[17742] = a[13] & g[9550];
assign g[25933] = b[13] & g[9550];
assign g[17743] = a[13] & g[9551];
assign g[25934] = b[13] & g[9551];
assign g[17744] = a[13] & g[9552];
assign g[25935] = b[13] & g[9552];
assign g[17745] = a[13] & g[9553];
assign g[25936] = b[13] & g[9553];
assign g[17746] = a[13] & g[9554];
assign g[25937] = b[13] & g[9554];
assign g[17747] = a[13] & g[9555];
assign g[25938] = b[13] & g[9555];
assign g[17748] = a[13] & g[9556];
assign g[25939] = b[13] & g[9556];
assign g[17749] = a[13] & g[9557];
assign g[25940] = b[13] & g[9557];
assign g[17750] = a[13] & g[9558];
assign g[25941] = b[13] & g[9558];
assign g[17751] = a[13] & g[9559];
assign g[25942] = b[13] & g[9559];
assign g[17752] = a[13] & g[9560];
assign g[25943] = b[13] & g[9560];
assign g[17753] = a[13] & g[9561];
assign g[25944] = b[13] & g[9561];
assign g[17754] = a[13] & g[9562];
assign g[25945] = b[13] & g[9562];
assign g[17755] = a[13] & g[9563];
assign g[25946] = b[13] & g[9563];
assign g[17756] = a[13] & g[9564];
assign g[25947] = b[13] & g[9564];
assign g[17757] = a[13] & g[9565];
assign g[25948] = b[13] & g[9565];
assign g[17758] = a[13] & g[9566];
assign g[25949] = b[13] & g[9566];
assign g[17759] = a[13] & g[9567];
assign g[25950] = b[13] & g[9567];
assign g[17760] = a[13] & g[9568];
assign g[25951] = b[13] & g[9568];
assign g[17761] = a[13] & g[9569];
assign g[25952] = b[13] & g[9569];
assign g[17762] = a[13] & g[9570];
assign g[25953] = b[13] & g[9570];
assign g[17763] = a[13] & g[9571];
assign g[25954] = b[13] & g[9571];
assign g[17764] = a[13] & g[9572];
assign g[25955] = b[13] & g[9572];
assign g[17765] = a[13] & g[9573];
assign g[25956] = b[13] & g[9573];
assign g[17766] = a[13] & g[9574];
assign g[25957] = b[13] & g[9574];
assign g[17767] = a[13] & g[9575];
assign g[25958] = b[13] & g[9575];
assign g[17768] = a[13] & g[9576];
assign g[25959] = b[13] & g[9576];
assign g[17769] = a[13] & g[9577];
assign g[25960] = b[13] & g[9577];
assign g[17770] = a[13] & g[9578];
assign g[25961] = b[13] & g[9578];
assign g[17771] = a[13] & g[9579];
assign g[25962] = b[13] & g[9579];
assign g[17772] = a[13] & g[9580];
assign g[25963] = b[13] & g[9580];
assign g[17773] = a[13] & g[9581];
assign g[25964] = b[13] & g[9581];
assign g[17774] = a[13] & g[9582];
assign g[25965] = b[13] & g[9582];
assign g[17775] = a[13] & g[9583];
assign g[25966] = b[13] & g[9583];
assign g[17776] = a[13] & g[9584];
assign g[25967] = b[13] & g[9584];
assign g[17777] = a[13] & g[9585];
assign g[25968] = b[13] & g[9585];
assign g[17778] = a[13] & g[9586];
assign g[25969] = b[13] & g[9586];
assign g[17779] = a[13] & g[9587];
assign g[25970] = b[13] & g[9587];
assign g[17780] = a[13] & g[9588];
assign g[25971] = b[13] & g[9588];
assign g[17781] = a[13] & g[9589];
assign g[25972] = b[13] & g[9589];
assign g[17782] = a[13] & g[9590];
assign g[25973] = b[13] & g[9590];
assign g[17783] = a[13] & g[9591];
assign g[25974] = b[13] & g[9591];
assign g[17784] = a[13] & g[9592];
assign g[25975] = b[13] & g[9592];
assign g[17785] = a[13] & g[9593];
assign g[25976] = b[13] & g[9593];
assign g[17786] = a[13] & g[9594];
assign g[25977] = b[13] & g[9594];
assign g[17787] = a[13] & g[9595];
assign g[25978] = b[13] & g[9595];
assign g[17788] = a[13] & g[9596];
assign g[25979] = b[13] & g[9596];
assign g[17789] = a[13] & g[9597];
assign g[25980] = b[13] & g[9597];
assign g[17790] = a[13] & g[9598];
assign g[25981] = b[13] & g[9598];
assign g[17791] = a[13] & g[9599];
assign g[25982] = b[13] & g[9599];
assign g[17792] = a[13] & g[9600];
assign g[25983] = b[13] & g[9600];
assign g[17793] = a[13] & g[9601];
assign g[25984] = b[13] & g[9601];
assign g[17794] = a[13] & g[9602];
assign g[25985] = b[13] & g[9602];
assign g[17795] = a[13] & g[9603];
assign g[25986] = b[13] & g[9603];
assign g[17796] = a[13] & g[9604];
assign g[25987] = b[13] & g[9604];
assign g[17797] = a[13] & g[9605];
assign g[25988] = b[13] & g[9605];
assign g[17798] = a[13] & g[9606];
assign g[25989] = b[13] & g[9606];
assign g[17799] = a[13] & g[9607];
assign g[25990] = b[13] & g[9607];
assign g[17800] = a[13] & g[9608];
assign g[25991] = b[13] & g[9608];
assign g[17801] = a[13] & g[9609];
assign g[25992] = b[13] & g[9609];
assign g[17802] = a[13] & g[9610];
assign g[25993] = b[13] & g[9610];
assign g[17803] = a[13] & g[9611];
assign g[25994] = b[13] & g[9611];
assign g[17804] = a[13] & g[9612];
assign g[25995] = b[13] & g[9612];
assign g[17805] = a[13] & g[9613];
assign g[25996] = b[13] & g[9613];
assign g[17806] = a[13] & g[9614];
assign g[25997] = b[13] & g[9614];
assign g[17807] = a[13] & g[9615];
assign g[25998] = b[13] & g[9615];
assign g[17808] = a[13] & g[9616];
assign g[25999] = b[13] & g[9616];
assign g[17809] = a[13] & g[9617];
assign g[26000] = b[13] & g[9617];
assign g[17810] = a[13] & g[9618];
assign g[26001] = b[13] & g[9618];
assign g[17811] = a[13] & g[9619];
assign g[26002] = b[13] & g[9619];
assign g[17812] = a[13] & g[9620];
assign g[26003] = b[13] & g[9620];
assign g[17813] = a[13] & g[9621];
assign g[26004] = b[13] & g[9621];
assign g[17814] = a[13] & g[9622];
assign g[26005] = b[13] & g[9622];
assign g[17815] = a[13] & g[9623];
assign g[26006] = b[13] & g[9623];
assign g[17816] = a[13] & g[9624];
assign g[26007] = b[13] & g[9624];
assign g[17817] = a[13] & g[9625];
assign g[26008] = b[13] & g[9625];
assign g[17818] = a[13] & g[9626];
assign g[26009] = b[13] & g[9626];
assign g[17819] = a[13] & g[9627];
assign g[26010] = b[13] & g[9627];
assign g[17820] = a[13] & g[9628];
assign g[26011] = b[13] & g[9628];
assign g[17821] = a[13] & g[9629];
assign g[26012] = b[13] & g[9629];
assign g[17822] = a[13] & g[9630];
assign g[26013] = b[13] & g[9630];
assign g[17823] = a[13] & g[9631];
assign g[26014] = b[13] & g[9631];
assign g[17824] = a[13] & g[9632];
assign g[26015] = b[13] & g[9632];
assign g[17825] = a[13] & g[9633];
assign g[26016] = b[13] & g[9633];
assign g[17826] = a[13] & g[9634];
assign g[26017] = b[13] & g[9634];
assign g[17827] = a[13] & g[9635];
assign g[26018] = b[13] & g[9635];
assign g[17828] = a[13] & g[9636];
assign g[26019] = b[13] & g[9636];
assign g[17829] = a[13] & g[9637];
assign g[26020] = b[13] & g[9637];
assign g[17830] = a[13] & g[9638];
assign g[26021] = b[13] & g[9638];
assign g[17831] = a[13] & g[9639];
assign g[26022] = b[13] & g[9639];
assign g[17832] = a[13] & g[9640];
assign g[26023] = b[13] & g[9640];
assign g[17833] = a[13] & g[9641];
assign g[26024] = b[13] & g[9641];
assign g[17834] = a[13] & g[9642];
assign g[26025] = b[13] & g[9642];
assign g[17835] = a[13] & g[9643];
assign g[26026] = b[13] & g[9643];
assign g[17836] = a[13] & g[9644];
assign g[26027] = b[13] & g[9644];
assign g[17837] = a[13] & g[9645];
assign g[26028] = b[13] & g[9645];
assign g[17838] = a[13] & g[9646];
assign g[26029] = b[13] & g[9646];
assign g[17839] = a[13] & g[9647];
assign g[26030] = b[13] & g[9647];
assign g[17840] = a[13] & g[9648];
assign g[26031] = b[13] & g[9648];
assign g[17841] = a[13] & g[9649];
assign g[26032] = b[13] & g[9649];
assign g[17842] = a[13] & g[9650];
assign g[26033] = b[13] & g[9650];
assign g[17843] = a[13] & g[9651];
assign g[26034] = b[13] & g[9651];
assign g[17844] = a[13] & g[9652];
assign g[26035] = b[13] & g[9652];
assign g[17845] = a[13] & g[9653];
assign g[26036] = b[13] & g[9653];
assign g[17846] = a[13] & g[9654];
assign g[26037] = b[13] & g[9654];
assign g[17847] = a[13] & g[9655];
assign g[26038] = b[13] & g[9655];
assign g[17848] = a[13] & g[9656];
assign g[26039] = b[13] & g[9656];
assign g[17849] = a[13] & g[9657];
assign g[26040] = b[13] & g[9657];
assign g[17850] = a[13] & g[9658];
assign g[26041] = b[13] & g[9658];
assign g[17851] = a[13] & g[9659];
assign g[26042] = b[13] & g[9659];
assign g[17852] = a[13] & g[9660];
assign g[26043] = b[13] & g[9660];
assign g[17853] = a[13] & g[9661];
assign g[26044] = b[13] & g[9661];
assign g[17854] = a[13] & g[9662];
assign g[26045] = b[13] & g[9662];
assign g[17855] = a[13] & g[9663];
assign g[26046] = b[13] & g[9663];
assign g[17856] = a[13] & g[9664];
assign g[26047] = b[13] & g[9664];
assign g[17857] = a[13] & g[9665];
assign g[26048] = b[13] & g[9665];
assign g[17858] = a[13] & g[9666];
assign g[26049] = b[13] & g[9666];
assign g[17859] = a[13] & g[9667];
assign g[26050] = b[13] & g[9667];
assign g[17860] = a[13] & g[9668];
assign g[26051] = b[13] & g[9668];
assign g[17861] = a[13] & g[9669];
assign g[26052] = b[13] & g[9669];
assign g[17862] = a[13] & g[9670];
assign g[26053] = b[13] & g[9670];
assign g[17863] = a[13] & g[9671];
assign g[26054] = b[13] & g[9671];
assign g[17864] = a[13] & g[9672];
assign g[26055] = b[13] & g[9672];
assign g[17865] = a[13] & g[9673];
assign g[26056] = b[13] & g[9673];
assign g[17866] = a[13] & g[9674];
assign g[26057] = b[13] & g[9674];
assign g[17867] = a[13] & g[9675];
assign g[26058] = b[13] & g[9675];
assign g[17868] = a[13] & g[9676];
assign g[26059] = b[13] & g[9676];
assign g[17869] = a[13] & g[9677];
assign g[26060] = b[13] & g[9677];
assign g[17870] = a[13] & g[9678];
assign g[26061] = b[13] & g[9678];
assign g[17871] = a[13] & g[9679];
assign g[26062] = b[13] & g[9679];
assign g[17872] = a[13] & g[9680];
assign g[26063] = b[13] & g[9680];
assign g[17873] = a[13] & g[9681];
assign g[26064] = b[13] & g[9681];
assign g[17874] = a[13] & g[9682];
assign g[26065] = b[13] & g[9682];
assign g[17875] = a[13] & g[9683];
assign g[26066] = b[13] & g[9683];
assign g[17876] = a[13] & g[9684];
assign g[26067] = b[13] & g[9684];
assign g[17877] = a[13] & g[9685];
assign g[26068] = b[13] & g[9685];
assign g[17878] = a[13] & g[9686];
assign g[26069] = b[13] & g[9686];
assign g[17879] = a[13] & g[9687];
assign g[26070] = b[13] & g[9687];
assign g[17880] = a[13] & g[9688];
assign g[26071] = b[13] & g[9688];
assign g[17881] = a[13] & g[9689];
assign g[26072] = b[13] & g[9689];
assign g[17882] = a[13] & g[9690];
assign g[26073] = b[13] & g[9690];
assign g[17883] = a[13] & g[9691];
assign g[26074] = b[13] & g[9691];
assign g[17884] = a[13] & g[9692];
assign g[26075] = b[13] & g[9692];
assign g[17885] = a[13] & g[9693];
assign g[26076] = b[13] & g[9693];
assign g[17886] = a[13] & g[9694];
assign g[26077] = b[13] & g[9694];
assign g[17887] = a[13] & g[9695];
assign g[26078] = b[13] & g[9695];
assign g[17888] = a[13] & g[9696];
assign g[26079] = b[13] & g[9696];
assign g[17889] = a[13] & g[9697];
assign g[26080] = b[13] & g[9697];
assign g[17890] = a[13] & g[9698];
assign g[26081] = b[13] & g[9698];
assign g[17891] = a[13] & g[9699];
assign g[26082] = b[13] & g[9699];
assign g[17892] = a[13] & g[9700];
assign g[26083] = b[13] & g[9700];
assign g[17893] = a[13] & g[9701];
assign g[26084] = b[13] & g[9701];
assign g[17894] = a[13] & g[9702];
assign g[26085] = b[13] & g[9702];
assign g[17895] = a[13] & g[9703];
assign g[26086] = b[13] & g[9703];
assign g[17896] = a[13] & g[9704];
assign g[26087] = b[13] & g[9704];
assign g[17897] = a[13] & g[9705];
assign g[26088] = b[13] & g[9705];
assign g[17898] = a[13] & g[9706];
assign g[26089] = b[13] & g[9706];
assign g[17899] = a[13] & g[9707];
assign g[26090] = b[13] & g[9707];
assign g[17900] = a[13] & g[9708];
assign g[26091] = b[13] & g[9708];
assign g[17901] = a[13] & g[9709];
assign g[26092] = b[13] & g[9709];
assign g[17902] = a[13] & g[9710];
assign g[26093] = b[13] & g[9710];
assign g[17903] = a[13] & g[9711];
assign g[26094] = b[13] & g[9711];
assign g[17904] = a[13] & g[9712];
assign g[26095] = b[13] & g[9712];
assign g[17905] = a[13] & g[9713];
assign g[26096] = b[13] & g[9713];
assign g[17906] = a[13] & g[9714];
assign g[26097] = b[13] & g[9714];
assign g[17907] = a[13] & g[9715];
assign g[26098] = b[13] & g[9715];
assign g[17908] = a[13] & g[9716];
assign g[26099] = b[13] & g[9716];
assign g[17909] = a[13] & g[9717];
assign g[26100] = b[13] & g[9717];
assign g[17910] = a[13] & g[9718];
assign g[26101] = b[13] & g[9718];
assign g[17911] = a[13] & g[9719];
assign g[26102] = b[13] & g[9719];
assign g[17912] = a[13] & g[9720];
assign g[26103] = b[13] & g[9720];
assign g[17913] = a[13] & g[9721];
assign g[26104] = b[13] & g[9721];
assign g[17914] = a[13] & g[9722];
assign g[26105] = b[13] & g[9722];
assign g[17915] = a[13] & g[9723];
assign g[26106] = b[13] & g[9723];
assign g[17916] = a[13] & g[9724];
assign g[26107] = b[13] & g[9724];
assign g[17917] = a[13] & g[9725];
assign g[26108] = b[13] & g[9725];
assign g[17918] = a[13] & g[9726];
assign g[26109] = b[13] & g[9726];
assign g[17919] = a[13] & g[9727];
assign g[26110] = b[13] & g[9727];
assign g[17920] = a[13] & g[9728];
assign g[26111] = b[13] & g[9728];
assign g[17921] = a[13] & g[9729];
assign g[26112] = b[13] & g[9729];
assign g[17922] = a[13] & g[9730];
assign g[26113] = b[13] & g[9730];
assign g[17923] = a[13] & g[9731];
assign g[26114] = b[13] & g[9731];
assign g[17924] = a[13] & g[9732];
assign g[26115] = b[13] & g[9732];
assign g[17925] = a[13] & g[9733];
assign g[26116] = b[13] & g[9733];
assign g[17926] = a[13] & g[9734];
assign g[26117] = b[13] & g[9734];
assign g[17927] = a[13] & g[9735];
assign g[26118] = b[13] & g[9735];
assign g[17928] = a[13] & g[9736];
assign g[26119] = b[13] & g[9736];
assign g[17929] = a[13] & g[9737];
assign g[26120] = b[13] & g[9737];
assign g[17930] = a[13] & g[9738];
assign g[26121] = b[13] & g[9738];
assign g[17931] = a[13] & g[9739];
assign g[26122] = b[13] & g[9739];
assign g[17932] = a[13] & g[9740];
assign g[26123] = b[13] & g[9740];
assign g[17933] = a[13] & g[9741];
assign g[26124] = b[13] & g[9741];
assign g[17934] = a[13] & g[9742];
assign g[26125] = b[13] & g[9742];
assign g[17935] = a[13] & g[9743];
assign g[26126] = b[13] & g[9743];
assign g[17936] = a[13] & g[9744];
assign g[26127] = b[13] & g[9744];
assign g[17937] = a[13] & g[9745];
assign g[26128] = b[13] & g[9745];
assign g[17938] = a[13] & g[9746];
assign g[26129] = b[13] & g[9746];
assign g[17939] = a[13] & g[9747];
assign g[26130] = b[13] & g[9747];
assign g[17940] = a[13] & g[9748];
assign g[26131] = b[13] & g[9748];
assign g[17941] = a[13] & g[9749];
assign g[26132] = b[13] & g[9749];
assign g[17942] = a[13] & g[9750];
assign g[26133] = b[13] & g[9750];
assign g[17943] = a[13] & g[9751];
assign g[26134] = b[13] & g[9751];
assign g[17944] = a[13] & g[9752];
assign g[26135] = b[13] & g[9752];
assign g[17945] = a[13] & g[9753];
assign g[26136] = b[13] & g[9753];
assign g[17946] = a[13] & g[9754];
assign g[26137] = b[13] & g[9754];
assign g[17947] = a[13] & g[9755];
assign g[26138] = b[13] & g[9755];
assign g[17948] = a[13] & g[9756];
assign g[26139] = b[13] & g[9756];
assign g[17949] = a[13] & g[9757];
assign g[26140] = b[13] & g[9757];
assign g[17950] = a[13] & g[9758];
assign g[26141] = b[13] & g[9758];
assign g[17951] = a[13] & g[9759];
assign g[26142] = b[13] & g[9759];
assign g[17952] = a[13] & g[9760];
assign g[26143] = b[13] & g[9760];
assign g[17953] = a[13] & g[9761];
assign g[26144] = b[13] & g[9761];
assign g[17954] = a[13] & g[9762];
assign g[26145] = b[13] & g[9762];
assign g[17955] = a[13] & g[9763];
assign g[26146] = b[13] & g[9763];
assign g[17956] = a[13] & g[9764];
assign g[26147] = b[13] & g[9764];
assign g[17957] = a[13] & g[9765];
assign g[26148] = b[13] & g[9765];
assign g[17958] = a[13] & g[9766];
assign g[26149] = b[13] & g[9766];
assign g[17959] = a[13] & g[9767];
assign g[26150] = b[13] & g[9767];
assign g[17960] = a[13] & g[9768];
assign g[26151] = b[13] & g[9768];
assign g[17961] = a[13] & g[9769];
assign g[26152] = b[13] & g[9769];
assign g[17962] = a[13] & g[9770];
assign g[26153] = b[13] & g[9770];
assign g[17963] = a[13] & g[9771];
assign g[26154] = b[13] & g[9771];
assign g[17964] = a[13] & g[9772];
assign g[26155] = b[13] & g[9772];
assign g[17965] = a[13] & g[9773];
assign g[26156] = b[13] & g[9773];
assign g[17966] = a[13] & g[9774];
assign g[26157] = b[13] & g[9774];
assign g[17967] = a[13] & g[9775];
assign g[26158] = b[13] & g[9775];
assign g[17968] = a[13] & g[9776];
assign g[26159] = b[13] & g[9776];
assign g[17969] = a[13] & g[9777];
assign g[26160] = b[13] & g[9777];
assign g[17970] = a[13] & g[9778];
assign g[26161] = b[13] & g[9778];
assign g[17971] = a[13] & g[9779];
assign g[26162] = b[13] & g[9779];
assign g[17972] = a[13] & g[9780];
assign g[26163] = b[13] & g[9780];
assign g[17973] = a[13] & g[9781];
assign g[26164] = b[13] & g[9781];
assign g[17974] = a[13] & g[9782];
assign g[26165] = b[13] & g[9782];
assign g[17975] = a[13] & g[9783];
assign g[26166] = b[13] & g[9783];
assign g[17976] = a[13] & g[9784];
assign g[26167] = b[13] & g[9784];
assign g[17977] = a[13] & g[9785];
assign g[26168] = b[13] & g[9785];
assign g[17978] = a[13] & g[9786];
assign g[26169] = b[13] & g[9786];
assign g[17979] = a[13] & g[9787];
assign g[26170] = b[13] & g[9787];
assign g[17980] = a[13] & g[9788];
assign g[26171] = b[13] & g[9788];
assign g[17981] = a[13] & g[9789];
assign g[26172] = b[13] & g[9789];
assign g[17982] = a[13] & g[9790];
assign g[26173] = b[13] & g[9790];
assign g[17983] = a[13] & g[9791];
assign g[26174] = b[13] & g[9791];
assign g[17984] = a[13] & g[9792];
assign g[26175] = b[13] & g[9792];
assign g[17985] = a[13] & g[9793];
assign g[26176] = b[13] & g[9793];
assign g[17986] = a[13] & g[9794];
assign g[26177] = b[13] & g[9794];
assign g[17987] = a[13] & g[9795];
assign g[26178] = b[13] & g[9795];
assign g[17988] = a[13] & g[9796];
assign g[26179] = b[13] & g[9796];
assign g[17989] = a[13] & g[9797];
assign g[26180] = b[13] & g[9797];
assign g[17990] = a[13] & g[9798];
assign g[26181] = b[13] & g[9798];
assign g[17991] = a[13] & g[9799];
assign g[26182] = b[13] & g[9799];
assign g[17992] = a[13] & g[9800];
assign g[26183] = b[13] & g[9800];
assign g[17993] = a[13] & g[9801];
assign g[26184] = b[13] & g[9801];
assign g[17994] = a[13] & g[9802];
assign g[26185] = b[13] & g[9802];
assign g[17995] = a[13] & g[9803];
assign g[26186] = b[13] & g[9803];
assign g[17996] = a[13] & g[9804];
assign g[26187] = b[13] & g[9804];
assign g[17997] = a[13] & g[9805];
assign g[26188] = b[13] & g[9805];
assign g[17998] = a[13] & g[9806];
assign g[26189] = b[13] & g[9806];
assign g[17999] = a[13] & g[9807];
assign g[26190] = b[13] & g[9807];
assign g[18000] = a[13] & g[9808];
assign g[26191] = b[13] & g[9808];
assign g[18001] = a[13] & g[9809];
assign g[26192] = b[13] & g[9809];
assign g[18002] = a[13] & g[9810];
assign g[26193] = b[13] & g[9810];
assign g[18003] = a[13] & g[9811];
assign g[26194] = b[13] & g[9811];
assign g[18004] = a[13] & g[9812];
assign g[26195] = b[13] & g[9812];
assign g[18005] = a[13] & g[9813];
assign g[26196] = b[13] & g[9813];
assign g[18006] = a[13] & g[9814];
assign g[26197] = b[13] & g[9814];
assign g[18007] = a[13] & g[9815];
assign g[26198] = b[13] & g[9815];
assign g[18008] = a[13] & g[9816];
assign g[26199] = b[13] & g[9816];
assign g[18009] = a[13] & g[9817];
assign g[26200] = b[13] & g[9817];
assign g[18010] = a[13] & g[9818];
assign g[26201] = b[13] & g[9818];
assign g[18011] = a[13] & g[9819];
assign g[26202] = b[13] & g[9819];
assign g[18012] = a[13] & g[9820];
assign g[26203] = b[13] & g[9820];
assign g[18013] = a[13] & g[9821];
assign g[26204] = b[13] & g[9821];
assign g[18014] = a[13] & g[9822];
assign g[26205] = b[13] & g[9822];
assign g[18015] = a[13] & g[9823];
assign g[26206] = b[13] & g[9823];
assign g[18016] = a[13] & g[9824];
assign g[26207] = b[13] & g[9824];
assign g[18017] = a[13] & g[9825];
assign g[26208] = b[13] & g[9825];
assign g[18018] = a[13] & g[9826];
assign g[26209] = b[13] & g[9826];
assign g[18019] = a[13] & g[9827];
assign g[26210] = b[13] & g[9827];
assign g[18020] = a[13] & g[9828];
assign g[26211] = b[13] & g[9828];
assign g[18021] = a[13] & g[9829];
assign g[26212] = b[13] & g[9829];
assign g[18022] = a[13] & g[9830];
assign g[26213] = b[13] & g[9830];
assign g[18023] = a[13] & g[9831];
assign g[26214] = b[13] & g[9831];
assign g[18024] = a[13] & g[9832];
assign g[26215] = b[13] & g[9832];
assign g[18025] = a[13] & g[9833];
assign g[26216] = b[13] & g[9833];
assign g[18026] = a[13] & g[9834];
assign g[26217] = b[13] & g[9834];
assign g[18027] = a[13] & g[9835];
assign g[26218] = b[13] & g[9835];
assign g[18028] = a[13] & g[9836];
assign g[26219] = b[13] & g[9836];
assign g[18029] = a[13] & g[9837];
assign g[26220] = b[13] & g[9837];
assign g[18030] = a[13] & g[9838];
assign g[26221] = b[13] & g[9838];
assign g[18031] = a[13] & g[9839];
assign g[26222] = b[13] & g[9839];
assign g[18032] = a[13] & g[9840];
assign g[26223] = b[13] & g[9840];
assign g[18033] = a[13] & g[9841];
assign g[26224] = b[13] & g[9841];
assign g[18034] = a[13] & g[9842];
assign g[26225] = b[13] & g[9842];
assign g[18035] = a[13] & g[9843];
assign g[26226] = b[13] & g[9843];
assign g[18036] = a[13] & g[9844];
assign g[26227] = b[13] & g[9844];
assign g[18037] = a[13] & g[9845];
assign g[26228] = b[13] & g[9845];
assign g[18038] = a[13] & g[9846];
assign g[26229] = b[13] & g[9846];
assign g[18039] = a[13] & g[9847];
assign g[26230] = b[13] & g[9847];
assign g[18040] = a[13] & g[9848];
assign g[26231] = b[13] & g[9848];
assign g[18041] = a[13] & g[9849];
assign g[26232] = b[13] & g[9849];
assign g[18042] = a[13] & g[9850];
assign g[26233] = b[13] & g[9850];
assign g[18043] = a[13] & g[9851];
assign g[26234] = b[13] & g[9851];
assign g[18044] = a[13] & g[9852];
assign g[26235] = b[13] & g[9852];
assign g[18045] = a[13] & g[9853];
assign g[26236] = b[13] & g[9853];
assign g[18046] = a[13] & g[9854];
assign g[26237] = b[13] & g[9854];
assign g[18047] = a[13] & g[9855];
assign g[26238] = b[13] & g[9855];
assign g[18048] = a[13] & g[9856];
assign g[26239] = b[13] & g[9856];
assign g[18049] = a[13] & g[9857];
assign g[26240] = b[13] & g[9857];
assign g[18050] = a[13] & g[9858];
assign g[26241] = b[13] & g[9858];
assign g[18051] = a[13] & g[9859];
assign g[26242] = b[13] & g[9859];
assign g[18052] = a[13] & g[9860];
assign g[26243] = b[13] & g[9860];
assign g[18053] = a[13] & g[9861];
assign g[26244] = b[13] & g[9861];
assign g[18054] = a[13] & g[9862];
assign g[26245] = b[13] & g[9862];
assign g[18055] = a[13] & g[9863];
assign g[26246] = b[13] & g[9863];
assign g[18056] = a[13] & g[9864];
assign g[26247] = b[13] & g[9864];
assign g[18057] = a[13] & g[9865];
assign g[26248] = b[13] & g[9865];
assign g[18058] = a[13] & g[9866];
assign g[26249] = b[13] & g[9866];
assign g[18059] = a[13] & g[9867];
assign g[26250] = b[13] & g[9867];
assign g[18060] = a[13] & g[9868];
assign g[26251] = b[13] & g[9868];
assign g[18061] = a[13] & g[9869];
assign g[26252] = b[13] & g[9869];
assign g[18062] = a[13] & g[9870];
assign g[26253] = b[13] & g[9870];
assign g[18063] = a[13] & g[9871];
assign g[26254] = b[13] & g[9871];
assign g[18064] = a[13] & g[9872];
assign g[26255] = b[13] & g[9872];
assign g[18065] = a[13] & g[9873];
assign g[26256] = b[13] & g[9873];
assign g[18066] = a[13] & g[9874];
assign g[26257] = b[13] & g[9874];
assign g[18067] = a[13] & g[9875];
assign g[26258] = b[13] & g[9875];
assign g[18068] = a[13] & g[9876];
assign g[26259] = b[13] & g[9876];
assign g[18069] = a[13] & g[9877];
assign g[26260] = b[13] & g[9877];
assign g[18070] = a[13] & g[9878];
assign g[26261] = b[13] & g[9878];
assign g[18071] = a[13] & g[9879];
assign g[26262] = b[13] & g[9879];
assign g[18072] = a[13] & g[9880];
assign g[26263] = b[13] & g[9880];
assign g[18073] = a[13] & g[9881];
assign g[26264] = b[13] & g[9881];
assign g[18074] = a[13] & g[9882];
assign g[26265] = b[13] & g[9882];
assign g[18075] = a[13] & g[9883];
assign g[26266] = b[13] & g[9883];
assign g[18076] = a[13] & g[9884];
assign g[26267] = b[13] & g[9884];
assign g[18077] = a[13] & g[9885];
assign g[26268] = b[13] & g[9885];
assign g[18078] = a[13] & g[9886];
assign g[26269] = b[13] & g[9886];
assign g[18079] = a[13] & g[9887];
assign g[26270] = b[13] & g[9887];
assign g[18080] = a[13] & g[9888];
assign g[26271] = b[13] & g[9888];
assign g[18081] = a[13] & g[9889];
assign g[26272] = b[13] & g[9889];
assign g[18082] = a[13] & g[9890];
assign g[26273] = b[13] & g[9890];
assign g[18083] = a[13] & g[9891];
assign g[26274] = b[13] & g[9891];
assign g[18084] = a[13] & g[9892];
assign g[26275] = b[13] & g[9892];
assign g[18085] = a[13] & g[9893];
assign g[26276] = b[13] & g[9893];
assign g[18086] = a[13] & g[9894];
assign g[26277] = b[13] & g[9894];
assign g[18087] = a[13] & g[9895];
assign g[26278] = b[13] & g[9895];
assign g[18088] = a[13] & g[9896];
assign g[26279] = b[13] & g[9896];
assign g[18089] = a[13] & g[9897];
assign g[26280] = b[13] & g[9897];
assign g[18090] = a[13] & g[9898];
assign g[26281] = b[13] & g[9898];
assign g[18091] = a[13] & g[9899];
assign g[26282] = b[13] & g[9899];
assign g[18092] = a[13] & g[9900];
assign g[26283] = b[13] & g[9900];
assign g[18093] = a[13] & g[9901];
assign g[26284] = b[13] & g[9901];
assign g[18094] = a[13] & g[9902];
assign g[26285] = b[13] & g[9902];
assign g[18095] = a[13] & g[9903];
assign g[26286] = b[13] & g[9903];
assign g[18096] = a[13] & g[9904];
assign g[26287] = b[13] & g[9904];
assign g[18097] = a[13] & g[9905];
assign g[26288] = b[13] & g[9905];
assign g[18098] = a[13] & g[9906];
assign g[26289] = b[13] & g[9906];
assign g[18099] = a[13] & g[9907];
assign g[26290] = b[13] & g[9907];
assign g[18100] = a[13] & g[9908];
assign g[26291] = b[13] & g[9908];
assign g[18101] = a[13] & g[9909];
assign g[26292] = b[13] & g[9909];
assign g[18102] = a[13] & g[9910];
assign g[26293] = b[13] & g[9910];
assign g[18103] = a[13] & g[9911];
assign g[26294] = b[13] & g[9911];
assign g[18104] = a[13] & g[9912];
assign g[26295] = b[13] & g[9912];
assign g[18105] = a[13] & g[9913];
assign g[26296] = b[13] & g[9913];
assign g[18106] = a[13] & g[9914];
assign g[26297] = b[13] & g[9914];
assign g[18107] = a[13] & g[9915];
assign g[26298] = b[13] & g[9915];
assign g[18108] = a[13] & g[9916];
assign g[26299] = b[13] & g[9916];
assign g[18109] = a[13] & g[9917];
assign g[26300] = b[13] & g[9917];
assign g[18110] = a[13] & g[9918];
assign g[26301] = b[13] & g[9918];
assign g[18111] = a[13] & g[9919];
assign g[26302] = b[13] & g[9919];
assign g[18112] = a[13] & g[9920];
assign g[26303] = b[13] & g[9920];
assign g[18113] = a[13] & g[9921];
assign g[26304] = b[13] & g[9921];
assign g[18114] = a[13] & g[9922];
assign g[26305] = b[13] & g[9922];
assign g[18115] = a[13] & g[9923];
assign g[26306] = b[13] & g[9923];
assign g[18116] = a[13] & g[9924];
assign g[26307] = b[13] & g[9924];
assign g[18117] = a[13] & g[9925];
assign g[26308] = b[13] & g[9925];
assign g[18118] = a[13] & g[9926];
assign g[26309] = b[13] & g[9926];
assign g[18119] = a[13] & g[9927];
assign g[26310] = b[13] & g[9927];
assign g[18120] = a[13] & g[9928];
assign g[26311] = b[13] & g[9928];
assign g[18121] = a[13] & g[9929];
assign g[26312] = b[13] & g[9929];
assign g[18122] = a[13] & g[9930];
assign g[26313] = b[13] & g[9930];
assign g[18123] = a[13] & g[9931];
assign g[26314] = b[13] & g[9931];
assign g[18124] = a[13] & g[9932];
assign g[26315] = b[13] & g[9932];
assign g[18125] = a[13] & g[9933];
assign g[26316] = b[13] & g[9933];
assign g[18126] = a[13] & g[9934];
assign g[26317] = b[13] & g[9934];
assign g[18127] = a[13] & g[9935];
assign g[26318] = b[13] & g[9935];
assign g[18128] = a[13] & g[9936];
assign g[26319] = b[13] & g[9936];
assign g[18129] = a[13] & g[9937];
assign g[26320] = b[13] & g[9937];
assign g[18130] = a[13] & g[9938];
assign g[26321] = b[13] & g[9938];
assign g[18131] = a[13] & g[9939];
assign g[26322] = b[13] & g[9939];
assign g[18132] = a[13] & g[9940];
assign g[26323] = b[13] & g[9940];
assign g[18133] = a[13] & g[9941];
assign g[26324] = b[13] & g[9941];
assign g[18134] = a[13] & g[9942];
assign g[26325] = b[13] & g[9942];
assign g[18135] = a[13] & g[9943];
assign g[26326] = b[13] & g[9943];
assign g[18136] = a[13] & g[9944];
assign g[26327] = b[13] & g[9944];
assign g[18137] = a[13] & g[9945];
assign g[26328] = b[13] & g[9945];
assign g[18138] = a[13] & g[9946];
assign g[26329] = b[13] & g[9946];
assign g[18139] = a[13] & g[9947];
assign g[26330] = b[13] & g[9947];
assign g[18140] = a[13] & g[9948];
assign g[26331] = b[13] & g[9948];
assign g[18141] = a[13] & g[9949];
assign g[26332] = b[13] & g[9949];
assign g[18142] = a[13] & g[9950];
assign g[26333] = b[13] & g[9950];
assign g[18143] = a[13] & g[9951];
assign g[26334] = b[13] & g[9951];
assign g[18144] = a[13] & g[9952];
assign g[26335] = b[13] & g[9952];
assign g[18145] = a[13] & g[9953];
assign g[26336] = b[13] & g[9953];
assign g[18146] = a[13] & g[9954];
assign g[26337] = b[13] & g[9954];
assign g[18147] = a[13] & g[9955];
assign g[26338] = b[13] & g[9955];
assign g[18148] = a[13] & g[9956];
assign g[26339] = b[13] & g[9956];
assign g[18149] = a[13] & g[9957];
assign g[26340] = b[13] & g[9957];
assign g[18150] = a[13] & g[9958];
assign g[26341] = b[13] & g[9958];
assign g[18151] = a[13] & g[9959];
assign g[26342] = b[13] & g[9959];
assign g[18152] = a[13] & g[9960];
assign g[26343] = b[13] & g[9960];
assign g[18153] = a[13] & g[9961];
assign g[26344] = b[13] & g[9961];
assign g[18154] = a[13] & g[9962];
assign g[26345] = b[13] & g[9962];
assign g[18155] = a[13] & g[9963];
assign g[26346] = b[13] & g[9963];
assign g[18156] = a[13] & g[9964];
assign g[26347] = b[13] & g[9964];
assign g[18157] = a[13] & g[9965];
assign g[26348] = b[13] & g[9965];
assign g[18158] = a[13] & g[9966];
assign g[26349] = b[13] & g[9966];
assign g[18159] = a[13] & g[9967];
assign g[26350] = b[13] & g[9967];
assign g[18160] = a[13] & g[9968];
assign g[26351] = b[13] & g[9968];
assign g[18161] = a[13] & g[9969];
assign g[26352] = b[13] & g[9969];
assign g[18162] = a[13] & g[9970];
assign g[26353] = b[13] & g[9970];
assign g[18163] = a[13] & g[9971];
assign g[26354] = b[13] & g[9971];
assign g[18164] = a[13] & g[9972];
assign g[26355] = b[13] & g[9972];
assign g[18165] = a[13] & g[9973];
assign g[26356] = b[13] & g[9973];
assign g[18166] = a[13] & g[9974];
assign g[26357] = b[13] & g[9974];
assign g[18167] = a[13] & g[9975];
assign g[26358] = b[13] & g[9975];
assign g[18168] = a[13] & g[9976];
assign g[26359] = b[13] & g[9976];
assign g[18169] = a[13] & g[9977];
assign g[26360] = b[13] & g[9977];
assign g[18170] = a[13] & g[9978];
assign g[26361] = b[13] & g[9978];
assign g[18171] = a[13] & g[9979];
assign g[26362] = b[13] & g[9979];
assign g[18172] = a[13] & g[9980];
assign g[26363] = b[13] & g[9980];
assign g[18173] = a[13] & g[9981];
assign g[26364] = b[13] & g[9981];
assign g[18174] = a[13] & g[9982];
assign g[26365] = b[13] & g[9982];
assign g[18175] = a[13] & g[9983];
assign g[26366] = b[13] & g[9983];
assign g[18176] = a[13] & g[9984];
assign g[26367] = b[13] & g[9984];
assign g[18177] = a[13] & g[9985];
assign g[26368] = b[13] & g[9985];
assign g[18178] = a[13] & g[9986];
assign g[26369] = b[13] & g[9986];
assign g[18179] = a[13] & g[9987];
assign g[26370] = b[13] & g[9987];
assign g[18180] = a[13] & g[9988];
assign g[26371] = b[13] & g[9988];
assign g[18181] = a[13] & g[9989];
assign g[26372] = b[13] & g[9989];
assign g[18182] = a[13] & g[9990];
assign g[26373] = b[13] & g[9990];
assign g[18183] = a[13] & g[9991];
assign g[26374] = b[13] & g[9991];
assign g[18184] = a[13] & g[9992];
assign g[26375] = b[13] & g[9992];
assign g[18185] = a[13] & g[9993];
assign g[26376] = b[13] & g[9993];
assign g[18186] = a[13] & g[9994];
assign g[26377] = b[13] & g[9994];
assign g[18187] = a[13] & g[9995];
assign g[26378] = b[13] & g[9995];
assign g[18188] = a[13] & g[9996];
assign g[26379] = b[13] & g[9996];
assign g[18189] = a[13] & g[9997];
assign g[26380] = b[13] & g[9997];
assign g[18190] = a[13] & g[9998];
assign g[26381] = b[13] & g[9998];
assign g[18191] = a[13] & g[9999];
assign g[26382] = b[13] & g[9999];
assign g[18192] = a[13] & g[10000];
assign g[26383] = b[13] & g[10000];
assign g[18193] = a[13] & g[10001];
assign g[26384] = b[13] & g[10001];
assign g[18194] = a[13] & g[10002];
assign g[26385] = b[13] & g[10002];
assign g[18195] = a[13] & g[10003];
assign g[26386] = b[13] & g[10003];
assign g[18196] = a[13] & g[10004];
assign g[26387] = b[13] & g[10004];
assign g[18197] = a[13] & g[10005];
assign g[26388] = b[13] & g[10005];
assign g[18198] = a[13] & g[10006];
assign g[26389] = b[13] & g[10006];
assign g[18199] = a[13] & g[10007];
assign g[26390] = b[13] & g[10007];
assign g[18200] = a[13] & g[10008];
assign g[26391] = b[13] & g[10008];
assign g[18201] = a[13] & g[10009];
assign g[26392] = b[13] & g[10009];
assign g[18202] = a[13] & g[10010];
assign g[26393] = b[13] & g[10010];
assign g[18203] = a[13] & g[10011];
assign g[26394] = b[13] & g[10011];
assign g[18204] = a[13] & g[10012];
assign g[26395] = b[13] & g[10012];
assign g[18205] = a[13] & g[10013];
assign g[26396] = b[13] & g[10013];
assign g[18206] = a[13] & g[10014];
assign g[26397] = b[13] & g[10014];
assign g[18207] = a[13] & g[10015];
assign g[26398] = b[13] & g[10015];
assign g[18208] = a[13] & g[10016];
assign g[26399] = b[13] & g[10016];
assign g[18209] = a[13] & g[10017];
assign g[26400] = b[13] & g[10017];
assign g[18210] = a[13] & g[10018];
assign g[26401] = b[13] & g[10018];
assign g[18211] = a[13] & g[10019];
assign g[26402] = b[13] & g[10019];
assign g[18212] = a[13] & g[10020];
assign g[26403] = b[13] & g[10020];
assign g[18213] = a[13] & g[10021];
assign g[26404] = b[13] & g[10021];
assign g[18214] = a[13] & g[10022];
assign g[26405] = b[13] & g[10022];
assign g[18215] = a[13] & g[10023];
assign g[26406] = b[13] & g[10023];
assign g[18216] = a[13] & g[10024];
assign g[26407] = b[13] & g[10024];
assign g[18217] = a[13] & g[10025];
assign g[26408] = b[13] & g[10025];
assign g[18218] = a[13] & g[10026];
assign g[26409] = b[13] & g[10026];
assign g[18219] = a[13] & g[10027];
assign g[26410] = b[13] & g[10027];
assign g[18220] = a[13] & g[10028];
assign g[26411] = b[13] & g[10028];
assign g[18221] = a[13] & g[10029];
assign g[26412] = b[13] & g[10029];
assign g[18222] = a[13] & g[10030];
assign g[26413] = b[13] & g[10030];
assign g[18223] = a[13] & g[10031];
assign g[26414] = b[13] & g[10031];
assign g[18224] = a[13] & g[10032];
assign g[26415] = b[13] & g[10032];
assign g[18225] = a[13] & g[10033];
assign g[26416] = b[13] & g[10033];
assign g[18226] = a[13] & g[10034];
assign g[26417] = b[13] & g[10034];
assign g[18227] = a[13] & g[10035];
assign g[26418] = b[13] & g[10035];
assign g[18228] = a[13] & g[10036];
assign g[26419] = b[13] & g[10036];
assign g[18229] = a[13] & g[10037];
assign g[26420] = b[13] & g[10037];
assign g[18230] = a[13] & g[10038];
assign g[26421] = b[13] & g[10038];
assign g[18231] = a[13] & g[10039];
assign g[26422] = b[13] & g[10039];
assign g[18232] = a[13] & g[10040];
assign g[26423] = b[13] & g[10040];
assign g[18233] = a[13] & g[10041];
assign g[26424] = b[13] & g[10041];
assign g[18234] = a[13] & g[10042];
assign g[26425] = b[13] & g[10042];
assign g[18235] = a[13] & g[10043];
assign g[26426] = b[13] & g[10043];
assign g[18236] = a[13] & g[10044];
assign g[26427] = b[13] & g[10044];
assign g[18237] = a[13] & g[10045];
assign g[26428] = b[13] & g[10045];
assign g[18238] = a[13] & g[10046];
assign g[26429] = b[13] & g[10046];
assign g[18239] = a[13] & g[10047];
assign g[26430] = b[13] & g[10047];
assign g[18240] = a[13] & g[10048];
assign g[26431] = b[13] & g[10048];
assign g[18241] = a[13] & g[10049];
assign g[26432] = b[13] & g[10049];
assign g[18242] = a[13] & g[10050];
assign g[26433] = b[13] & g[10050];
assign g[18243] = a[13] & g[10051];
assign g[26434] = b[13] & g[10051];
assign g[18244] = a[13] & g[10052];
assign g[26435] = b[13] & g[10052];
assign g[18245] = a[13] & g[10053];
assign g[26436] = b[13] & g[10053];
assign g[18246] = a[13] & g[10054];
assign g[26437] = b[13] & g[10054];
assign g[18247] = a[13] & g[10055];
assign g[26438] = b[13] & g[10055];
assign g[18248] = a[13] & g[10056];
assign g[26439] = b[13] & g[10056];
assign g[18249] = a[13] & g[10057];
assign g[26440] = b[13] & g[10057];
assign g[18250] = a[13] & g[10058];
assign g[26441] = b[13] & g[10058];
assign g[18251] = a[13] & g[10059];
assign g[26442] = b[13] & g[10059];
assign g[18252] = a[13] & g[10060];
assign g[26443] = b[13] & g[10060];
assign g[18253] = a[13] & g[10061];
assign g[26444] = b[13] & g[10061];
assign g[18254] = a[13] & g[10062];
assign g[26445] = b[13] & g[10062];
assign g[18255] = a[13] & g[10063];
assign g[26446] = b[13] & g[10063];
assign g[18256] = a[13] & g[10064];
assign g[26447] = b[13] & g[10064];
assign g[18257] = a[13] & g[10065];
assign g[26448] = b[13] & g[10065];
assign g[18258] = a[13] & g[10066];
assign g[26449] = b[13] & g[10066];
assign g[18259] = a[13] & g[10067];
assign g[26450] = b[13] & g[10067];
assign g[18260] = a[13] & g[10068];
assign g[26451] = b[13] & g[10068];
assign g[18261] = a[13] & g[10069];
assign g[26452] = b[13] & g[10069];
assign g[18262] = a[13] & g[10070];
assign g[26453] = b[13] & g[10070];
assign g[18263] = a[13] & g[10071];
assign g[26454] = b[13] & g[10071];
assign g[18264] = a[13] & g[10072];
assign g[26455] = b[13] & g[10072];
assign g[18265] = a[13] & g[10073];
assign g[26456] = b[13] & g[10073];
assign g[18266] = a[13] & g[10074];
assign g[26457] = b[13] & g[10074];
assign g[18267] = a[13] & g[10075];
assign g[26458] = b[13] & g[10075];
assign g[18268] = a[13] & g[10076];
assign g[26459] = b[13] & g[10076];
assign g[18269] = a[13] & g[10077];
assign g[26460] = b[13] & g[10077];
assign g[18270] = a[13] & g[10078];
assign g[26461] = b[13] & g[10078];
assign g[18271] = a[13] & g[10079];
assign g[26462] = b[13] & g[10079];
assign g[18272] = a[13] & g[10080];
assign g[26463] = b[13] & g[10080];
assign g[18273] = a[13] & g[10081];
assign g[26464] = b[13] & g[10081];
assign g[18274] = a[13] & g[10082];
assign g[26465] = b[13] & g[10082];
assign g[18275] = a[13] & g[10083];
assign g[26466] = b[13] & g[10083];
assign g[18276] = a[13] & g[10084];
assign g[26467] = b[13] & g[10084];
assign g[18277] = a[13] & g[10085];
assign g[26468] = b[13] & g[10085];
assign g[18278] = a[13] & g[10086];
assign g[26469] = b[13] & g[10086];
assign g[18279] = a[13] & g[10087];
assign g[26470] = b[13] & g[10087];
assign g[18280] = a[13] & g[10088];
assign g[26471] = b[13] & g[10088];
assign g[18281] = a[13] & g[10089];
assign g[26472] = b[13] & g[10089];
assign g[18282] = a[13] & g[10090];
assign g[26473] = b[13] & g[10090];
assign g[18283] = a[13] & g[10091];
assign g[26474] = b[13] & g[10091];
assign g[18284] = a[13] & g[10092];
assign g[26475] = b[13] & g[10092];
assign g[18285] = a[13] & g[10093];
assign g[26476] = b[13] & g[10093];
assign g[18286] = a[13] & g[10094];
assign g[26477] = b[13] & g[10094];
assign g[18287] = a[13] & g[10095];
assign g[26478] = b[13] & g[10095];
assign g[18288] = a[13] & g[10096];
assign g[26479] = b[13] & g[10096];
assign g[18289] = a[13] & g[10097];
assign g[26480] = b[13] & g[10097];
assign g[18290] = a[13] & g[10098];
assign g[26481] = b[13] & g[10098];
assign g[18291] = a[13] & g[10099];
assign g[26482] = b[13] & g[10099];
assign g[18292] = a[13] & g[10100];
assign g[26483] = b[13] & g[10100];
assign g[18293] = a[13] & g[10101];
assign g[26484] = b[13] & g[10101];
assign g[18294] = a[13] & g[10102];
assign g[26485] = b[13] & g[10102];
assign g[18295] = a[13] & g[10103];
assign g[26486] = b[13] & g[10103];
assign g[18296] = a[13] & g[10104];
assign g[26487] = b[13] & g[10104];
assign g[18297] = a[13] & g[10105];
assign g[26488] = b[13] & g[10105];
assign g[18298] = a[13] & g[10106];
assign g[26489] = b[13] & g[10106];
assign g[18299] = a[13] & g[10107];
assign g[26490] = b[13] & g[10107];
assign g[18300] = a[13] & g[10108];
assign g[26491] = b[13] & g[10108];
assign g[18301] = a[13] & g[10109];
assign g[26492] = b[13] & g[10109];
assign g[18302] = a[13] & g[10110];
assign g[26493] = b[13] & g[10110];
assign g[18303] = a[13] & g[10111];
assign g[26494] = b[13] & g[10111];
assign g[18304] = a[13] & g[10112];
assign g[26495] = b[13] & g[10112];
assign g[18305] = a[13] & g[10113];
assign g[26496] = b[13] & g[10113];
assign g[18306] = a[13] & g[10114];
assign g[26497] = b[13] & g[10114];
assign g[18307] = a[13] & g[10115];
assign g[26498] = b[13] & g[10115];
assign g[18308] = a[13] & g[10116];
assign g[26499] = b[13] & g[10116];
assign g[18309] = a[13] & g[10117];
assign g[26500] = b[13] & g[10117];
assign g[18310] = a[13] & g[10118];
assign g[26501] = b[13] & g[10118];
assign g[18311] = a[13] & g[10119];
assign g[26502] = b[13] & g[10119];
assign g[18312] = a[13] & g[10120];
assign g[26503] = b[13] & g[10120];
assign g[18313] = a[13] & g[10121];
assign g[26504] = b[13] & g[10121];
assign g[18314] = a[13] & g[10122];
assign g[26505] = b[13] & g[10122];
assign g[18315] = a[13] & g[10123];
assign g[26506] = b[13] & g[10123];
assign g[18316] = a[13] & g[10124];
assign g[26507] = b[13] & g[10124];
assign g[18317] = a[13] & g[10125];
assign g[26508] = b[13] & g[10125];
assign g[18318] = a[13] & g[10126];
assign g[26509] = b[13] & g[10126];
assign g[18319] = a[13] & g[10127];
assign g[26510] = b[13] & g[10127];
assign g[18320] = a[13] & g[10128];
assign g[26511] = b[13] & g[10128];
assign g[18321] = a[13] & g[10129];
assign g[26512] = b[13] & g[10129];
assign g[18322] = a[13] & g[10130];
assign g[26513] = b[13] & g[10130];
assign g[18323] = a[13] & g[10131];
assign g[26514] = b[13] & g[10131];
assign g[18324] = a[13] & g[10132];
assign g[26515] = b[13] & g[10132];
assign g[18325] = a[13] & g[10133];
assign g[26516] = b[13] & g[10133];
assign g[18326] = a[13] & g[10134];
assign g[26517] = b[13] & g[10134];
assign g[18327] = a[13] & g[10135];
assign g[26518] = b[13] & g[10135];
assign g[18328] = a[13] & g[10136];
assign g[26519] = b[13] & g[10136];
assign g[18329] = a[13] & g[10137];
assign g[26520] = b[13] & g[10137];
assign g[18330] = a[13] & g[10138];
assign g[26521] = b[13] & g[10138];
assign g[18331] = a[13] & g[10139];
assign g[26522] = b[13] & g[10139];
assign g[18332] = a[13] & g[10140];
assign g[26523] = b[13] & g[10140];
assign g[18333] = a[13] & g[10141];
assign g[26524] = b[13] & g[10141];
assign g[18334] = a[13] & g[10142];
assign g[26525] = b[13] & g[10142];
assign g[18335] = a[13] & g[10143];
assign g[26526] = b[13] & g[10143];
assign g[18336] = a[13] & g[10144];
assign g[26527] = b[13] & g[10144];
assign g[18337] = a[13] & g[10145];
assign g[26528] = b[13] & g[10145];
assign g[18338] = a[13] & g[10146];
assign g[26529] = b[13] & g[10146];
assign g[18339] = a[13] & g[10147];
assign g[26530] = b[13] & g[10147];
assign g[18340] = a[13] & g[10148];
assign g[26531] = b[13] & g[10148];
assign g[18341] = a[13] & g[10149];
assign g[26532] = b[13] & g[10149];
assign g[18342] = a[13] & g[10150];
assign g[26533] = b[13] & g[10150];
assign g[18343] = a[13] & g[10151];
assign g[26534] = b[13] & g[10151];
assign g[18344] = a[13] & g[10152];
assign g[26535] = b[13] & g[10152];
assign g[18345] = a[13] & g[10153];
assign g[26536] = b[13] & g[10153];
assign g[18346] = a[13] & g[10154];
assign g[26537] = b[13] & g[10154];
assign g[18347] = a[13] & g[10155];
assign g[26538] = b[13] & g[10155];
assign g[18348] = a[13] & g[10156];
assign g[26539] = b[13] & g[10156];
assign g[18349] = a[13] & g[10157];
assign g[26540] = b[13] & g[10157];
assign g[18350] = a[13] & g[10158];
assign g[26541] = b[13] & g[10158];
assign g[18351] = a[13] & g[10159];
assign g[26542] = b[13] & g[10159];
assign g[18352] = a[13] & g[10160];
assign g[26543] = b[13] & g[10160];
assign g[18353] = a[13] & g[10161];
assign g[26544] = b[13] & g[10161];
assign g[18354] = a[13] & g[10162];
assign g[26545] = b[13] & g[10162];
assign g[18355] = a[13] & g[10163];
assign g[26546] = b[13] & g[10163];
assign g[18356] = a[13] & g[10164];
assign g[26547] = b[13] & g[10164];
assign g[18357] = a[13] & g[10165];
assign g[26548] = b[13] & g[10165];
assign g[18358] = a[13] & g[10166];
assign g[26549] = b[13] & g[10166];
assign g[18359] = a[13] & g[10167];
assign g[26550] = b[13] & g[10167];
assign g[18360] = a[13] & g[10168];
assign g[26551] = b[13] & g[10168];
assign g[18361] = a[13] & g[10169];
assign g[26552] = b[13] & g[10169];
assign g[18362] = a[13] & g[10170];
assign g[26553] = b[13] & g[10170];
assign g[18363] = a[13] & g[10171];
assign g[26554] = b[13] & g[10171];
assign g[18364] = a[13] & g[10172];
assign g[26555] = b[13] & g[10172];
assign g[18365] = a[13] & g[10173];
assign g[26556] = b[13] & g[10173];
assign g[18366] = a[13] & g[10174];
assign g[26557] = b[13] & g[10174];
assign g[18367] = a[13] & g[10175];
assign g[26558] = b[13] & g[10175];
assign g[18368] = a[13] & g[10176];
assign g[26559] = b[13] & g[10176];
assign g[18369] = a[13] & g[10177];
assign g[26560] = b[13] & g[10177];
assign g[18370] = a[13] & g[10178];
assign g[26561] = b[13] & g[10178];
assign g[18371] = a[13] & g[10179];
assign g[26562] = b[13] & g[10179];
assign g[18372] = a[13] & g[10180];
assign g[26563] = b[13] & g[10180];
assign g[18373] = a[13] & g[10181];
assign g[26564] = b[13] & g[10181];
assign g[18374] = a[13] & g[10182];
assign g[26565] = b[13] & g[10182];
assign g[18375] = a[13] & g[10183];
assign g[26566] = b[13] & g[10183];
assign g[18376] = a[13] & g[10184];
assign g[26567] = b[13] & g[10184];
assign g[18377] = a[13] & g[10185];
assign g[26568] = b[13] & g[10185];
assign g[18378] = a[13] & g[10186];
assign g[26569] = b[13] & g[10186];
assign g[18379] = a[13] & g[10187];
assign g[26570] = b[13] & g[10187];
assign g[18380] = a[13] & g[10188];
assign g[26571] = b[13] & g[10188];
assign g[18381] = a[13] & g[10189];
assign g[26572] = b[13] & g[10189];
assign g[18382] = a[13] & g[10190];
assign g[26573] = b[13] & g[10190];
assign g[18383] = a[13] & g[10191];
assign g[26574] = b[13] & g[10191];
assign g[18384] = a[13] & g[10192];
assign g[26575] = b[13] & g[10192];
assign g[18385] = a[13] & g[10193];
assign g[26576] = b[13] & g[10193];
assign g[18386] = a[13] & g[10194];
assign g[26577] = b[13] & g[10194];
assign g[18387] = a[13] & g[10195];
assign g[26578] = b[13] & g[10195];
assign g[18388] = a[13] & g[10196];
assign g[26579] = b[13] & g[10196];
assign g[18389] = a[13] & g[10197];
assign g[26580] = b[13] & g[10197];
assign g[18390] = a[13] & g[10198];
assign g[26581] = b[13] & g[10198];
assign g[18391] = a[13] & g[10199];
assign g[26582] = b[13] & g[10199];
assign g[18392] = a[13] & g[10200];
assign g[26583] = b[13] & g[10200];
assign g[18393] = a[13] & g[10201];
assign g[26584] = b[13] & g[10201];
assign g[18394] = a[13] & g[10202];
assign g[26585] = b[13] & g[10202];
assign g[18395] = a[13] & g[10203];
assign g[26586] = b[13] & g[10203];
assign g[18396] = a[13] & g[10204];
assign g[26587] = b[13] & g[10204];
assign g[18397] = a[13] & g[10205];
assign g[26588] = b[13] & g[10205];
assign g[18398] = a[13] & g[10206];
assign g[26589] = b[13] & g[10206];
assign g[18399] = a[13] & g[10207];
assign g[26590] = b[13] & g[10207];
assign g[18400] = a[13] & g[10208];
assign g[26591] = b[13] & g[10208];
assign g[18401] = a[13] & g[10209];
assign g[26592] = b[13] & g[10209];
assign g[18402] = a[13] & g[10210];
assign g[26593] = b[13] & g[10210];
assign g[18403] = a[13] & g[10211];
assign g[26594] = b[13] & g[10211];
assign g[18404] = a[13] & g[10212];
assign g[26595] = b[13] & g[10212];
assign g[18405] = a[13] & g[10213];
assign g[26596] = b[13] & g[10213];
assign g[18406] = a[13] & g[10214];
assign g[26597] = b[13] & g[10214];
assign g[18407] = a[13] & g[10215];
assign g[26598] = b[13] & g[10215];
assign g[18408] = a[13] & g[10216];
assign g[26599] = b[13] & g[10216];
assign g[18409] = a[13] & g[10217];
assign g[26600] = b[13] & g[10217];
assign g[18410] = a[13] & g[10218];
assign g[26601] = b[13] & g[10218];
assign g[18411] = a[13] & g[10219];
assign g[26602] = b[13] & g[10219];
assign g[18412] = a[13] & g[10220];
assign g[26603] = b[13] & g[10220];
assign g[18413] = a[13] & g[10221];
assign g[26604] = b[13] & g[10221];
assign g[18414] = a[13] & g[10222];
assign g[26605] = b[13] & g[10222];
assign g[18415] = a[13] & g[10223];
assign g[26606] = b[13] & g[10223];
assign g[18416] = a[13] & g[10224];
assign g[26607] = b[13] & g[10224];
assign g[18417] = a[13] & g[10225];
assign g[26608] = b[13] & g[10225];
assign g[18418] = a[13] & g[10226];
assign g[26609] = b[13] & g[10226];
assign g[18419] = a[13] & g[10227];
assign g[26610] = b[13] & g[10227];
assign g[18420] = a[13] & g[10228];
assign g[26611] = b[13] & g[10228];
assign g[18421] = a[13] & g[10229];
assign g[26612] = b[13] & g[10229];
assign g[18422] = a[13] & g[10230];
assign g[26613] = b[13] & g[10230];
assign g[18423] = a[13] & g[10231];
assign g[26614] = b[13] & g[10231];
assign g[18424] = a[13] & g[10232];
assign g[26615] = b[13] & g[10232];
assign g[18425] = a[13] & g[10233];
assign g[26616] = b[13] & g[10233];
assign g[18426] = a[13] & g[10234];
assign g[26617] = b[13] & g[10234];
assign g[18427] = a[13] & g[10235];
assign g[26618] = b[13] & g[10235];
assign g[18428] = a[13] & g[10236];
assign g[26619] = b[13] & g[10236];
assign g[18429] = a[13] & g[10237];
assign g[26620] = b[13] & g[10237];
assign g[18430] = a[13] & g[10238];
assign g[26621] = b[13] & g[10238];
assign g[18431] = a[13] & g[10239];
assign g[26622] = b[13] & g[10239];
assign g[18432] = a[13] & g[10240];
assign g[26623] = b[13] & g[10240];
assign g[18433] = a[13] & g[10241];
assign g[26624] = b[13] & g[10241];
assign g[18434] = a[13] & g[10242];
assign g[26625] = b[13] & g[10242];
assign g[18435] = a[13] & g[10243];
assign g[26626] = b[13] & g[10243];
assign g[18436] = a[13] & g[10244];
assign g[26627] = b[13] & g[10244];
assign g[18437] = a[13] & g[10245];
assign g[26628] = b[13] & g[10245];
assign g[18438] = a[13] & g[10246];
assign g[26629] = b[13] & g[10246];
assign g[18439] = a[13] & g[10247];
assign g[26630] = b[13] & g[10247];
assign g[18440] = a[13] & g[10248];
assign g[26631] = b[13] & g[10248];
assign g[18441] = a[13] & g[10249];
assign g[26632] = b[13] & g[10249];
assign g[18442] = a[13] & g[10250];
assign g[26633] = b[13] & g[10250];
assign g[18443] = a[13] & g[10251];
assign g[26634] = b[13] & g[10251];
assign g[18444] = a[13] & g[10252];
assign g[26635] = b[13] & g[10252];
assign g[18445] = a[13] & g[10253];
assign g[26636] = b[13] & g[10253];
assign g[18446] = a[13] & g[10254];
assign g[26637] = b[13] & g[10254];
assign g[18447] = a[13] & g[10255];
assign g[26638] = b[13] & g[10255];
assign g[18448] = a[13] & g[10256];
assign g[26639] = b[13] & g[10256];
assign g[18449] = a[13] & g[10257];
assign g[26640] = b[13] & g[10257];
assign g[18450] = a[13] & g[10258];
assign g[26641] = b[13] & g[10258];
assign g[18451] = a[13] & g[10259];
assign g[26642] = b[13] & g[10259];
assign g[18452] = a[13] & g[10260];
assign g[26643] = b[13] & g[10260];
assign g[18453] = a[13] & g[10261];
assign g[26644] = b[13] & g[10261];
assign g[18454] = a[13] & g[10262];
assign g[26645] = b[13] & g[10262];
assign g[18455] = a[13] & g[10263];
assign g[26646] = b[13] & g[10263];
assign g[18456] = a[13] & g[10264];
assign g[26647] = b[13] & g[10264];
assign g[18457] = a[13] & g[10265];
assign g[26648] = b[13] & g[10265];
assign g[18458] = a[13] & g[10266];
assign g[26649] = b[13] & g[10266];
assign g[18459] = a[13] & g[10267];
assign g[26650] = b[13] & g[10267];
assign g[18460] = a[13] & g[10268];
assign g[26651] = b[13] & g[10268];
assign g[18461] = a[13] & g[10269];
assign g[26652] = b[13] & g[10269];
assign g[18462] = a[13] & g[10270];
assign g[26653] = b[13] & g[10270];
assign g[18463] = a[13] & g[10271];
assign g[26654] = b[13] & g[10271];
assign g[18464] = a[13] & g[10272];
assign g[26655] = b[13] & g[10272];
assign g[18465] = a[13] & g[10273];
assign g[26656] = b[13] & g[10273];
assign g[18466] = a[13] & g[10274];
assign g[26657] = b[13] & g[10274];
assign g[18467] = a[13] & g[10275];
assign g[26658] = b[13] & g[10275];
assign g[18468] = a[13] & g[10276];
assign g[26659] = b[13] & g[10276];
assign g[18469] = a[13] & g[10277];
assign g[26660] = b[13] & g[10277];
assign g[18470] = a[13] & g[10278];
assign g[26661] = b[13] & g[10278];
assign g[18471] = a[13] & g[10279];
assign g[26662] = b[13] & g[10279];
assign g[18472] = a[13] & g[10280];
assign g[26663] = b[13] & g[10280];
assign g[18473] = a[13] & g[10281];
assign g[26664] = b[13] & g[10281];
assign g[18474] = a[13] & g[10282];
assign g[26665] = b[13] & g[10282];
assign g[18475] = a[13] & g[10283];
assign g[26666] = b[13] & g[10283];
assign g[18476] = a[13] & g[10284];
assign g[26667] = b[13] & g[10284];
assign g[18477] = a[13] & g[10285];
assign g[26668] = b[13] & g[10285];
assign g[18478] = a[13] & g[10286];
assign g[26669] = b[13] & g[10286];
assign g[18479] = a[13] & g[10287];
assign g[26670] = b[13] & g[10287];
assign g[18480] = a[13] & g[10288];
assign g[26671] = b[13] & g[10288];
assign g[18481] = a[13] & g[10289];
assign g[26672] = b[13] & g[10289];
assign g[18482] = a[13] & g[10290];
assign g[26673] = b[13] & g[10290];
assign g[18483] = a[13] & g[10291];
assign g[26674] = b[13] & g[10291];
assign g[18484] = a[13] & g[10292];
assign g[26675] = b[13] & g[10292];
assign g[18485] = a[13] & g[10293];
assign g[26676] = b[13] & g[10293];
assign g[18486] = a[13] & g[10294];
assign g[26677] = b[13] & g[10294];
assign g[18487] = a[13] & g[10295];
assign g[26678] = b[13] & g[10295];
assign g[18488] = a[13] & g[10296];
assign g[26679] = b[13] & g[10296];
assign g[18489] = a[13] & g[10297];
assign g[26680] = b[13] & g[10297];
assign g[18490] = a[13] & g[10298];
assign g[26681] = b[13] & g[10298];
assign g[18491] = a[13] & g[10299];
assign g[26682] = b[13] & g[10299];
assign g[18492] = a[13] & g[10300];
assign g[26683] = b[13] & g[10300];
assign g[18493] = a[13] & g[10301];
assign g[26684] = b[13] & g[10301];
assign g[18494] = a[13] & g[10302];
assign g[26685] = b[13] & g[10302];
assign g[18495] = a[13] & g[10303];
assign g[26686] = b[13] & g[10303];
assign g[18496] = a[13] & g[10304];
assign g[26687] = b[13] & g[10304];
assign g[18497] = a[13] & g[10305];
assign g[26688] = b[13] & g[10305];
assign g[18498] = a[13] & g[10306];
assign g[26689] = b[13] & g[10306];
assign g[18499] = a[13] & g[10307];
assign g[26690] = b[13] & g[10307];
assign g[18500] = a[13] & g[10308];
assign g[26691] = b[13] & g[10308];
assign g[18501] = a[13] & g[10309];
assign g[26692] = b[13] & g[10309];
assign g[18502] = a[13] & g[10310];
assign g[26693] = b[13] & g[10310];
assign g[18503] = a[13] & g[10311];
assign g[26694] = b[13] & g[10311];
assign g[18504] = a[13] & g[10312];
assign g[26695] = b[13] & g[10312];
assign g[18505] = a[13] & g[10313];
assign g[26696] = b[13] & g[10313];
assign g[18506] = a[13] & g[10314];
assign g[26697] = b[13] & g[10314];
assign g[18507] = a[13] & g[10315];
assign g[26698] = b[13] & g[10315];
assign g[18508] = a[13] & g[10316];
assign g[26699] = b[13] & g[10316];
assign g[18509] = a[13] & g[10317];
assign g[26700] = b[13] & g[10317];
assign g[18510] = a[13] & g[10318];
assign g[26701] = b[13] & g[10318];
assign g[18511] = a[13] & g[10319];
assign g[26702] = b[13] & g[10319];
assign g[18512] = a[13] & g[10320];
assign g[26703] = b[13] & g[10320];
assign g[18513] = a[13] & g[10321];
assign g[26704] = b[13] & g[10321];
assign g[18514] = a[13] & g[10322];
assign g[26705] = b[13] & g[10322];
assign g[18515] = a[13] & g[10323];
assign g[26706] = b[13] & g[10323];
assign g[18516] = a[13] & g[10324];
assign g[26707] = b[13] & g[10324];
assign g[18517] = a[13] & g[10325];
assign g[26708] = b[13] & g[10325];
assign g[18518] = a[13] & g[10326];
assign g[26709] = b[13] & g[10326];
assign g[18519] = a[13] & g[10327];
assign g[26710] = b[13] & g[10327];
assign g[18520] = a[13] & g[10328];
assign g[26711] = b[13] & g[10328];
assign g[18521] = a[13] & g[10329];
assign g[26712] = b[13] & g[10329];
assign g[18522] = a[13] & g[10330];
assign g[26713] = b[13] & g[10330];
assign g[18523] = a[13] & g[10331];
assign g[26714] = b[13] & g[10331];
assign g[18524] = a[13] & g[10332];
assign g[26715] = b[13] & g[10332];
assign g[18525] = a[13] & g[10333];
assign g[26716] = b[13] & g[10333];
assign g[18526] = a[13] & g[10334];
assign g[26717] = b[13] & g[10334];
assign g[18527] = a[13] & g[10335];
assign g[26718] = b[13] & g[10335];
assign g[18528] = a[13] & g[10336];
assign g[26719] = b[13] & g[10336];
assign g[18529] = a[13] & g[10337];
assign g[26720] = b[13] & g[10337];
assign g[18530] = a[13] & g[10338];
assign g[26721] = b[13] & g[10338];
assign g[18531] = a[13] & g[10339];
assign g[26722] = b[13] & g[10339];
assign g[18532] = a[13] & g[10340];
assign g[26723] = b[13] & g[10340];
assign g[18533] = a[13] & g[10341];
assign g[26724] = b[13] & g[10341];
assign g[18534] = a[13] & g[10342];
assign g[26725] = b[13] & g[10342];
assign g[18535] = a[13] & g[10343];
assign g[26726] = b[13] & g[10343];
assign g[18536] = a[13] & g[10344];
assign g[26727] = b[13] & g[10344];
assign g[18537] = a[13] & g[10345];
assign g[26728] = b[13] & g[10345];
assign g[18538] = a[13] & g[10346];
assign g[26729] = b[13] & g[10346];
assign g[18539] = a[13] & g[10347];
assign g[26730] = b[13] & g[10347];
assign g[18540] = a[13] & g[10348];
assign g[26731] = b[13] & g[10348];
assign g[18541] = a[13] & g[10349];
assign g[26732] = b[13] & g[10349];
assign g[18542] = a[13] & g[10350];
assign g[26733] = b[13] & g[10350];
assign g[18543] = a[13] & g[10351];
assign g[26734] = b[13] & g[10351];
assign g[18544] = a[13] & g[10352];
assign g[26735] = b[13] & g[10352];
assign g[18545] = a[13] & g[10353];
assign g[26736] = b[13] & g[10353];
assign g[18546] = a[13] & g[10354];
assign g[26737] = b[13] & g[10354];
assign g[18547] = a[13] & g[10355];
assign g[26738] = b[13] & g[10355];
assign g[18548] = a[13] & g[10356];
assign g[26739] = b[13] & g[10356];
assign g[18549] = a[13] & g[10357];
assign g[26740] = b[13] & g[10357];
assign g[18550] = a[13] & g[10358];
assign g[26741] = b[13] & g[10358];
assign g[18551] = a[13] & g[10359];
assign g[26742] = b[13] & g[10359];
assign g[18552] = a[13] & g[10360];
assign g[26743] = b[13] & g[10360];
assign g[18553] = a[13] & g[10361];
assign g[26744] = b[13] & g[10361];
assign g[18554] = a[13] & g[10362];
assign g[26745] = b[13] & g[10362];
assign g[18555] = a[13] & g[10363];
assign g[26746] = b[13] & g[10363];
assign g[18556] = a[13] & g[10364];
assign g[26747] = b[13] & g[10364];
assign g[18557] = a[13] & g[10365];
assign g[26748] = b[13] & g[10365];
assign g[18558] = a[13] & g[10366];
assign g[26749] = b[13] & g[10366];
assign g[18559] = a[13] & g[10367];
assign g[26750] = b[13] & g[10367];
assign g[18560] = a[13] & g[10368];
assign g[26751] = b[13] & g[10368];
assign g[18561] = a[13] & g[10369];
assign g[26752] = b[13] & g[10369];
assign g[18562] = a[13] & g[10370];
assign g[26753] = b[13] & g[10370];
assign g[18563] = a[13] & g[10371];
assign g[26754] = b[13] & g[10371];
assign g[18564] = a[13] & g[10372];
assign g[26755] = b[13] & g[10372];
assign g[18565] = a[13] & g[10373];
assign g[26756] = b[13] & g[10373];
assign g[18566] = a[13] & g[10374];
assign g[26757] = b[13] & g[10374];
assign g[18567] = a[13] & g[10375];
assign g[26758] = b[13] & g[10375];
assign g[18568] = a[13] & g[10376];
assign g[26759] = b[13] & g[10376];
assign g[18569] = a[13] & g[10377];
assign g[26760] = b[13] & g[10377];
assign g[18570] = a[13] & g[10378];
assign g[26761] = b[13] & g[10378];
assign g[18571] = a[13] & g[10379];
assign g[26762] = b[13] & g[10379];
assign g[18572] = a[13] & g[10380];
assign g[26763] = b[13] & g[10380];
assign g[18573] = a[13] & g[10381];
assign g[26764] = b[13] & g[10381];
assign g[18574] = a[13] & g[10382];
assign g[26765] = b[13] & g[10382];
assign g[18575] = a[13] & g[10383];
assign g[26766] = b[13] & g[10383];
assign g[18576] = a[13] & g[10384];
assign g[26767] = b[13] & g[10384];
assign g[18577] = a[13] & g[10385];
assign g[26768] = b[13] & g[10385];
assign g[18578] = a[13] & g[10386];
assign g[26769] = b[13] & g[10386];
assign g[18579] = a[13] & g[10387];
assign g[26770] = b[13] & g[10387];
assign g[18580] = a[13] & g[10388];
assign g[26771] = b[13] & g[10388];
assign g[18581] = a[13] & g[10389];
assign g[26772] = b[13] & g[10389];
assign g[18582] = a[13] & g[10390];
assign g[26773] = b[13] & g[10390];
assign g[18583] = a[13] & g[10391];
assign g[26774] = b[13] & g[10391];
assign g[18584] = a[13] & g[10392];
assign g[26775] = b[13] & g[10392];
assign g[18585] = a[13] & g[10393];
assign g[26776] = b[13] & g[10393];
assign g[18586] = a[13] & g[10394];
assign g[26777] = b[13] & g[10394];
assign g[18587] = a[13] & g[10395];
assign g[26778] = b[13] & g[10395];
assign g[18588] = a[13] & g[10396];
assign g[26779] = b[13] & g[10396];
assign g[18589] = a[13] & g[10397];
assign g[26780] = b[13] & g[10397];
assign g[18590] = a[13] & g[10398];
assign g[26781] = b[13] & g[10398];
assign g[18591] = a[13] & g[10399];
assign g[26782] = b[13] & g[10399];
assign g[18592] = a[13] & g[10400];
assign g[26783] = b[13] & g[10400];
assign g[18593] = a[13] & g[10401];
assign g[26784] = b[13] & g[10401];
assign g[18594] = a[13] & g[10402];
assign g[26785] = b[13] & g[10402];
assign g[18595] = a[13] & g[10403];
assign g[26786] = b[13] & g[10403];
assign g[18596] = a[13] & g[10404];
assign g[26787] = b[13] & g[10404];
assign g[18597] = a[13] & g[10405];
assign g[26788] = b[13] & g[10405];
assign g[18598] = a[13] & g[10406];
assign g[26789] = b[13] & g[10406];
assign g[18599] = a[13] & g[10407];
assign g[26790] = b[13] & g[10407];
assign g[18600] = a[13] & g[10408];
assign g[26791] = b[13] & g[10408];
assign g[18601] = a[13] & g[10409];
assign g[26792] = b[13] & g[10409];
assign g[18602] = a[13] & g[10410];
assign g[26793] = b[13] & g[10410];
assign g[18603] = a[13] & g[10411];
assign g[26794] = b[13] & g[10411];
assign g[18604] = a[13] & g[10412];
assign g[26795] = b[13] & g[10412];
assign g[18605] = a[13] & g[10413];
assign g[26796] = b[13] & g[10413];
assign g[18606] = a[13] & g[10414];
assign g[26797] = b[13] & g[10414];
assign g[18607] = a[13] & g[10415];
assign g[26798] = b[13] & g[10415];
assign g[18608] = a[13] & g[10416];
assign g[26799] = b[13] & g[10416];
assign g[18609] = a[13] & g[10417];
assign g[26800] = b[13] & g[10417];
assign g[18610] = a[13] & g[10418];
assign g[26801] = b[13] & g[10418];
assign g[18611] = a[13] & g[10419];
assign g[26802] = b[13] & g[10419];
assign g[18612] = a[13] & g[10420];
assign g[26803] = b[13] & g[10420];
assign g[18613] = a[13] & g[10421];
assign g[26804] = b[13] & g[10421];
assign g[18614] = a[13] & g[10422];
assign g[26805] = b[13] & g[10422];
assign g[18615] = a[13] & g[10423];
assign g[26806] = b[13] & g[10423];
assign g[18616] = a[13] & g[10424];
assign g[26807] = b[13] & g[10424];
assign g[18617] = a[13] & g[10425];
assign g[26808] = b[13] & g[10425];
assign g[18618] = a[13] & g[10426];
assign g[26809] = b[13] & g[10426];
assign g[18619] = a[13] & g[10427];
assign g[26810] = b[13] & g[10427];
assign g[18620] = a[13] & g[10428];
assign g[26811] = b[13] & g[10428];
assign g[18621] = a[13] & g[10429];
assign g[26812] = b[13] & g[10429];
assign g[18622] = a[13] & g[10430];
assign g[26813] = b[13] & g[10430];
assign g[18623] = a[13] & g[10431];
assign g[26814] = b[13] & g[10431];
assign g[18624] = a[13] & g[10432];
assign g[26815] = b[13] & g[10432];
assign g[18625] = a[13] & g[10433];
assign g[26816] = b[13] & g[10433];
assign g[18626] = a[13] & g[10434];
assign g[26817] = b[13] & g[10434];
assign g[18627] = a[13] & g[10435];
assign g[26818] = b[13] & g[10435];
assign g[18628] = a[13] & g[10436];
assign g[26819] = b[13] & g[10436];
assign g[18629] = a[13] & g[10437];
assign g[26820] = b[13] & g[10437];
assign g[18630] = a[13] & g[10438];
assign g[26821] = b[13] & g[10438];
assign g[18631] = a[13] & g[10439];
assign g[26822] = b[13] & g[10439];
assign g[18632] = a[13] & g[10440];
assign g[26823] = b[13] & g[10440];
assign g[18633] = a[13] & g[10441];
assign g[26824] = b[13] & g[10441];
assign g[18634] = a[13] & g[10442];
assign g[26825] = b[13] & g[10442];
assign g[18635] = a[13] & g[10443];
assign g[26826] = b[13] & g[10443];
assign g[18636] = a[13] & g[10444];
assign g[26827] = b[13] & g[10444];
assign g[18637] = a[13] & g[10445];
assign g[26828] = b[13] & g[10445];
assign g[18638] = a[13] & g[10446];
assign g[26829] = b[13] & g[10446];
assign g[18639] = a[13] & g[10447];
assign g[26830] = b[13] & g[10447];
assign g[18640] = a[13] & g[10448];
assign g[26831] = b[13] & g[10448];
assign g[18641] = a[13] & g[10449];
assign g[26832] = b[13] & g[10449];
assign g[18642] = a[13] & g[10450];
assign g[26833] = b[13] & g[10450];
assign g[18643] = a[13] & g[10451];
assign g[26834] = b[13] & g[10451];
assign g[18644] = a[13] & g[10452];
assign g[26835] = b[13] & g[10452];
assign g[18645] = a[13] & g[10453];
assign g[26836] = b[13] & g[10453];
assign g[18646] = a[13] & g[10454];
assign g[26837] = b[13] & g[10454];
assign g[18647] = a[13] & g[10455];
assign g[26838] = b[13] & g[10455];
assign g[18648] = a[13] & g[10456];
assign g[26839] = b[13] & g[10456];
assign g[18649] = a[13] & g[10457];
assign g[26840] = b[13] & g[10457];
assign g[18650] = a[13] & g[10458];
assign g[26841] = b[13] & g[10458];
assign g[18651] = a[13] & g[10459];
assign g[26842] = b[13] & g[10459];
assign g[18652] = a[13] & g[10460];
assign g[26843] = b[13] & g[10460];
assign g[18653] = a[13] & g[10461];
assign g[26844] = b[13] & g[10461];
assign g[18654] = a[13] & g[10462];
assign g[26845] = b[13] & g[10462];
assign g[18655] = a[13] & g[10463];
assign g[26846] = b[13] & g[10463];
assign g[18656] = a[13] & g[10464];
assign g[26847] = b[13] & g[10464];
assign g[18657] = a[13] & g[10465];
assign g[26848] = b[13] & g[10465];
assign g[18658] = a[13] & g[10466];
assign g[26849] = b[13] & g[10466];
assign g[18659] = a[13] & g[10467];
assign g[26850] = b[13] & g[10467];
assign g[18660] = a[13] & g[10468];
assign g[26851] = b[13] & g[10468];
assign g[18661] = a[13] & g[10469];
assign g[26852] = b[13] & g[10469];
assign g[18662] = a[13] & g[10470];
assign g[26853] = b[13] & g[10470];
assign g[18663] = a[13] & g[10471];
assign g[26854] = b[13] & g[10471];
assign g[18664] = a[13] & g[10472];
assign g[26855] = b[13] & g[10472];
assign g[18665] = a[13] & g[10473];
assign g[26856] = b[13] & g[10473];
assign g[18666] = a[13] & g[10474];
assign g[26857] = b[13] & g[10474];
assign g[18667] = a[13] & g[10475];
assign g[26858] = b[13] & g[10475];
assign g[18668] = a[13] & g[10476];
assign g[26859] = b[13] & g[10476];
assign g[18669] = a[13] & g[10477];
assign g[26860] = b[13] & g[10477];
assign g[18670] = a[13] & g[10478];
assign g[26861] = b[13] & g[10478];
assign g[18671] = a[13] & g[10479];
assign g[26862] = b[13] & g[10479];
assign g[18672] = a[13] & g[10480];
assign g[26863] = b[13] & g[10480];
assign g[18673] = a[13] & g[10481];
assign g[26864] = b[13] & g[10481];
assign g[18674] = a[13] & g[10482];
assign g[26865] = b[13] & g[10482];
assign g[18675] = a[13] & g[10483];
assign g[26866] = b[13] & g[10483];
assign g[18676] = a[13] & g[10484];
assign g[26867] = b[13] & g[10484];
assign g[18677] = a[13] & g[10485];
assign g[26868] = b[13] & g[10485];
assign g[18678] = a[13] & g[10486];
assign g[26869] = b[13] & g[10486];
assign g[18679] = a[13] & g[10487];
assign g[26870] = b[13] & g[10487];
assign g[18680] = a[13] & g[10488];
assign g[26871] = b[13] & g[10488];
assign g[18681] = a[13] & g[10489];
assign g[26872] = b[13] & g[10489];
assign g[18682] = a[13] & g[10490];
assign g[26873] = b[13] & g[10490];
assign g[18683] = a[13] & g[10491];
assign g[26874] = b[13] & g[10491];
assign g[18684] = a[13] & g[10492];
assign g[26875] = b[13] & g[10492];
assign g[18685] = a[13] & g[10493];
assign g[26876] = b[13] & g[10493];
assign g[18686] = a[13] & g[10494];
assign g[26877] = b[13] & g[10494];
assign g[18687] = a[13] & g[10495];
assign g[26878] = b[13] & g[10495];
assign g[18688] = a[13] & g[10496];
assign g[26879] = b[13] & g[10496];
assign g[18689] = a[13] & g[10497];
assign g[26880] = b[13] & g[10497];
assign g[18690] = a[13] & g[10498];
assign g[26881] = b[13] & g[10498];
assign g[18691] = a[13] & g[10499];
assign g[26882] = b[13] & g[10499];
assign g[18692] = a[13] & g[10500];
assign g[26883] = b[13] & g[10500];
assign g[18693] = a[13] & g[10501];
assign g[26884] = b[13] & g[10501];
assign g[18694] = a[13] & g[10502];
assign g[26885] = b[13] & g[10502];
assign g[18695] = a[13] & g[10503];
assign g[26886] = b[13] & g[10503];
assign g[18696] = a[13] & g[10504];
assign g[26887] = b[13] & g[10504];
assign g[18697] = a[13] & g[10505];
assign g[26888] = b[13] & g[10505];
assign g[18698] = a[13] & g[10506];
assign g[26889] = b[13] & g[10506];
assign g[18699] = a[13] & g[10507];
assign g[26890] = b[13] & g[10507];
assign g[18700] = a[13] & g[10508];
assign g[26891] = b[13] & g[10508];
assign g[18701] = a[13] & g[10509];
assign g[26892] = b[13] & g[10509];
assign g[18702] = a[13] & g[10510];
assign g[26893] = b[13] & g[10510];
assign g[18703] = a[13] & g[10511];
assign g[26894] = b[13] & g[10511];
assign g[18704] = a[13] & g[10512];
assign g[26895] = b[13] & g[10512];
assign g[18705] = a[13] & g[10513];
assign g[26896] = b[13] & g[10513];
assign g[18706] = a[13] & g[10514];
assign g[26897] = b[13] & g[10514];
assign g[18707] = a[13] & g[10515];
assign g[26898] = b[13] & g[10515];
assign g[18708] = a[13] & g[10516];
assign g[26899] = b[13] & g[10516];
assign g[18709] = a[13] & g[10517];
assign g[26900] = b[13] & g[10517];
assign g[18710] = a[13] & g[10518];
assign g[26901] = b[13] & g[10518];
assign g[18711] = a[13] & g[10519];
assign g[26902] = b[13] & g[10519];
assign g[18712] = a[13] & g[10520];
assign g[26903] = b[13] & g[10520];
assign g[18713] = a[13] & g[10521];
assign g[26904] = b[13] & g[10521];
assign g[18714] = a[13] & g[10522];
assign g[26905] = b[13] & g[10522];
assign g[18715] = a[13] & g[10523];
assign g[26906] = b[13] & g[10523];
assign g[18716] = a[13] & g[10524];
assign g[26907] = b[13] & g[10524];
assign g[18717] = a[13] & g[10525];
assign g[26908] = b[13] & g[10525];
assign g[18718] = a[13] & g[10526];
assign g[26909] = b[13] & g[10526];
assign g[18719] = a[13] & g[10527];
assign g[26910] = b[13] & g[10527];
assign g[18720] = a[13] & g[10528];
assign g[26911] = b[13] & g[10528];
assign g[18721] = a[13] & g[10529];
assign g[26912] = b[13] & g[10529];
assign g[18722] = a[13] & g[10530];
assign g[26913] = b[13] & g[10530];
assign g[18723] = a[13] & g[10531];
assign g[26914] = b[13] & g[10531];
assign g[18724] = a[13] & g[10532];
assign g[26915] = b[13] & g[10532];
assign g[18725] = a[13] & g[10533];
assign g[26916] = b[13] & g[10533];
assign g[18726] = a[13] & g[10534];
assign g[26917] = b[13] & g[10534];
assign g[18727] = a[13] & g[10535];
assign g[26918] = b[13] & g[10535];
assign g[18728] = a[13] & g[10536];
assign g[26919] = b[13] & g[10536];
assign g[18729] = a[13] & g[10537];
assign g[26920] = b[13] & g[10537];
assign g[18730] = a[13] & g[10538];
assign g[26921] = b[13] & g[10538];
assign g[18731] = a[13] & g[10539];
assign g[26922] = b[13] & g[10539];
assign g[18732] = a[13] & g[10540];
assign g[26923] = b[13] & g[10540];
assign g[18733] = a[13] & g[10541];
assign g[26924] = b[13] & g[10541];
assign g[18734] = a[13] & g[10542];
assign g[26925] = b[13] & g[10542];
assign g[18735] = a[13] & g[10543];
assign g[26926] = b[13] & g[10543];
assign g[18736] = a[13] & g[10544];
assign g[26927] = b[13] & g[10544];
assign g[18737] = a[13] & g[10545];
assign g[26928] = b[13] & g[10545];
assign g[18738] = a[13] & g[10546];
assign g[26929] = b[13] & g[10546];
assign g[18739] = a[13] & g[10547];
assign g[26930] = b[13] & g[10547];
assign g[18740] = a[13] & g[10548];
assign g[26931] = b[13] & g[10548];
assign g[18741] = a[13] & g[10549];
assign g[26932] = b[13] & g[10549];
assign g[18742] = a[13] & g[10550];
assign g[26933] = b[13] & g[10550];
assign g[18743] = a[13] & g[10551];
assign g[26934] = b[13] & g[10551];
assign g[18744] = a[13] & g[10552];
assign g[26935] = b[13] & g[10552];
assign g[18745] = a[13] & g[10553];
assign g[26936] = b[13] & g[10553];
assign g[18746] = a[13] & g[10554];
assign g[26937] = b[13] & g[10554];
assign g[18747] = a[13] & g[10555];
assign g[26938] = b[13] & g[10555];
assign g[18748] = a[13] & g[10556];
assign g[26939] = b[13] & g[10556];
assign g[18749] = a[13] & g[10557];
assign g[26940] = b[13] & g[10557];
assign g[18750] = a[13] & g[10558];
assign g[26941] = b[13] & g[10558];
assign g[18751] = a[13] & g[10559];
assign g[26942] = b[13] & g[10559];
assign g[18752] = a[13] & g[10560];
assign g[26943] = b[13] & g[10560];
assign g[18753] = a[13] & g[10561];
assign g[26944] = b[13] & g[10561];
assign g[18754] = a[13] & g[10562];
assign g[26945] = b[13] & g[10562];
assign g[18755] = a[13] & g[10563];
assign g[26946] = b[13] & g[10563];
assign g[18756] = a[13] & g[10564];
assign g[26947] = b[13] & g[10564];
assign g[18757] = a[13] & g[10565];
assign g[26948] = b[13] & g[10565];
assign g[18758] = a[13] & g[10566];
assign g[26949] = b[13] & g[10566];
assign g[18759] = a[13] & g[10567];
assign g[26950] = b[13] & g[10567];
assign g[18760] = a[13] & g[10568];
assign g[26951] = b[13] & g[10568];
assign g[18761] = a[13] & g[10569];
assign g[26952] = b[13] & g[10569];
assign g[18762] = a[13] & g[10570];
assign g[26953] = b[13] & g[10570];
assign g[18763] = a[13] & g[10571];
assign g[26954] = b[13] & g[10571];
assign g[18764] = a[13] & g[10572];
assign g[26955] = b[13] & g[10572];
assign g[18765] = a[13] & g[10573];
assign g[26956] = b[13] & g[10573];
assign g[18766] = a[13] & g[10574];
assign g[26957] = b[13] & g[10574];
assign g[18767] = a[13] & g[10575];
assign g[26958] = b[13] & g[10575];
assign g[18768] = a[13] & g[10576];
assign g[26959] = b[13] & g[10576];
assign g[18769] = a[13] & g[10577];
assign g[26960] = b[13] & g[10577];
assign g[18770] = a[13] & g[10578];
assign g[26961] = b[13] & g[10578];
assign g[18771] = a[13] & g[10579];
assign g[26962] = b[13] & g[10579];
assign g[18772] = a[13] & g[10580];
assign g[26963] = b[13] & g[10580];
assign g[18773] = a[13] & g[10581];
assign g[26964] = b[13] & g[10581];
assign g[18774] = a[13] & g[10582];
assign g[26965] = b[13] & g[10582];
assign g[18775] = a[13] & g[10583];
assign g[26966] = b[13] & g[10583];
assign g[18776] = a[13] & g[10584];
assign g[26967] = b[13] & g[10584];
assign g[18777] = a[13] & g[10585];
assign g[26968] = b[13] & g[10585];
assign g[18778] = a[13] & g[10586];
assign g[26969] = b[13] & g[10586];
assign g[18779] = a[13] & g[10587];
assign g[26970] = b[13] & g[10587];
assign g[18780] = a[13] & g[10588];
assign g[26971] = b[13] & g[10588];
assign g[18781] = a[13] & g[10589];
assign g[26972] = b[13] & g[10589];
assign g[18782] = a[13] & g[10590];
assign g[26973] = b[13] & g[10590];
assign g[18783] = a[13] & g[10591];
assign g[26974] = b[13] & g[10591];
assign g[18784] = a[13] & g[10592];
assign g[26975] = b[13] & g[10592];
assign g[18785] = a[13] & g[10593];
assign g[26976] = b[13] & g[10593];
assign g[18786] = a[13] & g[10594];
assign g[26977] = b[13] & g[10594];
assign g[18787] = a[13] & g[10595];
assign g[26978] = b[13] & g[10595];
assign g[18788] = a[13] & g[10596];
assign g[26979] = b[13] & g[10596];
assign g[18789] = a[13] & g[10597];
assign g[26980] = b[13] & g[10597];
assign g[18790] = a[13] & g[10598];
assign g[26981] = b[13] & g[10598];
assign g[18791] = a[13] & g[10599];
assign g[26982] = b[13] & g[10599];
assign g[18792] = a[13] & g[10600];
assign g[26983] = b[13] & g[10600];
assign g[18793] = a[13] & g[10601];
assign g[26984] = b[13] & g[10601];
assign g[18794] = a[13] & g[10602];
assign g[26985] = b[13] & g[10602];
assign g[18795] = a[13] & g[10603];
assign g[26986] = b[13] & g[10603];
assign g[18796] = a[13] & g[10604];
assign g[26987] = b[13] & g[10604];
assign g[18797] = a[13] & g[10605];
assign g[26988] = b[13] & g[10605];
assign g[18798] = a[13] & g[10606];
assign g[26989] = b[13] & g[10606];
assign g[18799] = a[13] & g[10607];
assign g[26990] = b[13] & g[10607];
assign g[18800] = a[13] & g[10608];
assign g[26991] = b[13] & g[10608];
assign g[18801] = a[13] & g[10609];
assign g[26992] = b[13] & g[10609];
assign g[18802] = a[13] & g[10610];
assign g[26993] = b[13] & g[10610];
assign g[18803] = a[13] & g[10611];
assign g[26994] = b[13] & g[10611];
assign g[18804] = a[13] & g[10612];
assign g[26995] = b[13] & g[10612];
assign g[18805] = a[13] & g[10613];
assign g[26996] = b[13] & g[10613];
assign g[18806] = a[13] & g[10614];
assign g[26997] = b[13] & g[10614];
assign g[18807] = a[13] & g[10615];
assign g[26998] = b[13] & g[10615];
assign g[18808] = a[13] & g[10616];
assign g[26999] = b[13] & g[10616];
assign g[18809] = a[13] & g[10617];
assign g[27000] = b[13] & g[10617];
assign g[18810] = a[13] & g[10618];
assign g[27001] = b[13] & g[10618];
assign g[18811] = a[13] & g[10619];
assign g[27002] = b[13] & g[10619];
assign g[18812] = a[13] & g[10620];
assign g[27003] = b[13] & g[10620];
assign g[18813] = a[13] & g[10621];
assign g[27004] = b[13] & g[10621];
assign g[18814] = a[13] & g[10622];
assign g[27005] = b[13] & g[10622];
assign g[18815] = a[13] & g[10623];
assign g[27006] = b[13] & g[10623];
assign g[18816] = a[13] & g[10624];
assign g[27007] = b[13] & g[10624];
assign g[18817] = a[13] & g[10625];
assign g[27008] = b[13] & g[10625];
assign g[18818] = a[13] & g[10626];
assign g[27009] = b[13] & g[10626];
assign g[18819] = a[13] & g[10627];
assign g[27010] = b[13] & g[10627];
assign g[18820] = a[13] & g[10628];
assign g[27011] = b[13] & g[10628];
assign g[18821] = a[13] & g[10629];
assign g[27012] = b[13] & g[10629];
assign g[18822] = a[13] & g[10630];
assign g[27013] = b[13] & g[10630];
assign g[18823] = a[13] & g[10631];
assign g[27014] = b[13] & g[10631];
assign g[18824] = a[13] & g[10632];
assign g[27015] = b[13] & g[10632];
assign g[18825] = a[13] & g[10633];
assign g[27016] = b[13] & g[10633];
assign g[18826] = a[13] & g[10634];
assign g[27017] = b[13] & g[10634];
assign g[18827] = a[13] & g[10635];
assign g[27018] = b[13] & g[10635];
assign g[18828] = a[13] & g[10636];
assign g[27019] = b[13] & g[10636];
assign g[18829] = a[13] & g[10637];
assign g[27020] = b[13] & g[10637];
assign g[18830] = a[13] & g[10638];
assign g[27021] = b[13] & g[10638];
assign g[18831] = a[13] & g[10639];
assign g[27022] = b[13] & g[10639];
assign g[18832] = a[13] & g[10640];
assign g[27023] = b[13] & g[10640];
assign g[18833] = a[13] & g[10641];
assign g[27024] = b[13] & g[10641];
assign g[18834] = a[13] & g[10642];
assign g[27025] = b[13] & g[10642];
assign g[18835] = a[13] & g[10643];
assign g[27026] = b[13] & g[10643];
assign g[18836] = a[13] & g[10644];
assign g[27027] = b[13] & g[10644];
assign g[18837] = a[13] & g[10645];
assign g[27028] = b[13] & g[10645];
assign g[18838] = a[13] & g[10646];
assign g[27029] = b[13] & g[10646];
assign g[18839] = a[13] & g[10647];
assign g[27030] = b[13] & g[10647];
assign g[18840] = a[13] & g[10648];
assign g[27031] = b[13] & g[10648];
assign g[18841] = a[13] & g[10649];
assign g[27032] = b[13] & g[10649];
assign g[18842] = a[13] & g[10650];
assign g[27033] = b[13] & g[10650];
assign g[18843] = a[13] & g[10651];
assign g[27034] = b[13] & g[10651];
assign g[18844] = a[13] & g[10652];
assign g[27035] = b[13] & g[10652];
assign g[18845] = a[13] & g[10653];
assign g[27036] = b[13] & g[10653];
assign g[18846] = a[13] & g[10654];
assign g[27037] = b[13] & g[10654];
assign g[18847] = a[13] & g[10655];
assign g[27038] = b[13] & g[10655];
assign g[18848] = a[13] & g[10656];
assign g[27039] = b[13] & g[10656];
assign g[18849] = a[13] & g[10657];
assign g[27040] = b[13] & g[10657];
assign g[18850] = a[13] & g[10658];
assign g[27041] = b[13] & g[10658];
assign g[18851] = a[13] & g[10659];
assign g[27042] = b[13] & g[10659];
assign g[18852] = a[13] & g[10660];
assign g[27043] = b[13] & g[10660];
assign g[18853] = a[13] & g[10661];
assign g[27044] = b[13] & g[10661];
assign g[18854] = a[13] & g[10662];
assign g[27045] = b[13] & g[10662];
assign g[18855] = a[13] & g[10663];
assign g[27046] = b[13] & g[10663];
assign g[18856] = a[13] & g[10664];
assign g[27047] = b[13] & g[10664];
assign g[18857] = a[13] & g[10665];
assign g[27048] = b[13] & g[10665];
assign g[18858] = a[13] & g[10666];
assign g[27049] = b[13] & g[10666];
assign g[18859] = a[13] & g[10667];
assign g[27050] = b[13] & g[10667];
assign g[18860] = a[13] & g[10668];
assign g[27051] = b[13] & g[10668];
assign g[18861] = a[13] & g[10669];
assign g[27052] = b[13] & g[10669];
assign g[18862] = a[13] & g[10670];
assign g[27053] = b[13] & g[10670];
assign g[18863] = a[13] & g[10671];
assign g[27054] = b[13] & g[10671];
assign g[18864] = a[13] & g[10672];
assign g[27055] = b[13] & g[10672];
assign g[18865] = a[13] & g[10673];
assign g[27056] = b[13] & g[10673];
assign g[18866] = a[13] & g[10674];
assign g[27057] = b[13] & g[10674];
assign g[18867] = a[13] & g[10675];
assign g[27058] = b[13] & g[10675];
assign g[18868] = a[13] & g[10676];
assign g[27059] = b[13] & g[10676];
assign g[18869] = a[13] & g[10677];
assign g[27060] = b[13] & g[10677];
assign g[18870] = a[13] & g[10678];
assign g[27061] = b[13] & g[10678];
assign g[18871] = a[13] & g[10679];
assign g[27062] = b[13] & g[10679];
assign g[18872] = a[13] & g[10680];
assign g[27063] = b[13] & g[10680];
assign g[18873] = a[13] & g[10681];
assign g[27064] = b[13] & g[10681];
assign g[18874] = a[13] & g[10682];
assign g[27065] = b[13] & g[10682];
assign g[18875] = a[13] & g[10683];
assign g[27066] = b[13] & g[10683];
assign g[18876] = a[13] & g[10684];
assign g[27067] = b[13] & g[10684];
assign g[18877] = a[13] & g[10685];
assign g[27068] = b[13] & g[10685];
assign g[18878] = a[13] & g[10686];
assign g[27069] = b[13] & g[10686];
assign g[18879] = a[13] & g[10687];
assign g[27070] = b[13] & g[10687];
assign g[18880] = a[13] & g[10688];
assign g[27071] = b[13] & g[10688];
assign g[18881] = a[13] & g[10689];
assign g[27072] = b[13] & g[10689];
assign g[18882] = a[13] & g[10690];
assign g[27073] = b[13] & g[10690];
assign g[18883] = a[13] & g[10691];
assign g[27074] = b[13] & g[10691];
assign g[18884] = a[13] & g[10692];
assign g[27075] = b[13] & g[10692];
assign g[18885] = a[13] & g[10693];
assign g[27076] = b[13] & g[10693];
assign g[18886] = a[13] & g[10694];
assign g[27077] = b[13] & g[10694];
assign g[18887] = a[13] & g[10695];
assign g[27078] = b[13] & g[10695];
assign g[18888] = a[13] & g[10696];
assign g[27079] = b[13] & g[10696];
assign g[18889] = a[13] & g[10697];
assign g[27080] = b[13] & g[10697];
assign g[18890] = a[13] & g[10698];
assign g[27081] = b[13] & g[10698];
assign g[18891] = a[13] & g[10699];
assign g[27082] = b[13] & g[10699];
assign g[18892] = a[13] & g[10700];
assign g[27083] = b[13] & g[10700];
assign g[18893] = a[13] & g[10701];
assign g[27084] = b[13] & g[10701];
assign g[18894] = a[13] & g[10702];
assign g[27085] = b[13] & g[10702];
assign g[18895] = a[13] & g[10703];
assign g[27086] = b[13] & g[10703];
assign g[18896] = a[13] & g[10704];
assign g[27087] = b[13] & g[10704];
assign g[18897] = a[13] & g[10705];
assign g[27088] = b[13] & g[10705];
assign g[18898] = a[13] & g[10706];
assign g[27089] = b[13] & g[10706];
assign g[18899] = a[13] & g[10707];
assign g[27090] = b[13] & g[10707];
assign g[18900] = a[13] & g[10708];
assign g[27091] = b[13] & g[10708];
assign g[18901] = a[13] & g[10709];
assign g[27092] = b[13] & g[10709];
assign g[18902] = a[13] & g[10710];
assign g[27093] = b[13] & g[10710];
assign g[18903] = a[13] & g[10711];
assign g[27094] = b[13] & g[10711];
assign g[18904] = a[13] & g[10712];
assign g[27095] = b[13] & g[10712];
assign g[18905] = a[13] & g[10713];
assign g[27096] = b[13] & g[10713];
assign g[18906] = a[13] & g[10714];
assign g[27097] = b[13] & g[10714];
assign g[18907] = a[13] & g[10715];
assign g[27098] = b[13] & g[10715];
assign g[18908] = a[13] & g[10716];
assign g[27099] = b[13] & g[10716];
assign g[18909] = a[13] & g[10717];
assign g[27100] = b[13] & g[10717];
assign g[18910] = a[13] & g[10718];
assign g[27101] = b[13] & g[10718];
assign g[18911] = a[13] & g[10719];
assign g[27102] = b[13] & g[10719];
assign g[18912] = a[13] & g[10720];
assign g[27103] = b[13] & g[10720];
assign g[18913] = a[13] & g[10721];
assign g[27104] = b[13] & g[10721];
assign g[18914] = a[13] & g[10722];
assign g[27105] = b[13] & g[10722];
assign g[18915] = a[13] & g[10723];
assign g[27106] = b[13] & g[10723];
assign g[18916] = a[13] & g[10724];
assign g[27107] = b[13] & g[10724];
assign g[18917] = a[13] & g[10725];
assign g[27108] = b[13] & g[10725];
assign g[18918] = a[13] & g[10726];
assign g[27109] = b[13] & g[10726];
assign g[18919] = a[13] & g[10727];
assign g[27110] = b[13] & g[10727];
assign g[18920] = a[13] & g[10728];
assign g[27111] = b[13] & g[10728];
assign g[18921] = a[13] & g[10729];
assign g[27112] = b[13] & g[10729];
assign g[18922] = a[13] & g[10730];
assign g[27113] = b[13] & g[10730];
assign g[18923] = a[13] & g[10731];
assign g[27114] = b[13] & g[10731];
assign g[18924] = a[13] & g[10732];
assign g[27115] = b[13] & g[10732];
assign g[18925] = a[13] & g[10733];
assign g[27116] = b[13] & g[10733];
assign g[18926] = a[13] & g[10734];
assign g[27117] = b[13] & g[10734];
assign g[18927] = a[13] & g[10735];
assign g[27118] = b[13] & g[10735];
assign g[18928] = a[13] & g[10736];
assign g[27119] = b[13] & g[10736];
assign g[18929] = a[13] & g[10737];
assign g[27120] = b[13] & g[10737];
assign g[18930] = a[13] & g[10738];
assign g[27121] = b[13] & g[10738];
assign g[18931] = a[13] & g[10739];
assign g[27122] = b[13] & g[10739];
assign g[18932] = a[13] & g[10740];
assign g[27123] = b[13] & g[10740];
assign g[18933] = a[13] & g[10741];
assign g[27124] = b[13] & g[10741];
assign g[18934] = a[13] & g[10742];
assign g[27125] = b[13] & g[10742];
assign g[18935] = a[13] & g[10743];
assign g[27126] = b[13] & g[10743];
assign g[18936] = a[13] & g[10744];
assign g[27127] = b[13] & g[10744];
assign g[18937] = a[13] & g[10745];
assign g[27128] = b[13] & g[10745];
assign g[18938] = a[13] & g[10746];
assign g[27129] = b[13] & g[10746];
assign g[18939] = a[13] & g[10747];
assign g[27130] = b[13] & g[10747];
assign g[18940] = a[13] & g[10748];
assign g[27131] = b[13] & g[10748];
assign g[18941] = a[13] & g[10749];
assign g[27132] = b[13] & g[10749];
assign g[18942] = a[13] & g[10750];
assign g[27133] = b[13] & g[10750];
assign g[18943] = a[13] & g[10751];
assign g[27134] = b[13] & g[10751];
assign g[18944] = a[13] & g[10752];
assign g[27135] = b[13] & g[10752];
assign g[18945] = a[13] & g[10753];
assign g[27136] = b[13] & g[10753];
assign g[18946] = a[13] & g[10754];
assign g[27137] = b[13] & g[10754];
assign g[18947] = a[13] & g[10755];
assign g[27138] = b[13] & g[10755];
assign g[18948] = a[13] & g[10756];
assign g[27139] = b[13] & g[10756];
assign g[18949] = a[13] & g[10757];
assign g[27140] = b[13] & g[10757];
assign g[18950] = a[13] & g[10758];
assign g[27141] = b[13] & g[10758];
assign g[18951] = a[13] & g[10759];
assign g[27142] = b[13] & g[10759];
assign g[18952] = a[13] & g[10760];
assign g[27143] = b[13] & g[10760];
assign g[18953] = a[13] & g[10761];
assign g[27144] = b[13] & g[10761];
assign g[18954] = a[13] & g[10762];
assign g[27145] = b[13] & g[10762];
assign g[18955] = a[13] & g[10763];
assign g[27146] = b[13] & g[10763];
assign g[18956] = a[13] & g[10764];
assign g[27147] = b[13] & g[10764];
assign g[18957] = a[13] & g[10765];
assign g[27148] = b[13] & g[10765];
assign g[18958] = a[13] & g[10766];
assign g[27149] = b[13] & g[10766];
assign g[18959] = a[13] & g[10767];
assign g[27150] = b[13] & g[10767];
assign g[18960] = a[13] & g[10768];
assign g[27151] = b[13] & g[10768];
assign g[18961] = a[13] & g[10769];
assign g[27152] = b[13] & g[10769];
assign g[18962] = a[13] & g[10770];
assign g[27153] = b[13] & g[10770];
assign g[18963] = a[13] & g[10771];
assign g[27154] = b[13] & g[10771];
assign g[18964] = a[13] & g[10772];
assign g[27155] = b[13] & g[10772];
assign g[18965] = a[13] & g[10773];
assign g[27156] = b[13] & g[10773];
assign g[18966] = a[13] & g[10774];
assign g[27157] = b[13] & g[10774];
assign g[18967] = a[13] & g[10775];
assign g[27158] = b[13] & g[10775];
assign g[18968] = a[13] & g[10776];
assign g[27159] = b[13] & g[10776];
assign g[18969] = a[13] & g[10777];
assign g[27160] = b[13] & g[10777];
assign g[18970] = a[13] & g[10778];
assign g[27161] = b[13] & g[10778];
assign g[18971] = a[13] & g[10779];
assign g[27162] = b[13] & g[10779];
assign g[18972] = a[13] & g[10780];
assign g[27163] = b[13] & g[10780];
assign g[18973] = a[13] & g[10781];
assign g[27164] = b[13] & g[10781];
assign g[18974] = a[13] & g[10782];
assign g[27165] = b[13] & g[10782];
assign g[18975] = a[13] & g[10783];
assign g[27166] = b[13] & g[10783];
assign g[18976] = a[13] & g[10784];
assign g[27167] = b[13] & g[10784];
assign g[18977] = a[13] & g[10785];
assign g[27168] = b[13] & g[10785];
assign g[18978] = a[13] & g[10786];
assign g[27169] = b[13] & g[10786];
assign g[18979] = a[13] & g[10787];
assign g[27170] = b[13] & g[10787];
assign g[18980] = a[13] & g[10788];
assign g[27171] = b[13] & g[10788];
assign g[18981] = a[13] & g[10789];
assign g[27172] = b[13] & g[10789];
assign g[18982] = a[13] & g[10790];
assign g[27173] = b[13] & g[10790];
assign g[18983] = a[13] & g[10791];
assign g[27174] = b[13] & g[10791];
assign g[18984] = a[13] & g[10792];
assign g[27175] = b[13] & g[10792];
assign g[18985] = a[13] & g[10793];
assign g[27176] = b[13] & g[10793];
assign g[18986] = a[13] & g[10794];
assign g[27177] = b[13] & g[10794];
assign g[18987] = a[13] & g[10795];
assign g[27178] = b[13] & g[10795];
assign g[18988] = a[13] & g[10796];
assign g[27179] = b[13] & g[10796];
assign g[18989] = a[13] & g[10797];
assign g[27180] = b[13] & g[10797];
assign g[18990] = a[13] & g[10798];
assign g[27181] = b[13] & g[10798];
assign g[18991] = a[13] & g[10799];
assign g[27182] = b[13] & g[10799];
assign g[18992] = a[13] & g[10800];
assign g[27183] = b[13] & g[10800];
assign g[18993] = a[13] & g[10801];
assign g[27184] = b[13] & g[10801];
assign g[18994] = a[13] & g[10802];
assign g[27185] = b[13] & g[10802];
assign g[18995] = a[13] & g[10803];
assign g[27186] = b[13] & g[10803];
assign g[18996] = a[13] & g[10804];
assign g[27187] = b[13] & g[10804];
assign g[18997] = a[13] & g[10805];
assign g[27188] = b[13] & g[10805];
assign g[18998] = a[13] & g[10806];
assign g[27189] = b[13] & g[10806];
assign g[18999] = a[13] & g[10807];
assign g[27190] = b[13] & g[10807];
assign g[19000] = a[13] & g[10808];
assign g[27191] = b[13] & g[10808];
assign g[19001] = a[13] & g[10809];
assign g[27192] = b[13] & g[10809];
assign g[19002] = a[13] & g[10810];
assign g[27193] = b[13] & g[10810];
assign g[19003] = a[13] & g[10811];
assign g[27194] = b[13] & g[10811];
assign g[19004] = a[13] & g[10812];
assign g[27195] = b[13] & g[10812];
assign g[19005] = a[13] & g[10813];
assign g[27196] = b[13] & g[10813];
assign g[19006] = a[13] & g[10814];
assign g[27197] = b[13] & g[10814];
assign g[19007] = a[13] & g[10815];
assign g[27198] = b[13] & g[10815];
assign g[19008] = a[13] & g[10816];
assign g[27199] = b[13] & g[10816];
assign g[19009] = a[13] & g[10817];
assign g[27200] = b[13] & g[10817];
assign g[19010] = a[13] & g[10818];
assign g[27201] = b[13] & g[10818];
assign g[19011] = a[13] & g[10819];
assign g[27202] = b[13] & g[10819];
assign g[19012] = a[13] & g[10820];
assign g[27203] = b[13] & g[10820];
assign g[19013] = a[13] & g[10821];
assign g[27204] = b[13] & g[10821];
assign g[19014] = a[13] & g[10822];
assign g[27205] = b[13] & g[10822];
assign g[19015] = a[13] & g[10823];
assign g[27206] = b[13] & g[10823];
assign g[19016] = a[13] & g[10824];
assign g[27207] = b[13] & g[10824];
assign g[19017] = a[13] & g[10825];
assign g[27208] = b[13] & g[10825];
assign g[19018] = a[13] & g[10826];
assign g[27209] = b[13] & g[10826];
assign g[19019] = a[13] & g[10827];
assign g[27210] = b[13] & g[10827];
assign g[19020] = a[13] & g[10828];
assign g[27211] = b[13] & g[10828];
assign g[19021] = a[13] & g[10829];
assign g[27212] = b[13] & g[10829];
assign g[19022] = a[13] & g[10830];
assign g[27213] = b[13] & g[10830];
assign g[19023] = a[13] & g[10831];
assign g[27214] = b[13] & g[10831];
assign g[19024] = a[13] & g[10832];
assign g[27215] = b[13] & g[10832];
assign g[19025] = a[13] & g[10833];
assign g[27216] = b[13] & g[10833];
assign g[19026] = a[13] & g[10834];
assign g[27217] = b[13] & g[10834];
assign g[19027] = a[13] & g[10835];
assign g[27218] = b[13] & g[10835];
assign g[19028] = a[13] & g[10836];
assign g[27219] = b[13] & g[10836];
assign g[19029] = a[13] & g[10837];
assign g[27220] = b[13] & g[10837];
assign g[19030] = a[13] & g[10838];
assign g[27221] = b[13] & g[10838];
assign g[19031] = a[13] & g[10839];
assign g[27222] = b[13] & g[10839];
assign g[19032] = a[13] & g[10840];
assign g[27223] = b[13] & g[10840];
assign g[19033] = a[13] & g[10841];
assign g[27224] = b[13] & g[10841];
assign g[19034] = a[13] & g[10842];
assign g[27225] = b[13] & g[10842];
assign g[19035] = a[13] & g[10843];
assign g[27226] = b[13] & g[10843];
assign g[19036] = a[13] & g[10844];
assign g[27227] = b[13] & g[10844];
assign g[19037] = a[13] & g[10845];
assign g[27228] = b[13] & g[10845];
assign g[19038] = a[13] & g[10846];
assign g[27229] = b[13] & g[10846];
assign g[19039] = a[13] & g[10847];
assign g[27230] = b[13] & g[10847];
assign g[19040] = a[13] & g[10848];
assign g[27231] = b[13] & g[10848];
assign g[19041] = a[13] & g[10849];
assign g[27232] = b[13] & g[10849];
assign g[19042] = a[13] & g[10850];
assign g[27233] = b[13] & g[10850];
assign g[19043] = a[13] & g[10851];
assign g[27234] = b[13] & g[10851];
assign g[19044] = a[13] & g[10852];
assign g[27235] = b[13] & g[10852];
assign g[19045] = a[13] & g[10853];
assign g[27236] = b[13] & g[10853];
assign g[19046] = a[13] & g[10854];
assign g[27237] = b[13] & g[10854];
assign g[19047] = a[13] & g[10855];
assign g[27238] = b[13] & g[10855];
assign g[19048] = a[13] & g[10856];
assign g[27239] = b[13] & g[10856];
assign g[19049] = a[13] & g[10857];
assign g[27240] = b[13] & g[10857];
assign g[19050] = a[13] & g[10858];
assign g[27241] = b[13] & g[10858];
assign g[19051] = a[13] & g[10859];
assign g[27242] = b[13] & g[10859];
assign g[19052] = a[13] & g[10860];
assign g[27243] = b[13] & g[10860];
assign g[19053] = a[13] & g[10861];
assign g[27244] = b[13] & g[10861];
assign g[19054] = a[13] & g[10862];
assign g[27245] = b[13] & g[10862];
assign g[19055] = a[13] & g[10863];
assign g[27246] = b[13] & g[10863];
assign g[19056] = a[13] & g[10864];
assign g[27247] = b[13] & g[10864];
assign g[19057] = a[13] & g[10865];
assign g[27248] = b[13] & g[10865];
assign g[19058] = a[13] & g[10866];
assign g[27249] = b[13] & g[10866];
assign g[19059] = a[13] & g[10867];
assign g[27250] = b[13] & g[10867];
assign g[19060] = a[13] & g[10868];
assign g[27251] = b[13] & g[10868];
assign g[19061] = a[13] & g[10869];
assign g[27252] = b[13] & g[10869];
assign g[19062] = a[13] & g[10870];
assign g[27253] = b[13] & g[10870];
assign g[19063] = a[13] & g[10871];
assign g[27254] = b[13] & g[10871];
assign g[19064] = a[13] & g[10872];
assign g[27255] = b[13] & g[10872];
assign g[19065] = a[13] & g[10873];
assign g[27256] = b[13] & g[10873];
assign g[19066] = a[13] & g[10874];
assign g[27257] = b[13] & g[10874];
assign g[19067] = a[13] & g[10875];
assign g[27258] = b[13] & g[10875];
assign g[19068] = a[13] & g[10876];
assign g[27259] = b[13] & g[10876];
assign g[19069] = a[13] & g[10877];
assign g[27260] = b[13] & g[10877];
assign g[19070] = a[13] & g[10878];
assign g[27261] = b[13] & g[10878];
assign g[19071] = a[13] & g[10879];
assign g[27262] = b[13] & g[10879];
assign g[19072] = a[13] & g[10880];
assign g[27263] = b[13] & g[10880];
assign g[19073] = a[13] & g[10881];
assign g[27264] = b[13] & g[10881];
assign g[19074] = a[13] & g[10882];
assign g[27265] = b[13] & g[10882];
assign g[19075] = a[13] & g[10883];
assign g[27266] = b[13] & g[10883];
assign g[19076] = a[13] & g[10884];
assign g[27267] = b[13] & g[10884];
assign g[19077] = a[13] & g[10885];
assign g[27268] = b[13] & g[10885];
assign g[19078] = a[13] & g[10886];
assign g[27269] = b[13] & g[10886];
assign g[19079] = a[13] & g[10887];
assign g[27270] = b[13] & g[10887];
assign g[19080] = a[13] & g[10888];
assign g[27271] = b[13] & g[10888];
assign g[19081] = a[13] & g[10889];
assign g[27272] = b[13] & g[10889];
assign g[19082] = a[13] & g[10890];
assign g[27273] = b[13] & g[10890];
assign g[19083] = a[13] & g[10891];
assign g[27274] = b[13] & g[10891];
assign g[19084] = a[13] & g[10892];
assign g[27275] = b[13] & g[10892];
assign g[19085] = a[13] & g[10893];
assign g[27276] = b[13] & g[10893];
assign g[19086] = a[13] & g[10894];
assign g[27277] = b[13] & g[10894];
assign g[19087] = a[13] & g[10895];
assign g[27278] = b[13] & g[10895];
assign g[19088] = a[13] & g[10896];
assign g[27279] = b[13] & g[10896];
assign g[19089] = a[13] & g[10897];
assign g[27280] = b[13] & g[10897];
assign g[19090] = a[13] & g[10898];
assign g[27281] = b[13] & g[10898];
assign g[19091] = a[13] & g[10899];
assign g[27282] = b[13] & g[10899];
assign g[19092] = a[13] & g[10900];
assign g[27283] = b[13] & g[10900];
assign g[19093] = a[13] & g[10901];
assign g[27284] = b[13] & g[10901];
assign g[19094] = a[13] & g[10902];
assign g[27285] = b[13] & g[10902];
assign g[19095] = a[13] & g[10903];
assign g[27286] = b[13] & g[10903];
assign g[19096] = a[13] & g[10904];
assign g[27287] = b[13] & g[10904];
assign g[19097] = a[13] & g[10905];
assign g[27288] = b[13] & g[10905];
assign g[19098] = a[13] & g[10906];
assign g[27289] = b[13] & g[10906];
assign g[19099] = a[13] & g[10907];
assign g[27290] = b[13] & g[10907];
assign g[19100] = a[13] & g[10908];
assign g[27291] = b[13] & g[10908];
assign g[19101] = a[13] & g[10909];
assign g[27292] = b[13] & g[10909];
assign g[19102] = a[13] & g[10910];
assign g[27293] = b[13] & g[10910];
assign g[19103] = a[13] & g[10911];
assign g[27294] = b[13] & g[10911];
assign g[19104] = a[13] & g[10912];
assign g[27295] = b[13] & g[10912];
assign g[19105] = a[13] & g[10913];
assign g[27296] = b[13] & g[10913];
assign g[19106] = a[13] & g[10914];
assign g[27297] = b[13] & g[10914];
assign g[19107] = a[13] & g[10915];
assign g[27298] = b[13] & g[10915];
assign g[19108] = a[13] & g[10916];
assign g[27299] = b[13] & g[10916];
assign g[19109] = a[13] & g[10917];
assign g[27300] = b[13] & g[10917];
assign g[19110] = a[13] & g[10918];
assign g[27301] = b[13] & g[10918];
assign g[19111] = a[13] & g[10919];
assign g[27302] = b[13] & g[10919];
assign g[19112] = a[13] & g[10920];
assign g[27303] = b[13] & g[10920];
assign g[19113] = a[13] & g[10921];
assign g[27304] = b[13] & g[10921];
assign g[19114] = a[13] & g[10922];
assign g[27305] = b[13] & g[10922];
assign g[19115] = a[13] & g[10923];
assign g[27306] = b[13] & g[10923];
assign g[19116] = a[13] & g[10924];
assign g[27307] = b[13] & g[10924];
assign g[19117] = a[13] & g[10925];
assign g[27308] = b[13] & g[10925];
assign g[19118] = a[13] & g[10926];
assign g[27309] = b[13] & g[10926];
assign g[19119] = a[13] & g[10927];
assign g[27310] = b[13] & g[10927];
assign g[19120] = a[13] & g[10928];
assign g[27311] = b[13] & g[10928];
assign g[19121] = a[13] & g[10929];
assign g[27312] = b[13] & g[10929];
assign g[19122] = a[13] & g[10930];
assign g[27313] = b[13] & g[10930];
assign g[19123] = a[13] & g[10931];
assign g[27314] = b[13] & g[10931];
assign g[19124] = a[13] & g[10932];
assign g[27315] = b[13] & g[10932];
assign g[19125] = a[13] & g[10933];
assign g[27316] = b[13] & g[10933];
assign g[19126] = a[13] & g[10934];
assign g[27317] = b[13] & g[10934];
assign g[19127] = a[13] & g[10935];
assign g[27318] = b[13] & g[10935];
assign g[19128] = a[13] & g[10936];
assign g[27319] = b[13] & g[10936];
assign g[19129] = a[13] & g[10937];
assign g[27320] = b[13] & g[10937];
assign g[19130] = a[13] & g[10938];
assign g[27321] = b[13] & g[10938];
assign g[19131] = a[13] & g[10939];
assign g[27322] = b[13] & g[10939];
assign g[19132] = a[13] & g[10940];
assign g[27323] = b[13] & g[10940];
assign g[19133] = a[13] & g[10941];
assign g[27324] = b[13] & g[10941];
assign g[19134] = a[13] & g[10942];
assign g[27325] = b[13] & g[10942];
assign g[19135] = a[13] & g[10943];
assign g[27326] = b[13] & g[10943];
assign g[19136] = a[13] & g[10944];
assign g[27327] = b[13] & g[10944];
assign g[19137] = a[13] & g[10945];
assign g[27328] = b[13] & g[10945];
assign g[19138] = a[13] & g[10946];
assign g[27329] = b[13] & g[10946];
assign g[19139] = a[13] & g[10947];
assign g[27330] = b[13] & g[10947];
assign g[19140] = a[13] & g[10948];
assign g[27331] = b[13] & g[10948];
assign g[19141] = a[13] & g[10949];
assign g[27332] = b[13] & g[10949];
assign g[19142] = a[13] & g[10950];
assign g[27333] = b[13] & g[10950];
assign g[19143] = a[13] & g[10951];
assign g[27334] = b[13] & g[10951];
assign g[19144] = a[13] & g[10952];
assign g[27335] = b[13] & g[10952];
assign g[19145] = a[13] & g[10953];
assign g[27336] = b[13] & g[10953];
assign g[19146] = a[13] & g[10954];
assign g[27337] = b[13] & g[10954];
assign g[19147] = a[13] & g[10955];
assign g[27338] = b[13] & g[10955];
assign g[19148] = a[13] & g[10956];
assign g[27339] = b[13] & g[10956];
assign g[19149] = a[13] & g[10957];
assign g[27340] = b[13] & g[10957];
assign g[19150] = a[13] & g[10958];
assign g[27341] = b[13] & g[10958];
assign g[19151] = a[13] & g[10959];
assign g[27342] = b[13] & g[10959];
assign g[19152] = a[13] & g[10960];
assign g[27343] = b[13] & g[10960];
assign g[19153] = a[13] & g[10961];
assign g[27344] = b[13] & g[10961];
assign g[19154] = a[13] & g[10962];
assign g[27345] = b[13] & g[10962];
assign g[19155] = a[13] & g[10963];
assign g[27346] = b[13] & g[10963];
assign g[19156] = a[13] & g[10964];
assign g[27347] = b[13] & g[10964];
assign g[19157] = a[13] & g[10965];
assign g[27348] = b[13] & g[10965];
assign g[19158] = a[13] & g[10966];
assign g[27349] = b[13] & g[10966];
assign g[19159] = a[13] & g[10967];
assign g[27350] = b[13] & g[10967];
assign g[19160] = a[13] & g[10968];
assign g[27351] = b[13] & g[10968];
assign g[19161] = a[13] & g[10969];
assign g[27352] = b[13] & g[10969];
assign g[19162] = a[13] & g[10970];
assign g[27353] = b[13] & g[10970];
assign g[19163] = a[13] & g[10971];
assign g[27354] = b[13] & g[10971];
assign g[19164] = a[13] & g[10972];
assign g[27355] = b[13] & g[10972];
assign g[19165] = a[13] & g[10973];
assign g[27356] = b[13] & g[10973];
assign g[19166] = a[13] & g[10974];
assign g[27357] = b[13] & g[10974];
assign g[19167] = a[13] & g[10975];
assign g[27358] = b[13] & g[10975];
assign g[19168] = a[13] & g[10976];
assign g[27359] = b[13] & g[10976];
assign g[19169] = a[13] & g[10977];
assign g[27360] = b[13] & g[10977];
assign g[19170] = a[13] & g[10978];
assign g[27361] = b[13] & g[10978];
assign g[19171] = a[13] & g[10979];
assign g[27362] = b[13] & g[10979];
assign g[19172] = a[13] & g[10980];
assign g[27363] = b[13] & g[10980];
assign g[19173] = a[13] & g[10981];
assign g[27364] = b[13] & g[10981];
assign g[19174] = a[13] & g[10982];
assign g[27365] = b[13] & g[10982];
assign g[19175] = a[13] & g[10983];
assign g[27366] = b[13] & g[10983];
assign g[19176] = a[13] & g[10984];
assign g[27367] = b[13] & g[10984];
assign g[19177] = a[13] & g[10985];
assign g[27368] = b[13] & g[10985];
assign g[19178] = a[13] & g[10986];
assign g[27369] = b[13] & g[10986];
assign g[19179] = a[13] & g[10987];
assign g[27370] = b[13] & g[10987];
assign g[19180] = a[13] & g[10988];
assign g[27371] = b[13] & g[10988];
assign g[19181] = a[13] & g[10989];
assign g[27372] = b[13] & g[10989];
assign g[19182] = a[13] & g[10990];
assign g[27373] = b[13] & g[10990];
assign g[19183] = a[13] & g[10991];
assign g[27374] = b[13] & g[10991];
assign g[19184] = a[13] & g[10992];
assign g[27375] = b[13] & g[10992];
assign g[19185] = a[13] & g[10993];
assign g[27376] = b[13] & g[10993];
assign g[19186] = a[13] & g[10994];
assign g[27377] = b[13] & g[10994];
assign g[19187] = a[13] & g[10995];
assign g[27378] = b[13] & g[10995];
assign g[19188] = a[13] & g[10996];
assign g[27379] = b[13] & g[10996];
assign g[19189] = a[13] & g[10997];
assign g[27380] = b[13] & g[10997];
assign g[19190] = a[13] & g[10998];
assign g[27381] = b[13] & g[10998];
assign g[19191] = a[13] & g[10999];
assign g[27382] = b[13] & g[10999];
assign g[19192] = a[13] & g[11000];
assign g[27383] = b[13] & g[11000];
assign g[19193] = a[13] & g[11001];
assign g[27384] = b[13] & g[11001];
assign g[19194] = a[13] & g[11002];
assign g[27385] = b[13] & g[11002];
assign g[19195] = a[13] & g[11003];
assign g[27386] = b[13] & g[11003];
assign g[19196] = a[13] & g[11004];
assign g[27387] = b[13] & g[11004];
assign g[19197] = a[13] & g[11005];
assign g[27388] = b[13] & g[11005];
assign g[19198] = a[13] & g[11006];
assign g[27389] = b[13] & g[11006];
assign g[19199] = a[13] & g[11007];
assign g[27390] = b[13] & g[11007];
assign g[19200] = a[13] & g[11008];
assign g[27391] = b[13] & g[11008];
assign g[19201] = a[13] & g[11009];
assign g[27392] = b[13] & g[11009];
assign g[19202] = a[13] & g[11010];
assign g[27393] = b[13] & g[11010];
assign g[19203] = a[13] & g[11011];
assign g[27394] = b[13] & g[11011];
assign g[19204] = a[13] & g[11012];
assign g[27395] = b[13] & g[11012];
assign g[19205] = a[13] & g[11013];
assign g[27396] = b[13] & g[11013];
assign g[19206] = a[13] & g[11014];
assign g[27397] = b[13] & g[11014];
assign g[19207] = a[13] & g[11015];
assign g[27398] = b[13] & g[11015];
assign g[19208] = a[13] & g[11016];
assign g[27399] = b[13] & g[11016];
assign g[19209] = a[13] & g[11017];
assign g[27400] = b[13] & g[11017];
assign g[19210] = a[13] & g[11018];
assign g[27401] = b[13] & g[11018];
assign g[19211] = a[13] & g[11019];
assign g[27402] = b[13] & g[11019];
assign g[19212] = a[13] & g[11020];
assign g[27403] = b[13] & g[11020];
assign g[19213] = a[13] & g[11021];
assign g[27404] = b[13] & g[11021];
assign g[19214] = a[13] & g[11022];
assign g[27405] = b[13] & g[11022];
assign g[19215] = a[13] & g[11023];
assign g[27406] = b[13] & g[11023];
assign g[19216] = a[13] & g[11024];
assign g[27407] = b[13] & g[11024];
assign g[19217] = a[13] & g[11025];
assign g[27408] = b[13] & g[11025];
assign g[19218] = a[13] & g[11026];
assign g[27409] = b[13] & g[11026];
assign g[19219] = a[13] & g[11027];
assign g[27410] = b[13] & g[11027];
assign g[19220] = a[13] & g[11028];
assign g[27411] = b[13] & g[11028];
assign g[19221] = a[13] & g[11029];
assign g[27412] = b[13] & g[11029];
assign g[19222] = a[13] & g[11030];
assign g[27413] = b[13] & g[11030];
assign g[19223] = a[13] & g[11031];
assign g[27414] = b[13] & g[11031];
assign g[19224] = a[13] & g[11032];
assign g[27415] = b[13] & g[11032];
assign g[19225] = a[13] & g[11033];
assign g[27416] = b[13] & g[11033];
assign g[19226] = a[13] & g[11034];
assign g[27417] = b[13] & g[11034];
assign g[19227] = a[13] & g[11035];
assign g[27418] = b[13] & g[11035];
assign g[19228] = a[13] & g[11036];
assign g[27419] = b[13] & g[11036];
assign g[19229] = a[13] & g[11037];
assign g[27420] = b[13] & g[11037];
assign g[19230] = a[13] & g[11038];
assign g[27421] = b[13] & g[11038];
assign g[19231] = a[13] & g[11039];
assign g[27422] = b[13] & g[11039];
assign g[19232] = a[13] & g[11040];
assign g[27423] = b[13] & g[11040];
assign g[19233] = a[13] & g[11041];
assign g[27424] = b[13] & g[11041];
assign g[19234] = a[13] & g[11042];
assign g[27425] = b[13] & g[11042];
assign g[19235] = a[13] & g[11043];
assign g[27426] = b[13] & g[11043];
assign g[19236] = a[13] & g[11044];
assign g[27427] = b[13] & g[11044];
assign g[19237] = a[13] & g[11045];
assign g[27428] = b[13] & g[11045];
assign g[19238] = a[13] & g[11046];
assign g[27429] = b[13] & g[11046];
assign g[19239] = a[13] & g[11047];
assign g[27430] = b[13] & g[11047];
assign g[19240] = a[13] & g[11048];
assign g[27431] = b[13] & g[11048];
assign g[19241] = a[13] & g[11049];
assign g[27432] = b[13] & g[11049];
assign g[19242] = a[13] & g[11050];
assign g[27433] = b[13] & g[11050];
assign g[19243] = a[13] & g[11051];
assign g[27434] = b[13] & g[11051];
assign g[19244] = a[13] & g[11052];
assign g[27435] = b[13] & g[11052];
assign g[19245] = a[13] & g[11053];
assign g[27436] = b[13] & g[11053];
assign g[19246] = a[13] & g[11054];
assign g[27437] = b[13] & g[11054];
assign g[19247] = a[13] & g[11055];
assign g[27438] = b[13] & g[11055];
assign g[19248] = a[13] & g[11056];
assign g[27439] = b[13] & g[11056];
assign g[19249] = a[13] & g[11057];
assign g[27440] = b[13] & g[11057];
assign g[19250] = a[13] & g[11058];
assign g[27441] = b[13] & g[11058];
assign g[19251] = a[13] & g[11059];
assign g[27442] = b[13] & g[11059];
assign g[19252] = a[13] & g[11060];
assign g[27443] = b[13] & g[11060];
assign g[19253] = a[13] & g[11061];
assign g[27444] = b[13] & g[11061];
assign g[19254] = a[13] & g[11062];
assign g[27445] = b[13] & g[11062];
assign g[19255] = a[13] & g[11063];
assign g[27446] = b[13] & g[11063];
assign g[19256] = a[13] & g[11064];
assign g[27447] = b[13] & g[11064];
assign g[19257] = a[13] & g[11065];
assign g[27448] = b[13] & g[11065];
assign g[19258] = a[13] & g[11066];
assign g[27449] = b[13] & g[11066];
assign g[19259] = a[13] & g[11067];
assign g[27450] = b[13] & g[11067];
assign g[19260] = a[13] & g[11068];
assign g[27451] = b[13] & g[11068];
assign g[19261] = a[13] & g[11069];
assign g[27452] = b[13] & g[11069];
assign g[19262] = a[13] & g[11070];
assign g[27453] = b[13] & g[11070];
assign g[19263] = a[13] & g[11071];
assign g[27454] = b[13] & g[11071];
assign g[19264] = a[13] & g[11072];
assign g[27455] = b[13] & g[11072];
assign g[19265] = a[13] & g[11073];
assign g[27456] = b[13] & g[11073];
assign g[19266] = a[13] & g[11074];
assign g[27457] = b[13] & g[11074];
assign g[19267] = a[13] & g[11075];
assign g[27458] = b[13] & g[11075];
assign g[19268] = a[13] & g[11076];
assign g[27459] = b[13] & g[11076];
assign g[19269] = a[13] & g[11077];
assign g[27460] = b[13] & g[11077];
assign g[19270] = a[13] & g[11078];
assign g[27461] = b[13] & g[11078];
assign g[19271] = a[13] & g[11079];
assign g[27462] = b[13] & g[11079];
assign g[19272] = a[13] & g[11080];
assign g[27463] = b[13] & g[11080];
assign g[19273] = a[13] & g[11081];
assign g[27464] = b[13] & g[11081];
assign g[19274] = a[13] & g[11082];
assign g[27465] = b[13] & g[11082];
assign g[19275] = a[13] & g[11083];
assign g[27466] = b[13] & g[11083];
assign g[19276] = a[13] & g[11084];
assign g[27467] = b[13] & g[11084];
assign g[19277] = a[13] & g[11085];
assign g[27468] = b[13] & g[11085];
assign g[19278] = a[13] & g[11086];
assign g[27469] = b[13] & g[11086];
assign g[19279] = a[13] & g[11087];
assign g[27470] = b[13] & g[11087];
assign g[19280] = a[13] & g[11088];
assign g[27471] = b[13] & g[11088];
assign g[19281] = a[13] & g[11089];
assign g[27472] = b[13] & g[11089];
assign g[19282] = a[13] & g[11090];
assign g[27473] = b[13] & g[11090];
assign g[19283] = a[13] & g[11091];
assign g[27474] = b[13] & g[11091];
assign g[19284] = a[13] & g[11092];
assign g[27475] = b[13] & g[11092];
assign g[19285] = a[13] & g[11093];
assign g[27476] = b[13] & g[11093];
assign g[19286] = a[13] & g[11094];
assign g[27477] = b[13] & g[11094];
assign g[19287] = a[13] & g[11095];
assign g[27478] = b[13] & g[11095];
assign g[19288] = a[13] & g[11096];
assign g[27479] = b[13] & g[11096];
assign g[19289] = a[13] & g[11097];
assign g[27480] = b[13] & g[11097];
assign g[19290] = a[13] & g[11098];
assign g[27481] = b[13] & g[11098];
assign g[19291] = a[13] & g[11099];
assign g[27482] = b[13] & g[11099];
assign g[19292] = a[13] & g[11100];
assign g[27483] = b[13] & g[11100];
assign g[19293] = a[13] & g[11101];
assign g[27484] = b[13] & g[11101];
assign g[19294] = a[13] & g[11102];
assign g[27485] = b[13] & g[11102];
assign g[19295] = a[13] & g[11103];
assign g[27486] = b[13] & g[11103];
assign g[19296] = a[13] & g[11104];
assign g[27487] = b[13] & g[11104];
assign g[19297] = a[13] & g[11105];
assign g[27488] = b[13] & g[11105];
assign g[19298] = a[13] & g[11106];
assign g[27489] = b[13] & g[11106];
assign g[19299] = a[13] & g[11107];
assign g[27490] = b[13] & g[11107];
assign g[19300] = a[13] & g[11108];
assign g[27491] = b[13] & g[11108];
assign g[19301] = a[13] & g[11109];
assign g[27492] = b[13] & g[11109];
assign g[19302] = a[13] & g[11110];
assign g[27493] = b[13] & g[11110];
assign g[19303] = a[13] & g[11111];
assign g[27494] = b[13] & g[11111];
assign g[19304] = a[13] & g[11112];
assign g[27495] = b[13] & g[11112];
assign g[19305] = a[13] & g[11113];
assign g[27496] = b[13] & g[11113];
assign g[19306] = a[13] & g[11114];
assign g[27497] = b[13] & g[11114];
assign g[19307] = a[13] & g[11115];
assign g[27498] = b[13] & g[11115];
assign g[19308] = a[13] & g[11116];
assign g[27499] = b[13] & g[11116];
assign g[19309] = a[13] & g[11117];
assign g[27500] = b[13] & g[11117];
assign g[19310] = a[13] & g[11118];
assign g[27501] = b[13] & g[11118];
assign g[19311] = a[13] & g[11119];
assign g[27502] = b[13] & g[11119];
assign g[19312] = a[13] & g[11120];
assign g[27503] = b[13] & g[11120];
assign g[19313] = a[13] & g[11121];
assign g[27504] = b[13] & g[11121];
assign g[19314] = a[13] & g[11122];
assign g[27505] = b[13] & g[11122];
assign g[19315] = a[13] & g[11123];
assign g[27506] = b[13] & g[11123];
assign g[19316] = a[13] & g[11124];
assign g[27507] = b[13] & g[11124];
assign g[19317] = a[13] & g[11125];
assign g[27508] = b[13] & g[11125];
assign g[19318] = a[13] & g[11126];
assign g[27509] = b[13] & g[11126];
assign g[19319] = a[13] & g[11127];
assign g[27510] = b[13] & g[11127];
assign g[19320] = a[13] & g[11128];
assign g[27511] = b[13] & g[11128];
assign g[19321] = a[13] & g[11129];
assign g[27512] = b[13] & g[11129];
assign g[19322] = a[13] & g[11130];
assign g[27513] = b[13] & g[11130];
assign g[19323] = a[13] & g[11131];
assign g[27514] = b[13] & g[11131];
assign g[19324] = a[13] & g[11132];
assign g[27515] = b[13] & g[11132];
assign g[19325] = a[13] & g[11133];
assign g[27516] = b[13] & g[11133];
assign g[19326] = a[13] & g[11134];
assign g[27517] = b[13] & g[11134];
assign g[19327] = a[13] & g[11135];
assign g[27518] = b[13] & g[11135];
assign g[19328] = a[13] & g[11136];
assign g[27519] = b[13] & g[11136];
assign g[19329] = a[13] & g[11137];
assign g[27520] = b[13] & g[11137];
assign g[19330] = a[13] & g[11138];
assign g[27521] = b[13] & g[11138];
assign g[19331] = a[13] & g[11139];
assign g[27522] = b[13] & g[11139];
assign g[19332] = a[13] & g[11140];
assign g[27523] = b[13] & g[11140];
assign g[19333] = a[13] & g[11141];
assign g[27524] = b[13] & g[11141];
assign g[19334] = a[13] & g[11142];
assign g[27525] = b[13] & g[11142];
assign g[19335] = a[13] & g[11143];
assign g[27526] = b[13] & g[11143];
assign g[19336] = a[13] & g[11144];
assign g[27527] = b[13] & g[11144];
assign g[19337] = a[13] & g[11145];
assign g[27528] = b[13] & g[11145];
assign g[19338] = a[13] & g[11146];
assign g[27529] = b[13] & g[11146];
assign g[19339] = a[13] & g[11147];
assign g[27530] = b[13] & g[11147];
assign g[19340] = a[13] & g[11148];
assign g[27531] = b[13] & g[11148];
assign g[19341] = a[13] & g[11149];
assign g[27532] = b[13] & g[11149];
assign g[19342] = a[13] & g[11150];
assign g[27533] = b[13] & g[11150];
assign g[19343] = a[13] & g[11151];
assign g[27534] = b[13] & g[11151];
assign g[19344] = a[13] & g[11152];
assign g[27535] = b[13] & g[11152];
assign g[19345] = a[13] & g[11153];
assign g[27536] = b[13] & g[11153];
assign g[19346] = a[13] & g[11154];
assign g[27537] = b[13] & g[11154];
assign g[19347] = a[13] & g[11155];
assign g[27538] = b[13] & g[11155];
assign g[19348] = a[13] & g[11156];
assign g[27539] = b[13] & g[11156];
assign g[19349] = a[13] & g[11157];
assign g[27540] = b[13] & g[11157];
assign g[19350] = a[13] & g[11158];
assign g[27541] = b[13] & g[11158];
assign g[19351] = a[13] & g[11159];
assign g[27542] = b[13] & g[11159];
assign g[19352] = a[13] & g[11160];
assign g[27543] = b[13] & g[11160];
assign g[19353] = a[13] & g[11161];
assign g[27544] = b[13] & g[11161];
assign g[19354] = a[13] & g[11162];
assign g[27545] = b[13] & g[11162];
assign g[19355] = a[13] & g[11163];
assign g[27546] = b[13] & g[11163];
assign g[19356] = a[13] & g[11164];
assign g[27547] = b[13] & g[11164];
assign g[19357] = a[13] & g[11165];
assign g[27548] = b[13] & g[11165];
assign g[19358] = a[13] & g[11166];
assign g[27549] = b[13] & g[11166];
assign g[19359] = a[13] & g[11167];
assign g[27550] = b[13] & g[11167];
assign g[19360] = a[13] & g[11168];
assign g[27551] = b[13] & g[11168];
assign g[19361] = a[13] & g[11169];
assign g[27552] = b[13] & g[11169];
assign g[19362] = a[13] & g[11170];
assign g[27553] = b[13] & g[11170];
assign g[19363] = a[13] & g[11171];
assign g[27554] = b[13] & g[11171];
assign g[19364] = a[13] & g[11172];
assign g[27555] = b[13] & g[11172];
assign g[19365] = a[13] & g[11173];
assign g[27556] = b[13] & g[11173];
assign g[19366] = a[13] & g[11174];
assign g[27557] = b[13] & g[11174];
assign g[19367] = a[13] & g[11175];
assign g[27558] = b[13] & g[11175];
assign g[19368] = a[13] & g[11176];
assign g[27559] = b[13] & g[11176];
assign g[19369] = a[13] & g[11177];
assign g[27560] = b[13] & g[11177];
assign g[19370] = a[13] & g[11178];
assign g[27561] = b[13] & g[11178];
assign g[19371] = a[13] & g[11179];
assign g[27562] = b[13] & g[11179];
assign g[19372] = a[13] & g[11180];
assign g[27563] = b[13] & g[11180];
assign g[19373] = a[13] & g[11181];
assign g[27564] = b[13] & g[11181];
assign g[19374] = a[13] & g[11182];
assign g[27565] = b[13] & g[11182];
assign g[19375] = a[13] & g[11183];
assign g[27566] = b[13] & g[11183];
assign g[19376] = a[13] & g[11184];
assign g[27567] = b[13] & g[11184];
assign g[19377] = a[13] & g[11185];
assign g[27568] = b[13] & g[11185];
assign g[19378] = a[13] & g[11186];
assign g[27569] = b[13] & g[11186];
assign g[19379] = a[13] & g[11187];
assign g[27570] = b[13] & g[11187];
assign g[19380] = a[13] & g[11188];
assign g[27571] = b[13] & g[11188];
assign g[19381] = a[13] & g[11189];
assign g[27572] = b[13] & g[11189];
assign g[19382] = a[13] & g[11190];
assign g[27573] = b[13] & g[11190];
assign g[19383] = a[13] & g[11191];
assign g[27574] = b[13] & g[11191];
assign g[19384] = a[13] & g[11192];
assign g[27575] = b[13] & g[11192];
assign g[19385] = a[13] & g[11193];
assign g[27576] = b[13] & g[11193];
assign g[19386] = a[13] & g[11194];
assign g[27577] = b[13] & g[11194];
assign g[19387] = a[13] & g[11195];
assign g[27578] = b[13] & g[11195];
assign g[19388] = a[13] & g[11196];
assign g[27579] = b[13] & g[11196];
assign g[19389] = a[13] & g[11197];
assign g[27580] = b[13] & g[11197];
assign g[19390] = a[13] & g[11198];
assign g[27581] = b[13] & g[11198];
assign g[19391] = a[13] & g[11199];
assign g[27582] = b[13] & g[11199];
assign g[19392] = a[13] & g[11200];
assign g[27583] = b[13] & g[11200];
assign g[19393] = a[13] & g[11201];
assign g[27584] = b[13] & g[11201];
assign g[19394] = a[13] & g[11202];
assign g[27585] = b[13] & g[11202];
assign g[19395] = a[13] & g[11203];
assign g[27586] = b[13] & g[11203];
assign g[19396] = a[13] & g[11204];
assign g[27587] = b[13] & g[11204];
assign g[19397] = a[13] & g[11205];
assign g[27588] = b[13] & g[11205];
assign g[19398] = a[13] & g[11206];
assign g[27589] = b[13] & g[11206];
assign g[19399] = a[13] & g[11207];
assign g[27590] = b[13] & g[11207];
assign g[19400] = a[13] & g[11208];
assign g[27591] = b[13] & g[11208];
assign g[19401] = a[13] & g[11209];
assign g[27592] = b[13] & g[11209];
assign g[19402] = a[13] & g[11210];
assign g[27593] = b[13] & g[11210];
assign g[19403] = a[13] & g[11211];
assign g[27594] = b[13] & g[11211];
assign g[19404] = a[13] & g[11212];
assign g[27595] = b[13] & g[11212];
assign g[19405] = a[13] & g[11213];
assign g[27596] = b[13] & g[11213];
assign g[19406] = a[13] & g[11214];
assign g[27597] = b[13] & g[11214];
assign g[19407] = a[13] & g[11215];
assign g[27598] = b[13] & g[11215];
assign g[19408] = a[13] & g[11216];
assign g[27599] = b[13] & g[11216];
assign g[19409] = a[13] & g[11217];
assign g[27600] = b[13] & g[11217];
assign g[19410] = a[13] & g[11218];
assign g[27601] = b[13] & g[11218];
assign g[19411] = a[13] & g[11219];
assign g[27602] = b[13] & g[11219];
assign g[19412] = a[13] & g[11220];
assign g[27603] = b[13] & g[11220];
assign g[19413] = a[13] & g[11221];
assign g[27604] = b[13] & g[11221];
assign g[19414] = a[13] & g[11222];
assign g[27605] = b[13] & g[11222];
assign g[19415] = a[13] & g[11223];
assign g[27606] = b[13] & g[11223];
assign g[19416] = a[13] & g[11224];
assign g[27607] = b[13] & g[11224];
assign g[19417] = a[13] & g[11225];
assign g[27608] = b[13] & g[11225];
assign g[19418] = a[13] & g[11226];
assign g[27609] = b[13] & g[11226];
assign g[19419] = a[13] & g[11227];
assign g[27610] = b[13] & g[11227];
assign g[19420] = a[13] & g[11228];
assign g[27611] = b[13] & g[11228];
assign g[19421] = a[13] & g[11229];
assign g[27612] = b[13] & g[11229];
assign g[19422] = a[13] & g[11230];
assign g[27613] = b[13] & g[11230];
assign g[19423] = a[13] & g[11231];
assign g[27614] = b[13] & g[11231];
assign g[19424] = a[13] & g[11232];
assign g[27615] = b[13] & g[11232];
assign g[19425] = a[13] & g[11233];
assign g[27616] = b[13] & g[11233];
assign g[19426] = a[13] & g[11234];
assign g[27617] = b[13] & g[11234];
assign g[19427] = a[13] & g[11235];
assign g[27618] = b[13] & g[11235];
assign g[19428] = a[13] & g[11236];
assign g[27619] = b[13] & g[11236];
assign g[19429] = a[13] & g[11237];
assign g[27620] = b[13] & g[11237];
assign g[19430] = a[13] & g[11238];
assign g[27621] = b[13] & g[11238];
assign g[19431] = a[13] & g[11239];
assign g[27622] = b[13] & g[11239];
assign g[19432] = a[13] & g[11240];
assign g[27623] = b[13] & g[11240];
assign g[19433] = a[13] & g[11241];
assign g[27624] = b[13] & g[11241];
assign g[19434] = a[13] & g[11242];
assign g[27625] = b[13] & g[11242];
assign g[19435] = a[13] & g[11243];
assign g[27626] = b[13] & g[11243];
assign g[19436] = a[13] & g[11244];
assign g[27627] = b[13] & g[11244];
assign g[19437] = a[13] & g[11245];
assign g[27628] = b[13] & g[11245];
assign g[19438] = a[13] & g[11246];
assign g[27629] = b[13] & g[11246];
assign g[19439] = a[13] & g[11247];
assign g[27630] = b[13] & g[11247];
assign g[19440] = a[13] & g[11248];
assign g[27631] = b[13] & g[11248];
assign g[19441] = a[13] & g[11249];
assign g[27632] = b[13] & g[11249];
assign g[19442] = a[13] & g[11250];
assign g[27633] = b[13] & g[11250];
assign g[19443] = a[13] & g[11251];
assign g[27634] = b[13] & g[11251];
assign g[19444] = a[13] & g[11252];
assign g[27635] = b[13] & g[11252];
assign g[19445] = a[13] & g[11253];
assign g[27636] = b[13] & g[11253];
assign g[19446] = a[13] & g[11254];
assign g[27637] = b[13] & g[11254];
assign g[19447] = a[13] & g[11255];
assign g[27638] = b[13] & g[11255];
assign g[19448] = a[13] & g[11256];
assign g[27639] = b[13] & g[11256];
assign g[19449] = a[13] & g[11257];
assign g[27640] = b[13] & g[11257];
assign g[19450] = a[13] & g[11258];
assign g[27641] = b[13] & g[11258];
assign g[19451] = a[13] & g[11259];
assign g[27642] = b[13] & g[11259];
assign g[19452] = a[13] & g[11260];
assign g[27643] = b[13] & g[11260];
assign g[19453] = a[13] & g[11261];
assign g[27644] = b[13] & g[11261];
assign g[19454] = a[13] & g[11262];
assign g[27645] = b[13] & g[11262];
assign g[19455] = a[13] & g[11263];
assign g[27646] = b[13] & g[11263];
assign g[19456] = a[13] & g[11264];
assign g[27647] = b[13] & g[11264];
assign g[19457] = a[13] & g[11265];
assign g[27648] = b[13] & g[11265];
assign g[19458] = a[13] & g[11266];
assign g[27649] = b[13] & g[11266];
assign g[19459] = a[13] & g[11267];
assign g[27650] = b[13] & g[11267];
assign g[19460] = a[13] & g[11268];
assign g[27651] = b[13] & g[11268];
assign g[19461] = a[13] & g[11269];
assign g[27652] = b[13] & g[11269];
assign g[19462] = a[13] & g[11270];
assign g[27653] = b[13] & g[11270];
assign g[19463] = a[13] & g[11271];
assign g[27654] = b[13] & g[11271];
assign g[19464] = a[13] & g[11272];
assign g[27655] = b[13] & g[11272];
assign g[19465] = a[13] & g[11273];
assign g[27656] = b[13] & g[11273];
assign g[19466] = a[13] & g[11274];
assign g[27657] = b[13] & g[11274];
assign g[19467] = a[13] & g[11275];
assign g[27658] = b[13] & g[11275];
assign g[19468] = a[13] & g[11276];
assign g[27659] = b[13] & g[11276];
assign g[19469] = a[13] & g[11277];
assign g[27660] = b[13] & g[11277];
assign g[19470] = a[13] & g[11278];
assign g[27661] = b[13] & g[11278];
assign g[19471] = a[13] & g[11279];
assign g[27662] = b[13] & g[11279];
assign g[19472] = a[13] & g[11280];
assign g[27663] = b[13] & g[11280];
assign g[19473] = a[13] & g[11281];
assign g[27664] = b[13] & g[11281];
assign g[19474] = a[13] & g[11282];
assign g[27665] = b[13] & g[11282];
assign g[19475] = a[13] & g[11283];
assign g[27666] = b[13] & g[11283];
assign g[19476] = a[13] & g[11284];
assign g[27667] = b[13] & g[11284];
assign g[19477] = a[13] & g[11285];
assign g[27668] = b[13] & g[11285];
assign g[19478] = a[13] & g[11286];
assign g[27669] = b[13] & g[11286];
assign g[19479] = a[13] & g[11287];
assign g[27670] = b[13] & g[11287];
assign g[19480] = a[13] & g[11288];
assign g[27671] = b[13] & g[11288];
assign g[19481] = a[13] & g[11289];
assign g[27672] = b[13] & g[11289];
assign g[19482] = a[13] & g[11290];
assign g[27673] = b[13] & g[11290];
assign g[19483] = a[13] & g[11291];
assign g[27674] = b[13] & g[11291];
assign g[19484] = a[13] & g[11292];
assign g[27675] = b[13] & g[11292];
assign g[19485] = a[13] & g[11293];
assign g[27676] = b[13] & g[11293];
assign g[19486] = a[13] & g[11294];
assign g[27677] = b[13] & g[11294];
assign g[19487] = a[13] & g[11295];
assign g[27678] = b[13] & g[11295];
assign g[19488] = a[13] & g[11296];
assign g[27679] = b[13] & g[11296];
assign g[19489] = a[13] & g[11297];
assign g[27680] = b[13] & g[11297];
assign g[19490] = a[13] & g[11298];
assign g[27681] = b[13] & g[11298];
assign g[19491] = a[13] & g[11299];
assign g[27682] = b[13] & g[11299];
assign g[19492] = a[13] & g[11300];
assign g[27683] = b[13] & g[11300];
assign g[19493] = a[13] & g[11301];
assign g[27684] = b[13] & g[11301];
assign g[19494] = a[13] & g[11302];
assign g[27685] = b[13] & g[11302];
assign g[19495] = a[13] & g[11303];
assign g[27686] = b[13] & g[11303];
assign g[19496] = a[13] & g[11304];
assign g[27687] = b[13] & g[11304];
assign g[19497] = a[13] & g[11305];
assign g[27688] = b[13] & g[11305];
assign g[19498] = a[13] & g[11306];
assign g[27689] = b[13] & g[11306];
assign g[19499] = a[13] & g[11307];
assign g[27690] = b[13] & g[11307];
assign g[19500] = a[13] & g[11308];
assign g[27691] = b[13] & g[11308];
assign g[19501] = a[13] & g[11309];
assign g[27692] = b[13] & g[11309];
assign g[19502] = a[13] & g[11310];
assign g[27693] = b[13] & g[11310];
assign g[19503] = a[13] & g[11311];
assign g[27694] = b[13] & g[11311];
assign g[19504] = a[13] & g[11312];
assign g[27695] = b[13] & g[11312];
assign g[19505] = a[13] & g[11313];
assign g[27696] = b[13] & g[11313];
assign g[19506] = a[13] & g[11314];
assign g[27697] = b[13] & g[11314];
assign g[19507] = a[13] & g[11315];
assign g[27698] = b[13] & g[11315];
assign g[19508] = a[13] & g[11316];
assign g[27699] = b[13] & g[11316];
assign g[19509] = a[13] & g[11317];
assign g[27700] = b[13] & g[11317];
assign g[19510] = a[13] & g[11318];
assign g[27701] = b[13] & g[11318];
assign g[19511] = a[13] & g[11319];
assign g[27702] = b[13] & g[11319];
assign g[19512] = a[13] & g[11320];
assign g[27703] = b[13] & g[11320];
assign g[19513] = a[13] & g[11321];
assign g[27704] = b[13] & g[11321];
assign g[19514] = a[13] & g[11322];
assign g[27705] = b[13] & g[11322];
assign g[19515] = a[13] & g[11323];
assign g[27706] = b[13] & g[11323];
assign g[19516] = a[13] & g[11324];
assign g[27707] = b[13] & g[11324];
assign g[19517] = a[13] & g[11325];
assign g[27708] = b[13] & g[11325];
assign g[19518] = a[13] & g[11326];
assign g[27709] = b[13] & g[11326];
assign g[19519] = a[13] & g[11327];
assign g[27710] = b[13] & g[11327];
assign g[19520] = a[13] & g[11328];
assign g[27711] = b[13] & g[11328];
assign g[19521] = a[13] & g[11329];
assign g[27712] = b[13] & g[11329];
assign g[19522] = a[13] & g[11330];
assign g[27713] = b[13] & g[11330];
assign g[19523] = a[13] & g[11331];
assign g[27714] = b[13] & g[11331];
assign g[19524] = a[13] & g[11332];
assign g[27715] = b[13] & g[11332];
assign g[19525] = a[13] & g[11333];
assign g[27716] = b[13] & g[11333];
assign g[19526] = a[13] & g[11334];
assign g[27717] = b[13] & g[11334];
assign g[19527] = a[13] & g[11335];
assign g[27718] = b[13] & g[11335];
assign g[19528] = a[13] & g[11336];
assign g[27719] = b[13] & g[11336];
assign g[19529] = a[13] & g[11337];
assign g[27720] = b[13] & g[11337];
assign g[19530] = a[13] & g[11338];
assign g[27721] = b[13] & g[11338];
assign g[19531] = a[13] & g[11339];
assign g[27722] = b[13] & g[11339];
assign g[19532] = a[13] & g[11340];
assign g[27723] = b[13] & g[11340];
assign g[19533] = a[13] & g[11341];
assign g[27724] = b[13] & g[11341];
assign g[19534] = a[13] & g[11342];
assign g[27725] = b[13] & g[11342];
assign g[19535] = a[13] & g[11343];
assign g[27726] = b[13] & g[11343];
assign g[19536] = a[13] & g[11344];
assign g[27727] = b[13] & g[11344];
assign g[19537] = a[13] & g[11345];
assign g[27728] = b[13] & g[11345];
assign g[19538] = a[13] & g[11346];
assign g[27729] = b[13] & g[11346];
assign g[19539] = a[13] & g[11347];
assign g[27730] = b[13] & g[11347];
assign g[19540] = a[13] & g[11348];
assign g[27731] = b[13] & g[11348];
assign g[19541] = a[13] & g[11349];
assign g[27732] = b[13] & g[11349];
assign g[19542] = a[13] & g[11350];
assign g[27733] = b[13] & g[11350];
assign g[19543] = a[13] & g[11351];
assign g[27734] = b[13] & g[11351];
assign g[19544] = a[13] & g[11352];
assign g[27735] = b[13] & g[11352];
assign g[19545] = a[13] & g[11353];
assign g[27736] = b[13] & g[11353];
assign g[19546] = a[13] & g[11354];
assign g[27737] = b[13] & g[11354];
assign g[19547] = a[13] & g[11355];
assign g[27738] = b[13] & g[11355];
assign g[19548] = a[13] & g[11356];
assign g[27739] = b[13] & g[11356];
assign g[19549] = a[13] & g[11357];
assign g[27740] = b[13] & g[11357];
assign g[19550] = a[13] & g[11358];
assign g[27741] = b[13] & g[11358];
assign g[19551] = a[13] & g[11359];
assign g[27742] = b[13] & g[11359];
assign g[19552] = a[13] & g[11360];
assign g[27743] = b[13] & g[11360];
assign g[19553] = a[13] & g[11361];
assign g[27744] = b[13] & g[11361];
assign g[19554] = a[13] & g[11362];
assign g[27745] = b[13] & g[11362];
assign g[19555] = a[13] & g[11363];
assign g[27746] = b[13] & g[11363];
assign g[19556] = a[13] & g[11364];
assign g[27747] = b[13] & g[11364];
assign g[19557] = a[13] & g[11365];
assign g[27748] = b[13] & g[11365];
assign g[19558] = a[13] & g[11366];
assign g[27749] = b[13] & g[11366];
assign g[19559] = a[13] & g[11367];
assign g[27750] = b[13] & g[11367];
assign g[19560] = a[13] & g[11368];
assign g[27751] = b[13] & g[11368];
assign g[19561] = a[13] & g[11369];
assign g[27752] = b[13] & g[11369];
assign g[19562] = a[13] & g[11370];
assign g[27753] = b[13] & g[11370];
assign g[19563] = a[13] & g[11371];
assign g[27754] = b[13] & g[11371];
assign g[19564] = a[13] & g[11372];
assign g[27755] = b[13] & g[11372];
assign g[19565] = a[13] & g[11373];
assign g[27756] = b[13] & g[11373];
assign g[19566] = a[13] & g[11374];
assign g[27757] = b[13] & g[11374];
assign g[19567] = a[13] & g[11375];
assign g[27758] = b[13] & g[11375];
assign g[19568] = a[13] & g[11376];
assign g[27759] = b[13] & g[11376];
assign g[19569] = a[13] & g[11377];
assign g[27760] = b[13] & g[11377];
assign g[19570] = a[13] & g[11378];
assign g[27761] = b[13] & g[11378];
assign g[19571] = a[13] & g[11379];
assign g[27762] = b[13] & g[11379];
assign g[19572] = a[13] & g[11380];
assign g[27763] = b[13] & g[11380];
assign g[19573] = a[13] & g[11381];
assign g[27764] = b[13] & g[11381];
assign g[19574] = a[13] & g[11382];
assign g[27765] = b[13] & g[11382];
assign g[19575] = a[13] & g[11383];
assign g[27766] = b[13] & g[11383];
assign g[19576] = a[13] & g[11384];
assign g[27767] = b[13] & g[11384];
assign g[19577] = a[13] & g[11385];
assign g[27768] = b[13] & g[11385];
assign g[19578] = a[13] & g[11386];
assign g[27769] = b[13] & g[11386];
assign g[19579] = a[13] & g[11387];
assign g[27770] = b[13] & g[11387];
assign g[19580] = a[13] & g[11388];
assign g[27771] = b[13] & g[11388];
assign g[19581] = a[13] & g[11389];
assign g[27772] = b[13] & g[11389];
assign g[19582] = a[13] & g[11390];
assign g[27773] = b[13] & g[11390];
assign g[19583] = a[13] & g[11391];
assign g[27774] = b[13] & g[11391];
assign g[19584] = a[13] & g[11392];
assign g[27775] = b[13] & g[11392];
assign g[19585] = a[13] & g[11393];
assign g[27776] = b[13] & g[11393];
assign g[19586] = a[13] & g[11394];
assign g[27777] = b[13] & g[11394];
assign g[19587] = a[13] & g[11395];
assign g[27778] = b[13] & g[11395];
assign g[19588] = a[13] & g[11396];
assign g[27779] = b[13] & g[11396];
assign g[19589] = a[13] & g[11397];
assign g[27780] = b[13] & g[11397];
assign g[19590] = a[13] & g[11398];
assign g[27781] = b[13] & g[11398];
assign g[19591] = a[13] & g[11399];
assign g[27782] = b[13] & g[11399];
assign g[19592] = a[13] & g[11400];
assign g[27783] = b[13] & g[11400];
assign g[19593] = a[13] & g[11401];
assign g[27784] = b[13] & g[11401];
assign g[19594] = a[13] & g[11402];
assign g[27785] = b[13] & g[11402];
assign g[19595] = a[13] & g[11403];
assign g[27786] = b[13] & g[11403];
assign g[19596] = a[13] & g[11404];
assign g[27787] = b[13] & g[11404];
assign g[19597] = a[13] & g[11405];
assign g[27788] = b[13] & g[11405];
assign g[19598] = a[13] & g[11406];
assign g[27789] = b[13] & g[11406];
assign g[19599] = a[13] & g[11407];
assign g[27790] = b[13] & g[11407];
assign g[19600] = a[13] & g[11408];
assign g[27791] = b[13] & g[11408];
assign g[19601] = a[13] & g[11409];
assign g[27792] = b[13] & g[11409];
assign g[19602] = a[13] & g[11410];
assign g[27793] = b[13] & g[11410];
assign g[19603] = a[13] & g[11411];
assign g[27794] = b[13] & g[11411];
assign g[19604] = a[13] & g[11412];
assign g[27795] = b[13] & g[11412];
assign g[19605] = a[13] & g[11413];
assign g[27796] = b[13] & g[11413];
assign g[19606] = a[13] & g[11414];
assign g[27797] = b[13] & g[11414];
assign g[19607] = a[13] & g[11415];
assign g[27798] = b[13] & g[11415];
assign g[19608] = a[13] & g[11416];
assign g[27799] = b[13] & g[11416];
assign g[19609] = a[13] & g[11417];
assign g[27800] = b[13] & g[11417];
assign g[19610] = a[13] & g[11418];
assign g[27801] = b[13] & g[11418];
assign g[19611] = a[13] & g[11419];
assign g[27802] = b[13] & g[11419];
assign g[19612] = a[13] & g[11420];
assign g[27803] = b[13] & g[11420];
assign g[19613] = a[13] & g[11421];
assign g[27804] = b[13] & g[11421];
assign g[19614] = a[13] & g[11422];
assign g[27805] = b[13] & g[11422];
assign g[19615] = a[13] & g[11423];
assign g[27806] = b[13] & g[11423];
assign g[19616] = a[13] & g[11424];
assign g[27807] = b[13] & g[11424];
assign g[19617] = a[13] & g[11425];
assign g[27808] = b[13] & g[11425];
assign g[19618] = a[13] & g[11426];
assign g[27809] = b[13] & g[11426];
assign g[19619] = a[13] & g[11427];
assign g[27810] = b[13] & g[11427];
assign g[19620] = a[13] & g[11428];
assign g[27811] = b[13] & g[11428];
assign g[19621] = a[13] & g[11429];
assign g[27812] = b[13] & g[11429];
assign g[19622] = a[13] & g[11430];
assign g[27813] = b[13] & g[11430];
assign g[19623] = a[13] & g[11431];
assign g[27814] = b[13] & g[11431];
assign g[19624] = a[13] & g[11432];
assign g[27815] = b[13] & g[11432];
assign g[19625] = a[13] & g[11433];
assign g[27816] = b[13] & g[11433];
assign g[19626] = a[13] & g[11434];
assign g[27817] = b[13] & g[11434];
assign g[19627] = a[13] & g[11435];
assign g[27818] = b[13] & g[11435];
assign g[19628] = a[13] & g[11436];
assign g[27819] = b[13] & g[11436];
assign g[19629] = a[13] & g[11437];
assign g[27820] = b[13] & g[11437];
assign g[19630] = a[13] & g[11438];
assign g[27821] = b[13] & g[11438];
assign g[19631] = a[13] & g[11439];
assign g[27822] = b[13] & g[11439];
assign g[19632] = a[13] & g[11440];
assign g[27823] = b[13] & g[11440];
assign g[19633] = a[13] & g[11441];
assign g[27824] = b[13] & g[11441];
assign g[19634] = a[13] & g[11442];
assign g[27825] = b[13] & g[11442];
assign g[19635] = a[13] & g[11443];
assign g[27826] = b[13] & g[11443];
assign g[19636] = a[13] & g[11444];
assign g[27827] = b[13] & g[11444];
assign g[19637] = a[13] & g[11445];
assign g[27828] = b[13] & g[11445];
assign g[19638] = a[13] & g[11446];
assign g[27829] = b[13] & g[11446];
assign g[19639] = a[13] & g[11447];
assign g[27830] = b[13] & g[11447];
assign g[19640] = a[13] & g[11448];
assign g[27831] = b[13] & g[11448];
assign g[19641] = a[13] & g[11449];
assign g[27832] = b[13] & g[11449];
assign g[19642] = a[13] & g[11450];
assign g[27833] = b[13] & g[11450];
assign g[19643] = a[13] & g[11451];
assign g[27834] = b[13] & g[11451];
assign g[19644] = a[13] & g[11452];
assign g[27835] = b[13] & g[11452];
assign g[19645] = a[13] & g[11453];
assign g[27836] = b[13] & g[11453];
assign g[19646] = a[13] & g[11454];
assign g[27837] = b[13] & g[11454];
assign g[19647] = a[13] & g[11455];
assign g[27838] = b[13] & g[11455];
assign g[19648] = a[13] & g[11456];
assign g[27839] = b[13] & g[11456];
assign g[19649] = a[13] & g[11457];
assign g[27840] = b[13] & g[11457];
assign g[19650] = a[13] & g[11458];
assign g[27841] = b[13] & g[11458];
assign g[19651] = a[13] & g[11459];
assign g[27842] = b[13] & g[11459];
assign g[19652] = a[13] & g[11460];
assign g[27843] = b[13] & g[11460];
assign g[19653] = a[13] & g[11461];
assign g[27844] = b[13] & g[11461];
assign g[19654] = a[13] & g[11462];
assign g[27845] = b[13] & g[11462];
assign g[19655] = a[13] & g[11463];
assign g[27846] = b[13] & g[11463];
assign g[19656] = a[13] & g[11464];
assign g[27847] = b[13] & g[11464];
assign g[19657] = a[13] & g[11465];
assign g[27848] = b[13] & g[11465];
assign g[19658] = a[13] & g[11466];
assign g[27849] = b[13] & g[11466];
assign g[19659] = a[13] & g[11467];
assign g[27850] = b[13] & g[11467];
assign g[19660] = a[13] & g[11468];
assign g[27851] = b[13] & g[11468];
assign g[19661] = a[13] & g[11469];
assign g[27852] = b[13] & g[11469];
assign g[19662] = a[13] & g[11470];
assign g[27853] = b[13] & g[11470];
assign g[19663] = a[13] & g[11471];
assign g[27854] = b[13] & g[11471];
assign g[19664] = a[13] & g[11472];
assign g[27855] = b[13] & g[11472];
assign g[19665] = a[13] & g[11473];
assign g[27856] = b[13] & g[11473];
assign g[19666] = a[13] & g[11474];
assign g[27857] = b[13] & g[11474];
assign g[19667] = a[13] & g[11475];
assign g[27858] = b[13] & g[11475];
assign g[19668] = a[13] & g[11476];
assign g[27859] = b[13] & g[11476];
assign g[19669] = a[13] & g[11477];
assign g[27860] = b[13] & g[11477];
assign g[19670] = a[13] & g[11478];
assign g[27861] = b[13] & g[11478];
assign g[19671] = a[13] & g[11479];
assign g[27862] = b[13] & g[11479];
assign g[19672] = a[13] & g[11480];
assign g[27863] = b[13] & g[11480];
assign g[19673] = a[13] & g[11481];
assign g[27864] = b[13] & g[11481];
assign g[19674] = a[13] & g[11482];
assign g[27865] = b[13] & g[11482];
assign g[19675] = a[13] & g[11483];
assign g[27866] = b[13] & g[11483];
assign g[19676] = a[13] & g[11484];
assign g[27867] = b[13] & g[11484];
assign g[19677] = a[13] & g[11485];
assign g[27868] = b[13] & g[11485];
assign g[19678] = a[13] & g[11486];
assign g[27869] = b[13] & g[11486];
assign g[19679] = a[13] & g[11487];
assign g[27870] = b[13] & g[11487];
assign g[19680] = a[13] & g[11488];
assign g[27871] = b[13] & g[11488];
assign g[19681] = a[13] & g[11489];
assign g[27872] = b[13] & g[11489];
assign g[19682] = a[13] & g[11490];
assign g[27873] = b[13] & g[11490];
assign g[19683] = a[13] & g[11491];
assign g[27874] = b[13] & g[11491];
assign g[19684] = a[13] & g[11492];
assign g[27875] = b[13] & g[11492];
assign g[19685] = a[13] & g[11493];
assign g[27876] = b[13] & g[11493];
assign g[19686] = a[13] & g[11494];
assign g[27877] = b[13] & g[11494];
assign g[19687] = a[13] & g[11495];
assign g[27878] = b[13] & g[11495];
assign g[19688] = a[13] & g[11496];
assign g[27879] = b[13] & g[11496];
assign g[19689] = a[13] & g[11497];
assign g[27880] = b[13] & g[11497];
assign g[19690] = a[13] & g[11498];
assign g[27881] = b[13] & g[11498];
assign g[19691] = a[13] & g[11499];
assign g[27882] = b[13] & g[11499];
assign g[19692] = a[13] & g[11500];
assign g[27883] = b[13] & g[11500];
assign g[19693] = a[13] & g[11501];
assign g[27884] = b[13] & g[11501];
assign g[19694] = a[13] & g[11502];
assign g[27885] = b[13] & g[11502];
assign g[19695] = a[13] & g[11503];
assign g[27886] = b[13] & g[11503];
assign g[19696] = a[13] & g[11504];
assign g[27887] = b[13] & g[11504];
assign g[19697] = a[13] & g[11505];
assign g[27888] = b[13] & g[11505];
assign g[19698] = a[13] & g[11506];
assign g[27889] = b[13] & g[11506];
assign g[19699] = a[13] & g[11507];
assign g[27890] = b[13] & g[11507];
assign g[19700] = a[13] & g[11508];
assign g[27891] = b[13] & g[11508];
assign g[19701] = a[13] & g[11509];
assign g[27892] = b[13] & g[11509];
assign g[19702] = a[13] & g[11510];
assign g[27893] = b[13] & g[11510];
assign g[19703] = a[13] & g[11511];
assign g[27894] = b[13] & g[11511];
assign g[19704] = a[13] & g[11512];
assign g[27895] = b[13] & g[11512];
assign g[19705] = a[13] & g[11513];
assign g[27896] = b[13] & g[11513];
assign g[19706] = a[13] & g[11514];
assign g[27897] = b[13] & g[11514];
assign g[19707] = a[13] & g[11515];
assign g[27898] = b[13] & g[11515];
assign g[19708] = a[13] & g[11516];
assign g[27899] = b[13] & g[11516];
assign g[19709] = a[13] & g[11517];
assign g[27900] = b[13] & g[11517];
assign g[19710] = a[13] & g[11518];
assign g[27901] = b[13] & g[11518];
assign g[19711] = a[13] & g[11519];
assign g[27902] = b[13] & g[11519];
assign g[19712] = a[13] & g[11520];
assign g[27903] = b[13] & g[11520];
assign g[19713] = a[13] & g[11521];
assign g[27904] = b[13] & g[11521];
assign g[19714] = a[13] & g[11522];
assign g[27905] = b[13] & g[11522];
assign g[19715] = a[13] & g[11523];
assign g[27906] = b[13] & g[11523];
assign g[19716] = a[13] & g[11524];
assign g[27907] = b[13] & g[11524];
assign g[19717] = a[13] & g[11525];
assign g[27908] = b[13] & g[11525];
assign g[19718] = a[13] & g[11526];
assign g[27909] = b[13] & g[11526];
assign g[19719] = a[13] & g[11527];
assign g[27910] = b[13] & g[11527];
assign g[19720] = a[13] & g[11528];
assign g[27911] = b[13] & g[11528];
assign g[19721] = a[13] & g[11529];
assign g[27912] = b[13] & g[11529];
assign g[19722] = a[13] & g[11530];
assign g[27913] = b[13] & g[11530];
assign g[19723] = a[13] & g[11531];
assign g[27914] = b[13] & g[11531];
assign g[19724] = a[13] & g[11532];
assign g[27915] = b[13] & g[11532];
assign g[19725] = a[13] & g[11533];
assign g[27916] = b[13] & g[11533];
assign g[19726] = a[13] & g[11534];
assign g[27917] = b[13] & g[11534];
assign g[19727] = a[13] & g[11535];
assign g[27918] = b[13] & g[11535];
assign g[19728] = a[13] & g[11536];
assign g[27919] = b[13] & g[11536];
assign g[19729] = a[13] & g[11537];
assign g[27920] = b[13] & g[11537];
assign g[19730] = a[13] & g[11538];
assign g[27921] = b[13] & g[11538];
assign g[19731] = a[13] & g[11539];
assign g[27922] = b[13] & g[11539];
assign g[19732] = a[13] & g[11540];
assign g[27923] = b[13] & g[11540];
assign g[19733] = a[13] & g[11541];
assign g[27924] = b[13] & g[11541];
assign g[19734] = a[13] & g[11542];
assign g[27925] = b[13] & g[11542];
assign g[19735] = a[13] & g[11543];
assign g[27926] = b[13] & g[11543];
assign g[19736] = a[13] & g[11544];
assign g[27927] = b[13] & g[11544];
assign g[19737] = a[13] & g[11545];
assign g[27928] = b[13] & g[11545];
assign g[19738] = a[13] & g[11546];
assign g[27929] = b[13] & g[11546];
assign g[19739] = a[13] & g[11547];
assign g[27930] = b[13] & g[11547];
assign g[19740] = a[13] & g[11548];
assign g[27931] = b[13] & g[11548];
assign g[19741] = a[13] & g[11549];
assign g[27932] = b[13] & g[11549];
assign g[19742] = a[13] & g[11550];
assign g[27933] = b[13] & g[11550];
assign g[19743] = a[13] & g[11551];
assign g[27934] = b[13] & g[11551];
assign g[19744] = a[13] & g[11552];
assign g[27935] = b[13] & g[11552];
assign g[19745] = a[13] & g[11553];
assign g[27936] = b[13] & g[11553];
assign g[19746] = a[13] & g[11554];
assign g[27937] = b[13] & g[11554];
assign g[19747] = a[13] & g[11555];
assign g[27938] = b[13] & g[11555];
assign g[19748] = a[13] & g[11556];
assign g[27939] = b[13] & g[11556];
assign g[19749] = a[13] & g[11557];
assign g[27940] = b[13] & g[11557];
assign g[19750] = a[13] & g[11558];
assign g[27941] = b[13] & g[11558];
assign g[19751] = a[13] & g[11559];
assign g[27942] = b[13] & g[11559];
assign g[19752] = a[13] & g[11560];
assign g[27943] = b[13] & g[11560];
assign g[19753] = a[13] & g[11561];
assign g[27944] = b[13] & g[11561];
assign g[19754] = a[13] & g[11562];
assign g[27945] = b[13] & g[11562];
assign g[19755] = a[13] & g[11563];
assign g[27946] = b[13] & g[11563];
assign g[19756] = a[13] & g[11564];
assign g[27947] = b[13] & g[11564];
assign g[19757] = a[13] & g[11565];
assign g[27948] = b[13] & g[11565];
assign g[19758] = a[13] & g[11566];
assign g[27949] = b[13] & g[11566];
assign g[19759] = a[13] & g[11567];
assign g[27950] = b[13] & g[11567];
assign g[19760] = a[13] & g[11568];
assign g[27951] = b[13] & g[11568];
assign g[19761] = a[13] & g[11569];
assign g[27952] = b[13] & g[11569];
assign g[19762] = a[13] & g[11570];
assign g[27953] = b[13] & g[11570];
assign g[19763] = a[13] & g[11571];
assign g[27954] = b[13] & g[11571];
assign g[19764] = a[13] & g[11572];
assign g[27955] = b[13] & g[11572];
assign g[19765] = a[13] & g[11573];
assign g[27956] = b[13] & g[11573];
assign g[19766] = a[13] & g[11574];
assign g[27957] = b[13] & g[11574];
assign g[19767] = a[13] & g[11575];
assign g[27958] = b[13] & g[11575];
assign g[19768] = a[13] & g[11576];
assign g[27959] = b[13] & g[11576];
assign g[19769] = a[13] & g[11577];
assign g[27960] = b[13] & g[11577];
assign g[19770] = a[13] & g[11578];
assign g[27961] = b[13] & g[11578];
assign g[19771] = a[13] & g[11579];
assign g[27962] = b[13] & g[11579];
assign g[19772] = a[13] & g[11580];
assign g[27963] = b[13] & g[11580];
assign g[19773] = a[13] & g[11581];
assign g[27964] = b[13] & g[11581];
assign g[19774] = a[13] & g[11582];
assign g[27965] = b[13] & g[11582];
assign g[19775] = a[13] & g[11583];
assign g[27966] = b[13] & g[11583];
assign g[19776] = a[13] & g[11584];
assign g[27967] = b[13] & g[11584];
assign g[19777] = a[13] & g[11585];
assign g[27968] = b[13] & g[11585];
assign g[19778] = a[13] & g[11586];
assign g[27969] = b[13] & g[11586];
assign g[19779] = a[13] & g[11587];
assign g[27970] = b[13] & g[11587];
assign g[19780] = a[13] & g[11588];
assign g[27971] = b[13] & g[11588];
assign g[19781] = a[13] & g[11589];
assign g[27972] = b[13] & g[11589];
assign g[19782] = a[13] & g[11590];
assign g[27973] = b[13] & g[11590];
assign g[19783] = a[13] & g[11591];
assign g[27974] = b[13] & g[11591];
assign g[19784] = a[13] & g[11592];
assign g[27975] = b[13] & g[11592];
assign g[19785] = a[13] & g[11593];
assign g[27976] = b[13] & g[11593];
assign g[19786] = a[13] & g[11594];
assign g[27977] = b[13] & g[11594];
assign g[19787] = a[13] & g[11595];
assign g[27978] = b[13] & g[11595];
assign g[19788] = a[13] & g[11596];
assign g[27979] = b[13] & g[11596];
assign g[19789] = a[13] & g[11597];
assign g[27980] = b[13] & g[11597];
assign g[19790] = a[13] & g[11598];
assign g[27981] = b[13] & g[11598];
assign g[19791] = a[13] & g[11599];
assign g[27982] = b[13] & g[11599];
assign g[19792] = a[13] & g[11600];
assign g[27983] = b[13] & g[11600];
assign g[19793] = a[13] & g[11601];
assign g[27984] = b[13] & g[11601];
assign g[19794] = a[13] & g[11602];
assign g[27985] = b[13] & g[11602];
assign g[19795] = a[13] & g[11603];
assign g[27986] = b[13] & g[11603];
assign g[19796] = a[13] & g[11604];
assign g[27987] = b[13] & g[11604];
assign g[19797] = a[13] & g[11605];
assign g[27988] = b[13] & g[11605];
assign g[19798] = a[13] & g[11606];
assign g[27989] = b[13] & g[11606];
assign g[19799] = a[13] & g[11607];
assign g[27990] = b[13] & g[11607];
assign g[19800] = a[13] & g[11608];
assign g[27991] = b[13] & g[11608];
assign g[19801] = a[13] & g[11609];
assign g[27992] = b[13] & g[11609];
assign g[19802] = a[13] & g[11610];
assign g[27993] = b[13] & g[11610];
assign g[19803] = a[13] & g[11611];
assign g[27994] = b[13] & g[11611];
assign g[19804] = a[13] & g[11612];
assign g[27995] = b[13] & g[11612];
assign g[19805] = a[13] & g[11613];
assign g[27996] = b[13] & g[11613];
assign g[19806] = a[13] & g[11614];
assign g[27997] = b[13] & g[11614];
assign g[19807] = a[13] & g[11615];
assign g[27998] = b[13] & g[11615];
assign g[19808] = a[13] & g[11616];
assign g[27999] = b[13] & g[11616];
assign g[19809] = a[13] & g[11617];
assign g[28000] = b[13] & g[11617];
assign g[19810] = a[13] & g[11618];
assign g[28001] = b[13] & g[11618];
assign g[19811] = a[13] & g[11619];
assign g[28002] = b[13] & g[11619];
assign g[19812] = a[13] & g[11620];
assign g[28003] = b[13] & g[11620];
assign g[19813] = a[13] & g[11621];
assign g[28004] = b[13] & g[11621];
assign g[19814] = a[13] & g[11622];
assign g[28005] = b[13] & g[11622];
assign g[19815] = a[13] & g[11623];
assign g[28006] = b[13] & g[11623];
assign g[19816] = a[13] & g[11624];
assign g[28007] = b[13] & g[11624];
assign g[19817] = a[13] & g[11625];
assign g[28008] = b[13] & g[11625];
assign g[19818] = a[13] & g[11626];
assign g[28009] = b[13] & g[11626];
assign g[19819] = a[13] & g[11627];
assign g[28010] = b[13] & g[11627];
assign g[19820] = a[13] & g[11628];
assign g[28011] = b[13] & g[11628];
assign g[19821] = a[13] & g[11629];
assign g[28012] = b[13] & g[11629];
assign g[19822] = a[13] & g[11630];
assign g[28013] = b[13] & g[11630];
assign g[19823] = a[13] & g[11631];
assign g[28014] = b[13] & g[11631];
assign g[19824] = a[13] & g[11632];
assign g[28015] = b[13] & g[11632];
assign g[19825] = a[13] & g[11633];
assign g[28016] = b[13] & g[11633];
assign g[19826] = a[13] & g[11634];
assign g[28017] = b[13] & g[11634];
assign g[19827] = a[13] & g[11635];
assign g[28018] = b[13] & g[11635];
assign g[19828] = a[13] & g[11636];
assign g[28019] = b[13] & g[11636];
assign g[19829] = a[13] & g[11637];
assign g[28020] = b[13] & g[11637];
assign g[19830] = a[13] & g[11638];
assign g[28021] = b[13] & g[11638];
assign g[19831] = a[13] & g[11639];
assign g[28022] = b[13] & g[11639];
assign g[19832] = a[13] & g[11640];
assign g[28023] = b[13] & g[11640];
assign g[19833] = a[13] & g[11641];
assign g[28024] = b[13] & g[11641];
assign g[19834] = a[13] & g[11642];
assign g[28025] = b[13] & g[11642];
assign g[19835] = a[13] & g[11643];
assign g[28026] = b[13] & g[11643];
assign g[19836] = a[13] & g[11644];
assign g[28027] = b[13] & g[11644];
assign g[19837] = a[13] & g[11645];
assign g[28028] = b[13] & g[11645];
assign g[19838] = a[13] & g[11646];
assign g[28029] = b[13] & g[11646];
assign g[19839] = a[13] & g[11647];
assign g[28030] = b[13] & g[11647];
assign g[19840] = a[13] & g[11648];
assign g[28031] = b[13] & g[11648];
assign g[19841] = a[13] & g[11649];
assign g[28032] = b[13] & g[11649];
assign g[19842] = a[13] & g[11650];
assign g[28033] = b[13] & g[11650];
assign g[19843] = a[13] & g[11651];
assign g[28034] = b[13] & g[11651];
assign g[19844] = a[13] & g[11652];
assign g[28035] = b[13] & g[11652];
assign g[19845] = a[13] & g[11653];
assign g[28036] = b[13] & g[11653];
assign g[19846] = a[13] & g[11654];
assign g[28037] = b[13] & g[11654];
assign g[19847] = a[13] & g[11655];
assign g[28038] = b[13] & g[11655];
assign g[19848] = a[13] & g[11656];
assign g[28039] = b[13] & g[11656];
assign g[19849] = a[13] & g[11657];
assign g[28040] = b[13] & g[11657];
assign g[19850] = a[13] & g[11658];
assign g[28041] = b[13] & g[11658];
assign g[19851] = a[13] & g[11659];
assign g[28042] = b[13] & g[11659];
assign g[19852] = a[13] & g[11660];
assign g[28043] = b[13] & g[11660];
assign g[19853] = a[13] & g[11661];
assign g[28044] = b[13] & g[11661];
assign g[19854] = a[13] & g[11662];
assign g[28045] = b[13] & g[11662];
assign g[19855] = a[13] & g[11663];
assign g[28046] = b[13] & g[11663];
assign g[19856] = a[13] & g[11664];
assign g[28047] = b[13] & g[11664];
assign g[19857] = a[13] & g[11665];
assign g[28048] = b[13] & g[11665];
assign g[19858] = a[13] & g[11666];
assign g[28049] = b[13] & g[11666];
assign g[19859] = a[13] & g[11667];
assign g[28050] = b[13] & g[11667];
assign g[19860] = a[13] & g[11668];
assign g[28051] = b[13] & g[11668];
assign g[19861] = a[13] & g[11669];
assign g[28052] = b[13] & g[11669];
assign g[19862] = a[13] & g[11670];
assign g[28053] = b[13] & g[11670];
assign g[19863] = a[13] & g[11671];
assign g[28054] = b[13] & g[11671];
assign g[19864] = a[13] & g[11672];
assign g[28055] = b[13] & g[11672];
assign g[19865] = a[13] & g[11673];
assign g[28056] = b[13] & g[11673];
assign g[19866] = a[13] & g[11674];
assign g[28057] = b[13] & g[11674];
assign g[19867] = a[13] & g[11675];
assign g[28058] = b[13] & g[11675];
assign g[19868] = a[13] & g[11676];
assign g[28059] = b[13] & g[11676];
assign g[19869] = a[13] & g[11677];
assign g[28060] = b[13] & g[11677];
assign g[19870] = a[13] & g[11678];
assign g[28061] = b[13] & g[11678];
assign g[19871] = a[13] & g[11679];
assign g[28062] = b[13] & g[11679];
assign g[19872] = a[13] & g[11680];
assign g[28063] = b[13] & g[11680];
assign g[19873] = a[13] & g[11681];
assign g[28064] = b[13] & g[11681];
assign g[19874] = a[13] & g[11682];
assign g[28065] = b[13] & g[11682];
assign g[19875] = a[13] & g[11683];
assign g[28066] = b[13] & g[11683];
assign g[19876] = a[13] & g[11684];
assign g[28067] = b[13] & g[11684];
assign g[19877] = a[13] & g[11685];
assign g[28068] = b[13] & g[11685];
assign g[19878] = a[13] & g[11686];
assign g[28069] = b[13] & g[11686];
assign g[19879] = a[13] & g[11687];
assign g[28070] = b[13] & g[11687];
assign g[19880] = a[13] & g[11688];
assign g[28071] = b[13] & g[11688];
assign g[19881] = a[13] & g[11689];
assign g[28072] = b[13] & g[11689];
assign g[19882] = a[13] & g[11690];
assign g[28073] = b[13] & g[11690];
assign g[19883] = a[13] & g[11691];
assign g[28074] = b[13] & g[11691];
assign g[19884] = a[13] & g[11692];
assign g[28075] = b[13] & g[11692];
assign g[19885] = a[13] & g[11693];
assign g[28076] = b[13] & g[11693];
assign g[19886] = a[13] & g[11694];
assign g[28077] = b[13] & g[11694];
assign g[19887] = a[13] & g[11695];
assign g[28078] = b[13] & g[11695];
assign g[19888] = a[13] & g[11696];
assign g[28079] = b[13] & g[11696];
assign g[19889] = a[13] & g[11697];
assign g[28080] = b[13] & g[11697];
assign g[19890] = a[13] & g[11698];
assign g[28081] = b[13] & g[11698];
assign g[19891] = a[13] & g[11699];
assign g[28082] = b[13] & g[11699];
assign g[19892] = a[13] & g[11700];
assign g[28083] = b[13] & g[11700];
assign g[19893] = a[13] & g[11701];
assign g[28084] = b[13] & g[11701];
assign g[19894] = a[13] & g[11702];
assign g[28085] = b[13] & g[11702];
assign g[19895] = a[13] & g[11703];
assign g[28086] = b[13] & g[11703];
assign g[19896] = a[13] & g[11704];
assign g[28087] = b[13] & g[11704];
assign g[19897] = a[13] & g[11705];
assign g[28088] = b[13] & g[11705];
assign g[19898] = a[13] & g[11706];
assign g[28089] = b[13] & g[11706];
assign g[19899] = a[13] & g[11707];
assign g[28090] = b[13] & g[11707];
assign g[19900] = a[13] & g[11708];
assign g[28091] = b[13] & g[11708];
assign g[19901] = a[13] & g[11709];
assign g[28092] = b[13] & g[11709];
assign g[19902] = a[13] & g[11710];
assign g[28093] = b[13] & g[11710];
assign g[19903] = a[13] & g[11711];
assign g[28094] = b[13] & g[11711];
assign g[19904] = a[13] & g[11712];
assign g[28095] = b[13] & g[11712];
assign g[19905] = a[13] & g[11713];
assign g[28096] = b[13] & g[11713];
assign g[19906] = a[13] & g[11714];
assign g[28097] = b[13] & g[11714];
assign g[19907] = a[13] & g[11715];
assign g[28098] = b[13] & g[11715];
assign g[19908] = a[13] & g[11716];
assign g[28099] = b[13] & g[11716];
assign g[19909] = a[13] & g[11717];
assign g[28100] = b[13] & g[11717];
assign g[19910] = a[13] & g[11718];
assign g[28101] = b[13] & g[11718];
assign g[19911] = a[13] & g[11719];
assign g[28102] = b[13] & g[11719];
assign g[19912] = a[13] & g[11720];
assign g[28103] = b[13] & g[11720];
assign g[19913] = a[13] & g[11721];
assign g[28104] = b[13] & g[11721];
assign g[19914] = a[13] & g[11722];
assign g[28105] = b[13] & g[11722];
assign g[19915] = a[13] & g[11723];
assign g[28106] = b[13] & g[11723];
assign g[19916] = a[13] & g[11724];
assign g[28107] = b[13] & g[11724];
assign g[19917] = a[13] & g[11725];
assign g[28108] = b[13] & g[11725];
assign g[19918] = a[13] & g[11726];
assign g[28109] = b[13] & g[11726];
assign g[19919] = a[13] & g[11727];
assign g[28110] = b[13] & g[11727];
assign g[19920] = a[13] & g[11728];
assign g[28111] = b[13] & g[11728];
assign g[19921] = a[13] & g[11729];
assign g[28112] = b[13] & g[11729];
assign g[19922] = a[13] & g[11730];
assign g[28113] = b[13] & g[11730];
assign g[19923] = a[13] & g[11731];
assign g[28114] = b[13] & g[11731];
assign g[19924] = a[13] & g[11732];
assign g[28115] = b[13] & g[11732];
assign g[19925] = a[13] & g[11733];
assign g[28116] = b[13] & g[11733];
assign g[19926] = a[13] & g[11734];
assign g[28117] = b[13] & g[11734];
assign g[19927] = a[13] & g[11735];
assign g[28118] = b[13] & g[11735];
assign g[19928] = a[13] & g[11736];
assign g[28119] = b[13] & g[11736];
assign g[19929] = a[13] & g[11737];
assign g[28120] = b[13] & g[11737];
assign g[19930] = a[13] & g[11738];
assign g[28121] = b[13] & g[11738];
assign g[19931] = a[13] & g[11739];
assign g[28122] = b[13] & g[11739];
assign g[19932] = a[13] & g[11740];
assign g[28123] = b[13] & g[11740];
assign g[19933] = a[13] & g[11741];
assign g[28124] = b[13] & g[11741];
assign g[19934] = a[13] & g[11742];
assign g[28125] = b[13] & g[11742];
assign g[19935] = a[13] & g[11743];
assign g[28126] = b[13] & g[11743];
assign g[19936] = a[13] & g[11744];
assign g[28127] = b[13] & g[11744];
assign g[19937] = a[13] & g[11745];
assign g[28128] = b[13] & g[11745];
assign g[19938] = a[13] & g[11746];
assign g[28129] = b[13] & g[11746];
assign g[19939] = a[13] & g[11747];
assign g[28130] = b[13] & g[11747];
assign g[19940] = a[13] & g[11748];
assign g[28131] = b[13] & g[11748];
assign g[19941] = a[13] & g[11749];
assign g[28132] = b[13] & g[11749];
assign g[19942] = a[13] & g[11750];
assign g[28133] = b[13] & g[11750];
assign g[19943] = a[13] & g[11751];
assign g[28134] = b[13] & g[11751];
assign g[19944] = a[13] & g[11752];
assign g[28135] = b[13] & g[11752];
assign g[19945] = a[13] & g[11753];
assign g[28136] = b[13] & g[11753];
assign g[19946] = a[13] & g[11754];
assign g[28137] = b[13] & g[11754];
assign g[19947] = a[13] & g[11755];
assign g[28138] = b[13] & g[11755];
assign g[19948] = a[13] & g[11756];
assign g[28139] = b[13] & g[11756];
assign g[19949] = a[13] & g[11757];
assign g[28140] = b[13] & g[11757];
assign g[19950] = a[13] & g[11758];
assign g[28141] = b[13] & g[11758];
assign g[19951] = a[13] & g[11759];
assign g[28142] = b[13] & g[11759];
assign g[19952] = a[13] & g[11760];
assign g[28143] = b[13] & g[11760];
assign g[19953] = a[13] & g[11761];
assign g[28144] = b[13] & g[11761];
assign g[19954] = a[13] & g[11762];
assign g[28145] = b[13] & g[11762];
assign g[19955] = a[13] & g[11763];
assign g[28146] = b[13] & g[11763];
assign g[19956] = a[13] & g[11764];
assign g[28147] = b[13] & g[11764];
assign g[19957] = a[13] & g[11765];
assign g[28148] = b[13] & g[11765];
assign g[19958] = a[13] & g[11766];
assign g[28149] = b[13] & g[11766];
assign g[19959] = a[13] & g[11767];
assign g[28150] = b[13] & g[11767];
assign g[19960] = a[13] & g[11768];
assign g[28151] = b[13] & g[11768];
assign g[19961] = a[13] & g[11769];
assign g[28152] = b[13] & g[11769];
assign g[19962] = a[13] & g[11770];
assign g[28153] = b[13] & g[11770];
assign g[19963] = a[13] & g[11771];
assign g[28154] = b[13] & g[11771];
assign g[19964] = a[13] & g[11772];
assign g[28155] = b[13] & g[11772];
assign g[19965] = a[13] & g[11773];
assign g[28156] = b[13] & g[11773];
assign g[19966] = a[13] & g[11774];
assign g[28157] = b[13] & g[11774];
assign g[19967] = a[13] & g[11775];
assign g[28158] = b[13] & g[11775];
assign g[19968] = a[13] & g[11776];
assign g[28159] = b[13] & g[11776];
assign g[19969] = a[13] & g[11777];
assign g[28160] = b[13] & g[11777];
assign g[19970] = a[13] & g[11778];
assign g[28161] = b[13] & g[11778];
assign g[19971] = a[13] & g[11779];
assign g[28162] = b[13] & g[11779];
assign g[19972] = a[13] & g[11780];
assign g[28163] = b[13] & g[11780];
assign g[19973] = a[13] & g[11781];
assign g[28164] = b[13] & g[11781];
assign g[19974] = a[13] & g[11782];
assign g[28165] = b[13] & g[11782];
assign g[19975] = a[13] & g[11783];
assign g[28166] = b[13] & g[11783];
assign g[19976] = a[13] & g[11784];
assign g[28167] = b[13] & g[11784];
assign g[19977] = a[13] & g[11785];
assign g[28168] = b[13] & g[11785];
assign g[19978] = a[13] & g[11786];
assign g[28169] = b[13] & g[11786];
assign g[19979] = a[13] & g[11787];
assign g[28170] = b[13] & g[11787];
assign g[19980] = a[13] & g[11788];
assign g[28171] = b[13] & g[11788];
assign g[19981] = a[13] & g[11789];
assign g[28172] = b[13] & g[11789];
assign g[19982] = a[13] & g[11790];
assign g[28173] = b[13] & g[11790];
assign g[19983] = a[13] & g[11791];
assign g[28174] = b[13] & g[11791];
assign g[19984] = a[13] & g[11792];
assign g[28175] = b[13] & g[11792];
assign g[19985] = a[13] & g[11793];
assign g[28176] = b[13] & g[11793];
assign g[19986] = a[13] & g[11794];
assign g[28177] = b[13] & g[11794];
assign g[19987] = a[13] & g[11795];
assign g[28178] = b[13] & g[11795];
assign g[19988] = a[13] & g[11796];
assign g[28179] = b[13] & g[11796];
assign g[19989] = a[13] & g[11797];
assign g[28180] = b[13] & g[11797];
assign g[19990] = a[13] & g[11798];
assign g[28181] = b[13] & g[11798];
assign g[19991] = a[13] & g[11799];
assign g[28182] = b[13] & g[11799];
assign g[19992] = a[13] & g[11800];
assign g[28183] = b[13] & g[11800];
assign g[19993] = a[13] & g[11801];
assign g[28184] = b[13] & g[11801];
assign g[19994] = a[13] & g[11802];
assign g[28185] = b[13] & g[11802];
assign g[19995] = a[13] & g[11803];
assign g[28186] = b[13] & g[11803];
assign g[19996] = a[13] & g[11804];
assign g[28187] = b[13] & g[11804];
assign g[19997] = a[13] & g[11805];
assign g[28188] = b[13] & g[11805];
assign g[19998] = a[13] & g[11806];
assign g[28189] = b[13] & g[11806];
assign g[19999] = a[13] & g[11807];
assign g[28190] = b[13] & g[11807];
assign g[20000] = a[13] & g[11808];
assign g[28191] = b[13] & g[11808];
assign g[20001] = a[13] & g[11809];
assign g[28192] = b[13] & g[11809];
assign g[20002] = a[13] & g[11810];
assign g[28193] = b[13] & g[11810];
assign g[20003] = a[13] & g[11811];
assign g[28194] = b[13] & g[11811];
assign g[20004] = a[13] & g[11812];
assign g[28195] = b[13] & g[11812];
assign g[20005] = a[13] & g[11813];
assign g[28196] = b[13] & g[11813];
assign g[20006] = a[13] & g[11814];
assign g[28197] = b[13] & g[11814];
assign g[20007] = a[13] & g[11815];
assign g[28198] = b[13] & g[11815];
assign g[20008] = a[13] & g[11816];
assign g[28199] = b[13] & g[11816];
assign g[20009] = a[13] & g[11817];
assign g[28200] = b[13] & g[11817];
assign g[20010] = a[13] & g[11818];
assign g[28201] = b[13] & g[11818];
assign g[20011] = a[13] & g[11819];
assign g[28202] = b[13] & g[11819];
assign g[20012] = a[13] & g[11820];
assign g[28203] = b[13] & g[11820];
assign g[20013] = a[13] & g[11821];
assign g[28204] = b[13] & g[11821];
assign g[20014] = a[13] & g[11822];
assign g[28205] = b[13] & g[11822];
assign g[20015] = a[13] & g[11823];
assign g[28206] = b[13] & g[11823];
assign g[20016] = a[13] & g[11824];
assign g[28207] = b[13] & g[11824];
assign g[20017] = a[13] & g[11825];
assign g[28208] = b[13] & g[11825];
assign g[20018] = a[13] & g[11826];
assign g[28209] = b[13] & g[11826];
assign g[20019] = a[13] & g[11827];
assign g[28210] = b[13] & g[11827];
assign g[20020] = a[13] & g[11828];
assign g[28211] = b[13] & g[11828];
assign g[20021] = a[13] & g[11829];
assign g[28212] = b[13] & g[11829];
assign g[20022] = a[13] & g[11830];
assign g[28213] = b[13] & g[11830];
assign g[20023] = a[13] & g[11831];
assign g[28214] = b[13] & g[11831];
assign g[20024] = a[13] & g[11832];
assign g[28215] = b[13] & g[11832];
assign g[20025] = a[13] & g[11833];
assign g[28216] = b[13] & g[11833];
assign g[20026] = a[13] & g[11834];
assign g[28217] = b[13] & g[11834];
assign g[20027] = a[13] & g[11835];
assign g[28218] = b[13] & g[11835];
assign g[20028] = a[13] & g[11836];
assign g[28219] = b[13] & g[11836];
assign g[20029] = a[13] & g[11837];
assign g[28220] = b[13] & g[11837];
assign g[20030] = a[13] & g[11838];
assign g[28221] = b[13] & g[11838];
assign g[20031] = a[13] & g[11839];
assign g[28222] = b[13] & g[11839];
assign g[20032] = a[13] & g[11840];
assign g[28223] = b[13] & g[11840];
assign g[20033] = a[13] & g[11841];
assign g[28224] = b[13] & g[11841];
assign g[20034] = a[13] & g[11842];
assign g[28225] = b[13] & g[11842];
assign g[20035] = a[13] & g[11843];
assign g[28226] = b[13] & g[11843];
assign g[20036] = a[13] & g[11844];
assign g[28227] = b[13] & g[11844];
assign g[20037] = a[13] & g[11845];
assign g[28228] = b[13] & g[11845];
assign g[20038] = a[13] & g[11846];
assign g[28229] = b[13] & g[11846];
assign g[20039] = a[13] & g[11847];
assign g[28230] = b[13] & g[11847];
assign g[20040] = a[13] & g[11848];
assign g[28231] = b[13] & g[11848];
assign g[20041] = a[13] & g[11849];
assign g[28232] = b[13] & g[11849];
assign g[20042] = a[13] & g[11850];
assign g[28233] = b[13] & g[11850];
assign g[20043] = a[13] & g[11851];
assign g[28234] = b[13] & g[11851];
assign g[20044] = a[13] & g[11852];
assign g[28235] = b[13] & g[11852];
assign g[20045] = a[13] & g[11853];
assign g[28236] = b[13] & g[11853];
assign g[20046] = a[13] & g[11854];
assign g[28237] = b[13] & g[11854];
assign g[20047] = a[13] & g[11855];
assign g[28238] = b[13] & g[11855];
assign g[20048] = a[13] & g[11856];
assign g[28239] = b[13] & g[11856];
assign g[20049] = a[13] & g[11857];
assign g[28240] = b[13] & g[11857];
assign g[20050] = a[13] & g[11858];
assign g[28241] = b[13] & g[11858];
assign g[20051] = a[13] & g[11859];
assign g[28242] = b[13] & g[11859];
assign g[20052] = a[13] & g[11860];
assign g[28243] = b[13] & g[11860];
assign g[20053] = a[13] & g[11861];
assign g[28244] = b[13] & g[11861];
assign g[20054] = a[13] & g[11862];
assign g[28245] = b[13] & g[11862];
assign g[20055] = a[13] & g[11863];
assign g[28246] = b[13] & g[11863];
assign g[20056] = a[13] & g[11864];
assign g[28247] = b[13] & g[11864];
assign g[20057] = a[13] & g[11865];
assign g[28248] = b[13] & g[11865];
assign g[20058] = a[13] & g[11866];
assign g[28249] = b[13] & g[11866];
assign g[20059] = a[13] & g[11867];
assign g[28250] = b[13] & g[11867];
assign g[20060] = a[13] & g[11868];
assign g[28251] = b[13] & g[11868];
assign g[20061] = a[13] & g[11869];
assign g[28252] = b[13] & g[11869];
assign g[20062] = a[13] & g[11870];
assign g[28253] = b[13] & g[11870];
assign g[20063] = a[13] & g[11871];
assign g[28254] = b[13] & g[11871];
assign g[20064] = a[13] & g[11872];
assign g[28255] = b[13] & g[11872];
assign g[20065] = a[13] & g[11873];
assign g[28256] = b[13] & g[11873];
assign g[20066] = a[13] & g[11874];
assign g[28257] = b[13] & g[11874];
assign g[20067] = a[13] & g[11875];
assign g[28258] = b[13] & g[11875];
assign g[20068] = a[13] & g[11876];
assign g[28259] = b[13] & g[11876];
assign g[20069] = a[13] & g[11877];
assign g[28260] = b[13] & g[11877];
assign g[20070] = a[13] & g[11878];
assign g[28261] = b[13] & g[11878];
assign g[20071] = a[13] & g[11879];
assign g[28262] = b[13] & g[11879];
assign g[20072] = a[13] & g[11880];
assign g[28263] = b[13] & g[11880];
assign g[20073] = a[13] & g[11881];
assign g[28264] = b[13] & g[11881];
assign g[20074] = a[13] & g[11882];
assign g[28265] = b[13] & g[11882];
assign g[20075] = a[13] & g[11883];
assign g[28266] = b[13] & g[11883];
assign g[20076] = a[13] & g[11884];
assign g[28267] = b[13] & g[11884];
assign g[20077] = a[13] & g[11885];
assign g[28268] = b[13] & g[11885];
assign g[20078] = a[13] & g[11886];
assign g[28269] = b[13] & g[11886];
assign g[20079] = a[13] & g[11887];
assign g[28270] = b[13] & g[11887];
assign g[20080] = a[13] & g[11888];
assign g[28271] = b[13] & g[11888];
assign g[20081] = a[13] & g[11889];
assign g[28272] = b[13] & g[11889];
assign g[20082] = a[13] & g[11890];
assign g[28273] = b[13] & g[11890];
assign g[20083] = a[13] & g[11891];
assign g[28274] = b[13] & g[11891];
assign g[20084] = a[13] & g[11892];
assign g[28275] = b[13] & g[11892];
assign g[20085] = a[13] & g[11893];
assign g[28276] = b[13] & g[11893];
assign g[20086] = a[13] & g[11894];
assign g[28277] = b[13] & g[11894];
assign g[20087] = a[13] & g[11895];
assign g[28278] = b[13] & g[11895];
assign g[20088] = a[13] & g[11896];
assign g[28279] = b[13] & g[11896];
assign g[20089] = a[13] & g[11897];
assign g[28280] = b[13] & g[11897];
assign g[20090] = a[13] & g[11898];
assign g[28281] = b[13] & g[11898];
assign g[20091] = a[13] & g[11899];
assign g[28282] = b[13] & g[11899];
assign g[20092] = a[13] & g[11900];
assign g[28283] = b[13] & g[11900];
assign g[20093] = a[13] & g[11901];
assign g[28284] = b[13] & g[11901];
assign g[20094] = a[13] & g[11902];
assign g[28285] = b[13] & g[11902];
assign g[20095] = a[13] & g[11903];
assign g[28286] = b[13] & g[11903];
assign g[20096] = a[13] & g[11904];
assign g[28287] = b[13] & g[11904];
assign g[20097] = a[13] & g[11905];
assign g[28288] = b[13] & g[11905];
assign g[20098] = a[13] & g[11906];
assign g[28289] = b[13] & g[11906];
assign g[20099] = a[13] & g[11907];
assign g[28290] = b[13] & g[11907];
assign g[20100] = a[13] & g[11908];
assign g[28291] = b[13] & g[11908];
assign g[20101] = a[13] & g[11909];
assign g[28292] = b[13] & g[11909];
assign g[20102] = a[13] & g[11910];
assign g[28293] = b[13] & g[11910];
assign g[20103] = a[13] & g[11911];
assign g[28294] = b[13] & g[11911];
assign g[20104] = a[13] & g[11912];
assign g[28295] = b[13] & g[11912];
assign g[20105] = a[13] & g[11913];
assign g[28296] = b[13] & g[11913];
assign g[20106] = a[13] & g[11914];
assign g[28297] = b[13] & g[11914];
assign g[20107] = a[13] & g[11915];
assign g[28298] = b[13] & g[11915];
assign g[20108] = a[13] & g[11916];
assign g[28299] = b[13] & g[11916];
assign g[20109] = a[13] & g[11917];
assign g[28300] = b[13] & g[11917];
assign g[20110] = a[13] & g[11918];
assign g[28301] = b[13] & g[11918];
assign g[20111] = a[13] & g[11919];
assign g[28302] = b[13] & g[11919];
assign g[20112] = a[13] & g[11920];
assign g[28303] = b[13] & g[11920];
assign g[20113] = a[13] & g[11921];
assign g[28304] = b[13] & g[11921];
assign g[20114] = a[13] & g[11922];
assign g[28305] = b[13] & g[11922];
assign g[20115] = a[13] & g[11923];
assign g[28306] = b[13] & g[11923];
assign g[20116] = a[13] & g[11924];
assign g[28307] = b[13] & g[11924];
assign g[20117] = a[13] & g[11925];
assign g[28308] = b[13] & g[11925];
assign g[20118] = a[13] & g[11926];
assign g[28309] = b[13] & g[11926];
assign g[20119] = a[13] & g[11927];
assign g[28310] = b[13] & g[11927];
assign g[20120] = a[13] & g[11928];
assign g[28311] = b[13] & g[11928];
assign g[20121] = a[13] & g[11929];
assign g[28312] = b[13] & g[11929];
assign g[20122] = a[13] & g[11930];
assign g[28313] = b[13] & g[11930];
assign g[20123] = a[13] & g[11931];
assign g[28314] = b[13] & g[11931];
assign g[20124] = a[13] & g[11932];
assign g[28315] = b[13] & g[11932];
assign g[20125] = a[13] & g[11933];
assign g[28316] = b[13] & g[11933];
assign g[20126] = a[13] & g[11934];
assign g[28317] = b[13] & g[11934];
assign g[20127] = a[13] & g[11935];
assign g[28318] = b[13] & g[11935];
assign g[20128] = a[13] & g[11936];
assign g[28319] = b[13] & g[11936];
assign g[20129] = a[13] & g[11937];
assign g[28320] = b[13] & g[11937];
assign g[20130] = a[13] & g[11938];
assign g[28321] = b[13] & g[11938];
assign g[20131] = a[13] & g[11939];
assign g[28322] = b[13] & g[11939];
assign g[20132] = a[13] & g[11940];
assign g[28323] = b[13] & g[11940];
assign g[20133] = a[13] & g[11941];
assign g[28324] = b[13] & g[11941];
assign g[20134] = a[13] & g[11942];
assign g[28325] = b[13] & g[11942];
assign g[20135] = a[13] & g[11943];
assign g[28326] = b[13] & g[11943];
assign g[20136] = a[13] & g[11944];
assign g[28327] = b[13] & g[11944];
assign g[20137] = a[13] & g[11945];
assign g[28328] = b[13] & g[11945];
assign g[20138] = a[13] & g[11946];
assign g[28329] = b[13] & g[11946];
assign g[20139] = a[13] & g[11947];
assign g[28330] = b[13] & g[11947];
assign g[20140] = a[13] & g[11948];
assign g[28331] = b[13] & g[11948];
assign g[20141] = a[13] & g[11949];
assign g[28332] = b[13] & g[11949];
assign g[20142] = a[13] & g[11950];
assign g[28333] = b[13] & g[11950];
assign g[20143] = a[13] & g[11951];
assign g[28334] = b[13] & g[11951];
assign g[20144] = a[13] & g[11952];
assign g[28335] = b[13] & g[11952];
assign g[20145] = a[13] & g[11953];
assign g[28336] = b[13] & g[11953];
assign g[20146] = a[13] & g[11954];
assign g[28337] = b[13] & g[11954];
assign g[20147] = a[13] & g[11955];
assign g[28338] = b[13] & g[11955];
assign g[20148] = a[13] & g[11956];
assign g[28339] = b[13] & g[11956];
assign g[20149] = a[13] & g[11957];
assign g[28340] = b[13] & g[11957];
assign g[20150] = a[13] & g[11958];
assign g[28341] = b[13] & g[11958];
assign g[20151] = a[13] & g[11959];
assign g[28342] = b[13] & g[11959];
assign g[20152] = a[13] & g[11960];
assign g[28343] = b[13] & g[11960];
assign g[20153] = a[13] & g[11961];
assign g[28344] = b[13] & g[11961];
assign g[20154] = a[13] & g[11962];
assign g[28345] = b[13] & g[11962];
assign g[20155] = a[13] & g[11963];
assign g[28346] = b[13] & g[11963];
assign g[20156] = a[13] & g[11964];
assign g[28347] = b[13] & g[11964];
assign g[20157] = a[13] & g[11965];
assign g[28348] = b[13] & g[11965];
assign g[20158] = a[13] & g[11966];
assign g[28349] = b[13] & g[11966];
assign g[20159] = a[13] & g[11967];
assign g[28350] = b[13] & g[11967];
assign g[20160] = a[13] & g[11968];
assign g[28351] = b[13] & g[11968];
assign g[20161] = a[13] & g[11969];
assign g[28352] = b[13] & g[11969];
assign g[20162] = a[13] & g[11970];
assign g[28353] = b[13] & g[11970];
assign g[20163] = a[13] & g[11971];
assign g[28354] = b[13] & g[11971];
assign g[20164] = a[13] & g[11972];
assign g[28355] = b[13] & g[11972];
assign g[20165] = a[13] & g[11973];
assign g[28356] = b[13] & g[11973];
assign g[20166] = a[13] & g[11974];
assign g[28357] = b[13] & g[11974];
assign g[20167] = a[13] & g[11975];
assign g[28358] = b[13] & g[11975];
assign g[20168] = a[13] & g[11976];
assign g[28359] = b[13] & g[11976];
assign g[20169] = a[13] & g[11977];
assign g[28360] = b[13] & g[11977];
assign g[20170] = a[13] & g[11978];
assign g[28361] = b[13] & g[11978];
assign g[20171] = a[13] & g[11979];
assign g[28362] = b[13] & g[11979];
assign g[20172] = a[13] & g[11980];
assign g[28363] = b[13] & g[11980];
assign g[20173] = a[13] & g[11981];
assign g[28364] = b[13] & g[11981];
assign g[20174] = a[13] & g[11982];
assign g[28365] = b[13] & g[11982];
assign g[20175] = a[13] & g[11983];
assign g[28366] = b[13] & g[11983];
assign g[20176] = a[13] & g[11984];
assign g[28367] = b[13] & g[11984];
assign g[20177] = a[13] & g[11985];
assign g[28368] = b[13] & g[11985];
assign g[20178] = a[13] & g[11986];
assign g[28369] = b[13] & g[11986];
assign g[20179] = a[13] & g[11987];
assign g[28370] = b[13] & g[11987];
assign g[20180] = a[13] & g[11988];
assign g[28371] = b[13] & g[11988];
assign g[20181] = a[13] & g[11989];
assign g[28372] = b[13] & g[11989];
assign g[20182] = a[13] & g[11990];
assign g[28373] = b[13] & g[11990];
assign g[20183] = a[13] & g[11991];
assign g[28374] = b[13] & g[11991];
assign g[20184] = a[13] & g[11992];
assign g[28375] = b[13] & g[11992];
assign g[20185] = a[13] & g[11993];
assign g[28376] = b[13] & g[11993];
assign g[20186] = a[13] & g[11994];
assign g[28377] = b[13] & g[11994];
assign g[20187] = a[13] & g[11995];
assign g[28378] = b[13] & g[11995];
assign g[20188] = a[13] & g[11996];
assign g[28379] = b[13] & g[11996];
assign g[20189] = a[13] & g[11997];
assign g[28380] = b[13] & g[11997];
assign g[20190] = a[13] & g[11998];
assign g[28381] = b[13] & g[11998];
assign g[20191] = a[13] & g[11999];
assign g[28382] = b[13] & g[11999];
assign g[20192] = a[13] & g[12000];
assign g[28383] = b[13] & g[12000];
assign g[20193] = a[13] & g[12001];
assign g[28384] = b[13] & g[12001];
assign g[20194] = a[13] & g[12002];
assign g[28385] = b[13] & g[12002];
assign g[20195] = a[13] & g[12003];
assign g[28386] = b[13] & g[12003];
assign g[20196] = a[13] & g[12004];
assign g[28387] = b[13] & g[12004];
assign g[20197] = a[13] & g[12005];
assign g[28388] = b[13] & g[12005];
assign g[20198] = a[13] & g[12006];
assign g[28389] = b[13] & g[12006];
assign g[20199] = a[13] & g[12007];
assign g[28390] = b[13] & g[12007];
assign g[20200] = a[13] & g[12008];
assign g[28391] = b[13] & g[12008];
assign g[20201] = a[13] & g[12009];
assign g[28392] = b[13] & g[12009];
assign g[20202] = a[13] & g[12010];
assign g[28393] = b[13] & g[12010];
assign g[20203] = a[13] & g[12011];
assign g[28394] = b[13] & g[12011];
assign g[20204] = a[13] & g[12012];
assign g[28395] = b[13] & g[12012];
assign g[20205] = a[13] & g[12013];
assign g[28396] = b[13] & g[12013];
assign g[20206] = a[13] & g[12014];
assign g[28397] = b[13] & g[12014];
assign g[20207] = a[13] & g[12015];
assign g[28398] = b[13] & g[12015];
assign g[20208] = a[13] & g[12016];
assign g[28399] = b[13] & g[12016];
assign g[20209] = a[13] & g[12017];
assign g[28400] = b[13] & g[12017];
assign g[20210] = a[13] & g[12018];
assign g[28401] = b[13] & g[12018];
assign g[20211] = a[13] & g[12019];
assign g[28402] = b[13] & g[12019];
assign g[20212] = a[13] & g[12020];
assign g[28403] = b[13] & g[12020];
assign g[20213] = a[13] & g[12021];
assign g[28404] = b[13] & g[12021];
assign g[20214] = a[13] & g[12022];
assign g[28405] = b[13] & g[12022];
assign g[20215] = a[13] & g[12023];
assign g[28406] = b[13] & g[12023];
assign g[20216] = a[13] & g[12024];
assign g[28407] = b[13] & g[12024];
assign g[20217] = a[13] & g[12025];
assign g[28408] = b[13] & g[12025];
assign g[20218] = a[13] & g[12026];
assign g[28409] = b[13] & g[12026];
assign g[20219] = a[13] & g[12027];
assign g[28410] = b[13] & g[12027];
assign g[20220] = a[13] & g[12028];
assign g[28411] = b[13] & g[12028];
assign g[20221] = a[13] & g[12029];
assign g[28412] = b[13] & g[12029];
assign g[20222] = a[13] & g[12030];
assign g[28413] = b[13] & g[12030];
assign g[20223] = a[13] & g[12031];
assign g[28414] = b[13] & g[12031];
assign g[20224] = a[13] & g[12032];
assign g[28415] = b[13] & g[12032];
assign g[20225] = a[13] & g[12033];
assign g[28416] = b[13] & g[12033];
assign g[20226] = a[13] & g[12034];
assign g[28417] = b[13] & g[12034];
assign g[20227] = a[13] & g[12035];
assign g[28418] = b[13] & g[12035];
assign g[20228] = a[13] & g[12036];
assign g[28419] = b[13] & g[12036];
assign g[20229] = a[13] & g[12037];
assign g[28420] = b[13] & g[12037];
assign g[20230] = a[13] & g[12038];
assign g[28421] = b[13] & g[12038];
assign g[20231] = a[13] & g[12039];
assign g[28422] = b[13] & g[12039];
assign g[20232] = a[13] & g[12040];
assign g[28423] = b[13] & g[12040];
assign g[20233] = a[13] & g[12041];
assign g[28424] = b[13] & g[12041];
assign g[20234] = a[13] & g[12042];
assign g[28425] = b[13] & g[12042];
assign g[20235] = a[13] & g[12043];
assign g[28426] = b[13] & g[12043];
assign g[20236] = a[13] & g[12044];
assign g[28427] = b[13] & g[12044];
assign g[20237] = a[13] & g[12045];
assign g[28428] = b[13] & g[12045];
assign g[20238] = a[13] & g[12046];
assign g[28429] = b[13] & g[12046];
assign g[20239] = a[13] & g[12047];
assign g[28430] = b[13] & g[12047];
assign g[20240] = a[13] & g[12048];
assign g[28431] = b[13] & g[12048];
assign g[20241] = a[13] & g[12049];
assign g[28432] = b[13] & g[12049];
assign g[20242] = a[13] & g[12050];
assign g[28433] = b[13] & g[12050];
assign g[20243] = a[13] & g[12051];
assign g[28434] = b[13] & g[12051];
assign g[20244] = a[13] & g[12052];
assign g[28435] = b[13] & g[12052];
assign g[20245] = a[13] & g[12053];
assign g[28436] = b[13] & g[12053];
assign g[20246] = a[13] & g[12054];
assign g[28437] = b[13] & g[12054];
assign g[20247] = a[13] & g[12055];
assign g[28438] = b[13] & g[12055];
assign g[20248] = a[13] & g[12056];
assign g[28439] = b[13] & g[12056];
assign g[20249] = a[13] & g[12057];
assign g[28440] = b[13] & g[12057];
assign g[20250] = a[13] & g[12058];
assign g[28441] = b[13] & g[12058];
assign g[20251] = a[13] & g[12059];
assign g[28442] = b[13] & g[12059];
assign g[20252] = a[13] & g[12060];
assign g[28443] = b[13] & g[12060];
assign g[20253] = a[13] & g[12061];
assign g[28444] = b[13] & g[12061];
assign g[20254] = a[13] & g[12062];
assign g[28445] = b[13] & g[12062];
assign g[20255] = a[13] & g[12063];
assign g[28446] = b[13] & g[12063];
assign g[20256] = a[13] & g[12064];
assign g[28447] = b[13] & g[12064];
assign g[20257] = a[13] & g[12065];
assign g[28448] = b[13] & g[12065];
assign g[20258] = a[13] & g[12066];
assign g[28449] = b[13] & g[12066];
assign g[20259] = a[13] & g[12067];
assign g[28450] = b[13] & g[12067];
assign g[20260] = a[13] & g[12068];
assign g[28451] = b[13] & g[12068];
assign g[20261] = a[13] & g[12069];
assign g[28452] = b[13] & g[12069];
assign g[20262] = a[13] & g[12070];
assign g[28453] = b[13] & g[12070];
assign g[20263] = a[13] & g[12071];
assign g[28454] = b[13] & g[12071];
assign g[20264] = a[13] & g[12072];
assign g[28455] = b[13] & g[12072];
assign g[20265] = a[13] & g[12073];
assign g[28456] = b[13] & g[12073];
assign g[20266] = a[13] & g[12074];
assign g[28457] = b[13] & g[12074];
assign g[20267] = a[13] & g[12075];
assign g[28458] = b[13] & g[12075];
assign g[20268] = a[13] & g[12076];
assign g[28459] = b[13] & g[12076];
assign g[20269] = a[13] & g[12077];
assign g[28460] = b[13] & g[12077];
assign g[20270] = a[13] & g[12078];
assign g[28461] = b[13] & g[12078];
assign g[20271] = a[13] & g[12079];
assign g[28462] = b[13] & g[12079];
assign g[20272] = a[13] & g[12080];
assign g[28463] = b[13] & g[12080];
assign g[20273] = a[13] & g[12081];
assign g[28464] = b[13] & g[12081];
assign g[20274] = a[13] & g[12082];
assign g[28465] = b[13] & g[12082];
assign g[20275] = a[13] & g[12083];
assign g[28466] = b[13] & g[12083];
assign g[20276] = a[13] & g[12084];
assign g[28467] = b[13] & g[12084];
assign g[20277] = a[13] & g[12085];
assign g[28468] = b[13] & g[12085];
assign g[20278] = a[13] & g[12086];
assign g[28469] = b[13] & g[12086];
assign g[20279] = a[13] & g[12087];
assign g[28470] = b[13] & g[12087];
assign g[20280] = a[13] & g[12088];
assign g[28471] = b[13] & g[12088];
assign g[20281] = a[13] & g[12089];
assign g[28472] = b[13] & g[12089];
assign g[20282] = a[13] & g[12090];
assign g[28473] = b[13] & g[12090];
assign g[20283] = a[13] & g[12091];
assign g[28474] = b[13] & g[12091];
assign g[20284] = a[13] & g[12092];
assign g[28475] = b[13] & g[12092];
assign g[20285] = a[13] & g[12093];
assign g[28476] = b[13] & g[12093];
assign g[20286] = a[13] & g[12094];
assign g[28477] = b[13] & g[12094];
assign g[20287] = a[13] & g[12095];
assign g[28478] = b[13] & g[12095];
assign g[20288] = a[13] & g[12096];
assign g[28479] = b[13] & g[12096];
assign g[20289] = a[13] & g[12097];
assign g[28480] = b[13] & g[12097];
assign g[20290] = a[13] & g[12098];
assign g[28481] = b[13] & g[12098];
assign g[20291] = a[13] & g[12099];
assign g[28482] = b[13] & g[12099];
assign g[20292] = a[13] & g[12100];
assign g[28483] = b[13] & g[12100];
assign g[20293] = a[13] & g[12101];
assign g[28484] = b[13] & g[12101];
assign g[20294] = a[13] & g[12102];
assign g[28485] = b[13] & g[12102];
assign g[20295] = a[13] & g[12103];
assign g[28486] = b[13] & g[12103];
assign g[20296] = a[13] & g[12104];
assign g[28487] = b[13] & g[12104];
assign g[20297] = a[13] & g[12105];
assign g[28488] = b[13] & g[12105];
assign g[20298] = a[13] & g[12106];
assign g[28489] = b[13] & g[12106];
assign g[20299] = a[13] & g[12107];
assign g[28490] = b[13] & g[12107];
assign g[20300] = a[13] & g[12108];
assign g[28491] = b[13] & g[12108];
assign g[20301] = a[13] & g[12109];
assign g[28492] = b[13] & g[12109];
assign g[20302] = a[13] & g[12110];
assign g[28493] = b[13] & g[12110];
assign g[20303] = a[13] & g[12111];
assign g[28494] = b[13] & g[12111];
assign g[20304] = a[13] & g[12112];
assign g[28495] = b[13] & g[12112];
assign g[20305] = a[13] & g[12113];
assign g[28496] = b[13] & g[12113];
assign g[20306] = a[13] & g[12114];
assign g[28497] = b[13] & g[12114];
assign g[20307] = a[13] & g[12115];
assign g[28498] = b[13] & g[12115];
assign g[20308] = a[13] & g[12116];
assign g[28499] = b[13] & g[12116];
assign g[20309] = a[13] & g[12117];
assign g[28500] = b[13] & g[12117];
assign g[20310] = a[13] & g[12118];
assign g[28501] = b[13] & g[12118];
assign g[20311] = a[13] & g[12119];
assign g[28502] = b[13] & g[12119];
assign g[20312] = a[13] & g[12120];
assign g[28503] = b[13] & g[12120];
assign g[20313] = a[13] & g[12121];
assign g[28504] = b[13] & g[12121];
assign g[20314] = a[13] & g[12122];
assign g[28505] = b[13] & g[12122];
assign g[20315] = a[13] & g[12123];
assign g[28506] = b[13] & g[12123];
assign g[20316] = a[13] & g[12124];
assign g[28507] = b[13] & g[12124];
assign g[20317] = a[13] & g[12125];
assign g[28508] = b[13] & g[12125];
assign g[20318] = a[13] & g[12126];
assign g[28509] = b[13] & g[12126];
assign g[20319] = a[13] & g[12127];
assign g[28510] = b[13] & g[12127];
assign g[20320] = a[13] & g[12128];
assign g[28511] = b[13] & g[12128];
assign g[20321] = a[13] & g[12129];
assign g[28512] = b[13] & g[12129];
assign g[20322] = a[13] & g[12130];
assign g[28513] = b[13] & g[12130];
assign g[20323] = a[13] & g[12131];
assign g[28514] = b[13] & g[12131];
assign g[20324] = a[13] & g[12132];
assign g[28515] = b[13] & g[12132];
assign g[20325] = a[13] & g[12133];
assign g[28516] = b[13] & g[12133];
assign g[20326] = a[13] & g[12134];
assign g[28517] = b[13] & g[12134];
assign g[20327] = a[13] & g[12135];
assign g[28518] = b[13] & g[12135];
assign g[20328] = a[13] & g[12136];
assign g[28519] = b[13] & g[12136];
assign g[20329] = a[13] & g[12137];
assign g[28520] = b[13] & g[12137];
assign g[20330] = a[13] & g[12138];
assign g[28521] = b[13] & g[12138];
assign g[20331] = a[13] & g[12139];
assign g[28522] = b[13] & g[12139];
assign g[20332] = a[13] & g[12140];
assign g[28523] = b[13] & g[12140];
assign g[20333] = a[13] & g[12141];
assign g[28524] = b[13] & g[12141];
assign g[20334] = a[13] & g[12142];
assign g[28525] = b[13] & g[12142];
assign g[20335] = a[13] & g[12143];
assign g[28526] = b[13] & g[12143];
assign g[20336] = a[13] & g[12144];
assign g[28527] = b[13] & g[12144];
assign g[20337] = a[13] & g[12145];
assign g[28528] = b[13] & g[12145];
assign g[20338] = a[13] & g[12146];
assign g[28529] = b[13] & g[12146];
assign g[20339] = a[13] & g[12147];
assign g[28530] = b[13] & g[12147];
assign g[20340] = a[13] & g[12148];
assign g[28531] = b[13] & g[12148];
assign g[20341] = a[13] & g[12149];
assign g[28532] = b[13] & g[12149];
assign g[20342] = a[13] & g[12150];
assign g[28533] = b[13] & g[12150];
assign g[20343] = a[13] & g[12151];
assign g[28534] = b[13] & g[12151];
assign g[20344] = a[13] & g[12152];
assign g[28535] = b[13] & g[12152];
assign g[20345] = a[13] & g[12153];
assign g[28536] = b[13] & g[12153];
assign g[20346] = a[13] & g[12154];
assign g[28537] = b[13] & g[12154];
assign g[20347] = a[13] & g[12155];
assign g[28538] = b[13] & g[12155];
assign g[20348] = a[13] & g[12156];
assign g[28539] = b[13] & g[12156];
assign g[20349] = a[13] & g[12157];
assign g[28540] = b[13] & g[12157];
assign g[20350] = a[13] & g[12158];
assign g[28541] = b[13] & g[12158];
assign g[20351] = a[13] & g[12159];
assign g[28542] = b[13] & g[12159];
assign g[20352] = a[13] & g[12160];
assign g[28543] = b[13] & g[12160];
assign g[20353] = a[13] & g[12161];
assign g[28544] = b[13] & g[12161];
assign g[20354] = a[13] & g[12162];
assign g[28545] = b[13] & g[12162];
assign g[20355] = a[13] & g[12163];
assign g[28546] = b[13] & g[12163];
assign g[20356] = a[13] & g[12164];
assign g[28547] = b[13] & g[12164];
assign g[20357] = a[13] & g[12165];
assign g[28548] = b[13] & g[12165];
assign g[20358] = a[13] & g[12166];
assign g[28549] = b[13] & g[12166];
assign g[20359] = a[13] & g[12167];
assign g[28550] = b[13] & g[12167];
assign g[20360] = a[13] & g[12168];
assign g[28551] = b[13] & g[12168];
assign g[20361] = a[13] & g[12169];
assign g[28552] = b[13] & g[12169];
assign g[20362] = a[13] & g[12170];
assign g[28553] = b[13] & g[12170];
assign g[20363] = a[13] & g[12171];
assign g[28554] = b[13] & g[12171];
assign g[20364] = a[13] & g[12172];
assign g[28555] = b[13] & g[12172];
assign g[20365] = a[13] & g[12173];
assign g[28556] = b[13] & g[12173];
assign g[20366] = a[13] & g[12174];
assign g[28557] = b[13] & g[12174];
assign g[20367] = a[13] & g[12175];
assign g[28558] = b[13] & g[12175];
assign g[20368] = a[13] & g[12176];
assign g[28559] = b[13] & g[12176];
assign g[20369] = a[13] & g[12177];
assign g[28560] = b[13] & g[12177];
assign g[20370] = a[13] & g[12178];
assign g[28561] = b[13] & g[12178];
assign g[20371] = a[13] & g[12179];
assign g[28562] = b[13] & g[12179];
assign g[20372] = a[13] & g[12180];
assign g[28563] = b[13] & g[12180];
assign g[20373] = a[13] & g[12181];
assign g[28564] = b[13] & g[12181];
assign g[20374] = a[13] & g[12182];
assign g[28565] = b[13] & g[12182];
assign g[20375] = a[13] & g[12183];
assign g[28566] = b[13] & g[12183];
assign g[20376] = a[13] & g[12184];
assign g[28567] = b[13] & g[12184];
assign g[20377] = a[13] & g[12185];
assign g[28568] = b[13] & g[12185];
assign g[20378] = a[13] & g[12186];
assign g[28569] = b[13] & g[12186];
assign g[20379] = a[13] & g[12187];
assign g[28570] = b[13] & g[12187];
assign g[20380] = a[13] & g[12188];
assign g[28571] = b[13] & g[12188];
assign g[20381] = a[13] & g[12189];
assign g[28572] = b[13] & g[12189];
assign g[20382] = a[13] & g[12190];
assign g[28573] = b[13] & g[12190];
assign g[20383] = a[13] & g[12191];
assign g[28574] = b[13] & g[12191];
assign g[20384] = a[13] & g[12192];
assign g[28575] = b[13] & g[12192];
assign g[20385] = a[13] & g[12193];
assign g[28576] = b[13] & g[12193];
assign g[20386] = a[13] & g[12194];
assign g[28577] = b[13] & g[12194];
assign g[20387] = a[13] & g[12195];
assign g[28578] = b[13] & g[12195];
assign g[20388] = a[13] & g[12196];
assign g[28579] = b[13] & g[12196];
assign g[20389] = a[13] & g[12197];
assign g[28580] = b[13] & g[12197];
assign g[20390] = a[13] & g[12198];
assign g[28581] = b[13] & g[12198];
assign g[20391] = a[13] & g[12199];
assign g[28582] = b[13] & g[12199];
assign g[20392] = a[13] & g[12200];
assign g[28583] = b[13] & g[12200];
assign g[20393] = a[13] & g[12201];
assign g[28584] = b[13] & g[12201];
assign g[20394] = a[13] & g[12202];
assign g[28585] = b[13] & g[12202];
assign g[20395] = a[13] & g[12203];
assign g[28586] = b[13] & g[12203];
assign g[20396] = a[13] & g[12204];
assign g[28587] = b[13] & g[12204];
assign g[20397] = a[13] & g[12205];
assign g[28588] = b[13] & g[12205];
assign g[20398] = a[13] & g[12206];
assign g[28589] = b[13] & g[12206];
assign g[20399] = a[13] & g[12207];
assign g[28590] = b[13] & g[12207];
assign g[20400] = a[13] & g[12208];
assign g[28591] = b[13] & g[12208];
assign g[20401] = a[13] & g[12209];
assign g[28592] = b[13] & g[12209];
assign g[20402] = a[13] & g[12210];
assign g[28593] = b[13] & g[12210];
assign g[20403] = a[13] & g[12211];
assign g[28594] = b[13] & g[12211];
assign g[20404] = a[13] & g[12212];
assign g[28595] = b[13] & g[12212];
assign g[20405] = a[13] & g[12213];
assign g[28596] = b[13] & g[12213];
assign g[20406] = a[13] & g[12214];
assign g[28597] = b[13] & g[12214];
assign g[20407] = a[13] & g[12215];
assign g[28598] = b[13] & g[12215];
assign g[20408] = a[13] & g[12216];
assign g[28599] = b[13] & g[12216];
assign g[20409] = a[13] & g[12217];
assign g[28600] = b[13] & g[12217];
assign g[20410] = a[13] & g[12218];
assign g[28601] = b[13] & g[12218];
assign g[20411] = a[13] & g[12219];
assign g[28602] = b[13] & g[12219];
assign g[20412] = a[13] & g[12220];
assign g[28603] = b[13] & g[12220];
assign g[20413] = a[13] & g[12221];
assign g[28604] = b[13] & g[12221];
assign g[20414] = a[13] & g[12222];
assign g[28605] = b[13] & g[12222];
assign g[20415] = a[13] & g[12223];
assign g[28606] = b[13] & g[12223];
assign g[20416] = a[13] & g[12224];
assign g[28607] = b[13] & g[12224];
assign g[20417] = a[13] & g[12225];
assign g[28608] = b[13] & g[12225];
assign g[20418] = a[13] & g[12226];
assign g[28609] = b[13] & g[12226];
assign g[20419] = a[13] & g[12227];
assign g[28610] = b[13] & g[12227];
assign g[20420] = a[13] & g[12228];
assign g[28611] = b[13] & g[12228];
assign g[20421] = a[13] & g[12229];
assign g[28612] = b[13] & g[12229];
assign g[20422] = a[13] & g[12230];
assign g[28613] = b[13] & g[12230];
assign g[20423] = a[13] & g[12231];
assign g[28614] = b[13] & g[12231];
assign g[20424] = a[13] & g[12232];
assign g[28615] = b[13] & g[12232];
assign g[20425] = a[13] & g[12233];
assign g[28616] = b[13] & g[12233];
assign g[20426] = a[13] & g[12234];
assign g[28617] = b[13] & g[12234];
assign g[20427] = a[13] & g[12235];
assign g[28618] = b[13] & g[12235];
assign g[20428] = a[13] & g[12236];
assign g[28619] = b[13] & g[12236];
assign g[20429] = a[13] & g[12237];
assign g[28620] = b[13] & g[12237];
assign g[20430] = a[13] & g[12238];
assign g[28621] = b[13] & g[12238];
assign g[20431] = a[13] & g[12239];
assign g[28622] = b[13] & g[12239];
assign g[20432] = a[13] & g[12240];
assign g[28623] = b[13] & g[12240];
assign g[20433] = a[13] & g[12241];
assign g[28624] = b[13] & g[12241];
assign g[20434] = a[13] & g[12242];
assign g[28625] = b[13] & g[12242];
assign g[20435] = a[13] & g[12243];
assign g[28626] = b[13] & g[12243];
assign g[20436] = a[13] & g[12244];
assign g[28627] = b[13] & g[12244];
assign g[20437] = a[13] & g[12245];
assign g[28628] = b[13] & g[12245];
assign g[20438] = a[13] & g[12246];
assign g[28629] = b[13] & g[12246];
assign g[20439] = a[13] & g[12247];
assign g[28630] = b[13] & g[12247];
assign g[20440] = a[13] & g[12248];
assign g[28631] = b[13] & g[12248];
assign g[20441] = a[13] & g[12249];
assign g[28632] = b[13] & g[12249];
assign g[20442] = a[13] & g[12250];
assign g[28633] = b[13] & g[12250];
assign g[20443] = a[13] & g[12251];
assign g[28634] = b[13] & g[12251];
assign g[20444] = a[13] & g[12252];
assign g[28635] = b[13] & g[12252];
assign g[20445] = a[13] & g[12253];
assign g[28636] = b[13] & g[12253];
assign g[20446] = a[13] & g[12254];
assign g[28637] = b[13] & g[12254];
assign g[20447] = a[13] & g[12255];
assign g[28638] = b[13] & g[12255];
assign g[20448] = a[13] & g[12256];
assign g[28639] = b[13] & g[12256];
assign g[20449] = a[13] & g[12257];
assign g[28640] = b[13] & g[12257];
assign g[20450] = a[13] & g[12258];
assign g[28641] = b[13] & g[12258];
assign g[20451] = a[13] & g[12259];
assign g[28642] = b[13] & g[12259];
assign g[20452] = a[13] & g[12260];
assign g[28643] = b[13] & g[12260];
assign g[20453] = a[13] & g[12261];
assign g[28644] = b[13] & g[12261];
assign g[20454] = a[13] & g[12262];
assign g[28645] = b[13] & g[12262];
assign g[20455] = a[13] & g[12263];
assign g[28646] = b[13] & g[12263];
assign g[20456] = a[13] & g[12264];
assign g[28647] = b[13] & g[12264];
assign g[20457] = a[13] & g[12265];
assign g[28648] = b[13] & g[12265];
assign g[20458] = a[13] & g[12266];
assign g[28649] = b[13] & g[12266];
assign g[20459] = a[13] & g[12267];
assign g[28650] = b[13] & g[12267];
assign g[20460] = a[13] & g[12268];
assign g[28651] = b[13] & g[12268];
assign g[20461] = a[13] & g[12269];
assign g[28652] = b[13] & g[12269];
assign g[20462] = a[13] & g[12270];
assign g[28653] = b[13] & g[12270];
assign g[20463] = a[13] & g[12271];
assign g[28654] = b[13] & g[12271];
assign g[20464] = a[13] & g[12272];
assign g[28655] = b[13] & g[12272];
assign g[20465] = a[13] & g[12273];
assign g[28656] = b[13] & g[12273];
assign g[20466] = a[13] & g[12274];
assign g[28657] = b[13] & g[12274];
assign g[20467] = a[13] & g[12275];
assign g[28658] = b[13] & g[12275];
assign g[20468] = a[13] & g[12276];
assign g[28659] = b[13] & g[12276];
assign g[20469] = a[13] & g[12277];
assign g[28660] = b[13] & g[12277];
assign g[20470] = a[13] & g[12278];
assign g[28661] = b[13] & g[12278];
assign g[20471] = a[13] & g[12279];
assign g[28662] = b[13] & g[12279];
assign g[20472] = a[13] & g[12280];
assign g[28663] = b[13] & g[12280];
assign g[20473] = a[13] & g[12281];
assign g[28664] = b[13] & g[12281];
assign g[20474] = a[13] & g[12282];
assign g[28665] = b[13] & g[12282];
assign g[20475] = a[13] & g[12283];
assign g[28666] = b[13] & g[12283];
assign g[20476] = a[13] & g[12284];
assign g[28667] = b[13] & g[12284];
assign g[20477] = a[13] & g[12285];
assign g[28668] = b[13] & g[12285];
assign g[20478] = a[13] & g[12286];
assign g[28669] = b[13] & g[12286];
assign g[20479] = a[13] & g[12287];
assign g[28670] = b[13] & g[12287];
assign g[20480] = a[13] & g[12288];
assign g[28671] = b[13] & g[12288];
assign g[20481] = a[13] & g[12289];
assign g[28672] = b[13] & g[12289];
assign g[20482] = a[13] & g[12290];
assign g[28673] = b[13] & g[12290];
assign g[20483] = a[13] & g[12291];
assign g[28674] = b[13] & g[12291];
assign g[20484] = a[13] & g[12292];
assign g[28675] = b[13] & g[12292];
assign g[20485] = a[13] & g[12293];
assign g[28676] = b[13] & g[12293];
assign g[20486] = a[13] & g[12294];
assign g[28677] = b[13] & g[12294];
assign g[20487] = a[13] & g[12295];
assign g[28678] = b[13] & g[12295];
assign g[20488] = a[13] & g[12296];
assign g[28679] = b[13] & g[12296];
assign g[20489] = a[13] & g[12297];
assign g[28680] = b[13] & g[12297];
assign g[20490] = a[13] & g[12298];
assign g[28681] = b[13] & g[12298];
assign g[20491] = a[13] & g[12299];
assign g[28682] = b[13] & g[12299];
assign g[20492] = a[13] & g[12300];
assign g[28683] = b[13] & g[12300];
assign g[20493] = a[13] & g[12301];
assign g[28684] = b[13] & g[12301];
assign g[20494] = a[13] & g[12302];
assign g[28685] = b[13] & g[12302];
assign g[20495] = a[13] & g[12303];
assign g[28686] = b[13] & g[12303];
assign g[20496] = a[13] & g[12304];
assign g[28687] = b[13] & g[12304];
assign g[20497] = a[13] & g[12305];
assign g[28688] = b[13] & g[12305];
assign g[20498] = a[13] & g[12306];
assign g[28689] = b[13] & g[12306];
assign g[20499] = a[13] & g[12307];
assign g[28690] = b[13] & g[12307];
assign g[20500] = a[13] & g[12308];
assign g[28691] = b[13] & g[12308];
assign g[20501] = a[13] & g[12309];
assign g[28692] = b[13] & g[12309];
assign g[20502] = a[13] & g[12310];
assign g[28693] = b[13] & g[12310];
assign g[20503] = a[13] & g[12311];
assign g[28694] = b[13] & g[12311];
assign g[20504] = a[13] & g[12312];
assign g[28695] = b[13] & g[12312];
assign g[20505] = a[13] & g[12313];
assign g[28696] = b[13] & g[12313];
assign g[20506] = a[13] & g[12314];
assign g[28697] = b[13] & g[12314];
assign g[20507] = a[13] & g[12315];
assign g[28698] = b[13] & g[12315];
assign g[20508] = a[13] & g[12316];
assign g[28699] = b[13] & g[12316];
assign g[20509] = a[13] & g[12317];
assign g[28700] = b[13] & g[12317];
assign g[20510] = a[13] & g[12318];
assign g[28701] = b[13] & g[12318];
assign g[20511] = a[13] & g[12319];
assign g[28702] = b[13] & g[12319];
assign g[20512] = a[13] & g[12320];
assign g[28703] = b[13] & g[12320];
assign g[20513] = a[13] & g[12321];
assign g[28704] = b[13] & g[12321];
assign g[20514] = a[13] & g[12322];
assign g[28705] = b[13] & g[12322];
assign g[20515] = a[13] & g[12323];
assign g[28706] = b[13] & g[12323];
assign g[20516] = a[13] & g[12324];
assign g[28707] = b[13] & g[12324];
assign g[20517] = a[13] & g[12325];
assign g[28708] = b[13] & g[12325];
assign g[20518] = a[13] & g[12326];
assign g[28709] = b[13] & g[12326];
assign g[20519] = a[13] & g[12327];
assign g[28710] = b[13] & g[12327];
assign g[20520] = a[13] & g[12328];
assign g[28711] = b[13] & g[12328];
assign g[20521] = a[13] & g[12329];
assign g[28712] = b[13] & g[12329];
assign g[20522] = a[13] & g[12330];
assign g[28713] = b[13] & g[12330];
assign g[20523] = a[13] & g[12331];
assign g[28714] = b[13] & g[12331];
assign g[20524] = a[13] & g[12332];
assign g[28715] = b[13] & g[12332];
assign g[20525] = a[13] & g[12333];
assign g[28716] = b[13] & g[12333];
assign g[20526] = a[13] & g[12334];
assign g[28717] = b[13] & g[12334];
assign g[20527] = a[13] & g[12335];
assign g[28718] = b[13] & g[12335];
assign g[20528] = a[13] & g[12336];
assign g[28719] = b[13] & g[12336];
assign g[20529] = a[13] & g[12337];
assign g[28720] = b[13] & g[12337];
assign g[20530] = a[13] & g[12338];
assign g[28721] = b[13] & g[12338];
assign g[20531] = a[13] & g[12339];
assign g[28722] = b[13] & g[12339];
assign g[20532] = a[13] & g[12340];
assign g[28723] = b[13] & g[12340];
assign g[20533] = a[13] & g[12341];
assign g[28724] = b[13] & g[12341];
assign g[20534] = a[13] & g[12342];
assign g[28725] = b[13] & g[12342];
assign g[20535] = a[13] & g[12343];
assign g[28726] = b[13] & g[12343];
assign g[20536] = a[13] & g[12344];
assign g[28727] = b[13] & g[12344];
assign g[20537] = a[13] & g[12345];
assign g[28728] = b[13] & g[12345];
assign g[20538] = a[13] & g[12346];
assign g[28729] = b[13] & g[12346];
assign g[20539] = a[13] & g[12347];
assign g[28730] = b[13] & g[12347];
assign g[20540] = a[13] & g[12348];
assign g[28731] = b[13] & g[12348];
assign g[20541] = a[13] & g[12349];
assign g[28732] = b[13] & g[12349];
assign g[20542] = a[13] & g[12350];
assign g[28733] = b[13] & g[12350];
assign g[20543] = a[13] & g[12351];
assign g[28734] = b[13] & g[12351];
assign g[20544] = a[13] & g[12352];
assign g[28735] = b[13] & g[12352];
assign g[20545] = a[13] & g[12353];
assign g[28736] = b[13] & g[12353];
assign g[20546] = a[13] & g[12354];
assign g[28737] = b[13] & g[12354];
assign g[20547] = a[13] & g[12355];
assign g[28738] = b[13] & g[12355];
assign g[20548] = a[13] & g[12356];
assign g[28739] = b[13] & g[12356];
assign g[20549] = a[13] & g[12357];
assign g[28740] = b[13] & g[12357];
assign g[20550] = a[13] & g[12358];
assign g[28741] = b[13] & g[12358];
assign g[20551] = a[13] & g[12359];
assign g[28742] = b[13] & g[12359];
assign g[20552] = a[13] & g[12360];
assign g[28743] = b[13] & g[12360];
assign g[20553] = a[13] & g[12361];
assign g[28744] = b[13] & g[12361];
assign g[20554] = a[13] & g[12362];
assign g[28745] = b[13] & g[12362];
assign g[20555] = a[13] & g[12363];
assign g[28746] = b[13] & g[12363];
assign g[20556] = a[13] & g[12364];
assign g[28747] = b[13] & g[12364];
assign g[20557] = a[13] & g[12365];
assign g[28748] = b[13] & g[12365];
assign g[20558] = a[13] & g[12366];
assign g[28749] = b[13] & g[12366];
assign g[20559] = a[13] & g[12367];
assign g[28750] = b[13] & g[12367];
assign g[20560] = a[13] & g[12368];
assign g[28751] = b[13] & g[12368];
assign g[20561] = a[13] & g[12369];
assign g[28752] = b[13] & g[12369];
assign g[20562] = a[13] & g[12370];
assign g[28753] = b[13] & g[12370];
assign g[20563] = a[13] & g[12371];
assign g[28754] = b[13] & g[12371];
assign g[20564] = a[13] & g[12372];
assign g[28755] = b[13] & g[12372];
assign g[20565] = a[13] & g[12373];
assign g[28756] = b[13] & g[12373];
assign g[20566] = a[13] & g[12374];
assign g[28757] = b[13] & g[12374];
assign g[20567] = a[13] & g[12375];
assign g[28758] = b[13] & g[12375];
assign g[20568] = a[13] & g[12376];
assign g[28759] = b[13] & g[12376];
assign g[20569] = a[13] & g[12377];
assign g[28760] = b[13] & g[12377];
assign g[20570] = a[13] & g[12378];
assign g[28761] = b[13] & g[12378];
assign g[20571] = a[13] & g[12379];
assign g[28762] = b[13] & g[12379];
assign g[20572] = a[13] & g[12380];
assign g[28763] = b[13] & g[12380];
assign g[20573] = a[13] & g[12381];
assign g[28764] = b[13] & g[12381];
assign g[20574] = a[13] & g[12382];
assign g[28765] = b[13] & g[12382];
assign g[20575] = a[13] & g[12383];
assign g[28766] = b[13] & g[12383];
assign g[20576] = a[13] & g[12384];
assign g[28767] = b[13] & g[12384];
assign g[20577] = a[13] & g[12385];
assign g[28768] = b[13] & g[12385];
assign g[20578] = a[13] & g[12386];
assign g[28769] = b[13] & g[12386];
assign g[20579] = a[13] & g[12387];
assign g[28770] = b[13] & g[12387];
assign g[20580] = a[13] & g[12388];
assign g[28771] = b[13] & g[12388];
assign g[20581] = a[13] & g[12389];
assign g[28772] = b[13] & g[12389];
assign g[20582] = a[13] & g[12390];
assign g[28773] = b[13] & g[12390];
assign g[20583] = a[13] & g[12391];
assign g[28774] = b[13] & g[12391];
assign g[20584] = a[13] & g[12392];
assign g[28775] = b[13] & g[12392];
assign g[20585] = a[13] & g[12393];
assign g[28776] = b[13] & g[12393];
assign g[20586] = a[13] & g[12394];
assign g[28777] = b[13] & g[12394];
assign g[20587] = a[13] & g[12395];
assign g[28778] = b[13] & g[12395];
assign g[20588] = a[13] & g[12396];
assign g[28779] = b[13] & g[12396];
assign g[20589] = a[13] & g[12397];
assign g[28780] = b[13] & g[12397];
assign g[20590] = a[13] & g[12398];
assign g[28781] = b[13] & g[12398];
assign g[20591] = a[13] & g[12399];
assign g[28782] = b[13] & g[12399];
assign g[20592] = a[13] & g[12400];
assign g[28783] = b[13] & g[12400];
assign g[20593] = a[13] & g[12401];
assign g[28784] = b[13] & g[12401];
assign g[20594] = a[13] & g[12402];
assign g[28785] = b[13] & g[12402];
assign g[20595] = a[13] & g[12403];
assign g[28786] = b[13] & g[12403];
assign g[20596] = a[13] & g[12404];
assign g[28787] = b[13] & g[12404];
assign g[20597] = a[13] & g[12405];
assign g[28788] = b[13] & g[12405];
assign g[20598] = a[13] & g[12406];
assign g[28789] = b[13] & g[12406];
assign g[20599] = a[13] & g[12407];
assign g[28790] = b[13] & g[12407];
assign g[20600] = a[13] & g[12408];
assign g[28791] = b[13] & g[12408];
assign g[20601] = a[13] & g[12409];
assign g[28792] = b[13] & g[12409];
assign g[20602] = a[13] & g[12410];
assign g[28793] = b[13] & g[12410];
assign g[20603] = a[13] & g[12411];
assign g[28794] = b[13] & g[12411];
assign g[20604] = a[13] & g[12412];
assign g[28795] = b[13] & g[12412];
assign g[20605] = a[13] & g[12413];
assign g[28796] = b[13] & g[12413];
assign g[20606] = a[13] & g[12414];
assign g[28797] = b[13] & g[12414];
assign g[20607] = a[13] & g[12415];
assign g[28798] = b[13] & g[12415];
assign g[20608] = a[13] & g[12416];
assign g[28799] = b[13] & g[12416];
assign g[20609] = a[13] & g[12417];
assign g[28800] = b[13] & g[12417];
assign g[20610] = a[13] & g[12418];
assign g[28801] = b[13] & g[12418];
assign g[20611] = a[13] & g[12419];
assign g[28802] = b[13] & g[12419];
assign g[20612] = a[13] & g[12420];
assign g[28803] = b[13] & g[12420];
assign g[20613] = a[13] & g[12421];
assign g[28804] = b[13] & g[12421];
assign g[20614] = a[13] & g[12422];
assign g[28805] = b[13] & g[12422];
assign g[20615] = a[13] & g[12423];
assign g[28806] = b[13] & g[12423];
assign g[20616] = a[13] & g[12424];
assign g[28807] = b[13] & g[12424];
assign g[20617] = a[13] & g[12425];
assign g[28808] = b[13] & g[12425];
assign g[20618] = a[13] & g[12426];
assign g[28809] = b[13] & g[12426];
assign g[20619] = a[13] & g[12427];
assign g[28810] = b[13] & g[12427];
assign g[20620] = a[13] & g[12428];
assign g[28811] = b[13] & g[12428];
assign g[20621] = a[13] & g[12429];
assign g[28812] = b[13] & g[12429];
assign g[20622] = a[13] & g[12430];
assign g[28813] = b[13] & g[12430];
assign g[20623] = a[13] & g[12431];
assign g[28814] = b[13] & g[12431];
assign g[20624] = a[13] & g[12432];
assign g[28815] = b[13] & g[12432];
assign g[20625] = a[13] & g[12433];
assign g[28816] = b[13] & g[12433];
assign g[20626] = a[13] & g[12434];
assign g[28817] = b[13] & g[12434];
assign g[20627] = a[13] & g[12435];
assign g[28818] = b[13] & g[12435];
assign g[20628] = a[13] & g[12436];
assign g[28819] = b[13] & g[12436];
assign g[20629] = a[13] & g[12437];
assign g[28820] = b[13] & g[12437];
assign g[20630] = a[13] & g[12438];
assign g[28821] = b[13] & g[12438];
assign g[20631] = a[13] & g[12439];
assign g[28822] = b[13] & g[12439];
assign g[20632] = a[13] & g[12440];
assign g[28823] = b[13] & g[12440];
assign g[20633] = a[13] & g[12441];
assign g[28824] = b[13] & g[12441];
assign g[20634] = a[13] & g[12442];
assign g[28825] = b[13] & g[12442];
assign g[20635] = a[13] & g[12443];
assign g[28826] = b[13] & g[12443];
assign g[20636] = a[13] & g[12444];
assign g[28827] = b[13] & g[12444];
assign g[20637] = a[13] & g[12445];
assign g[28828] = b[13] & g[12445];
assign g[20638] = a[13] & g[12446];
assign g[28829] = b[13] & g[12446];
assign g[20639] = a[13] & g[12447];
assign g[28830] = b[13] & g[12447];
assign g[20640] = a[13] & g[12448];
assign g[28831] = b[13] & g[12448];
assign g[20641] = a[13] & g[12449];
assign g[28832] = b[13] & g[12449];
assign g[20642] = a[13] & g[12450];
assign g[28833] = b[13] & g[12450];
assign g[20643] = a[13] & g[12451];
assign g[28834] = b[13] & g[12451];
assign g[20644] = a[13] & g[12452];
assign g[28835] = b[13] & g[12452];
assign g[20645] = a[13] & g[12453];
assign g[28836] = b[13] & g[12453];
assign g[20646] = a[13] & g[12454];
assign g[28837] = b[13] & g[12454];
assign g[20647] = a[13] & g[12455];
assign g[28838] = b[13] & g[12455];
assign g[20648] = a[13] & g[12456];
assign g[28839] = b[13] & g[12456];
assign g[20649] = a[13] & g[12457];
assign g[28840] = b[13] & g[12457];
assign g[20650] = a[13] & g[12458];
assign g[28841] = b[13] & g[12458];
assign g[20651] = a[13] & g[12459];
assign g[28842] = b[13] & g[12459];
assign g[20652] = a[13] & g[12460];
assign g[28843] = b[13] & g[12460];
assign g[20653] = a[13] & g[12461];
assign g[28844] = b[13] & g[12461];
assign g[20654] = a[13] & g[12462];
assign g[28845] = b[13] & g[12462];
assign g[20655] = a[13] & g[12463];
assign g[28846] = b[13] & g[12463];
assign g[20656] = a[13] & g[12464];
assign g[28847] = b[13] & g[12464];
assign g[20657] = a[13] & g[12465];
assign g[28848] = b[13] & g[12465];
assign g[20658] = a[13] & g[12466];
assign g[28849] = b[13] & g[12466];
assign g[20659] = a[13] & g[12467];
assign g[28850] = b[13] & g[12467];
assign g[20660] = a[13] & g[12468];
assign g[28851] = b[13] & g[12468];
assign g[20661] = a[13] & g[12469];
assign g[28852] = b[13] & g[12469];
assign g[20662] = a[13] & g[12470];
assign g[28853] = b[13] & g[12470];
assign g[20663] = a[13] & g[12471];
assign g[28854] = b[13] & g[12471];
assign g[20664] = a[13] & g[12472];
assign g[28855] = b[13] & g[12472];
assign g[20665] = a[13] & g[12473];
assign g[28856] = b[13] & g[12473];
assign g[20666] = a[13] & g[12474];
assign g[28857] = b[13] & g[12474];
assign g[20667] = a[13] & g[12475];
assign g[28858] = b[13] & g[12475];
assign g[20668] = a[13] & g[12476];
assign g[28859] = b[13] & g[12476];
assign g[20669] = a[13] & g[12477];
assign g[28860] = b[13] & g[12477];
assign g[20670] = a[13] & g[12478];
assign g[28861] = b[13] & g[12478];
assign g[20671] = a[13] & g[12479];
assign g[28862] = b[13] & g[12479];
assign g[20672] = a[13] & g[12480];
assign g[28863] = b[13] & g[12480];
assign g[20673] = a[13] & g[12481];
assign g[28864] = b[13] & g[12481];
assign g[20674] = a[13] & g[12482];
assign g[28865] = b[13] & g[12482];
assign g[20675] = a[13] & g[12483];
assign g[28866] = b[13] & g[12483];
assign g[20676] = a[13] & g[12484];
assign g[28867] = b[13] & g[12484];
assign g[20677] = a[13] & g[12485];
assign g[28868] = b[13] & g[12485];
assign g[20678] = a[13] & g[12486];
assign g[28869] = b[13] & g[12486];
assign g[20679] = a[13] & g[12487];
assign g[28870] = b[13] & g[12487];
assign g[20680] = a[13] & g[12488];
assign g[28871] = b[13] & g[12488];
assign g[20681] = a[13] & g[12489];
assign g[28872] = b[13] & g[12489];
assign g[20682] = a[13] & g[12490];
assign g[28873] = b[13] & g[12490];
assign g[20683] = a[13] & g[12491];
assign g[28874] = b[13] & g[12491];
assign g[20684] = a[13] & g[12492];
assign g[28875] = b[13] & g[12492];
assign g[20685] = a[13] & g[12493];
assign g[28876] = b[13] & g[12493];
assign g[20686] = a[13] & g[12494];
assign g[28877] = b[13] & g[12494];
assign g[20687] = a[13] & g[12495];
assign g[28878] = b[13] & g[12495];
assign g[20688] = a[13] & g[12496];
assign g[28879] = b[13] & g[12496];
assign g[20689] = a[13] & g[12497];
assign g[28880] = b[13] & g[12497];
assign g[20690] = a[13] & g[12498];
assign g[28881] = b[13] & g[12498];
assign g[20691] = a[13] & g[12499];
assign g[28882] = b[13] & g[12499];
assign g[20692] = a[13] & g[12500];
assign g[28883] = b[13] & g[12500];
assign g[20693] = a[13] & g[12501];
assign g[28884] = b[13] & g[12501];
assign g[20694] = a[13] & g[12502];
assign g[28885] = b[13] & g[12502];
assign g[20695] = a[13] & g[12503];
assign g[28886] = b[13] & g[12503];
assign g[20696] = a[13] & g[12504];
assign g[28887] = b[13] & g[12504];
assign g[20697] = a[13] & g[12505];
assign g[28888] = b[13] & g[12505];
assign g[20698] = a[13] & g[12506];
assign g[28889] = b[13] & g[12506];
assign g[20699] = a[13] & g[12507];
assign g[28890] = b[13] & g[12507];
assign g[20700] = a[13] & g[12508];
assign g[28891] = b[13] & g[12508];
assign g[20701] = a[13] & g[12509];
assign g[28892] = b[13] & g[12509];
assign g[20702] = a[13] & g[12510];
assign g[28893] = b[13] & g[12510];
assign g[20703] = a[13] & g[12511];
assign g[28894] = b[13] & g[12511];
assign g[20704] = a[13] & g[12512];
assign g[28895] = b[13] & g[12512];
assign g[20705] = a[13] & g[12513];
assign g[28896] = b[13] & g[12513];
assign g[20706] = a[13] & g[12514];
assign g[28897] = b[13] & g[12514];
assign g[20707] = a[13] & g[12515];
assign g[28898] = b[13] & g[12515];
assign g[20708] = a[13] & g[12516];
assign g[28899] = b[13] & g[12516];
assign g[20709] = a[13] & g[12517];
assign g[28900] = b[13] & g[12517];
assign g[20710] = a[13] & g[12518];
assign g[28901] = b[13] & g[12518];
assign g[20711] = a[13] & g[12519];
assign g[28902] = b[13] & g[12519];
assign g[20712] = a[13] & g[12520];
assign g[28903] = b[13] & g[12520];
assign g[20713] = a[13] & g[12521];
assign g[28904] = b[13] & g[12521];
assign g[20714] = a[13] & g[12522];
assign g[28905] = b[13] & g[12522];
assign g[20715] = a[13] & g[12523];
assign g[28906] = b[13] & g[12523];
assign g[20716] = a[13] & g[12524];
assign g[28907] = b[13] & g[12524];
assign g[20717] = a[13] & g[12525];
assign g[28908] = b[13] & g[12525];
assign g[20718] = a[13] & g[12526];
assign g[28909] = b[13] & g[12526];
assign g[20719] = a[13] & g[12527];
assign g[28910] = b[13] & g[12527];
assign g[20720] = a[13] & g[12528];
assign g[28911] = b[13] & g[12528];
assign g[20721] = a[13] & g[12529];
assign g[28912] = b[13] & g[12529];
assign g[20722] = a[13] & g[12530];
assign g[28913] = b[13] & g[12530];
assign g[20723] = a[13] & g[12531];
assign g[28914] = b[13] & g[12531];
assign g[20724] = a[13] & g[12532];
assign g[28915] = b[13] & g[12532];
assign g[20725] = a[13] & g[12533];
assign g[28916] = b[13] & g[12533];
assign g[20726] = a[13] & g[12534];
assign g[28917] = b[13] & g[12534];
assign g[20727] = a[13] & g[12535];
assign g[28918] = b[13] & g[12535];
assign g[20728] = a[13] & g[12536];
assign g[28919] = b[13] & g[12536];
assign g[20729] = a[13] & g[12537];
assign g[28920] = b[13] & g[12537];
assign g[20730] = a[13] & g[12538];
assign g[28921] = b[13] & g[12538];
assign g[20731] = a[13] & g[12539];
assign g[28922] = b[13] & g[12539];
assign g[20732] = a[13] & g[12540];
assign g[28923] = b[13] & g[12540];
assign g[20733] = a[13] & g[12541];
assign g[28924] = b[13] & g[12541];
assign g[20734] = a[13] & g[12542];
assign g[28925] = b[13] & g[12542];
assign g[20735] = a[13] & g[12543];
assign g[28926] = b[13] & g[12543];
assign g[20736] = a[13] & g[12544];
assign g[28927] = b[13] & g[12544];
assign g[20737] = a[13] & g[12545];
assign g[28928] = b[13] & g[12545];
assign g[20738] = a[13] & g[12546];
assign g[28929] = b[13] & g[12546];
assign g[20739] = a[13] & g[12547];
assign g[28930] = b[13] & g[12547];
assign g[20740] = a[13] & g[12548];
assign g[28931] = b[13] & g[12548];
assign g[20741] = a[13] & g[12549];
assign g[28932] = b[13] & g[12549];
assign g[20742] = a[13] & g[12550];
assign g[28933] = b[13] & g[12550];
assign g[20743] = a[13] & g[12551];
assign g[28934] = b[13] & g[12551];
assign g[20744] = a[13] & g[12552];
assign g[28935] = b[13] & g[12552];
assign g[20745] = a[13] & g[12553];
assign g[28936] = b[13] & g[12553];
assign g[20746] = a[13] & g[12554];
assign g[28937] = b[13] & g[12554];
assign g[20747] = a[13] & g[12555];
assign g[28938] = b[13] & g[12555];
assign g[20748] = a[13] & g[12556];
assign g[28939] = b[13] & g[12556];
assign g[20749] = a[13] & g[12557];
assign g[28940] = b[13] & g[12557];
assign g[20750] = a[13] & g[12558];
assign g[28941] = b[13] & g[12558];
assign g[20751] = a[13] & g[12559];
assign g[28942] = b[13] & g[12559];
assign g[20752] = a[13] & g[12560];
assign g[28943] = b[13] & g[12560];
assign g[20753] = a[13] & g[12561];
assign g[28944] = b[13] & g[12561];
assign g[20754] = a[13] & g[12562];
assign g[28945] = b[13] & g[12562];
assign g[20755] = a[13] & g[12563];
assign g[28946] = b[13] & g[12563];
assign g[20756] = a[13] & g[12564];
assign g[28947] = b[13] & g[12564];
assign g[20757] = a[13] & g[12565];
assign g[28948] = b[13] & g[12565];
assign g[20758] = a[13] & g[12566];
assign g[28949] = b[13] & g[12566];
assign g[20759] = a[13] & g[12567];
assign g[28950] = b[13] & g[12567];
assign g[20760] = a[13] & g[12568];
assign g[28951] = b[13] & g[12568];
assign g[20761] = a[13] & g[12569];
assign g[28952] = b[13] & g[12569];
assign g[20762] = a[13] & g[12570];
assign g[28953] = b[13] & g[12570];
assign g[20763] = a[13] & g[12571];
assign g[28954] = b[13] & g[12571];
assign g[20764] = a[13] & g[12572];
assign g[28955] = b[13] & g[12572];
assign g[20765] = a[13] & g[12573];
assign g[28956] = b[13] & g[12573];
assign g[20766] = a[13] & g[12574];
assign g[28957] = b[13] & g[12574];
assign g[20767] = a[13] & g[12575];
assign g[28958] = b[13] & g[12575];
assign g[20768] = a[13] & g[12576];
assign g[28959] = b[13] & g[12576];
assign g[20769] = a[13] & g[12577];
assign g[28960] = b[13] & g[12577];
assign g[20770] = a[13] & g[12578];
assign g[28961] = b[13] & g[12578];
assign g[20771] = a[13] & g[12579];
assign g[28962] = b[13] & g[12579];
assign g[20772] = a[13] & g[12580];
assign g[28963] = b[13] & g[12580];
assign g[20773] = a[13] & g[12581];
assign g[28964] = b[13] & g[12581];
assign g[20774] = a[13] & g[12582];
assign g[28965] = b[13] & g[12582];
assign g[20775] = a[13] & g[12583];
assign g[28966] = b[13] & g[12583];
assign g[20776] = a[13] & g[12584];
assign g[28967] = b[13] & g[12584];
assign g[20777] = a[13] & g[12585];
assign g[28968] = b[13] & g[12585];
assign g[20778] = a[13] & g[12586];
assign g[28969] = b[13] & g[12586];
assign g[20779] = a[13] & g[12587];
assign g[28970] = b[13] & g[12587];
assign g[20780] = a[13] & g[12588];
assign g[28971] = b[13] & g[12588];
assign g[20781] = a[13] & g[12589];
assign g[28972] = b[13] & g[12589];
assign g[20782] = a[13] & g[12590];
assign g[28973] = b[13] & g[12590];
assign g[20783] = a[13] & g[12591];
assign g[28974] = b[13] & g[12591];
assign g[20784] = a[13] & g[12592];
assign g[28975] = b[13] & g[12592];
assign g[20785] = a[13] & g[12593];
assign g[28976] = b[13] & g[12593];
assign g[20786] = a[13] & g[12594];
assign g[28977] = b[13] & g[12594];
assign g[20787] = a[13] & g[12595];
assign g[28978] = b[13] & g[12595];
assign g[20788] = a[13] & g[12596];
assign g[28979] = b[13] & g[12596];
assign g[20789] = a[13] & g[12597];
assign g[28980] = b[13] & g[12597];
assign g[20790] = a[13] & g[12598];
assign g[28981] = b[13] & g[12598];
assign g[20791] = a[13] & g[12599];
assign g[28982] = b[13] & g[12599];
assign g[20792] = a[13] & g[12600];
assign g[28983] = b[13] & g[12600];
assign g[20793] = a[13] & g[12601];
assign g[28984] = b[13] & g[12601];
assign g[20794] = a[13] & g[12602];
assign g[28985] = b[13] & g[12602];
assign g[20795] = a[13] & g[12603];
assign g[28986] = b[13] & g[12603];
assign g[20796] = a[13] & g[12604];
assign g[28987] = b[13] & g[12604];
assign g[20797] = a[13] & g[12605];
assign g[28988] = b[13] & g[12605];
assign g[20798] = a[13] & g[12606];
assign g[28989] = b[13] & g[12606];
assign g[20799] = a[13] & g[12607];
assign g[28990] = b[13] & g[12607];
assign g[20800] = a[13] & g[12608];
assign g[28991] = b[13] & g[12608];
assign g[20801] = a[13] & g[12609];
assign g[28992] = b[13] & g[12609];
assign g[20802] = a[13] & g[12610];
assign g[28993] = b[13] & g[12610];
assign g[20803] = a[13] & g[12611];
assign g[28994] = b[13] & g[12611];
assign g[20804] = a[13] & g[12612];
assign g[28995] = b[13] & g[12612];
assign g[20805] = a[13] & g[12613];
assign g[28996] = b[13] & g[12613];
assign g[20806] = a[13] & g[12614];
assign g[28997] = b[13] & g[12614];
assign g[20807] = a[13] & g[12615];
assign g[28998] = b[13] & g[12615];
assign g[20808] = a[13] & g[12616];
assign g[28999] = b[13] & g[12616];
assign g[20809] = a[13] & g[12617];
assign g[29000] = b[13] & g[12617];
assign g[20810] = a[13] & g[12618];
assign g[29001] = b[13] & g[12618];
assign g[20811] = a[13] & g[12619];
assign g[29002] = b[13] & g[12619];
assign g[20812] = a[13] & g[12620];
assign g[29003] = b[13] & g[12620];
assign g[20813] = a[13] & g[12621];
assign g[29004] = b[13] & g[12621];
assign g[20814] = a[13] & g[12622];
assign g[29005] = b[13] & g[12622];
assign g[20815] = a[13] & g[12623];
assign g[29006] = b[13] & g[12623];
assign g[20816] = a[13] & g[12624];
assign g[29007] = b[13] & g[12624];
assign g[20817] = a[13] & g[12625];
assign g[29008] = b[13] & g[12625];
assign g[20818] = a[13] & g[12626];
assign g[29009] = b[13] & g[12626];
assign g[20819] = a[13] & g[12627];
assign g[29010] = b[13] & g[12627];
assign g[20820] = a[13] & g[12628];
assign g[29011] = b[13] & g[12628];
assign g[20821] = a[13] & g[12629];
assign g[29012] = b[13] & g[12629];
assign g[20822] = a[13] & g[12630];
assign g[29013] = b[13] & g[12630];
assign g[20823] = a[13] & g[12631];
assign g[29014] = b[13] & g[12631];
assign g[20824] = a[13] & g[12632];
assign g[29015] = b[13] & g[12632];
assign g[20825] = a[13] & g[12633];
assign g[29016] = b[13] & g[12633];
assign g[20826] = a[13] & g[12634];
assign g[29017] = b[13] & g[12634];
assign g[20827] = a[13] & g[12635];
assign g[29018] = b[13] & g[12635];
assign g[20828] = a[13] & g[12636];
assign g[29019] = b[13] & g[12636];
assign g[20829] = a[13] & g[12637];
assign g[29020] = b[13] & g[12637];
assign g[20830] = a[13] & g[12638];
assign g[29021] = b[13] & g[12638];
assign g[20831] = a[13] & g[12639];
assign g[29022] = b[13] & g[12639];
assign g[20832] = a[13] & g[12640];
assign g[29023] = b[13] & g[12640];
assign g[20833] = a[13] & g[12641];
assign g[29024] = b[13] & g[12641];
assign g[20834] = a[13] & g[12642];
assign g[29025] = b[13] & g[12642];
assign g[20835] = a[13] & g[12643];
assign g[29026] = b[13] & g[12643];
assign g[20836] = a[13] & g[12644];
assign g[29027] = b[13] & g[12644];
assign g[20837] = a[13] & g[12645];
assign g[29028] = b[13] & g[12645];
assign g[20838] = a[13] & g[12646];
assign g[29029] = b[13] & g[12646];
assign g[20839] = a[13] & g[12647];
assign g[29030] = b[13] & g[12647];
assign g[20840] = a[13] & g[12648];
assign g[29031] = b[13] & g[12648];
assign g[20841] = a[13] & g[12649];
assign g[29032] = b[13] & g[12649];
assign g[20842] = a[13] & g[12650];
assign g[29033] = b[13] & g[12650];
assign g[20843] = a[13] & g[12651];
assign g[29034] = b[13] & g[12651];
assign g[20844] = a[13] & g[12652];
assign g[29035] = b[13] & g[12652];
assign g[20845] = a[13] & g[12653];
assign g[29036] = b[13] & g[12653];
assign g[20846] = a[13] & g[12654];
assign g[29037] = b[13] & g[12654];
assign g[20847] = a[13] & g[12655];
assign g[29038] = b[13] & g[12655];
assign g[20848] = a[13] & g[12656];
assign g[29039] = b[13] & g[12656];
assign g[20849] = a[13] & g[12657];
assign g[29040] = b[13] & g[12657];
assign g[20850] = a[13] & g[12658];
assign g[29041] = b[13] & g[12658];
assign g[20851] = a[13] & g[12659];
assign g[29042] = b[13] & g[12659];
assign g[20852] = a[13] & g[12660];
assign g[29043] = b[13] & g[12660];
assign g[20853] = a[13] & g[12661];
assign g[29044] = b[13] & g[12661];
assign g[20854] = a[13] & g[12662];
assign g[29045] = b[13] & g[12662];
assign g[20855] = a[13] & g[12663];
assign g[29046] = b[13] & g[12663];
assign g[20856] = a[13] & g[12664];
assign g[29047] = b[13] & g[12664];
assign g[20857] = a[13] & g[12665];
assign g[29048] = b[13] & g[12665];
assign g[20858] = a[13] & g[12666];
assign g[29049] = b[13] & g[12666];
assign g[20859] = a[13] & g[12667];
assign g[29050] = b[13] & g[12667];
assign g[20860] = a[13] & g[12668];
assign g[29051] = b[13] & g[12668];
assign g[20861] = a[13] & g[12669];
assign g[29052] = b[13] & g[12669];
assign g[20862] = a[13] & g[12670];
assign g[29053] = b[13] & g[12670];
assign g[20863] = a[13] & g[12671];
assign g[29054] = b[13] & g[12671];
assign g[20864] = a[13] & g[12672];
assign g[29055] = b[13] & g[12672];
assign g[20865] = a[13] & g[12673];
assign g[29056] = b[13] & g[12673];
assign g[20866] = a[13] & g[12674];
assign g[29057] = b[13] & g[12674];
assign g[20867] = a[13] & g[12675];
assign g[29058] = b[13] & g[12675];
assign g[20868] = a[13] & g[12676];
assign g[29059] = b[13] & g[12676];
assign g[20869] = a[13] & g[12677];
assign g[29060] = b[13] & g[12677];
assign g[20870] = a[13] & g[12678];
assign g[29061] = b[13] & g[12678];
assign g[20871] = a[13] & g[12679];
assign g[29062] = b[13] & g[12679];
assign g[20872] = a[13] & g[12680];
assign g[29063] = b[13] & g[12680];
assign g[20873] = a[13] & g[12681];
assign g[29064] = b[13] & g[12681];
assign g[20874] = a[13] & g[12682];
assign g[29065] = b[13] & g[12682];
assign g[20875] = a[13] & g[12683];
assign g[29066] = b[13] & g[12683];
assign g[20876] = a[13] & g[12684];
assign g[29067] = b[13] & g[12684];
assign g[20877] = a[13] & g[12685];
assign g[29068] = b[13] & g[12685];
assign g[20878] = a[13] & g[12686];
assign g[29069] = b[13] & g[12686];
assign g[20879] = a[13] & g[12687];
assign g[29070] = b[13] & g[12687];
assign g[20880] = a[13] & g[12688];
assign g[29071] = b[13] & g[12688];
assign g[20881] = a[13] & g[12689];
assign g[29072] = b[13] & g[12689];
assign g[20882] = a[13] & g[12690];
assign g[29073] = b[13] & g[12690];
assign g[20883] = a[13] & g[12691];
assign g[29074] = b[13] & g[12691];
assign g[20884] = a[13] & g[12692];
assign g[29075] = b[13] & g[12692];
assign g[20885] = a[13] & g[12693];
assign g[29076] = b[13] & g[12693];
assign g[20886] = a[13] & g[12694];
assign g[29077] = b[13] & g[12694];
assign g[20887] = a[13] & g[12695];
assign g[29078] = b[13] & g[12695];
assign g[20888] = a[13] & g[12696];
assign g[29079] = b[13] & g[12696];
assign g[20889] = a[13] & g[12697];
assign g[29080] = b[13] & g[12697];
assign g[20890] = a[13] & g[12698];
assign g[29081] = b[13] & g[12698];
assign g[20891] = a[13] & g[12699];
assign g[29082] = b[13] & g[12699];
assign g[20892] = a[13] & g[12700];
assign g[29083] = b[13] & g[12700];
assign g[20893] = a[13] & g[12701];
assign g[29084] = b[13] & g[12701];
assign g[20894] = a[13] & g[12702];
assign g[29085] = b[13] & g[12702];
assign g[20895] = a[13] & g[12703];
assign g[29086] = b[13] & g[12703];
assign g[20896] = a[13] & g[12704];
assign g[29087] = b[13] & g[12704];
assign g[20897] = a[13] & g[12705];
assign g[29088] = b[13] & g[12705];
assign g[20898] = a[13] & g[12706];
assign g[29089] = b[13] & g[12706];
assign g[20899] = a[13] & g[12707];
assign g[29090] = b[13] & g[12707];
assign g[20900] = a[13] & g[12708];
assign g[29091] = b[13] & g[12708];
assign g[20901] = a[13] & g[12709];
assign g[29092] = b[13] & g[12709];
assign g[20902] = a[13] & g[12710];
assign g[29093] = b[13] & g[12710];
assign g[20903] = a[13] & g[12711];
assign g[29094] = b[13] & g[12711];
assign g[20904] = a[13] & g[12712];
assign g[29095] = b[13] & g[12712];
assign g[20905] = a[13] & g[12713];
assign g[29096] = b[13] & g[12713];
assign g[20906] = a[13] & g[12714];
assign g[29097] = b[13] & g[12714];
assign g[20907] = a[13] & g[12715];
assign g[29098] = b[13] & g[12715];
assign g[20908] = a[13] & g[12716];
assign g[29099] = b[13] & g[12716];
assign g[20909] = a[13] & g[12717];
assign g[29100] = b[13] & g[12717];
assign g[20910] = a[13] & g[12718];
assign g[29101] = b[13] & g[12718];
assign g[20911] = a[13] & g[12719];
assign g[29102] = b[13] & g[12719];
assign g[20912] = a[13] & g[12720];
assign g[29103] = b[13] & g[12720];
assign g[20913] = a[13] & g[12721];
assign g[29104] = b[13] & g[12721];
assign g[20914] = a[13] & g[12722];
assign g[29105] = b[13] & g[12722];
assign g[20915] = a[13] & g[12723];
assign g[29106] = b[13] & g[12723];
assign g[20916] = a[13] & g[12724];
assign g[29107] = b[13] & g[12724];
assign g[20917] = a[13] & g[12725];
assign g[29108] = b[13] & g[12725];
assign g[20918] = a[13] & g[12726];
assign g[29109] = b[13] & g[12726];
assign g[20919] = a[13] & g[12727];
assign g[29110] = b[13] & g[12727];
assign g[20920] = a[13] & g[12728];
assign g[29111] = b[13] & g[12728];
assign g[20921] = a[13] & g[12729];
assign g[29112] = b[13] & g[12729];
assign g[20922] = a[13] & g[12730];
assign g[29113] = b[13] & g[12730];
assign g[20923] = a[13] & g[12731];
assign g[29114] = b[13] & g[12731];
assign g[20924] = a[13] & g[12732];
assign g[29115] = b[13] & g[12732];
assign g[20925] = a[13] & g[12733];
assign g[29116] = b[13] & g[12733];
assign g[20926] = a[13] & g[12734];
assign g[29117] = b[13] & g[12734];
assign g[20927] = a[13] & g[12735];
assign g[29118] = b[13] & g[12735];
assign g[20928] = a[13] & g[12736];
assign g[29119] = b[13] & g[12736];
assign g[20929] = a[13] & g[12737];
assign g[29120] = b[13] & g[12737];
assign g[20930] = a[13] & g[12738];
assign g[29121] = b[13] & g[12738];
assign g[20931] = a[13] & g[12739];
assign g[29122] = b[13] & g[12739];
assign g[20932] = a[13] & g[12740];
assign g[29123] = b[13] & g[12740];
assign g[20933] = a[13] & g[12741];
assign g[29124] = b[13] & g[12741];
assign g[20934] = a[13] & g[12742];
assign g[29125] = b[13] & g[12742];
assign g[20935] = a[13] & g[12743];
assign g[29126] = b[13] & g[12743];
assign g[20936] = a[13] & g[12744];
assign g[29127] = b[13] & g[12744];
assign g[20937] = a[13] & g[12745];
assign g[29128] = b[13] & g[12745];
assign g[20938] = a[13] & g[12746];
assign g[29129] = b[13] & g[12746];
assign g[20939] = a[13] & g[12747];
assign g[29130] = b[13] & g[12747];
assign g[20940] = a[13] & g[12748];
assign g[29131] = b[13] & g[12748];
assign g[20941] = a[13] & g[12749];
assign g[29132] = b[13] & g[12749];
assign g[20942] = a[13] & g[12750];
assign g[29133] = b[13] & g[12750];
assign g[20943] = a[13] & g[12751];
assign g[29134] = b[13] & g[12751];
assign g[20944] = a[13] & g[12752];
assign g[29135] = b[13] & g[12752];
assign g[20945] = a[13] & g[12753];
assign g[29136] = b[13] & g[12753];
assign g[20946] = a[13] & g[12754];
assign g[29137] = b[13] & g[12754];
assign g[20947] = a[13] & g[12755];
assign g[29138] = b[13] & g[12755];
assign g[20948] = a[13] & g[12756];
assign g[29139] = b[13] & g[12756];
assign g[20949] = a[13] & g[12757];
assign g[29140] = b[13] & g[12757];
assign g[20950] = a[13] & g[12758];
assign g[29141] = b[13] & g[12758];
assign g[20951] = a[13] & g[12759];
assign g[29142] = b[13] & g[12759];
assign g[20952] = a[13] & g[12760];
assign g[29143] = b[13] & g[12760];
assign g[20953] = a[13] & g[12761];
assign g[29144] = b[13] & g[12761];
assign g[20954] = a[13] & g[12762];
assign g[29145] = b[13] & g[12762];
assign g[20955] = a[13] & g[12763];
assign g[29146] = b[13] & g[12763];
assign g[20956] = a[13] & g[12764];
assign g[29147] = b[13] & g[12764];
assign g[20957] = a[13] & g[12765];
assign g[29148] = b[13] & g[12765];
assign g[20958] = a[13] & g[12766];
assign g[29149] = b[13] & g[12766];
assign g[20959] = a[13] & g[12767];
assign g[29150] = b[13] & g[12767];
assign g[20960] = a[13] & g[12768];
assign g[29151] = b[13] & g[12768];
assign g[20961] = a[13] & g[12769];
assign g[29152] = b[13] & g[12769];
assign g[20962] = a[13] & g[12770];
assign g[29153] = b[13] & g[12770];
assign g[20963] = a[13] & g[12771];
assign g[29154] = b[13] & g[12771];
assign g[20964] = a[13] & g[12772];
assign g[29155] = b[13] & g[12772];
assign g[20965] = a[13] & g[12773];
assign g[29156] = b[13] & g[12773];
assign g[20966] = a[13] & g[12774];
assign g[29157] = b[13] & g[12774];
assign g[20967] = a[13] & g[12775];
assign g[29158] = b[13] & g[12775];
assign g[20968] = a[13] & g[12776];
assign g[29159] = b[13] & g[12776];
assign g[20969] = a[13] & g[12777];
assign g[29160] = b[13] & g[12777];
assign g[20970] = a[13] & g[12778];
assign g[29161] = b[13] & g[12778];
assign g[20971] = a[13] & g[12779];
assign g[29162] = b[13] & g[12779];
assign g[20972] = a[13] & g[12780];
assign g[29163] = b[13] & g[12780];
assign g[20973] = a[13] & g[12781];
assign g[29164] = b[13] & g[12781];
assign g[20974] = a[13] & g[12782];
assign g[29165] = b[13] & g[12782];
assign g[20975] = a[13] & g[12783];
assign g[29166] = b[13] & g[12783];
assign g[20976] = a[13] & g[12784];
assign g[29167] = b[13] & g[12784];
assign g[20977] = a[13] & g[12785];
assign g[29168] = b[13] & g[12785];
assign g[20978] = a[13] & g[12786];
assign g[29169] = b[13] & g[12786];
assign g[20979] = a[13] & g[12787];
assign g[29170] = b[13] & g[12787];
assign g[20980] = a[13] & g[12788];
assign g[29171] = b[13] & g[12788];
assign g[20981] = a[13] & g[12789];
assign g[29172] = b[13] & g[12789];
assign g[20982] = a[13] & g[12790];
assign g[29173] = b[13] & g[12790];
assign g[20983] = a[13] & g[12791];
assign g[29174] = b[13] & g[12791];
assign g[20984] = a[13] & g[12792];
assign g[29175] = b[13] & g[12792];
assign g[20985] = a[13] & g[12793];
assign g[29176] = b[13] & g[12793];
assign g[20986] = a[13] & g[12794];
assign g[29177] = b[13] & g[12794];
assign g[20987] = a[13] & g[12795];
assign g[29178] = b[13] & g[12795];
assign g[20988] = a[13] & g[12796];
assign g[29179] = b[13] & g[12796];
assign g[20989] = a[13] & g[12797];
assign g[29180] = b[13] & g[12797];
assign g[20990] = a[13] & g[12798];
assign g[29181] = b[13] & g[12798];
assign g[20991] = a[13] & g[12799];
assign g[29182] = b[13] & g[12799];
assign g[20992] = a[13] & g[12800];
assign g[29183] = b[13] & g[12800];
assign g[20993] = a[13] & g[12801];
assign g[29184] = b[13] & g[12801];
assign g[20994] = a[13] & g[12802];
assign g[29185] = b[13] & g[12802];
assign g[20995] = a[13] & g[12803];
assign g[29186] = b[13] & g[12803];
assign g[20996] = a[13] & g[12804];
assign g[29187] = b[13] & g[12804];
assign g[20997] = a[13] & g[12805];
assign g[29188] = b[13] & g[12805];
assign g[20998] = a[13] & g[12806];
assign g[29189] = b[13] & g[12806];
assign g[20999] = a[13] & g[12807];
assign g[29190] = b[13] & g[12807];
assign g[21000] = a[13] & g[12808];
assign g[29191] = b[13] & g[12808];
assign g[21001] = a[13] & g[12809];
assign g[29192] = b[13] & g[12809];
assign g[21002] = a[13] & g[12810];
assign g[29193] = b[13] & g[12810];
assign g[21003] = a[13] & g[12811];
assign g[29194] = b[13] & g[12811];
assign g[21004] = a[13] & g[12812];
assign g[29195] = b[13] & g[12812];
assign g[21005] = a[13] & g[12813];
assign g[29196] = b[13] & g[12813];
assign g[21006] = a[13] & g[12814];
assign g[29197] = b[13] & g[12814];
assign g[21007] = a[13] & g[12815];
assign g[29198] = b[13] & g[12815];
assign g[21008] = a[13] & g[12816];
assign g[29199] = b[13] & g[12816];
assign g[21009] = a[13] & g[12817];
assign g[29200] = b[13] & g[12817];
assign g[21010] = a[13] & g[12818];
assign g[29201] = b[13] & g[12818];
assign g[21011] = a[13] & g[12819];
assign g[29202] = b[13] & g[12819];
assign g[21012] = a[13] & g[12820];
assign g[29203] = b[13] & g[12820];
assign g[21013] = a[13] & g[12821];
assign g[29204] = b[13] & g[12821];
assign g[21014] = a[13] & g[12822];
assign g[29205] = b[13] & g[12822];
assign g[21015] = a[13] & g[12823];
assign g[29206] = b[13] & g[12823];
assign g[21016] = a[13] & g[12824];
assign g[29207] = b[13] & g[12824];
assign g[21017] = a[13] & g[12825];
assign g[29208] = b[13] & g[12825];
assign g[21018] = a[13] & g[12826];
assign g[29209] = b[13] & g[12826];
assign g[21019] = a[13] & g[12827];
assign g[29210] = b[13] & g[12827];
assign g[21020] = a[13] & g[12828];
assign g[29211] = b[13] & g[12828];
assign g[21021] = a[13] & g[12829];
assign g[29212] = b[13] & g[12829];
assign g[21022] = a[13] & g[12830];
assign g[29213] = b[13] & g[12830];
assign g[21023] = a[13] & g[12831];
assign g[29214] = b[13] & g[12831];
assign g[21024] = a[13] & g[12832];
assign g[29215] = b[13] & g[12832];
assign g[21025] = a[13] & g[12833];
assign g[29216] = b[13] & g[12833];
assign g[21026] = a[13] & g[12834];
assign g[29217] = b[13] & g[12834];
assign g[21027] = a[13] & g[12835];
assign g[29218] = b[13] & g[12835];
assign g[21028] = a[13] & g[12836];
assign g[29219] = b[13] & g[12836];
assign g[21029] = a[13] & g[12837];
assign g[29220] = b[13] & g[12837];
assign g[21030] = a[13] & g[12838];
assign g[29221] = b[13] & g[12838];
assign g[21031] = a[13] & g[12839];
assign g[29222] = b[13] & g[12839];
assign g[21032] = a[13] & g[12840];
assign g[29223] = b[13] & g[12840];
assign g[21033] = a[13] & g[12841];
assign g[29224] = b[13] & g[12841];
assign g[21034] = a[13] & g[12842];
assign g[29225] = b[13] & g[12842];
assign g[21035] = a[13] & g[12843];
assign g[29226] = b[13] & g[12843];
assign g[21036] = a[13] & g[12844];
assign g[29227] = b[13] & g[12844];
assign g[21037] = a[13] & g[12845];
assign g[29228] = b[13] & g[12845];
assign g[21038] = a[13] & g[12846];
assign g[29229] = b[13] & g[12846];
assign g[21039] = a[13] & g[12847];
assign g[29230] = b[13] & g[12847];
assign g[21040] = a[13] & g[12848];
assign g[29231] = b[13] & g[12848];
assign g[21041] = a[13] & g[12849];
assign g[29232] = b[13] & g[12849];
assign g[21042] = a[13] & g[12850];
assign g[29233] = b[13] & g[12850];
assign g[21043] = a[13] & g[12851];
assign g[29234] = b[13] & g[12851];
assign g[21044] = a[13] & g[12852];
assign g[29235] = b[13] & g[12852];
assign g[21045] = a[13] & g[12853];
assign g[29236] = b[13] & g[12853];
assign g[21046] = a[13] & g[12854];
assign g[29237] = b[13] & g[12854];
assign g[21047] = a[13] & g[12855];
assign g[29238] = b[13] & g[12855];
assign g[21048] = a[13] & g[12856];
assign g[29239] = b[13] & g[12856];
assign g[21049] = a[13] & g[12857];
assign g[29240] = b[13] & g[12857];
assign g[21050] = a[13] & g[12858];
assign g[29241] = b[13] & g[12858];
assign g[21051] = a[13] & g[12859];
assign g[29242] = b[13] & g[12859];
assign g[21052] = a[13] & g[12860];
assign g[29243] = b[13] & g[12860];
assign g[21053] = a[13] & g[12861];
assign g[29244] = b[13] & g[12861];
assign g[21054] = a[13] & g[12862];
assign g[29245] = b[13] & g[12862];
assign g[21055] = a[13] & g[12863];
assign g[29246] = b[13] & g[12863];
assign g[21056] = a[13] & g[12864];
assign g[29247] = b[13] & g[12864];
assign g[21057] = a[13] & g[12865];
assign g[29248] = b[13] & g[12865];
assign g[21058] = a[13] & g[12866];
assign g[29249] = b[13] & g[12866];
assign g[21059] = a[13] & g[12867];
assign g[29250] = b[13] & g[12867];
assign g[21060] = a[13] & g[12868];
assign g[29251] = b[13] & g[12868];
assign g[21061] = a[13] & g[12869];
assign g[29252] = b[13] & g[12869];
assign g[21062] = a[13] & g[12870];
assign g[29253] = b[13] & g[12870];
assign g[21063] = a[13] & g[12871];
assign g[29254] = b[13] & g[12871];
assign g[21064] = a[13] & g[12872];
assign g[29255] = b[13] & g[12872];
assign g[21065] = a[13] & g[12873];
assign g[29256] = b[13] & g[12873];
assign g[21066] = a[13] & g[12874];
assign g[29257] = b[13] & g[12874];
assign g[21067] = a[13] & g[12875];
assign g[29258] = b[13] & g[12875];
assign g[21068] = a[13] & g[12876];
assign g[29259] = b[13] & g[12876];
assign g[21069] = a[13] & g[12877];
assign g[29260] = b[13] & g[12877];
assign g[21070] = a[13] & g[12878];
assign g[29261] = b[13] & g[12878];
assign g[21071] = a[13] & g[12879];
assign g[29262] = b[13] & g[12879];
assign g[21072] = a[13] & g[12880];
assign g[29263] = b[13] & g[12880];
assign g[21073] = a[13] & g[12881];
assign g[29264] = b[13] & g[12881];
assign g[21074] = a[13] & g[12882];
assign g[29265] = b[13] & g[12882];
assign g[21075] = a[13] & g[12883];
assign g[29266] = b[13] & g[12883];
assign g[21076] = a[13] & g[12884];
assign g[29267] = b[13] & g[12884];
assign g[21077] = a[13] & g[12885];
assign g[29268] = b[13] & g[12885];
assign g[21078] = a[13] & g[12886];
assign g[29269] = b[13] & g[12886];
assign g[21079] = a[13] & g[12887];
assign g[29270] = b[13] & g[12887];
assign g[21080] = a[13] & g[12888];
assign g[29271] = b[13] & g[12888];
assign g[21081] = a[13] & g[12889];
assign g[29272] = b[13] & g[12889];
assign g[21082] = a[13] & g[12890];
assign g[29273] = b[13] & g[12890];
assign g[21083] = a[13] & g[12891];
assign g[29274] = b[13] & g[12891];
assign g[21084] = a[13] & g[12892];
assign g[29275] = b[13] & g[12892];
assign g[21085] = a[13] & g[12893];
assign g[29276] = b[13] & g[12893];
assign g[21086] = a[13] & g[12894];
assign g[29277] = b[13] & g[12894];
assign g[21087] = a[13] & g[12895];
assign g[29278] = b[13] & g[12895];
assign g[21088] = a[13] & g[12896];
assign g[29279] = b[13] & g[12896];
assign g[21089] = a[13] & g[12897];
assign g[29280] = b[13] & g[12897];
assign g[21090] = a[13] & g[12898];
assign g[29281] = b[13] & g[12898];
assign g[21091] = a[13] & g[12899];
assign g[29282] = b[13] & g[12899];
assign g[21092] = a[13] & g[12900];
assign g[29283] = b[13] & g[12900];
assign g[21093] = a[13] & g[12901];
assign g[29284] = b[13] & g[12901];
assign g[21094] = a[13] & g[12902];
assign g[29285] = b[13] & g[12902];
assign g[21095] = a[13] & g[12903];
assign g[29286] = b[13] & g[12903];
assign g[21096] = a[13] & g[12904];
assign g[29287] = b[13] & g[12904];
assign g[21097] = a[13] & g[12905];
assign g[29288] = b[13] & g[12905];
assign g[21098] = a[13] & g[12906];
assign g[29289] = b[13] & g[12906];
assign g[21099] = a[13] & g[12907];
assign g[29290] = b[13] & g[12907];
assign g[21100] = a[13] & g[12908];
assign g[29291] = b[13] & g[12908];
assign g[21101] = a[13] & g[12909];
assign g[29292] = b[13] & g[12909];
assign g[21102] = a[13] & g[12910];
assign g[29293] = b[13] & g[12910];
assign g[21103] = a[13] & g[12911];
assign g[29294] = b[13] & g[12911];
assign g[21104] = a[13] & g[12912];
assign g[29295] = b[13] & g[12912];
assign g[21105] = a[13] & g[12913];
assign g[29296] = b[13] & g[12913];
assign g[21106] = a[13] & g[12914];
assign g[29297] = b[13] & g[12914];
assign g[21107] = a[13] & g[12915];
assign g[29298] = b[13] & g[12915];
assign g[21108] = a[13] & g[12916];
assign g[29299] = b[13] & g[12916];
assign g[21109] = a[13] & g[12917];
assign g[29300] = b[13] & g[12917];
assign g[21110] = a[13] & g[12918];
assign g[29301] = b[13] & g[12918];
assign g[21111] = a[13] & g[12919];
assign g[29302] = b[13] & g[12919];
assign g[21112] = a[13] & g[12920];
assign g[29303] = b[13] & g[12920];
assign g[21113] = a[13] & g[12921];
assign g[29304] = b[13] & g[12921];
assign g[21114] = a[13] & g[12922];
assign g[29305] = b[13] & g[12922];
assign g[21115] = a[13] & g[12923];
assign g[29306] = b[13] & g[12923];
assign g[21116] = a[13] & g[12924];
assign g[29307] = b[13] & g[12924];
assign g[21117] = a[13] & g[12925];
assign g[29308] = b[13] & g[12925];
assign g[21118] = a[13] & g[12926];
assign g[29309] = b[13] & g[12926];
assign g[21119] = a[13] & g[12927];
assign g[29310] = b[13] & g[12927];
assign g[21120] = a[13] & g[12928];
assign g[29311] = b[13] & g[12928];
assign g[21121] = a[13] & g[12929];
assign g[29312] = b[13] & g[12929];
assign g[21122] = a[13] & g[12930];
assign g[29313] = b[13] & g[12930];
assign g[21123] = a[13] & g[12931];
assign g[29314] = b[13] & g[12931];
assign g[21124] = a[13] & g[12932];
assign g[29315] = b[13] & g[12932];
assign g[21125] = a[13] & g[12933];
assign g[29316] = b[13] & g[12933];
assign g[21126] = a[13] & g[12934];
assign g[29317] = b[13] & g[12934];
assign g[21127] = a[13] & g[12935];
assign g[29318] = b[13] & g[12935];
assign g[21128] = a[13] & g[12936];
assign g[29319] = b[13] & g[12936];
assign g[21129] = a[13] & g[12937];
assign g[29320] = b[13] & g[12937];
assign g[21130] = a[13] & g[12938];
assign g[29321] = b[13] & g[12938];
assign g[21131] = a[13] & g[12939];
assign g[29322] = b[13] & g[12939];
assign g[21132] = a[13] & g[12940];
assign g[29323] = b[13] & g[12940];
assign g[21133] = a[13] & g[12941];
assign g[29324] = b[13] & g[12941];
assign g[21134] = a[13] & g[12942];
assign g[29325] = b[13] & g[12942];
assign g[21135] = a[13] & g[12943];
assign g[29326] = b[13] & g[12943];
assign g[21136] = a[13] & g[12944];
assign g[29327] = b[13] & g[12944];
assign g[21137] = a[13] & g[12945];
assign g[29328] = b[13] & g[12945];
assign g[21138] = a[13] & g[12946];
assign g[29329] = b[13] & g[12946];
assign g[21139] = a[13] & g[12947];
assign g[29330] = b[13] & g[12947];
assign g[21140] = a[13] & g[12948];
assign g[29331] = b[13] & g[12948];
assign g[21141] = a[13] & g[12949];
assign g[29332] = b[13] & g[12949];
assign g[21142] = a[13] & g[12950];
assign g[29333] = b[13] & g[12950];
assign g[21143] = a[13] & g[12951];
assign g[29334] = b[13] & g[12951];
assign g[21144] = a[13] & g[12952];
assign g[29335] = b[13] & g[12952];
assign g[21145] = a[13] & g[12953];
assign g[29336] = b[13] & g[12953];
assign g[21146] = a[13] & g[12954];
assign g[29337] = b[13] & g[12954];
assign g[21147] = a[13] & g[12955];
assign g[29338] = b[13] & g[12955];
assign g[21148] = a[13] & g[12956];
assign g[29339] = b[13] & g[12956];
assign g[21149] = a[13] & g[12957];
assign g[29340] = b[13] & g[12957];
assign g[21150] = a[13] & g[12958];
assign g[29341] = b[13] & g[12958];
assign g[21151] = a[13] & g[12959];
assign g[29342] = b[13] & g[12959];
assign g[21152] = a[13] & g[12960];
assign g[29343] = b[13] & g[12960];
assign g[21153] = a[13] & g[12961];
assign g[29344] = b[13] & g[12961];
assign g[21154] = a[13] & g[12962];
assign g[29345] = b[13] & g[12962];
assign g[21155] = a[13] & g[12963];
assign g[29346] = b[13] & g[12963];
assign g[21156] = a[13] & g[12964];
assign g[29347] = b[13] & g[12964];
assign g[21157] = a[13] & g[12965];
assign g[29348] = b[13] & g[12965];
assign g[21158] = a[13] & g[12966];
assign g[29349] = b[13] & g[12966];
assign g[21159] = a[13] & g[12967];
assign g[29350] = b[13] & g[12967];
assign g[21160] = a[13] & g[12968];
assign g[29351] = b[13] & g[12968];
assign g[21161] = a[13] & g[12969];
assign g[29352] = b[13] & g[12969];
assign g[21162] = a[13] & g[12970];
assign g[29353] = b[13] & g[12970];
assign g[21163] = a[13] & g[12971];
assign g[29354] = b[13] & g[12971];
assign g[21164] = a[13] & g[12972];
assign g[29355] = b[13] & g[12972];
assign g[21165] = a[13] & g[12973];
assign g[29356] = b[13] & g[12973];
assign g[21166] = a[13] & g[12974];
assign g[29357] = b[13] & g[12974];
assign g[21167] = a[13] & g[12975];
assign g[29358] = b[13] & g[12975];
assign g[21168] = a[13] & g[12976];
assign g[29359] = b[13] & g[12976];
assign g[21169] = a[13] & g[12977];
assign g[29360] = b[13] & g[12977];
assign g[21170] = a[13] & g[12978];
assign g[29361] = b[13] & g[12978];
assign g[21171] = a[13] & g[12979];
assign g[29362] = b[13] & g[12979];
assign g[21172] = a[13] & g[12980];
assign g[29363] = b[13] & g[12980];
assign g[21173] = a[13] & g[12981];
assign g[29364] = b[13] & g[12981];
assign g[21174] = a[13] & g[12982];
assign g[29365] = b[13] & g[12982];
assign g[21175] = a[13] & g[12983];
assign g[29366] = b[13] & g[12983];
assign g[21176] = a[13] & g[12984];
assign g[29367] = b[13] & g[12984];
assign g[21177] = a[13] & g[12985];
assign g[29368] = b[13] & g[12985];
assign g[21178] = a[13] & g[12986];
assign g[29369] = b[13] & g[12986];
assign g[21179] = a[13] & g[12987];
assign g[29370] = b[13] & g[12987];
assign g[21180] = a[13] & g[12988];
assign g[29371] = b[13] & g[12988];
assign g[21181] = a[13] & g[12989];
assign g[29372] = b[13] & g[12989];
assign g[21182] = a[13] & g[12990];
assign g[29373] = b[13] & g[12990];
assign g[21183] = a[13] & g[12991];
assign g[29374] = b[13] & g[12991];
assign g[21184] = a[13] & g[12992];
assign g[29375] = b[13] & g[12992];
assign g[21185] = a[13] & g[12993];
assign g[29376] = b[13] & g[12993];
assign g[21186] = a[13] & g[12994];
assign g[29377] = b[13] & g[12994];
assign g[21187] = a[13] & g[12995];
assign g[29378] = b[13] & g[12995];
assign g[21188] = a[13] & g[12996];
assign g[29379] = b[13] & g[12996];
assign g[21189] = a[13] & g[12997];
assign g[29380] = b[13] & g[12997];
assign g[21190] = a[13] & g[12998];
assign g[29381] = b[13] & g[12998];
assign g[21191] = a[13] & g[12999];
assign g[29382] = b[13] & g[12999];
assign g[21192] = a[13] & g[13000];
assign g[29383] = b[13] & g[13000];
assign g[21193] = a[13] & g[13001];
assign g[29384] = b[13] & g[13001];
assign g[21194] = a[13] & g[13002];
assign g[29385] = b[13] & g[13002];
assign g[21195] = a[13] & g[13003];
assign g[29386] = b[13] & g[13003];
assign g[21196] = a[13] & g[13004];
assign g[29387] = b[13] & g[13004];
assign g[21197] = a[13] & g[13005];
assign g[29388] = b[13] & g[13005];
assign g[21198] = a[13] & g[13006];
assign g[29389] = b[13] & g[13006];
assign g[21199] = a[13] & g[13007];
assign g[29390] = b[13] & g[13007];
assign g[21200] = a[13] & g[13008];
assign g[29391] = b[13] & g[13008];
assign g[21201] = a[13] & g[13009];
assign g[29392] = b[13] & g[13009];
assign g[21202] = a[13] & g[13010];
assign g[29393] = b[13] & g[13010];
assign g[21203] = a[13] & g[13011];
assign g[29394] = b[13] & g[13011];
assign g[21204] = a[13] & g[13012];
assign g[29395] = b[13] & g[13012];
assign g[21205] = a[13] & g[13013];
assign g[29396] = b[13] & g[13013];
assign g[21206] = a[13] & g[13014];
assign g[29397] = b[13] & g[13014];
assign g[21207] = a[13] & g[13015];
assign g[29398] = b[13] & g[13015];
assign g[21208] = a[13] & g[13016];
assign g[29399] = b[13] & g[13016];
assign g[21209] = a[13] & g[13017];
assign g[29400] = b[13] & g[13017];
assign g[21210] = a[13] & g[13018];
assign g[29401] = b[13] & g[13018];
assign g[21211] = a[13] & g[13019];
assign g[29402] = b[13] & g[13019];
assign g[21212] = a[13] & g[13020];
assign g[29403] = b[13] & g[13020];
assign g[21213] = a[13] & g[13021];
assign g[29404] = b[13] & g[13021];
assign g[21214] = a[13] & g[13022];
assign g[29405] = b[13] & g[13022];
assign g[21215] = a[13] & g[13023];
assign g[29406] = b[13] & g[13023];
assign g[21216] = a[13] & g[13024];
assign g[29407] = b[13] & g[13024];
assign g[21217] = a[13] & g[13025];
assign g[29408] = b[13] & g[13025];
assign g[21218] = a[13] & g[13026];
assign g[29409] = b[13] & g[13026];
assign g[21219] = a[13] & g[13027];
assign g[29410] = b[13] & g[13027];
assign g[21220] = a[13] & g[13028];
assign g[29411] = b[13] & g[13028];
assign g[21221] = a[13] & g[13029];
assign g[29412] = b[13] & g[13029];
assign g[21222] = a[13] & g[13030];
assign g[29413] = b[13] & g[13030];
assign g[21223] = a[13] & g[13031];
assign g[29414] = b[13] & g[13031];
assign g[21224] = a[13] & g[13032];
assign g[29415] = b[13] & g[13032];
assign g[21225] = a[13] & g[13033];
assign g[29416] = b[13] & g[13033];
assign g[21226] = a[13] & g[13034];
assign g[29417] = b[13] & g[13034];
assign g[21227] = a[13] & g[13035];
assign g[29418] = b[13] & g[13035];
assign g[21228] = a[13] & g[13036];
assign g[29419] = b[13] & g[13036];
assign g[21229] = a[13] & g[13037];
assign g[29420] = b[13] & g[13037];
assign g[21230] = a[13] & g[13038];
assign g[29421] = b[13] & g[13038];
assign g[21231] = a[13] & g[13039];
assign g[29422] = b[13] & g[13039];
assign g[21232] = a[13] & g[13040];
assign g[29423] = b[13] & g[13040];
assign g[21233] = a[13] & g[13041];
assign g[29424] = b[13] & g[13041];
assign g[21234] = a[13] & g[13042];
assign g[29425] = b[13] & g[13042];
assign g[21235] = a[13] & g[13043];
assign g[29426] = b[13] & g[13043];
assign g[21236] = a[13] & g[13044];
assign g[29427] = b[13] & g[13044];
assign g[21237] = a[13] & g[13045];
assign g[29428] = b[13] & g[13045];
assign g[21238] = a[13] & g[13046];
assign g[29429] = b[13] & g[13046];
assign g[21239] = a[13] & g[13047];
assign g[29430] = b[13] & g[13047];
assign g[21240] = a[13] & g[13048];
assign g[29431] = b[13] & g[13048];
assign g[21241] = a[13] & g[13049];
assign g[29432] = b[13] & g[13049];
assign g[21242] = a[13] & g[13050];
assign g[29433] = b[13] & g[13050];
assign g[21243] = a[13] & g[13051];
assign g[29434] = b[13] & g[13051];
assign g[21244] = a[13] & g[13052];
assign g[29435] = b[13] & g[13052];
assign g[21245] = a[13] & g[13053];
assign g[29436] = b[13] & g[13053];
assign g[21246] = a[13] & g[13054];
assign g[29437] = b[13] & g[13054];
assign g[21247] = a[13] & g[13055];
assign g[29438] = b[13] & g[13055];
assign g[21248] = a[13] & g[13056];
assign g[29439] = b[13] & g[13056];
assign g[21249] = a[13] & g[13057];
assign g[29440] = b[13] & g[13057];
assign g[21250] = a[13] & g[13058];
assign g[29441] = b[13] & g[13058];
assign g[21251] = a[13] & g[13059];
assign g[29442] = b[13] & g[13059];
assign g[21252] = a[13] & g[13060];
assign g[29443] = b[13] & g[13060];
assign g[21253] = a[13] & g[13061];
assign g[29444] = b[13] & g[13061];
assign g[21254] = a[13] & g[13062];
assign g[29445] = b[13] & g[13062];
assign g[21255] = a[13] & g[13063];
assign g[29446] = b[13] & g[13063];
assign g[21256] = a[13] & g[13064];
assign g[29447] = b[13] & g[13064];
assign g[21257] = a[13] & g[13065];
assign g[29448] = b[13] & g[13065];
assign g[21258] = a[13] & g[13066];
assign g[29449] = b[13] & g[13066];
assign g[21259] = a[13] & g[13067];
assign g[29450] = b[13] & g[13067];
assign g[21260] = a[13] & g[13068];
assign g[29451] = b[13] & g[13068];
assign g[21261] = a[13] & g[13069];
assign g[29452] = b[13] & g[13069];
assign g[21262] = a[13] & g[13070];
assign g[29453] = b[13] & g[13070];
assign g[21263] = a[13] & g[13071];
assign g[29454] = b[13] & g[13071];
assign g[21264] = a[13] & g[13072];
assign g[29455] = b[13] & g[13072];
assign g[21265] = a[13] & g[13073];
assign g[29456] = b[13] & g[13073];
assign g[21266] = a[13] & g[13074];
assign g[29457] = b[13] & g[13074];
assign g[21267] = a[13] & g[13075];
assign g[29458] = b[13] & g[13075];
assign g[21268] = a[13] & g[13076];
assign g[29459] = b[13] & g[13076];
assign g[21269] = a[13] & g[13077];
assign g[29460] = b[13] & g[13077];
assign g[21270] = a[13] & g[13078];
assign g[29461] = b[13] & g[13078];
assign g[21271] = a[13] & g[13079];
assign g[29462] = b[13] & g[13079];
assign g[21272] = a[13] & g[13080];
assign g[29463] = b[13] & g[13080];
assign g[21273] = a[13] & g[13081];
assign g[29464] = b[13] & g[13081];
assign g[21274] = a[13] & g[13082];
assign g[29465] = b[13] & g[13082];
assign g[21275] = a[13] & g[13083];
assign g[29466] = b[13] & g[13083];
assign g[21276] = a[13] & g[13084];
assign g[29467] = b[13] & g[13084];
assign g[21277] = a[13] & g[13085];
assign g[29468] = b[13] & g[13085];
assign g[21278] = a[13] & g[13086];
assign g[29469] = b[13] & g[13086];
assign g[21279] = a[13] & g[13087];
assign g[29470] = b[13] & g[13087];
assign g[21280] = a[13] & g[13088];
assign g[29471] = b[13] & g[13088];
assign g[21281] = a[13] & g[13089];
assign g[29472] = b[13] & g[13089];
assign g[21282] = a[13] & g[13090];
assign g[29473] = b[13] & g[13090];
assign g[21283] = a[13] & g[13091];
assign g[29474] = b[13] & g[13091];
assign g[21284] = a[13] & g[13092];
assign g[29475] = b[13] & g[13092];
assign g[21285] = a[13] & g[13093];
assign g[29476] = b[13] & g[13093];
assign g[21286] = a[13] & g[13094];
assign g[29477] = b[13] & g[13094];
assign g[21287] = a[13] & g[13095];
assign g[29478] = b[13] & g[13095];
assign g[21288] = a[13] & g[13096];
assign g[29479] = b[13] & g[13096];
assign g[21289] = a[13] & g[13097];
assign g[29480] = b[13] & g[13097];
assign g[21290] = a[13] & g[13098];
assign g[29481] = b[13] & g[13098];
assign g[21291] = a[13] & g[13099];
assign g[29482] = b[13] & g[13099];
assign g[21292] = a[13] & g[13100];
assign g[29483] = b[13] & g[13100];
assign g[21293] = a[13] & g[13101];
assign g[29484] = b[13] & g[13101];
assign g[21294] = a[13] & g[13102];
assign g[29485] = b[13] & g[13102];
assign g[21295] = a[13] & g[13103];
assign g[29486] = b[13] & g[13103];
assign g[21296] = a[13] & g[13104];
assign g[29487] = b[13] & g[13104];
assign g[21297] = a[13] & g[13105];
assign g[29488] = b[13] & g[13105];
assign g[21298] = a[13] & g[13106];
assign g[29489] = b[13] & g[13106];
assign g[21299] = a[13] & g[13107];
assign g[29490] = b[13] & g[13107];
assign g[21300] = a[13] & g[13108];
assign g[29491] = b[13] & g[13108];
assign g[21301] = a[13] & g[13109];
assign g[29492] = b[13] & g[13109];
assign g[21302] = a[13] & g[13110];
assign g[29493] = b[13] & g[13110];
assign g[21303] = a[13] & g[13111];
assign g[29494] = b[13] & g[13111];
assign g[21304] = a[13] & g[13112];
assign g[29495] = b[13] & g[13112];
assign g[21305] = a[13] & g[13113];
assign g[29496] = b[13] & g[13113];
assign g[21306] = a[13] & g[13114];
assign g[29497] = b[13] & g[13114];
assign g[21307] = a[13] & g[13115];
assign g[29498] = b[13] & g[13115];
assign g[21308] = a[13] & g[13116];
assign g[29499] = b[13] & g[13116];
assign g[21309] = a[13] & g[13117];
assign g[29500] = b[13] & g[13117];
assign g[21310] = a[13] & g[13118];
assign g[29501] = b[13] & g[13118];
assign g[21311] = a[13] & g[13119];
assign g[29502] = b[13] & g[13119];
assign g[21312] = a[13] & g[13120];
assign g[29503] = b[13] & g[13120];
assign g[21313] = a[13] & g[13121];
assign g[29504] = b[13] & g[13121];
assign g[21314] = a[13] & g[13122];
assign g[29505] = b[13] & g[13122];
assign g[21315] = a[13] & g[13123];
assign g[29506] = b[13] & g[13123];
assign g[21316] = a[13] & g[13124];
assign g[29507] = b[13] & g[13124];
assign g[21317] = a[13] & g[13125];
assign g[29508] = b[13] & g[13125];
assign g[21318] = a[13] & g[13126];
assign g[29509] = b[13] & g[13126];
assign g[21319] = a[13] & g[13127];
assign g[29510] = b[13] & g[13127];
assign g[21320] = a[13] & g[13128];
assign g[29511] = b[13] & g[13128];
assign g[21321] = a[13] & g[13129];
assign g[29512] = b[13] & g[13129];
assign g[21322] = a[13] & g[13130];
assign g[29513] = b[13] & g[13130];
assign g[21323] = a[13] & g[13131];
assign g[29514] = b[13] & g[13131];
assign g[21324] = a[13] & g[13132];
assign g[29515] = b[13] & g[13132];
assign g[21325] = a[13] & g[13133];
assign g[29516] = b[13] & g[13133];
assign g[21326] = a[13] & g[13134];
assign g[29517] = b[13] & g[13134];
assign g[21327] = a[13] & g[13135];
assign g[29518] = b[13] & g[13135];
assign g[21328] = a[13] & g[13136];
assign g[29519] = b[13] & g[13136];
assign g[21329] = a[13] & g[13137];
assign g[29520] = b[13] & g[13137];
assign g[21330] = a[13] & g[13138];
assign g[29521] = b[13] & g[13138];
assign g[21331] = a[13] & g[13139];
assign g[29522] = b[13] & g[13139];
assign g[21332] = a[13] & g[13140];
assign g[29523] = b[13] & g[13140];
assign g[21333] = a[13] & g[13141];
assign g[29524] = b[13] & g[13141];
assign g[21334] = a[13] & g[13142];
assign g[29525] = b[13] & g[13142];
assign g[21335] = a[13] & g[13143];
assign g[29526] = b[13] & g[13143];
assign g[21336] = a[13] & g[13144];
assign g[29527] = b[13] & g[13144];
assign g[21337] = a[13] & g[13145];
assign g[29528] = b[13] & g[13145];
assign g[21338] = a[13] & g[13146];
assign g[29529] = b[13] & g[13146];
assign g[21339] = a[13] & g[13147];
assign g[29530] = b[13] & g[13147];
assign g[21340] = a[13] & g[13148];
assign g[29531] = b[13] & g[13148];
assign g[21341] = a[13] & g[13149];
assign g[29532] = b[13] & g[13149];
assign g[21342] = a[13] & g[13150];
assign g[29533] = b[13] & g[13150];
assign g[21343] = a[13] & g[13151];
assign g[29534] = b[13] & g[13151];
assign g[21344] = a[13] & g[13152];
assign g[29535] = b[13] & g[13152];
assign g[21345] = a[13] & g[13153];
assign g[29536] = b[13] & g[13153];
assign g[21346] = a[13] & g[13154];
assign g[29537] = b[13] & g[13154];
assign g[21347] = a[13] & g[13155];
assign g[29538] = b[13] & g[13155];
assign g[21348] = a[13] & g[13156];
assign g[29539] = b[13] & g[13156];
assign g[21349] = a[13] & g[13157];
assign g[29540] = b[13] & g[13157];
assign g[21350] = a[13] & g[13158];
assign g[29541] = b[13] & g[13158];
assign g[21351] = a[13] & g[13159];
assign g[29542] = b[13] & g[13159];
assign g[21352] = a[13] & g[13160];
assign g[29543] = b[13] & g[13160];
assign g[21353] = a[13] & g[13161];
assign g[29544] = b[13] & g[13161];
assign g[21354] = a[13] & g[13162];
assign g[29545] = b[13] & g[13162];
assign g[21355] = a[13] & g[13163];
assign g[29546] = b[13] & g[13163];
assign g[21356] = a[13] & g[13164];
assign g[29547] = b[13] & g[13164];
assign g[21357] = a[13] & g[13165];
assign g[29548] = b[13] & g[13165];
assign g[21358] = a[13] & g[13166];
assign g[29549] = b[13] & g[13166];
assign g[21359] = a[13] & g[13167];
assign g[29550] = b[13] & g[13167];
assign g[21360] = a[13] & g[13168];
assign g[29551] = b[13] & g[13168];
assign g[21361] = a[13] & g[13169];
assign g[29552] = b[13] & g[13169];
assign g[21362] = a[13] & g[13170];
assign g[29553] = b[13] & g[13170];
assign g[21363] = a[13] & g[13171];
assign g[29554] = b[13] & g[13171];
assign g[21364] = a[13] & g[13172];
assign g[29555] = b[13] & g[13172];
assign g[21365] = a[13] & g[13173];
assign g[29556] = b[13] & g[13173];
assign g[21366] = a[13] & g[13174];
assign g[29557] = b[13] & g[13174];
assign g[21367] = a[13] & g[13175];
assign g[29558] = b[13] & g[13175];
assign g[21368] = a[13] & g[13176];
assign g[29559] = b[13] & g[13176];
assign g[21369] = a[13] & g[13177];
assign g[29560] = b[13] & g[13177];
assign g[21370] = a[13] & g[13178];
assign g[29561] = b[13] & g[13178];
assign g[21371] = a[13] & g[13179];
assign g[29562] = b[13] & g[13179];
assign g[21372] = a[13] & g[13180];
assign g[29563] = b[13] & g[13180];
assign g[21373] = a[13] & g[13181];
assign g[29564] = b[13] & g[13181];
assign g[21374] = a[13] & g[13182];
assign g[29565] = b[13] & g[13182];
assign g[21375] = a[13] & g[13183];
assign g[29566] = b[13] & g[13183];
assign g[21376] = a[13] & g[13184];
assign g[29567] = b[13] & g[13184];
assign g[21377] = a[13] & g[13185];
assign g[29568] = b[13] & g[13185];
assign g[21378] = a[13] & g[13186];
assign g[29569] = b[13] & g[13186];
assign g[21379] = a[13] & g[13187];
assign g[29570] = b[13] & g[13187];
assign g[21380] = a[13] & g[13188];
assign g[29571] = b[13] & g[13188];
assign g[21381] = a[13] & g[13189];
assign g[29572] = b[13] & g[13189];
assign g[21382] = a[13] & g[13190];
assign g[29573] = b[13] & g[13190];
assign g[21383] = a[13] & g[13191];
assign g[29574] = b[13] & g[13191];
assign g[21384] = a[13] & g[13192];
assign g[29575] = b[13] & g[13192];
assign g[21385] = a[13] & g[13193];
assign g[29576] = b[13] & g[13193];
assign g[21386] = a[13] & g[13194];
assign g[29577] = b[13] & g[13194];
assign g[21387] = a[13] & g[13195];
assign g[29578] = b[13] & g[13195];
assign g[21388] = a[13] & g[13196];
assign g[29579] = b[13] & g[13196];
assign g[21389] = a[13] & g[13197];
assign g[29580] = b[13] & g[13197];
assign g[21390] = a[13] & g[13198];
assign g[29581] = b[13] & g[13198];
assign g[21391] = a[13] & g[13199];
assign g[29582] = b[13] & g[13199];
assign g[21392] = a[13] & g[13200];
assign g[29583] = b[13] & g[13200];
assign g[21393] = a[13] & g[13201];
assign g[29584] = b[13] & g[13201];
assign g[21394] = a[13] & g[13202];
assign g[29585] = b[13] & g[13202];
assign g[21395] = a[13] & g[13203];
assign g[29586] = b[13] & g[13203];
assign g[21396] = a[13] & g[13204];
assign g[29587] = b[13] & g[13204];
assign g[21397] = a[13] & g[13205];
assign g[29588] = b[13] & g[13205];
assign g[21398] = a[13] & g[13206];
assign g[29589] = b[13] & g[13206];
assign g[21399] = a[13] & g[13207];
assign g[29590] = b[13] & g[13207];
assign g[21400] = a[13] & g[13208];
assign g[29591] = b[13] & g[13208];
assign g[21401] = a[13] & g[13209];
assign g[29592] = b[13] & g[13209];
assign g[21402] = a[13] & g[13210];
assign g[29593] = b[13] & g[13210];
assign g[21403] = a[13] & g[13211];
assign g[29594] = b[13] & g[13211];
assign g[21404] = a[13] & g[13212];
assign g[29595] = b[13] & g[13212];
assign g[21405] = a[13] & g[13213];
assign g[29596] = b[13] & g[13213];
assign g[21406] = a[13] & g[13214];
assign g[29597] = b[13] & g[13214];
assign g[21407] = a[13] & g[13215];
assign g[29598] = b[13] & g[13215];
assign g[21408] = a[13] & g[13216];
assign g[29599] = b[13] & g[13216];
assign g[21409] = a[13] & g[13217];
assign g[29600] = b[13] & g[13217];
assign g[21410] = a[13] & g[13218];
assign g[29601] = b[13] & g[13218];
assign g[21411] = a[13] & g[13219];
assign g[29602] = b[13] & g[13219];
assign g[21412] = a[13] & g[13220];
assign g[29603] = b[13] & g[13220];
assign g[21413] = a[13] & g[13221];
assign g[29604] = b[13] & g[13221];
assign g[21414] = a[13] & g[13222];
assign g[29605] = b[13] & g[13222];
assign g[21415] = a[13] & g[13223];
assign g[29606] = b[13] & g[13223];
assign g[21416] = a[13] & g[13224];
assign g[29607] = b[13] & g[13224];
assign g[21417] = a[13] & g[13225];
assign g[29608] = b[13] & g[13225];
assign g[21418] = a[13] & g[13226];
assign g[29609] = b[13] & g[13226];
assign g[21419] = a[13] & g[13227];
assign g[29610] = b[13] & g[13227];
assign g[21420] = a[13] & g[13228];
assign g[29611] = b[13] & g[13228];
assign g[21421] = a[13] & g[13229];
assign g[29612] = b[13] & g[13229];
assign g[21422] = a[13] & g[13230];
assign g[29613] = b[13] & g[13230];
assign g[21423] = a[13] & g[13231];
assign g[29614] = b[13] & g[13231];
assign g[21424] = a[13] & g[13232];
assign g[29615] = b[13] & g[13232];
assign g[21425] = a[13] & g[13233];
assign g[29616] = b[13] & g[13233];
assign g[21426] = a[13] & g[13234];
assign g[29617] = b[13] & g[13234];
assign g[21427] = a[13] & g[13235];
assign g[29618] = b[13] & g[13235];
assign g[21428] = a[13] & g[13236];
assign g[29619] = b[13] & g[13236];
assign g[21429] = a[13] & g[13237];
assign g[29620] = b[13] & g[13237];
assign g[21430] = a[13] & g[13238];
assign g[29621] = b[13] & g[13238];
assign g[21431] = a[13] & g[13239];
assign g[29622] = b[13] & g[13239];
assign g[21432] = a[13] & g[13240];
assign g[29623] = b[13] & g[13240];
assign g[21433] = a[13] & g[13241];
assign g[29624] = b[13] & g[13241];
assign g[21434] = a[13] & g[13242];
assign g[29625] = b[13] & g[13242];
assign g[21435] = a[13] & g[13243];
assign g[29626] = b[13] & g[13243];
assign g[21436] = a[13] & g[13244];
assign g[29627] = b[13] & g[13244];
assign g[21437] = a[13] & g[13245];
assign g[29628] = b[13] & g[13245];
assign g[21438] = a[13] & g[13246];
assign g[29629] = b[13] & g[13246];
assign g[21439] = a[13] & g[13247];
assign g[29630] = b[13] & g[13247];
assign g[21440] = a[13] & g[13248];
assign g[29631] = b[13] & g[13248];
assign g[21441] = a[13] & g[13249];
assign g[29632] = b[13] & g[13249];
assign g[21442] = a[13] & g[13250];
assign g[29633] = b[13] & g[13250];
assign g[21443] = a[13] & g[13251];
assign g[29634] = b[13] & g[13251];
assign g[21444] = a[13] & g[13252];
assign g[29635] = b[13] & g[13252];
assign g[21445] = a[13] & g[13253];
assign g[29636] = b[13] & g[13253];
assign g[21446] = a[13] & g[13254];
assign g[29637] = b[13] & g[13254];
assign g[21447] = a[13] & g[13255];
assign g[29638] = b[13] & g[13255];
assign g[21448] = a[13] & g[13256];
assign g[29639] = b[13] & g[13256];
assign g[21449] = a[13] & g[13257];
assign g[29640] = b[13] & g[13257];
assign g[21450] = a[13] & g[13258];
assign g[29641] = b[13] & g[13258];
assign g[21451] = a[13] & g[13259];
assign g[29642] = b[13] & g[13259];
assign g[21452] = a[13] & g[13260];
assign g[29643] = b[13] & g[13260];
assign g[21453] = a[13] & g[13261];
assign g[29644] = b[13] & g[13261];
assign g[21454] = a[13] & g[13262];
assign g[29645] = b[13] & g[13262];
assign g[21455] = a[13] & g[13263];
assign g[29646] = b[13] & g[13263];
assign g[21456] = a[13] & g[13264];
assign g[29647] = b[13] & g[13264];
assign g[21457] = a[13] & g[13265];
assign g[29648] = b[13] & g[13265];
assign g[21458] = a[13] & g[13266];
assign g[29649] = b[13] & g[13266];
assign g[21459] = a[13] & g[13267];
assign g[29650] = b[13] & g[13267];
assign g[21460] = a[13] & g[13268];
assign g[29651] = b[13] & g[13268];
assign g[21461] = a[13] & g[13269];
assign g[29652] = b[13] & g[13269];
assign g[21462] = a[13] & g[13270];
assign g[29653] = b[13] & g[13270];
assign g[21463] = a[13] & g[13271];
assign g[29654] = b[13] & g[13271];
assign g[21464] = a[13] & g[13272];
assign g[29655] = b[13] & g[13272];
assign g[21465] = a[13] & g[13273];
assign g[29656] = b[13] & g[13273];
assign g[21466] = a[13] & g[13274];
assign g[29657] = b[13] & g[13274];
assign g[21467] = a[13] & g[13275];
assign g[29658] = b[13] & g[13275];
assign g[21468] = a[13] & g[13276];
assign g[29659] = b[13] & g[13276];
assign g[21469] = a[13] & g[13277];
assign g[29660] = b[13] & g[13277];
assign g[21470] = a[13] & g[13278];
assign g[29661] = b[13] & g[13278];
assign g[21471] = a[13] & g[13279];
assign g[29662] = b[13] & g[13279];
assign g[21472] = a[13] & g[13280];
assign g[29663] = b[13] & g[13280];
assign g[21473] = a[13] & g[13281];
assign g[29664] = b[13] & g[13281];
assign g[21474] = a[13] & g[13282];
assign g[29665] = b[13] & g[13282];
assign g[21475] = a[13] & g[13283];
assign g[29666] = b[13] & g[13283];
assign g[21476] = a[13] & g[13284];
assign g[29667] = b[13] & g[13284];
assign g[21477] = a[13] & g[13285];
assign g[29668] = b[13] & g[13285];
assign g[21478] = a[13] & g[13286];
assign g[29669] = b[13] & g[13286];
assign g[21479] = a[13] & g[13287];
assign g[29670] = b[13] & g[13287];
assign g[21480] = a[13] & g[13288];
assign g[29671] = b[13] & g[13288];
assign g[21481] = a[13] & g[13289];
assign g[29672] = b[13] & g[13289];
assign g[21482] = a[13] & g[13290];
assign g[29673] = b[13] & g[13290];
assign g[21483] = a[13] & g[13291];
assign g[29674] = b[13] & g[13291];
assign g[21484] = a[13] & g[13292];
assign g[29675] = b[13] & g[13292];
assign g[21485] = a[13] & g[13293];
assign g[29676] = b[13] & g[13293];
assign g[21486] = a[13] & g[13294];
assign g[29677] = b[13] & g[13294];
assign g[21487] = a[13] & g[13295];
assign g[29678] = b[13] & g[13295];
assign g[21488] = a[13] & g[13296];
assign g[29679] = b[13] & g[13296];
assign g[21489] = a[13] & g[13297];
assign g[29680] = b[13] & g[13297];
assign g[21490] = a[13] & g[13298];
assign g[29681] = b[13] & g[13298];
assign g[21491] = a[13] & g[13299];
assign g[29682] = b[13] & g[13299];
assign g[21492] = a[13] & g[13300];
assign g[29683] = b[13] & g[13300];
assign g[21493] = a[13] & g[13301];
assign g[29684] = b[13] & g[13301];
assign g[21494] = a[13] & g[13302];
assign g[29685] = b[13] & g[13302];
assign g[21495] = a[13] & g[13303];
assign g[29686] = b[13] & g[13303];
assign g[21496] = a[13] & g[13304];
assign g[29687] = b[13] & g[13304];
assign g[21497] = a[13] & g[13305];
assign g[29688] = b[13] & g[13305];
assign g[21498] = a[13] & g[13306];
assign g[29689] = b[13] & g[13306];
assign g[21499] = a[13] & g[13307];
assign g[29690] = b[13] & g[13307];
assign g[21500] = a[13] & g[13308];
assign g[29691] = b[13] & g[13308];
assign g[21501] = a[13] & g[13309];
assign g[29692] = b[13] & g[13309];
assign g[21502] = a[13] & g[13310];
assign g[29693] = b[13] & g[13310];
assign g[21503] = a[13] & g[13311];
assign g[29694] = b[13] & g[13311];
assign g[21504] = a[13] & g[13312];
assign g[29695] = b[13] & g[13312];
assign g[21505] = a[13] & g[13313];
assign g[29696] = b[13] & g[13313];
assign g[21506] = a[13] & g[13314];
assign g[29697] = b[13] & g[13314];
assign g[21507] = a[13] & g[13315];
assign g[29698] = b[13] & g[13315];
assign g[21508] = a[13] & g[13316];
assign g[29699] = b[13] & g[13316];
assign g[21509] = a[13] & g[13317];
assign g[29700] = b[13] & g[13317];
assign g[21510] = a[13] & g[13318];
assign g[29701] = b[13] & g[13318];
assign g[21511] = a[13] & g[13319];
assign g[29702] = b[13] & g[13319];
assign g[21512] = a[13] & g[13320];
assign g[29703] = b[13] & g[13320];
assign g[21513] = a[13] & g[13321];
assign g[29704] = b[13] & g[13321];
assign g[21514] = a[13] & g[13322];
assign g[29705] = b[13] & g[13322];
assign g[21515] = a[13] & g[13323];
assign g[29706] = b[13] & g[13323];
assign g[21516] = a[13] & g[13324];
assign g[29707] = b[13] & g[13324];
assign g[21517] = a[13] & g[13325];
assign g[29708] = b[13] & g[13325];
assign g[21518] = a[13] & g[13326];
assign g[29709] = b[13] & g[13326];
assign g[21519] = a[13] & g[13327];
assign g[29710] = b[13] & g[13327];
assign g[21520] = a[13] & g[13328];
assign g[29711] = b[13] & g[13328];
assign g[21521] = a[13] & g[13329];
assign g[29712] = b[13] & g[13329];
assign g[21522] = a[13] & g[13330];
assign g[29713] = b[13] & g[13330];
assign g[21523] = a[13] & g[13331];
assign g[29714] = b[13] & g[13331];
assign g[21524] = a[13] & g[13332];
assign g[29715] = b[13] & g[13332];
assign g[21525] = a[13] & g[13333];
assign g[29716] = b[13] & g[13333];
assign g[21526] = a[13] & g[13334];
assign g[29717] = b[13] & g[13334];
assign g[21527] = a[13] & g[13335];
assign g[29718] = b[13] & g[13335];
assign g[21528] = a[13] & g[13336];
assign g[29719] = b[13] & g[13336];
assign g[21529] = a[13] & g[13337];
assign g[29720] = b[13] & g[13337];
assign g[21530] = a[13] & g[13338];
assign g[29721] = b[13] & g[13338];
assign g[21531] = a[13] & g[13339];
assign g[29722] = b[13] & g[13339];
assign g[21532] = a[13] & g[13340];
assign g[29723] = b[13] & g[13340];
assign g[21533] = a[13] & g[13341];
assign g[29724] = b[13] & g[13341];
assign g[21534] = a[13] & g[13342];
assign g[29725] = b[13] & g[13342];
assign g[21535] = a[13] & g[13343];
assign g[29726] = b[13] & g[13343];
assign g[21536] = a[13] & g[13344];
assign g[29727] = b[13] & g[13344];
assign g[21537] = a[13] & g[13345];
assign g[29728] = b[13] & g[13345];
assign g[21538] = a[13] & g[13346];
assign g[29729] = b[13] & g[13346];
assign g[21539] = a[13] & g[13347];
assign g[29730] = b[13] & g[13347];
assign g[21540] = a[13] & g[13348];
assign g[29731] = b[13] & g[13348];
assign g[21541] = a[13] & g[13349];
assign g[29732] = b[13] & g[13349];
assign g[21542] = a[13] & g[13350];
assign g[29733] = b[13] & g[13350];
assign g[21543] = a[13] & g[13351];
assign g[29734] = b[13] & g[13351];
assign g[21544] = a[13] & g[13352];
assign g[29735] = b[13] & g[13352];
assign g[21545] = a[13] & g[13353];
assign g[29736] = b[13] & g[13353];
assign g[21546] = a[13] & g[13354];
assign g[29737] = b[13] & g[13354];
assign g[21547] = a[13] & g[13355];
assign g[29738] = b[13] & g[13355];
assign g[21548] = a[13] & g[13356];
assign g[29739] = b[13] & g[13356];
assign g[21549] = a[13] & g[13357];
assign g[29740] = b[13] & g[13357];
assign g[21550] = a[13] & g[13358];
assign g[29741] = b[13] & g[13358];
assign g[21551] = a[13] & g[13359];
assign g[29742] = b[13] & g[13359];
assign g[21552] = a[13] & g[13360];
assign g[29743] = b[13] & g[13360];
assign g[21553] = a[13] & g[13361];
assign g[29744] = b[13] & g[13361];
assign g[21554] = a[13] & g[13362];
assign g[29745] = b[13] & g[13362];
assign g[21555] = a[13] & g[13363];
assign g[29746] = b[13] & g[13363];
assign g[21556] = a[13] & g[13364];
assign g[29747] = b[13] & g[13364];
assign g[21557] = a[13] & g[13365];
assign g[29748] = b[13] & g[13365];
assign g[21558] = a[13] & g[13366];
assign g[29749] = b[13] & g[13366];
assign g[21559] = a[13] & g[13367];
assign g[29750] = b[13] & g[13367];
assign g[21560] = a[13] & g[13368];
assign g[29751] = b[13] & g[13368];
assign g[21561] = a[13] & g[13369];
assign g[29752] = b[13] & g[13369];
assign g[21562] = a[13] & g[13370];
assign g[29753] = b[13] & g[13370];
assign g[21563] = a[13] & g[13371];
assign g[29754] = b[13] & g[13371];
assign g[21564] = a[13] & g[13372];
assign g[29755] = b[13] & g[13372];
assign g[21565] = a[13] & g[13373];
assign g[29756] = b[13] & g[13373];
assign g[21566] = a[13] & g[13374];
assign g[29757] = b[13] & g[13374];
assign g[21567] = a[13] & g[13375];
assign g[29758] = b[13] & g[13375];
assign g[21568] = a[13] & g[13376];
assign g[29759] = b[13] & g[13376];
assign g[21569] = a[13] & g[13377];
assign g[29760] = b[13] & g[13377];
assign g[21570] = a[13] & g[13378];
assign g[29761] = b[13] & g[13378];
assign g[21571] = a[13] & g[13379];
assign g[29762] = b[13] & g[13379];
assign g[21572] = a[13] & g[13380];
assign g[29763] = b[13] & g[13380];
assign g[21573] = a[13] & g[13381];
assign g[29764] = b[13] & g[13381];
assign g[21574] = a[13] & g[13382];
assign g[29765] = b[13] & g[13382];
assign g[21575] = a[13] & g[13383];
assign g[29766] = b[13] & g[13383];
assign g[21576] = a[13] & g[13384];
assign g[29767] = b[13] & g[13384];
assign g[21577] = a[13] & g[13385];
assign g[29768] = b[13] & g[13385];
assign g[21578] = a[13] & g[13386];
assign g[29769] = b[13] & g[13386];
assign g[21579] = a[13] & g[13387];
assign g[29770] = b[13] & g[13387];
assign g[21580] = a[13] & g[13388];
assign g[29771] = b[13] & g[13388];
assign g[21581] = a[13] & g[13389];
assign g[29772] = b[13] & g[13389];
assign g[21582] = a[13] & g[13390];
assign g[29773] = b[13] & g[13390];
assign g[21583] = a[13] & g[13391];
assign g[29774] = b[13] & g[13391];
assign g[21584] = a[13] & g[13392];
assign g[29775] = b[13] & g[13392];
assign g[21585] = a[13] & g[13393];
assign g[29776] = b[13] & g[13393];
assign g[21586] = a[13] & g[13394];
assign g[29777] = b[13] & g[13394];
assign g[21587] = a[13] & g[13395];
assign g[29778] = b[13] & g[13395];
assign g[21588] = a[13] & g[13396];
assign g[29779] = b[13] & g[13396];
assign g[21589] = a[13] & g[13397];
assign g[29780] = b[13] & g[13397];
assign g[21590] = a[13] & g[13398];
assign g[29781] = b[13] & g[13398];
assign g[21591] = a[13] & g[13399];
assign g[29782] = b[13] & g[13399];
assign g[21592] = a[13] & g[13400];
assign g[29783] = b[13] & g[13400];
assign g[21593] = a[13] & g[13401];
assign g[29784] = b[13] & g[13401];
assign g[21594] = a[13] & g[13402];
assign g[29785] = b[13] & g[13402];
assign g[21595] = a[13] & g[13403];
assign g[29786] = b[13] & g[13403];
assign g[21596] = a[13] & g[13404];
assign g[29787] = b[13] & g[13404];
assign g[21597] = a[13] & g[13405];
assign g[29788] = b[13] & g[13405];
assign g[21598] = a[13] & g[13406];
assign g[29789] = b[13] & g[13406];
assign g[21599] = a[13] & g[13407];
assign g[29790] = b[13] & g[13407];
assign g[21600] = a[13] & g[13408];
assign g[29791] = b[13] & g[13408];
assign g[21601] = a[13] & g[13409];
assign g[29792] = b[13] & g[13409];
assign g[21602] = a[13] & g[13410];
assign g[29793] = b[13] & g[13410];
assign g[21603] = a[13] & g[13411];
assign g[29794] = b[13] & g[13411];
assign g[21604] = a[13] & g[13412];
assign g[29795] = b[13] & g[13412];
assign g[21605] = a[13] & g[13413];
assign g[29796] = b[13] & g[13413];
assign g[21606] = a[13] & g[13414];
assign g[29797] = b[13] & g[13414];
assign g[21607] = a[13] & g[13415];
assign g[29798] = b[13] & g[13415];
assign g[21608] = a[13] & g[13416];
assign g[29799] = b[13] & g[13416];
assign g[21609] = a[13] & g[13417];
assign g[29800] = b[13] & g[13417];
assign g[21610] = a[13] & g[13418];
assign g[29801] = b[13] & g[13418];
assign g[21611] = a[13] & g[13419];
assign g[29802] = b[13] & g[13419];
assign g[21612] = a[13] & g[13420];
assign g[29803] = b[13] & g[13420];
assign g[21613] = a[13] & g[13421];
assign g[29804] = b[13] & g[13421];
assign g[21614] = a[13] & g[13422];
assign g[29805] = b[13] & g[13422];
assign g[21615] = a[13] & g[13423];
assign g[29806] = b[13] & g[13423];
assign g[21616] = a[13] & g[13424];
assign g[29807] = b[13] & g[13424];
assign g[21617] = a[13] & g[13425];
assign g[29808] = b[13] & g[13425];
assign g[21618] = a[13] & g[13426];
assign g[29809] = b[13] & g[13426];
assign g[21619] = a[13] & g[13427];
assign g[29810] = b[13] & g[13427];
assign g[21620] = a[13] & g[13428];
assign g[29811] = b[13] & g[13428];
assign g[21621] = a[13] & g[13429];
assign g[29812] = b[13] & g[13429];
assign g[21622] = a[13] & g[13430];
assign g[29813] = b[13] & g[13430];
assign g[21623] = a[13] & g[13431];
assign g[29814] = b[13] & g[13431];
assign g[21624] = a[13] & g[13432];
assign g[29815] = b[13] & g[13432];
assign g[21625] = a[13] & g[13433];
assign g[29816] = b[13] & g[13433];
assign g[21626] = a[13] & g[13434];
assign g[29817] = b[13] & g[13434];
assign g[21627] = a[13] & g[13435];
assign g[29818] = b[13] & g[13435];
assign g[21628] = a[13] & g[13436];
assign g[29819] = b[13] & g[13436];
assign g[21629] = a[13] & g[13437];
assign g[29820] = b[13] & g[13437];
assign g[21630] = a[13] & g[13438];
assign g[29821] = b[13] & g[13438];
assign g[21631] = a[13] & g[13439];
assign g[29822] = b[13] & g[13439];
assign g[21632] = a[13] & g[13440];
assign g[29823] = b[13] & g[13440];
assign g[21633] = a[13] & g[13441];
assign g[29824] = b[13] & g[13441];
assign g[21634] = a[13] & g[13442];
assign g[29825] = b[13] & g[13442];
assign g[21635] = a[13] & g[13443];
assign g[29826] = b[13] & g[13443];
assign g[21636] = a[13] & g[13444];
assign g[29827] = b[13] & g[13444];
assign g[21637] = a[13] & g[13445];
assign g[29828] = b[13] & g[13445];
assign g[21638] = a[13] & g[13446];
assign g[29829] = b[13] & g[13446];
assign g[21639] = a[13] & g[13447];
assign g[29830] = b[13] & g[13447];
assign g[21640] = a[13] & g[13448];
assign g[29831] = b[13] & g[13448];
assign g[21641] = a[13] & g[13449];
assign g[29832] = b[13] & g[13449];
assign g[21642] = a[13] & g[13450];
assign g[29833] = b[13] & g[13450];
assign g[21643] = a[13] & g[13451];
assign g[29834] = b[13] & g[13451];
assign g[21644] = a[13] & g[13452];
assign g[29835] = b[13] & g[13452];
assign g[21645] = a[13] & g[13453];
assign g[29836] = b[13] & g[13453];
assign g[21646] = a[13] & g[13454];
assign g[29837] = b[13] & g[13454];
assign g[21647] = a[13] & g[13455];
assign g[29838] = b[13] & g[13455];
assign g[21648] = a[13] & g[13456];
assign g[29839] = b[13] & g[13456];
assign g[21649] = a[13] & g[13457];
assign g[29840] = b[13] & g[13457];
assign g[21650] = a[13] & g[13458];
assign g[29841] = b[13] & g[13458];
assign g[21651] = a[13] & g[13459];
assign g[29842] = b[13] & g[13459];
assign g[21652] = a[13] & g[13460];
assign g[29843] = b[13] & g[13460];
assign g[21653] = a[13] & g[13461];
assign g[29844] = b[13] & g[13461];
assign g[21654] = a[13] & g[13462];
assign g[29845] = b[13] & g[13462];
assign g[21655] = a[13] & g[13463];
assign g[29846] = b[13] & g[13463];
assign g[21656] = a[13] & g[13464];
assign g[29847] = b[13] & g[13464];
assign g[21657] = a[13] & g[13465];
assign g[29848] = b[13] & g[13465];
assign g[21658] = a[13] & g[13466];
assign g[29849] = b[13] & g[13466];
assign g[21659] = a[13] & g[13467];
assign g[29850] = b[13] & g[13467];
assign g[21660] = a[13] & g[13468];
assign g[29851] = b[13] & g[13468];
assign g[21661] = a[13] & g[13469];
assign g[29852] = b[13] & g[13469];
assign g[21662] = a[13] & g[13470];
assign g[29853] = b[13] & g[13470];
assign g[21663] = a[13] & g[13471];
assign g[29854] = b[13] & g[13471];
assign g[21664] = a[13] & g[13472];
assign g[29855] = b[13] & g[13472];
assign g[21665] = a[13] & g[13473];
assign g[29856] = b[13] & g[13473];
assign g[21666] = a[13] & g[13474];
assign g[29857] = b[13] & g[13474];
assign g[21667] = a[13] & g[13475];
assign g[29858] = b[13] & g[13475];
assign g[21668] = a[13] & g[13476];
assign g[29859] = b[13] & g[13476];
assign g[21669] = a[13] & g[13477];
assign g[29860] = b[13] & g[13477];
assign g[21670] = a[13] & g[13478];
assign g[29861] = b[13] & g[13478];
assign g[21671] = a[13] & g[13479];
assign g[29862] = b[13] & g[13479];
assign g[21672] = a[13] & g[13480];
assign g[29863] = b[13] & g[13480];
assign g[21673] = a[13] & g[13481];
assign g[29864] = b[13] & g[13481];
assign g[21674] = a[13] & g[13482];
assign g[29865] = b[13] & g[13482];
assign g[21675] = a[13] & g[13483];
assign g[29866] = b[13] & g[13483];
assign g[21676] = a[13] & g[13484];
assign g[29867] = b[13] & g[13484];
assign g[21677] = a[13] & g[13485];
assign g[29868] = b[13] & g[13485];
assign g[21678] = a[13] & g[13486];
assign g[29869] = b[13] & g[13486];
assign g[21679] = a[13] & g[13487];
assign g[29870] = b[13] & g[13487];
assign g[21680] = a[13] & g[13488];
assign g[29871] = b[13] & g[13488];
assign g[21681] = a[13] & g[13489];
assign g[29872] = b[13] & g[13489];
assign g[21682] = a[13] & g[13490];
assign g[29873] = b[13] & g[13490];
assign g[21683] = a[13] & g[13491];
assign g[29874] = b[13] & g[13491];
assign g[21684] = a[13] & g[13492];
assign g[29875] = b[13] & g[13492];
assign g[21685] = a[13] & g[13493];
assign g[29876] = b[13] & g[13493];
assign g[21686] = a[13] & g[13494];
assign g[29877] = b[13] & g[13494];
assign g[21687] = a[13] & g[13495];
assign g[29878] = b[13] & g[13495];
assign g[21688] = a[13] & g[13496];
assign g[29879] = b[13] & g[13496];
assign g[21689] = a[13] & g[13497];
assign g[29880] = b[13] & g[13497];
assign g[21690] = a[13] & g[13498];
assign g[29881] = b[13] & g[13498];
assign g[21691] = a[13] & g[13499];
assign g[29882] = b[13] & g[13499];
assign g[21692] = a[13] & g[13500];
assign g[29883] = b[13] & g[13500];
assign g[21693] = a[13] & g[13501];
assign g[29884] = b[13] & g[13501];
assign g[21694] = a[13] & g[13502];
assign g[29885] = b[13] & g[13502];
assign g[21695] = a[13] & g[13503];
assign g[29886] = b[13] & g[13503];
assign g[21696] = a[13] & g[13504];
assign g[29887] = b[13] & g[13504];
assign g[21697] = a[13] & g[13505];
assign g[29888] = b[13] & g[13505];
assign g[21698] = a[13] & g[13506];
assign g[29889] = b[13] & g[13506];
assign g[21699] = a[13] & g[13507];
assign g[29890] = b[13] & g[13507];
assign g[21700] = a[13] & g[13508];
assign g[29891] = b[13] & g[13508];
assign g[21701] = a[13] & g[13509];
assign g[29892] = b[13] & g[13509];
assign g[21702] = a[13] & g[13510];
assign g[29893] = b[13] & g[13510];
assign g[21703] = a[13] & g[13511];
assign g[29894] = b[13] & g[13511];
assign g[21704] = a[13] & g[13512];
assign g[29895] = b[13] & g[13512];
assign g[21705] = a[13] & g[13513];
assign g[29896] = b[13] & g[13513];
assign g[21706] = a[13] & g[13514];
assign g[29897] = b[13] & g[13514];
assign g[21707] = a[13] & g[13515];
assign g[29898] = b[13] & g[13515];
assign g[21708] = a[13] & g[13516];
assign g[29899] = b[13] & g[13516];
assign g[21709] = a[13] & g[13517];
assign g[29900] = b[13] & g[13517];
assign g[21710] = a[13] & g[13518];
assign g[29901] = b[13] & g[13518];
assign g[21711] = a[13] & g[13519];
assign g[29902] = b[13] & g[13519];
assign g[21712] = a[13] & g[13520];
assign g[29903] = b[13] & g[13520];
assign g[21713] = a[13] & g[13521];
assign g[29904] = b[13] & g[13521];
assign g[21714] = a[13] & g[13522];
assign g[29905] = b[13] & g[13522];
assign g[21715] = a[13] & g[13523];
assign g[29906] = b[13] & g[13523];
assign g[21716] = a[13] & g[13524];
assign g[29907] = b[13] & g[13524];
assign g[21717] = a[13] & g[13525];
assign g[29908] = b[13] & g[13525];
assign g[21718] = a[13] & g[13526];
assign g[29909] = b[13] & g[13526];
assign g[21719] = a[13] & g[13527];
assign g[29910] = b[13] & g[13527];
assign g[21720] = a[13] & g[13528];
assign g[29911] = b[13] & g[13528];
assign g[21721] = a[13] & g[13529];
assign g[29912] = b[13] & g[13529];
assign g[21722] = a[13] & g[13530];
assign g[29913] = b[13] & g[13530];
assign g[21723] = a[13] & g[13531];
assign g[29914] = b[13] & g[13531];
assign g[21724] = a[13] & g[13532];
assign g[29915] = b[13] & g[13532];
assign g[21725] = a[13] & g[13533];
assign g[29916] = b[13] & g[13533];
assign g[21726] = a[13] & g[13534];
assign g[29917] = b[13] & g[13534];
assign g[21727] = a[13] & g[13535];
assign g[29918] = b[13] & g[13535];
assign g[21728] = a[13] & g[13536];
assign g[29919] = b[13] & g[13536];
assign g[21729] = a[13] & g[13537];
assign g[29920] = b[13] & g[13537];
assign g[21730] = a[13] & g[13538];
assign g[29921] = b[13] & g[13538];
assign g[21731] = a[13] & g[13539];
assign g[29922] = b[13] & g[13539];
assign g[21732] = a[13] & g[13540];
assign g[29923] = b[13] & g[13540];
assign g[21733] = a[13] & g[13541];
assign g[29924] = b[13] & g[13541];
assign g[21734] = a[13] & g[13542];
assign g[29925] = b[13] & g[13542];
assign g[21735] = a[13] & g[13543];
assign g[29926] = b[13] & g[13543];
assign g[21736] = a[13] & g[13544];
assign g[29927] = b[13] & g[13544];
assign g[21737] = a[13] & g[13545];
assign g[29928] = b[13] & g[13545];
assign g[21738] = a[13] & g[13546];
assign g[29929] = b[13] & g[13546];
assign g[21739] = a[13] & g[13547];
assign g[29930] = b[13] & g[13547];
assign g[21740] = a[13] & g[13548];
assign g[29931] = b[13] & g[13548];
assign g[21741] = a[13] & g[13549];
assign g[29932] = b[13] & g[13549];
assign g[21742] = a[13] & g[13550];
assign g[29933] = b[13] & g[13550];
assign g[21743] = a[13] & g[13551];
assign g[29934] = b[13] & g[13551];
assign g[21744] = a[13] & g[13552];
assign g[29935] = b[13] & g[13552];
assign g[21745] = a[13] & g[13553];
assign g[29936] = b[13] & g[13553];
assign g[21746] = a[13] & g[13554];
assign g[29937] = b[13] & g[13554];
assign g[21747] = a[13] & g[13555];
assign g[29938] = b[13] & g[13555];
assign g[21748] = a[13] & g[13556];
assign g[29939] = b[13] & g[13556];
assign g[21749] = a[13] & g[13557];
assign g[29940] = b[13] & g[13557];
assign g[21750] = a[13] & g[13558];
assign g[29941] = b[13] & g[13558];
assign g[21751] = a[13] & g[13559];
assign g[29942] = b[13] & g[13559];
assign g[21752] = a[13] & g[13560];
assign g[29943] = b[13] & g[13560];
assign g[21753] = a[13] & g[13561];
assign g[29944] = b[13] & g[13561];
assign g[21754] = a[13] & g[13562];
assign g[29945] = b[13] & g[13562];
assign g[21755] = a[13] & g[13563];
assign g[29946] = b[13] & g[13563];
assign g[21756] = a[13] & g[13564];
assign g[29947] = b[13] & g[13564];
assign g[21757] = a[13] & g[13565];
assign g[29948] = b[13] & g[13565];
assign g[21758] = a[13] & g[13566];
assign g[29949] = b[13] & g[13566];
assign g[21759] = a[13] & g[13567];
assign g[29950] = b[13] & g[13567];
assign g[21760] = a[13] & g[13568];
assign g[29951] = b[13] & g[13568];
assign g[21761] = a[13] & g[13569];
assign g[29952] = b[13] & g[13569];
assign g[21762] = a[13] & g[13570];
assign g[29953] = b[13] & g[13570];
assign g[21763] = a[13] & g[13571];
assign g[29954] = b[13] & g[13571];
assign g[21764] = a[13] & g[13572];
assign g[29955] = b[13] & g[13572];
assign g[21765] = a[13] & g[13573];
assign g[29956] = b[13] & g[13573];
assign g[21766] = a[13] & g[13574];
assign g[29957] = b[13] & g[13574];
assign g[21767] = a[13] & g[13575];
assign g[29958] = b[13] & g[13575];
assign g[21768] = a[13] & g[13576];
assign g[29959] = b[13] & g[13576];
assign g[21769] = a[13] & g[13577];
assign g[29960] = b[13] & g[13577];
assign g[21770] = a[13] & g[13578];
assign g[29961] = b[13] & g[13578];
assign g[21771] = a[13] & g[13579];
assign g[29962] = b[13] & g[13579];
assign g[21772] = a[13] & g[13580];
assign g[29963] = b[13] & g[13580];
assign g[21773] = a[13] & g[13581];
assign g[29964] = b[13] & g[13581];
assign g[21774] = a[13] & g[13582];
assign g[29965] = b[13] & g[13582];
assign g[21775] = a[13] & g[13583];
assign g[29966] = b[13] & g[13583];
assign g[21776] = a[13] & g[13584];
assign g[29967] = b[13] & g[13584];
assign g[21777] = a[13] & g[13585];
assign g[29968] = b[13] & g[13585];
assign g[21778] = a[13] & g[13586];
assign g[29969] = b[13] & g[13586];
assign g[21779] = a[13] & g[13587];
assign g[29970] = b[13] & g[13587];
assign g[21780] = a[13] & g[13588];
assign g[29971] = b[13] & g[13588];
assign g[21781] = a[13] & g[13589];
assign g[29972] = b[13] & g[13589];
assign g[21782] = a[13] & g[13590];
assign g[29973] = b[13] & g[13590];
assign g[21783] = a[13] & g[13591];
assign g[29974] = b[13] & g[13591];
assign g[21784] = a[13] & g[13592];
assign g[29975] = b[13] & g[13592];
assign g[21785] = a[13] & g[13593];
assign g[29976] = b[13] & g[13593];
assign g[21786] = a[13] & g[13594];
assign g[29977] = b[13] & g[13594];
assign g[21787] = a[13] & g[13595];
assign g[29978] = b[13] & g[13595];
assign g[21788] = a[13] & g[13596];
assign g[29979] = b[13] & g[13596];
assign g[21789] = a[13] & g[13597];
assign g[29980] = b[13] & g[13597];
assign g[21790] = a[13] & g[13598];
assign g[29981] = b[13] & g[13598];
assign g[21791] = a[13] & g[13599];
assign g[29982] = b[13] & g[13599];
assign g[21792] = a[13] & g[13600];
assign g[29983] = b[13] & g[13600];
assign g[21793] = a[13] & g[13601];
assign g[29984] = b[13] & g[13601];
assign g[21794] = a[13] & g[13602];
assign g[29985] = b[13] & g[13602];
assign g[21795] = a[13] & g[13603];
assign g[29986] = b[13] & g[13603];
assign g[21796] = a[13] & g[13604];
assign g[29987] = b[13] & g[13604];
assign g[21797] = a[13] & g[13605];
assign g[29988] = b[13] & g[13605];
assign g[21798] = a[13] & g[13606];
assign g[29989] = b[13] & g[13606];
assign g[21799] = a[13] & g[13607];
assign g[29990] = b[13] & g[13607];
assign g[21800] = a[13] & g[13608];
assign g[29991] = b[13] & g[13608];
assign g[21801] = a[13] & g[13609];
assign g[29992] = b[13] & g[13609];
assign g[21802] = a[13] & g[13610];
assign g[29993] = b[13] & g[13610];
assign g[21803] = a[13] & g[13611];
assign g[29994] = b[13] & g[13611];
assign g[21804] = a[13] & g[13612];
assign g[29995] = b[13] & g[13612];
assign g[21805] = a[13] & g[13613];
assign g[29996] = b[13] & g[13613];
assign g[21806] = a[13] & g[13614];
assign g[29997] = b[13] & g[13614];
assign g[21807] = a[13] & g[13615];
assign g[29998] = b[13] & g[13615];
assign g[21808] = a[13] & g[13616];
assign g[29999] = b[13] & g[13616];
assign g[21809] = a[13] & g[13617];
assign g[30000] = b[13] & g[13617];
assign g[21810] = a[13] & g[13618];
assign g[30001] = b[13] & g[13618];
assign g[21811] = a[13] & g[13619];
assign g[30002] = b[13] & g[13619];
assign g[21812] = a[13] & g[13620];
assign g[30003] = b[13] & g[13620];
assign g[21813] = a[13] & g[13621];
assign g[30004] = b[13] & g[13621];
assign g[21814] = a[13] & g[13622];
assign g[30005] = b[13] & g[13622];
assign g[21815] = a[13] & g[13623];
assign g[30006] = b[13] & g[13623];
assign g[21816] = a[13] & g[13624];
assign g[30007] = b[13] & g[13624];
assign g[21817] = a[13] & g[13625];
assign g[30008] = b[13] & g[13625];
assign g[21818] = a[13] & g[13626];
assign g[30009] = b[13] & g[13626];
assign g[21819] = a[13] & g[13627];
assign g[30010] = b[13] & g[13627];
assign g[21820] = a[13] & g[13628];
assign g[30011] = b[13] & g[13628];
assign g[21821] = a[13] & g[13629];
assign g[30012] = b[13] & g[13629];
assign g[21822] = a[13] & g[13630];
assign g[30013] = b[13] & g[13630];
assign g[21823] = a[13] & g[13631];
assign g[30014] = b[13] & g[13631];
assign g[21824] = a[13] & g[13632];
assign g[30015] = b[13] & g[13632];
assign g[21825] = a[13] & g[13633];
assign g[30016] = b[13] & g[13633];
assign g[21826] = a[13] & g[13634];
assign g[30017] = b[13] & g[13634];
assign g[21827] = a[13] & g[13635];
assign g[30018] = b[13] & g[13635];
assign g[21828] = a[13] & g[13636];
assign g[30019] = b[13] & g[13636];
assign g[21829] = a[13] & g[13637];
assign g[30020] = b[13] & g[13637];
assign g[21830] = a[13] & g[13638];
assign g[30021] = b[13] & g[13638];
assign g[21831] = a[13] & g[13639];
assign g[30022] = b[13] & g[13639];
assign g[21832] = a[13] & g[13640];
assign g[30023] = b[13] & g[13640];
assign g[21833] = a[13] & g[13641];
assign g[30024] = b[13] & g[13641];
assign g[21834] = a[13] & g[13642];
assign g[30025] = b[13] & g[13642];
assign g[21835] = a[13] & g[13643];
assign g[30026] = b[13] & g[13643];
assign g[21836] = a[13] & g[13644];
assign g[30027] = b[13] & g[13644];
assign g[21837] = a[13] & g[13645];
assign g[30028] = b[13] & g[13645];
assign g[21838] = a[13] & g[13646];
assign g[30029] = b[13] & g[13646];
assign g[21839] = a[13] & g[13647];
assign g[30030] = b[13] & g[13647];
assign g[21840] = a[13] & g[13648];
assign g[30031] = b[13] & g[13648];
assign g[21841] = a[13] & g[13649];
assign g[30032] = b[13] & g[13649];
assign g[21842] = a[13] & g[13650];
assign g[30033] = b[13] & g[13650];
assign g[21843] = a[13] & g[13651];
assign g[30034] = b[13] & g[13651];
assign g[21844] = a[13] & g[13652];
assign g[30035] = b[13] & g[13652];
assign g[21845] = a[13] & g[13653];
assign g[30036] = b[13] & g[13653];
assign g[21846] = a[13] & g[13654];
assign g[30037] = b[13] & g[13654];
assign g[21847] = a[13] & g[13655];
assign g[30038] = b[13] & g[13655];
assign g[21848] = a[13] & g[13656];
assign g[30039] = b[13] & g[13656];
assign g[21849] = a[13] & g[13657];
assign g[30040] = b[13] & g[13657];
assign g[21850] = a[13] & g[13658];
assign g[30041] = b[13] & g[13658];
assign g[21851] = a[13] & g[13659];
assign g[30042] = b[13] & g[13659];
assign g[21852] = a[13] & g[13660];
assign g[30043] = b[13] & g[13660];
assign g[21853] = a[13] & g[13661];
assign g[30044] = b[13] & g[13661];
assign g[21854] = a[13] & g[13662];
assign g[30045] = b[13] & g[13662];
assign g[21855] = a[13] & g[13663];
assign g[30046] = b[13] & g[13663];
assign g[21856] = a[13] & g[13664];
assign g[30047] = b[13] & g[13664];
assign g[21857] = a[13] & g[13665];
assign g[30048] = b[13] & g[13665];
assign g[21858] = a[13] & g[13666];
assign g[30049] = b[13] & g[13666];
assign g[21859] = a[13] & g[13667];
assign g[30050] = b[13] & g[13667];
assign g[21860] = a[13] & g[13668];
assign g[30051] = b[13] & g[13668];
assign g[21861] = a[13] & g[13669];
assign g[30052] = b[13] & g[13669];
assign g[21862] = a[13] & g[13670];
assign g[30053] = b[13] & g[13670];
assign g[21863] = a[13] & g[13671];
assign g[30054] = b[13] & g[13671];
assign g[21864] = a[13] & g[13672];
assign g[30055] = b[13] & g[13672];
assign g[21865] = a[13] & g[13673];
assign g[30056] = b[13] & g[13673];
assign g[21866] = a[13] & g[13674];
assign g[30057] = b[13] & g[13674];
assign g[21867] = a[13] & g[13675];
assign g[30058] = b[13] & g[13675];
assign g[21868] = a[13] & g[13676];
assign g[30059] = b[13] & g[13676];
assign g[21869] = a[13] & g[13677];
assign g[30060] = b[13] & g[13677];
assign g[21870] = a[13] & g[13678];
assign g[30061] = b[13] & g[13678];
assign g[21871] = a[13] & g[13679];
assign g[30062] = b[13] & g[13679];
assign g[21872] = a[13] & g[13680];
assign g[30063] = b[13] & g[13680];
assign g[21873] = a[13] & g[13681];
assign g[30064] = b[13] & g[13681];
assign g[21874] = a[13] & g[13682];
assign g[30065] = b[13] & g[13682];
assign g[21875] = a[13] & g[13683];
assign g[30066] = b[13] & g[13683];
assign g[21876] = a[13] & g[13684];
assign g[30067] = b[13] & g[13684];
assign g[21877] = a[13] & g[13685];
assign g[30068] = b[13] & g[13685];
assign g[21878] = a[13] & g[13686];
assign g[30069] = b[13] & g[13686];
assign g[21879] = a[13] & g[13687];
assign g[30070] = b[13] & g[13687];
assign g[21880] = a[13] & g[13688];
assign g[30071] = b[13] & g[13688];
assign g[21881] = a[13] & g[13689];
assign g[30072] = b[13] & g[13689];
assign g[21882] = a[13] & g[13690];
assign g[30073] = b[13] & g[13690];
assign g[21883] = a[13] & g[13691];
assign g[30074] = b[13] & g[13691];
assign g[21884] = a[13] & g[13692];
assign g[30075] = b[13] & g[13692];
assign g[21885] = a[13] & g[13693];
assign g[30076] = b[13] & g[13693];
assign g[21886] = a[13] & g[13694];
assign g[30077] = b[13] & g[13694];
assign g[21887] = a[13] & g[13695];
assign g[30078] = b[13] & g[13695];
assign g[21888] = a[13] & g[13696];
assign g[30079] = b[13] & g[13696];
assign g[21889] = a[13] & g[13697];
assign g[30080] = b[13] & g[13697];
assign g[21890] = a[13] & g[13698];
assign g[30081] = b[13] & g[13698];
assign g[21891] = a[13] & g[13699];
assign g[30082] = b[13] & g[13699];
assign g[21892] = a[13] & g[13700];
assign g[30083] = b[13] & g[13700];
assign g[21893] = a[13] & g[13701];
assign g[30084] = b[13] & g[13701];
assign g[21894] = a[13] & g[13702];
assign g[30085] = b[13] & g[13702];
assign g[21895] = a[13] & g[13703];
assign g[30086] = b[13] & g[13703];
assign g[21896] = a[13] & g[13704];
assign g[30087] = b[13] & g[13704];
assign g[21897] = a[13] & g[13705];
assign g[30088] = b[13] & g[13705];
assign g[21898] = a[13] & g[13706];
assign g[30089] = b[13] & g[13706];
assign g[21899] = a[13] & g[13707];
assign g[30090] = b[13] & g[13707];
assign g[21900] = a[13] & g[13708];
assign g[30091] = b[13] & g[13708];
assign g[21901] = a[13] & g[13709];
assign g[30092] = b[13] & g[13709];
assign g[21902] = a[13] & g[13710];
assign g[30093] = b[13] & g[13710];
assign g[21903] = a[13] & g[13711];
assign g[30094] = b[13] & g[13711];
assign g[21904] = a[13] & g[13712];
assign g[30095] = b[13] & g[13712];
assign g[21905] = a[13] & g[13713];
assign g[30096] = b[13] & g[13713];
assign g[21906] = a[13] & g[13714];
assign g[30097] = b[13] & g[13714];
assign g[21907] = a[13] & g[13715];
assign g[30098] = b[13] & g[13715];
assign g[21908] = a[13] & g[13716];
assign g[30099] = b[13] & g[13716];
assign g[21909] = a[13] & g[13717];
assign g[30100] = b[13] & g[13717];
assign g[21910] = a[13] & g[13718];
assign g[30101] = b[13] & g[13718];
assign g[21911] = a[13] & g[13719];
assign g[30102] = b[13] & g[13719];
assign g[21912] = a[13] & g[13720];
assign g[30103] = b[13] & g[13720];
assign g[21913] = a[13] & g[13721];
assign g[30104] = b[13] & g[13721];
assign g[21914] = a[13] & g[13722];
assign g[30105] = b[13] & g[13722];
assign g[21915] = a[13] & g[13723];
assign g[30106] = b[13] & g[13723];
assign g[21916] = a[13] & g[13724];
assign g[30107] = b[13] & g[13724];
assign g[21917] = a[13] & g[13725];
assign g[30108] = b[13] & g[13725];
assign g[21918] = a[13] & g[13726];
assign g[30109] = b[13] & g[13726];
assign g[21919] = a[13] & g[13727];
assign g[30110] = b[13] & g[13727];
assign g[21920] = a[13] & g[13728];
assign g[30111] = b[13] & g[13728];
assign g[21921] = a[13] & g[13729];
assign g[30112] = b[13] & g[13729];
assign g[21922] = a[13] & g[13730];
assign g[30113] = b[13] & g[13730];
assign g[21923] = a[13] & g[13731];
assign g[30114] = b[13] & g[13731];
assign g[21924] = a[13] & g[13732];
assign g[30115] = b[13] & g[13732];
assign g[21925] = a[13] & g[13733];
assign g[30116] = b[13] & g[13733];
assign g[21926] = a[13] & g[13734];
assign g[30117] = b[13] & g[13734];
assign g[21927] = a[13] & g[13735];
assign g[30118] = b[13] & g[13735];
assign g[21928] = a[13] & g[13736];
assign g[30119] = b[13] & g[13736];
assign g[21929] = a[13] & g[13737];
assign g[30120] = b[13] & g[13737];
assign g[21930] = a[13] & g[13738];
assign g[30121] = b[13] & g[13738];
assign g[21931] = a[13] & g[13739];
assign g[30122] = b[13] & g[13739];
assign g[21932] = a[13] & g[13740];
assign g[30123] = b[13] & g[13740];
assign g[21933] = a[13] & g[13741];
assign g[30124] = b[13] & g[13741];
assign g[21934] = a[13] & g[13742];
assign g[30125] = b[13] & g[13742];
assign g[21935] = a[13] & g[13743];
assign g[30126] = b[13] & g[13743];
assign g[21936] = a[13] & g[13744];
assign g[30127] = b[13] & g[13744];
assign g[21937] = a[13] & g[13745];
assign g[30128] = b[13] & g[13745];
assign g[21938] = a[13] & g[13746];
assign g[30129] = b[13] & g[13746];
assign g[21939] = a[13] & g[13747];
assign g[30130] = b[13] & g[13747];
assign g[21940] = a[13] & g[13748];
assign g[30131] = b[13] & g[13748];
assign g[21941] = a[13] & g[13749];
assign g[30132] = b[13] & g[13749];
assign g[21942] = a[13] & g[13750];
assign g[30133] = b[13] & g[13750];
assign g[21943] = a[13] & g[13751];
assign g[30134] = b[13] & g[13751];
assign g[21944] = a[13] & g[13752];
assign g[30135] = b[13] & g[13752];
assign g[21945] = a[13] & g[13753];
assign g[30136] = b[13] & g[13753];
assign g[21946] = a[13] & g[13754];
assign g[30137] = b[13] & g[13754];
assign g[21947] = a[13] & g[13755];
assign g[30138] = b[13] & g[13755];
assign g[21948] = a[13] & g[13756];
assign g[30139] = b[13] & g[13756];
assign g[21949] = a[13] & g[13757];
assign g[30140] = b[13] & g[13757];
assign g[21950] = a[13] & g[13758];
assign g[30141] = b[13] & g[13758];
assign g[21951] = a[13] & g[13759];
assign g[30142] = b[13] & g[13759];
assign g[21952] = a[13] & g[13760];
assign g[30143] = b[13] & g[13760];
assign g[21953] = a[13] & g[13761];
assign g[30144] = b[13] & g[13761];
assign g[21954] = a[13] & g[13762];
assign g[30145] = b[13] & g[13762];
assign g[21955] = a[13] & g[13763];
assign g[30146] = b[13] & g[13763];
assign g[21956] = a[13] & g[13764];
assign g[30147] = b[13] & g[13764];
assign g[21957] = a[13] & g[13765];
assign g[30148] = b[13] & g[13765];
assign g[21958] = a[13] & g[13766];
assign g[30149] = b[13] & g[13766];
assign g[21959] = a[13] & g[13767];
assign g[30150] = b[13] & g[13767];
assign g[21960] = a[13] & g[13768];
assign g[30151] = b[13] & g[13768];
assign g[21961] = a[13] & g[13769];
assign g[30152] = b[13] & g[13769];
assign g[21962] = a[13] & g[13770];
assign g[30153] = b[13] & g[13770];
assign g[21963] = a[13] & g[13771];
assign g[30154] = b[13] & g[13771];
assign g[21964] = a[13] & g[13772];
assign g[30155] = b[13] & g[13772];
assign g[21965] = a[13] & g[13773];
assign g[30156] = b[13] & g[13773];
assign g[21966] = a[13] & g[13774];
assign g[30157] = b[13] & g[13774];
assign g[21967] = a[13] & g[13775];
assign g[30158] = b[13] & g[13775];
assign g[21968] = a[13] & g[13776];
assign g[30159] = b[13] & g[13776];
assign g[21969] = a[13] & g[13777];
assign g[30160] = b[13] & g[13777];
assign g[21970] = a[13] & g[13778];
assign g[30161] = b[13] & g[13778];
assign g[21971] = a[13] & g[13779];
assign g[30162] = b[13] & g[13779];
assign g[21972] = a[13] & g[13780];
assign g[30163] = b[13] & g[13780];
assign g[21973] = a[13] & g[13781];
assign g[30164] = b[13] & g[13781];
assign g[21974] = a[13] & g[13782];
assign g[30165] = b[13] & g[13782];
assign g[21975] = a[13] & g[13783];
assign g[30166] = b[13] & g[13783];
assign g[21976] = a[13] & g[13784];
assign g[30167] = b[13] & g[13784];
assign g[21977] = a[13] & g[13785];
assign g[30168] = b[13] & g[13785];
assign g[21978] = a[13] & g[13786];
assign g[30169] = b[13] & g[13786];
assign g[21979] = a[13] & g[13787];
assign g[30170] = b[13] & g[13787];
assign g[21980] = a[13] & g[13788];
assign g[30171] = b[13] & g[13788];
assign g[21981] = a[13] & g[13789];
assign g[30172] = b[13] & g[13789];
assign g[21982] = a[13] & g[13790];
assign g[30173] = b[13] & g[13790];
assign g[21983] = a[13] & g[13791];
assign g[30174] = b[13] & g[13791];
assign g[21984] = a[13] & g[13792];
assign g[30175] = b[13] & g[13792];
assign g[21985] = a[13] & g[13793];
assign g[30176] = b[13] & g[13793];
assign g[21986] = a[13] & g[13794];
assign g[30177] = b[13] & g[13794];
assign g[21987] = a[13] & g[13795];
assign g[30178] = b[13] & g[13795];
assign g[21988] = a[13] & g[13796];
assign g[30179] = b[13] & g[13796];
assign g[21989] = a[13] & g[13797];
assign g[30180] = b[13] & g[13797];
assign g[21990] = a[13] & g[13798];
assign g[30181] = b[13] & g[13798];
assign g[21991] = a[13] & g[13799];
assign g[30182] = b[13] & g[13799];
assign g[21992] = a[13] & g[13800];
assign g[30183] = b[13] & g[13800];
assign g[21993] = a[13] & g[13801];
assign g[30184] = b[13] & g[13801];
assign g[21994] = a[13] & g[13802];
assign g[30185] = b[13] & g[13802];
assign g[21995] = a[13] & g[13803];
assign g[30186] = b[13] & g[13803];
assign g[21996] = a[13] & g[13804];
assign g[30187] = b[13] & g[13804];
assign g[21997] = a[13] & g[13805];
assign g[30188] = b[13] & g[13805];
assign g[21998] = a[13] & g[13806];
assign g[30189] = b[13] & g[13806];
assign g[21999] = a[13] & g[13807];
assign g[30190] = b[13] & g[13807];
assign g[22000] = a[13] & g[13808];
assign g[30191] = b[13] & g[13808];
assign g[22001] = a[13] & g[13809];
assign g[30192] = b[13] & g[13809];
assign g[22002] = a[13] & g[13810];
assign g[30193] = b[13] & g[13810];
assign g[22003] = a[13] & g[13811];
assign g[30194] = b[13] & g[13811];
assign g[22004] = a[13] & g[13812];
assign g[30195] = b[13] & g[13812];
assign g[22005] = a[13] & g[13813];
assign g[30196] = b[13] & g[13813];
assign g[22006] = a[13] & g[13814];
assign g[30197] = b[13] & g[13814];
assign g[22007] = a[13] & g[13815];
assign g[30198] = b[13] & g[13815];
assign g[22008] = a[13] & g[13816];
assign g[30199] = b[13] & g[13816];
assign g[22009] = a[13] & g[13817];
assign g[30200] = b[13] & g[13817];
assign g[22010] = a[13] & g[13818];
assign g[30201] = b[13] & g[13818];
assign g[22011] = a[13] & g[13819];
assign g[30202] = b[13] & g[13819];
assign g[22012] = a[13] & g[13820];
assign g[30203] = b[13] & g[13820];
assign g[22013] = a[13] & g[13821];
assign g[30204] = b[13] & g[13821];
assign g[22014] = a[13] & g[13822];
assign g[30205] = b[13] & g[13822];
assign g[22015] = a[13] & g[13823];
assign g[30206] = b[13] & g[13823];
assign g[22016] = a[13] & g[13824];
assign g[30207] = b[13] & g[13824];
assign g[22017] = a[13] & g[13825];
assign g[30208] = b[13] & g[13825];
assign g[22018] = a[13] & g[13826];
assign g[30209] = b[13] & g[13826];
assign g[22019] = a[13] & g[13827];
assign g[30210] = b[13] & g[13827];
assign g[22020] = a[13] & g[13828];
assign g[30211] = b[13] & g[13828];
assign g[22021] = a[13] & g[13829];
assign g[30212] = b[13] & g[13829];
assign g[22022] = a[13] & g[13830];
assign g[30213] = b[13] & g[13830];
assign g[22023] = a[13] & g[13831];
assign g[30214] = b[13] & g[13831];
assign g[22024] = a[13] & g[13832];
assign g[30215] = b[13] & g[13832];
assign g[22025] = a[13] & g[13833];
assign g[30216] = b[13] & g[13833];
assign g[22026] = a[13] & g[13834];
assign g[30217] = b[13] & g[13834];
assign g[22027] = a[13] & g[13835];
assign g[30218] = b[13] & g[13835];
assign g[22028] = a[13] & g[13836];
assign g[30219] = b[13] & g[13836];
assign g[22029] = a[13] & g[13837];
assign g[30220] = b[13] & g[13837];
assign g[22030] = a[13] & g[13838];
assign g[30221] = b[13] & g[13838];
assign g[22031] = a[13] & g[13839];
assign g[30222] = b[13] & g[13839];
assign g[22032] = a[13] & g[13840];
assign g[30223] = b[13] & g[13840];
assign g[22033] = a[13] & g[13841];
assign g[30224] = b[13] & g[13841];
assign g[22034] = a[13] & g[13842];
assign g[30225] = b[13] & g[13842];
assign g[22035] = a[13] & g[13843];
assign g[30226] = b[13] & g[13843];
assign g[22036] = a[13] & g[13844];
assign g[30227] = b[13] & g[13844];
assign g[22037] = a[13] & g[13845];
assign g[30228] = b[13] & g[13845];
assign g[22038] = a[13] & g[13846];
assign g[30229] = b[13] & g[13846];
assign g[22039] = a[13] & g[13847];
assign g[30230] = b[13] & g[13847];
assign g[22040] = a[13] & g[13848];
assign g[30231] = b[13] & g[13848];
assign g[22041] = a[13] & g[13849];
assign g[30232] = b[13] & g[13849];
assign g[22042] = a[13] & g[13850];
assign g[30233] = b[13] & g[13850];
assign g[22043] = a[13] & g[13851];
assign g[30234] = b[13] & g[13851];
assign g[22044] = a[13] & g[13852];
assign g[30235] = b[13] & g[13852];
assign g[22045] = a[13] & g[13853];
assign g[30236] = b[13] & g[13853];
assign g[22046] = a[13] & g[13854];
assign g[30237] = b[13] & g[13854];
assign g[22047] = a[13] & g[13855];
assign g[30238] = b[13] & g[13855];
assign g[22048] = a[13] & g[13856];
assign g[30239] = b[13] & g[13856];
assign g[22049] = a[13] & g[13857];
assign g[30240] = b[13] & g[13857];
assign g[22050] = a[13] & g[13858];
assign g[30241] = b[13] & g[13858];
assign g[22051] = a[13] & g[13859];
assign g[30242] = b[13] & g[13859];
assign g[22052] = a[13] & g[13860];
assign g[30243] = b[13] & g[13860];
assign g[22053] = a[13] & g[13861];
assign g[30244] = b[13] & g[13861];
assign g[22054] = a[13] & g[13862];
assign g[30245] = b[13] & g[13862];
assign g[22055] = a[13] & g[13863];
assign g[30246] = b[13] & g[13863];
assign g[22056] = a[13] & g[13864];
assign g[30247] = b[13] & g[13864];
assign g[22057] = a[13] & g[13865];
assign g[30248] = b[13] & g[13865];
assign g[22058] = a[13] & g[13866];
assign g[30249] = b[13] & g[13866];
assign g[22059] = a[13] & g[13867];
assign g[30250] = b[13] & g[13867];
assign g[22060] = a[13] & g[13868];
assign g[30251] = b[13] & g[13868];
assign g[22061] = a[13] & g[13869];
assign g[30252] = b[13] & g[13869];
assign g[22062] = a[13] & g[13870];
assign g[30253] = b[13] & g[13870];
assign g[22063] = a[13] & g[13871];
assign g[30254] = b[13] & g[13871];
assign g[22064] = a[13] & g[13872];
assign g[30255] = b[13] & g[13872];
assign g[22065] = a[13] & g[13873];
assign g[30256] = b[13] & g[13873];
assign g[22066] = a[13] & g[13874];
assign g[30257] = b[13] & g[13874];
assign g[22067] = a[13] & g[13875];
assign g[30258] = b[13] & g[13875];
assign g[22068] = a[13] & g[13876];
assign g[30259] = b[13] & g[13876];
assign g[22069] = a[13] & g[13877];
assign g[30260] = b[13] & g[13877];
assign g[22070] = a[13] & g[13878];
assign g[30261] = b[13] & g[13878];
assign g[22071] = a[13] & g[13879];
assign g[30262] = b[13] & g[13879];
assign g[22072] = a[13] & g[13880];
assign g[30263] = b[13] & g[13880];
assign g[22073] = a[13] & g[13881];
assign g[30264] = b[13] & g[13881];
assign g[22074] = a[13] & g[13882];
assign g[30265] = b[13] & g[13882];
assign g[22075] = a[13] & g[13883];
assign g[30266] = b[13] & g[13883];
assign g[22076] = a[13] & g[13884];
assign g[30267] = b[13] & g[13884];
assign g[22077] = a[13] & g[13885];
assign g[30268] = b[13] & g[13885];
assign g[22078] = a[13] & g[13886];
assign g[30269] = b[13] & g[13886];
assign g[22079] = a[13] & g[13887];
assign g[30270] = b[13] & g[13887];
assign g[22080] = a[13] & g[13888];
assign g[30271] = b[13] & g[13888];
assign g[22081] = a[13] & g[13889];
assign g[30272] = b[13] & g[13889];
assign g[22082] = a[13] & g[13890];
assign g[30273] = b[13] & g[13890];
assign g[22083] = a[13] & g[13891];
assign g[30274] = b[13] & g[13891];
assign g[22084] = a[13] & g[13892];
assign g[30275] = b[13] & g[13892];
assign g[22085] = a[13] & g[13893];
assign g[30276] = b[13] & g[13893];
assign g[22086] = a[13] & g[13894];
assign g[30277] = b[13] & g[13894];
assign g[22087] = a[13] & g[13895];
assign g[30278] = b[13] & g[13895];
assign g[22088] = a[13] & g[13896];
assign g[30279] = b[13] & g[13896];
assign g[22089] = a[13] & g[13897];
assign g[30280] = b[13] & g[13897];
assign g[22090] = a[13] & g[13898];
assign g[30281] = b[13] & g[13898];
assign g[22091] = a[13] & g[13899];
assign g[30282] = b[13] & g[13899];
assign g[22092] = a[13] & g[13900];
assign g[30283] = b[13] & g[13900];
assign g[22093] = a[13] & g[13901];
assign g[30284] = b[13] & g[13901];
assign g[22094] = a[13] & g[13902];
assign g[30285] = b[13] & g[13902];
assign g[22095] = a[13] & g[13903];
assign g[30286] = b[13] & g[13903];
assign g[22096] = a[13] & g[13904];
assign g[30287] = b[13] & g[13904];
assign g[22097] = a[13] & g[13905];
assign g[30288] = b[13] & g[13905];
assign g[22098] = a[13] & g[13906];
assign g[30289] = b[13] & g[13906];
assign g[22099] = a[13] & g[13907];
assign g[30290] = b[13] & g[13907];
assign g[22100] = a[13] & g[13908];
assign g[30291] = b[13] & g[13908];
assign g[22101] = a[13] & g[13909];
assign g[30292] = b[13] & g[13909];
assign g[22102] = a[13] & g[13910];
assign g[30293] = b[13] & g[13910];
assign g[22103] = a[13] & g[13911];
assign g[30294] = b[13] & g[13911];
assign g[22104] = a[13] & g[13912];
assign g[30295] = b[13] & g[13912];
assign g[22105] = a[13] & g[13913];
assign g[30296] = b[13] & g[13913];
assign g[22106] = a[13] & g[13914];
assign g[30297] = b[13] & g[13914];
assign g[22107] = a[13] & g[13915];
assign g[30298] = b[13] & g[13915];
assign g[22108] = a[13] & g[13916];
assign g[30299] = b[13] & g[13916];
assign g[22109] = a[13] & g[13917];
assign g[30300] = b[13] & g[13917];
assign g[22110] = a[13] & g[13918];
assign g[30301] = b[13] & g[13918];
assign g[22111] = a[13] & g[13919];
assign g[30302] = b[13] & g[13919];
assign g[22112] = a[13] & g[13920];
assign g[30303] = b[13] & g[13920];
assign g[22113] = a[13] & g[13921];
assign g[30304] = b[13] & g[13921];
assign g[22114] = a[13] & g[13922];
assign g[30305] = b[13] & g[13922];
assign g[22115] = a[13] & g[13923];
assign g[30306] = b[13] & g[13923];
assign g[22116] = a[13] & g[13924];
assign g[30307] = b[13] & g[13924];
assign g[22117] = a[13] & g[13925];
assign g[30308] = b[13] & g[13925];
assign g[22118] = a[13] & g[13926];
assign g[30309] = b[13] & g[13926];
assign g[22119] = a[13] & g[13927];
assign g[30310] = b[13] & g[13927];
assign g[22120] = a[13] & g[13928];
assign g[30311] = b[13] & g[13928];
assign g[22121] = a[13] & g[13929];
assign g[30312] = b[13] & g[13929];
assign g[22122] = a[13] & g[13930];
assign g[30313] = b[13] & g[13930];
assign g[22123] = a[13] & g[13931];
assign g[30314] = b[13] & g[13931];
assign g[22124] = a[13] & g[13932];
assign g[30315] = b[13] & g[13932];
assign g[22125] = a[13] & g[13933];
assign g[30316] = b[13] & g[13933];
assign g[22126] = a[13] & g[13934];
assign g[30317] = b[13] & g[13934];
assign g[22127] = a[13] & g[13935];
assign g[30318] = b[13] & g[13935];
assign g[22128] = a[13] & g[13936];
assign g[30319] = b[13] & g[13936];
assign g[22129] = a[13] & g[13937];
assign g[30320] = b[13] & g[13937];
assign g[22130] = a[13] & g[13938];
assign g[30321] = b[13] & g[13938];
assign g[22131] = a[13] & g[13939];
assign g[30322] = b[13] & g[13939];
assign g[22132] = a[13] & g[13940];
assign g[30323] = b[13] & g[13940];
assign g[22133] = a[13] & g[13941];
assign g[30324] = b[13] & g[13941];
assign g[22134] = a[13] & g[13942];
assign g[30325] = b[13] & g[13942];
assign g[22135] = a[13] & g[13943];
assign g[30326] = b[13] & g[13943];
assign g[22136] = a[13] & g[13944];
assign g[30327] = b[13] & g[13944];
assign g[22137] = a[13] & g[13945];
assign g[30328] = b[13] & g[13945];
assign g[22138] = a[13] & g[13946];
assign g[30329] = b[13] & g[13946];
assign g[22139] = a[13] & g[13947];
assign g[30330] = b[13] & g[13947];
assign g[22140] = a[13] & g[13948];
assign g[30331] = b[13] & g[13948];
assign g[22141] = a[13] & g[13949];
assign g[30332] = b[13] & g[13949];
assign g[22142] = a[13] & g[13950];
assign g[30333] = b[13] & g[13950];
assign g[22143] = a[13] & g[13951];
assign g[30334] = b[13] & g[13951];
assign g[22144] = a[13] & g[13952];
assign g[30335] = b[13] & g[13952];
assign g[22145] = a[13] & g[13953];
assign g[30336] = b[13] & g[13953];
assign g[22146] = a[13] & g[13954];
assign g[30337] = b[13] & g[13954];
assign g[22147] = a[13] & g[13955];
assign g[30338] = b[13] & g[13955];
assign g[22148] = a[13] & g[13956];
assign g[30339] = b[13] & g[13956];
assign g[22149] = a[13] & g[13957];
assign g[30340] = b[13] & g[13957];
assign g[22150] = a[13] & g[13958];
assign g[30341] = b[13] & g[13958];
assign g[22151] = a[13] & g[13959];
assign g[30342] = b[13] & g[13959];
assign g[22152] = a[13] & g[13960];
assign g[30343] = b[13] & g[13960];
assign g[22153] = a[13] & g[13961];
assign g[30344] = b[13] & g[13961];
assign g[22154] = a[13] & g[13962];
assign g[30345] = b[13] & g[13962];
assign g[22155] = a[13] & g[13963];
assign g[30346] = b[13] & g[13963];
assign g[22156] = a[13] & g[13964];
assign g[30347] = b[13] & g[13964];
assign g[22157] = a[13] & g[13965];
assign g[30348] = b[13] & g[13965];
assign g[22158] = a[13] & g[13966];
assign g[30349] = b[13] & g[13966];
assign g[22159] = a[13] & g[13967];
assign g[30350] = b[13] & g[13967];
assign g[22160] = a[13] & g[13968];
assign g[30351] = b[13] & g[13968];
assign g[22161] = a[13] & g[13969];
assign g[30352] = b[13] & g[13969];
assign g[22162] = a[13] & g[13970];
assign g[30353] = b[13] & g[13970];
assign g[22163] = a[13] & g[13971];
assign g[30354] = b[13] & g[13971];
assign g[22164] = a[13] & g[13972];
assign g[30355] = b[13] & g[13972];
assign g[22165] = a[13] & g[13973];
assign g[30356] = b[13] & g[13973];
assign g[22166] = a[13] & g[13974];
assign g[30357] = b[13] & g[13974];
assign g[22167] = a[13] & g[13975];
assign g[30358] = b[13] & g[13975];
assign g[22168] = a[13] & g[13976];
assign g[30359] = b[13] & g[13976];
assign g[22169] = a[13] & g[13977];
assign g[30360] = b[13] & g[13977];
assign g[22170] = a[13] & g[13978];
assign g[30361] = b[13] & g[13978];
assign g[22171] = a[13] & g[13979];
assign g[30362] = b[13] & g[13979];
assign g[22172] = a[13] & g[13980];
assign g[30363] = b[13] & g[13980];
assign g[22173] = a[13] & g[13981];
assign g[30364] = b[13] & g[13981];
assign g[22174] = a[13] & g[13982];
assign g[30365] = b[13] & g[13982];
assign g[22175] = a[13] & g[13983];
assign g[30366] = b[13] & g[13983];
assign g[22176] = a[13] & g[13984];
assign g[30367] = b[13] & g[13984];
assign g[22177] = a[13] & g[13985];
assign g[30368] = b[13] & g[13985];
assign g[22178] = a[13] & g[13986];
assign g[30369] = b[13] & g[13986];
assign g[22179] = a[13] & g[13987];
assign g[30370] = b[13] & g[13987];
assign g[22180] = a[13] & g[13988];
assign g[30371] = b[13] & g[13988];
assign g[22181] = a[13] & g[13989];
assign g[30372] = b[13] & g[13989];
assign g[22182] = a[13] & g[13990];
assign g[30373] = b[13] & g[13990];
assign g[22183] = a[13] & g[13991];
assign g[30374] = b[13] & g[13991];
assign g[22184] = a[13] & g[13992];
assign g[30375] = b[13] & g[13992];
assign g[22185] = a[13] & g[13993];
assign g[30376] = b[13] & g[13993];
assign g[22186] = a[13] & g[13994];
assign g[30377] = b[13] & g[13994];
assign g[22187] = a[13] & g[13995];
assign g[30378] = b[13] & g[13995];
assign g[22188] = a[13] & g[13996];
assign g[30379] = b[13] & g[13996];
assign g[22189] = a[13] & g[13997];
assign g[30380] = b[13] & g[13997];
assign g[22190] = a[13] & g[13998];
assign g[30381] = b[13] & g[13998];
assign g[22191] = a[13] & g[13999];
assign g[30382] = b[13] & g[13999];
assign g[22192] = a[13] & g[14000];
assign g[30383] = b[13] & g[14000];
assign g[22193] = a[13] & g[14001];
assign g[30384] = b[13] & g[14001];
assign g[22194] = a[13] & g[14002];
assign g[30385] = b[13] & g[14002];
assign g[22195] = a[13] & g[14003];
assign g[30386] = b[13] & g[14003];
assign g[22196] = a[13] & g[14004];
assign g[30387] = b[13] & g[14004];
assign g[22197] = a[13] & g[14005];
assign g[30388] = b[13] & g[14005];
assign g[22198] = a[13] & g[14006];
assign g[30389] = b[13] & g[14006];
assign g[22199] = a[13] & g[14007];
assign g[30390] = b[13] & g[14007];
assign g[22200] = a[13] & g[14008];
assign g[30391] = b[13] & g[14008];
assign g[22201] = a[13] & g[14009];
assign g[30392] = b[13] & g[14009];
assign g[22202] = a[13] & g[14010];
assign g[30393] = b[13] & g[14010];
assign g[22203] = a[13] & g[14011];
assign g[30394] = b[13] & g[14011];
assign g[22204] = a[13] & g[14012];
assign g[30395] = b[13] & g[14012];
assign g[22205] = a[13] & g[14013];
assign g[30396] = b[13] & g[14013];
assign g[22206] = a[13] & g[14014];
assign g[30397] = b[13] & g[14014];
assign g[22207] = a[13] & g[14015];
assign g[30398] = b[13] & g[14015];
assign g[22208] = a[13] & g[14016];
assign g[30399] = b[13] & g[14016];
assign g[22209] = a[13] & g[14017];
assign g[30400] = b[13] & g[14017];
assign g[22210] = a[13] & g[14018];
assign g[30401] = b[13] & g[14018];
assign g[22211] = a[13] & g[14019];
assign g[30402] = b[13] & g[14019];
assign g[22212] = a[13] & g[14020];
assign g[30403] = b[13] & g[14020];
assign g[22213] = a[13] & g[14021];
assign g[30404] = b[13] & g[14021];
assign g[22214] = a[13] & g[14022];
assign g[30405] = b[13] & g[14022];
assign g[22215] = a[13] & g[14023];
assign g[30406] = b[13] & g[14023];
assign g[22216] = a[13] & g[14024];
assign g[30407] = b[13] & g[14024];
assign g[22217] = a[13] & g[14025];
assign g[30408] = b[13] & g[14025];
assign g[22218] = a[13] & g[14026];
assign g[30409] = b[13] & g[14026];
assign g[22219] = a[13] & g[14027];
assign g[30410] = b[13] & g[14027];
assign g[22220] = a[13] & g[14028];
assign g[30411] = b[13] & g[14028];
assign g[22221] = a[13] & g[14029];
assign g[30412] = b[13] & g[14029];
assign g[22222] = a[13] & g[14030];
assign g[30413] = b[13] & g[14030];
assign g[22223] = a[13] & g[14031];
assign g[30414] = b[13] & g[14031];
assign g[22224] = a[13] & g[14032];
assign g[30415] = b[13] & g[14032];
assign g[22225] = a[13] & g[14033];
assign g[30416] = b[13] & g[14033];
assign g[22226] = a[13] & g[14034];
assign g[30417] = b[13] & g[14034];
assign g[22227] = a[13] & g[14035];
assign g[30418] = b[13] & g[14035];
assign g[22228] = a[13] & g[14036];
assign g[30419] = b[13] & g[14036];
assign g[22229] = a[13] & g[14037];
assign g[30420] = b[13] & g[14037];
assign g[22230] = a[13] & g[14038];
assign g[30421] = b[13] & g[14038];
assign g[22231] = a[13] & g[14039];
assign g[30422] = b[13] & g[14039];
assign g[22232] = a[13] & g[14040];
assign g[30423] = b[13] & g[14040];
assign g[22233] = a[13] & g[14041];
assign g[30424] = b[13] & g[14041];
assign g[22234] = a[13] & g[14042];
assign g[30425] = b[13] & g[14042];
assign g[22235] = a[13] & g[14043];
assign g[30426] = b[13] & g[14043];
assign g[22236] = a[13] & g[14044];
assign g[30427] = b[13] & g[14044];
assign g[22237] = a[13] & g[14045];
assign g[30428] = b[13] & g[14045];
assign g[22238] = a[13] & g[14046];
assign g[30429] = b[13] & g[14046];
assign g[22239] = a[13] & g[14047];
assign g[30430] = b[13] & g[14047];
assign g[22240] = a[13] & g[14048];
assign g[30431] = b[13] & g[14048];
assign g[22241] = a[13] & g[14049];
assign g[30432] = b[13] & g[14049];
assign g[22242] = a[13] & g[14050];
assign g[30433] = b[13] & g[14050];
assign g[22243] = a[13] & g[14051];
assign g[30434] = b[13] & g[14051];
assign g[22244] = a[13] & g[14052];
assign g[30435] = b[13] & g[14052];
assign g[22245] = a[13] & g[14053];
assign g[30436] = b[13] & g[14053];
assign g[22246] = a[13] & g[14054];
assign g[30437] = b[13] & g[14054];
assign g[22247] = a[13] & g[14055];
assign g[30438] = b[13] & g[14055];
assign g[22248] = a[13] & g[14056];
assign g[30439] = b[13] & g[14056];
assign g[22249] = a[13] & g[14057];
assign g[30440] = b[13] & g[14057];
assign g[22250] = a[13] & g[14058];
assign g[30441] = b[13] & g[14058];
assign g[22251] = a[13] & g[14059];
assign g[30442] = b[13] & g[14059];
assign g[22252] = a[13] & g[14060];
assign g[30443] = b[13] & g[14060];
assign g[22253] = a[13] & g[14061];
assign g[30444] = b[13] & g[14061];
assign g[22254] = a[13] & g[14062];
assign g[30445] = b[13] & g[14062];
assign g[22255] = a[13] & g[14063];
assign g[30446] = b[13] & g[14063];
assign g[22256] = a[13] & g[14064];
assign g[30447] = b[13] & g[14064];
assign g[22257] = a[13] & g[14065];
assign g[30448] = b[13] & g[14065];
assign g[22258] = a[13] & g[14066];
assign g[30449] = b[13] & g[14066];
assign g[22259] = a[13] & g[14067];
assign g[30450] = b[13] & g[14067];
assign g[22260] = a[13] & g[14068];
assign g[30451] = b[13] & g[14068];
assign g[22261] = a[13] & g[14069];
assign g[30452] = b[13] & g[14069];
assign g[22262] = a[13] & g[14070];
assign g[30453] = b[13] & g[14070];
assign g[22263] = a[13] & g[14071];
assign g[30454] = b[13] & g[14071];
assign g[22264] = a[13] & g[14072];
assign g[30455] = b[13] & g[14072];
assign g[22265] = a[13] & g[14073];
assign g[30456] = b[13] & g[14073];
assign g[22266] = a[13] & g[14074];
assign g[30457] = b[13] & g[14074];
assign g[22267] = a[13] & g[14075];
assign g[30458] = b[13] & g[14075];
assign g[22268] = a[13] & g[14076];
assign g[30459] = b[13] & g[14076];
assign g[22269] = a[13] & g[14077];
assign g[30460] = b[13] & g[14077];
assign g[22270] = a[13] & g[14078];
assign g[30461] = b[13] & g[14078];
assign g[22271] = a[13] & g[14079];
assign g[30462] = b[13] & g[14079];
assign g[22272] = a[13] & g[14080];
assign g[30463] = b[13] & g[14080];
assign g[22273] = a[13] & g[14081];
assign g[30464] = b[13] & g[14081];
assign g[22274] = a[13] & g[14082];
assign g[30465] = b[13] & g[14082];
assign g[22275] = a[13] & g[14083];
assign g[30466] = b[13] & g[14083];
assign g[22276] = a[13] & g[14084];
assign g[30467] = b[13] & g[14084];
assign g[22277] = a[13] & g[14085];
assign g[30468] = b[13] & g[14085];
assign g[22278] = a[13] & g[14086];
assign g[30469] = b[13] & g[14086];
assign g[22279] = a[13] & g[14087];
assign g[30470] = b[13] & g[14087];
assign g[22280] = a[13] & g[14088];
assign g[30471] = b[13] & g[14088];
assign g[22281] = a[13] & g[14089];
assign g[30472] = b[13] & g[14089];
assign g[22282] = a[13] & g[14090];
assign g[30473] = b[13] & g[14090];
assign g[22283] = a[13] & g[14091];
assign g[30474] = b[13] & g[14091];
assign g[22284] = a[13] & g[14092];
assign g[30475] = b[13] & g[14092];
assign g[22285] = a[13] & g[14093];
assign g[30476] = b[13] & g[14093];
assign g[22286] = a[13] & g[14094];
assign g[30477] = b[13] & g[14094];
assign g[22287] = a[13] & g[14095];
assign g[30478] = b[13] & g[14095];
assign g[22288] = a[13] & g[14096];
assign g[30479] = b[13] & g[14096];
assign g[22289] = a[13] & g[14097];
assign g[30480] = b[13] & g[14097];
assign g[22290] = a[13] & g[14098];
assign g[30481] = b[13] & g[14098];
assign g[22291] = a[13] & g[14099];
assign g[30482] = b[13] & g[14099];
assign g[22292] = a[13] & g[14100];
assign g[30483] = b[13] & g[14100];
assign g[22293] = a[13] & g[14101];
assign g[30484] = b[13] & g[14101];
assign g[22294] = a[13] & g[14102];
assign g[30485] = b[13] & g[14102];
assign g[22295] = a[13] & g[14103];
assign g[30486] = b[13] & g[14103];
assign g[22296] = a[13] & g[14104];
assign g[30487] = b[13] & g[14104];
assign g[22297] = a[13] & g[14105];
assign g[30488] = b[13] & g[14105];
assign g[22298] = a[13] & g[14106];
assign g[30489] = b[13] & g[14106];
assign g[22299] = a[13] & g[14107];
assign g[30490] = b[13] & g[14107];
assign g[22300] = a[13] & g[14108];
assign g[30491] = b[13] & g[14108];
assign g[22301] = a[13] & g[14109];
assign g[30492] = b[13] & g[14109];
assign g[22302] = a[13] & g[14110];
assign g[30493] = b[13] & g[14110];
assign g[22303] = a[13] & g[14111];
assign g[30494] = b[13] & g[14111];
assign g[22304] = a[13] & g[14112];
assign g[30495] = b[13] & g[14112];
assign g[22305] = a[13] & g[14113];
assign g[30496] = b[13] & g[14113];
assign g[22306] = a[13] & g[14114];
assign g[30497] = b[13] & g[14114];
assign g[22307] = a[13] & g[14115];
assign g[30498] = b[13] & g[14115];
assign g[22308] = a[13] & g[14116];
assign g[30499] = b[13] & g[14116];
assign g[22309] = a[13] & g[14117];
assign g[30500] = b[13] & g[14117];
assign g[22310] = a[13] & g[14118];
assign g[30501] = b[13] & g[14118];
assign g[22311] = a[13] & g[14119];
assign g[30502] = b[13] & g[14119];
assign g[22312] = a[13] & g[14120];
assign g[30503] = b[13] & g[14120];
assign g[22313] = a[13] & g[14121];
assign g[30504] = b[13] & g[14121];
assign g[22314] = a[13] & g[14122];
assign g[30505] = b[13] & g[14122];
assign g[22315] = a[13] & g[14123];
assign g[30506] = b[13] & g[14123];
assign g[22316] = a[13] & g[14124];
assign g[30507] = b[13] & g[14124];
assign g[22317] = a[13] & g[14125];
assign g[30508] = b[13] & g[14125];
assign g[22318] = a[13] & g[14126];
assign g[30509] = b[13] & g[14126];
assign g[22319] = a[13] & g[14127];
assign g[30510] = b[13] & g[14127];
assign g[22320] = a[13] & g[14128];
assign g[30511] = b[13] & g[14128];
assign g[22321] = a[13] & g[14129];
assign g[30512] = b[13] & g[14129];
assign g[22322] = a[13] & g[14130];
assign g[30513] = b[13] & g[14130];
assign g[22323] = a[13] & g[14131];
assign g[30514] = b[13] & g[14131];
assign g[22324] = a[13] & g[14132];
assign g[30515] = b[13] & g[14132];
assign g[22325] = a[13] & g[14133];
assign g[30516] = b[13] & g[14133];
assign g[22326] = a[13] & g[14134];
assign g[30517] = b[13] & g[14134];
assign g[22327] = a[13] & g[14135];
assign g[30518] = b[13] & g[14135];
assign g[22328] = a[13] & g[14136];
assign g[30519] = b[13] & g[14136];
assign g[22329] = a[13] & g[14137];
assign g[30520] = b[13] & g[14137];
assign g[22330] = a[13] & g[14138];
assign g[30521] = b[13] & g[14138];
assign g[22331] = a[13] & g[14139];
assign g[30522] = b[13] & g[14139];
assign g[22332] = a[13] & g[14140];
assign g[30523] = b[13] & g[14140];
assign g[22333] = a[13] & g[14141];
assign g[30524] = b[13] & g[14141];
assign g[22334] = a[13] & g[14142];
assign g[30525] = b[13] & g[14142];
assign g[22335] = a[13] & g[14143];
assign g[30526] = b[13] & g[14143];
assign g[22336] = a[13] & g[14144];
assign g[30527] = b[13] & g[14144];
assign g[22337] = a[13] & g[14145];
assign g[30528] = b[13] & g[14145];
assign g[22338] = a[13] & g[14146];
assign g[30529] = b[13] & g[14146];
assign g[22339] = a[13] & g[14147];
assign g[30530] = b[13] & g[14147];
assign g[22340] = a[13] & g[14148];
assign g[30531] = b[13] & g[14148];
assign g[22341] = a[13] & g[14149];
assign g[30532] = b[13] & g[14149];
assign g[22342] = a[13] & g[14150];
assign g[30533] = b[13] & g[14150];
assign g[22343] = a[13] & g[14151];
assign g[30534] = b[13] & g[14151];
assign g[22344] = a[13] & g[14152];
assign g[30535] = b[13] & g[14152];
assign g[22345] = a[13] & g[14153];
assign g[30536] = b[13] & g[14153];
assign g[22346] = a[13] & g[14154];
assign g[30537] = b[13] & g[14154];
assign g[22347] = a[13] & g[14155];
assign g[30538] = b[13] & g[14155];
assign g[22348] = a[13] & g[14156];
assign g[30539] = b[13] & g[14156];
assign g[22349] = a[13] & g[14157];
assign g[30540] = b[13] & g[14157];
assign g[22350] = a[13] & g[14158];
assign g[30541] = b[13] & g[14158];
assign g[22351] = a[13] & g[14159];
assign g[30542] = b[13] & g[14159];
assign g[22352] = a[13] & g[14160];
assign g[30543] = b[13] & g[14160];
assign g[22353] = a[13] & g[14161];
assign g[30544] = b[13] & g[14161];
assign g[22354] = a[13] & g[14162];
assign g[30545] = b[13] & g[14162];
assign g[22355] = a[13] & g[14163];
assign g[30546] = b[13] & g[14163];
assign g[22356] = a[13] & g[14164];
assign g[30547] = b[13] & g[14164];
assign g[22357] = a[13] & g[14165];
assign g[30548] = b[13] & g[14165];
assign g[22358] = a[13] & g[14166];
assign g[30549] = b[13] & g[14166];
assign g[22359] = a[13] & g[14167];
assign g[30550] = b[13] & g[14167];
assign g[22360] = a[13] & g[14168];
assign g[30551] = b[13] & g[14168];
assign g[22361] = a[13] & g[14169];
assign g[30552] = b[13] & g[14169];
assign g[22362] = a[13] & g[14170];
assign g[30553] = b[13] & g[14170];
assign g[22363] = a[13] & g[14171];
assign g[30554] = b[13] & g[14171];
assign g[22364] = a[13] & g[14172];
assign g[30555] = b[13] & g[14172];
assign g[22365] = a[13] & g[14173];
assign g[30556] = b[13] & g[14173];
assign g[22366] = a[13] & g[14174];
assign g[30557] = b[13] & g[14174];
assign g[22367] = a[13] & g[14175];
assign g[30558] = b[13] & g[14175];
assign g[22368] = a[13] & g[14176];
assign g[30559] = b[13] & g[14176];
assign g[22369] = a[13] & g[14177];
assign g[30560] = b[13] & g[14177];
assign g[22370] = a[13] & g[14178];
assign g[30561] = b[13] & g[14178];
assign g[22371] = a[13] & g[14179];
assign g[30562] = b[13] & g[14179];
assign g[22372] = a[13] & g[14180];
assign g[30563] = b[13] & g[14180];
assign g[22373] = a[13] & g[14181];
assign g[30564] = b[13] & g[14181];
assign g[22374] = a[13] & g[14182];
assign g[30565] = b[13] & g[14182];
assign g[22375] = a[13] & g[14183];
assign g[30566] = b[13] & g[14183];
assign g[22376] = a[13] & g[14184];
assign g[30567] = b[13] & g[14184];
assign g[22377] = a[13] & g[14185];
assign g[30568] = b[13] & g[14185];
assign g[22378] = a[13] & g[14186];
assign g[30569] = b[13] & g[14186];
assign g[22379] = a[13] & g[14187];
assign g[30570] = b[13] & g[14187];
assign g[22380] = a[13] & g[14188];
assign g[30571] = b[13] & g[14188];
assign g[22381] = a[13] & g[14189];
assign g[30572] = b[13] & g[14189];
assign g[22382] = a[13] & g[14190];
assign g[30573] = b[13] & g[14190];
assign g[22383] = a[13] & g[14191];
assign g[30574] = b[13] & g[14191];
assign g[22384] = a[13] & g[14192];
assign g[30575] = b[13] & g[14192];
assign g[22385] = a[13] & g[14193];
assign g[30576] = b[13] & g[14193];
assign g[22386] = a[13] & g[14194];
assign g[30577] = b[13] & g[14194];
assign g[22387] = a[13] & g[14195];
assign g[30578] = b[13] & g[14195];
assign g[22388] = a[13] & g[14196];
assign g[30579] = b[13] & g[14196];
assign g[22389] = a[13] & g[14197];
assign g[30580] = b[13] & g[14197];
assign g[22390] = a[13] & g[14198];
assign g[30581] = b[13] & g[14198];
assign g[22391] = a[13] & g[14199];
assign g[30582] = b[13] & g[14199];
assign g[22392] = a[13] & g[14200];
assign g[30583] = b[13] & g[14200];
assign g[22393] = a[13] & g[14201];
assign g[30584] = b[13] & g[14201];
assign g[22394] = a[13] & g[14202];
assign g[30585] = b[13] & g[14202];
assign g[22395] = a[13] & g[14203];
assign g[30586] = b[13] & g[14203];
assign g[22396] = a[13] & g[14204];
assign g[30587] = b[13] & g[14204];
assign g[22397] = a[13] & g[14205];
assign g[30588] = b[13] & g[14205];
assign g[22398] = a[13] & g[14206];
assign g[30589] = b[13] & g[14206];
assign g[22399] = a[13] & g[14207];
assign g[30590] = b[13] & g[14207];
assign g[22400] = a[13] & g[14208];
assign g[30591] = b[13] & g[14208];
assign g[22401] = a[13] & g[14209];
assign g[30592] = b[13] & g[14209];
assign g[22402] = a[13] & g[14210];
assign g[30593] = b[13] & g[14210];
assign g[22403] = a[13] & g[14211];
assign g[30594] = b[13] & g[14211];
assign g[22404] = a[13] & g[14212];
assign g[30595] = b[13] & g[14212];
assign g[22405] = a[13] & g[14213];
assign g[30596] = b[13] & g[14213];
assign g[22406] = a[13] & g[14214];
assign g[30597] = b[13] & g[14214];
assign g[22407] = a[13] & g[14215];
assign g[30598] = b[13] & g[14215];
assign g[22408] = a[13] & g[14216];
assign g[30599] = b[13] & g[14216];
assign g[22409] = a[13] & g[14217];
assign g[30600] = b[13] & g[14217];
assign g[22410] = a[13] & g[14218];
assign g[30601] = b[13] & g[14218];
assign g[22411] = a[13] & g[14219];
assign g[30602] = b[13] & g[14219];
assign g[22412] = a[13] & g[14220];
assign g[30603] = b[13] & g[14220];
assign g[22413] = a[13] & g[14221];
assign g[30604] = b[13] & g[14221];
assign g[22414] = a[13] & g[14222];
assign g[30605] = b[13] & g[14222];
assign g[22415] = a[13] & g[14223];
assign g[30606] = b[13] & g[14223];
assign g[22416] = a[13] & g[14224];
assign g[30607] = b[13] & g[14224];
assign g[22417] = a[13] & g[14225];
assign g[30608] = b[13] & g[14225];
assign g[22418] = a[13] & g[14226];
assign g[30609] = b[13] & g[14226];
assign g[22419] = a[13] & g[14227];
assign g[30610] = b[13] & g[14227];
assign g[22420] = a[13] & g[14228];
assign g[30611] = b[13] & g[14228];
assign g[22421] = a[13] & g[14229];
assign g[30612] = b[13] & g[14229];
assign g[22422] = a[13] & g[14230];
assign g[30613] = b[13] & g[14230];
assign g[22423] = a[13] & g[14231];
assign g[30614] = b[13] & g[14231];
assign g[22424] = a[13] & g[14232];
assign g[30615] = b[13] & g[14232];
assign g[22425] = a[13] & g[14233];
assign g[30616] = b[13] & g[14233];
assign g[22426] = a[13] & g[14234];
assign g[30617] = b[13] & g[14234];
assign g[22427] = a[13] & g[14235];
assign g[30618] = b[13] & g[14235];
assign g[22428] = a[13] & g[14236];
assign g[30619] = b[13] & g[14236];
assign g[22429] = a[13] & g[14237];
assign g[30620] = b[13] & g[14237];
assign g[22430] = a[13] & g[14238];
assign g[30621] = b[13] & g[14238];
assign g[22431] = a[13] & g[14239];
assign g[30622] = b[13] & g[14239];
assign g[22432] = a[13] & g[14240];
assign g[30623] = b[13] & g[14240];
assign g[22433] = a[13] & g[14241];
assign g[30624] = b[13] & g[14241];
assign g[22434] = a[13] & g[14242];
assign g[30625] = b[13] & g[14242];
assign g[22435] = a[13] & g[14243];
assign g[30626] = b[13] & g[14243];
assign g[22436] = a[13] & g[14244];
assign g[30627] = b[13] & g[14244];
assign g[22437] = a[13] & g[14245];
assign g[30628] = b[13] & g[14245];
assign g[22438] = a[13] & g[14246];
assign g[30629] = b[13] & g[14246];
assign g[22439] = a[13] & g[14247];
assign g[30630] = b[13] & g[14247];
assign g[22440] = a[13] & g[14248];
assign g[30631] = b[13] & g[14248];
assign g[22441] = a[13] & g[14249];
assign g[30632] = b[13] & g[14249];
assign g[22442] = a[13] & g[14250];
assign g[30633] = b[13] & g[14250];
assign g[22443] = a[13] & g[14251];
assign g[30634] = b[13] & g[14251];
assign g[22444] = a[13] & g[14252];
assign g[30635] = b[13] & g[14252];
assign g[22445] = a[13] & g[14253];
assign g[30636] = b[13] & g[14253];
assign g[22446] = a[13] & g[14254];
assign g[30637] = b[13] & g[14254];
assign g[22447] = a[13] & g[14255];
assign g[30638] = b[13] & g[14255];
assign g[22448] = a[13] & g[14256];
assign g[30639] = b[13] & g[14256];
assign g[22449] = a[13] & g[14257];
assign g[30640] = b[13] & g[14257];
assign g[22450] = a[13] & g[14258];
assign g[30641] = b[13] & g[14258];
assign g[22451] = a[13] & g[14259];
assign g[30642] = b[13] & g[14259];
assign g[22452] = a[13] & g[14260];
assign g[30643] = b[13] & g[14260];
assign g[22453] = a[13] & g[14261];
assign g[30644] = b[13] & g[14261];
assign g[22454] = a[13] & g[14262];
assign g[30645] = b[13] & g[14262];
assign g[22455] = a[13] & g[14263];
assign g[30646] = b[13] & g[14263];
assign g[22456] = a[13] & g[14264];
assign g[30647] = b[13] & g[14264];
assign g[22457] = a[13] & g[14265];
assign g[30648] = b[13] & g[14265];
assign g[22458] = a[13] & g[14266];
assign g[30649] = b[13] & g[14266];
assign g[22459] = a[13] & g[14267];
assign g[30650] = b[13] & g[14267];
assign g[22460] = a[13] & g[14268];
assign g[30651] = b[13] & g[14268];
assign g[22461] = a[13] & g[14269];
assign g[30652] = b[13] & g[14269];
assign g[22462] = a[13] & g[14270];
assign g[30653] = b[13] & g[14270];
assign g[22463] = a[13] & g[14271];
assign g[30654] = b[13] & g[14271];
assign g[22464] = a[13] & g[14272];
assign g[30655] = b[13] & g[14272];
assign g[22465] = a[13] & g[14273];
assign g[30656] = b[13] & g[14273];
assign g[22466] = a[13] & g[14274];
assign g[30657] = b[13] & g[14274];
assign g[22467] = a[13] & g[14275];
assign g[30658] = b[13] & g[14275];
assign g[22468] = a[13] & g[14276];
assign g[30659] = b[13] & g[14276];
assign g[22469] = a[13] & g[14277];
assign g[30660] = b[13] & g[14277];
assign g[22470] = a[13] & g[14278];
assign g[30661] = b[13] & g[14278];
assign g[22471] = a[13] & g[14279];
assign g[30662] = b[13] & g[14279];
assign g[22472] = a[13] & g[14280];
assign g[30663] = b[13] & g[14280];
assign g[22473] = a[13] & g[14281];
assign g[30664] = b[13] & g[14281];
assign g[22474] = a[13] & g[14282];
assign g[30665] = b[13] & g[14282];
assign g[22475] = a[13] & g[14283];
assign g[30666] = b[13] & g[14283];
assign g[22476] = a[13] & g[14284];
assign g[30667] = b[13] & g[14284];
assign g[22477] = a[13] & g[14285];
assign g[30668] = b[13] & g[14285];
assign g[22478] = a[13] & g[14286];
assign g[30669] = b[13] & g[14286];
assign g[22479] = a[13] & g[14287];
assign g[30670] = b[13] & g[14287];
assign g[22480] = a[13] & g[14288];
assign g[30671] = b[13] & g[14288];
assign g[22481] = a[13] & g[14289];
assign g[30672] = b[13] & g[14289];
assign g[22482] = a[13] & g[14290];
assign g[30673] = b[13] & g[14290];
assign g[22483] = a[13] & g[14291];
assign g[30674] = b[13] & g[14291];
assign g[22484] = a[13] & g[14292];
assign g[30675] = b[13] & g[14292];
assign g[22485] = a[13] & g[14293];
assign g[30676] = b[13] & g[14293];
assign g[22486] = a[13] & g[14294];
assign g[30677] = b[13] & g[14294];
assign g[22487] = a[13] & g[14295];
assign g[30678] = b[13] & g[14295];
assign g[22488] = a[13] & g[14296];
assign g[30679] = b[13] & g[14296];
assign g[22489] = a[13] & g[14297];
assign g[30680] = b[13] & g[14297];
assign g[22490] = a[13] & g[14298];
assign g[30681] = b[13] & g[14298];
assign g[22491] = a[13] & g[14299];
assign g[30682] = b[13] & g[14299];
assign g[22492] = a[13] & g[14300];
assign g[30683] = b[13] & g[14300];
assign g[22493] = a[13] & g[14301];
assign g[30684] = b[13] & g[14301];
assign g[22494] = a[13] & g[14302];
assign g[30685] = b[13] & g[14302];
assign g[22495] = a[13] & g[14303];
assign g[30686] = b[13] & g[14303];
assign g[22496] = a[13] & g[14304];
assign g[30687] = b[13] & g[14304];
assign g[22497] = a[13] & g[14305];
assign g[30688] = b[13] & g[14305];
assign g[22498] = a[13] & g[14306];
assign g[30689] = b[13] & g[14306];
assign g[22499] = a[13] & g[14307];
assign g[30690] = b[13] & g[14307];
assign g[22500] = a[13] & g[14308];
assign g[30691] = b[13] & g[14308];
assign g[22501] = a[13] & g[14309];
assign g[30692] = b[13] & g[14309];
assign g[22502] = a[13] & g[14310];
assign g[30693] = b[13] & g[14310];
assign g[22503] = a[13] & g[14311];
assign g[30694] = b[13] & g[14311];
assign g[22504] = a[13] & g[14312];
assign g[30695] = b[13] & g[14312];
assign g[22505] = a[13] & g[14313];
assign g[30696] = b[13] & g[14313];
assign g[22506] = a[13] & g[14314];
assign g[30697] = b[13] & g[14314];
assign g[22507] = a[13] & g[14315];
assign g[30698] = b[13] & g[14315];
assign g[22508] = a[13] & g[14316];
assign g[30699] = b[13] & g[14316];
assign g[22509] = a[13] & g[14317];
assign g[30700] = b[13] & g[14317];
assign g[22510] = a[13] & g[14318];
assign g[30701] = b[13] & g[14318];
assign g[22511] = a[13] & g[14319];
assign g[30702] = b[13] & g[14319];
assign g[22512] = a[13] & g[14320];
assign g[30703] = b[13] & g[14320];
assign g[22513] = a[13] & g[14321];
assign g[30704] = b[13] & g[14321];
assign g[22514] = a[13] & g[14322];
assign g[30705] = b[13] & g[14322];
assign g[22515] = a[13] & g[14323];
assign g[30706] = b[13] & g[14323];
assign g[22516] = a[13] & g[14324];
assign g[30707] = b[13] & g[14324];
assign g[22517] = a[13] & g[14325];
assign g[30708] = b[13] & g[14325];
assign g[22518] = a[13] & g[14326];
assign g[30709] = b[13] & g[14326];
assign g[22519] = a[13] & g[14327];
assign g[30710] = b[13] & g[14327];
assign g[22520] = a[13] & g[14328];
assign g[30711] = b[13] & g[14328];
assign g[22521] = a[13] & g[14329];
assign g[30712] = b[13] & g[14329];
assign g[22522] = a[13] & g[14330];
assign g[30713] = b[13] & g[14330];
assign g[22523] = a[13] & g[14331];
assign g[30714] = b[13] & g[14331];
assign g[22524] = a[13] & g[14332];
assign g[30715] = b[13] & g[14332];
assign g[22525] = a[13] & g[14333];
assign g[30716] = b[13] & g[14333];
assign g[22526] = a[13] & g[14334];
assign g[30717] = b[13] & g[14334];
assign g[22527] = a[13] & g[14335];
assign g[30718] = b[13] & g[14335];
assign g[22528] = a[13] & g[14336];
assign g[30719] = b[13] & g[14336];
assign g[22529] = a[13] & g[14337];
assign g[30720] = b[13] & g[14337];
assign g[22530] = a[13] & g[14338];
assign g[30721] = b[13] & g[14338];
assign g[22531] = a[13] & g[14339];
assign g[30722] = b[13] & g[14339];
assign g[22532] = a[13] & g[14340];
assign g[30723] = b[13] & g[14340];
assign g[22533] = a[13] & g[14341];
assign g[30724] = b[13] & g[14341];
assign g[22534] = a[13] & g[14342];
assign g[30725] = b[13] & g[14342];
assign g[22535] = a[13] & g[14343];
assign g[30726] = b[13] & g[14343];
assign g[22536] = a[13] & g[14344];
assign g[30727] = b[13] & g[14344];
assign g[22537] = a[13] & g[14345];
assign g[30728] = b[13] & g[14345];
assign g[22538] = a[13] & g[14346];
assign g[30729] = b[13] & g[14346];
assign g[22539] = a[13] & g[14347];
assign g[30730] = b[13] & g[14347];
assign g[22540] = a[13] & g[14348];
assign g[30731] = b[13] & g[14348];
assign g[22541] = a[13] & g[14349];
assign g[30732] = b[13] & g[14349];
assign g[22542] = a[13] & g[14350];
assign g[30733] = b[13] & g[14350];
assign g[22543] = a[13] & g[14351];
assign g[30734] = b[13] & g[14351];
assign g[22544] = a[13] & g[14352];
assign g[30735] = b[13] & g[14352];
assign g[22545] = a[13] & g[14353];
assign g[30736] = b[13] & g[14353];
assign g[22546] = a[13] & g[14354];
assign g[30737] = b[13] & g[14354];
assign g[22547] = a[13] & g[14355];
assign g[30738] = b[13] & g[14355];
assign g[22548] = a[13] & g[14356];
assign g[30739] = b[13] & g[14356];
assign g[22549] = a[13] & g[14357];
assign g[30740] = b[13] & g[14357];
assign g[22550] = a[13] & g[14358];
assign g[30741] = b[13] & g[14358];
assign g[22551] = a[13] & g[14359];
assign g[30742] = b[13] & g[14359];
assign g[22552] = a[13] & g[14360];
assign g[30743] = b[13] & g[14360];
assign g[22553] = a[13] & g[14361];
assign g[30744] = b[13] & g[14361];
assign g[22554] = a[13] & g[14362];
assign g[30745] = b[13] & g[14362];
assign g[22555] = a[13] & g[14363];
assign g[30746] = b[13] & g[14363];
assign g[22556] = a[13] & g[14364];
assign g[30747] = b[13] & g[14364];
assign g[22557] = a[13] & g[14365];
assign g[30748] = b[13] & g[14365];
assign g[22558] = a[13] & g[14366];
assign g[30749] = b[13] & g[14366];
assign g[22559] = a[13] & g[14367];
assign g[30750] = b[13] & g[14367];
assign g[22560] = a[13] & g[14368];
assign g[30751] = b[13] & g[14368];
assign g[22561] = a[13] & g[14369];
assign g[30752] = b[13] & g[14369];
assign g[22562] = a[13] & g[14370];
assign g[30753] = b[13] & g[14370];
assign g[22563] = a[13] & g[14371];
assign g[30754] = b[13] & g[14371];
assign g[22564] = a[13] & g[14372];
assign g[30755] = b[13] & g[14372];
assign g[22565] = a[13] & g[14373];
assign g[30756] = b[13] & g[14373];
assign g[22566] = a[13] & g[14374];
assign g[30757] = b[13] & g[14374];
assign g[22567] = a[13] & g[14375];
assign g[30758] = b[13] & g[14375];
assign g[22568] = a[13] & g[14376];
assign g[30759] = b[13] & g[14376];
assign g[22569] = a[13] & g[14377];
assign g[30760] = b[13] & g[14377];
assign g[22570] = a[13] & g[14378];
assign g[30761] = b[13] & g[14378];
assign g[22571] = a[13] & g[14379];
assign g[30762] = b[13] & g[14379];
assign g[22572] = a[13] & g[14380];
assign g[30763] = b[13] & g[14380];
assign g[22573] = a[13] & g[14381];
assign g[30764] = b[13] & g[14381];
assign g[22574] = a[13] & g[14382];
assign g[30765] = b[13] & g[14382];
assign g[22575] = a[13] & g[14383];
assign g[30766] = b[13] & g[14383];
assign g[22576] = a[13] & g[14384];
assign g[30767] = b[13] & g[14384];
assign g[22577] = a[13] & g[14385];
assign g[30768] = b[13] & g[14385];
assign g[22578] = a[13] & g[14386];
assign g[30769] = b[13] & g[14386];
assign g[22579] = a[13] & g[14387];
assign g[30770] = b[13] & g[14387];
assign g[22580] = a[13] & g[14388];
assign g[30771] = b[13] & g[14388];
assign g[22581] = a[13] & g[14389];
assign g[30772] = b[13] & g[14389];
assign g[22582] = a[13] & g[14390];
assign g[30773] = b[13] & g[14390];
assign g[22583] = a[13] & g[14391];
assign g[30774] = b[13] & g[14391];
assign g[22584] = a[13] & g[14392];
assign g[30775] = b[13] & g[14392];
assign g[22585] = a[13] & g[14393];
assign g[30776] = b[13] & g[14393];
assign g[22586] = a[13] & g[14394];
assign g[30777] = b[13] & g[14394];
assign g[22587] = a[13] & g[14395];
assign g[30778] = b[13] & g[14395];
assign g[22588] = a[13] & g[14396];
assign g[30779] = b[13] & g[14396];
assign g[22589] = a[13] & g[14397];
assign g[30780] = b[13] & g[14397];
assign g[22590] = a[13] & g[14398];
assign g[30781] = b[13] & g[14398];
assign g[22591] = a[13] & g[14399];
assign g[30782] = b[13] & g[14399];
assign g[22592] = a[13] & g[14400];
assign g[30783] = b[13] & g[14400];
assign g[22593] = a[13] & g[14401];
assign g[30784] = b[13] & g[14401];
assign g[22594] = a[13] & g[14402];
assign g[30785] = b[13] & g[14402];
assign g[22595] = a[13] & g[14403];
assign g[30786] = b[13] & g[14403];
assign g[22596] = a[13] & g[14404];
assign g[30787] = b[13] & g[14404];
assign g[22597] = a[13] & g[14405];
assign g[30788] = b[13] & g[14405];
assign g[22598] = a[13] & g[14406];
assign g[30789] = b[13] & g[14406];
assign g[22599] = a[13] & g[14407];
assign g[30790] = b[13] & g[14407];
assign g[22600] = a[13] & g[14408];
assign g[30791] = b[13] & g[14408];
assign g[22601] = a[13] & g[14409];
assign g[30792] = b[13] & g[14409];
assign g[22602] = a[13] & g[14410];
assign g[30793] = b[13] & g[14410];
assign g[22603] = a[13] & g[14411];
assign g[30794] = b[13] & g[14411];
assign g[22604] = a[13] & g[14412];
assign g[30795] = b[13] & g[14412];
assign g[22605] = a[13] & g[14413];
assign g[30796] = b[13] & g[14413];
assign g[22606] = a[13] & g[14414];
assign g[30797] = b[13] & g[14414];
assign g[22607] = a[13] & g[14415];
assign g[30798] = b[13] & g[14415];
assign g[22608] = a[13] & g[14416];
assign g[30799] = b[13] & g[14416];
assign g[22609] = a[13] & g[14417];
assign g[30800] = b[13] & g[14417];
assign g[22610] = a[13] & g[14418];
assign g[30801] = b[13] & g[14418];
assign g[22611] = a[13] & g[14419];
assign g[30802] = b[13] & g[14419];
assign g[22612] = a[13] & g[14420];
assign g[30803] = b[13] & g[14420];
assign g[22613] = a[13] & g[14421];
assign g[30804] = b[13] & g[14421];
assign g[22614] = a[13] & g[14422];
assign g[30805] = b[13] & g[14422];
assign g[22615] = a[13] & g[14423];
assign g[30806] = b[13] & g[14423];
assign g[22616] = a[13] & g[14424];
assign g[30807] = b[13] & g[14424];
assign g[22617] = a[13] & g[14425];
assign g[30808] = b[13] & g[14425];
assign g[22618] = a[13] & g[14426];
assign g[30809] = b[13] & g[14426];
assign g[22619] = a[13] & g[14427];
assign g[30810] = b[13] & g[14427];
assign g[22620] = a[13] & g[14428];
assign g[30811] = b[13] & g[14428];
assign g[22621] = a[13] & g[14429];
assign g[30812] = b[13] & g[14429];
assign g[22622] = a[13] & g[14430];
assign g[30813] = b[13] & g[14430];
assign g[22623] = a[13] & g[14431];
assign g[30814] = b[13] & g[14431];
assign g[22624] = a[13] & g[14432];
assign g[30815] = b[13] & g[14432];
assign g[22625] = a[13] & g[14433];
assign g[30816] = b[13] & g[14433];
assign g[22626] = a[13] & g[14434];
assign g[30817] = b[13] & g[14434];
assign g[22627] = a[13] & g[14435];
assign g[30818] = b[13] & g[14435];
assign g[22628] = a[13] & g[14436];
assign g[30819] = b[13] & g[14436];
assign g[22629] = a[13] & g[14437];
assign g[30820] = b[13] & g[14437];
assign g[22630] = a[13] & g[14438];
assign g[30821] = b[13] & g[14438];
assign g[22631] = a[13] & g[14439];
assign g[30822] = b[13] & g[14439];
assign g[22632] = a[13] & g[14440];
assign g[30823] = b[13] & g[14440];
assign g[22633] = a[13] & g[14441];
assign g[30824] = b[13] & g[14441];
assign g[22634] = a[13] & g[14442];
assign g[30825] = b[13] & g[14442];
assign g[22635] = a[13] & g[14443];
assign g[30826] = b[13] & g[14443];
assign g[22636] = a[13] & g[14444];
assign g[30827] = b[13] & g[14444];
assign g[22637] = a[13] & g[14445];
assign g[30828] = b[13] & g[14445];
assign g[22638] = a[13] & g[14446];
assign g[30829] = b[13] & g[14446];
assign g[22639] = a[13] & g[14447];
assign g[30830] = b[13] & g[14447];
assign g[22640] = a[13] & g[14448];
assign g[30831] = b[13] & g[14448];
assign g[22641] = a[13] & g[14449];
assign g[30832] = b[13] & g[14449];
assign g[22642] = a[13] & g[14450];
assign g[30833] = b[13] & g[14450];
assign g[22643] = a[13] & g[14451];
assign g[30834] = b[13] & g[14451];
assign g[22644] = a[13] & g[14452];
assign g[30835] = b[13] & g[14452];
assign g[22645] = a[13] & g[14453];
assign g[30836] = b[13] & g[14453];
assign g[22646] = a[13] & g[14454];
assign g[30837] = b[13] & g[14454];
assign g[22647] = a[13] & g[14455];
assign g[30838] = b[13] & g[14455];
assign g[22648] = a[13] & g[14456];
assign g[30839] = b[13] & g[14456];
assign g[22649] = a[13] & g[14457];
assign g[30840] = b[13] & g[14457];
assign g[22650] = a[13] & g[14458];
assign g[30841] = b[13] & g[14458];
assign g[22651] = a[13] & g[14459];
assign g[30842] = b[13] & g[14459];
assign g[22652] = a[13] & g[14460];
assign g[30843] = b[13] & g[14460];
assign g[22653] = a[13] & g[14461];
assign g[30844] = b[13] & g[14461];
assign g[22654] = a[13] & g[14462];
assign g[30845] = b[13] & g[14462];
assign g[22655] = a[13] & g[14463];
assign g[30846] = b[13] & g[14463];
assign g[22656] = a[13] & g[14464];
assign g[30847] = b[13] & g[14464];
assign g[22657] = a[13] & g[14465];
assign g[30848] = b[13] & g[14465];
assign g[22658] = a[13] & g[14466];
assign g[30849] = b[13] & g[14466];
assign g[22659] = a[13] & g[14467];
assign g[30850] = b[13] & g[14467];
assign g[22660] = a[13] & g[14468];
assign g[30851] = b[13] & g[14468];
assign g[22661] = a[13] & g[14469];
assign g[30852] = b[13] & g[14469];
assign g[22662] = a[13] & g[14470];
assign g[30853] = b[13] & g[14470];
assign g[22663] = a[13] & g[14471];
assign g[30854] = b[13] & g[14471];
assign g[22664] = a[13] & g[14472];
assign g[30855] = b[13] & g[14472];
assign g[22665] = a[13] & g[14473];
assign g[30856] = b[13] & g[14473];
assign g[22666] = a[13] & g[14474];
assign g[30857] = b[13] & g[14474];
assign g[22667] = a[13] & g[14475];
assign g[30858] = b[13] & g[14475];
assign g[22668] = a[13] & g[14476];
assign g[30859] = b[13] & g[14476];
assign g[22669] = a[13] & g[14477];
assign g[30860] = b[13] & g[14477];
assign g[22670] = a[13] & g[14478];
assign g[30861] = b[13] & g[14478];
assign g[22671] = a[13] & g[14479];
assign g[30862] = b[13] & g[14479];
assign g[22672] = a[13] & g[14480];
assign g[30863] = b[13] & g[14480];
assign g[22673] = a[13] & g[14481];
assign g[30864] = b[13] & g[14481];
assign g[22674] = a[13] & g[14482];
assign g[30865] = b[13] & g[14482];
assign g[22675] = a[13] & g[14483];
assign g[30866] = b[13] & g[14483];
assign g[22676] = a[13] & g[14484];
assign g[30867] = b[13] & g[14484];
assign g[22677] = a[13] & g[14485];
assign g[30868] = b[13] & g[14485];
assign g[22678] = a[13] & g[14486];
assign g[30869] = b[13] & g[14486];
assign g[22679] = a[13] & g[14487];
assign g[30870] = b[13] & g[14487];
assign g[22680] = a[13] & g[14488];
assign g[30871] = b[13] & g[14488];
assign g[22681] = a[13] & g[14489];
assign g[30872] = b[13] & g[14489];
assign g[22682] = a[13] & g[14490];
assign g[30873] = b[13] & g[14490];
assign g[22683] = a[13] & g[14491];
assign g[30874] = b[13] & g[14491];
assign g[22684] = a[13] & g[14492];
assign g[30875] = b[13] & g[14492];
assign g[22685] = a[13] & g[14493];
assign g[30876] = b[13] & g[14493];
assign g[22686] = a[13] & g[14494];
assign g[30877] = b[13] & g[14494];
assign g[22687] = a[13] & g[14495];
assign g[30878] = b[13] & g[14495];
assign g[22688] = a[13] & g[14496];
assign g[30879] = b[13] & g[14496];
assign g[22689] = a[13] & g[14497];
assign g[30880] = b[13] & g[14497];
assign g[22690] = a[13] & g[14498];
assign g[30881] = b[13] & g[14498];
assign g[22691] = a[13] & g[14499];
assign g[30882] = b[13] & g[14499];
assign g[22692] = a[13] & g[14500];
assign g[30883] = b[13] & g[14500];
assign g[22693] = a[13] & g[14501];
assign g[30884] = b[13] & g[14501];
assign g[22694] = a[13] & g[14502];
assign g[30885] = b[13] & g[14502];
assign g[22695] = a[13] & g[14503];
assign g[30886] = b[13] & g[14503];
assign g[22696] = a[13] & g[14504];
assign g[30887] = b[13] & g[14504];
assign g[22697] = a[13] & g[14505];
assign g[30888] = b[13] & g[14505];
assign g[22698] = a[13] & g[14506];
assign g[30889] = b[13] & g[14506];
assign g[22699] = a[13] & g[14507];
assign g[30890] = b[13] & g[14507];
assign g[22700] = a[13] & g[14508];
assign g[30891] = b[13] & g[14508];
assign g[22701] = a[13] & g[14509];
assign g[30892] = b[13] & g[14509];
assign g[22702] = a[13] & g[14510];
assign g[30893] = b[13] & g[14510];
assign g[22703] = a[13] & g[14511];
assign g[30894] = b[13] & g[14511];
assign g[22704] = a[13] & g[14512];
assign g[30895] = b[13] & g[14512];
assign g[22705] = a[13] & g[14513];
assign g[30896] = b[13] & g[14513];
assign g[22706] = a[13] & g[14514];
assign g[30897] = b[13] & g[14514];
assign g[22707] = a[13] & g[14515];
assign g[30898] = b[13] & g[14515];
assign g[22708] = a[13] & g[14516];
assign g[30899] = b[13] & g[14516];
assign g[22709] = a[13] & g[14517];
assign g[30900] = b[13] & g[14517];
assign g[22710] = a[13] & g[14518];
assign g[30901] = b[13] & g[14518];
assign g[22711] = a[13] & g[14519];
assign g[30902] = b[13] & g[14519];
assign g[22712] = a[13] & g[14520];
assign g[30903] = b[13] & g[14520];
assign g[22713] = a[13] & g[14521];
assign g[30904] = b[13] & g[14521];
assign g[22714] = a[13] & g[14522];
assign g[30905] = b[13] & g[14522];
assign g[22715] = a[13] & g[14523];
assign g[30906] = b[13] & g[14523];
assign g[22716] = a[13] & g[14524];
assign g[30907] = b[13] & g[14524];
assign g[22717] = a[13] & g[14525];
assign g[30908] = b[13] & g[14525];
assign g[22718] = a[13] & g[14526];
assign g[30909] = b[13] & g[14526];
assign g[22719] = a[13] & g[14527];
assign g[30910] = b[13] & g[14527];
assign g[22720] = a[13] & g[14528];
assign g[30911] = b[13] & g[14528];
assign g[22721] = a[13] & g[14529];
assign g[30912] = b[13] & g[14529];
assign g[22722] = a[13] & g[14530];
assign g[30913] = b[13] & g[14530];
assign g[22723] = a[13] & g[14531];
assign g[30914] = b[13] & g[14531];
assign g[22724] = a[13] & g[14532];
assign g[30915] = b[13] & g[14532];
assign g[22725] = a[13] & g[14533];
assign g[30916] = b[13] & g[14533];
assign g[22726] = a[13] & g[14534];
assign g[30917] = b[13] & g[14534];
assign g[22727] = a[13] & g[14535];
assign g[30918] = b[13] & g[14535];
assign g[22728] = a[13] & g[14536];
assign g[30919] = b[13] & g[14536];
assign g[22729] = a[13] & g[14537];
assign g[30920] = b[13] & g[14537];
assign g[22730] = a[13] & g[14538];
assign g[30921] = b[13] & g[14538];
assign g[22731] = a[13] & g[14539];
assign g[30922] = b[13] & g[14539];
assign g[22732] = a[13] & g[14540];
assign g[30923] = b[13] & g[14540];
assign g[22733] = a[13] & g[14541];
assign g[30924] = b[13] & g[14541];
assign g[22734] = a[13] & g[14542];
assign g[30925] = b[13] & g[14542];
assign g[22735] = a[13] & g[14543];
assign g[30926] = b[13] & g[14543];
assign g[22736] = a[13] & g[14544];
assign g[30927] = b[13] & g[14544];
assign g[22737] = a[13] & g[14545];
assign g[30928] = b[13] & g[14545];
assign g[22738] = a[13] & g[14546];
assign g[30929] = b[13] & g[14546];
assign g[22739] = a[13] & g[14547];
assign g[30930] = b[13] & g[14547];
assign g[22740] = a[13] & g[14548];
assign g[30931] = b[13] & g[14548];
assign g[22741] = a[13] & g[14549];
assign g[30932] = b[13] & g[14549];
assign g[22742] = a[13] & g[14550];
assign g[30933] = b[13] & g[14550];
assign g[22743] = a[13] & g[14551];
assign g[30934] = b[13] & g[14551];
assign g[22744] = a[13] & g[14552];
assign g[30935] = b[13] & g[14552];
assign g[22745] = a[13] & g[14553];
assign g[30936] = b[13] & g[14553];
assign g[22746] = a[13] & g[14554];
assign g[30937] = b[13] & g[14554];
assign g[22747] = a[13] & g[14555];
assign g[30938] = b[13] & g[14555];
assign g[22748] = a[13] & g[14556];
assign g[30939] = b[13] & g[14556];
assign g[22749] = a[13] & g[14557];
assign g[30940] = b[13] & g[14557];
assign g[22750] = a[13] & g[14558];
assign g[30941] = b[13] & g[14558];
assign g[22751] = a[13] & g[14559];
assign g[30942] = b[13] & g[14559];
assign g[22752] = a[13] & g[14560];
assign g[30943] = b[13] & g[14560];
assign g[22753] = a[13] & g[14561];
assign g[30944] = b[13] & g[14561];
assign g[22754] = a[13] & g[14562];
assign g[30945] = b[13] & g[14562];
assign g[22755] = a[13] & g[14563];
assign g[30946] = b[13] & g[14563];
assign g[22756] = a[13] & g[14564];
assign g[30947] = b[13] & g[14564];
assign g[22757] = a[13] & g[14565];
assign g[30948] = b[13] & g[14565];
assign g[22758] = a[13] & g[14566];
assign g[30949] = b[13] & g[14566];
assign g[22759] = a[13] & g[14567];
assign g[30950] = b[13] & g[14567];
assign g[22760] = a[13] & g[14568];
assign g[30951] = b[13] & g[14568];
assign g[22761] = a[13] & g[14569];
assign g[30952] = b[13] & g[14569];
assign g[22762] = a[13] & g[14570];
assign g[30953] = b[13] & g[14570];
assign g[22763] = a[13] & g[14571];
assign g[30954] = b[13] & g[14571];
assign g[22764] = a[13] & g[14572];
assign g[30955] = b[13] & g[14572];
assign g[22765] = a[13] & g[14573];
assign g[30956] = b[13] & g[14573];
assign g[22766] = a[13] & g[14574];
assign g[30957] = b[13] & g[14574];
assign g[22767] = a[13] & g[14575];
assign g[30958] = b[13] & g[14575];
assign g[22768] = a[13] & g[14576];
assign g[30959] = b[13] & g[14576];
assign g[22769] = a[13] & g[14577];
assign g[30960] = b[13] & g[14577];
assign g[22770] = a[13] & g[14578];
assign g[30961] = b[13] & g[14578];
assign g[22771] = a[13] & g[14579];
assign g[30962] = b[13] & g[14579];
assign g[22772] = a[13] & g[14580];
assign g[30963] = b[13] & g[14580];
assign g[22773] = a[13] & g[14581];
assign g[30964] = b[13] & g[14581];
assign g[22774] = a[13] & g[14582];
assign g[30965] = b[13] & g[14582];
assign g[22775] = a[13] & g[14583];
assign g[30966] = b[13] & g[14583];
assign g[22776] = a[13] & g[14584];
assign g[30967] = b[13] & g[14584];
assign g[22777] = a[13] & g[14585];
assign g[30968] = b[13] & g[14585];
assign g[22778] = a[13] & g[14586];
assign g[30969] = b[13] & g[14586];
assign g[22779] = a[13] & g[14587];
assign g[30970] = b[13] & g[14587];
assign g[22780] = a[13] & g[14588];
assign g[30971] = b[13] & g[14588];
assign g[22781] = a[13] & g[14589];
assign g[30972] = b[13] & g[14589];
assign g[22782] = a[13] & g[14590];
assign g[30973] = b[13] & g[14590];
assign g[22783] = a[13] & g[14591];
assign g[30974] = b[13] & g[14591];
assign g[22784] = a[13] & g[14592];
assign g[30975] = b[13] & g[14592];
assign g[22785] = a[13] & g[14593];
assign g[30976] = b[13] & g[14593];
assign g[22786] = a[13] & g[14594];
assign g[30977] = b[13] & g[14594];
assign g[22787] = a[13] & g[14595];
assign g[30978] = b[13] & g[14595];
assign g[22788] = a[13] & g[14596];
assign g[30979] = b[13] & g[14596];
assign g[22789] = a[13] & g[14597];
assign g[30980] = b[13] & g[14597];
assign g[22790] = a[13] & g[14598];
assign g[30981] = b[13] & g[14598];
assign g[22791] = a[13] & g[14599];
assign g[30982] = b[13] & g[14599];
assign g[22792] = a[13] & g[14600];
assign g[30983] = b[13] & g[14600];
assign g[22793] = a[13] & g[14601];
assign g[30984] = b[13] & g[14601];
assign g[22794] = a[13] & g[14602];
assign g[30985] = b[13] & g[14602];
assign g[22795] = a[13] & g[14603];
assign g[30986] = b[13] & g[14603];
assign g[22796] = a[13] & g[14604];
assign g[30987] = b[13] & g[14604];
assign g[22797] = a[13] & g[14605];
assign g[30988] = b[13] & g[14605];
assign g[22798] = a[13] & g[14606];
assign g[30989] = b[13] & g[14606];
assign g[22799] = a[13] & g[14607];
assign g[30990] = b[13] & g[14607];
assign g[22800] = a[13] & g[14608];
assign g[30991] = b[13] & g[14608];
assign g[22801] = a[13] & g[14609];
assign g[30992] = b[13] & g[14609];
assign g[22802] = a[13] & g[14610];
assign g[30993] = b[13] & g[14610];
assign g[22803] = a[13] & g[14611];
assign g[30994] = b[13] & g[14611];
assign g[22804] = a[13] & g[14612];
assign g[30995] = b[13] & g[14612];
assign g[22805] = a[13] & g[14613];
assign g[30996] = b[13] & g[14613];
assign g[22806] = a[13] & g[14614];
assign g[30997] = b[13] & g[14614];
assign g[22807] = a[13] & g[14615];
assign g[30998] = b[13] & g[14615];
assign g[22808] = a[13] & g[14616];
assign g[30999] = b[13] & g[14616];
assign g[22809] = a[13] & g[14617];
assign g[31000] = b[13] & g[14617];
assign g[22810] = a[13] & g[14618];
assign g[31001] = b[13] & g[14618];
assign g[22811] = a[13] & g[14619];
assign g[31002] = b[13] & g[14619];
assign g[22812] = a[13] & g[14620];
assign g[31003] = b[13] & g[14620];
assign g[22813] = a[13] & g[14621];
assign g[31004] = b[13] & g[14621];
assign g[22814] = a[13] & g[14622];
assign g[31005] = b[13] & g[14622];
assign g[22815] = a[13] & g[14623];
assign g[31006] = b[13] & g[14623];
assign g[22816] = a[13] & g[14624];
assign g[31007] = b[13] & g[14624];
assign g[22817] = a[13] & g[14625];
assign g[31008] = b[13] & g[14625];
assign g[22818] = a[13] & g[14626];
assign g[31009] = b[13] & g[14626];
assign g[22819] = a[13] & g[14627];
assign g[31010] = b[13] & g[14627];
assign g[22820] = a[13] & g[14628];
assign g[31011] = b[13] & g[14628];
assign g[22821] = a[13] & g[14629];
assign g[31012] = b[13] & g[14629];
assign g[22822] = a[13] & g[14630];
assign g[31013] = b[13] & g[14630];
assign g[22823] = a[13] & g[14631];
assign g[31014] = b[13] & g[14631];
assign g[22824] = a[13] & g[14632];
assign g[31015] = b[13] & g[14632];
assign g[22825] = a[13] & g[14633];
assign g[31016] = b[13] & g[14633];
assign g[22826] = a[13] & g[14634];
assign g[31017] = b[13] & g[14634];
assign g[22827] = a[13] & g[14635];
assign g[31018] = b[13] & g[14635];
assign g[22828] = a[13] & g[14636];
assign g[31019] = b[13] & g[14636];
assign g[22829] = a[13] & g[14637];
assign g[31020] = b[13] & g[14637];
assign g[22830] = a[13] & g[14638];
assign g[31021] = b[13] & g[14638];
assign g[22831] = a[13] & g[14639];
assign g[31022] = b[13] & g[14639];
assign g[22832] = a[13] & g[14640];
assign g[31023] = b[13] & g[14640];
assign g[22833] = a[13] & g[14641];
assign g[31024] = b[13] & g[14641];
assign g[22834] = a[13] & g[14642];
assign g[31025] = b[13] & g[14642];
assign g[22835] = a[13] & g[14643];
assign g[31026] = b[13] & g[14643];
assign g[22836] = a[13] & g[14644];
assign g[31027] = b[13] & g[14644];
assign g[22837] = a[13] & g[14645];
assign g[31028] = b[13] & g[14645];
assign g[22838] = a[13] & g[14646];
assign g[31029] = b[13] & g[14646];
assign g[22839] = a[13] & g[14647];
assign g[31030] = b[13] & g[14647];
assign g[22840] = a[13] & g[14648];
assign g[31031] = b[13] & g[14648];
assign g[22841] = a[13] & g[14649];
assign g[31032] = b[13] & g[14649];
assign g[22842] = a[13] & g[14650];
assign g[31033] = b[13] & g[14650];
assign g[22843] = a[13] & g[14651];
assign g[31034] = b[13] & g[14651];
assign g[22844] = a[13] & g[14652];
assign g[31035] = b[13] & g[14652];
assign g[22845] = a[13] & g[14653];
assign g[31036] = b[13] & g[14653];
assign g[22846] = a[13] & g[14654];
assign g[31037] = b[13] & g[14654];
assign g[22847] = a[13] & g[14655];
assign g[31038] = b[13] & g[14655];
assign g[22848] = a[13] & g[14656];
assign g[31039] = b[13] & g[14656];
assign g[22849] = a[13] & g[14657];
assign g[31040] = b[13] & g[14657];
assign g[22850] = a[13] & g[14658];
assign g[31041] = b[13] & g[14658];
assign g[22851] = a[13] & g[14659];
assign g[31042] = b[13] & g[14659];
assign g[22852] = a[13] & g[14660];
assign g[31043] = b[13] & g[14660];
assign g[22853] = a[13] & g[14661];
assign g[31044] = b[13] & g[14661];
assign g[22854] = a[13] & g[14662];
assign g[31045] = b[13] & g[14662];
assign g[22855] = a[13] & g[14663];
assign g[31046] = b[13] & g[14663];
assign g[22856] = a[13] & g[14664];
assign g[31047] = b[13] & g[14664];
assign g[22857] = a[13] & g[14665];
assign g[31048] = b[13] & g[14665];
assign g[22858] = a[13] & g[14666];
assign g[31049] = b[13] & g[14666];
assign g[22859] = a[13] & g[14667];
assign g[31050] = b[13] & g[14667];
assign g[22860] = a[13] & g[14668];
assign g[31051] = b[13] & g[14668];
assign g[22861] = a[13] & g[14669];
assign g[31052] = b[13] & g[14669];
assign g[22862] = a[13] & g[14670];
assign g[31053] = b[13] & g[14670];
assign g[22863] = a[13] & g[14671];
assign g[31054] = b[13] & g[14671];
assign g[22864] = a[13] & g[14672];
assign g[31055] = b[13] & g[14672];
assign g[22865] = a[13] & g[14673];
assign g[31056] = b[13] & g[14673];
assign g[22866] = a[13] & g[14674];
assign g[31057] = b[13] & g[14674];
assign g[22867] = a[13] & g[14675];
assign g[31058] = b[13] & g[14675];
assign g[22868] = a[13] & g[14676];
assign g[31059] = b[13] & g[14676];
assign g[22869] = a[13] & g[14677];
assign g[31060] = b[13] & g[14677];
assign g[22870] = a[13] & g[14678];
assign g[31061] = b[13] & g[14678];
assign g[22871] = a[13] & g[14679];
assign g[31062] = b[13] & g[14679];
assign g[22872] = a[13] & g[14680];
assign g[31063] = b[13] & g[14680];
assign g[22873] = a[13] & g[14681];
assign g[31064] = b[13] & g[14681];
assign g[22874] = a[13] & g[14682];
assign g[31065] = b[13] & g[14682];
assign g[22875] = a[13] & g[14683];
assign g[31066] = b[13] & g[14683];
assign g[22876] = a[13] & g[14684];
assign g[31067] = b[13] & g[14684];
assign g[22877] = a[13] & g[14685];
assign g[31068] = b[13] & g[14685];
assign g[22878] = a[13] & g[14686];
assign g[31069] = b[13] & g[14686];
assign g[22879] = a[13] & g[14687];
assign g[31070] = b[13] & g[14687];
assign g[22880] = a[13] & g[14688];
assign g[31071] = b[13] & g[14688];
assign g[22881] = a[13] & g[14689];
assign g[31072] = b[13] & g[14689];
assign g[22882] = a[13] & g[14690];
assign g[31073] = b[13] & g[14690];
assign g[22883] = a[13] & g[14691];
assign g[31074] = b[13] & g[14691];
assign g[22884] = a[13] & g[14692];
assign g[31075] = b[13] & g[14692];
assign g[22885] = a[13] & g[14693];
assign g[31076] = b[13] & g[14693];
assign g[22886] = a[13] & g[14694];
assign g[31077] = b[13] & g[14694];
assign g[22887] = a[13] & g[14695];
assign g[31078] = b[13] & g[14695];
assign g[22888] = a[13] & g[14696];
assign g[31079] = b[13] & g[14696];
assign g[22889] = a[13] & g[14697];
assign g[31080] = b[13] & g[14697];
assign g[22890] = a[13] & g[14698];
assign g[31081] = b[13] & g[14698];
assign g[22891] = a[13] & g[14699];
assign g[31082] = b[13] & g[14699];
assign g[22892] = a[13] & g[14700];
assign g[31083] = b[13] & g[14700];
assign g[22893] = a[13] & g[14701];
assign g[31084] = b[13] & g[14701];
assign g[22894] = a[13] & g[14702];
assign g[31085] = b[13] & g[14702];
assign g[22895] = a[13] & g[14703];
assign g[31086] = b[13] & g[14703];
assign g[22896] = a[13] & g[14704];
assign g[31087] = b[13] & g[14704];
assign g[22897] = a[13] & g[14705];
assign g[31088] = b[13] & g[14705];
assign g[22898] = a[13] & g[14706];
assign g[31089] = b[13] & g[14706];
assign g[22899] = a[13] & g[14707];
assign g[31090] = b[13] & g[14707];
assign g[22900] = a[13] & g[14708];
assign g[31091] = b[13] & g[14708];
assign g[22901] = a[13] & g[14709];
assign g[31092] = b[13] & g[14709];
assign g[22902] = a[13] & g[14710];
assign g[31093] = b[13] & g[14710];
assign g[22903] = a[13] & g[14711];
assign g[31094] = b[13] & g[14711];
assign g[22904] = a[13] & g[14712];
assign g[31095] = b[13] & g[14712];
assign g[22905] = a[13] & g[14713];
assign g[31096] = b[13] & g[14713];
assign g[22906] = a[13] & g[14714];
assign g[31097] = b[13] & g[14714];
assign g[22907] = a[13] & g[14715];
assign g[31098] = b[13] & g[14715];
assign g[22908] = a[13] & g[14716];
assign g[31099] = b[13] & g[14716];
assign g[22909] = a[13] & g[14717];
assign g[31100] = b[13] & g[14717];
assign g[22910] = a[13] & g[14718];
assign g[31101] = b[13] & g[14718];
assign g[22911] = a[13] & g[14719];
assign g[31102] = b[13] & g[14719];
assign g[22912] = a[13] & g[14720];
assign g[31103] = b[13] & g[14720];
assign g[22913] = a[13] & g[14721];
assign g[31104] = b[13] & g[14721];
assign g[22914] = a[13] & g[14722];
assign g[31105] = b[13] & g[14722];
assign g[22915] = a[13] & g[14723];
assign g[31106] = b[13] & g[14723];
assign g[22916] = a[13] & g[14724];
assign g[31107] = b[13] & g[14724];
assign g[22917] = a[13] & g[14725];
assign g[31108] = b[13] & g[14725];
assign g[22918] = a[13] & g[14726];
assign g[31109] = b[13] & g[14726];
assign g[22919] = a[13] & g[14727];
assign g[31110] = b[13] & g[14727];
assign g[22920] = a[13] & g[14728];
assign g[31111] = b[13] & g[14728];
assign g[22921] = a[13] & g[14729];
assign g[31112] = b[13] & g[14729];
assign g[22922] = a[13] & g[14730];
assign g[31113] = b[13] & g[14730];
assign g[22923] = a[13] & g[14731];
assign g[31114] = b[13] & g[14731];
assign g[22924] = a[13] & g[14732];
assign g[31115] = b[13] & g[14732];
assign g[22925] = a[13] & g[14733];
assign g[31116] = b[13] & g[14733];
assign g[22926] = a[13] & g[14734];
assign g[31117] = b[13] & g[14734];
assign g[22927] = a[13] & g[14735];
assign g[31118] = b[13] & g[14735];
assign g[22928] = a[13] & g[14736];
assign g[31119] = b[13] & g[14736];
assign g[22929] = a[13] & g[14737];
assign g[31120] = b[13] & g[14737];
assign g[22930] = a[13] & g[14738];
assign g[31121] = b[13] & g[14738];
assign g[22931] = a[13] & g[14739];
assign g[31122] = b[13] & g[14739];
assign g[22932] = a[13] & g[14740];
assign g[31123] = b[13] & g[14740];
assign g[22933] = a[13] & g[14741];
assign g[31124] = b[13] & g[14741];
assign g[22934] = a[13] & g[14742];
assign g[31125] = b[13] & g[14742];
assign g[22935] = a[13] & g[14743];
assign g[31126] = b[13] & g[14743];
assign g[22936] = a[13] & g[14744];
assign g[31127] = b[13] & g[14744];
assign g[22937] = a[13] & g[14745];
assign g[31128] = b[13] & g[14745];
assign g[22938] = a[13] & g[14746];
assign g[31129] = b[13] & g[14746];
assign g[22939] = a[13] & g[14747];
assign g[31130] = b[13] & g[14747];
assign g[22940] = a[13] & g[14748];
assign g[31131] = b[13] & g[14748];
assign g[22941] = a[13] & g[14749];
assign g[31132] = b[13] & g[14749];
assign g[22942] = a[13] & g[14750];
assign g[31133] = b[13] & g[14750];
assign g[22943] = a[13] & g[14751];
assign g[31134] = b[13] & g[14751];
assign g[22944] = a[13] & g[14752];
assign g[31135] = b[13] & g[14752];
assign g[22945] = a[13] & g[14753];
assign g[31136] = b[13] & g[14753];
assign g[22946] = a[13] & g[14754];
assign g[31137] = b[13] & g[14754];
assign g[22947] = a[13] & g[14755];
assign g[31138] = b[13] & g[14755];
assign g[22948] = a[13] & g[14756];
assign g[31139] = b[13] & g[14756];
assign g[22949] = a[13] & g[14757];
assign g[31140] = b[13] & g[14757];
assign g[22950] = a[13] & g[14758];
assign g[31141] = b[13] & g[14758];
assign g[22951] = a[13] & g[14759];
assign g[31142] = b[13] & g[14759];
assign g[22952] = a[13] & g[14760];
assign g[31143] = b[13] & g[14760];
assign g[22953] = a[13] & g[14761];
assign g[31144] = b[13] & g[14761];
assign g[22954] = a[13] & g[14762];
assign g[31145] = b[13] & g[14762];
assign g[22955] = a[13] & g[14763];
assign g[31146] = b[13] & g[14763];
assign g[22956] = a[13] & g[14764];
assign g[31147] = b[13] & g[14764];
assign g[22957] = a[13] & g[14765];
assign g[31148] = b[13] & g[14765];
assign g[22958] = a[13] & g[14766];
assign g[31149] = b[13] & g[14766];
assign g[22959] = a[13] & g[14767];
assign g[31150] = b[13] & g[14767];
assign g[22960] = a[13] & g[14768];
assign g[31151] = b[13] & g[14768];
assign g[22961] = a[13] & g[14769];
assign g[31152] = b[13] & g[14769];
assign g[22962] = a[13] & g[14770];
assign g[31153] = b[13] & g[14770];
assign g[22963] = a[13] & g[14771];
assign g[31154] = b[13] & g[14771];
assign g[22964] = a[13] & g[14772];
assign g[31155] = b[13] & g[14772];
assign g[22965] = a[13] & g[14773];
assign g[31156] = b[13] & g[14773];
assign g[22966] = a[13] & g[14774];
assign g[31157] = b[13] & g[14774];
assign g[22967] = a[13] & g[14775];
assign g[31158] = b[13] & g[14775];
assign g[22968] = a[13] & g[14776];
assign g[31159] = b[13] & g[14776];
assign g[22969] = a[13] & g[14777];
assign g[31160] = b[13] & g[14777];
assign g[22970] = a[13] & g[14778];
assign g[31161] = b[13] & g[14778];
assign g[22971] = a[13] & g[14779];
assign g[31162] = b[13] & g[14779];
assign g[22972] = a[13] & g[14780];
assign g[31163] = b[13] & g[14780];
assign g[22973] = a[13] & g[14781];
assign g[31164] = b[13] & g[14781];
assign g[22974] = a[13] & g[14782];
assign g[31165] = b[13] & g[14782];
assign g[22975] = a[13] & g[14783];
assign g[31166] = b[13] & g[14783];
assign g[22976] = a[13] & g[14784];
assign g[31167] = b[13] & g[14784];
assign g[22977] = a[13] & g[14785];
assign g[31168] = b[13] & g[14785];
assign g[22978] = a[13] & g[14786];
assign g[31169] = b[13] & g[14786];
assign g[22979] = a[13] & g[14787];
assign g[31170] = b[13] & g[14787];
assign g[22980] = a[13] & g[14788];
assign g[31171] = b[13] & g[14788];
assign g[22981] = a[13] & g[14789];
assign g[31172] = b[13] & g[14789];
assign g[22982] = a[13] & g[14790];
assign g[31173] = b[13] & g[14790];
assign g[22983] = a[13] & g[14791];
assign g[31174] = b[13] & g[14791];
assign g[22984] = a[13] & g[14792];
assign g[31175] = b[13] & g[14792];
assign g[22985] = a[13] & g[14793];
assign g[31176] = b[13] & g[14793];
assign g[22986] = a[13] & g[14794];
assign g[31177] = b[13] & g[14794];
assign g[22987] = a[13] & g[14795];
assign g[31178] = b[13] & g[14795];
assign g[22988] = a[13] & g[14796];
assign g[31179] = b[13] & g[14796];
assign g[22989] = a[13] & g[14797];
assign g[31180] = b[13] & g[14797];
assign g[22990] = a[13] & g[14798];
assign g[31181] = b[13] & g[14798];
assign g[22991] = a[13] & g[14799];
assign g[31182] = b[13] & g[14799];
assign g[22992] = a[13] & g[14800];
assign g[31183] = b[13] & g[14800];
assign g[22993] = a[13] & g[14801];
assign g[31184] = b[13] & g[14801];
assign g[22994] = a[13] & g[14802];
assign g[31185] = b[13] & g[14802];
assign g[22995] = a[13] & g[14803];
assign g[31186] = b[13] & g[14803];
assign g[22996] = a[13] & g[14804];
assign g[31187] = b[13] & g[14804];
assign g[22997] = a[13] & g[14805];
assign g[31188] = b[13] & g[14805];
assign g[22998] = a[13] & g[14806];
assign g[31189] = b[13] & g[14806];
assign g[22999] = a[13] & g[14807];
assign g[31190] = b[13] & g[14807];
assign g[23000] = a[13] & g[14808];
assign g[31191] = b[13] & g[14808];
assign g[23001] = a[13] & g[14809];
assign g[31192] = b[13] & g[14809];
assign g[23002] = a[13] & g[14810];
assign g[31193] = b[13] & g[14810];
assign g[23003] = a[13] & g[14811];
assign g[31194] = b[13] & g[14811];
assign g[23004] = a[13] & g[14812];
assign g[31195] = b[13] & g[14812];
assign g[23005] = a[13] & g[14813];
assign g[31196] = b[13] & g[14813];
assign g[23006] = a[13] & g[14814];
assign g[31197] = b[13] & g[14814];
assign g[23007] = a[13] & g[14815];
assign g[31198] = b[13] & g[14815];
assign g[23008] = a[13] & g[14816];
assign g[31199] = b[13] & g[14816];
assign g[23009] = a[13] & g[14817];
assign g[31200] = b[13] & g[14817];
assign g[23010] = a[13] & g[14818];
assign g[31201] = b[13] & g[14818];
assign g[23011] = a[13] & g[14819];
assign g[31202] = b[13] & g[14819];
assign g[23012] = a[13] & g[14820];
assign g[31203] = b[13] & g[14820];
assign g[23013] = a[13] & g[14821];
assign g[31204] = b[13] & g[14821];
assign g[23014] = a[13] & g[14822];
assign g[31205] = b[13] & g[14822];
assign g[23015] = a[13] & g[14823];
assign g[31206] = b[13] & g[14823];
assign g[23016] = a[13] & g[14824];
assign g[31207] = b[13] & g[14824];
assign g[23017] = a[13] & g[14825];
assign g[31208] = b[13] & g[14825];
assign g[23018] = a[13] & g[14826];
assign g[31209] = b[13] & g[14826];
assign g[23019] = a[13] & g[14827];
assign g[31210] = b[13] & g[14827];
assign g[23020] = a[13] & g[14828];
assign g[31211] = b[13] & g[14828];
assign g[23021] = a[13] & g[14829];
assign g[31212] = b[13] & g[14829];
assign g[23022] = a[13] & g[14830];
assign g[31213] = b[13] & g[14830];
assign g[23023] = a[13] & g[14831];
assign g[31214] = b[13] & g[14831];
assign g[23024] = a[13] & g[14832];
assign g[31215] = b[13] & g[14832];
assign g[23025] = a[13] & g[14833];
assign g[31216] = b[13] & g[14833];
assign g[23026] = a[13] & g[14834];
assign g[31217] = b[13] & g[14834];
assign g[23027] = a[13] & g[14835];
assign g[31218] = b[13] & g[14835];
assign g[23028] = a[13] & g[14836];
assign g[31219] = b[13] & g[14836];
assign g[23029] = a[13] & g[14837];
assign g[31220] = b[13] & g[14837];
assign g[23030] = a[13] & g[14838];
assign g[31221] = b[13] & g[14838];
assign g[23031] = a[13] & g[14839];
assign g[31222] = b[13] & g[14839];
assign g[23032] = a[13] & g[14840];
assign g[31223] = b[13] & g[14840];
assign g[23033] = a[13] & g[14841];
assign g[31224] = b[13] & g[14841];
assign g[23034] = a[13] & g[14842];
assign g[31225] = b[13] & g[14842];
assign g[23035] = a[13] & g[14843];
assign g[31226] = b[13] & g[14843];
assign g[23036] = a[13] & g[14844];
assign g[31227] = b[13] & g[14844];
assign g[23037] = a[13] & g[14845];
assign g[31228] = b[13] & g[14845];
assign g[23038] = a[13] & g[14846];
assign g[31229] = b[13] & g[14846];
assign g[23039] = a[13] & g[14847];
assign g[31230] = b[13] & g[14847];
assign g[23040] = a[13] & g[14848];
assign g[31231] = b[13] & g[14848];
assign g[23041] = a[13] & g[14849];
assign g[31232] = b[13] & g[14849];
assign g[23042] = a[13] & g[14850];
assign g[31233] = b[13] & g[14850];
assign g[23043] = a[13] & g[14851];
assign g[31234] = b[13] & g[14851];
assign g[23044] = a[13] & g[14852];
assign g[31235] = b[13] & g[14852];
assign g[23045] = a[13] & g[14853];
assign g[31236] = b[13] & g[14853];
assign g[23046] = a[13] & g[14854];
assign g[31237] = b[13] & g[14854];
assign g[23047] = a[13] & g[14855];
assign g[31238] = b[13] & g[14855];
assign g[23048] = a[13] & g[14856];
assign g[31239] = b[13] & g[14856];
assign g[23049] = a[13] & g[14857];
assign g[31240] = b[13] & g[14857];
assign g[23050] = a[13] & g[14858];
assign g[31241] = b[13] & g[14858];
assign g[23051] = a[13] & g[14859];
assign g[31242] = b[13] & g[14859];
assign g[23052] = a[13] & g[14860];
assign g[31243] = b[13] & g[14860];
assign g[23053] = a[13] & g[14861];
assign g[31244] = b[13] & g[14861];
assign g[23054] = a[13] & g[14862];
assign g[31245] = b[13] & g[14862];
assign g[23055] = a[13] & g[14863];
assign g[31246] = b[13] & g[14863];
assign g[23056] = a[13] & g[14864];
assign g[31247] = b[13] & g[14864];
assign g[23057] = a[13] & g[14865];
assign g[31248] = b[13] & g[14865];
assign g[23058] = a[13] & g[14866];
assign g[31249] = b[13] & g[14866];
assign g[23059] = a[13] & g[14867];
assign g[31250] = b[13] & g[14867];
assign g[23060] = a[13] & g[14868];
assign g[31251] = b[13] & g[14868];
assign g[23061] = a[13] & g[14869];
assign g[31252] = b[13] & g[14869];
assign g[23062] = a[13] & g[14870];
assign g[31253] = b[13] & g[14870];
assign g[23063] = a[13] & g[14871];
assign g[31254] = b[13] & g[14871];
assign g[23064] = a[13] & g[14872];
assign g[31255] = b[13] & g[14872];
assign g[23065] = a[13] & g[14873];
assign g[31256] = b[13] & g[14873];
assign g[23066] = a[13] & g[14874];
assign g[31257] = b[13] & g[14874];
assign g[23067] = a[13] & g[14875];
assign g[31258] = b[13] & g[14875];
assign g[23068] = a[13] & g[14876];
assign g[31259] = b[13] & g[14876];
assign g[23069] = a[13] & g[14877];
assign g[31260] = b[13] & g[14877];
assign g[23070] = a[13] & g[14878];
assign g[31261] = b[13] & g[14878];
assign g[23071] = a[13] & g[14879];
assign g[31262] = b[13] & g[14879];
assign g[23072] = a[13] & g[14880];
assign g[31263] = b[13] & g[14880];
assign g[23073] = a[13] & g[14881];
assign g[31264] = b[13] & g[14881];
assign g[23074] = a[13] & g[14882];
assign g[31265] = b[13] & g[14882];
assign g[23075] = a[13] & g[14883];
assign g[31266] = b[13] & g[14883];
assign g[23076] = a[13] & g[14884];
assign g[31267] = b[13] & g[14884];
assign g[23077] = a[13] & g[14885];
assign g[31268] = b[13] & g[14885];
assign g[23078] = a[13] & g[14886];
assign g[31269] = b[13] & g[14886];
assign g[23079] = a[13] & g[14887];
assign g[31270] = b[13] & g[14887];
assign g[23080] = a[13] & g[14888];
assign g[31271] = b[13] & g[14888];
assign g[23081] = a[13] & g[14889];
assign g[31272] = b[13] & g[14889];
assign g[23082] = a[13] & g[14890];
assign g[31273] = b[13] & g[14890];
assign g[23083] = a[13] & g[14891];
assign g[31274] = b[13] & g[14891];
assign g[23084] = a[13] & g[14892];
assign g[31275] = b[13] & g[14892];
assign g[23085] = a[13] & g[14893];
assign g[31276] = b[13] & g[14893];
assign g[23086] = a[13] & g[14894];
assign g[31277] = b[13] & g[14894];
assign g[23087] = a[13] & g[14895];
assign g[31278] = b[13] & g[14895];
assign g[23088] = a[13] & g[14896];
assign g[31279] = b[13] & g[14896];
assign g[23089] = a[13] & g[14897];
assign g[31280] = b[13] & g[14897];
assign g[23090] = a[13] & g[14898];
assign g[31281] = b[13] & g[14898];
assign g[23091] = a[13] & g[14899];
assign g[31282] = b[13] & g[14899];
assign g[23092] = a[13] & g[14900];
assign g[31283] = b[13] & g[14900];
assign g[23093] = a[13] & g[14901];
assign g[31284] = b[13] & g[14901];
assign g[23094] = a[13] & g[14902];
assign g[31285] = b[13] & g[14902];
assign g[23095] = a[13] & g[14903];
assign g[31286] = b[13] & g[14903];
assign g[23096] = a[13] & g[14904];
assign g[31287] = b[13] & g[14904];
assign g[23097] = a[13] & g[14905];
assign g[31288] = b[13] & g[14905];
assign g[23098] = a[13] & g[14906];
assign g[31289] = b[13] & g[14906];
assign g[23099] = a[13] & g[14907];
assign g[31290] = b[13] & g[14907];
assign g[23100] = a[13] & g[14908];
assign g[31291] = b[13] & g[14908];
assign g[23101] = a[13] & g[14909];
assign g[31292] = b[13] & g[14909];
assign g[23102] = a[13] & g[14910];
assign g[31293] = b[13] & g[14910];
assign g[23103] = a[13] & g[14911];
assign g[31294] = b[13] & g[14911];
assign g[23104] = a[13] & g[14912];
assign g[31295] = b[13] & g[14912];
assign g[23105] = a[13] & g[14913];
assign g[31296] = b[13] & g[14913];
assign g[23106] = a[13] & g[14914];
assign g[31297] = b[13] & g[14914];
assign g[23107] = a[13] & g[14915];
assign g[31298] = b[13] & g[14915];
assign g[23108] = a[13] & g[14916];
assign g[31299] = b[13] & g[14916];
assign g[23109] = a[13] & g[14917];
assign g[31300] = b[13] & g[14917];
assign g[23110] = a[13] & g[14918];
assign g[31301] = b[13] & g[14918];
assign g[23111] = a[13] & g[14919];
assign g[31302] = b[13] & g[14919];
assign g[23112] = a[13] & g[14920];
assign g[31303] = b[13] & g[14920];
assign g[23113] = a[13] & g[14921];
assign g[31304] = b[13] & g[14921];
assign g[23114] = a[13] & g[14922];
assign g[31305] = b[13] & g[14922];
assign g[23115] = a[13] & g[14923];
assign g[31306] = b[13] & g[14923];
assign g[23116] = a[13] & g[14924];
assign g[31307] = b[13] & g[14924];
assign g[23117] = a[13] & g[14925];
assign g[31308] = b[13] & g[14925];
assign g[23118] = a[13] & g[14926];
assign g[31309] = b[13] & g[14926];
assign g[23119] = a[13] & g[14927];
assign g[31310] = b[13] & g[14927];
assign g[23120] = a[13] & g[14928];
assign g[31311] = b[13] & g[14928];
assign g[23121] = a[13] & g[14929];
assign g[31312] = b[13] & g[14929];
assign g[23122] = a[13] & g[14930];
assign g[31313] = b[13] & g[14930];
assign g[23123] = a[13] & g[14931];
assign g[31314] = b[13] & g[14931];
assign g[23124] = a[13] & g[14932];
assign g[31315] = b[13] & g[14932];
assign g[23125] = a[13] & g[14933];
assign g[31316] = b[13] & g[14933];
assign g[23126] = a[13] & g[14934];
assign g[31317] = b[13] & g[14934];
assign g[23127] = a[13] & g[14935];
assign g[31318] = b[13] & g[14935];
assign g[23128] = a[13] & g[14936];
assign g[31319] = b[13] & g[14936];
assign g[23129] = a[13] & g[14937];
assign g[31320] = b[13] & g[14937];
assign g[23130] = a[13] & g[14938];
assign g[31321] = b[13] & g[14938];
assign g[23131] = a[13] & g[14939];
assign g[31322] = b[13] & g[14939];
assign g[23132] = a[13] & g[14940];
assign g[31323] = b[13] & g[14940];
assign g[23133] = a[13] & g[14941];
assign g[31324] = b[13] & g[14941];
assign g[23134] = a[13] & g[14942];
assign g[31325] = b[13] & g[14942];
assign g[23135] = a[13] & g[14943];
assign g[31326] = b[13] & g[14943];
assign g[23136] = a[13] & g[14944];
assign g[31327] = b[13] & g[14944];
assign g[23137] = a[13] & g[14945];
assign g[31328] = b[13] & g[14945];
assign g[23138] = a[13] & g[14946];
assign g[31329] = b[13] & g[14946];
assign g[23139] = a[13] & g[14947];
assign g[31330] = b[13] & g[14947];
assign g[23140] = a[13] & g[14948];
assign g[31331] = b[13] & g[14948];
assign g[23141] = a[13] & g[14949];
assign g[31332] = b[13] & g[14949];
assign g[23142] = a[13] & g[14950];
assign g[31333] = b[13] & g[14950];
assign g[23143] = a[13] & g[14951];
assign g[31334] = b[13] & g[14951];
assign g[23144] = a[13] & g[14952];
assign g[31335] = b[13] & g[14952];
assign g[23145] = a[13] & g[14953];
assign g[31336] = b[13] & g[14953];
assign g[23146] = a[13] & g[14954];
assign g[31337] = b[13] & g[14954];
assign g[23147] = a[13] & g[14955];
assign g[31338] = b[13] & g[14955];
assign g[23148] = a[13] & g[14956];
assign g[31339] = b[13] & g[14956];
assign g[23149] = a[13] & g[14957];
assign g[31340] = b[13] & g[14957];
assign g[23150] = a[13] & g[14958];
assign g[31341] = b[13] & g[14958];
assign g[23151] = a[13] & g[14959];
assign g[31342] = b[13] & g[14959];
assign g[23152] = a[13] & g[14960];
assign g[31343] = b[13] & g[14960];
assign g[23153] = a[13] & g[14961];
assign g[31344] = b[13] & g[14961];
assign g[23154] = a[13] & g[14962];
assign g[31345] = b[13] & g[14962];
assign g[23155] = a[13] & g[14963];
assign g[31346] = b[13] & g[14963];
assign g[23156] = a[13] & g[14964];
assign g[31347] = b[13] & g[14964];
assign g[23157] = a[13] & g[14965];
assign g[31348] = b[13] & g[14965];
assign g[23158] = a[13] & g[14966];
assign g[31349] = b[13] & g[14966];
assign g[23159] = a[13] & g[14967];
assign g[31350] = b[13] & g[14967];
assign g[23160] = a[13] & g[14968];
assign g[31351] = b[13] & g[14968];
assign g[23161] = a[13] & g[14969];
assign g[31352] = b[13] & g[14969];
assign g[23162] = a[13] & g[14970];
assign g[31353] = b[13] & g[14970];
assign g[23163] = a[13] & g[14971];
assign g[31354] = b[13] & g[14971];
assign g[23164] = a[13] & g[14972];
assign g[31355] = b[13] & g[14972];
assign g[23165] = a[13] & g[14973];
assign g[31356] = b[13] & g[14973];
assign g[23166] = a[13] & g[14974];
assign g[31357] = b[13] & g[14974];
assign g[23167] = a[13] & g[14975];
assign g[31358] = b[13] & g[14975];
assign g[23168] = a[13] & g[14976];
assign g[31359] = b[13] & g[14976];
assign g[23169] = a[13] & g[14977];
assign g[31360] = b[13] & g[14977];
assign g[23170] = a[13] & g[14978];
assign g[31361] = b[13] & g[14978];
assign g[23171] = a[13] & g[14979];
assign g[31362] = b[13] & g[14979];
assign g[23172] = a[13] & g[14980];
assign g[31363] = b[13] & g[14980];
assign g[23173] = a[13] & g[14981];
assign g[31364] = b[13] & g[14981];
assign g[23174] = a[13] & g[14982];
assign g[31365] = b[13] & g[14982];
assign g[23175] = a[13] & g[14983];
assign g[31366] = b[13] & g[14983];
assign g[23176] = a[13] & g[14984];
assign g[31367] = b[13] & g[14984];
assign g[23177] = a[13] & g[14985];
assign g[31368] = b[13] & g[14985];
assign g[23178] = a[13] & g[14986];
assign g[31369] = b[13] & g[14986];
assign g[23179] = a[13] & g[14987];
assign g[31370] = b[13] & g[14987];
assign g[23180] = a[13] & g[14988];
assign g[31371] = b[13] & g[14988];
assign g[23181] = a[13] & g[14989];
assign g[31372] = b[13] & g[14989];
assign g[23182] = a[13] & g[14990];
assign g[31373] = b[13] & g[14990];
assign g[23183] = a[13] & g[14991];
assign g[31374] = b[13] & g[14991];
assign g[23184] = a[13] & g[14992];
assign g[31375] = b[13] & g[14992];
assign g[23185] = a[13] & g[14993];
assign g[31376] = b[13] & g[14993];
assign g[23186] = a[13] & g[14994];
assign g[31377] = b[13] & g[14994];
assign g[23187] = a[13] & g[14995];
assign g[31378] = b[13] & g[14995];
assign g[23188] = a[13] & g[14996];
assign g[31379] = b[13] & g[14996];
assign g[23189] = a[13] & g[14997];
assign g[31380] = b[13] & g[14997];
assign g[23190] = a[13] & g[14998];
assign g[31381] = b[13] & g[14998];
assign g[23191] = a[13] & g[14999];
assign g[31382] = b[13] & g[14999];
assign g[23192] = a[13] & g[15000];
assign g[31383] = b[13] & g[15000];
assign g[23193] = a[13] & g[15001];
assign g[31384] = b[13] & g[15001];
assign g[23194] = a[13] & g[15002];
assign g[31385] = b[13] & g[15002];
assign g[23195] = a[13] & g[15003];
assign g[31386] = b[13] & g[15003];
assign g[23196] = a[13] & g[15004];
assign g[31387] = b[13] & g[15004];
assign g[23197] = a[13] & g[15005];
assign g[31388] = b[13] & g[15005];
assign g[23198] = a[13] & g[15006];
assign g[31389] = b[13] & g[15006];
assign g[23199] = a[13] & g[15007];
assign g[31390] = b[13] & g[15007];
assign g[23200] = a[13] & g[15008];
assign g[31391] = b[13] & g[15008];
assign g[23201] = a[13] & g[15009];
assign g[31392] = b[13] & g[15009];
assign g[23202] = a[13] & g[15010];
assign g[31393] = b[13] & g[15010];
assign g[23203] = a[13] & g[15011];
assign g[31394] = b[13] & g[15011];
assign g[23204] = a[13] & g[15012];
assign g[31395] = b[13] & g[15012];
assign g[23205] = a[13] & g[15013];
assign g[31396] = b[13] & g[15013];
assign g[23206] = a[13] & g[15014];
assign g[31397] = b[13] & g[15014];
assign g[23207] = a[13] & g[15015];
assign g[31398] = b[13] & g[15015];
assign g[23208] = a[13] & g[15016];
assign g[31399] = b[13] & g[15016];
assign g[23209] = a[13] & g[15017];
assign g[31400] = b[13] & g[15017];
assign g[23210] = a[13] & g[15018];
assign g[31401] = b[13] & g[15018];
assign g[23211] = a[13] & g[15019];
assign g[31402] = b[13] & g[15019];
assign g[23212] = a[13] & g[15020];
assign g[31403] = b[13] & g[15020];
assign g[23213] = a[13] & g[15021];
assign g[31404] = b[13] & g[15021];
assign g[23214] = a[13] & g[15022];
assign g[31405] = b[13] & g[15022];
assign g[23215] = a[13] & g[15023];
assign g[31406] = b[13] & g[15023];
assign g[23216] = a[13] & g[15024];
assign g[31407] = b[13] & g[15024];
assign g[23217] = a[13] & g[15025];
assign g[31408] = b[13] & g[15025];
assign g[23218] = a[13] & g[15026];
assign g[31409] = b[13] & g[15026];
assign g[23219] = a[13] & g[15027];
assign g[31410] = b[13] & g[15027];
assign g[23220] = a[13] & g[15028];
assign g[31411] = b[13] & g[15028];
assign g[23221] = a[13] & g[15029];
assign g[31412] = b[13] & g[15029];
assign g[23222] = a[13] & g[15030];
assign g[31413] = b[13] & g[15030];
assign g[23223] = a[13] & g[15031];
assign g[31414] = b[13] & g[15031];
assign g[23224] = a[13] & g[15032];
assign g[31415] = b[13] & g[15032];
assign g[23225] = a[13] & g[15033];
assign g[31416] = b[13] & g[15033];
assign g[23226] = a[13] & g[15034];
assign g[31417] = b[13] & g[15034];
assign g[23227] = a[13] & g[15035];
assign g[31418] = b[13] & g[15035];
assign g[23228] = a[13] & g[15036];
assign g[31419] = b[13] & g[15036];
assign g[23229] = a[13] & g[15037];
assign g[31420] = b[13] & g[15037];
assign g[23230] = a[13] & g[15038];
assign g[31421] = b[13] & g[15038];
assign g[23231] = a[13] & g[15039];
assign g[31422] = b[13] & g[15039];
assign g[23232] = a[13] & g[15040];
assign g[31423] = b[13] & g[15040];
assign g[23233] = a[13] & g[15041];
assign g[31424] = b[13] & g[15041];
assign g[23234] = a[13] & g[15042];
assign g[31425] = b[13] & g[15042];
assign g[23235] = a[13] & g[15043];
assign g[31426] = b[13] & g[15043];
assign g[23236] = a[13] & g[15044];
assign g[31427] = b[13] & g[15044];
assign g[23237] = a[13] & g[15045];
assign g[31428] = b[13] & g[15045];
assign g[23238] = a[13] & g[15046];
assign g[31429] = b[13] & g[15046];
assign g[23239] = a[13] & g[15047];
assign g[31430] = b[13] & g[15047];
assign g[23240] = a[13] & g[15048];
assign g[31431] = b[13] & g[15048];
assign g[23241] = a[13] & g[15049];
assign g[31432] = b[13] & g[15049];
assign g[23242] = a[13] & g[15050];
assign g[31433] = b[13] & g[15050];
assign g[23243] = a[13] & g[15051];
assign g[31434] = b[13] & g[15051];
assign g[23244] = a[13] & g[15052];
assign g[31435] = b[13] & g[15052];
assign g[23245] = a[13] & g[15053];
assign g[31436] = b[13] & g[15053];
assign g[23246] = a[13] & g[15054];
assign g[31437] = b[13] & g[15054];
assign g[23247] = a[13] & g[15055];
assign g[31438] = b[13] & g[15055];
assign g[23248] = a[13] & g[15056];
assign g[31439] = b[13] & g[15056];
assign g[23249] = a[13] & g[15057];
assign g[31440] = b[13] & g[15057];
assign g[23250] = a[13] & g[15058];
assign g[31441] = b[13] & g[15058];
assign g[23251] = a[13] & g[15059];
assign g[31442] = b[13] & g[15059];
assign g[23252] = a[13] & g[15060];
assign g[31443] = b[13] & g[15060];
assign g[23253] = a[13] & g[15061];
assign g[31444] = b[13] & g[15061];
assign g[23254] = a[13] & g[15062];
assign g[31445] = b[13] & g[15062];
assign g[23255] = a[13] & g[15063];
assign g[31446] = b[13] & g[15063];
assign g[23256] = a[13] & g[15064];
assign g[31447] = b[13] & g[15064];
assign g[23257] = a[13] & g[15065];
assign g[31448] = b[13] & g[15065];
assign g[23258] = a[13] & g[15066];
assign g[31449] = b[13] & g[15066];
assign g[23259] = a[13] & g[15067];
assign g[31450] = b[13] & g[15067];
assign g[23260] = a[13] & g[15068];
assign g[31451] = b[13] & g[15068];
assign g[23261] = a[13] & g[15069];
assign g[31452] = b[13] & g[15069];
assign g[23262] = a[13] & g[15070];
assign g[31453] = b[13] & g[15070];
assign g[23263] = a[13] & g[15071];
assign g[31454] = b[13] & g[15071];
assign g[23264] = a[13] & g[15072];
assign g[31455] = b[13] & g[15072];
assign g[23265] = a[13] & g[15073];
assign g[31456] = b[13] & g[15073];
assign g[23266] = a[13] & g[15074];
assign g[31457] = b[13] & g[15074];
assign g[23267] = a[13] & g[15075];
assign g[31458] = b[13] & g[15075];
assign g[23268] = a[13] & g[15076];
assign g[31459] = b[13] & g[15076];
assign g[23269] = a[13] & g[15077];
assign g[31460] = b[13] & g[15077];
assign g[23270] = a[13] & g[15078];
assign g[31461] = b[13] & g[15078];
assign g[23271] = a[13] & g[15079];
assign g[31462] = b[13] & g[15079];
assign g[23272] = a[13] & g[15080];
assign g[31463] = b[13] & g[15080];
assign g[23273] = a[13] & g[15081];
assign g[31464] = b[13] & g[15081];
assign g[23274] = a[13] & g[15082];
assign g[31465] = b[13] & g[15082];
assign g[23275] = a[13] & g[15083];
assign g[31466] = b[13] & g[15083];
assign g[23276] = a[13] & g[15084];
assign g[31467] = b[13] & g[15084];
assign g[23277] = a[13] & g[15085];
assign g[31468] = b[13] & g[15085];
assign g[23278] = a[13] & g[15086];
assign g[31469] = b[13] & g[15086];
assign g[23279] = a[13] & g[15087];
assign g[31470] = b[13] & g[15087];
assign g[23280] = a[13] & g[15088];
assign g[31471] = b[13] & g[15088];
assign g[23281] = a[13] & g[15089];
assign g[31472] = b[13] & g[15089];
assign g[23282] = a[13] & g[15090];
assign g[31473] = b[13] & g[15090];
assign g[23283] = a[13] & g[15091];
assign g[31474] = b[13] & g[15091];
assign g[23284] = a[13] & g[15092];
assign g[31475] = b[13] & g[15092];
assign g[23285] = a[13] & g[15093];
assign g[31476] = b[13] & g[15093];
assign g[23286] = a[13] & g[15094];
assign g[31477] = b[13] & g[15094];
assign g[23287] = a[13] & g[15095];
assign g[31478] = b[13] & g[15095];
assign g[23288] = a[13] & g[15096];
assign g[31479] = b[13] & g[15096];
assign g[23289] = a[13] & g[15097];
assign g[31480] = b[13] & g[15097];
assign g[23290] = a[13] & g[15098];
assign g[31481] = b[13] & g[15098];
assign g[23291] = a[13] & g[15099];
assign g[31482] = b[13] & g[15099];
assign g[23292] = a[13] & g[15100];
assign g[31483] = b[13] & g[15100];
assign g[23293] = a[13] & g[15101];
assign g[31484] = b[13] & g[15101];
assign g[23294] = a[13] & g[15102];
assign g[31485] = b[13] & g[15102];
assign g[23295] = a[13] & g[15103];
assign g[31486] = b[13] & g[15103];
assign g[23296] = a[13] & g[15104];
assign g[31487] = b[13] & g[15104];
assign g[23297] = a[13] & g[15105];
assign g[31488] = b[13] & g[15105];
assign g[23298] = a[13] & g[15106];
assign g[31489] = b[13] & g[15106];
assign g[23299] = a[13] & g[15107];
assign g[31490] = b[13] & g[15107];
assign g[23300] = a[13] & g[15108];
assign g[31491] = b[13] & g[15108];
assign g[23301] = a[13] & g[15109];
assign g[31492] = b[13] & g[15109];
assign g[23302] = a[13] & g[15110];
assign g[31493] = b[13] & g[15110];
assign g[23303] = a[13] & g[15111];
assign g[31494] = b[13] & g[15111];
assign g[23304] = a[13] & g[15112];
assign g[31495] = b[13] & g[15112];
assign g[23305] = a[13] & g[15113];
assign g[31496] = b[13] & g[15113];
assign g[23306] = a[13] & g[15114];
assign g[31497] = b[13] & g[15114];
assign g[23307] = a[13] & g[15115];
assign g[31498] = b[13] & g[15115];
assign g[23308] = a[13] & g[15116];
assign g[31499] = b[13] & g[15116];
assign g[23309] = a[13] & g[15117];
assign g[31500] = b[13] & g[15117];
assign g[23310] = a[13] & g[15118];
assign g[31501] = b[13] & g[15118];
assign g[23311] = a[13] & g[15119];
assign g[31502] = b[13] & g[15119];
assign g[23312] = a[13] & g[15120];
assign g[31503] = b[13] & g[15120];
assign g[23313] = a[13] & g[15121];
assign g[31504] = b[13] & g[15121];
assign g[23314] = a[13] & g[15122];
assign g[31505] = b[13] & g[15122];
assign g[23315] = a[13] & g[15123];
assign g[31506] = b[13] & g[15123];
assign g[23316] = a[13] & g[15124];
assign g[31507] = b[13] & g[15124];
assign g[23317] = a[13] & g[15125];
assign g[31508] = b[13] & g[15125];
assign g[23318] = a[13] & g[15126];
assign g[31509] = b[13] & g[15126];
assign g[23319] = a[13] & g[15127];
assign g[31510] = b[13] & g[15127];
assign g[23320] = a[13] & g[15128];
assign g[31511] = b[13] & g[15128];
assign g[23321] = a[13] & g[15129];
assign g[31512] = b[13] & g[15129];
assign g[23322] = a[13] & g[15130];
assign g[31513] = b[13] & g[15130];
assign g[23323] = a[13] & g[15131];
assign g[31514] = b[13] & g[15131];
assign g[23324] = a[13] & g[15132];
assign g[31515] = b[13] & g[15132];
assign g[23325] = a[13] & g[15133];
assign g[31516] = b[13] & g[15133];
assign g[23326] = a[13] & g[15134];
assign g[31517] = b[13] & g[15134];
assign g[23327] = a[13] & g[15135];
assign g[31518] = b[13] & g[15135];
assign g[23328] = a[13] & g[15136];
assign g[31519] = b[13] & g[15136];
assign g[23329] = a[13] & g[15137];
assign g[31520] = b[13] & g[15137];
assign g[23330] = a[13] & g[15138];
assign g[31521] = b[13] & g[15138];
assign g[23331] = a[13] & g[15139];
assign g[31522] = b[13] & g[15139];
assign g[23332] = a[13] & g[15140];
assign g[31523] = b[13] & g[15140];
assign g[23333] = a[13] & g[15141];
assign g[31524] = b[13] & g[15141];
assign g[23334] = a[13] & g[15142];
assign g[31525] = b[13] & g[15142];
assign g[23335] = a[13] & g[15143];
assign g[31526] = b[13] & g[15143];
assign g[23336] = a[13] & g[15144];
assign g[31527] = b[13] & g[15144];
assign g[23337] = a[13] & g[15145];
assign g[31528] = b[13] & g[15145];
assign g[23338] = a[13] & g[15146];
assign g[31529] = b[13] & g[15146];
assign g[23339] = a[13] & g[15147];
assign g[31530] = b[13] & g[15147];
assign g[23340] = a[13] & g[15148];
assign g[31531] = b[13] & g[15148];
assign g[23341] = a[13] & g[15149];
assign g[31532] = b[13] & g[15149];
assign g[23342] = a[13] & g[15150];
assign g[31533] = b[13] & g[15150];
assign g[23343] = a[13] & g[15151];
assign g[31534] = b[13] & g[15151];
assign g[23344] = a[13] & g[15152];
assign g[31535] = b[13] & g[15152];
assign g[23345] = a[13] & g[15153];
assign g[31536] = b[13] & g[15153];
assign g[23346] = a[13] & g[15154];
assign g[31537] = b[13] & g[15154];
assign g[23347] = a[13] & g[15155];
assign g[31538] = b[13] & g[15155];
assign g[23348] = a[13] & g[15156];
assign g[31539] = b[13] & g[15156];
assign g[23349] = a[13] & g[15157];
assign g[31540] = b[13] & g[15157];
assign g[23350] = a[13] & g[15158];
assign g[31541] = b[13] & g[15158];
assign g[23351] = a[13] & g[15159];
assign g[31542] = b[13] & g[15159];
assign g[23352] = a[13] & g[15160];
assign g[31543] = b[13] & g[15160];
assign g[23353] = a[13] & g[15161];
assign g[31544] = b[13] & g[15161];
assign g[23354] = a[13] & g[15162];
assign g[31545] = b[13] & g[15162];
assign g[23355] = a[13] & g[15163];
assign g[31546] = b[13] & g[15163];
assign g[23356] = a[13] & g[15164];
assign g[31547] = b[13] & g[15164];
assign g[23357] = a[13] & g[15165];
assign g[31548] = b[13] & g[15165];
assign g[23358] = a[13] & g[15166];
assign g[31549] = b[13] & g[15166];
assign g[23359] = a[13] & g[15167];
assign g[31550] = b[13] & g[15167];
assign g[23360] = a[13] & g[15168];
assign g[31551] = b[13] & g[15168];
assign g[23361] = a[13] & g[15169];
assign g[31552] = b[13] & g[15169];
assign g[23362] = a[13] & g[15170];
assign g[31553] = b[13] & g[15170];
assign g[23363] = a[13] & g[15171];
assign g[31554] = b[13] & g[15171];
assign g[23364] = a[13] & g[15172];
assign g[31555] = b[13] & g[15172];
assign g[23365] = a[13] & g[15173];
assign g[31556] = b[13] & g[15173];
assign g[23366] = a[13] & g[15174];
assign g[31557] = b[13] & g[15174];
assign g[23367] = a[13] & g[15175];
assign g[31558] = b[13] & g[15175];
assign g[23368] = a[13] & g[15176];
assign g[31559] = b[13] & g[15176];
assign g[23369] = a[13] & g[15177];
assign g[31560] = b[13] & g[15177];
assign g[23370] = a[13] & g[15178];
assign g[31561] = b[13] & g[15178];
assign g[23371] = a[13] & g[15179];
assign g[31562] = b[13] & g[15179];
assign g[23372] = a[13] & g[15180];
assign g[31563] = b[13] & g[15180];
assign g[23373] = a[13] & g[15181];
assign g[31564] = b[13] & g[15181];
assign g[23374] = a[13] & g[15182];
assign g[31565] = b[13] & g[15182];
assign g[23375] = a[13] & g[15183];
assign g[31566] = b[13] & g[15183];
assign g[23376] = a[13] & g[15184];
assign g[31567] = b[13] & g[15184];
assign g[23377] = a[13] & g[15185];
assign g[31568] = b[13] & g[15185];
assign g[23378] = a[13] & g[15186];
assign g[31569] = b[13] & g[15186];
assign g[23379] = a[13] & g[15187];
assign g[31570] = b[13] & g[15187];
assign g[23380] = a[13] & g[15188];
assign g[31571] = b[13] & g[15188];
assign g[23381] = a[13] & g[15189];
assign g[31572] = b[13] & g[15189];
assign g[23382] = a[13] & g[15190];
assign g[31573] = b[13] & g[15190];
assign g[23383] = a[13] & g[15191];
assign g[31574] = b[13] & g[15191];
assign g[23384] = a[13] & g[15192];
assign g[31575] = b[13] & g[15192];
assign g[23385] = a[13] & g[15193];
assign g[31576] = b[13] & g[15193];
assign g[23386] = a[13] & g[15194];
assign g[31577] = b[13] & g[15194];
assign g[23387] = a[13] & g[15195];
assign g[31578] = b[13] & g[15195];
assign g[23388] = a[13] & g[15196];
assign g[31579] = b[13] & g[15196];
assign g[23389] = a[13] & g[15197];
assign g[31580] = b[13] & g[15197];
assign g[23390] = a[13] & g[15198];
assign g[31581] = b[13] & g[15198];
assign g[23391] = a[13] & g[15199];
assign g[31582] = b[13] & g[15199];
assign g[23392] = a[13] & g[15200];
assign g[31583] = b[13] & g[15200];
assign g[23393] = a[13] & g[15201];
assign g[31584] = b[13] & g[15201];
assign g[23394] = a[13] & g[15202];
assign g[31585] = b[13] & g[15202];
assign g[23395] = a[13] & g[15203];
assign g[31586] = b[13] & g[15203];
assign g[23396] = a[13] & g[15204];
assign g[31587] = b[13] & g[15204];
assign g[23397] = a[13] & g[15205];
assign g[31588] = b[13] & g[15205];
assign g[23398] = a[13] & g[15206];
assign g[31589] = b[13] & g[15206];
assign g[23399] = a[13] & g[15207];
assign g[31590] = b[13] & g[15207];
assign g[23400] = a[13] & g[15208];
assign g[31591] = b[13] & g[15208];
assign g[23401] = a[13] & g[15209];
assign g[31592] = b[13] & g[15209];
assign g[23402] = a[13] & g[15210];
assign g[31593] = b[13] & g[15210];
assign g[23403] = a[13] & g[15211];
assign g[31594] = b[13] & g[15211];
assign g[23404] = a[13] & g[15212];
assign g[31595] = b[13] & g[15212];
assign g[23405] = a[13] & g[15213];
assign g[31596] = b[13] & g[15213];
assign g[23406] = a[13] & g[15214];
assign g[31597] = b[13] & g[15214];
assign g[23407] = a[13] & g[15215];
assign g[31598] = b[13] & g[15215];
assign g[23408] = a[13] & g[15216];
assign g[31599] = b[13] & g[15216];
assign g[23409] = a[13] & g[15217];
assign g[31600] = b[13] & g[15217];
assign g[23410] = a[13] & g[15218];
assign g[31601] = b[13] & g[15218];
assign g[23411] = a[13] & g[15219];
assign g[31602] = b[13] & g[15219];
assign g[23412] = a[13] & g[15220];
assign g[31603] = b[13] & g[15220];
assign g[23413] = a[13] & g[15221];
assign g[31604] = b[13] & g[15221];
assign g[23414] = a[13] & g[15222];
assign g[31605] = b[13] & g[15222];
assign g[23415] = a[13] & g[15223];
assign g[31606] = b[13] & g[15223];
assign g[23416] = a[13] & g[15224];
assign g[31607] = b[13] & g[15224];
assign g[23417] = a[13] & g[15225];
assign g[31608] = b[13] & g[15225];
assign g[23418] = a[13] & g[15226];
assign g[31609] = b[13] & g[15226];
assign g[23419] = a[13] & g[15227];
assign g[31610] = b[13] & g[15227];
assign g[23420] = a[13] & g[15228];
assign g[31611] = b[13] & g[15228];
assign g[23421] = a[13] & g[15229];
assign g[31612] = b[13] & g[15229];
assign g[23422] = a[13] & g[15230];
assign g[31613] = b[13] & g[15230];
assign g[23423] = a[13] & g[15231];
assign g[31614] = b[13] & g[15231];
assign g[23424] = a[13] & g[15232];
assign g[31615] = b[13] & g[15232];
assign g[23425] = a[13] & g[15233];
assign g[31616] = b[13] & g[15233];
assign g[23426] = a[13] & g[15234];
assign g[31617] = b[13] & g[15234];
assign g[23427] = a[13] & g[15235];
assign g[31618] = b[13] & g[15235];
assign g[23428] = a[13] & g[15236];
assign g[31619] = b[13] & g[15236];
assign g[23429] = a[13] & g[15237];
assign g[31620] = b[13] & g[15237];
assign g[23430] = a[13] & g[15238];
assign g[31621] = b[13] & g[15238];
assign g[23431] = a[13] & g[15239];
assign g[31622] = b[13] & g[15239];
assign g[23432] = a[13] & g[15240];
assign g[31623] = b[13] & g[15240];
assign g[23433] = a[13] & g[15241];
assign g[31624] = b[13] & g[15241];
assign g[23434] = a[13] & g[15242];
assign g[31625] = b[13] & g[15242];
assign g[23435] = a[13] & g[15243];
assign g[31626] = b[13] & g[15243];
assign g[23436] = a[13] & g[15244];
assign g[31627] = b[13] & g[15244];
assign g[23437] = a[13] & g[15245];
assign g[31628] = b[13] & g[15245];
assign g[23438] = a[13] & g[15246];
assign g[31629] = b[13] & g[15246];
assign g[23439] = a[13] & g[15247];
assign g[31630] = b[13] & g[15247];
assign g[23440] = a[13] & g[15248];
assign g[31631] = b[13] & g[15248];
assign g[23441] = a[13] & g[15249];
assign g[31632] = b[13] & g[15249];
assign g[23442] = a[13] & g[15250];
assign g[31633] = b[13] & g[15250];
assign g[23443] = a[13] & g[15251];
assign g[31634] = b[13] & g[15251];
assign g[23444] = a[13] & g[15252];
assign g[31635] = b[13] & g[15252];
assign g[23445] = a[13] & g[15253];
assign g[31636] = b[13] & g[15253];
assign g[23446] = a[13] & g[15254];
assign g[31637] = b[13] & g[15254];
assign g[23447] = a[13] & g[15255];
assign g[31638] = b[13] & g[15255];
assign g[23448] = a[13] & g[15256];
assign g[31639] = b[13] & g[15256];
assign g[23449] = a[13] & g[15257];
assign g[31640] = b[13] & g[15257];
assign g[23450] = a[13] & g[15258];
assign g[31641] = b[13] & g[15258];
assign g[23451] = a[13] & g[15259];
assign g[31642] = b[13] & g[15259];
assign g[23452] = a[13] & g[15260];
assign g[31643] = b[13] & g[15260];
assign g[23453] = a[13] & g[15261];
assign g[31644] = b[13] & g[15261];
assign g[23454] = a[13] & g[15262];
assign g[31645] = b[13] & g[15262];
assign g[23455] = a[13] & g[15263];
assign g[31646] = b[13] & g[15263];
assign g[23456] = a[13] & g[15264];
assign g[31647] = b[13] & g[15264];
assign g[23457] = a[13] & g[15265];
assign g[31648] = b[13] & g[15265];
assign g[23458] = a[13] & g[15266];
assign g[31649] = b[13] & g[15266];
assign g[23459] = a[13] & g[15267];
assign g[31650] = b[13] & g[15267];
assign g[23460] = a[13] & g[15268];
assign g[31651] = b[13] & g[15268];
assign g[23461] = a[13] & g[15269];
assign g[31652] = b[13] & g[15269];
assign g[23462] = a[13] & g[15270];
assign g[31653] = b[13] & g[15270];
assign g[23463] = a[13] & g[15271];
assign g[31654] = b[13] & g[15271];
assign g[23464] = a[13] & g[15272];
assign g[31655] = b[13] & g[15272];
assign g[23465] = a[13] & g[15273];
assign g[31656] = b[13] & g[15273];
assign g[23466] = a[13] & g[15274];
assign g[31657] = b[13] & g[15274];
assign g[23467] = a[13] & g[15275];
assign g[31658] = b[13] & g[15275];
assign g[23468] = a[13] & g[15276];
assign g[31659] = b[13] & g[15276];
assign g[23469] = a[13] & g[15277];
assign g[31660] = b[13] & g[15277];
assign g[23470] = a[13] & g[15278];
assign g[31661] = b[13] & g[15278];
assign g[23471] = a[13] & g[15279];
assign g[31662] = b[13] & g[15279];
assign g[23472] = a[13] & g[15280];
assign g[31663] = b[13] & g[15280];
assign g[23473] = a[13] & g[15281];
assign g[31664] = b[13] & g[15281];
assign g[23474] = a[13] & g[15282];
assign g[31665] = b[13] & g[15282];
assign g[23475] = a[13] & g[15283];
assign g[31666] = b[13] & g[15283];
assign g[23476] = a[13] & g[15284];
assign g[31667] = b[13] & g[15284];
assign g[23477] = a[13] & g[15285];
assign g[31668] = b[13] & g[15285];
assign g[23478] = a[13] & g[15286];
assign g[31669] = b[13] & g[15286];
assign g[23479] = a[13] & g[15287];
assign g[31670] = b[13] & g[15287];
assign g[23480] = a[13] & g[15288];
assign g[31671] = b[13] & g[15288];
assign g[23481] = a[13] & g[15289];
assign g[31672] = b[13] & g[15289];
assign g[23482] = a[13] & g[15290];
assign g[31673] = b[13] & g[15290];
assign g[23483] = a[13] & g[15291];
assign g[31674] = b[13] & g[15291];
assign g[23484] = a[13] & g[15292];
assign g[31675] = b[13] & g[15292];
assign g[23485] = a[13] & g[15293];
assign g[31676] = b[13] & g[15293];
assign g[23486] = a[13] & g[15294];
assign g[31677] = b[13] & g[15294];
assign g[23487] = a[13] & g[15295];
assign g[31678] = b[13] & g[15295];
assign g[23488] = a[13] & g[15296];
assign g[31679] = b[13] & g[15296];
assign g[23489] = a[13] & g[15297];
assign g[31680] = b[13] & g[15297];
assign g[23490] = a[13] & g[15298];
assign g[31681] = b[13] & g[15298];
assign g[23491] = a[13] & g[15299];
assign g[31682] = b[13] & g[15299];
assign g[23492] = a[13] & g[15300];
assign g[31683] = b[13] & g[15300];
assign g[23493] = a[13] & g[15301];
assign g[31684] = b[13] & g[15301];
assign g[23494] = a[13] & g[15302];
assign g[31685] = b[13] & g[15302];
assign g[23495] = a[13] & g[15303];
assign g[31686] = b[13] & g[15303];
assign g[23496] = a[13] & g[15304];
assign g[31687] = b[13] & g[15304];
assign g[23497] = a[13] & g[15305];
assign g[31688] = b[13] & g[15305];
assign g[23498] = a[13] & g[15306];
assign g[31689] = b[13] & g[15306];
assign g[23499] = a[13] & g[15307];
assign g[31690] = b[13] & g[15307];
assign g[23500] = a[13] & g[15308];
assign g[31691] = b[13] & g[15308];
assign g[23501] = a[13] & g[15309];
assign g[31692] = b[13] & g[15309];
assign g[23502] = a[13] & g[15310];
assign g[31693] = b[13] & g[15310];
assign g[23503] = a[13] & g[15311];
assign g[31694] = b[13] & g[15311];
assign g[23504] = a[13] & g[15312];
assign g[31695] = b[13] & g[15312];
assign g[23505] = a[13] & g[15313];
assign g[31696] = b[13] & g[15313];
assign g[23506] = a[13] & g[15314];
assign g[31697] = b[13] & g[15314];
assign g[23507] = a[13] & g[15315];
assign g[31698] = b[13] & g[15315];
assign g[23508] = a[13] & g[15316];
assign g[31699] = b[13] & g[15316];
assign g[23509] = a[13] & g[15317];
assign g[31700] = b[13] & g[15317];
assign g[23510] = a[13] & g[15318];
assign g[31701] = b[13] & g[15318];
assign g[23511] = a[13] & g[15319];
assign g[31702] = b[13] & g[15319];
assign g[23512] = a[13] & g[15320];
assign g[31703] = b[13] & g[15320];
assign g[23513] = a[13] & g[15321];
assign g[31704] = b[13] & g[15321];
assign g[23514] = a[13] & g[15322];
assign g[31705] = b[13] & g[15322];
assign g[23515] = a[13] & g[15323];
assign g[31706] = b[13] & g[15323];
assign g[23516] = a[13] & g[15324];
assign g[31707] = b[13] & g[15324];
assign g[23517] = a[13] & g[15325];
assign g[31708] = b[13] & g[15325];
assign g[23518] = a[13] & g[15326];
assign g[31709] = b[13] & g[15326];
assign g[23519] = a[13] & g[15327];
assign g[31710] = b[13] & g[15327];
assign g[23520] = a[13] & g[15328];
assign g[31711] = b[13] & g[15328];
assign g[23521] = a[13] & g[15329];
assign g[31712] = b[13] & g[15329];
assign g[23522] = a[13] & g[15330];
assign g[31713] = b[13] & g[15330];
assign g[23523] = a[13] & g[15331];
assign g[31714] = b[13] & g[15331];
assign g[23524] = a[13] & g[15332];
assign g[31715] = b[13] & g[15332];
assign g[23525] = a[13] & g[15333];
assign g[31716] = b[13] & g[15333];
assign g[23526] = a[13] & g[15334];
assign g[31717] = b[13] & g[15334];
assign g[23527] = a[13] & g[15335];
assign g[31718] = b[13] & g[15335];
assign g[23528] = a[13] & g[15336];
assign g[31719] = b[13] & g[15336];
assign g[23529] = a[13] & g[15337];
assign g[31720] = b[13] & g[15337];
assign g[23530] = a[13] & g[15338];
assign g[31721] = b[13] & g[15338];
assign g[23531] = a[13] & g[15339];
assign g[31722] = b[13] & g[15339];
assign g[23532] = a[13] & g[15340];
assign g[31723] = b[13] & g[15340];
assign g[23533] = a[13] & g[15341];
assign g[31724] = b[13] & g[15341];
assign g[23534] = a[13] & g[15342];
assign g[31725] = b[13] & g[15342];
assign g[23535] = a[13] & g[15343];
assign g[31726] = b[13] & g[15343];
assign g[23536] = a[13] & g[15344];
assign g[31727] = b[13] & g[15344];
assign g[23537] = a[13] & g[15345];
assign g[31728] = b[13] & g[15345];
assign g[23538] = a[13] & g[15346];
assign g[31729] = b[13] & g[15346];
assign g[23539] = a[13] & g[15347];
assign g[31730] = b[13] & g[15347];
assign g[23540] = a[13] & g[15348];
assign g[31731] = b[13] & g[15348];
assign g[23541] = a[13] & g[15349];
assign g[31732] = b[13] & g[15349];
assign g[23542] = a[13] & g[15350];
assign g[31733] = b[13] & g[15350];
assign g[23543] = a[13] & g[15351];
assign g[31734] = b[13] & g[15351];
assign g[23544] = a[13] & g[15352];
assign g[31735] = b[13] & g[15352];
assign g[23545] = a[13] & g[15353];
assign g[31736] = b[13] & g[15353];
assign g[23546] = a[13] & g[15354];
assign g[31737] = b[13] & g[15354];
assign g[23547] = a[13] & g[15355];
assign g[31738] = b[13] & g[15355];
assign g[23548] = a[13] & g[15356];
assign g[31739] = b[13] & g[15356];
assign g[23549] = a[13] & g[15357];
assign g[31740] = b[13] & g[15357];
assign g[23550] = a[13] & g[15358];
assign g[31741] = b[13] & g[15358];
assign g[23551] = a[13] & g[15359];
assign g[31742] = b[13] & g[15359];
assign g[23552] = a[13] & g[15360];
assign g[31743] = b[13] & g[15360];
assign g[23553] = a[13] & g[15361];
assign g[31744] = b[13] & g[15361];
assign g[23554] = a[13] & g[15362];
assign g[31745] = b[13] & g[15362];
assign g[23555] = a[13] & g[15363];
assign g[31746] = b[13] & g[15363];
assign g[23556] = a[13] & g[15364];
assign g[31747] = b[13] & g[15364];
assign g[23557] = a[13] & g[15365];
assign g[31748] = b[13] & g[15365];
assign g[23558] = a[13] & g[15366];
assign g[31749] = b[13] & g[15366];
assign g[23559] = a[13] & g[15367];
assign g[31750] = b[13] & g[15367];
assign g[23560] = a[13] & g[15368];
assign g[31751] = b[13] & g[15368];
assign g[23561] = a[13] & g[15369];
assign g[31752] = b[13] & g[15369];
assign g[23562] = a[13] & g[15370];
assign g[31753] = b[13] & g[15370];
assign g[23563] = a[13] & g[15371];
assign g[31754] = b[13] & g[15371];
assign g[23564] = a[13] & g[15372];
assign g[31755] = b[13] & g[15372];
assign g[23565] = a[13] & g[15373];
assign g[31756] = b[13] & g[15373];
assign g[23566] = a[13] & g[15374];
assign g[31757] = b[13] & g[15374];
assign g[23567] = a[13] & g[15375];
assign g[31758] = b[13] & g[15375];
assign g[23568] = a[13] & g[15376];
assign g[31759] = b[13] & g[15376];
assign g[23569] = a[13] & g[15377];
assign g[31760] = b[13] & g[15377];
assign g[23570] = a[13] & g[15378];
assign g[31761] = b[13] & g[15378];
assign g[23571] = a[13] & g[15379];
assign g[31762] = b[13] & g[15379];
assign g[23572] = a[13] & g[15380];
assign g[31763] = b[13] & g[15380];
assign g[23573] = a[13] & g[15381];
assign g[31764] = b[13] & g[15381];
assign g[23574] = a[13] & g[15382];
assign g[31765] = b[13] & g[15382];
assign g[23575] = a[13] & g[15383];
assign g[31766] = b[13] & g[15383];
assign g[23576] = a[13] & g[15384];
assign g[31767] = b[13] & g[15384];
assign g[23577] = a[13] & g[15385];
assign g[31768] = b[13] & g[15385];
assign g[23578] = a[13] & g[15386];
assign g[31769] = b[13] & g[15386];
assign g[23579] = a[13] & g[15387];
assign g[31770] = b[13] & g[15387];
assign g[23580] = a[13] & g[15388];
assign g[31771] = b[13] & g[15388];
assign g[23581] = a[13] & g[15389];
assign g[31772] = b[13] & g[15389];
assign g[23582] = a[13] & g[15390];
assign g[31773] = b[13] & g[15390];
assign g[23583] = a[13] & g[15391];
assign g[31774] = b[13] & g[15391];
assign g[23584] = a[13] & g[15392];
assign g[31775] = b[13] & g[15392];
assign g[23585] = a[13] & g[15393];
assign g[31776] = b[13] & g[15393];
assign g[23586] = a[13] & g[15394];
assign g[31777] = b[13] & g[15394];
assign g[23587] = a[13] & g[15395];
assign g[31778] = b[13] & g[15395];
assign g[23588] = a[13] & g[15396];
assign g[31779] = b[13] & g[15396];
assign g[23589] = a[13] & g[15397];
assign g[31780] = b[13] & g[15397];
assign g[23590] = a[13] & g[15398];
assign g[31781] = b[13] & g[15398];
assign g[23591] = a[13] & g[15399];
assign g[31782] = b[13] & g[15399];
assign g[23592] = a[13] & g[15400];
assign g[31783] = b[13] & g[15400];
assign g[23593] = a[13] & g[15401];
assign g[31784] = b[13] & g[15401];
assign g[23594] = a[13] & g[15402];
assign g[31785] = b[13] & g[15402];
assign g[23595] = a[13] & g[15403];
assign g[31786] = b[13] & g[15403];
assign g[23596] = a[13] & g[15404];
assign g[31787] = b[13] & g[15404];
assign g[23597] = a[13] & g[15405];
assign g[31788] = b[13] & g[15405];
assign g[23598] = a[13] & g[15406];
assign g[31789] = b[13] & g[15406];
assign g[23599] = a[13] & g[15407];
assign g[31790] = b[13] & g[15407];
assign g[23600] = a[13] & g[15408];
assign g[31791] = b[13] & g[15408];
assign g[23601] = a[13] & g[15409];
assign g[31792] = b[13] & g[15409];
assign g[23602] = a[13] & g[15410];
assign g[31793] = b[13] & g[15410];
assign g[23603] = a[13] & g[15411];
assign g[31794] = b[13] & g[15411];
assign g[23604] = a[13] & g[15412];
assign g[31795] = b[13] & g[15412];
assign g[23605] = a[13] & g[15413];
assign g[31796] = b[13] & g[15413];
assign g[23606] = a[13] & g[15414];
assign g[31797] = b[13] & g[15414];
assign g[23607] = a[13] & g[15415];
assign g[31798] = b[13] & g[15415];
assign g[23608] = a[13] & g[15416];
assign g[31799] = b[13] & g[15416];
assign g[23609] = a[13] & g[15417];
assign g[31800] = b[13] & g[15417];
assign g[23610] = a[13] & g[15418];
assign g[31801] = b[13] & g[15418];
assign g[23611] = a[13] & g[15419];
assign g[31802] = b[13] & g[15419];
assign g[23612] = a[13] & g[15420];
assign g[31803] = b[13] & g[15420];
assign g[23613] = a[13] & g[15421];
assign g[31804] = b[13] & g[15421];
assign g[23614] = a[13] & g[15422];
assign g[31805] = b[13] & g[15422];
assign g[23615] = a[13] & g[15423];
assign g[31806] = b[13] & g[15423];
assign g[23616] = a[13] & g[15424];
assign g[31807] = b[13] & g[15424];
assign g[23617] = a[13] & g[15425];
assign g[31808] = b[13] & g[15425];
assign g[23618] = a[13] & g[15426];
assign g[31809] = b[13] & g[15426];
assign g[23619] = a[13] & g[15427];
assign g[31810] = b[13] & g[15427];
assign g[23620] = a[13] & g[15428];
assign g[31811] = b[13] & g[15428];
assign g[23621] = a[13] & g[15429];
assign g[31812] = b[13] & g[15429];
assign g[23622] = a[13] & g[15430];
assign g[31813] = b[13] & g[15430];
assign g[23623] = a[13] & g[15431];
assign g[31814] = b[13] & g[15431];
assign g[23624] = a[13] & g[15432];
assign g[31815] = b[13] & g[15432];
assign g[23625] = a[13] & g[15433];
assign g[31816] = b[13] & g[15433];
assign g[23626] = a[13] & g[15434];
assign g[31817] = b[13] & g[15434];
assign g[23627] = a[13] & g[15435];
assign g[31818] = b[13] & g[15435];
assign g[23628] = a[13] & g[15436];
assign g[31819] = b[13] & g[15436];
assign g[23629] = a[13] & g[15437];
assign g[31820] = b[13] & g[15437];
assign g[23630] = a[13] & g[15438];
assign g[31821] = b[13] & g[15438];
assign g[23631] = a[13] & g[15439];
assign g[31822] = b[13] & g[15439];
assign g[23632] = a[13] & g[15440];
assign g[31823] = b[13] & g[15440];
assign g[23633] = a[13] & g[15441];
assign g[31824] = b[13] & g[15441];
assign g[23634] = a[13] & g[15442];
assign g[31825] = b[13] & g[15442];
assign g[23635] = a[13] & g[15443];
assign g[31826] = b[13] & g[15443];
assign g[23636] = a[13] & g[15444];
assign g[31827] = b[13] & g[15444];
assign g[23637] = a[13] & g[15445];
assign g[31828] = b[13] & g[15445];
assign g[23638] = a[13] & g[15446];
assign g[31829] = b[13] & g[15446];
assign g[23639] = a[13] & g[15447];
assign g[31830] = b[13] & g[15447];
assign g[23640] = a[13] & g[15448];
assign g[31831] = b[13] & g[15448];
assign g[23641] = a[13] & g[15449];
assign g[31832] = b[13] & g[15449];
assign g[23642] = a[13] & g[15450];
assign g[31833] = b[13] & g[15450];
assign g[23643] = a[13] & g[15451];
assign g[31834] = b[13] & g[15451];
assign g[23644] = a[13] & g[15452];
assign g[31835] = b[13] & g[15452];
assign g[23645] = a[13] & g[15453];
assign g[31836] = b[13] & g[15453];
assign g[23646] = a[13] & g[15454];
assign g[31837] = b[13] & g[15454];
assign g[23647] = a[13] & g[15455];
assign g[31838] = b[13] & g[15455];
assign g[23648] = a[13] & g[15456];
assign g[31839] = b[13] & g[15456];
assign g[23649] = a[13] & g[15457];
assign g[31840] = b[13] & g[15457];
assign g[23650] = a[13] & g[15458];
assign g[31841] = b[13] & g[15458];
assign g[23651] = a[13] & g[15459];
assign g[31842] = b[13] & g[15459];
assign g[23652] = a[13] & g[15460];
assign g[31843] = b[13] & g[15460];
assign g[23653] = a[13] & g[15461];
assign g[31844] = b[13] & g[15461];
assign g[23654] = a[13] & g[15462];
assign g[31845] = b[13] & g[15462];
assign g[23655] = a[13] & g[15463];
assign g[31846] = b[13] & g[15463];
assign g[23656] = a[13] & g[15464];
assign g[31847] = b[13] & g[15464];
assign g[23657] = a[13] & g[15465];
assign g[31848] = b[13] & g[15465];
assign g[23658] = a[13] & g[15466];
assign g[31849] = b[13] & g[15466];
assign g[23659] = a[13] & g[15467];
assign g[31850] = b[13] & g[15467];
assign g[23660] = a[13] & g[15468];
assign g[31851] = b[13] & g[15468];
assign g[23661] = a[13] & g[15469];
assign g[31852] = b[13] & g[15469];
assign g[23662] = a[13] & g[15470];
assign g[31853] = b[13] & g[15470];
assign g[23663] = a[13] & g[15471];
assign g[31854] = b[13] & g[15471];
assign g[23664] = a[13] & g[15472];
assign g[31855] = b[13] & g[15472];
assign g[23665] = a[13] & g[15473];
assign g[31856] = b[13] & g[15473];
assign g[23666] = a[13] & g[15474];
assign g[31857] = b[13] & g[15474];
assign g[23667] = a[13] & g[15475];
assign g[31858] = b[13] & g[15475];
assign g[23668] = a[13] & g[15476];
assign g[31859] = b[13] & g[15476];
assign g[23669] = a[13] & g[15477];
assign g[31860] = b[13] & g[15477];
assign g[23670] = a[13] & g[15478];
assign g[31861] = b[13] & g[15478];
assign g[23671] = a[13] & g[15479];
assign g[31862] = b[13] & g[15479];
assign g[23672] = a[13] & g[15480];
assign g[31863] = b[13] & g[15480];
assign g[23673] = a[13] & g[15481];
assign g[31864] = b[13] & g[15481];
assign g[23674] = a[13] & g[15482];
assign g[31865] = b[13] & g[15482];
assign g[23675] = a[13] & g[15483];
assign g[31866] = b[13] & g[15483];
assign g[23676] = a[13] & g[15484];
assign g[31867] = b[13] & g[15484];
assign g[23677] = a[13] & g[15485];
assign g[31868] = b[13] & g[15485];
assign g[23678] = a[13] & g[15486];
assign g[31869] = b[13] & g[15486];
assign g[23679] = a[13] & g[15487];
assign g[31870] = b[13] & g[15487];
assign g[23680] = a[13] & g[15488];
assign g[31871] = b[13] & g[15488];
assign g[23681] = a[13] & g[15489];
assign g[31872] = b[13] & g[15489];
assign g[23682] = a[13] & g[15490];
assign g[31873] = b[13] & g[15490];
assign g[23683] = a[13] & g[15491];
assign g[31874] = b[13] & g[15491];
assign g[23684] = a[13] & g[15492];
assign g[31875] = b[13] & g[15492];
assign g[23685] = a[13] & g[15493];
assign g[31876] = b[13] & g[15493];
assign g[23686] = a[13] & g[15494];
assign g[31877] = b[13] & g[15494];
assign g[23687] = a[13] & g[15495];
assign g[31878] = b[13] & g[15495];
assign g[23688] = a[13] & g[15496];
assign g[31879] = b[13] & g[15496];
assign g[23689] = a[13] & g[15497];
assign g[31880] = b[13] & g[15497];
assign g[23690] = a[13] & g[15498];
assign g[31881] = b[13] & g[15498];
assign g[23691] = a[13] & g[15499];
assign g[31882] = b[13] & g[15499];
assign g[23692] = a[13] & g[15500];
assign g[31883] = b[13] & g[15500];
assign g[23693] = a[13] & g[15501];
assign g[31884] = b[13] & g[15501];
assign g[23694] = a[13] & g[15502];
assign g[31885] = b[13] & g[15502];
assign g[23695] = a[13] & g[15503];
assign g[31886] = b[13] & g[15503];
assign g[23696] = a[13] & g[15504];
assign g[31887] = b[13] & g[15504];
assign g[23697] = a[13] & g[15505];
assign g[31888] = b[13] & g[15505];
assign g[23698] = a[13] & g[15506];
assign g[31889] = b[13] & g[15506];
assign g[23699] = a[13] & g[15507];
assign g[31890] = b[13] & g[15507];
assign g[23700] = a[13] & g[15508];
assign g[31891] = b[13] & g[15508];
assign g[23701] = a[13] & g[15509];
assign g[31892] = b[13] & g[15509];
assign g[23702] = a[13] & g[15510];
assign g[31893] = b[13] & g[15510];
assign g[23703] = a[13] & g[15511];
assign g[31894] = b[13] & g[15511];
assign g[23704] = a[13] & g[15512];
assign g[31895] = b[13] & g[15512];
assign g[23705] = a[13] & g[15513];
assign g[31896] = b[13] & g[15513];
assign g[23706] = a[13] & g[15514];
assign g[31897] = b[13] & g[15514];
assign g[23707] = a[13] & g[15515];
assign g[31898] = b[13] & g[15515];
assign g[23708] = a[13] & g[15516];
assign g[31899] = b[13] & g[15516];
assign g[23709] = a[13] & g[15517];
assign g[31900] = b[13] & g[15517];
assign g[23710] = a[13] & g[15518];
assign g[31901] = b[13] & g[15518];
assign g[23711] = a[13] & g[15519];
assign g[31902] = b[13] & g[15519];
assign g[23712] = a[13] & g[15520];
assign g[31903] = b[13] & g[15520];
assign g[23713] = a[13] & g[15521];
assign g[31904] = b[13] & g[15521];
assign g[23714] = a[13] & g[15522];
assign g[31905] = b[13] & g[15522];
assign g[23715] = a[13] & g[15523];
assign g[31906] = b[13] & g[15523];
assign g[23716] = a[13] & g[15524];
assign g[31907] = b[13] & g[15524];
assign g[23717] = a[13] & g[15525];
assign g[31908] = b[13] & g[15525];
assign g[23718] = a[13] & g[15526];
assign g[31909] = b[13] & g[15526];
assign g[23719] = a[13] & g[15527];
assign g[31910] = b[13] & g[15527];
assign g[23720] = a[13] & g[15528];
assign g[31911] = b[13] & g[15528];
assign g[23721] = a[13] & g[15529];
assign g[31912] = b[13] & g[15529];
assign g[23722] = a[13] & g[15530];
assign g[31913] = b[13] & g[15530];
assign g[23723] = a[13] & g[15531];
assign g[31914] = b[13] & g[15531];
assign g[23724] = a[13] & g[15532];
assign g[31915] = b[13] & g[15532];
assign g[23725] = a[13] & g[15533];
assign g[31916] = b[13] & g[15533];
assign g[23726] = a[13] & g[15534];
assign g[31917] = b[13] & g[15534];
assign g[23727] = a[13] & g[15535];
assign g[31918] = b[13] & g[15535];
assign g[23728] = a[13] & g[15536];
assign g[31919] = b[13] & g[15536];
assign g[23729] = a[13] & g[15537];
assign g[31920] = b[13] & g[15537];
assign g[23730] = a[13] & g[15538];
assign g[31921] = b[13] & g[15538];
assign g[23731] = a[13] & g[15539];
assign g[31922] = b[13] & g[15539];
assign g[23732] = a[13] & g[15540];
assign g[31923] = b[13] & g[15540];
assign g[23733] = a[13] & g[15541];
assign g[31924] = b[13] & g[15541];
assign g[23734] = a[13] & g[15542];
assign g[31925] = b[13] & g[15542];
assign g[23735] = a[13] & g[15543];
assign g[31926] = b[13] & g[15543];
assign g[23736] = a[13] & g[15544];
assign g[31927] = b[13] & g[15544];
assign g[23737] = a[13] & g[15545];
assign g[31928] = b[13] & g[15545];
assign g[23738] = a[13] & g[15546];
assign g[31929] = b[13] & g[15546];
assign g[23739] = a[13] & g[15547];
assign g[31930] = b[13] & g[15547];
assign g[23740] = a[13] & g[15548];
assign g[31931] = b[13] & g[15548];
assign g[23741] = a[13] & g[15549];
assign g[31932] = b[13] & g[15549];
assign g[23742] = a[13] & g[15550];
assign g[31933] = b[13] & g[15550];
assign g[23743] = a[13] & g[15551];
assign g[31934] = b[13] & g[15551];
assign g[23744] = a[13] & g[15552];
assign g[31935] = b[13] & g[15552];
assign g[23745] = a[13] & g[15553];
assign g[31936] = b[13] & g[15553];
assign g[23746] = a[13] & g[15554];
assign g[31937] = b[13] & g[15554];
assign g[23747] = a[13] & g[15555];
assign g[31938] = b[13] & g[15555];
assign g[23748] = a[13] & g[15556];
assign g[31939] = b[13] & g[15556];
assign g[23749] = a[13] & g[15557];
assign g[31940] = b[13] & g[15557];
assign g[23750] = a[13] & g[15558];
assign g[31941] = b[13] & g[15558];
assign g[23751] = a[13] & g[15559];
assign g[31942] = b[13] & g[15559];
assign g[23752] = a[13] & g[15560];
assign g[31943] = b[13] & g[15560];
assign g[23753] = a[13] & g[15561];
assign g[31944] = b[13] & g[15561];
assign g[23754] = a[13] & g[15562];
assign g[31945] = b[13] & g[15562];
assign g[23755] = a[13] & g[15563];
assign g[31946] = b[13] & g[15563];
assign g[23756] = a[13] & g[15564];
assign g[31947] = b[13] & g[15564];
assign g[23757] = a[13] & g[15565];
assign g[31948] = b[13] & g[15565];
assign g[23758] = a[13] & g[15566];
assign g[31949] = b[13] & g[15566];
assign g[23759] = a[13] & g[15567];
assign g[31950] = b[13] & g[15567];
assign g[23760] = a[13] & g[15568];
assign g[31951] = b[13] & g[15568];
assign g[23761] = a[13] & g[15569];
assign g[31952] = b[13] & g[15569];
assign g[23762] = a[13] & g[15570];
assign g[31953] = b[13] & g[15570];
assign g[23763] = a[13] & g[15571];
assign g[31954] = b[13] & g[15571];
assign g[23764] = a[13] & g[15572];
assign g[31955] = b[13] & g[15572];
assign g[23765] = a[13] & g[15573];
assign g[31956] = b[13] & g[15573];
assign g[23766] = a[13] & g[15574];
assign g[31957] = b[13] & g[15574];
assign g[23767] = a[13] & g[15575];
assign g[31958] = b[13] & g[15575];
assign g[23768] = a[13] & g[15576];
assign g[31959] = b[13] & g[15576];
assign g[23769] = a[13] & g[15577];
assign g[31960] = b[13] & g[15577];
assign g[23770] = a[13] & g[15578];
assign g[31961] = b[13] & g[15578];
assign g[23771] = a[13] & g[15579];
assign g[31962] = b[13] & g[15579];
assign g[23772] = a[13] & g[15580];
assign g[31963] = b[13] & g[15580];
assign g[23773] = a[13] & g[15581];
assign g[31964] = b[13] & g[15581];
assign g[23774] = a[13] & g[15582];
assign g[31965] = b[13] & g[15582];
assign g[23775] = a[13] & g[15583];
assign g[31966] = b[13] & g[15583];
assign g[23776] = a[13] & g[15584];
assign g[31967] = b[13] & g[15584];
assign g[23777] = a[13] & g[15585];
assign g[31968] = b[13] & g[15585];
assign g[23778] = a[13] & g[15586];
assign g[31969] = b[13] & g[15586];
assign g[23779] = a[13] & g[15587];
assign g[31970] = b[13] & g[15587];
assign g[23780] = a[13] & g[15588];
assign g[31971] = b[13] & g[15588];
assign g[23781] = a[13] & g[15589];
assign g[31972] = b[13] & g[15589];
assign g[23782] = a[13] & g[15590];
assign g[31973] = b[13] & g[15590];
assign g[23783] = a[13] & g[15591];
assign g[31974] = b[13] & g[15591];
assign g[23784] = a[13] & g[15592];
assign g[31975] = b[13] & g[15592];
assign g[23785] = a[13] & g[15593];
assign g[31976] = b[13] & g[15593];
assign g[23786] = a[13] & g[15594];
assign g[31977] = b[13] & g[15594];
assign g[23787] = a[13] & g[15595];
assign g[31978] = b[13] & g[15595];
assign g[23788] = a[13] & g[15596];
assign g[31979] = b[13] & g[15596];
assign g[23789] = a[13] & g[15597];
assign g[31980] = b[13] & g[15597];
assign g[23790] = a[13] & g[15598];
assign g[31981] = b[13] & g[15598];
assign g[23791] = a[13] & g[15599];
assign g[31982] = b[13] & g[15599];
assign g[23792] = a[13] & g[15600];
assign g[31983] = b[13] & g[15600];
assign g[23793] = a[13] & g[15601];
assign g[31984] = b[13] & g[15601];
assign g[23794] = a[13] & g[15602];
assign g[31985] = b[13] & g[15602];
assign g[23795] = a[13] & g[15603];
assign g[31986] = b[13] & g[15603];
assign g[23796] = a[13] & g[15604];
assign g[31987] = b[13] & g[15604];
assign g[23797] = a[13] & g[15605];
assign g[31988] = b[13] & g[15605];
assign g[23798] = a[13] & g[15606];
assign g[31989] = b[13] & g[15606];
assign g[23799] = a[13] & g[15607];
assign g[31990] = b[13] & g[15607];
assign g[23800] = a[13] & g[15608];
assign g[31991] = b[13] & g[15608];
assign g[23801] = a[13] & g[15609];
assign g[31992] = b[13] & g[15609];
assign g[23802] = a[13] & g[15610];
assign g[31993] = b[13] & g[15610];
assign g[23803] = a[13] & g[15611];
assign g[31994] = b[13] & g[15611];
assign g[23804] = a[13] & g[15612];
assign g[31995] = b[13] & g[15612];
assign g[23805] = a[13] & g[15613];
assign g[31996] = b[13] & g[15613];
assign g[23806] = a[13] & g[15614];
assign g[31997] = b[13] & g[15614];
assign g[23807] = a[13] & g[15615];
assign g[31998] = b[13] & g[15615];
assign g[23808] = a[13] & g[15616];
assign g[31999] = b[13] & g[15616];
assign g[23809] = a[13] & g[15617];
assign g[32000] = b[13] & g[15617];
assign g[23810] = a[13] & g[15618];
assign g[32001] = b[13] & g[15618];
assign g[23811] = a[13] & g[15619];
assign g[32002] = b[13] & g[15619];
assign g[23812] = a[13] & g[15620];
assign g[32003] = b[13] & g[15620];
assign g[23813] = a[13] & g[15621];
assign g[32004] = b[13] & g[15621];
assign g[23814] = a[13] & g[15622];
assign g[32005] = b[13] & g[15622];
assign g[23815] = a[13] & g[15623];
assign g[32006] = b[13] & g[15623];
assign g[23816] = a[13] & g[15624];
assign g[32007] = b[13] & g[15624];
assign g[23817] = a[13] & g[15625];
assign g[32008] = b[13] & g[15625];
assign g[23818] = a[13] & g[15626];
assign g[32009] = b[13] & g[15626];
assign g[23819] = a[13] & g[15627];
assign g[32010] = b[13] & g[15627];
assign g[23820] = a[13] & g[15628];
assign g[32011] = b[13] & g[15628];
assign g[23821] = a[13] & g[15629];
assign g[32012] = b[13] & g[15629];
assign g[23822] = a[13] & g[15630];
assign g[32013] = b[13] & g[15630];
assign g[23823] = a[13] & g[15631];
assign g[32014] = b[13] & g[15631];
assign g[23824] = a[13] & g[15632];
assign g[32015] = b[13] & g[15632];
assign g[23825] = a[13] & g[15633];
assign g[32016] = b[13] & g[15633];
assign g[23826] = a[13] & g[15634];
assign g[32017] = b[13] & g[15634];
assign g[23827] = a[13] & g[15635];
assign g[32018] = b[13] & g[15635];
assign g[23828] = a[13] & g[15636];
assign g[32019] = b[13] & g[15636];
assign g[23829] = a[13] & g[15637];
assign g[32020] = b[13] & g[15637];
assign g[23830] = a[13] & g[15638];
assign g[32021] = b[13] & g[15638];
assign g[23831] = a[13] & g[15639];
assign g[32022] = b[13] & g[15639];
assign g[23832] = a[13] & g[15640];
assign g[32023] = b[13] & g[15640];
assign g[23833] = a[13] & g[15641];
assign g[32024] = b[13] & g[15641];
assign g[23834] = a[13] & g[15642];
assign g[32025] = b[13] & g[15642];
assign g[23835] = a[13] & g[15643];
assign g[32026] = b[13] & g[15643];
assign g[23836] = a[13] & g[15644];
assign g[32027] = b[13] & g[15644];
assign g[23837] = a[13] & g[15645];
assign g[32028] = b[13] & g[15645];
assign g[23838] = a[13] & g[15646];
assign g[32029] = b[13] & g[15646];
assign g[23839] = a[13] & g[15647];
assign g[32030] = b[13] & g[15647];
assign g[23840] = a[13] & g[15648];
assign g[32031] = b[13] & g[15648];
assign g[23841] = a[13] & g[15649];
assign g[32032] = b[13] & g[15649];
assign g[23842] = a[13] & g[15650];
assign g[32033] = b[13] & g[15650];
assign g[23843] = a[13] & g[15651];
assign g[32034] = b[13] & g[15651];
assign g[23844] = a[13] & g[15652];
assign g[32035] = b[13] & g[15652];
assign g[23845] = a[13] & g[15653];
assign g[32036] = b[13] & g[15653];
assign g[23846] = a[13] & g[15654];
assign g[32037] = b[13] & g[15654];
assign g[23847] = a[13] & g[15655];
assign g[32038] = b[13] & g[15655];
assign g[23848] = a[13] & g[15656];
assign g[32039] = b[13] & g[15656];
assign g[23849] = a[13] & g[15657];
assign g[32040] = b[13] & g[15657];
assign g[23850] = a[13] & g[15658];
assign g[32041] = b[13] & g[15658];
assign g[23851] = a[13] & g[15659];
assign g[32042] = b[13] & g[15659];
assign g[23852] = a[13] & g[15660];
assign g[32043] = b[13] & g[15660];
assign g[23853] = a[13] & g[15661];
assign g[32044] = b[13] & g[15661];
assign g[23854] = a[13] & g[15662];
assign g[32045] = b[13] & g[15662];
assign g[23855] = a[13] & g[15663];
assign g[32046] = b[13] & g[15663];
assign g[23856] = a[13] & g[15664];
assign g[32047] = b[13] & g[15664];
assign g[23857] = a[13] & g[15665];
assign g[32048] = b[13] & g[15665];
assign g[23858] = a[13] & g[15666];
assign g[32049] = b[13] & g[15666];
assign g[23859] = a[13] & g[15667];
assign g[32050] = b[13] & g[15667];
assign g[23860] = a[13] & g[15668];
assign g[32051] = b[13] & g[15668];
assign g[23861] = a[13] & g[15669];
assign g[32052] = b[13] & g[15669];
assign g[23862] = a[13] & g[15670];
assign g[32053] = b[13] & g[15670];
assign g[23863] = a[13] & g[15671];
assign g[32054] = b[13] & g[15671];
assign g[23864] = a[13] & g[15672];
assign g[32055] = b[13] & g[15672];
assign g[23865] = a[13] & g[15673];
assign g[32056] = b[13] & g[15673];
assign g[23866] = a[13] & g[15674];
assign g[32057] = b[13] & g[15674];
assign g[23867] = a[13] & g[15675];
assign g[32058] = b[13] & g[15675];
assign g[23868] = a[13] & g[15676];
assign g[32059] = b[13] & g[15676];
assign g[23869] = a[13] & g[15677];
assign g[32060] = b[13] & g[15677];
assign g[23870] = a[13] & g[15678];
assign g[32061] = b[13] & g[15678];
assign g[23871] = a[13] & g[15679];
assign g[32062] = b[13] & g[15679];
assign g[23872] = a[13] & g[15680];
assign g[32063] = b[13] & g[15680];
assign g[23873] = a[13] & g[15681];
assign g[32064] = b[13] & g[15681];
assign g[23874] = a[13] & g[15682];
assign g[32065] = b[13] & g[15682];
assign g[23875] = a[13] & g[15683];
assign g[32066] = b[13] & g[15683];
assign g[23876] = a[13] & g[15684];
assign g[32067] = b[13] & g[15684];
assign g[23877] = a[13] & g[15685];
assign g[32068] = b[13] & g[15685];
assign g[23878] = a[13] & g[15686];
assign g[32069] = b[13] & g[15686];
assign g[23879] = a[13] & g[15687];
assign g[32070] = b[13] & g[15687];
assign g[23880] = a[13] & g[15688];
assign g[32071] = b[13] & g[15688];
assign g[23881] = a[13] & g[15689];
assign g[32072] = b[13] & g[15689];
assign g[23882] = a[13] & g[15690];
assign g[32073] = b[13] & g[15690];
assign g[23883] = a[13] & g[15691];
assign g[32074] = b[13] & g[15691];
assign g[23884] = a[13] & g[15692];
assign g[32075] = b[13] & g[15692];
assign g[23885] = a[13] & g[15693];
assign g[32076] = b[13] & g[15693];
assign g[23886] = a[13] & g[15694];
assign g[32077] = b[13] & g[15694];
assign g[23887] = a[13] & g[15695];
assign g[32078] = b[13] & g[15695];
assign g[23888] = a[13] & g[15696];
assign g[32079] = b[13] & g[15696];
assign g[23889] = a[13] & g[15697];
assign g[32080] = b[13] & g[15697];
assign g[23890] = a[13] & g[15698];
assign g[32081] = b[13] & g[15698];
assign g[23891] = a[13] & g[15699];
assign g[32082] = b[13] & g[15699];
assign g[23892] = a[13] & g[15700];
assign g[32083] = b[13] & g[15700];
assign g[23893] = a[13] & g[15701];
assign g[32084] = b[13] & g[15701];
assign g[23894] = a[13] & g[15702];
assign g[32085] = b[13] & g[15702];
assign g[23895] = a[13] & g[15703];
assign g[32086] = b[13] & g[15703];
assign g[23896] = a[13] & g[15704];
assign g[32087] = b[13] & g[15704];
assign g[23897] = a[13] & g[15705];
assign g[32088] = b[13] & g[15705];
assign g[23898] = a[13] & g[15706];
assign g[32089] = b[13] & g[15706];
assign g[23899] = a[13] & g[15707];
assign g[32090] = b[13] & g[15707];
assign g[23900] = a[13] & g[15708];
assign g[32091] = b[13] & g[15708];
assign g[23901] = a[13] & g[15709];
assign g[32092] = b[13] & g[15709];
assign g[23902] = a[13] & g[15710];
assign g[32093] = b[13] & g[15710];
assign g[23903] = a[13] & g[15711];
assign g[32094] = b[13] & g[15711];
assign g[23904] = a[13] & g[15712];
assign g[32095] = b[13] & g[15712];
assign g[23905] = a[13] & g[15713];
assign g[32096] = b[13] & g[15713];
assign g[23906] = a[13] & g[15714];
assign g[32097] = b[13] & g[15714];
assign g[23907] = a[13] & g[15715];
assign g[32098] = b[13] & g[15715];
assign g[23908] = a[13] & g[15716];
assign g[32099] = b[13] & g[15716];
assign g[23909] = a[13] & g[15717];
assign g[32100] = b[13] & g[15717];
assign g[23910] = a[13] & g[15718];
assign g[32101] = b[13] & g[15718];
assign g[23911] = a[13] & g[15719];
assign g[32102] = b[13] & g[15719];
assign g[23912] = a[13] & g[15720];
assign g[32103] = b[13] & g[15720];
assign g[23913] = a[13] & g[15721];
assign g[32104] = b[13] & g[15721];
assign g[23914] = a[13] & g[15722];
assign g[32105] = b[13] & g[15722];
assign g[23915] = a[13] & g[15723];
assign g[32106] = b[13] & g[15723];
assign g[23916] = a[13] & g[15724];
assign g[32107] = b[13] & g[15724];
assign g[23917] = a[13] & g[15725];
assign g[32108] = b[13] & g[15725];
assign g[23918] = a[13] & g[15726];
assign g[32109] = b[13] & g[15726];
assign g[23919] = a[13] & g[15727];
assign g[32110] = b[13] & g[15727];
assign g[23920] = a[13] & g[15728];
assign g[32111] = b[13] & g[15728];
assign g[23921] = a[13] & g[15729];
assign g[32112] = b[13] & g[15729];
assign g[23922] = a[13] & g[15730];
assign g[32113] = b[13] & g[15730];
assign g[23923] = a[13] & g[15731];
assign g[32114] = b[13] & g[15731];
assign g[23924] = a[13] & g[15732];
assign g[32115] = b[13] & g[15732];
assign g[23925] = a[13] & g[15733];
assign g[32116] = b[13] & g[15733];
assign g[23926] = a[13] & g[15734];
assign g[32117] = b[13] & g[15734];
assign g[23927] = a[13] & g[15735];
assign g[32118] = b[13] & g[15735];
assign g[23928] = a[13] & g[15736];
assign g[32119] = b[13] & g[15736];
assign g[23929] = a[13] & g[15737];
assign g[32120] = b[13] & g[15737];
assign g[23930] = a[13] & g[15738];
assign g[32121] = b[13] & g[15738];
assign g[23931] = a[13] & g[15739];
assign g[32122] = b[13] & g[15739];
assign g[23932] = a[13] & g[15740];
assign g[32123] = b[13] & g[15740];
assign g[23933] = a[13] & g[15741];
assign g[32124] = b[13] & g[15741];
assign g[23934] = a[13] & g[15742];
assign g[32125] = b[13] & g[15742];
assign g[23935] = a[13] & g[15743];
assign g[32126] = b[13] & g[15743];
assign g[23936] = a[13] & g[15744];
assign g[32127] = b[13] & g[15744];
assign g[23937] = a[13] & g[15745];
assign g[32128] = b[13] & g[15745];
assign g[23938] = a[13] & g[15746];
assign g[32129] = b[13] & g[15746];
assign g[23939] = a[13] & g[15747];
assign g[32130] = b[13] & g[15747];
assign g[23940] = a[13] & g[15748];
assign g[32131] = b[13] & g[15748];
assign g[23941] = a[13] & g[15749];
assign g[32132] = b[13] & g[15749];
assign g[23942] = a[13] & g[15750];
assign g[32133] = b[13] & g[15750];
assign g[23943] = a[13] & g[15751];
assign g[32134] = b[13] & g[15751];
assign g[23944] = a[13] & g[15752];
assign g[32135] = b[13] & g[15752];
assign g[23945] = a[13] & g[15753];
assign g[32136] = b[13] & g[15753];
assign g[23946] = a[13] & g[15754];
assign g[32137] = b[13] & g[15754];
assign g[23947] = a[13] & g[15755];
assign g[32138] = b[13] & g[15755];
assign g[23948] = a[13] & g[15756];
assign g[32139] = b[13] & g[15756];
assign g[23949] = a[13] & g[15757];
assign g[32140] = b[13] & g[15757];
assign g[23950] = a[13] & g[15758];
assign g[32141] = b[13] & g[15758];
assign g[23951] = a[13] & g[15759];
assign g[32142] = b[13] & g[15759];
assign g[23952] = a[13] & g[15760];
assign g[32143] = b[13] & g[15760];
assign g[23953] = a[13] & g[15761];
assign g[32144] = b[13] & g[15761];
assign g[23954] = a[13] & g[15762];
assign g[32145] = b[13] & g[15762];
assign g[23955] = a[13] & g[15763];
assign g[32146] = b[13] & g[15763];
assign g[23956] = a[13] & g[15764];
assign g[32147] = b[13] & g[15764];
assign g[23957] = a[13] & g[15765];
assign g[32148] = b[13] & g[15765];
assign g[23958] = a[13] & g[15766];
assign g[32149] = b[13] & g[15766];
assign g[23959] = a[13] & g[15767];
assign g[32150] = b[13] & g[15767];
assign g[23960] = a[13] & g[15768];
assign g[32151] = b[13] & g[15768];
assign g[23961] = a[13] & g[15769];
assign g[32152] = b[13] & g[15769];
assign g[23962] = a[13] & g[15770];
assign g[32153] = b[13] & g[15770];
assign g[23963] = a[13] & g[15771];
assign g[32154] = b[13] & g[15771];
assign g[23964] = a[13] & g[15772];
assign g[32155] = b[13] & g[15772];
assign g[23965] = a[13] & g[15773];
assign g[32156] = b[13] & g[15773];
assign g[23966] = a[13] & g[15774];
assign g[32157] = b[13] & g[15774];
assign g[23967] = a[13] & g[15775];
assign g[32158] = b[13] & g[15775];
assign g[23968] = a[13] & g[15776];
assign g[32159] = b[13] & g[15776];
assign g[23969] = a[13] & g[15777];
assign g[32160] = b[13] & g[15777];
assign g[23970] = a[13] & g[15778];
assign g[32161] = b[13] & g[15778];
assign g[23971] = a[13] & g[15779];
assign g[32162] = b[13] & g[15779];
assign g[23972] = a[13] & g[15780];
assign g[32163] = b[13] & g[15780];
assign g[23973] = a[13] & g[15781];
assign g[32164] = b[13] & g[15781];
assign g[23974] = a[13] & g[15782];
assign g[32165] = b[13] & g[15782];
assign g[23975] = a[13] & g[15783];
assign g[32166] = b[13] & g[15783];
assign g[23976] = a[13] & g[15784];
assign g[32167] = b[13] & g[15784];
assign g[23977] = a[13] & g[15785];
assign g[32168] = b[13] & g[15785];
assign g[23978] = a[13] & g[15786];
assign g[32169] = b[13] & g[15786];
assign g[23979] = a[13] & g[15787];
assign g[32170] = b[13] & g[15787];
assign g[23980] = a[13] & g[15788];
assign g[32171] = b[13] & g[15788];
assign g[23981] = a[13] & g[15789];
assign g[32172] = b[13] & g[15789];
assign g[23982] = a[13] & g[15790];
assign g[32173] = b[13] & g[15790];
assign g[23983] = a[13] & g[15791];
assign g[32174] = b[13] & g[15791];
assign g[23984] = a[13] & g[15792];
assign g[32175] = b[13] & g[15792];
assign g[23985] = a[13] & g[15793];
assign g[32176] = b[13] & g[15793];
assign g[23986] = a[13] & g[15794];
assign g[32177] = b[13] & g[15794];
assign g[23987] = a[13] & g[15795];
assign g[32178] = b[13] & g[15795];
assign g[23988] = a[13] & g[15796];
assign g[32179] = b[13] & g[15796];
assign g[23989] = a[13] & g[15797];
assign g[32180] = b[13] & g[15797];
assign g[23990] = a[13] & g[15798];
assign g[32181] = b[13] & g[15798];
assign g[23991] = a[13] & g[15799];
assign g[32182] = b[13] & g[15799];
assign g[23992] = a[13] & g[15800];
assign g[32183] = b[13] & g[15800];
assign g[23993] = a[13] & g[15801];
assign g[32184] = b[13] & g[15801];
assign g[23994] = a[13] & g[15802];
assign g[32185] = b[13] & g[15802];
assign g[23995] = a[13] & g[15803];
assign g[32186] = b[13] & g[15803];
assign g[23996] = a[13] & g[15804];
assign g[32187] = b[13] & g[15804];
assign g[23997] = a[13] & g[15805];
assign g[32188] = b[13] & g[15805];
assign g[23998] = a[13] & g[15806];
assign g[32189] = b[13] & g[15806];
assign g[23999] = a[13] & g[15807];
assign g[32190] = b[13] & g[15807];
assign g[24000] = a[13] & g[15808];
assign g[32191] = b[13] & g[15808];
assign g[24001] = a[13] & g[15809];
assign g[32192] = b[13] & g[15809];
assign g[24002] = a[13] & g[15810];
assign g[32193] = b[13] & g[15810];
assign g[24003] = a[13] & g[15811];
assign g[32194] = b[13] & g[15811];
assign g[24004] = a[13] & g[15812];
assign g[32195] = b[13] & g[15812];
assign g[24005] = a[13] & g[15813];
assign g[32196] = b[13] & g[15813];
assign g[24006] = a[13] & g[15814];
assign g[32197] = b[13] & g[15814];
assign g[24007] = a[13] & g[15815];
assign g[32198] = b[13] & g[15815];
assign g[24008] = a[13] & g[15816];
assign g[32199] = b[13] & g[15816];
assign g[24009] = a[13] & g[15817];
assign g[32200] = b[13] & g[15817];
assign g[24010] = a[13] & g[15818];
assign g[32201] = b[13] & g[15818];
assign g[24011] = a[13] & g[15819];
assign g[32202] = b[13] & g[15819];
assign g[24012] = a[13] & g[15820];
assign g[32203] = b[13] & g[15820];
assign g[24013] = a[13] & g[15821];
assign g[32204] = b[13] & g[15821];
assign g[24014] = a[13] & g[15822];
assign g[32205] = b[13] & g[15822];
assign g[24015] = a[13] & g[15823];
assign g[32206] = b[13] & g[15823];
assign g[24016] = a[13] & g[15824];
assign g[32207] = b[13] & g[15824];
assign g[24017] = a[13] & g[15825];
assign g[32208] = b[13] & g[15825];
assign g[24018] = a[13] & g[15826];
assign g[32209] = b[13] & g[15826];
assign g[24019] = a[13] & g[15827];
assign g[32210] = b[13] & g[15827];
assign g[24020] = a[13] & g[15828];
assign g[32211] = b[13] & g[15828];
assign g[24021] = a[13] & g[15829];
assign g[32212] = b[13] & g[15829];
assign g[24022] = a[13] & g[15830];
assign g[32213] = b[13] & g[15830];
assign g[24023] = a[13] & g[15831];
assign g[32214] = b[13] & g[15831];
assign g[24024] = a[13] & g[15832];
assign g[32215] = b[13] & g[15832];
assign g[24025] = a[13] & g[15833];
assign g[32216] = b[13] & g[15833];
assign g[24026] = a[13] & g[15834];
assign g[32217] = b[13] & g[15834];
assign g[24027] = a[13] & g[15835];
assign g[32218] = b[13] & g[15835];
assign g[24028] = a[13] & g[15836];
assign g[32219] = b[13] & g[15836];
assign g[24029] = a[13] & g[15837];
assign g[32220] = b[13] & g[15837];
assign g[24030] = a[13] & g[15838];
assign g[32221] = b[13] & g[15838];
assign g[24031] = a[13] & g[15839];
assign g[32222] = b[13] & g[15839];
assign g[24032] = a[13] & g[15840];
assign g[32223] = b[13] & g[15840];
assign g[24033] = a[13] & g[15841];
assign g[32224] = b[13] & g[15841];
assign g[24034] = a[13] & g[15842];
assign g[32225] = b[13] & g[15842];
assign g[24035] = a[13] & g[15843];
assign g[32226] = b[13] & g[15843];
assign g[24036] = a[13] & g[15844];
assign g[32227] = b[13] & g[15844];
assign g[24037] = a[13] & g[15845];
assign g[32228] = b[13] & g[15845];
assign g[24038] = a[13] & g[15846];
assign g[32229] = b[13] & g[15846];
assign g[24039] = a[13] & g[15847];
assign g[32230] = b[13] & g[15847];
assign g[24040] = a[13] & g[15848];
assign g[32231] = b[13] & g[15848];
assign g[24041] = a[13] & g[15849];
assign g[32232] = b[13] & g[15849];
assign g[24042] = a[13] & g[15850];
assign g[32233] = b[13] & g[15850];
assign g[24043] = a[13] & g[15851];
assign g[32234] = b[13] & g[15851];
assign g[24044] = a[13] & g[15852];
assign g[32235] = b[13] & g[15852];
assign g[24045] = a[13] & g[15853];
assign g[32236] = b[13] & g[15853];
assign g[24046] = a[13] & g[15854];
assign g[32237] = b[13] & g[15854];
assign g[24047] = a[13] & g[15855];
assign g[32238] = b[13] & g[15855];
assign g[24048] = a[13] & g[15856];
assign g[32239] = b[13] & g[15856];
assign g[24049] = a[13] & g[15857];
assign g[32240] = b[13] & g[15857];
assign g[24050] = a[13] & g[15858];
assign g[32241] = b[13] & g[15858];
assign g[24051] = a[13] & g[15859];
assign g[32242] = b[13] & g[15859];
assign g[24052] = a[13] & g[15860];
assign g[32243] = b[13] & g[15860];
assign g[24053] = a[13] & g[15861];
assign g[32244] = b[13] & g[15861];
assign g[24054] = a[13] & g[15862];
assign g[32245] = b[13] & g[15862];
assign g[24055] = a[13] & g[15863];
assign g[32246] = b[13] & g[15863];
assign g[24056] = a[13] & g[15864];
assign g[32247] = b[13] & g[15864];
assign g[24057] = a[13] & g[15865];
assign g[32248] = b[13] & g[15865];
assign g[24058] = a[13] & g[15866];
assign g[32249] = b[13] & g[15866];
assign g[24059] = a[13] & g[15867];
assign g[32250] = b[13] & g[15867];
assign g[24060] = a[13] & g[15868];
assign g[32251] = b[13] & g[15868];
assign g[24061] = a[13] & g[15869];
assign g[32252] = b[13] & g[15869];
assign g[24062] = a[13] & g[15870];
assign g[32253] = b[13] & g[15870];
assign g[24063] = a[13] & g[15871];
assign g[32254] = b[13] & g[15871];
assign g[24064] = a[13] & g[15872];
assign g[32255] = b[13] & g[15872];
assign g[24065] = a[13] & g[15873];
assign g[32256] = b[13] & g[15873];
assign g[24066] = a[13] & g[15874];
assign g[32257] = b[13] & g[15874];
assign g[24067] = a[13] & g[15875];
assign g[32258] = b[13] & g[15875];
assign g[24068] = a[13] & g[15876];
assign g[32259] = b[13] & g[15876];
assign g[24069] = a[13] & g[15877];
assign g[32260] = b[13] & g[15877];
assign g[24070] = a[13] & g[15878];
assign g[32261] = b[13] & g[15878];
assign g[24071] = a[13] & g[15879];
assign g[32262] = b[13] & g[15879];
assign g[24072] = a[13] & g[15880];
assign g[32263] = b[13] & g[15880];
assign g[24073] = a[13] & g[15881];
assign g[32264] = b[13] & g[15881];
assign g[24074] = a[13] & g[15882];
assign g[32265] = b[13] & g[15882];
assign g[24075] = a[13] & g[15883];
assign g[32266] = b[13] & g[15883];
assign g[24076] = a[13] & g[15884];
assign g[32267] = b[13] & g[15884];
assign g[24077] = a[13] & g[15885];
assign g[32268] = b[13] & g[15885];
assign g[24078] = a[13] & g[15886];
assign g[32269] = b[13] & g[15886];
assign g[24079] = a[13] & g[15887];
assign g[32270] = b[13] & g[15887];
assign g[24080] = a[13] & g[15888];
assign g[32271] = b[13] & g[15888];
assign g[24081] = a[13] & g[15889];
assign g[32272] = b[13] & g[15889];
assign g[24082] = a[13] & g[15890];
assign g[32273] = b[13] & g[15890];
assign g[24083] = a[13] & g[15891];
assign g[32274] = b[13] & g[15891];
assign g[24084] = a[13] & g[15892];
assign g[32275] = b[13] & g[15892];
assign g[24085] = a[13] & g[15893];
assign g[32276] = b[13] & g[15893];
assign g[24086] = a[13] & g[15894];
assign g[32277] = b[13] & g[15894];
assign g[24087] = a[13] & g[15895];
assign g[32278] = b[13] & g[15895];
assign g[24088] = a[13] & g[15896];
assign g[32279] = b[13] & g[15896];
assign g[24089] = a[13] & g[15897];
assign g[32280] = b[13] & g[15897];
assign g[24090] = a[13] & g[15898];
assign g[32281] = b[13] & g[15898];
assign g[24091] = a[13] & g[15899];
assign g[32282] = b[13] & g[15899];
assign g[24092] = a[13] & g[15900];
assign g[32283] = b[13] & g[15900];
assign g[24093] = a[13] & g[15901];
assign g[32284] = b[13] & g[15901];
assign g[24094] = a[13] & g[15902];
assign g[32285] = b[13] & g[15902];
assign g[24095] = a[13] & g[15903];
assign g[32286] = b[13] & g[15903];
assign g[24096] = a[13] & g[15904];
assign g[32287] = b[13] & g[15904];
assign g[24097] = a[13] & g[15905];
assign g[32288] = b[13] & g[15905];
assign g[24098] = a[13] & g[15906];
assign g[32289] = b[13] & g[15906];
assign g[24099] = a[13] & g[15907];
assign g[32290] = b[13] & g[15907];
assign g[24100] = a[13] & g[15908];
assign g[32291] = b[13] & g[15908];
assign g[24101] = a[13] & g[15909];
assign g[32292] = b[13] & g[15909];
assign g[24102] = a[13] & g[15910];
assign g[32293] = b[13] & g[15910];
assign g[24103] = a[13] & g[15911];
assign g[32294] = b[13] & g[15911];
assign g[24104] = a[13] & g[15912];
assign g[32295] = b[13] & g[15912];
assign g[24105] = a[13] & g[15913];
assign g[32296] = b[13] & g[15913];
assign g[24106] = a[13] & g[15914];
assign g[32297] = b[13] & g[15914];
assign g[24107] = a[13] & g[15915];
assign g[32298] = b[13] & g[15915];
assign g[24108] = a[13] & g[15916];
assign g[32299] = b[13] & g[15916];
assign g[24109] = a[13] & g[15917];
assign g[32300] = b[13] & g[15917];
assign g[24110] = a[13] & g[15918];
assign g[32301] = b[13] & g[15918];
assign g[24111] = a[13] & g[15919];
assign g[32302] = b[13] & g[15919];
assign g[24112] = a[13] & g[15920];
assign g[32303] = b[13] & g[15920];
assign g[24113] = a[13] & g[15921];
assign g[32304] = b[13] & g[15921];
assign g[24114] = a[13] & g[15922];
assign g[32305] = b[13] & g[15922];
assign g[24115] = a[13] & g[15923];
assign g[32306] = b[13] & g[15923];
assign g[24116] = a[13] & g[15924];
assign g[32307] = b[13] & g[15924];
assign g[24117] = a[13] & g[15925];
assign g[32308] = b[13] & g[15925];
assign g[24118] = a[13] & g[15926];
assign g[32309] = b[13] & g[15926];
assign g[24119] = a[13] & g[15927];
assign g[32310] = b[13] & g[15927];
assign g[24120] = a[13] & g[15928];
assign g[32311] = b[13] & g[15928];
assign g[24121] = a[13] & g[15929];
assign g[32312] = b[13] & g[15929];
assign g[24122] = a[13] & g[15930];
assign g[32313] = b[13] & g[15930];
assign g[24123] = a[13] & g[15931];
assign g[32314] = b[13] & g[15931];
assign g[24124] = a[13] & g[15932];
assign g[32315] = b[13] & g[15932];
assign g[24125] = a[13] & g[15933];
assign g[32316] = b[13] & g[15933];
assign g[24126] = a[13] & g[15934];
assign g[32317] = b[13] & g[15934];
assign g[24127] = a[13] & g[15935];
assign g[32318] = b[13] & g[15935];
assign g[24128] = a[13] & g[15936];
assign g[32319] = b[13] & g[15936];
assign g[24129] = a[13] & g[15937];
assign g[32320] = b[13] & g[15937];
assign g[24130] = a[13] & g[15938];
assign g[32321] = b[13] & g[15938];
assign g[24131] = a[13] & g[15939];
assign g[32322] = b[13] & g[15939];
assign g[24132] = a[13] & g[15940];
assign g[32323] = b[13] & g[15940];
assign g[24133] = a[13] & g[15941];
assign g[32324] = b[13] & g[15941];
assign g[24134] = a[13] & g[15942];
assign g[32325] = b[13] & g[15942];
assign g[24135] = a[13] & g[15943];
assign g[32326] = b[13] & g[15943];
assign g[24136] = a[13] & g[15944];
assign g[32327] = b[13] & g[15944];
assign g[24137] = a[13] & g[15945];
assign g[32328] = b[13] & g[15945];
assign g[24138] = a[13] & g[15946];
assign g[32329] = b[13] & g[15946];
assign g[24139] = a[13] & g[15947];
assign g[32330] = b[13] & g[15947];
assign g[24140] = a[13] & g[15948];
assign g[32331] = b[13] & g[15948];
assign g[24141] = a[13] & g[15949];
assign g[32332] = b[13] & g[15949];
assign g[24142] = a[13] & g[15950];
assign g[32333] = b[13] & g[15950];
assign g[24143] = a[13] & g[15951];
assign g[32334] = b[13] & g[15951];
assign g[24144] = a[13] & g[15952];
assign g[32335] = b[13] & g[15952];
assign g[24145] = a[13] & g[15953];
assign g[32336] = b[13] & g[15953];
assign g[24146] = a[13] & g[15954];
assign g[32337] = b[13] & g[15954];
assign g[24147] = a[13] & g[15955];
assign g[32338] = b[13] & g[15955];
assign g[24148] = a[13] & g[15956];
assign g[32339] = b[13] & g[15956];
assign g[24149] = a[13] & g[15957];
assign g[32340] = b[13] & g[15957];
assign g[24150] = a[13] & g[15958];
assign g[32341] = b[13] & g[15958];
assign g[24151] = a[13] & g[15959];
assign g[32342] = b[13] & g[15959];
assign g[24152] = a[13] & g[15960];
assign g[32343] = b[13] & g[15960];
assign g[24153] = a[13] & g[15961];
assign g[32344] = b[13] & g[15961];
assign g[24154] = a[13] & g[15962];
assign g[32345] = b[13] & g[15962];
assign g[24155] = a[13] & g[15963];
assign g[32346] = b[13] & g[15963];
assign g[24156] = a[13] & g[15964];
assign g[32347] = b[13] & g[15964];
assign g[24157] = a[13] & g[15965];
assign g[32348] = b[13] & g[15965];
assign g[24158] = a[13] & g[15966];
assign g[32349] = b[13] & g[15966];
assign g[24159] = a[13] & g[15967];
assign g[32350] = b[13] & g[15967];
assign g[24160] = a[13] & g[15968];
assign g[32351] = b[13] & g[15968];
assign g[24161] = a[13] & g[15969];
assign g[32352] = b[13] & g[15969];
assign g[24162] = a[13] & g[15970];
assign g[32353] = b[13] & g[15970];
assign g[24163] = a[13] & g[15971];
assign g[32354] = b[13] & g[15971];
assign g[24164] = a[13] & g[15972];
assign g[32355] = b[13] & g[15972];
assign g[24165] = a[13] & g[15973];
assign g[32356] = b[13] & g[15973];
assign g[24166] = a[13] & g[15974];
assign g[32357] = b[13] & g[15974];
assign g[24167] = a[13] & g[15975];
assign g[32358] = b[13] & g[15975];
assign g[24168] = a[13] & g[15976];
assign g[32359] = b[13] & g[15976];
assign g[24169] = a[13] & g[15977];
assign g[32360] = b[13] & g[15977];
assign g[24170] = a[13] & g[15978];
assign g[32361] = b[13] & g[15978];
assign g[24171] = a[13] & g[15979];
assign g[32362] = b[13] & g[15979];
assign g[24172] = a[13] & g[15980];
assign g[32363] = b[13] & g[15980];
assign g[24173] = a[13] & g[15981];
assign g[32364] = b[13] & g[15981];
assign g[24174] = a[13] & g[15982];
assign g[32365] = b[13] & g[15982];
assign g[24175] = a[13] & g[15983];
assign g[32366] = b[13] & g[15983];
assign g[24176] = a[13] & g[15984];
assign g[32367] = b[13] & g[15984];
assign g[24177] = a[13] & g[15985];
assign g[32368] = b[13] & g[15985];
assign g[24178] = a[13] & g[15986];
assign g[32369] = b[13] & g[15986];
assign g[24179] = a[13] & g[15987];
assign g[32370] = b[13] & g[15987];
assign g[24180] = a[13] & g[15988];
assign g[32371] = b[13] & g[15988];
assign g[24181] = a[13] & g[15989];
assign g[32372] = b[13] & g[15989];
assign g[24182] = a[13] & g[15990];
assign g[32373] = b[13] & g[15990];
assign g[24183] = a[13] & g[15991];
assign g[32374] = b[13] & g[15991];
assign g[24184] = a[13] & g[15992];
assign g[32375] = b[13] & g[15992];
assign g[24185] = a[13] & g[15993];
assign g[32376] = b[13] & g[15993];
assign g[24186] = a[13] & g[15994];
assign g[32377] = b[13] & g[15994];
assign g[24187] = a[13] & g[15995];
assign g[32378] = b[13] & g[15995];
assign g[24188] = a[13] & g[15996];
assign g[32379] = b[13] & g[15996];
assign g[24189] = a[13] & g[15997];
assign g[32380] = b[13] & g[15997];
assign g[24190] = a[13] & g[15998];
assign g[32381] = b[13] & g[15998];
assign g[24191] = a[13] & g[15999];
assign g[32382] = b[13] & g[15999];
assign g[24192] = a[13] & g[16000];
assign g[32383] = b[13] & g[16000];
assign g[24193] = a[13] & g[16001];
assign g[32384] = b[13] & g[16001];
assign g[24194] = a[13] & g[16002];
assign g[32385] = b[13] & g[16002];
assign g[24195] = a[13] & g[16003];
assign g[32386] = b[13] & g[16003];
assign g[24196] = a[13] & g[16004];
assign g[32387] = b[13] & g[16004];
assign g[24197] = a[13] & g[16005];
assign g[32388] = b[13] & g[16005];
assign g[24198] = a[13] & g[16006];
assign g[32389] = b[13] & g[16006];
assign g[24199] = a[13] & g[16007];
assign g[32390] = b[13] & g[16007];
assign g[24200] = a[13] & g[16008];
assign g[32391] = b[13] & g[16008];
assign g[24201] = a[13] & g[16009];
assign g[32392] = b[13] & g[16009];
assign g[24202] = a[13] & g[16010];
assign g[32393] = b[13] & g[16010];
assign g[24203] = a[13] & g[16011];
assign g[32394] = b[13] & g[16011];
assign g[24204] = a[13] & g[16012];
assign g[32395] = b[13] & g[16012];
assign g[24205] = a[13] & g[16013];
assign g[32396] = b[13] & g[16013];
assign g[24206] = a[13] & g[16014];
assign g[32397] = b[13] & g[16014];
assign g[24207] = a[13] & g[16015];
assign g[32398] = b[13] & g[16015];
assign g[24208] = a[13] & g[16016];
assign g[32399] = b[13] & g[16016];
assign g[24209] = a[13] & g[16017];
assign g[32400] = b[13] & g[16017];
assign g[24210] = a[13] & g[16018];
assign g[32401] = b[13] & g[16018];
assign g[24211] = a[13] & g[16019];
assign g[32402] = b[13] & g[16019];
assign g[24212] = a[13] & g[16020];
assign g[32403] = b[13] & g[16020];
assign g[24213] = a[13] & g[16021];
assign g[32404] = b[13] & g[16021];
assign g[24214] = a[13] & g[16022];
assign g[32405] = b[13] & g[16022];
assign g[24215] = a[13] & g[16023];
assign g[32406] = b[13] & g[16023];
assign g[24216] = a[13] & g[16024];
assign g[32407] = b[13] & g[16024];
assign g[24217] = a[13] & g[16025];
assign g[32408] = b[13] & g[16025];
assign g[24218] = a[13] & g[16026];
assign g[32409] = b[13] & g[16026];
assign g[24219] = a[13] & g[16027];
assign g[32410] = b[13] & g[16027];
assign g[24220] = a[13] & g[16028];
assign g[32411] = b[13] & g[16028];
assign g[24221] = a[13] & g[16029];
assign g[32412] = b[13] & g[16029];
assign g[24222] = a[13] & g[16030];
assign g[32413] = b[13] & g[16030];
assign g[24223] = a[13] & g[16031];
assign g[32414] = b[13] & g[16031];
assign g[24224] = a[13] & g[16032];
assign g[32415] = b[13] & g[16032];
assign g[24225] = a[13] & g[16033];
assign g[32416] = b[13] & g[16033];
assign g[24226] = a[13] & g[16034];
assign g[32417] = b[13] & g[16034];
assign g[24227] = a[13] & g[16035];
assign g[32418] = b[13] & g[16035];
assign g[24228] = a[13] & g[16036];
assign g[32419] = b[13] & g[16036];
assign g[24229] = a[13] & g[16037];
assign g[32420] = b[13] & g[16037];
assign g[24230] = a[13] & g[16038];
assign g[32421] = b[13] & g[16038];
assign g[24231] = a[13] & g[16039];
assign g[32422] = b[13] & g[16039];
assign g[24232] = a[13] & g[16040];
assign g[32423] = b[13] & g[16040];
assign g[24233] = a[13] & g[16041];
assign g[32424] = b[13] & g[16041];
assign g[24234] = a[13] & g[16042];
assign g[32425] = b[13] & g[16042];
assign g[24235] = a[13] & g[16043];
assign g[32426] = b[13] & g[16043];
assign g[24236] = a[13] & g[16044];
assign g[32427] = b[13] & g[16044];
assign g[24237] = a[13] & g[16045];
assign g[32428] = b[13] & g[16045];
assign g[24238] = a[13] & g[16046];
assign g[32429] = b[13] & g[16046];
assign g[24239] = a[13] & g[16047];
assign g[32430] = b[13] & g[16047];
assign g[24240] = a[13] & g[16048];
assign g[32431] = b[13] & g[16048];
assign g[24241] = a[13] & g[16049];
assign g[32432] = b[13] & g[16049];
assign g[24242] = a[13] & g[16050];
assign g[32433] = b[13] & g[16050];
assign g[24243] = a[13] & g[16051];
assign g[32434] = b[13] & g[16051];
assign g[24244] = a[13] & g[16052];
assign g[32435] = b[13] & g[16052];
assign g[24245] = a[13] & g[16053];
assign g[32436] = b[13] & g[16053];
assign g[24246] = a[13] & g[16054];
assign g[32437] = b[13] & g[16054];
assign g[24247] = a[13] & g[16055];
assign g[32438] = b[13] & g[16055];
assign g[24248] = a[13] & g[16056];
assign g[32439] = b[13] & g[16056];
assign g[24249] = a[13] & g[16057];
assign g[32440] = b[13] & g[16057];
assign g[24250] = a[13] & g[16058];
assign g[32441] = b[13] & g[16058];
assign g[24251] = a[13] & g[16059];
assign g[32442] = b[13] & g[16059];
assign g[24252] = a[13] & g[16060];
assign g[32443] = b[13] & g[16060];
assign g[24253] = a[13] & g[16061];
assign g[32444] = b[13] & g[16061];
assign g[24254] = a[13] & g[16062];
assign g[32445] = b[13] & g[16062];
assign g[24255] = a[13] & g[16063];
assign g[32446] = b[13] & g[16063];
assign g[24256] = a[13] & g[16064];
assign g[32447] = b[13] & g[16064];
assign g[24257] = a[13] & g[16065];
assign g[32448] = b[13] & g[16065];
assign g[24258] = a[13] & g[16066];
assign g[32449] = b[13] & g[16066];
assign g[24259] = a[13] & g[16067];
assign g[32450] = b[13] & g[16067];
assign g[24260] = a[13] & g[16068];
assign g[32451] = b[13] & g[16068];
assign g[24261] = a[13] & g[16069];
assign g[32452] = b[13] & g[16069];
assign g[24262] = a[13] & g[16070];
assign g[32453] = b[13] & g[16070];
assign g[24263] = a[13] & g[16071];
assign g[32454] = b[13] & g[16071];
assign g[24264] = a[13] & g[16072];
assign g[32455] = b[13] & g[16072];
assign g[24265] = a[13] & g[16073];
assign g[32456] = b[13] & g[16073];
assign g[24266] = a[13] & g[16074];
assign g[32457] = b[13] & g[16074];
assign g[24267] = a[13] & g[16075];
assign g[32458] = b[13] & g[16075];
assign g[24268] = a[13] & g[16076];
assign g[32459] = b[13] & g[16076];
assign g[24269] = a[13] & g[16077];
assign g[32460] = b[13] & g[16077];
assign g[24270] = a[13] & g[16078];
assign g[32461] = b[13] & g[16078];
assign g[24271] = a[13] & g[16079];
assign g[32462] = b[13] & g[16079];
assign g[24272] = a[13] & g[16080];
assign g[32463] = b[13] & g[16080];
assign g[24273] = a[13] & g[16081];
assign g[32464] = b[13] & g[16081];
assign g[24274] = a[13] & g[16082];
assign g[32465] = b[13] & g[16082];
assign g[24275] = a[13] & g[16083];
assign g[32466] = b[13] & g[16083];
assign g[24276] = a[13] & g[16084];
assign g[32467] = b[13] & g[16084];
assign g[24277] = a[13] & g[16085];
assign g[32468] = b[13] & g[16085];
assign g[24278] = a[13] & g[16086];
assign g[32469] = b[13] & g[16086];
assign g[24279] = a[13] & g[16087];
assign g[32470] = b[13] & g[16087];
assign g[24280] = a[13] & g[16088];
assign g[32471] = b[13] & g[16088];
assign g[24281] = a[13] & g[16089];
assign g[32472] = b[13] & g[16089];
assign g[24282] = a[13] & g[16090];
assign g[32473] = b[13] & g[16090];
assign g[24283] = a[13] & g[16091];
assign g[32474] = b[13] & g[16091];
assign g[24284] = a[13] & g[16092];
assign g[32475] = b[13] & g[16092];
assign g[24285] = a[13] & g[16093];
assign g[32476] = b[13] & g[16093];
assign g[24286] = a[13] & g[16094];
assign g[32477] = b[13] & g[16094];
assign g[24287] = a[13] & g[16095];
assign g[32478] = b[13] & g[16095];
assign g[24288] = a[13] & g[16096];
assign g[32479] = b[13] & g[16096];
assign g[24289] = a[13] & g[16097];
assign g[32480] = b[13] & g[16097];
assign g[24290] = a[13] & g[16098];
assign g[32481] = b[13] & g[16098];
assign g[24291] = a[13] & g[16099];
assign g[32482] = b[13] & g[16099];
assign g[24292] = a[13] & g[16100];
assign g[32483] = b[13] & g[16100];
assign g[24293] = a[13] & g[16101];
assign g[32484] = b[13] & g[16101];
assign g[24294] = a[13] & g[16102];
assign g[32485] = b[13] & g[16102];
assign g[24295] = a[13] & g[16103];
assign g[32486] = b[13] & g[16103];
assign g[24296] = a[13] & g[16104];
assign g[32487] = b[13] & g[16104];
assign g[24297] = a[13] & g[16105];
assign g[32488] = b[13] & g[16105];
assign g[24298] = a[13] & g[16106];
assign g[32489] = b[13] & g[16106];
assign g[24299] = a[13] & g[16107];
assign g[32490] = b[13] & g[16107];
assign g[24300] = a[13] & g[16108];
assign g[32491] = b[13] & g[16108];
assign g[24301] = a[13] & g[16109];
assign g[32492] = b[13] & g[16109];
assign g[24302] = a[13] & g[16110];
assign g[32493] = b[13] & g[16110];
assign g[24303] = a[13] & g[16111];
assign g[32494] = b[13] & g[16111];
assign g[24304] = a[13] & g[16112];
assign g[32495] = b[13] & g[16112];
assign g[24305] = a[13] & g[16113];
assign g[32496] = b[13] & g[16113];
assign g[24306] = a[13] & g[16114];
assign g[32497] = b[13] & g[16114];
assign g[24307] = a[13] & g[16115];
assign g[32498] = b[13] & g[16115];
assign g[24308] = a[13] & g[16116];
assign g[32499] = b[13] & g[16116];
assign g[24309] = a[13] & g[16117];
assign g[32500] = b[13] & g[16117];
assign g[24310] = a[13] & g[16118];
assign g[32501] = b[13] & g[16118];
assign g[24311] = a[13] & g[16119];
assign g[32502] = b[13] & g[16119];
assign g[24312] = a[13] & g[16120];
assign g[32503] = b[13] & g[16120];
assign g[24313] = a[13] & g[16121];
assign g[32504] = b[13] & g[16121];
assign g[24314] = a[13] & g[16122];
assign g[32505] = b[13] & g[16122];
assign g[24315] = a[13] & g[16123];
assign g[32506] = b[13] & g[16123];
assign g[24316] = a[13] & g[16124];
assign g[32507] = b[13] & g[16124];
assign g[24317] = a[13] & g[16125];
assign g[32508] = b[13] & g[16125];
assign g[24318] = a[13] & g[16126];
assign g[32509] = b[13] & g[16126];
assign g[24319] = a[13] & g[16127];
assign g[32510] = b[13] & g[16127];
assign g[24320] = a[13] & g[16128];
assign g[32511] = b[13] & g[16128];
assign g[24321] = a[13] & g[16129];
assign g[32512] = b[13] & g[16129];
assign g[24322] = a[13] & g[16130];
assign g[32513] = b[13] & g[16130];
assign g[24323] = a[13] & g[16131];
assign g[32514] = b[13] & g[16131];
assign g[24324] = a[13] & g[16132];
assign g[32515] = b[13] & g[16132];
assign g[24325] = a[13] & g[16133];
assign g[32516] = b[13] & g[16133];
assign g[24326] = a[13] & g[16134];
assign g[32517] = b[13] & g[16134];
assign g[24327] = a[13] & g[16135];
assign g[32518] = b[13] & g[16135];
assign g[24328] = a[13] & g[16136];
assign g[32519] = b[13] & g[16136];
assign g[24329] = a[13] & g[16137];
assign g[32520] = b[13] & g[16137];
assign g[24330] = a[13] & g[16138];
assign g[32521] = b[13] & g[16138];
assign g[24331] = a[13] & g[16139];
assign g[32522] = b[13] & g[16139];
assign g[24332] = a[13] & g[16140];
assign g[32523] = b[13] & g[16140];
assign g[24333] = a[13] & g[16141];
assign g[32524] = b[13] & g[16141];
assign g[24334] = a[13] & g[16142];
assign g[32525] = b[13] & g[16142];
assign g[24335] = a[13] & g[16143];
assign g[32526] = b[13] & g[16143];
assign g[24336] = a[13] & g[16144];
assign g[32527] = b[13] & g[16144];
assign g[24337] = a[13] & g[16145];
assign g[32528] = b[13] & g[16145];
assign g[24338] = a[13] & g[16146];
assign g[32529] = b[13] & g[16146];
assign g[24339] = a[13] & g[16147];
assign g[32530] = b[13] & g[16147];
assign g[24340] = a[13] & g[16148];
assign g[32531] = b[13] & g[16148];
assign g[24341] = a[13] & g[16149];
assign g[32532] = b[13] & g[16149];
assign g[24342] = a[13] & g[16150];
assign g[32533] = b[13] & g[16150];
assign g[24343] = a[13] & g[16151];
assign g[32534] = b[13] & g[16151];
assign g[24344] = a[13] & g[16152];
assign g[32535] = b[13] & g[16152];
assign g[24345] = a[13] & g[16153];
assign g[32536] = b[13] & g[16153];
assign g[24346] = a[13] & g[16154];
assign g[32537] = b[13] & g[16154];
assign g[24347] = a[13] & g[16155];
assign g[32538] = b[13] & g[16155];
assign g[24348] = a[13] & g[16156];
assign g[32539] = b[13] & g[16156];
assign g[24349] = a[13] & g[16157];
assign g[32540] = b[13] & g[16157];
assign g[24350] = a[13] & g[16158];
assign g[32541] = b[13] & g[16158];
assign g[24351] = a[13] & g[16159];
assign g[32542] = b[13] & g[16159];
assign g[24352] = a[13] & g[16160];
assign g[32543] = b[13] & g[16160];
assign g[24353] = a[13] & g[16161];
assign g[32544] = b[13] & g[16161];
assign g[24354] = a[13] & g[16162];
assign g[32545] = b[13] & g[16162];
assign g[24355] = a[13] & g[16163];
assign g[32546] = b[13] & g[16163];
assign g[24356] = a[13] & g[16164];
assign g[32547] = b[13] & g[16164];
assign g[24357] = a[13] & g[16165];
assign g[32548] = b[13] & g[16165];
assign g[24358] = a[13] & g[16166];
assign g[32549] = b[13] & g[16166];
assign g[24359] = a[13] & g[16167];
assign g[32550] = b[13] & g[16167];
assign g[24360] = a[13] & g[16168];
assign g[32551] = b[13] & g[16168];
assign g[24361] = a[13] & g[16169];
assign g[32552] = b[13] & g[16169];
assign g[24362] = a[13] & g[16170];
assign g[32553] = b[13] & g[16170];
assign g[24363] = a[13] & g[16171];
assign g[32554] = b[13] & g[16171];
assign g[24364] = a[13] & g[16172];
assign g[32555] = b[13] & g[16172];
assign g[24365] = a[13] & g[16173];
assign g[32556] = b[13] & g[16173];
assign g[24366] = a[13] & g[16174];
assign g[32557] = b[13] & g[16174];
assign g[24367] = a[13] & g[16175];
assign g[32558] = b[13] & g[16175];
assign g[24368] = a[13] & g[16176];
assign g[32559] = b[13] & g[16176];
assign g[24369] = a[13] & g[16177];
assign g[32560] = b[13] & g[16177];
assign g[24370] = a[13] & g[16178];
assign g[32561] = b[13] & g[16178];
assign g[24371] = a[13] & g[16179];
assign g[32562] = b[13] & g[16179];
assign g[24372] = a[13] & g[16180];
assign g[32563] = b[13] & g[16180];
assign g[24373] = a[13] & g[16181];
assign g[32564] = b[13] & g[16181];
assign g[24374] = a[13] & g[16182];
assign g[32565] = b[13] & g[16182];
assign g[24375] = a[13] & g[16183];
assign g[32566] = b[13] & g[16183];
assign g[24376] = a[13] & g[16184];
assign g[32567] = b[13] & g[16184];
assign g[24377] = a[13] & g[16185];
assign g[32568] = b[13] & g[16185];
assign g[24378] = a[13] & g[16186];
assign g[32569] = b[13] & g[16186];
assign g[24379] = a[13] & g[16187];
assign g[32570] = b[13] & g[16187];
assign g[24380] = a[13] & g[16188];
assign g[32571] = b[13] & g[16188];
assign g[24381] = a[13] & g[16189];
assign g[32572] = b[13] & g[16189];
assign g[24382] = a[13] & g[16190];
assign g[32573] = b[13] & g[16190];
assign g[24383] = a[13] & g[16191];
assign g[32574] = b[13] & g[16191];
assign g[24384] = a[13] & g[16192];
assign g[32575] = b[13] & g[16192];
assign g[24385] = a[13] & g[16193];
assign g[32576] = b[13] & g[16193];
assign g[24386] = a[13] & g[16194];
assign g[32577] = b[13] & g[16194];
assign g[24387] = a[13] & g[16195];
assign g[32578] = b[13] & g[16195];
assign g[24388] = a[13] & g[16196];
assign g[32579] = b[13] & g[16196];
assign g[24389] = a[13] & g[16197];
assign g[32580] = b[13] & g[16197];
assign g[24390] = a[13] & g[16198];
assign g[32581] = b[13] & g[16198];
assign g[24391] = a[13] & g[16199];
assign g[32582] = b[13] & g[16199];
assign g[24392] = a[13] & g[16200];
assign g[32583] = b[13] & g[16200];
assign g[24393] = a[13] & g[16201];
assign g[32584] = b[13] & g[16201];
assign g[24394] = a[13] & g[16202];
assign g[32585] = b[13] & g[16202];
assign g[24395] = a[13] & g[16203];
assign g[32586] = b[13] & g[16203];
assign g[24396] = a[13] & g[16204];
assign g[32587] = b[13] & g[16204];
assign g[24397] = a[13] & g[16205];
assign g[32588] = b[13] & g[16205];
assign g[24398] = a[13] & g[16206];
assign g[32589] = b[13] & g[16206];
assign g[24399] = a[13] & g[16207];
assign g[32590] = b[13] & g[16207];
assign g[24400] = a[13] & g[16208];
assign g[32591] = b[13] & g[16208];
assign g[24401] = a[13] & g[16209];
assign g[32592] = b[13] & g[16209];
assign g[24402] = a[13] & g[16210];
assign g[32593] = b[13] & g[16210];
assign g[24403] = a[13] & g[16211];
assign g[32594] = b[13] & g[16211];
assign g[24404] = a[13] & g[16212];
assign g[32595] = b[13] & g[16212];
assign g[24405] = a[13] & g[16213];
assign g[32596] = b[13] & g[16213];
assign g[24406] = a[13] & g[16214];
assign g[32597] = b[13] & g[16214];
assign g[24407] = a[13] & g[16215];
assign g[32598] = b[13] & g[16215];
assign g[24408] = a[13] & g[16216];
assign g[32599] = b[13] & g[16216];
assign g[24409] = a[13] & g[16217];
assign g[32600] = b[13] & g[16217];
assign g[24410] = a[13] & g[16218];
assign g[32601] = b[13] & g[16218];
assign g[24411] = a[13] & g[16219];
assign g[32602] = b[13] & g[16219];
assign g[24412] = a[13] & g[16220];
assign g[32603] = b[13] & g[16220];
assign g[24413] = a[13] & g[16221];
assign g[32604] = b[13] & g[16221];
assign g[24414] = a[13] & g[16222];
assign g[32605] = b[13] & g[16222];
assign g[24415] = a[13] & g[16223];
assign g[32606] = b[13] & g[16223];
assign g[24416] = a[13] & g[16224];
assign g[32607] = b[13] & g[16224];
assign g[24417] = a[13] & g[16225];
assign g[32608] = b[13] & g[16225];
assign g[24418] = a[13] & g[16226];
assign g[32609] = b[13] & g[16226];
assign g[24419] = a[13] & g[16227];
assign g[32610] = b[13] & g[16227];
assign g[24420] = a[13] & g[16228];
assign g[32611] = b[13] & g[16228];
assign g[24421] = a[13] & g[16229];
assign g[32612] = b[13] & g[16229];
assign g[24422] = a[13] & g[16230];
assign g[32613] = b[13] & g[16230];
assign g[24423] = a[13] & g[16231];
assign g[32614] = b[13] & g[16231];
assign g[24424] = a[13] & g[16232];
assign g[32615] = b[13] & g[16232];
assign g[24425] = a[13] & g[16233];
assign g[32616] = b[13] & g[16233];
assign g[24426] = a[13] & g[16234];
assign g[32617] = b[13] & g[16234];
assign g[24427] = a[13] & g[16235];
assign g[32618] = b[13] & g[16235];
assign g[24428] = a[13] & g[16236];
assign g[32619] = b[13] & g[16236];
assign g[24429] = a[13] & g[16237];
assign g[32620] = b[13] & g[16237];
assign g[24430] = a[13] & g[16238];
assign g[32621] = b[13] & g[16238];
assign g[24431] = a[13] & g[16239];
assign g[32622] = b[13] & g[16239];
assign g[24432] = a[13] & g[16240];
assign g[32623] = b[13] & g[16240];
assign g[24433] = a[13] & g[16241];
assign g[32624] = b[13] & g[16241];
assign g[24434] = a[13] & g[16242];
assign g[32625] = b[13] & g[16242];
assign g[24435] = a[13] & g[16243];
assign g[32626] = b[13] & g[16243];
assign g[24436] = a[13] & g[16244];
assign g[32627] = b[13] & g[16244];
assign g[24437] = a[13] & g[16245];
assign g[32628] = b[13] & g[16245];
assign g[24438] = a[13] & g[16246];
assign g[32629] = b[13] & g[16246];
assign g[24439] = a[13] & g[16247];
assign g[32630] = b[13] & g[16247];
assign g[24440] = a[13] & g[16248];
assign g[32631] = b[13] & g[16248];
assign g[24441] = a[13] & g[16249];
assign g[32632] = b[13] & g[16249];
assign g[24442] = a[13] & g[16250];
assign g[32633] = b[13] & g[16250];
assign g[24443] = a[13] & g[16251];
assign g[32634] = b[13] & g[16251];
assign g[24444] = a[13] & g[16252];
assign g[32635] = b[13] & g[16252];
assign g[24445] = a[13] & g[16253];
assign g[32636] = b[13] & g[16253];
assign g[24446] = a[13] & g[16254];
assign g[32637] = b[13] & g[16254];
assign g[24447] = a[13] & g[16255];
assign g[32638] = b[13] & g[16255];
assign g[24448] = a[13] & g[16256];
assign g[32639] = b[13] & g[16256];
assign g[24449] = a[13] & g[16257];
assign g[32640] = b[13] & g[16257];
assign g[24450] = a[13] & g[16258];
assign g[32641] = b[13] & g[16258];
assign g[24451] = a[13] & g[16259];
assign g[32642] = b[13] & g[16259];
assign g[24452] = a[13] & g[16260];
assign g[32643] = b[13] & g[16260];
assign g[24453] = a[13] & g[16261];
assign g[32644] = b[13] & g[16261];
assign g[24454] = a[13] & g[16262];
assign g[32645] = b[13] & g[16262];
assign g[24455] = a[13] & g[16263];
assign g[32646] = b[13] & g[16263];
assign g[24456] = a[13] & g[16264];
assign g[32647] = b[13] & g[16264];
assign g[24457] = a[13] & g[16265];
assign g[32648] = b[13] & g[16265];
assign g[24458] = a[13] & g[16266];
assign g[32649] = b[13] & g[16266];
assign g[24459] = a[13] & g[16267];
assign g[32650] = b[13] & g[16267];
assign g[24460] = a[13] & g[16268];
assign g[32651] = b[13] & g[16268];
assign g[24461] = a[13] & g[16269];
assign g[32652] = b[13] & g[16269];
assign g[24462] = a[13] & g[16270];
assign g[32653] = b[13] & g[16270];
assign g[24463] = a[13] & g[16271];
assign g[32654] = b[13] & g[16271];
assign g[24464] = a[13] & g[16272];
assign g[32655] = b[13] & g[16272];
assign g[24465] = a[13] & g[16273];
assign g[32656] = b[13] & g[16273];
assign g[24466] = a[13] & g[16274];
assign g[32657] = b[13] & g[16274];
assign g[24467] = a[13] & g[16275];
assign g[32658] = b[13] & g[16275];
assign g[24468] = a[13] & g[16276];
assign g[32659] = b[13] & g[16276];
assign g[24469] = a[13] & g[16277];
assign g[32660] = b[13] & g[16277];
assign g[24470] = a[13] & g[16278];
assign g[32661] = b[13] & g[16278];
assign g[24471] = a[13] & g[16279];
assign g[32662] = b[13] & g[16279];
assign g[24472] = a[13] & g[16280];
assign g[32663] = b[13] & g[16280];
assign g[24473] = a[13] & g[16281];
assign g[32664] = b[13] & g[16281];
assign g[24474] = a[13] & g[16282];
assign g[32665] = b[13] & g[16282];
assign g[24475] = a[13] & g[16283];
assign g[32666] = b[13] & g[16283];
assign g[24476] = a[13] & g[16284];
assign g[32667] = b[13] & g[16284];
assign g[24477] = a[13] & g[16285];
assign g[32668] = b[13] & g[16285];
assign g[24478] = a[13] & g[16286];
assign g[32669] = b[13] & g[16286];
assign g[24479] = a[13] & g[16287];
assign g[32670] = b[13] & g[16287];
assign g[24480] = a[13] & g[16288];
assign g[32671] = b[13] & g[16288];
assign g[24481] = a[13] & g[16289];
assign g[32672] = b[13] & g[16289];
assign g[24482] = a[13] & g[16290];
assign g[32673] = b[13] & g[16290];
assign g[24483] = a[13] & g[16291];
assign g[32674] = b[13] & g[16291];
assign g[24484] = a[13] & g[16292];
assign g[32675] = b[13] & g[16292];
assign g[24485] = a[13] & g[16293];
assign g[32676] = b[13] & g[16293];
assign g[24486] = a[13] & g[16294];
assign g[32677] = b[13] & g[16294];
assign g[24487] = a[13] & g[16295];
assign g[32678] = b[13] & g[16295];
assign g[24488] = a[13] & g[16296];
assign g[32679] = b[13] & g[16296];
assign g[24489] = a[13] & g[16297];
assign g[32680] = b[13] & g[16297];
assign g[24490] = a[13] & g[16298];
assign g[32681] = b[13] & g[16298];
assign g[24491] = a[13] & g[16299];
assign g[32682] = b[13] & g[16299];
assign g[24492] = a[13] & g[16300];
assign g[32683] = b[13] & g[16300];
assign g[24493] = a[13] & g[16301];
assign g[32684] = b[13] & g[16301];
assign g[24494] = a[13] & g[16302];
assign g[32685] = b[13] & g[16302];
assign g[24495] = a[13] & g[16303];
assign g[32686] = b[13] & g[16303];
assign g[24496] = a[13] & g[16304];
assign g[32687] = b[13] & g[16304];
assign g[24497] = a[13] & g[16305];
assign g[32688] = b[13] & g[16305];
assign g[24498] = a[13] & g[16306];
assign g[32689] = b[13] & g[16306];
assign g[24499] = a[13] & g[16307];
assign g[32690] = b[13] & g[16307];
assign g[24500] = a[13] & g[16308];
assign g[32691] = b[13] & g[16308];
assign g[24501] = a[13] & g[16309];
assign g[32692] = b[13] & g[16309];
assign g[24502] = a[13] & g[16310];
assign g[32693] = b[13] & g[16310];
assign g[24503] = a[13] & g[16311];
assign g[32694] = b[13] & g[16311];
assign g[24504] = a[13] & g[16312];
assign g[32695] = b[13] & g[16312];
assign g[24505] = a[13] & g[16313];
assign g[32696] = b[13] & g[16313];
assign g[24506] = a[13] & g[16314];
assign g[32697] = b[13] & g[16314];
assign g[24507] = a[13] & g[16315];
assign g[32698] = b[13] & g[16315];
assign g[24508] = a[13] & g[16316];
assign g[32699] = b[13] & g[16316];
assign g[24509] = a[13] & g[16317];
assign g[32700] = b[13] & g[16317];
assign g[24510] = a[13] & g[16318];
assign g[32701] = b[13] & g[16318];
assign g[24511] = a[13] & g[16319];
assign g[32702] = b[13] & g[16319];
assign g[24512] = a[13] & g[16320];
assign g[32703] = b[13] & g[16320];
assign g[24513] = a[13] & g[16321];
assign g[32704] = b[13] & g[16321];
assign g[24514] = a[13] & g[16322];
assign g[32705] = b[13] & g[16322];
assign g[24515] = a[13] & g[16323];
assign g[32706] = b[13] & g[16323];
assign g[24516] = a[13] & g[16324];
assign g[32707] = b[13] & g[16324];
assign g[24517] = a[13] & g[16325];
assign g[32708] = b[13] & g[16325];
assign g[24518] = a[13] & g[16326];
assign g[32709] = b[13] & g[16326];
assign g[24519] = a[13] & g[16327];
assign g[32710] = b[13] & g[16327];
assign g[24520] = a[13] & g[16328];
assign g[32711] = b[13] & g[16328];
assign g[24521] = a[13] & g[16329];
assign g[32712] = b[13] & g[16329];
assign g[24522] = a[13] & g[16330];
assign g[32713] = b[13] & g[16330];
assign g[24523] = a[13] & g[16331];
assign g[32714] = b[13] & g[16331];
assign g[24524] = a[13] & g[16332];
assign g[32715] = b[13] & g[16332];
assign g[24525] = a[13] & g[16333];
assign g[32716] = b[13] & g[16333];
assign g[24526] = a[13] & g[16334];
assign g[32717] = b[13] & g[16334];
assign g[24527] = a[13] & g[16335];
assign g[32718] = b[13] & g[16335];
assign g[24528] = a[13] & g[16336];
assign g[32719] = b[13] & g[16336];
assign g[24529] = a[13] & g[16337];
assign g[32720] = b[13] & g[16337];
assign g[24530] = a[13] & g[16338];
assign g[32721] = b[13] & g[16338];
assign g[24531] = a[13] & g[16339];
assign g[32722] = b[13] & g[16339];
assign g[24532] = a[13] & g[16340];
assign g[32723] = b[13] & g[16340];
assign g[24533] = a[13] & g[16341];
assign g[32724] = b[13] & g[16341];
assign g[24534] = a[13] & g[16342];
assign g[32725] = b[13] & g[16342];
assign g[24535] = a[13] & g[16343];
assign g[32726] = b[13] & g[16343];
assign g[24536] = a[13] & g[16344];
assign g[32727] = b[13] & g[16344];
assign g[24537] = a[13] & g[16345];
assign g[32728] = b[13] & g[16345];
assign g[24538] = a[13] & g[16346];
assign g[32729] = b[13] & g[16346];
assign g[24539] = a[13] & g[16347];
assign g[32730] = b[13] & g[16347];
assign g[24540] = a[13] & g[16348];
assign g[32731] = b[13] & g[16348];
assign g[24541] = a[13] & g[16349];
assign g[32732] = b[13] & g[16349];
assign g[24542] = a[13] & g[16350];
assign g[32733] = b[13] & g[16350];
assign g[24543] = a[13] & g[16351];
assign g[32734] = b[13] & g[16351];
assign g[24544] = a[13] & g[16352];
assign g[32735] = b[13] & g[16352];
assign g[24545] = a[13] & g[16353];
assign g[32736] = b[13] & g[16353];
assign g[24546] = a[13] & g[16354];
assign g[32737] = b[13] & g[16354];
assign g[24547] = a[13] & g[16355];
assign g[32738] = b[13] & g[16355];
assign g[24548] = a[13] & g[16356];
assign g[32739] = b[13] & g[16356];
assign g[24549] = a[13] & g[16357];
assign g[32740] = b[13] & g[16357];
assign g[24550] = a[13] & g[16358];
assign g[32741] = b[13] & g[16358];
assign g[24551] = a[13] & g[16359];
assign g[32742] = b[13] & g[16359];
assign g[24552] = a[13] & g[16360];
assign g[32743] = b[13] & g[16360];
assign g[24553] = a[13] & g[16361];
assign g[32744] = b[13] & g[16361];
assign g[24554] = a[13] & g[16362];
assign g[32745] = b[13] & g[16362];
assign g[24555] = a[13] & g[16363];
assign g[32746] = b[13] & g[16363];
assign g[24556] = a[13] & g[16364];
assign g[32747] = b[13] & g[16364];
assign g[24557] = a[13] & g[16365];
assign g[32748] = b[13] & g[16365];
assign g[24558] = a[13] & g[16366];
assign g[32749] = b[13] & g[16366];
assign g[24559] = a[13] & g[16367];
assign g[32750] = b[13] & g[16367];
assign g[24560] = a[13] & g[16368];
assign g[32751] = b[13] & g[16368];
//Assigning outputs for input bit 15
assign g[32752] = a[14] & b[14];
assign g[32753] = a[14] & g[16369];
assign g[49136] = b[14] & g[16369];
assign g[32754] = a[14] & g[16370];
assign g[49137] = b[14] & g[16370];
assign g[32755] = a[14] & g[16371];
assign g[49138] = b[14] & g[16371];
assign g[32756] = a[14] & g[16372];
assign g[49139] = b[14] & g[16372];
assign g[32757] = a[14] & g[16373];
assign g[49140] = b[14] & g[16373];
assign g[32758] = a[14] & g[16374];
assign g[49141] = b[14] & g[16374];
assign g[32759] = a[14] & g[16375];
assign g[49142] = b[14] & g[16375];
assign g[32760] = a[14] & g[16376];
assign g[49143] = b[14] & g[16376];
assign g[32761] = a[14] & g[16377];
assign g[49144] = b[14] & g[16377];
assign g[32762] = a[14] & g[16378];
assign g[49145] = b[14] & g[16378];
assign g[32763] = a[14] & g[16379];
assign g[49146] = b[14] & g[16379];
assign g[32764] = a[14] & g[16380];
assign g[49147] = b[14] & g[16380];
assign g[32765] = a[14] & g[16381];
assign g[49148] = b[14] & g[16381];
assign g[32766] = a[14] & g[16382];
assign g[49149] = b[14] & g[16382];
assign g[32767] = a[14] & g[16383];
assign g[49150] = b[14] & g[16383];
assign g[32768] = a[14] & g[16384];
assign g[49151] = b[14] & g[16384];
assign g[32769] = a[14] & g[16385];
assign g[49152] = b[14] & g[16385];
assign g[32770] = a[14] & g[16386];
assign g[49153] = b[14] & g[16386];
assign g[32771] = a[14] & g[16387];
assign g[49154] = b[14] & g[16387];
assign g[32772] = a[14] & g[16388];
assign g[49155] = b[14] & g[16388];
assign g[32773] = a[14] & g[16389];
assign g[49156] = b[14] & g[16389];
assign g[32774] = a[14] & g[16390];
assign g[49157] = b[14] & g[16390];
assign g[32775] = a[14] & g[16391];
assign g[49158] = b[14] & g[16391];
assign g[32776] = a[14] & g[16392];
assign g[49159] = b[14] & g[16392];
assign g[32777] = a[14] & g[16393];
assign g[49160] = b[14] & g[16393];
assign g[32778] = a[14] & g[16394];
assign g[49161] = b[14] & g[16394];
assign g[32779] = a[14] & g[16395];
assign g[49162] = b[14] & g[16395];
assign g[32780] = a[14] & g[16396];
assign g[49163] = b[14] & g[16396];
assign g[32781] = a[14] & g[16397];
assign g[49164] = b[14] & g[16397];
assign g[32782] = a[14] & g[16398];
assign g[49165] = b[14] & g[16398];
assign g[32783] = a[14] & g[16399];
assign g[49166] = b[14] & g[16399];
assign g[32784] = a[14] & g[16400];
assign g[49167] = b[14] & g[16400];
assign g[32785] = a[14] & g[16401];
assign g[49168] = b[14] & g[16401];
assign g[32786] = a[14] & g[16402];
assign g[49169] = b[14] & g[16402];
assign g[32787] = a[14] & g[16403];
assign g[49170] = b[14] & g[16403];
assign g[32788] = a[14] & g[16404];
assign g[49171] = b[14] & g[16404];
assign g[32789] = a[14] & g[16405];
assign g[49172] = b[14] & g[16405];
assign g[32790] = a[14] & g[16406];
assign g[49173] = b[14] & g[16406];
assign g[32791] = a[14] & g[16407];
assign g[49174] = b[14] & g[16407];
assign g[32792] = a[14] & g[16408];
assign g[49175] = b[14] & g[16408];
assign g[32793] = a[14] & g[16409];
assign g[49176] = b[14] & g[16409];
assign g[32794] = a[14] & g[16410];
assign g[49177] = b[14] & g[16410];
assign g[32795] = a[14] & g[16411];
assign g[49178] = b[14] & g[16411];
assign g[32796] = a[14] & g[16412];
assign g[49179] = b[14] & g[16412];
assign g[32797] = a[14] & g[16413];
assign g[49180] = b[14] & g[16413];
assign g[32798] = a[14] & g[16414];
assign g[49181] = b[14] & g[16414];
assign g[32799] = a[14] & g[16415];
assign g[49182] = b[14] & g[16415];
assign g[32800] = a[14] & g[16416];
assign g[49183] = b[14] & g[16416];
assign g[32801] = a[14] & g[16417];
assign g[49184] = b[14] & g[16417];
assign g[32802] = a[14] & g[16418];
assign g[49185] = b[14] & g[16418];
assign g[32803] = a[14] & g[16419];
assign g[49186] = b[14] & g[16419];
assign g[32804] = a[14] & g[16420];
assign g[49187] = b[14] & g[16420];
assign g[32805] = a[14] & g[16421];
assign g[49188] = b[14] & g[16421];
assign g[32806] = a[14] & g[16422];
assign g[49189] = b[14] & g[16422];
assign g[32807] = a[14] & g[16423];
assign g[49190] = b[14] & g[16423];
assign g[32808] = a[14] & g[16424];
assign g[49191] = b[14] & g[16424];
assign g[32809] = a[14] & g[16425];
assign g[49192] = b[14] & g[16425];
assign g[32810] = a[14] & g[16426];
assign g[49193] = b[14] & g[16426];
assign g[32811] = a[14] & g[16427];
assign g[49194] = b[14] & g[16427];
assign g[32812] = a[14] & g[16428];
assign g[49195] = b[14] & g[16428];
assign g[32813] = a[14] & g[16429];
assign g[49196] = b[14] & g[16429];
assign g[32814] = a[14] & g[16430];
assign g[49197] = b[14] & g[16430];
assign g[32815] = a[14] & g[16431];
assign g[49198] = b[14] & g[16431];
assign g[32816] = a[14] & g[16432];
assign g[49199] = b[14] & g[16432];
assign g[32817] = a[14] & g[16433];
assign g[49200] = b[14] & g[16433];
assign g[32818] = a[14] & g[16434];
assign g[49201] = b[14] & g[16434];
assign g[32819] = a[14] & g[16435];
assign g[49202] = b[14] & g[16435];
assign g[32820] = a[14] & g[16436];
assign g[49203] = b[14] & g[16436];
assign g[32821] = a[14] & g[16437];
assign g[49204] = b[14] & g[16437];
assign g[32822] = a[14] & g[16438];
assign g[49205] = b[14] & g[16438];
assign g[32823] = a[14] & g[16439];
assign g[49206] = b[14] & g[16439];
assign g[32824] = a[14] & g[16440];
assign g[49207] = b[14] & g[16440];
assign g[32825] = a[14] & g[16441];
assign g[49208] = b[14] & g[16441];
assign g[32826] = a[14] & g[16442];
assign g[49209] = b[14] & g[16442];
assign g[32827] = a[14] & g[16443];
assign g[49210] = b[14] & g[16443];
assign g[32828] = a[14] & g[16444];
assign g[49211] = b[14] & g[16444];
assign g[32829] = a[14] & g[16445];
assign g[49212] = b[14] & g[16445];
assign g[32830] = a[14] & g[16446];
assign g[49213] = b[14] & g[16446];
assign g[32831] = a[14] & g[16447];
assign g[49214] = b[14] & g[16447];
assign g[32832] = a[14] & g[16448];
assign g[49215] = b[14] & g[16448];
assign g[32833] = a[14] & g[16449];
assign g[49216] = b[14] & g[16449];
assign g[32834] = a[14] & g[16450];
assign g[49217] = b[14] & g[16450];
assign g[32835] = a[14] & g[16451];
assign g[49218] = b[14] & g[16451];
assign g[32836] = a[14] & g[16452];
assign g[49219] = b[14] & g[16452];
assign g[32837] = a[14] & g[16453];
assign g[49220] = b[14] & g[16453];
assign g[32838] = a[14] & g[16454];
assign g[49221] = b[14] & g[16454];
assign g[32839] = a[14] & g[16455];
assign g[49222] = b[14] & g[16455];
assign g[32840] = a[14] & g[16456];
assign g[49223] = b[14] & g[16456];
assign g[32841] = a[14] & g[16457];
assign g[49224] = b[14] & g[16457];
assign g[32842] = a[14] & g[16458];
assign g[49225] = b[14] & g[16458];
assign g[32843] = a[14] & g[16459];
assign g[49226] = b[14] & g[16459];
assign g[32844] = a[14] & g[16460];
assign g[49227] = b[14] & g[16460];
assign g[32845] = a[14] & g[16461];
assign g[49228] = b[14] & g[16461];
assign g[32846] = a[14] & g[16462];
assign g[49229] = b[14] & g[16462];
assign g[32847] = a[14] & g[16463];
assign g[49230] = b[14] & g[16463];
assign g[32848] = a[14] & g[16464];
assign g[49231] = b[14] & g[16464];
assign g[32849] = a[14] & g[16465];
assign g[49232] = b[14] & g[16465];
assign g[32850] = a[14] & g[16466];
assign g[49233] = b[14] & g[16466];
assign g[32851] = a[14] & g[16467];
assign g[49234] = b[14] & g[16467];
assign g[32852] = a[14] & g[16468];
assign g[49235] = b[14] & g[16468];
assign g[32853] = a[14] & g[16469];
assign g[49236] = b[14] & g[16469];
assign g[32854] = a[14] & g[16470];
assign g[49237] = b[14] & g[16470];
assign g[32855] = a[14] & g[16471];
assign g[49238] = b[14] & g[16471];
assign g[32856] = a[14] & g[16472];
assign g[49239] = b[14] & g[16472];
assign g[32857] = a[14] & g[16473];
assign g[49240] = b[14] & g[16473];
assign g[32858] = a[14] & g[16474];
assign g[49241] = b[14] & g[16474];
assign g[32859] = a[14] & g[16475];
assign g[49242] = b[14] & g[16475];
assign g[32860] = a[14] & g[16476];
assign g[49243] = b[14] & g[16476];
assign g[32861] = a[14] & g[16477];
assign g[49244] = b[14] & g[16477];
assign g[32862] = a[14] & g[16478];
assign g[49245] = b[14] & g[16478];
assign g[32863] = a[14] & g[16479];
assign g[49246] = b[14] & g[16479];
assign g[32864] = a[14] & g[16480];
assign g[49247] = b[14] & g[16480];
assign g[32865] = a[14] & g[16481];
assign g[49248] = b[14] & g[16481];
assign g[32866] = a[14] & g[16482];
assign g[49249] = b[14] & g[16482];
assign g[32867] = a[14] & g[16483];
assign g[49250] = b[14] & g[16483];
assign g[32868] = a[14] & g[16484];
assign g[49251] = b[14] & g[16484];
assign g[32869] = a[14] & g[16485];
assign g[49252] = b[14] & g[16485];
assign g[32870] = a[14] & g[16486];
assign g[49253] = b[14] & g[16486];
assign g[32871] = a[14] & g[16487];
assign g[49254] = b[14] & g[16487];
assign g[32872] = a[14] & g[16488];
assign g[49255] = b[14] & g[16488];
assign g[32873] = a[14] & g[16489];
assign g[49256] = b[14] & g[16489];
assign g[32874] = a[14] & g[16490];
assign g[49257] = b[14] & g[16490];
assign g[32875] = a[14] & g[16491];
assign g[49258] = b[14] & g[16491];
assign g[32876] = a[14] & g[16492];
assign g[49259] = b[14] & g[16492];
assign g[32877] = a[14] & g[16493];
assign g[49260] = b[14] & g[16493];
assign g[32878] = a[14] & g[16494];
assign g[49261] = b[14] & g[16494];
assign g[32879] = a[14] & g[16495];
assign g[49262] = b[14] & g[16495];
assign g[32880] = a[14] & g[16496];
assign g[49263] = b[14] & g[16496];
assign g[32881] = a[14] & g[16497];
assign g[49264] = b[14] & g[16497];
assign g[32882] = a[14] & g[16498];
assign g[49265] = b[14] & g[16498];
assign g[32883] = a[14] & g[16499];
assign g[49266] = b[14] & g[16499];
assign g[32884] = a[14] & g[16500];
assign g[49267] = b[14] & g[16500];
assign g[32885] = a[14] & g[16501];
assign g[49268] = b[14] & g[16501];
assign g[32886] = a[14] & g[16502];
assign g[49269] = b[14] & g[16502];
assign g[32887] = a[14] & g[16503];
assign g[49270] = b[14] & g[16503];
assign g[32888] = a[14] & g[16504];
assign g[49271] = b[14] & g[16504];
assign g[32889] = a[14] & g[16505];
assign g[49272] = b[14] & g[16505];
assign g[32890] = a[14] & g[16506];
assign g[49273] = b[14] & g[16506];
assign g[32891] = a[14] & g[16507];
assign g[49274] = b[14] & g[16507];
assign g[32892] = a[14] & g[16508];
assign g[49275] = b[14] & g[16508];
assign g[32893] = a[14] & g[16509];
assign g[49276] = b[14] & g[16509];
assign g[32894] = a[14] & g[16510];
assign g[49277] = b[14] & g[16510];
assign g[32895] = a[14] & g[16511];
assign g[49278] = b[14] & g[16511];
assign g[32896] = a[14] & g[16512];
assign g[49279] = b[14] & g[16512];
assign g[32897] = a[14] & g[16513];
assign g[49280] = b[14] & g[16513];
assign g[32898] = a[14] & g[16514];
assign g[49281] = b[14] & g[16514];
assign g[32899] = a[14] & g[16515];
assign g[49282] = b[14] & g[16515];
assign g[32900] = a[14] & g[16516];
assign g[49283] = b[14] & g[16516];
assign g[32901] = a[14] & g[16517];
assign g[49284] = b[14] & g[16517];
assign g[32902] = a[14] & g[16518];
assign g[49285] = b[14] & g[16518];
assign g[32903] = a[14] & g[16519];
assign g[49286] = b[14] & g[16519];
assign g[32904] = a[14] & g[16520];
assign g[49287] = b[14] & g[16520];
assign g[32905] = a[14] & g[16521];
assign g[49288] = b[14] & g[16521];
assign g[32906] = a[14] & g[16522];
assign g[49289] = b[14] & g[16522];
assign g[32907] = a[14] & g[16523];
assign g[49290] = b[14] & g[16523];
assign g[32908] = a[14] & g[16524];
assign g[49291] = b[14] & g[16524];
assign g[32909] = a[14] & g[16525];
assign g[49292] = b[14] & g[16525];
assign g[32910] = a[14] & g[16526];
assign g[49293] = b[14] & g[16526];
assign g[32911] = a[14] & g[16527];
assign g[49294] = b[14] & g[16527];
assign g[32912] = a[14] & g[16528];
assign g[49295] = b[14] & g[16528];
assign g[32913] = a[14] & g[16529];
assign g[49296] = b[14] & g[16529];
assign g[32914] = a[14] & g[16530];
assign g[49297] = b[14] & g[16530];
assign g[32915] = a[14] & g[16531];
assign g[49298] = b[14] & g[16531];
assign g[32916] = a[14] & g[16532];
assign g[49299] = b[14] & g[16532];
assign g[32917] = a[14] & g[16533];
assign g[49300] = b[14] & g[16533];
assign g[32918] = a[14] & g[16534];
assign g[49301] = b[14] & g[16534];
assign g[32919] = a[14] & g[16535];
assign g[49302] = b[14] & g[16535];
assign g[32920] = a[14] & g[16536];
assign g[49303] = b[14] & g[16536];
assign g[32921] = a[14] & g[16537];
assign g[49304] = b[14] & g[16537];
assign g[32922] = a[14] & g[16538];
assign g[49305] = b[14] & g[16538];
assign g[32923] = a[14] & g[16539];
assign g[49306] = b[14] & g[16539];
assign g[32924] = a[14] & g[16540];
assign g[49307] = b[14] & g[16540];
assign g[32925] = a[14] & g[16541];
assign g[49308] = b[14] & g[16541];
assign g[32926] = a[14] & g[16542];
assign g[49309] = b[14] & g[16542];
assign g[32927] = a[14] & g[16543];
assign g[49310] = b[14] & g[16543];
assign g[32928] = a[14] & g[16544];
assign g[49311] = b[14] & g[16544];
assign g[32929] = a[14] & g[16545];
assign g[49312] = b[14] & g[16545];
assign g[32930] = a[14] & g[16546];
assign g[49313] = b[14] & g[16546];
assign g[32931] = a[14] & g[16547];
assign g[49314] = b[14] & g[16547];
assign g[32932] = a[14] & g[16548];
assign g[49315] = b[14] & g[16548];
assign g[32933] = a[14] & g[16549];
assign g[49316] = b[14] & g[16549];
assign g[32934] = a[14] & g[16550];
assign g[49317] = b[14] & g[16550];
assign g[32935] = a[14] & g[16551];
assign g[49318] = b[14] & g[16551];
assign g[32936] = a[14] & g[16552];
assign g[49319] = b[14] & g[16552];
assign g[32937] = a[14] & g[16553];
assign g[49320] = b[14] & g[16553];
assign g[32938] = a[14] & g[16554];
assign g[49321] = b[14] & g[16554];
assign g[32939] = a[14] & g[16555];
assign g[49322] = b[14] & g[16555];
assign g[32940] = a[14] & g[16556];
assign g[49323] = b[14] & g[16556];
assign g[32941] = a[14] & g[16557];
assign g[49324] = b[14] & g[16557];
assign g[32942] = a[14] & g[16558];
assign g[49325] = b[14] & g[16558];
assign g[32943] = a[14] & g[16559];
assign g[49326] = b[14] & g[16559];
assign g[32944] = a[14] & g[16560];
assign g[49327] = b[14] & g[16560];
assign g[32945] = a[14] & g[16561];
assign g[49328] = b[14] & g[16561];
assign g[32946] = a[14] & g[16562];
assign g[49329] = b[14] & g[16562];
assign g[32947] = a[14] & g[16563];
assign g[49330] = b[14] & g[16563];
assign g[32948] = a[14] & g[16564];
assign g[49331] = b[14] & g[16564];
assign g[32949] = a[14] & g[16565];
assign g[49332] = b[14] & g[16565];
assign g[32950] = a[14] & g[16566];
assign g[49333] = b[14] & g[16566];
assign g[32951] = a[14] & g[16567];
assign g[49334] = b[14] & g[16567];
assign g[32952] = a[14] & g[16568];
assign g[49335] = b[14] & g[16568];
assign g[32953] = a[14] & g[16569];
assign g[49336] = b[14] & g[16569];
assign g[32954] = a[14] & g[16570];
assign g[49337] = b[14] & g[16570];
assign g[32955] = a[14] & g[16571];
assign g[49338] = b[14] & g[16571];
assign g[32956] = a[14] & g[16572];
assign g[49339] = b[14] & g[16572];
assign g[32957] = a[14] & g[16573];
assign g[49340] = b[14] & g[16573];
assign g[32958] = a[14] & g[16574];
assign g[49341] = b[14] & g[16574];
assign g[32959] = a[14] & g[16575];
assign g[49342] = b[14] & g[16575];
assign g[32960] = a[14] & g[16576];
assign g[49343] = b[14] & g[16576];
assign g[32961] = a[14] & g[16577];
assign g[49344] = b[14] & g[16577];
assign g[32962] = a[14] & g[16578];
assign g[49345] = b[14] & g[16578];
assign g[32963] = a[14] & g[16579];
assign g[49346] = b[14] & g[16579];
assign g[32964] = a[14] & g[16580];
assign g[49347] = b[14] & g[16580];
assign g[32965] = a[14] & g[16581];
assign g[49348] = b[14] & g[16581];
assign g[32966] = a[14] & g[16582];
assign g[49349] = b[14] & g[16582];
assign g[32967] = a[14] & g[16583];
assign g[49350] = b[14] & g[16583];
assign g[32968] = a[14] & g[16584];
assign g[49351] = b[14] & g[16584];
assign g[32969] = a[14] & g[16585];
assign g[49352] = b[14] & g[16585];
assign g[32970] = a[14] & g[16586];
assign g[49353] = b[14] & g[16586];
assign g[32971] = a[14] & g[16587];
assign g[49354] = b[14] & g[16587];
assign g[32972] = a[14] & g[16588];
assign g[49355] = b[14] & g[16588];
assign g[32973] = a[14] & g[16589];
assign g[49356] = b[14] & g[16589];
assign g[32974] = a[14] & g[16590];
assign g[49357] = b[14] & g[16590];
assign g[32975] = a[14] & g[16591];
assign g[49358] = b[14] & g[16591];
assign g[32976] = a[14] & g[16592];
assign g[49359] = b[14] & g[16592];
assign g[32977] = a[14] & g[16593];
assign g[49360] = b[14] & g[16593];
assign g[32978] = a[14] & g[16594];
assign g[49361] = b[14] & g[16594];
assign g[32979] = a[14] & g[16595];
assign g[49362] = b[14] & g[16595];
assign g[32980] = a[14] & g[16596];
assign g[49363] = b[14] & g[16596];
assign g[32981] = a[14] & g[16597];
assign g[49364] = b[14] & g[16597];
assign g[32982] = a[14] & g[16598];
assign g[49365] = b[14] & g[16598];
assign g[32983] = a[14] & g[16599];
assign g[49366] = b[14] & g[16599];
assign g[32984] = a[14] & g[16600];
assign g[49367] = b[14] & g[16600];
assign g[32985] = a[14] & g[16601];
assign g[49368] = b[14] & g[16601];
assign g[32986] = a[14] & g[16602];
assign g[49369] = b[14] & g[16602];
assign g[32987] = a[14] & g[16603];
assign g[49370] = b[14] & g[16603];
assign g[32988] = a[14] & g[16604];
assign g[49371] = b[14] & g[16604];
assign g[32989] = a[14] & g[16605];
assign g[49372] = b[14] & g[16605];
assign g[32990] = a[14] & g[16606];
assign g[49373] = b[14] & g[16606];
assign g[32991] = a[14] & g[16607];
assign g[49374] = b[14] & g[16607];
assign g[32992] = a[14] & g[16608];
assign g[49375] = b[14] & g[16608];
assign g[32993] = a[14] & g[16609];
assign g[49376] = b[14] & g[16609];
assign g[32994] = a[14] & g[16610];
assign g[49377] = b[14] & g[16610];
assign g[32995] = a[14] & g[16611];
assign g[49378] = b[14] & g[16611];
assign g[32996] = a[14] & g[16612];
assign g[49379] = b[14] & g[16612];
assign g[32997] = a[14] & g[16613];
assign g[49380] = b[14] & g[16613];
assign g[32998] = a[14] & g[16614];
assign g[49381] = b[14] & g[16614];
assign g[32999] = a[14] & g[16615];
assign g[49382] = b[14] & g[16615];
assign g[33000] = a[14] & g[16616];
assign g[49383] = b[14] & g[16616];
assign g[33001] = a[14] & g[16617];
assign g[49384] = b[14] & g[16617];
assign g[33002] = a[14] & g[16618];
assign g[49385] = b[14] & g[16618];
assign g[33003] = a[14] & g[16619];
assign g[49386] = b[14] & g[16619];
assign g[33004] = a[14] & g[16620];
assign g[49387] = b[14] & g[16620];
assign g[33005] = a[14] & g[16621];
assign g[49388] = b[14] & g[16621];
assign g[33006] = a[14] & g[16622];
assign g[49389] = b[14] & g[16622];
assign g[33007] = a[14] & g[16623];
assign g[49390] = b[14] & g[16623];
assign g[33008] = a[14] & g[16624];
assign g[49391] = b[14] & g[16624];
assign g[33009] = a[14] & g[16625];
assign g[49392] = b[14] & g[16625];
assign g[33010] = a[14] & g[16626];
assign g[49393] = b[14] & g[16626];
assign g[33011] = a[14] & g[16627];
assign g[49394] = b[14] & g[16627];
assign g[33012] = a[14] & g[16628];
assign g[49395] = b[14] & g[16628];
assign g[33013] = a[14] & g[16629];
assign g[49396] = b[14] & g[16629];
assign g[33014] = a[14] & g[16630];
assign g[49397] = b[14] & g[16630];
assign g[33015] = a[14] & g[16631];
assign g[49398] = b[14] & g[16631];
assign g[33016] = a[14] & g[16632];
assign g[49399] = b[14] & g[16632];
assign g[33017] = a[14] & g[16633];
assign g[49400] = b[14] & g[16633];
assign g[33018] = a[14] & g[16634];
assign g[49401] = b[14] & g[16634];
assign g[33019] = a[14] & g[16635];
assign g[49402] = b[14] & g[16635];
assign g[33020] = a[14] & g[16636];
assign g[49403] = b[14] & g[16636];
assign g[33021] = a[14] & g[16637];
assign g[49404] = b[14] & g[16637];
assign g[33022] = a[14] & g[16638];
assign g[49405] = b[14] & g[16638];
assign g[33023] = a[14] & g[16639];
assign g[49406] = b[14] & g[16639];
assign g[33024] = a[14] & g[16640];
assign g[49407] = b[14] & g[16640];
assign g[33025] = a[14] & g[16641];
assign g[49408] = b[14] & g[16641];
assign g[33026] = a[14] & g[16642];
assign g[49409] = b[14] & g[16642];
assign g[33027] = a[14] & g[16643];
assign g[49410] = b[14] & g[16643];
assign g[33028] = a[14] & g[16644];
assign g[49411] = b[14] & g[16644];
assign g[33029] = a[14] & g[16645];
assign g[49412] = b[14] & g[16645];
assign g[33030] = a[14] & g[16646];
assign g[49413] = b[14] & g[16646];
assign g[33031] = a[14] & g[16647];
assign g[49414] = b[14] & g[16647];
assign g[33032] = a[14] & g[16648];
assign g[49415] = b[14] & g[16648];
assign g[33033] = a[14] & g[16649];
assign g[49416] = b[14] & g[16649];
assign g[33034] = a[14] & g[16650];
assign g[49417] = b[14] & g[16650];
assign g[33035] = a[14] & g[16651];
assign g[49418] = b[14] & g[16651];
assign g[33036] = a[14] & g[16652];
assign g[49419] = b[14] & g[16652];
assign g[33037] = a[14] & g[16653];
assign g[49420] = b[14] & g[16653];
assign g[33038] = a[14] & g[16654];
assign g[49421] = b[14] & g[16654];
assign g[33039] = a[14] & g[16655];
assign g[49422] = b[14] & g[16655];
assign g[33040] = a[14] & g[16656];
assign g[49423] = b[14] & g[16656];
assign g[33041] = a[14] & g[16657];
assign g[49424] = b[14] & g[16657];
assign g[33042] = a[14] & g[16658];
assign g[49425] = b[14] & g[16658];
assign g[33043] = a[14] & g[16659];
assign g[49426] = b[14] & g[16659];
assign g[33044] = a[14] & g[16660];
assign g[49427] = b[14] & g[16660];
assign g[33045] = a[14] & g[16661];
assign g[49428] = b[14] & g[16661];
assign g[33046] = a[14] & g[16662];
assign g[49429] = b[14] & g[16662];
assign g[33047] = a[14] & g[16663];
assign g[49430] = b[14] & g[16663];
assign g[33048] = a[14] & g[16664];
assign g[49431] = b[14] & g[16664];
assign g[33049] = a[14] & g[16665];
assign g[49432] = b[14] & g[16665];
assign g[33050] = a[14] & g[16666];
assign g[49433] = b[14] & g[16666];
assign g[33051] = a[14] & g[16667];
assign g[49434] = b[14] & g[16667];
assign g[33052] = a[14] & g[16668];
assign g[49435] = b[14] & g[16668];
assign g[33053] = a[14] & g[16669];
assign g[49436] = b[14] & g[16669];
assign g[33054] = a[14] & g[16670];
assign g[49437] = b[14] & g[16670];
assign g[33055] = a[14] & g[16671];
assign g[49438] = b[14] & g[16671];
assign g[33056] = a[14] & g[16672];
assign g[49439] = b[14] & g[16672];
assign g[33057] = a[14] & g[16673];
assign g[49440] = b[14] & g[16673];
assign g[33058] = a[14] & g[16674];
assign g[49441] = b[14] & g[16674];
assign g[33059] = a[14] & g[16675];
assign g[49442] = b[14] & g[16675];
assign g[33060] = a[14] & g[16676];
assign g[49443] = b[14] & g[16676];
assign g[33061] = a[14] & g[16677];
assign g[49444] = b[14] & g[16677];
assign g[33062] = a[14] & g[16678];
assign g[49445] = b[14] & g[16678];
assign g[33063] = a[14] & g[16679];
assign g[49446] = b[14] & g[16679];
assign g[33064] = a[14] & g[16680];
assign g[49447] = b[14] & g[16680];
assign g[33065] = a[14] & g[16681];
assign g[49448] = b[14] & g[16681];
assign g[33066] = a[14] & g[16682];
assign g[49449] = b[14] & g[16682];
assign g[33067] = a[14] & g[16683];
assign g[49450] = b[14] & g[16683];
assign g[33068] = a[14] & g[16684];
assign g[49451] = b[14] & g[16684];
assign g[33069] = a[14] & g[16685];
assign g[49452] = b[14] & g[16685];
assign g[33070] = a[14] & g[16686];
assign g[49453] = b[14] & g[16686];
assign g[33071] = a[14] & g[16687];
assign g[49454] = b[14] & g[16687];
assign g[33072] = a[14] & g[16688];
assign g[49455] = b[14] & g[16688];
assign g[33073] = a[14] & g[16689];
assign g[49456] = b[14] & g[16689];
assign g[33074] = a[14] & g[16690];
assign g[49457] = b[14] & g[16690];
assign g[33075] = a[14] & g[16691];
assign g[49458] = b[14] & g[16691];
assign g[33076] = a[14] & g[16692];
assign g[49459] = b[14] & g[16692];
assign g[33077] = a[14] & g[16693];
assign g[49460] = b[14] & g[16693];
assign g[33078] = a[14] & g[16694];
assign g[49461] = b[14] & g[16694];
assign g[33079] = a[14] & g[16695];
assign g[49462] = b[14] & g[16695];
assign g[33080] = a[14] & g[16696];
assign g[49463] = b[14] & g[16696];
assign g[33081] = a[14] & g[16697];
assign g[49464] = b[14] & g[16697];
assign g[33082] = a[14] & g[16698];
assign g[49465] = b[14] & g[16698];
assign g[33083] = a[14] & g[16699];
assign g[49466] = b[14] & g[16699];
assign g[33084] = a[14] & g[16700];
assign g[49467] = b[14] & g[16700];
assign g[33085] = a[14] & g[16701];
assign g[49468] = b[14] & g[16701];
assign g[33086] = a[14] & g[16702];
assign g[49469] = b[14] & g[16702];
assign g[33087] = a[14] & g[16703];
assign g[49470] = b[14] & g[16703];
assign g[33088] = a[14] & g[16704];
assign g[49471] = b[14] & g[16704];
assign g[33089] = a[14] & g[16705];
assign g[49472] = b[14] & g[16705];
assign g[33090] = a[14] & g[16706];
assign g[49473] = b[14] & g[16706];
assign g[33091] = a[14] & g[16707];
assign g[49474] = b[14] & g[16707];
assign g[33092] = a[14] & g[16708];
assign g[49475] = b[14] & g[16708];
assign g[33093] = a[14] & g[16709];
assign g[49476] = b[14] & g[16709];
assign g[33094] = a[14] & g[16710];
assign g[49477] = b[14] & g[16710];
assign g[33095] = a[14] & g[16711];
assign g[49478] = b[14] & g[16711];
assign g[33096] = a[14] & g[16712];
assign g[49479] = b[14] & g[16712];
assign g[33097] = a[14] & g[16713];
assign g[49480] = b[14] & g[16713];
assign g[33098] = a[14] & g[16714];
assign g[49481] = b[14] & g[16714];
assign g[33099] = a[14] & g[16715];
assign g[49482] = b[14] & g[16715];
assign g[33100] = a[14] & g[16716];
assign g[49483] = b[14] & g[16716];
assign g[33101] = a[14] & g[16717];
assign g[49484] = b[14] & g[16717];
assign g[33102] = a[14] & g[16718];
assign g[49485] = b[14] & g[16718];
assign g[33103] = a[14] & g[16719];
assign g[49486] = b[14] & g[16719];
assign g[33104] = a[14] & g[16720];
assign g[49487] = b[14] & g[16720];
assign g[33105] = a[14] & g[16721];
assign g[49488] = b[14] & g[16721];
assign g[33106] = a[14] & g[16722];
assign g[49489] = b[14] & g[16722];
assign g[33107] = a[14] & g[16723];
assign g[49490] = b[14] & g[16723];
assign g[33108] = a[14] & g[16724];
assign g[49491] = b[14] & g[16724];
assign g[33109] = a[14] & g[16725];
assign g[49492] = b[14] & g[16725];
assign g[33110] = a[14] & g[16726];
assign g[49493] = b[14] & g[16726];
assign g[33111] = a[14] & g[16727];
assign g[49494] = b[14] & g[16727];
assign g[33112] = a[14] & g[16728];
assign g[49495] = b[14] & g[16728];
assign g[33113] = a[14] & g[16729];
assign g[49496] = b[14] & g[16729];
assign g[33114] = a[14] & g[16730];
assign g[49497] = b[14] & g[16730];
assign g[33115] = a[14] & g[16731];
assign g[49498] = b[14] & g[16731];
assign g[33116] = a[14] & g[16732];
assign g[49499] = b[14] & g[16732];
assign g[33117] = a[14] & g[16733];
assign g[49500] = b[14] & g[16733];
assign g[33118] = a[14] & g[16734];
assign g[49501] = b[14] & g[16734];
assign g[33119] = a[14] & g[16735];
assign g[49502] = b[14] & g[16735];
assign g[33120] = a[14] & g[16736];
assign g[49503] = b[14] & g[16736];
assign g[33121] = a[14] & g[16737];
assign g[49504] = b[14] & g[16737];
assign g[33122] = a[14] & g[16738];
assign g[49505] = b[14] & g[16738];
assign g[33123] = a[14] & g[16739];
assign g[49506] = b[14] & g[16739];
assign g[33124] = a[14] & g[16740];
assign g[49507] = b[14] & g[16740];
assign g[33125] = a[14] & g[16741];
assign g[49508] = b[14] & g[16741];
assign g[33126] = a[14] & g[16742];
assign g[49509] = b[14] & g[16742];
assign g[33127] = a[14] & g[16743];
assign g[49510] = b[14] & g[16743];
assign g[33128] = a[14] & g[16744];
assign g[49511] = b[14] & g[16744];
assign g[33129] = a[14] & g[16745];
assign g[49512] = b[14] & g[16745];
assign g[33130] = a[14] & g[16746];
assign g[49513] = b[14] & g[16746];
assign g[33131] = a[14] & g[16747];
assign g[49514] = b[14] & g[16747];
assign g[33132] = a[14] & g[16748];
assign g[49515] = b[14] & g[16748];
assign g[33133] = a[14] & g[16749];
assign g[49516] = b[14] & g[16749];
assign g[33134] = a[14] & g[16750];
assign g[49517] = b[14] & g[16750];
assign g[33135] = a[14] & g[16751];
assign g[49518] = b[14] & g[16751];
assign g[33136] = a[14] & g[16752];
assign g[49519] = b[14] & g[16752];
assign g[33137] = a[14] & g[16753];
assign g[49520] = b[14] & g[16753];
assign g[33138] = a[14] & g[16754];
assign g[49521] = b[14] & g[16754];
assign g[33139] = a[14] & g[16755];
assign g[49522] = b[14] & g[16755];
assign g[33140] = a[14] & g[16756];
assign g[49523] = b[14] & g[16756];
assign g[33141] = a[14] & g[16757];
assign g[49524] = b[14] & g[16757];
assign g[33142] = a[14] & g[16758];
assign g[49525] = b[14] & g[16758];
assign g[33143] = a[14] & g[16759];
assign g[49526] = b[14] & g[16759];
assign g[33144] = a[14] & g[16760];
assign g[49527] = b[14] & g[16760];
assign g[33145] = a[14] & g[16761];
assign g[49528] = b[14] & g[16761];
assign g[33146] = a[14] & g[16762];
assign g[49529] = b[14] & g[16762];
assign g[33147] = a[14] & g[16763];
assign g[49530] = b[14] & g[16763];
assign g[33148] = a[14] & g[16764];
assign g[49531] = b[14] & g[16764];
assign g[33149] = a[14] & g[16765];
assign g[49532] = b[14] & g[16765];
assign g[33150] = a[14] & g[16766];
assign g[49533] = b[14] & g[16766];
assign g[33151] = a[14] & g[16767];
assign g[49534] = b[14] & g[16767];
assign g[33152] = a[14] & g[16768];
assign g[49535] = b[14] & g[16768];
assign g[33153] = a[14] & g[16769];
assign g[49536] = b[14] & g[16769];
assign g[33154] = a[14] & g[16770];
assign g[49537] = b[14] & g[16770];
assign g[33155] = a[14] & g[16771];
assign g[49538] = b[14] & g[16771];
assign g[33156] = a[14] & g[16772];
assign g[49539] = b[14] & g[16772];
assign g[33157] = a[14] & g[16773];
assign g[49540] = b[14] & g[16773];
assign g[33158] = a[14] & g[16774];
assign g[49541] = b[14] & g[16774];
assign g[33159] = a[14] & g[16775];
assign g[49542] = b[14] & g[16775];
assign g[33160] = a[14] & g[16776];
assign g[49543] = b[14] & g[16776];
assign g[33161] = a[14] & g[16777];
assign g[49544] = b[14] & g[16777];
assign g[33162] = a[14] & g[16778];
assign g[49545] = b[14] & g[16778];
assign g[33163] = a[14] & g[16779];
assign g[49546] = b[14] & g[16779];
assign g[33164] = a[14] & g[16780];
assign g[49547] = b[14] & g[16780];
assign g[33165] = a[14] & g[16781];
assign g[49548] = b[14] & g[16781];
assign g[33166] = a[14] & g[16782];
assign g[49549] = b[14] & g[16782];
assign g[33167] = a[14] & g[16783];
assign g[49550] = b[14] & g[16783];
assign g[33168] = a[14] & g[16784];
assign g[49551] = b[14] & g[16784];
assign g[33169] = a[14] & g[16785];
assign g[49552] = b[14] & g[16785];
assign g[33170] = a[14] & g[16786];
assign g[49553] = b[14] & g[16786];
assign g[33171] = a[14] & g[16787];
assign g[49554] = b[14] & g[16787];
assign g[33172] = a[14] & g[16788];
assign g[49555] = b[14] & g[16788];
assign g[33173] = a[14] & g[16789];
assign g[49556] = b[14] & g[16789];
assign g[33174] = a[14] & g[16790];
assign g[49557] = b[14] & g[16790];
assign g[33175] = a[14] & g[16791];
assign g[49558] = b[14] & g[16791];
assign g[33176] = a[14] & g[16792];
assign g[49559] = b[14] & g[16792];
assign g[33177] = a[14] & g[16793];
assign g[49560] = b[14] & g[16793];
assign g[33178] = a[14] & g[16794];
assign g[49561] = b[14] & g[16794];
assign g[33179] = a[14] & g[16795];
assign g[49562] = b[14] & g[16795];
assign g[33180] = a[14] & g[16796];
assign g[49563] = b[14] & g[16796];
assign g[33181] = a[14] & g[16797];
assign g[49564] = b[14] & g[16797];
assign g[33182] = a[14] & g[16798];
assign g[49565] = b[14] & g[16798];
assign g[33183] = a[14] & g[16799];
assign g[49566] = b[14] & g[16799];
assign g[33184] = a[14] & g[16800];
assign g[49567] = b[14] & g[16800];
assign g[33185] = a[14] & g[16801];
assign g[49568] = b[14] & g[16801];
assign g[33186] = a[14] & g[16802];
assign g[49569] = b[14] & g[16802];
assign g[33187] = a[14] & g[16803];
assign g[49570] = b[14] & g[16803];
assign g[33188] = a[14] & g[16804];
assign g[49571] = b[14] & g[16804];
assign g[33189] = a[14] & g[16805];
assign g[49572] = b[14] & g[16805];
assign g[33190] = a[14] & g[16806];
assign g[49573] = b[14] & g[16806];
assign g[33191] = a[14] & g[16807];
assign g[49574] = b[14] & g[16807];
assign g[33192] = a[14] & g[16808];
assign g[49575] = b[14] & g[16808];
assign g[33193] = a[14] & g[16809];
assign g[49576] = b[14] & g[16809];
assign g[33194] = a[14] & g[16810];
assign g[49577] = b[14] & g[16810];
assign g[33195] = a[14] & g[16811];
assign g[49578] = b[14] & g[16811];
assign g[33196] = a[14] & g[16812];
assign g[49579] = b[14] & g[16812];
assign g[33197] = a[14] & g[16813];
assign g[49580] = b[14] & g[16813];
assign g[33198] = a[14] & g[16814];
assign g[49581] = b[14] & g[16814];
assign g[33199] = a[14] & g[16815];
assign g[49582] = b[14] & g[16815];
assign g[33200] = a[14] & g[16816];
assign g[49583] = b[14] & g[16816];
assign g[33201] = a[14] & g[16817];
assign g[49584] = b[14] & g[16817];
assign g[33202] = a[14] & g[16818];
assign g[49585] = b[14] & g[16818];
assign g[33203] = a[14] & g[16819];
assign g[49586] = b[14] & g[16819];
assign g[33204] = a[14] & g[16820];
assign g[49587] = b[14] & g[16820];
assign g[33205] = a[14] & g[16821];
assign g[49588] = b[14] & g[16821];
assign g[33206] = a[14] & g[16822];
assign g[49589] = b[14] & g[16822];
assign g[33207] = a[14] & g[16823];
assign g[49590] = b[14] & g[16823];
assign g[33208] = a[14] & g[16824];
assign g[49591] = b[14] & g[16824];
assign g[33209] = a[14] & g[16825];
assign g[49592] = b[14] & g[16825];
assign g[33210] = a[14] & g[16826];
assign g[49593] = b[14] & g[16826];
assign g[33211] = a[14] & g[16827];
assign g[49594] = b[14] & g[16827];
assign g[33212] = a[14] & g[16828];
assign g[49595] = b[14] & g[16828];
assign g[33213] = a[14] & g[16829];
assign g[49596] = b[14] & g[16829];
assign g[33214] = a[14] & g[16830];
assign g[49597] = b[14] & g[16830];
assign g[33215] = a[14] & g[16831];
assign g[49598] = b[14] & g[16831];
assign g[33216] = a[14] & g[16832];
assign g[49599] = b[14] & g[16832];
assign g[33217] = a[14] & g[16833];
assign g[49600] = b[14] & g[16833];
assign g[33218] = a[14] & g[16834];
assign g[49601] = b[14] & g[16834];
assign g[33219] = a[14] & g[16835];
assign g[49602] = b[14] & g[16835];
assign g[33220] = a[14] & g[16836];
assign g[49603] = b[14] & g[16836];
assign g[33221] = a[14] & g[16837];
assign g[49604] = b[14] & g[16837];
assign g[33222] = a[14] & g[16838];
assign g[49605] = b[14] & g[16838];
assign g[33223] = a[14] & g[16839];
assign g[49606] = b[14] & g[16839];
assign g[33224] = a[14] & g[16840];
assign g[49607] = b[14] & g[16840];
assign g[33225] = a[14] & g[16841];
assign g[49608] = b[14] & g[16841];
assign g[33226] = a[14] & g[16842];
assign g[49609] = b[14] & g[16842];
assign g[33227] = a[14] & g[16843];
assign g[49610] = b[14] & g[16843];
assign g[33228] = a[14] & g[16844];
assign g[49611] = b[14] & g[16844];
assign g[33229] = a[14] & g[16845];
assign g[49612] = b[14] & g[16845];
assign g[33230] = a[14] & g[16846];
assign g[49613] = b[14] & g[16846];
assign g[33231] = a[14] & g[16847];
assign g[49614] = b[14] & g[16847];
assign g[33232] = a[14] & g[16848];
assign g[49615] = b[14] & g[16848];
assign g[33233] = a[14] & g[16849];
assign g[49616] = b[14] & g[16849];
assign g[33234] = a[14] & g[16850];
assign g[49617] = b[14] & g[16850];
assign g[33235] = a[14] & g[16851];
assign g[49618] = b[14] & g[16851];
assign g[33236] = a[14] & g[16852];
assign g[49619] = b[14] & g[16852];
assign g[33237] = a[14] & g[16853];
assign g[49620] = b[14] & g[16853];
assign g[33238] = a[14] & g[16854];
assign g[49621] = b[14] & g[16854];
assign g[33239] = a[14] & g[16855];
assign g[49622] = b[14] & g[16855];
assign g[33240] = a[14] & g[16856];
assign g[49623] = b[14] & g[16856];
assign g[33241] = a[14] & g[16857];
assign g[49624] = b[14] & g[16857];
assign g[33242] = a[14] & g[16858];
assign g[49625] = b[14] & g[16858];
assign g[33243] = a[14] & g[16859];
assign g[49626] = b[14] & g[16859];
assign g[33244] = a[14] & g[16860];
assign g[49627] = b[14] & g[16860];
assign g[33245] = a[14] & g[16861];
assign g[49628] = b[14] & g[16861];
assign g[33246] = a[14] & g[16862];
assign g[49629] = b[14] & g[16862];
assign g[33247] = a[14] & g[16863];
assign g[49630] = b[14] & g[16863];
assign g[33248] = a[14] & g[16864];
assign g[49631] = b[14] & g[16864];
assign g[33249] = a[14] & g[16865];
assign g[49632] = b[14] & g[16865];
assign g[33250] = a[14] & g[16866];
assign g[49633] = b[14] & g[16866];
assign g[33251] = a[14] & g[16867];
assign g[49634] = b[14] & g[16867];
assign g[33252] = a[14] & g[16868];
assign g[49635] = b[14] & g[16868];
assign g[33253] = a[14] & g[16869];
assign g[49636] = b[14] & g[16869];
assign g[33254] = a[14] & g[16870];
assign g[49637] = b[14] & g[16870];
assign g[33255] = a[14] & g[16871];
assign g[49638] = b[14] & g[16871];
assign g[33256] = a[14] & g[16872];
assign g[49639] = b[14] & g[16872];
assign g[33257] = a[14] & g[16873];
assign g[49640] = b[14] & g[16873];
assign g[33258] = a[14] & g[16874];
assign g[49641] = b[14] & g[16874];
assign g[33259] = a[14] & g[16875];
assign g[49642] = b[14] & g[16875];
assign g[33260] = a[14] & g[16876];
assign g[49643] = b[14] & g[16876];
assign g[33261] = a[14] & g[16877];
assign g[49644] = b[14] & g[16877];
assign g[33262] = a[14] & g[16878];
assign g[49645] = b[14] & g[16878];
assign g[33263] = a[14] & g[16879];
assign g[49646] = b[14] & g[16879];
assign g[33264] = a[14] & g[16880];
assign g[49647] = b[14] & g[16880];
assign g[33265] = a[14] & g[16881];
assign g[49648] = b[14] & g[16881];
assign g[33266] = a[14] & g[16882];
assign g[49649] = b[14] & g[16882];
assign g[33267] = a[14] & g[16883];
assign g[49650] = b[14] & g[16883];
assign g[33268] = a[14] & g[16884];
assign g[49651] = b[14] & g[16884];
assign g[33269] = a[14] & g[16885];
assign g[49652] = b[14] & g[16885];
assign g[33270] = a[14] & g[16886];
assign g[49653] = b[14] & g[16886];
assign g[33271] = a[14] & g[16887];
assign g[49654] = b[14] & g[16887];
assign g[33272] = a[14] & g[16888];
assign g[49655] = b[14] & g[16888];
assign g[33273] = a[14] & g[16889];
assign g[49656] = b[14] & g[16889];
assign g[33274] = a[14] & g[16890];
assign g[49657] = b[14] & g[16890];
assign g[33275] = a[14] & g[16891];
assign g[49658] = b[14] & g[16891];
assign g[33276] = a[14] & g[16892];
assign g[49659] = b[14] & g[16892];
assign g[33277] = a[14] & g[16893];
assign g[49660] = b[14] & g[16893];
assign g[33278] = a[14] & g[16894];
assign g[49661] = b[14] & g[16894];
assign g[33279] = a[14] & g[16895];
assign g[49662] = b[14] & g[16895];
assign g[33280] = a[14] & g[16896];
assign g[49663] = b[14] & g[16896];
assign g[33281] = a[14] & g[16897];
assign g[49664] = b[14] & g[16897];
assign g[33282] = a[14] & g[16898];
assign g[49665] = b[14] & g[16898];
assign g[33283] = a[14] & g[16899];
assign g[49666] = b[14] & g[16899];
assign g[33284] = a[14] & g[16900];
assign g[49667] = b[14] & g[16900];
assign g[33285] = a[14] & g[16901];
assign g[49668] = b[14] & g[16901];
assign g[33286] = a[14] & g[16902];
assign g[49669] = b[14] & g[16902];
assign g[33287] = a[14] & g[16903];
assign g[49670] = b[14] & g[16903];
assign g[33288] = a[14] & g[16904];
assign g[49671] = b[14] & g[16904];
assign g[33289] = a[14] & g[16905];
assign g[49672] = b[14] & g[16905];
assign g[33290] = a[14] & g[16906];
assign g[49673] = b[14] & g[16906];
assign g[33291] = a[14] & g[16907];
assign g[49674] = b[14] & g[16907];
assign g[33292] = a[14] & g[16908];
assign g[49675] = b[14] & g[16908];
assign g[33293] = a[14] & g[16909];
assign g[49676] = b[14] & g[16909];
assign g[33294] = a[14] & g[16910];
assign g[49677] = b[14] & g[16910];
assign g[33295] = a[14] & g[16911];
assign g[49678] = b[14] & g[16911];
assign g[33296] = a[14] & g[16912];
assign g[49679] = b[14] & g[16912];
assign g[33297] = a[14] & g[16913];
assign g[49680] = b[14] & g[16913];
assign g[33298] = a[14] & g[16914];
assign g[49681] = b[14] & g[16914];
assign g[33299] = a[14] & g[16915];
assign g[49682] = b[14] & g[16915];
assign g[33300] = a[14] & g[16916];
assign g[49683] = b[14] & g[16916];
assign g[33301] = a[14] & g[16917];
assign g[49684] = b[14] & g[16917];
assign g[33302] = a[14] & g[16918];
assign g[49685] = b[14] & g[16918];
assign g[33303] = a[14] & g[16919];
assign g[49686] = b[14] & g[16919];
assign g[33304] = a[14] & g[16920];
assign g[49687] = b[14] & g[16920];
assign g[33305] = a[14] & g[16921];
assign g[49688] = b[14] & g[16921];
assign g[33306] = a[14] & g[16922];
assign g[49689] = b[14] & g[16922];
assign g[33307] = a[14] & g[16923];
assign g[49690] = b[14] & g[16923];
assign g[33308] = a[14] & g[16924];
assign g[49691] = b[14] & g[16924];
assign g[33309] = a[14] & g[16925];
assign g[49692] = b[14] & g[16925];
assign g[33310] = a[14] & g[16926];
assign g[49693] = b[14] & g[16926];
assign g[33311] = a[14] & g[16927];
assign g[49694] = b[14] & g[16927];
assign g[33312] = a[14] & g[16928];
assign g[49695] = b[14] & g[16928];
assign g[33313] = a[14] & g[16929];
assign g[49696] = b[14] & g[16929];
assign g[33314] = a[14] & g[16930];
assign g[49697] = b[14] & g[16930];
assign g[33315] = a[14] & g[16931];
assign g[49698] = b[14] & g[16931];
assign g[33316] = a[14] & g[16932];
assign g[49699] = b[14] & g[16932];
assign g[33317] = a[14] & g[16933];
assign g[49700] = b[14] & g[16933];
assign g[33318] = a[14] & g[16934];
assign g[49701] = b[14] & g[16934];
assign g[33319] = a[14] & g[16935];
assign g[49702] = b[14] & g[16935];
assign g[33320] = a[14] & g[16936];
assign g[49703] = b[14] & g[16936];
assign g[33321] = a[14] & g[16937];
assign g[49704] = b[14] & g[16937];
assign g[33322] = a[14] & g[16938];
assign g[49705] = b[14] & g[16938];
assign g[33323] = a[14] & g[16939];
assign g[49706] = b[14] & g[16939];
assign g[33324] = a[14] & g[16940];
assign g[49707] = b[14] & g[16940];
assign g[33325] = a[14] & g[16941];
assign g[49708] = b[14] & g[16941];
assign g[33326] = a[14] & g[16942];
assign g[49709] = b[14] & g[16942];
assign g[33327] = a[14] & g[16943];
assign g[49710] = b[14] & g[16943];
assign g[33328] = a[14] & g[16944];
assign g[49711] = b[14] & g[16944];
assign g[33329] = a[14] & g[16945];
assign g[49712] = b[14] & g[16945];
assign g[33330] = a[14] & g[16946];
assign g[49713] = b[14] & g[16946];
assign g[33331] = a[14] & g[16947];
assign g[49714] = b[14] & g[16947];
assign g[33332] = a[14] & g[16948];
assign g[49715] = b[14] & g[16948];
assign g[33333] = a[14] & g[16949];
assign g[49716] = b[14] & g[16949];
assign g[33334] = a[14] & g[16950];
assign g[49717] = b[14] & g[16950];
assign g[33335] = a[14] & g[16951];
assign g[49718] = b[14] & g[16951];
assign g[33336] = a[14] & g[16952];
assign g[49719] = b[14] & g[16952];
assign g[33337] = a[14] & g[16953];
assign g[49720] = b[14] & g[16953];
assign g[33338] = a[14] & g[16954];
assign g[49721] = b[14] & g[16954];
assign g[33339] = a[14] & g[16955];
assign g[49722] = b[14] & g[16955];
assign g[33340] = a[14] & g[16956];
assign g[49723] = b[14] & g[16956];
assign g[33341] = a[14] & g[16957];
assign g[49724] = b[14] & g[16957];
assign g[33342] = a[14] & g[16958];
assign g[49725] = b[14] & g[16958];
assign g[33343] = a[14] & g[16959];
assign g[49726] = b[14] & g[16959];
assign g[33344] = a[14] & g[16960];
assign g[49727] = b[14] & g[16960];
assign g[33345] = a[14] & g[16961];
assign g[49728] = b[14] & g[16961];
assign g[33346] = a[14] & g[16962];
assign g[49729] = b[14] & g[16962];
assign g[33347] = a[14] & g[16963];
assign g[49730] = b[14] & g[16963];
assign g[33348] = a[14] & g[16964];
assign g[49731] = b[14] & g[16964];
assign g[33349] = a[14] & g[16965];
assign g[49732] = b[14] & g[16965];
assign g[33350] = a[14] & g[16966];
assign g[49733] = b[14] & g[16966];
assign g[33351] = a[14] & g[16967];
assign g[49734] = b[14] & g[16967];
assign g[33352] = a[14] & g[16968];
assign g[49735] = b[14] & g[16968];
assign g[33353] = a[14] & g[16969];
assign g[49736] = b[14] & g[16969];
assign g[33354] = a[14] & g[16970];
assign g[49737] = b[14] & g[16970];
assign g[33355] = a[14] & g[16971];
assign g[49738] = b[14] & g[16971];
assign g[33356] = a[14] & g[16972];
assign g[49739] = b[14] & g[16972];
assign g[33357] = a[14] & g[16973];
assign g[49740] = b[14] & g[16973];
assign g[33358] = a[14] & g[16974];
assign g[49741] = b[14] & g[16974];
assign g[33359] = a[14] & g[16975];
assign g[49742] = b[14] & g[16975];
assign g[33360] = a[14] & g[16976];
assign g[49743] = b[14] & g[16976];
assign g[33361] = a[14] & g[16977];
assign g[49744] = b[14] & g[16977];
assign g[33362] = a[14] & g[16978];
assign g[49745] = b[14] & g[16978];
assign g[33363] = a[14] & g[16979];
assign g[49746] = b[14] & g[16979];
assign g[33364] = a[14] & g[16980];
assign g[49747] = b[14] & g[16980];
assign g[33365] = a[14] & g[16981];
assign g[49748] = b[14] & g[16981];
assign g[33366] = a[14] & g[16982];
assign g[49749] = b[14] & g[16982];
assign g[33367] = a[14] & g[16983];
assign g[49750] = b[14] & g[16983];
assign g[33368] = a[14] & g[16984];
assign g[49751] = b[14] & g[16984];
assign g[33369] = a[14] & g[16985];
assign g[49752] = b[14] & g[16985];
assign g[33370] = a[14] & g[16986];
assign g[49753] = b[14] & g[16986];
assign g[33371] = a[14] & g[16987];
assign g[49754] = b[14] & g[16987];
assign g[33372] = a[14] & g[16988];
assign g[49755] = b[14] & g[16988];
assign g[33373] = a[14] & g[16989];
assign g[49756] = b[14] & g[16989];
assign g[33374] = a[14] & g[16990];
assign g[49757] = b[14] & g[16990];
assign g[33375] = a[14] & g[16991];
assign g[49758] = b[14] & g[16991];
assign g[33376] = a[14] & g[16992];
assign g[49759] = b[14] & g[16992];
assign g[33377] = a[14] & g[16993];
assign g[49760] = b[14] & g[16993];
assign g[33378] = a[14] & g[16994];
assign g[49761] = b[14] & g[16994];
assign g[33379] = a[14] & g[16995];
assign g[49762] = b[14] & g[16995];
assign g[33380] = a[14] & g[16996];
assign g[49763] = b[14] & g[16996];
assign g[33381] = a[14] & g[16997];
assign g[49764] = b[14] & g[16997];
assign g[33382] = a[14] & g[16998];
assign g[49765] = b[14] & g[16998];
assign g[33383] = a[14] & g[16999];
assign g[49766] = b[14] & g[16999];
assign g[33384] = a[14] & g[17000];
assign g[49767] = b[14] & g[17000];
assign g[33385] = a[14] & g[17001];
assign g[49768] = b[14] & g[17001];
assign g[33386] = a[14] & g[17002];
assign g[49769] = b[14] & g[17002];
assign g[33387] = a[14] & g[17003];
assign g[49770] = b[14] & g[17003];
assign g[33388] = a[14] & g[17004];
assign g[49771] = b[14] & g[17004];
assign g[33389] = a[14] & g[17005];
assign g[49772] = b[14] & g[17005];
assign g[33390] = a[14] & g[17006];
assign g[49773] = b[14] & g[17006];
assign g[33391] = a[14] & g[17007];
assign g[49774] = b[14] & g[17007];
assign g[33392] = a[14] & g[17008];
assign g[49775] = b[14] & g[17008];
assign g[33393] = a[14] & g[17009];
assign g[49776] = b[14] & g[17009];
assign g[33394] = a[14] & g[17010];
assign g[49777] = b[14] & g[17010];
assign g[33395] = a[14] & g[17011];
assign g[49778] = b[14] & g[17011];
assign g[33396] = a[14] & g[17012];
assign g[49779] = b[14] & g[17012];
assign g[33397] = a[14] & g[17013];
assign g[49780] = b[14] & g[17013];
assign g[33398] = a[14] & g[17014];
assign g[49781] = b[14] & g[17014];
assign g[33399] = a[14] & g[17015];
assign g[49782] = b[14] & g[17015];
assign g[33400] = a[14] & g[17016];
assign g[49783] = b[14] & g[17016];
assign g[33401] = a[14] & g[17017];
assign g[49784] = b[14] & g[17017];
assign g[33402] = a[14] & g[17018];
assign g[49785] = b[14] & g[17018];
assign g[33403] = a[14] & g[17019];
assign g[49786] = b[14] & g[17019];
assign g[33404] = a[14] & g[17020];
assign g[49787] = b[14] & g[17020];
assign g[33405] = a[14] & g[17021];
assign g[49788] = b[14] & g[17021];
assign g[33406] = a[14] & g[17022];
assign g[49789] = b[14] & g[17022];
assign g[33407] = a[14] & g[17023];
assign g[49790] = b[14] & g[17023];
assign g[33408] = a[14] & g[17024];
assign g[49791] = b[14] & g[17024];
assign g[33409] = a[14] & g[17025];
assign g[49792] = b[14] & g[17025];
assign g[33410] = a[14] & g[17026];
assign g[49793] = b[14] & g[17026];
assign g[33411] = a[14] & g[17027];
assign g[49794] = b[14] & g[17027];
assign g[33412] = a[14] & g[17028];
assign g[49795] = b[14] & g[17028];
assign g[33413] = a[14] & g[17029];
assign g[49796] = b[14] & g[17029];
assign g[33414] = a[14] & g[17030];
assign g[49797] = b[14] & g[17030];
assign g[33415] = a[14] & g[17031];
assign g[49798] = b[14] & g[17031];
assign g[33416] = a[14] & g[17032];
assign g[49799] = b[14] & g[17032];
assign g[33417] = a[14] & g[17033];
assign g[49800] = b[14] & g[17033];
assign g[33418] = a[14] & g[17034];
assign g[49801] = b[14] & g[17034];
assign g[33419] = a[14] & g[17035];
assign g[49802] = b[14] & g[17035];
assign g[33420] = a[14] & g[17036];
assign g[49803] = b[14] & g[17036];
assign g[33421] = a[14] & g[17037];
assign g[49804] = b[14] & g[17037];
assign g[33422] = a[14] & g[17038];
assign g[49805] = b[14] & g[17038];
assign g[33423] = a[14] & g[17039];
assign g[49806] = b[14] & g[17039];
assign g[33424] = a[14] & g[17040];
assign g[49807] = b[14] & g[17040];
assign g[33425] = a[14] & g[17041];
assign g[49808] = b[14] & g[17041];
assign g[33426] = a[14] & g[17042];
assign g[49809] = b[14] & g[17042];
assign g[33427] = a[14] & g[17043];
assign g[49810] = b[14] & g[17043];
assign g[33428] = a[14] & g[17044];
assign g[49811] = b[14] & g[17044];
assign g[33429] = a[14] & g[17045];
assign g[49812] = b[14] & g[17045];
assign g[33430] = a[14] & g[17046];
assign g[49813] = b[14] & g[17046];
assign g[33431] = a[14] & g[17047];
assign g[49814] = b[14] & g[17047];
assign g[33432] = a[14] & g[17048];
assign g[49815] = b[14] & g[17048];
assign g[33433] = a[14] & g[17049];
assign g[49816] = b[14] & g[17049];
assign g[33434] = a[14] & g[17050];
assign g[49817] = b[14] & g[17050];
assign g[33435] = a[14] & g[17051];
assign g[49818] = b[14] & g[17051];
assign g[33436] = a[14] & g[17052];
assign g[49819] = b[14] & g[17052];
assign g[33437] = a[14] & g[17053];
assign g[49820] = b[14] & g[17053];
assign g[33438] = a[14] & g[17054];
assign g[49821] = b[14] & g[17054];
assign g[33439] = a[14] & g[17055];
assign g[49822] = b[14] & g[17055];
assign g[33440] = a[14] & g[17056];
assign g[49823] = b[14] & g[17056];
assign g[33441] = a[14] & g[17057];
assign g[49824] = b[14] & g[17057];
assign g[33442] = a[14] & g[17058];
assign g[49825] = b[14] & g[17058];
assign g[33443] = a[14] & g[17059];
assign g[49826] = b[14] & g[17059];
assign g[33444] = a[14] & g[17060];
assign g[49827] = b[14] & g[17060];
assign g[33445] = a[14] & g[17061];
assign g[49828] = b[14] & g[17061];
assign g[33446] = a[14] & g[17062];
assign g[49829] = b[14] & g[17062];
assign g[33447] = a[14] & g[17063];
assign g[49830] = b[14] & g[17063];
assign g[33448] = a[14] & g[17064];
assign g[49831] = b[14] & g[17064];
assign g[33449] = a[14] & g[17065];
assign g[49832] = b[14] & g[17065];
assign g[33450] = a[14] & g[17066];
assign g[49833] = b[14] & g[17066];
assign g[33451] = a[14] & g[17067];
assign g[49834] = b[14] & g[17067];
assign g[33452] = a[14] & g[17068];
assign g[49835] = b[14] & g[17068];
assign g[33453] = a[14] & g[17069];
assign g[49836] = b[14] & g[17069];
assign g[33454] = a[14] & g[17070];
assign g[49837] = b[14] & g[17070];
assign g[33455] = a[14] & g[17071];
assign g[49838] = b[14] & g[17071];
assign g[33456] = a[14] & g[17072];
assign g[49839] = b[14] & g[17072];
assign g[33457] = a[14] & g[17073];
assign g[49840] = b[14] & g[17073];
assign g[33458] = a[14] & g[17074];
assign g[49841] = b[14] & g[17074];
assign g[33459] = a[14] & g[17075];
assign g[49842] = b[14] & g[17075];
assign g[33460] = a[14] & g[17076];
assign g[49843] = b[14] & g[17076];
assign g[33461] = a[14] & g[17077];
assign g[49844] = b[14] & g[17077];
assign g[33462] = a[14] & g[17078];
assign g[49845] = b[14] & g[17078];
assign g[33463] = a[14] & g[17079];
assign g[49846] = b[14] & g[17079];
assign g[33464] = a[14] & g[17080];
assign g[49847] = b[14] & g[17080];
assign g[33465] = a[14] & g[17081];
assign g[49848] = b[14] & g[17081];
assign g[33466] = a[14] & g[17082];
assign g[49849] = b[14] & g[17082];
assign g[33467] = a[14] & g[17083];
assign g[49850] = b[14] & g[17083];
assign g[33468] = a[14] & g[17084];
assign g[49851] = b[14] & g[17084];
assign g[33469] = a[14] & g[17085];
assign g[49852] = b[14] & g[17085];
assign g[33470] = a[14] & g[17086];
assign g[49853] = b[14] & g[17086];
assign g[33471] = a[14] & g[17087];
assign g[49854] = b[14] & g[17087];
assign g[33472] = a[14] & g[17088];
assign g[49855] = b[14] & g[17088];
assign g[33473] = a[14] & g[17089];
assign g[49856] = b[14] & g[17089];
assign g[33474] = a[14] & g[17090];
assign g[49857] = b[14] & g[17090];
assign g[33475] = a[14] & g[17091];
assign g[49858] = b[14] & g[17091];
assign g[33476] = a[14] & g[17092];
assign g[49859] = b[14] & g[17092];
assign g[33477] = a[14] & g[17093];
assign g[49860] = b[14] & g[17093];
assign g[33478] = a[14] & g[17094];
assign g[49861] = b[14] & g[17094];
assign g[33479] = a[14] & g[17095];
assign g[49862] = b[14] & g[17095];
assign g[33480] = a[14] & g[17096];
assign g[49863] = b[14] & g[17096];
assign g[33481] = a[14] & g[17097];
assign g[49864] = b[14] & g[17097];
assign g[33482] = a[14] & g[17098];
assign g[49865] = b[14] & g[17098];
assign g[33483] = a[14] & g[17099];
assign g[49866] = b[14] & g[17099];
assign g[33484] = a[14] & g[17100];
assign g[49867] = b[14] & g[17100];
assign g[33485] = a[14] & g[17101];
assign g[49868] = b[14] & g[17101];
assign g[33486] = a[14] & g[17102];
assign g[49869] = b[14] & g[17102];
assign g[33487] = a[14] & g[17103];
assign g[49870] = b[14] & g[17103];
assign g[33488] = a[14] & g[17104];
assign g[49871] = b[14] & g[17104];
assign g[33489] = a[14] & g[17105];
assign g[49872] = b[14] & g[17105];
assign g[33490] = a[14] & g[17106];
assign g[49873] = b[14] & g[17106];
assign g[33491] = a[14] & g[17107];
assign g[49874] = b[14] & g[17107];
assign g[33492] = a[14] & g[17108];
assign g[49875] = b[14] & g[17108];
assign g[33493] = a[14] & g[17109];
assign g[49876] = b[14] & g[17109];
assign g[33494] = a[14] & g[17110];
assign g[49877] = b[14] & g[17110];
assign g[33495] = a[14] & g[17111];
assign g[49878] = b[14] & g[17111];
assign g[33496] = a[14] & g[17112];
assign g[49879] = b[14] & g[17112];
assign g[33497] = a[14] & g[17113];
assign g[49880] = b[14] & g[17113];
assign g[33498] = a[14] & g[17114];
assign g[49881] = b[14] & g[17114];
assign g[33499] = a[14] & g[17115];
assign g[49882] = b[14] & g[17115];
assign g[33500] = a[14] & g[17116];
assign g[49883] = b[14] & g[17116];
assign g[33501] = a[14] & g[17117];
assign g[49884] = b[14] & g[17117];
assign g[33502] = a[14] & g[17118];
assign g[49885] = b[14] & g[17118];
assign g[33503] = a[14] & g[17119];
assign g[49886] = b[14] & g[17119];
assign g[33504] = a[14] & g[17120];
assign g[49887] = b[14] & g[17120];
assign g[33505] = a[14] & g[17121];
assign g[49888] = b[14] & g[17121];
assign g[33506] = a[14] & g[17122];
assign g[49889] = b[14] & g[17122];
assign g[33507] = a[14] & g[17123];
assign g[49890] = b[14] & g[17123];
assign g[33508] = a[14] & g[17124];
assign g[49891] = b[14] & g[17124];
assign g[33509] = a[14] & g[17125];
assign g[49892] = b[14] & g[17125];
assign g[33510] = a[14] & g[17126];
assign g[49893] = b[14] & g[17126];
assign g[33511] = a[14] & g[17127];
assign g[49894] = b[14] & g[17127];
assign g[33512] = a[14] & g[17128];
assign g[49895] = b[14] & g[17128];
assign g[33513] = a[14] & g[17129];
assign g[49896] = b[14] & g[17129];
assign g[33514] = a[14] & g[17130];
assign g[49897] = b[14] & g[17130];
assign g[33515] = a[14] & g[17131];
assign g[49898] = b[14] & g[17131];
assign g[33516] = a[14] & g[17132];
assign g[49899] = b[14] & g[17132];
assign g[33517] = a[14] & g[17133];
assign g[49900] = b[14] & g[17133];
assign g[33518] = a[14] & g[17134];
assign g[49901] = b[14] & g[17134];
assign g[33519] = a[14] & g[17135];
assign g[49902] = b[14] & g[17135];
assign g[33520] = a[14] & g[17136];
assign g[49903] = b[14] & g[17136];
assign g[33521] = a[14] & g[17137];
assign g[49904] = b[14] & g[17137];
assign g[33522] = a[14] & g[17138];
assign g[49905] = b[14] & g[17138];
assign g[33523] = a[14] & g[17139];
assign g[49906] = b[14] & g[17139];
assign g[33524] = a[14] & g[17140];
assign g[49907] = b[14] & g[17140];
assign g[33525] = a[14] & g[17141];
assign g[49908] = b[14] & g[17141];
assign g[33526] = a[14] & g[17142];
assign g[49909] = b[14] & g[17142];
assign g[33527] = a[14] & g[17143];
assign g[49910] = b[14] & g[17143];
assign g[33528] = a[14] & g[17144];
assign g[49911] = b[14] & g[17144];
assign g[33529] = a[14] & g[17145];
assign g[49912] = b[14] & g[17145];
assign g[33530] = a[14] & g[17146];
assign g[49913] = b[14] & g[17146];
assign g[33531] = a[14] & g[17147];
assign g[49914] = b[14] & g[17147];
assign g[33532] = a[14] & g[17148];
assign g[49915] = b[14] & g[17148];
assign g[33533] = a[14] & g[17149];
assign g[49916] = b[14] & g[17149];
assign g[33534] = a[14] & g[17150];
assign g[49917] = b[14] & g[17150];
assign g[33535] = a[14] & g[17151];
assign g[49918] = b[14] & g[17151];
assign g[33536] = a[14] & g[17152];
assign g[49919] = b[14] & g[17152];
assign g[33537] = a[14] & g[17153];
assign g[49920] = b[14] & g[17153];
assign g[33538] = a[14] & g[17154];
assign g[49921] = b[14] & g[17154];
assign g[33539] = a[14] & g[17155];
assign g[49922] = b[14] & g[17155];
assign g[33540] = a[14] & g[17156];
assign g[49923] = b[14] & g[17156];
assign g[33541] = a[14] & g[17157];
assign g[49924] = b[14] & g[17157];
assign g[33542] = a[14] & g[17158];
assign g[49925] = b[14] & g[17158];
assign g[33543] = a[14] & g[17159];
assign g[49926] = b[14] & g[17159];
assign g[33544] = a[14] & g[17160];
assign g[49927] = b[14] & g[17160];
assign g[33545] = a[14] & g[17161];
assign g[49928] = b[14] & g[17161];
assign g[33546] = a[14] & g[17162];
assign g[49929] = b[14] & g[17162];
assign g[33547] = a[14] & g[17163];
assign g[49930] = b[14] & g[17163];
assign g[33548] = a[14] & g[17164];
assign g[49931] = b[14] & g[17164];
assign g[33549] = a[14] & g[17165];
assign g[49932] = b[14] & g[17165];
assign g[33550] = a[14] & g[17166];
assign g[49933] = b[14] & g[17166];
assign g[33551] = a[14] & g[17167];
assign g[49934] = b[14] & g[17167];
assign g[33552] = a[14] & g[17168];
assign g[49935] = b[14] & g[17168];
assign g[33553] = a[14] & g[17169];
assign g[49936] = b[14] & g[17169];
assign g[33554] = a[14] & g[17170];
assign g[49937] = b[14] & g[17170];
assign g[33555] = a[14] & g[17171];
assign g[49938] = b[14] & g[17171];
assign g[33556] = a[14] & g[17172];
assign g[49939] = b[14] & g[17172];
assign g[33557] = a[14] & g[17173];
assign g[49940] = b[14] & g[17173];
assign g[33558] = a[14] & g[17174];
assign g[49941] = b[14] & g[17174];
assign g[33559] = a[14] & g[17175];
assign g[49942] = b[14] & g[17175];
assign g[33560] = a[14] & g[17176];
assign g[49943] = b[14] & g[17176];
assign g[33561] = a[14] & g[17177];
assign g[49944] = b[14] & g[17177];
assign g[33562] = a[14] & g[17178];
assign g[49945] = b[14] & g[17178];
assign g[33563] = a[14] & g[17179];
assign g[49946] = b[14] & g[17179];
assign g[33564] = a[14] & g[17180];
assign g[49947] = b[14] & g[17180];
assign g[33565] = a[14] & g[17181];
assign g[49948] = b[14] & g[17181];
assign g[33566] = a[14] & g[17182];
assign g[49949] = b[14] & g[17182];
assign g[33567] = a[14] & g[17183];
assign g[49950] = b[14] & g[17183];
assign g[33568] = a[14] & g[17184];
assign g[49951] = b[14] & g[17184];
assign g[33569] = a[14] & g[17185];
assign g[49952] = b[14] & g[17185];
assign g[33570] = a[14] & g[17186];
assign g[49953] = b[14] & g[17186];
assign g[33571] = a[14] & g[17187];
assign g[49954] = b[14] & g[17187];
assign g[33572] = a[14] & g[17188];
assign g[49955] = b[14] & g[17188];
assign g[33573] = a[14] & g[17189];
assign g[49956] = b[14] & g[17189];
assign g[33574] = a[14] & g[17190];
assign g[49957] = b[14] & g[17190];
assign g[33575] = a[14] & g[17191];
assign g[49958] = b[14] & g[17191];
assign g[33576] = a[14] & g[17192];
assign g[49959] = b[14] & g[17192];
assign g[33577] = a[14] & g[17193];
assign g[49960] = b[14] & g[17193];
assign g[33578] = a[14] & g[17194];
assign g[49961] = b[14] & g[17194];
assign g[33579] = a[14] & g[17195];
assign g[49962] = b[14] & g[17195];
assign g[33580] = a[14] & g[17196];
assign g[49963] = b[14] & g[17196];
assign g[33581] = a[14] & g[17197];
assign g[49964] = b[14] & g[17197];
assign g[33582] = a[14] & g[17198];
assign g[49965] = b[14] & g[17198];
assign g[33583] = a[14] & g[17199];
assign g[49966] = b[14] & g[17199];
assign g[33584] = a[14] & g[17200];
assign g[49967] = b[14] & g[17200];
assign g[33585] = a[14] & g[17201];
assign g[49968] = b[14] & g[17201];
assign g[33586] = a[14] & g[17202];
assign g[49969] = b[14] & g[17202];
assign g[33587] = a[14] & g[17203];
assign g[49970] = b[14] & g[17203];
assign g[33588] = a[14] & g[17204];
assign g[49971] = b[14] & g[17204];
assign g[33589] = a[14] & g[17205];
assign g[49972] = b[14] & g[17205];
assign g[33590] = a[14] & g[17206];
assign g[49973] = b[14] & g[17206];
assign g[33591] = a[14] & g[17207];
assign g[49974] = b[14] & g[17207];
assign g[33592] = a[14] & g[17208];
assign g[49975] = b[14] & g[17208];
assign g[33593] = a[14] & g[17209];
assign g[49976] = b[14] & g[17209];
assign g[33594] = a[14] & g[17210];
assign g[49977] = b[14] & g[17210];
assign g[33595] = a[14] & g[17211];
assign g[49978] = b[14] & g[17211];
assign g[33596] = a[14] & g[17212];
assign g[49979] = b[14] & g[17212];
assign g[33597] = a[14] & g[17213];
assign g[49980] = b[14] & g[17213];
assign g[33598] = a[14] & g[17214];
assign g[49981] = b[14] & g[17214];
assign g[33599] = a[14] & g[17215];
assign g[49982] = b[14] & g[17215];
assign g[33600] = a[14] & g[17216];
assign g[49983] = b[14] & g[17216];
assign g[33601] = a[14] & g[17217];
assign g[49984] = b[14] & g[17217];
assign g[33602] = a[14] & g[17218];
assign g[49985] = b[14] & g[17218];
assign g[33603] = a[14] & g[17219];
assign g[49986] = b[14] & g[17219];
assign g[33604] = a[14] & g[17220];
assign g[49987] = b[14] & g[17220];
assign g[33605] = a[14] & g[17221];
assign g[49988] = b[14] & g[17221];
assign g[33606] = a[14] & g[17222];
assign g[49989] = b[14] & g[17222];
assign g[33607] = a[14] & g[17223];
assign g[49990] = b[14] & g[17223];
assign g[33608] = a[14] & g[17224];
assign g[49991] = b[14] & g[17224];
assign g[33609] = a[14] & g[17225];
assign g[49992] = b[14] & g[17225];
assign g[33610] = a[14] & g[17226];
assign g[49993] = b[14] & g[17226];
assign g[33611] = a[14] & g[17227];
assign g[49994] = b[14] & g[17227];
assign g[33612] = a[14] & g[17228];
assign g[49995] = b[14] & g[17228];
assign g[33613] = a[14] & g[17229];
assign g[49996] = b[14] & g[17229];
assign g[33614] = a[14] & g[17230];
assign g[49997] = b[14] & g[17230];
assign g[33615] = a[14] & g[17231];
assign g[49998] = b[14] & g[17231];
assign g[33616] = a[14] & g[17232];
assign g[49999] = b[14] & g[17232];
assign g[33617] = a[14] & g[17233];
assign g[50000] = b[14] & g[17233];
assign g[33618] = a[14] & g[17234];
assign g[50001] = b[14] & g[17234];
assign g[33619] = a[14] & g[17235];
assign g[50002] = b[14] & g[17235];
assign g[33620] = a[14] & g[17236];
assign g[50003] = b[14] & g[17236];
assign g[33621] = a[14] & g[17237];
assign g[50004] = b[14] & g[17237];
assign g[33622] = a[14] & g[17238];
assign g[50005] = b[14] & g[17238];
assign g[33623] = a[14] & g[17239];
assign g[50006] = b[14] & g[17239];
assign g[33624] = a[14] & g[17240];
assign g[50007] = b[14] & g[17240];
assign g[33625] = a[14] & g[17241];
assign g[50008] = b[14] & g[17241];
assign g[33626] = a[14] & g[17242];
assign g[50009] = b[14] & g[17242];
assign g[33627] = a[14] & g[17243];
assign g[50010] = b[14] & g[17243];
assign g[33628] = a[14] & g[17244];
assign g[50011] = b[14] & g[17244];
assign g[33629] = a[14] & g[17245];
assign g[50012] = b[14] & g[17245];
assign g[33630] = a[14] & g[17246];
assign g[50013] = b[14] & g[17246];
assign g[33631] = a[14] & g[17247];
assign g[50014] = b[14] & g[17247];
assign g[33632] = a[14] & g[17248];
assign g[50015] = b[14] & g[17248];
assign g[33633] = a[14] & g[17249];
assign g[50016] = b[14] & g[17249];
assign g[33634] = a[14] & g[17250];
assign g[50017] = b[14] & g[17250];
assign g[33635] = a[14] & g[17251];
assign g[50018] = b[14] & g[17251];
assign g[33636] = a[14] & g[17252];
assign g[50019] = b[14] & g[17252];
assign g[33637] = a[14] & g[17253];
assign g[50020] = b[14] & g[17253];
assign g[33638] = a[14] & g[17254];
assign g[50021] = b[14] & g[17254];
assign g[33639] = a[14] & g[17255];
assign g[50022] = b[14] & g[17255];
assign g[33640] = a[14] & g[17256];
assign g[50023] = b[14] & g[17256];
assign g[33641] = a[14] & g[17257];
assign g[50024] = b[14] & g[17257];
assign g[33642] = a[14] & g[17258];
assign g[50025] = b[14] & g[17258];
assign g[33643] = a[14] & g[17259];
assign g[50026] = b[14] & g[17259];
assign g[33644] = a[14] & g[17260];
assign g[50027] = b[14] & g[17260];
assign g[33645] = a[14] & g[17261];
assign g[50028] = b[14] & g[17261];
assign g[33646] = a[14] & g[17262];
assign g[50029] = b[14] & g[17262];
assign g[33647] = a[14] & g[17263];
assign g[50030] = b[14] & g[17263];
assign g[33648] = a[14] & g[17264];
assign g[50031] = b[14] & g[17264];
assign g[33649] = a[14] & g[17265];
assign g[50032] = b[14] & g[17265];
assign g[33650] = a[14] & g[17266];
assign g[50033] = b[14] & g[17266];
assign g[33651] = a[14] & g[17267];
assign g[50034] = b[14] & g[17267];
assign g[33652] = a[14] & g[17268];
assign g[50035] = b[14] & g[17268];
assign g[33653] = a[14] & g[17269];
assign g[50036] = b[14] & g[17269];
assign g[33654] = a[14] & g[17270];
assign g[50037] = b[14] & g[17270];
assign g[33655] = a[14] & g[17271];
assign g[50038] = b[14] & g[17271];
assign g[33656] = a[14] & g[17272];
assign g[50039] = b[14] & g[17272];
assign g[33657] = a[14] & g[17273];
assign g[50040] = b[14] & g[17273];
assign g[33658] = a[14] & g[17274];
assign g[50041] = b[14] & g[17274];
assign g[33659] = a[14] & g[17275];
assign g[50042] = b[14] & g[17275];
assign g[33660] = a[14] & g[17276];
assign g[50043] = b[14] & g[17276];
assign g[33661] = a[14] & g[17277];
assign g[50044] = b[14] & g[17277];
assign g[33662] = a[14] & g[17278];
assign g[50045] = b[14] & g[17278];
assign g[33663] = a[14] & g[17279];
assign g[50046] = b[14] & g[17279];
assign g[33664] = a[14] & g[17280];
assign g[50047] = b[14] & g[17280];
assign g[33665] = a[14] & g[17281];
assign g[50048] = b[14] & g[17281];
assign g[33666] = a[14] & g[17282];
assign g[50049] = b[14] & g[17282];
assign g[33667] = a[14] & g[17283];
assign g[50050] = b[14] & g[17283];
assign g[33668] = a[14] & g[17284];
assign g[50051] = b[14] & g[17284];
assign g[33669] = a[14] & g[17285];
assign g[50052] = b[14] & g[17285];
assign g[33670] = a[14] & g[17286];
assign g[50053] = b[14] & g[17286];
assign g[33671] = a[14] & g[17287];
assign g[50054] = b[14] & g[17287];
assign g[33672] = a[14] & g[17288];
assign g[50055] = b[14] & g[17288];
assign g[33673] = a[14] & g[17289];
assign g[50056] = b[14] & g[17289];
assign g[33674] = a[14] & g[17290];
assign g[50057] = b[14] & g[17290];
assign g[33675] = a[14] & g[17291];
assign g[50058] = b[14] & g[17291];
assign g[33676] = a[14] & g[17292];
assign g[50059] = b[14] & g[17292];
assign g[33677] = a[14] & g[17293];
assign g[50060] = b[14] & g[17293];
assign g[33678] = a[14] & g[17294];
assign g[50061] = b[14] & g[17294];
assign g[33679] = a[14] & g[17295];
assign g[50062] = b[14] & g[17295];
assign g[33680] = a[14] & g[17296];
assign g[50063] = b[14] & g[17296];
assign g[33681] = a[14] & g[17297];
assign g[50064] = b[14] & g[17297];
assign g[33682] = a[14] & g[17298];
assign g[50065] = b[14] & g[17298];
assign g[33683] = a[14] & g[17299];
assign g[50066] = b[14] & g[17299];
assign g[33684] = a[14] & g[17300];
assign g[50067] = b[14] & g[17300];
assign g[33685] = a[14] & g[17301];
assign g[50068] = b[14] & g[17301];
assign g[33686] = a[14] & g[17302];
assign g[50069] = b[14] & g[17302];
assign g[33687] = a[14] & g[17303];
assign g[50070] = b[14] & g[17303];
assign g[33688] = a[14] & g[17304];
assign g[50071] = b[14] & g[17304];
assign g[33689] = a[14] & g[17305];
assign g[50072] = b[14] & g[17305];
assign g[33690] = a[14] & g[17306];
assign g[50073] = b[14] & g[17306];
assign g[33691] = a[14] & g[17307];
assign g[50074] = b[14] & g[17307];
assign g[33692] = a[14] & g[17308];
assign g[50075] = b[14] & g[17308];
assign g[33693] = a[14] & g[17309];
assign g[50076] = b[14] & g[17309];
assign g[33694] = a[14] & g[17310];
assign g[50077] = b[14] & g[17310];
assign g[33695] = a[14] & g[17311];
assign g[50078] = b[14] & g[17311];
assign g[33696] = a[14] & g[17312];
assign g[50079] = b[14] & g[17312];
assign g[33697] = a[14] & g[17313];
assign g[50080] = b[14] & g[17313];
assign g[33698] = a[14] & g[17314];
assign g[50081] = b[14] & g[17314];
assign g[33699] = a[14] & g[17315];
assign g[50082] = b[14] & g[17315];
assign g[33700] = a[14] & g[17316];
assign g[50083] = b[14] & g[17316];
assign g[33701] = a[14] & g[17317];
assign g[50084] = b[14] & g[17317];
assign g[33702] = a[14] & g[17318];
assign g[50085] = b[14] & g[17318];
assign g[33703] = a[14] & g[17319];
assign g[50086] = b[14] & g[17319];
assign g[33704] = a[14] & g[17320];
assign g[50087] = b[14] & g[17320];
assign g[33705] = a[14] & g[17321];
assign g[50088] = b[14] & g[17321];
assign g[33706] = a[14] & g[17322];
assign g[50089] = b[14] & g[17322];
assign g[33707] = a[14] & g[17323];
assign g[50090] = b[14] & g[17323];
assign g[33708] = a[14] & g[17324];
assign g[50091] = b[14] & g[17324];
assign g[33709] = a[14] & g[17325];
assign g[50092] = b[14] & g[17325];
assign g[33710] = a[14] & g[17326];
assign g[50093] = b[14] & g[17326];
assign g[33711] = a[14] & g[17327];
assign g[50094] = b[14] & g[17327];
assign g[33712] = a[14] & g[17328];
assign g[50095] = b[14] & g[17328];
assign g[33713] = a[14] & g[17329];
assign g[50096] = b[14] & g[17329];
assign g[33714] = a[14] & g[17330];
assign g[50097] = b[14] & g[17330];
assign g[33715] = a[14] & g[17331];
assign g[50098] = b[14] & g[17331];
assign g[33716] = a[14] & g[17332];
assign g[50099] = b[14] & g[17332];
assign g[33717] = a[14] & g[17333];
assign g[50100] = b[14] & g[17333];
assign g[33718] = a[14] & g[17334];
assign g[50101] = b[14] & g[17334];
assign g[33719] = a[14] & g[17335];
assign g[50102] = b[14] & g[17335];
assign g[33720] = a[14] & g[17336];
assign g[50103] = b[14] & g[17336];
assign g[33721] = a[14] & g[17337];
assign g[50104] = b[14] & g[17337];
assign g[33722] = a[14] & g[17338];
assign g[50105] = b[14] & g[17338];
assign g[33723] = a[14] & g[17339];
assign g[50106] = b[14] & g[17339];
assign g[33724] = a[14] & g[17340];
assign g[50107] = b[14] & g[17340];
assign g[33725] = a[14] & g[17341];
assign g[50108] = b[14] & g[17341];
assign g[33726] = a[14] & g[17342];
assign g[50109] = b[14] & g[17342];
assign g[33727] = a[14] & g[17343];
assign g[50110] = b[14] & g[17343];
assign g[33728] = a[14] & g[17344];
assign g[50111] = b[14] & g[17344];
assign g[33729] = a[14] & g[17345];
assign g[50112] = b[14] & g[17345];
assign g[33730] = a[14] & g[17346];
assign g[50113] = b[14] & g[17346];
assign g[33731] = a[14] & g[17347];
assign g[50114] = b[14] & g[17347];
assign g[33732] = a[14] & g[17348];
assign g[50115] = b[14] & g[17348];
assign g[33733] = a[14] & g[17349];
assign g[50116] = b[14] & g[17349];
assign g[33734] = a[14] & g[17350];
assign g[50117] = b[14] & g[17350];
assign g[33735] = a[14] & g[17351];
assign g[50118] = b[14] & g[17351];
assign g[33736] = a[14] & g[17352];
assign g[50119] = b[14] & g[17352];
assign g[33737] = a[14] & g[17353];
assign g[50120] = b[14] & g[17353];
assign g[33738] = a[14] & g[17354];
assign g[50121] = b[14] & g[17354];
assign g[33739] = a[14] & g[17355];
assign g[50122] = b[14] & g[17355];
assign g[33740] = a[14] & g[17356];
assign g[50123] = b[14] & g[17356];
assign g[33741] = a[14] & g[17357];
assign g[50124] = b[14] & g[17357];
assign g[33742] = a[14] & g[17358];
assign g[50125] = b[14] & g[17358];
assign g[33743] = a[14] & g[17359];
assign g[50126] = b[14] & g[17359];
assign g[33744] = a[14] & g[17360];
assign g[50127] = b[14] & g[17360];
assign g[33745] = a[14] & g[17361];
assign g[50128] = b[14] & g[17361];
assign g[33746] = a[14] & g[17362];
assign g[50129] = b[14] & g[17362];
assign g[33747] = a[14] & g[17363];
assign g[50130] = b[14] & g[17363];
assign g[33748] = a[14] & g[17364];
assign g[50131] = b[14] & g[17364];
assign g[33749] = a[14] & g[17365];
assign g[50132] = b[14] & g[17365];
assign g[33750] = a[14] & g[17366];
assign g[50133] = b[14] & g[17366];
assign g[33751] = a[14] & g[17367];
assign g[50134] = b[14] & g[17367];
assign g[33752] = a[14] & g[17368];
assign g[50135] = b[14] & g[17368];
assign g[33753] = a[14] & g[17369];
assign g[50136] = b[14] & g[17369];
assign g[33754] = a[14] & g[17370];
assign g[50137] = b[14] & g[17370];
assign g[33755] = a[14] & g[17371];
assign g[50138] = b[14] & g[17371];
assign g[33756] = a[14] & g[17372];
assign g[50139] = b[14] & g[17372];
assign g[33757] = a[14] & g[17373];
assign g[50140] = b[14] & g[17373];
assign g[33758] = a[14] & g[17374];
assign g[50141] = b[14] & g[17374];
assign g[33759] = a[14] & g[17375];
assign g[50142] = b[14] & g[17375];
assign g[33760] = a[14] & g[17376];
assign g[50143] = b[14] & g[17376];
assign g[33761] = a[14] & g[17377];
assign g[50144] = b[14] & g[17377];
assign g[33762] = a[14] & g[17378];
assign g[50145] = b[14] & g[17378];
assign g[33763] = a[14] & g[17379];
assign g[50146] = b[14] & g[17379];
assign g[33764] = a[14] & g[17380];
assign g[50147] = b[14] & g[17380];
assign g[33765] = a[14] & g[17381];
assign g[50148] = b[14] & g[17381];
assign g[33766] = a[14] & g[17382];
assign g[50149] = b[14] & g[17382];
assign g[33767] = a[14] & g[17383];
assign g[50150] = b[14] & g[17383];
assign g[33768] = a[14] & g[17384];
assign g[50151] = b[14] & g[17384];
assign g[33769] = a[14] & g[17385];
assign g[50152] = b[14] & g[17385];
assign g[33770] = a[14] & g[17386];
assign g[50153] = b[14] & g[17386];
assign g[33771] = a[14] & g[17387];
assign g[50154] = b[14] & g[17387];
assign g[33772] = a[14] & g[17388];
assign g[50155] = b[14] & g[17388];
assign g[33773] = a[14] & g[17389];
assign g[50156] = b[14] & g[17389];
assign g[33774] = a[14] & g[17390];
assign g[50157] = b[14] & g[17390];
assign g[33775] = a[14] & g[17391];
assign g[50158] = b[14] & g[17391];
assign g[33776] = a[14] & g[17392];
assign g[50159] = b[14] & g[17392];
assign g[33777] = a[14] & g[17393];
assign g[50160] = b[14] & g[17393];
assign g[33778] = a[14] & g[17394];
assign g[50161] = b[14] & g[17394];
assign g[33779] = a[14] & g[17395];
assign g[50162] = b[14] & g[17395];
assign g[33780] = a[14] & g[17396];
assign g[50163] = b[14] & g[17396];
assign g[33781] = a[14] & g[17397];
assign g[50164] = b[14] & g[17397];
assign g[33782] = a[14] & g[17398];
assign g[50165] = b[14] & g[17398];
assign g[33783] = a[14] & g[17399];
assign g[50166] = b[14] & g[17399];
assign g[33784] = a[14] & g[17400];
assign g[50167] = b[14] & g[17400];
assign g[33785] = a[14] & g[17401];
assign g[50168] = b[14] & g[17401];
assign g[33786] = a[14] & g[17402];
assign g[50169] = b[14] & g[17402];
assign g[33787] = a[14] & g[17403];
assign g[50170] = b[14] & g[17403];
assign g[33788] = a[14] & g[17404];
assign g[50171] = b[14] & g[17404];
assign g[33789] = a[14] & g[17405];
assign g[50172] = b[14] & g[17405];
assign g[33790] = a[14] & g[17406];
assign g[50173] = b[14] & g[17406];
assign g[33791] = a[14] & g[17407];
assign g[50174] = b[14] & g[17407];
assign g[33792] = a[14] & g[17408];
assign g[50175] = b[14] & g[17408];
assign g[33793] = a[14] & g[17409];
assign g[50176] = b[14] & g[17409];
assign g[33794] = a[14] & g[17410];
assign g[50177] = b[14] & g[17410];
assign g[33795] = a[14] & g[17411];
assign g[50178] = b[14] & g[17411];
assign g[33796] = a[14] & g[17412];
assign g[50179] = b[14] & g[17412];
assign g[33797] = a[14] & g[17413];
assign g[50180] = b[14] & g[17413];
assign g[33798] = a[14] & g[17414];
assign g[50181] = b[14] & g[17414];
assign g[33799] = a[14] & g[17415];
assign g[50182] = b[14] & g[17415];
assign g[33800] = a[14] & g[17416];
assign g[50183] = b[14] & g[17416];
assign g[33801] = a[14] & g[17417];
assign g[50184] = b[14] & g[17417];
assign g[33802] = a[14] & g[17418];
assign g[50185] = b[14] & g[17418];
assign g[33803] = a[14] & g[17419];
assign g[50186] = b[14] & g[17419];
assign g[33804] = a[14] & g[17420];
assign g[50187] = b[14] & g[17420];
assign g[33805] = a[14] & g[17421];
assign g[50188] = b[14] & g[17421];
assign g[33806] = a[14] & g[17422];
assign g[50189] = b[14] & g[17422];
assign g[33807] = a[14] & g[17423];
assign g[50190] = b[14] & g[17423];
assign g[33808] = a[14] & g[17424];
assign g[50191] = b[14] & g[17424];
assign g[33809] = a[14] & g[17425];
assign g[50192] = b[14] & g[17425];
assign g[33810] = a[14] & g[17426];
assign g[50193] = b[14] & g[17426];
assign g[33811] = a[14] & g[17427];
assign g[50194] = b[14] & g[17427];
assign g[33812] = a[14] & g[17428];
assign g[50195] = b[14] & g[17428];
assign g[33813] = a[14] & g[17429];
assign g[50196] = b[14] & g[17429];
assign g[33814] = a[14] & g[17430];
assign g[50197] = b[14] & g[17430];
assign g[33815] = a[14] & g[17431];
assign g[50198] = b[14] & g[17431];
assign g[33816] = a[14] & g[17432];
assign g[50199] = b[14] & g[17432];
assign g[33817] = a[14] & g[17433];
assign g[50200] = b[14] & g[17433];
assign g[33818] = a[14] & g[17434];
assign g[50201] = b[14] & g[17434];
assign g[33819] = a[14] & g[17435];
assign g[50202] = b[14] & g[17435];
assign g[33820] = a[14] & g[17436];
assign g[50203] = b[14] & g[17436];
assign g[33821] = a[14] & g[17437];
assign g[50204] = b[14] & g[17437];
assign g[33822] = a[14] & g[17438];
assign g[50205] = b[14] & g[17438];
assign g[33823] = a[14] & g[17439];
assign g[50206] = b[14] & g[17439];
assign g[33824] = a[14] & g[17440];
assign g[50207] = b[14] & g[17440];
assign g[33825] = a[14] & g[17441];
assign g[50208] = b[14] & g[17441];
assign g[33826] = a[14] & g[17442];
assign g[50209] = b[14] & g[17442];
assign g[33827] = a[14] & g[17443];
assign g[50210] = b[14] & g[17443];
assign g[33828] = a[14] & g[17444];
assign g[50211] = b[14] & g[17444];
assign g[33829] = a[14] & g[17445];
assign g[50212] = b[14] & g[17445];
assign g[33830] = a[14] & g[17446];
assign g[50213] = b[14] & g[17446];
assign g[33831] = a[14] & g[17447];
assign g[50214] = b[14] & g[17447];
assign g[33832] = a[14] & g[17448];
assign g[50215] = b[14] & g[17448];
assign g[33833] = a[14] & g[17449];
assign g[50216] = b[14] & g[17449];
assign g[33834] = a[14] & g[17450];
assign g[50217] = b[14] & g[17450];
assign g[33835] = a[14] & g[17451];
assign g[50218] = b[14] & g[17451];
assign g[33836] = a[14] & g[17452];
assign g[50219] = b[14] & g[17452];
assign g[33837] = a[14] & g[17453];
assign g[50220] = b[14] & g[17453];
assign g[33838] = a[14] & g[17454];
assign g[50221] = b[14] & g[17454];
assign g[33839] = a[14] & g[17455];
assign g[50222] = b[14] & g[17455];
assign g[33840] = a[14] & g[17456];
assign g[50223] = b[14] & g[17456];
assign g[33841] = a[14] & g[17457];
assign g[50224] = b[14] & g[17457];
assign g[33842] = a[14] & g[17458];
assign g[50225] = b[14] & g[17458];
assign g[33843] = a[14] & g[17459];
assign g[50226] = b[14] & g[17459];
assign g[33844] = a[14] & g[17460];
assign g[50227] = b[14] & g[17460];
assign g[33845] = a[14] & g[17461];
assign g[50228] = b[14] & g[17461];
assign g[33846] = a[14] & g[17462];
assign g[50229] = b[14] & g[17462];
assign g[33847] = a[14] & g[17463];
assign g[50230] = b[14] & g[17463];
assign g[33848] = a[14] & g[17464];
assign g[50231] = b[14] & g[17464];
assign g[33849] = a[14] & g[17465];
assign g[50232] = b[14] & g[17465];
assign g[33850] = a[14] & g[17466];
assign g[50233] = b[14] & g[17466];
assign g[33851] = a[14] & g[17467];
assign g[50234] = b[14] & g[17467];
assign g[33852] = a[14] & g[17468];
assign g[50235] = b[14] & g[17468];
assign g[33853] = a[14] & g[17469];
assign g[50236] = b[14] & g[17469];
assign g[33854] = a[14] & g[17470];
assign g[50237] = b[14] & g[17470];
assign g[33855] = a[14] & g[17471];
assign g[50238] = b[14] & g[17471];
assign g[33856] = a[14] & g[17472];
assign g[50239] = b[14] & g[17472];
assign g[33857] = a[14] & g[17473];
assign g[50240] = b[14] & g[17473];
assign g[33858] = a[14] & g[17474];
assign g[50241] = b[14] & g[17474];
assign g[33859] = a[14] & g[17475];
assign g[50242] = b[14] & g[17475];
assign g[33860] = a[14] & g[17476];
assign g[50243] = b[14] & g[17476];
assign g[33861] = a[14] & g[17477];
assign g[50244] = b[14] & g[17477];
assign g[33862] = a[14] & g[17478];
assign g[50245] = b[14] & g[17478];
assign g[33863] = a[14] & g[17479];
assign g[50246] = b[14] & g[17479];
assign g[33864] = a[14] & g[17480];
assign g[50247] = b[14] & g[17480];
assign g[33865] = a[14] & g[17481];
assign g[50248] = b[14] & g[17481];
assign g[33866] = a[14] & g[17482];
assign g[50249] = b[14] & g[17482];
assign g[33867] = a[14] & g[17483];
assign g[50250] = b[14] & g[17483];
assign g[33868] = a[14] & g[17484];
assign g[50251] = b[14] & g[17484];
assign g[33869] = a[14] & g[17485];
assign g[50252] = b[14] & g[17485];
assign g[33870] = a[14] & g[17486];
assign g[50253] = b[14] & g[17486];
assign g[33871] = a[14] & g[17487];
assign g[50254] = b[14] & g[17487];
assign g[33872] = a[14] & g[17488];
assign g[50255] = b[14] & g[17488];
assign g[33873] = a[14] & g[17489];
assign g[50256] = b[14] & g[17489];
assign g[33874] = a[14] & g[17490];
assign g[50257] = b[14] & g[17490];
assign g[33875] = a[14] & g[17491];
assign g[50258] = b[14] & g[17491];
assign g[33876] = a[14] & g[17492];
assign g[50259] = b[14] & g[17492];
assign g[33877] = a[14] & g[17493];
assign g[50260] = b[14] & g[17493];
assign g[33878] = a[14] & g[17494];
assign g[50261] = b[14] & g[17494];
assign g[33879] = a[14] & g[17495];
assign g[50262] = b[14] & g[17495];
assign g[33880] = a[14] & g[17496];
assign g[50263] = b[14] & g[17496];
assign g[33881] = a[14] & g[17497];
assign g[50264] = b[14] & g[17497];
assign g[33882] = a[14] & g[17498];
assign g[50265] = b[14] & g[17498];
assign g[33883] = a[14] & g[17499];
assign g[50266] = b[14] & g[17499];
assign g[33884] = a[14] & g[17500];
assign g[50267] = b[14] & g[17500];
assign g[33885] = a[14] & g[17501];
assign g[50268] = b[14] & g[17501];
assign g[33886] = a[14] & g[17502];
assign g[50269] = b[14] & g[17502];
assign g[33887] = a[14] & g[17503];
assign g[50270] = b[14] & g[17503];
assign g[33888] = a[14] & g[17504];
assign g[50271] = b[14] & g[17504];
assign g[33889] = a[14] & g[17505];
assign g[50272] = b[14] & g[17505];
assign g[33890] = a[14] & g[17506];
assign g[50273] = b[14] & g[17506];
assign g[33891] = a[14] & g[17507];
assign g[50274] = b[14] & g[17507];
assign g[33892] = a[14] & g[17508];
assign g[50275] = b[14] & g[17508];
assign g[33893] = a[14] & g[17509];
assign g[50276] = b[14] & g[17509];
assign g[33894] = a[14] & g[17510];
assign g[50277] = b[14] & g[17510];
assign g[33895] = a[14] & g[17511];
assign g[50278] = b[14] & g[17511];
assign g[33896] = a[14] & g[17512];
assign g[50279] = b[14] & g[17512];
assign g[33897] = a[14] & g[17513];
assign g[50280] = b[14] & g[17513];
assign g[33898] = a[14] & g[17514];
assign g[50281] = b[14] & g[17514];
assign g[33899] = a[14] & g[17515];
assign g[50282] = b[14] & g[17515];
assign g[33900] = a[14] & g[17516];
assign g[50283] = b[14] & g[17516];
assign g[33901] = a[14] & g[17517];
assign g[50284] = b[14] & g[17517];
assign g[33902] = a[14] & g[17518];
assign g[50285] = b[14] & g[17518];
assign g[33903] = a[14] & g[17519];
assign g[50286] = b[14] & g[17519];
assign g[33904] = a[14] & g[17520];
assign g[50287] = b[14] & g[17520];
assign g[33905] = a[14] & g[17521];
assign g[50288] = b[14] & g[17521];
assign g[33906] = a[14] & g[17522];
assign g[50289] = b[14] & g[17522];
assign g[33907] = a[14] & g[17523];
assign g[50290] = b[14] & g[17523];
assign g[33908] = a[14] & g[17524];
assign g[50291] = b[14] & g[17524];
assign g[33909] = a[14] & g[17525];
assign g[50292] = b[14] & g[17525];
assign g[33910] = a[14] & g[17526];
assign g[50293] = b[14] & g[17526];
assign g[33911] = a[14] & g[17527];
assign g[50294] = b[14] & g[17527];
assign g[33912] = a[14] & g[17528];
assign g[50295] = b[14] & g[17528];
assign g[33913] = a[14] & g[17529];
assign g[50296] = b[14] & g[17529];
assign g[33914] = a[14] & g[17530];
assign g[50297] = b[14] & g[17530];
assign g[33915] = a[14] & g[17531];
assign g[50298] = b[14] & g[17531];
assign g[33916] = a[14] & g[17532];
assign g[50299] = b[14] & g[17532];
assign g[33917] = a[14] & g[17533];
assign g[50300] = b[14] & g[17533];
assign g[33918] = a[14] & g[17534];
assign g[50301] = b[14] & g[17534];
assign g[33919] = a[14] & g[17535];
assign g[50302] = b[14] & g[17535];
assign g[33920] = a[14] & g[17536];
assign g[50303] = b[14] & g[17536];
assign g[33921] = a[14] & g[17537];
assign g[50304] = b[14] & g[17537];
assign g[33922] = a[14] & g[17538];
assign g[50305] = b[14] & g[17538];
assign g[33923] = a[14] & g[17539];
assign g[50306] = b[14] & g[17539];
assign g[33924] = a[14] & g[17540];
assign g[50307] = b[14] & g[17540];
assign g[33925] = a[14] & g[17541];
assign g[50308] = b[14] & g[17541];
assign g[33926] = a[14] & g[17542];
assign g[50309] = b[14] & g[17542];
assign g[33927] = a[14] & g[17543];
assign g[50310] = b[14] & g[17543];
assign g[33928] = a[14] & g[17544];
assign g[50311] = b[14] & g[17544];
assign g[33929] = a[14] & g[17545];
assign g[50312] = b[14] & g[17545];
assign g[33930] = a[14] & g[17546];
assign g[50313] = b[14] & g[17546];
assign g[33931] = a[14] & g[17547];
assign g[50314] = b[14] & g[17547];
assign g[33932] = a[14] & g[17548];
assign g[50315] = b[14] & g[17548];
assign g[33933] = a[14] & g[17549];
assign g[50316] = b[14] & g[17549];
assign g[33934] = a[14] & g[17550];
assign g[50317] = b[14] & g[17550];
assign g[33935] = a[14] & g[17551];
assign g[50318] = b[14] & g[17551];
assign g[33936] = a[14] & g[17552];
assign g[50319] = b[14] & g[17552];
assign g[33937] = a[14] & g[17553];
assign g[50320] = b[14] & g[17553];
assign g[33938] = a[14] & g[17554];
assign g[50321] = b[14] & g[17554];
assign g[33939] = a[14] & g[17555];
assign g[50322] = b[14] & g[17555];
assign g[33940] = a[14] & g[17556];
assign g[50323] = b[14] & g[17556];
assign g[33941] = a[14] & g[17557];
assign g[50324] = b[14] & g[17557];
assign g[33942] = a[14] & g[17558];
assign g[50325] = b[14] & g[17558];
assign g[33943] = a[14] & g[17559];
assign g[50326] = b[14] & g[17559];
assign g[33944] = a[14] & g[17560];
assign g[50327] = b[14] & g[17560];
assign g[33945] = a[14] & g[17561];
assign g[50328] = b[14] & g[17561];
assign g[33946] = a[14] & g[17562];
assign g[50329] = b[14] & g[17562];
assign g[33947] = a[14] & g[17563];
assign g[50330] = b[14] & g[17563];
assign g[33948] = a[14] & g[17564];
assign g[50331] = b[14] & g[17564];
assign g[33949] = a[14] & g[17565];
assign g[50332] = b[14] & g[17565];
assign g[33950] = a[14] & g[17566];
assign g[50333] = b[14] & g[17566];
assign g[33951] = a[14] & g[17567];
assign g[50334] = b[14] & g[17567];
assign g[33952] = a[14] & g[17568];
assign g[50335] = b[14] & g[17568];
assign g[33953] = a[14] & g[17569];
assign g[50336] = b[14] & g[17569];
assign g[33954] = a[14] & g[17570];
assign g[50337] = b[14] & g[17570];
assign g[33955] = a[14] & g[17571];
assign g[50338] = b[14] & g[17571];
assign g[33956] = a[14] & g[17572];
assign g[50339] = b[14] & g[17572];
assign g[33957] = a[14] & g[17573];
assign g[50340] = b[14] & g[17573];
assign g[33958] = a[14] & g[17574];
assign g[50341] = b[14] & g[17574];
assign g[33959] = a[14] & g[17575];
assign g[50342] = b[14] & g[17575];
assign g[33960] = a[14] & g[17576];
assign g[50343] = b[14] & g[17576];
assign g[33961] = a[14] & g[17577];
assign g[50344] = b[14] & g[17577];
assign g[33962] = a[14] & g[17578];
assign g[50345] = b[14] & g[17578];
assign g[33963] = a[14] & g[17579];
assign g[50346] = b[14] & g[17579];
assign g[33964] = a[14] & g[17580];
assign g[50347] = b[14] & g[17580];
assign g[33965] = a[14] & g[17581];
assign g[50348] = b[14] & g[17581];
assign g[33966] = a[14] & g[17582];
assign g[50349] = b[14] & g[17582];
assign g[33967] = a[14] & g[17583];
assign g[50350] = b[14] & g[17583];
assign g[33968] = a[14] & g[17584];
assign g[50351] = b[14] & g[17584];
assign g[33969] = a[14] & g[17585];
assign g[50352] = b[14] & g[17585];
assign g[33970] = a[14] & g[17586];
assign g[50353] = b[14] & g[17586];
assign g[33971] = a[14] & g[17587];
assign g[50354] = b[14] & g[17587];
assign g[33972] = a[14] & g[17588];
assign g[50355] = b[14] & g[17588];
assign g[33973] = a[14] & g[17589];
assign g[50356] = b[14] & g[17589];
assign g[33974] = a[14] & g[17590];
assign g[50357] = b[14] & g[17590];
assign g[33975] = a[14] & g[17591];
assign g[50358] = b[14] & g[17591];
assign g[33976] = a[14] & g[17592];
assign g[50359] = b[14] & g[17592];
assign g[33977] = a[14] & g[17593];
assign g[50360] = b[14] & g[17593];
assign g[33978] = a[14] & g[17594];
assign g[50361] = b[14] & g[17594];
assign g[33979] = a[14] & g[17595];
assign g[50362] = b[14] & g[17595];
assign g[33980] = a[14] & g[17596];
assign g[50363] = b[14] & g[17596];
assign g[33981] = a[14] & g[17597];
assign g[50364] = b[14] & g[17597];
assign g[33982] = a[14] & g[17598];
assign g[50365] = b[14] & g[17598];
assign g[33983] = a[14] & g[17599];
assign g[50366] = b[14] & g[17599];
assign g[33984] = a[14] & g[17600];
assign g[50367] = b[14] & g[17600];
assign g[33985] = a[14] & g[17601];
assign g[50368] = b[14] & g[17601];
assign g[33986] = a[14] & g[17602];
assign g[50369] = b[14] & g[17602];
assign g[33987] = a[14] & g[17603];
assign g[50370] = b[14] & g[17603];
assign g[33988] = a[14] & g[17604];
assign g[50371] = b[14] & g[17604];
assign g[33989] = a[14] & g[17605];
assign g[50372] = b[14] & g[17605];
assign g[33990] = a[14] & g[17606];
assign g[50373] = b[14] & g[17606];
assign g[33991] = a[14] & g[17607];
assign g[50374] = b[14] & g[17607];
assign g[33992] = a[14] & g[17608];
assign g[50375] = b[14] & g[17608];
assign g[33993] = a[14] & g[17609];
assign g[50376] = b[14] & g[17609];
assign g[33994] = a[14] & g[17610];
assign g[50377] = b[14] & g[17610];
assign g[33995] = a[14] & g[17611];
assign g[50378] = b[14] & g[17611];
assign g[33996] = a[14] & g[17612];
assign g[50379] = b[14] & g[17612];
assign g[33997] = a[14] & g[17613];
assign g[50380] = b[14] & g[17613];
assign g[33998] = a[14] & g[17614];
assign g[50381] = b[14] & g[17614];
assign g[33999] = a[14] & g[17615];
assign g[50382] = b[14] & g[17615];
assign g[34000] = a[14] & g[17616];
assign g[50383] = b[14] & g[17616];
assign g[34001] = a[14] & g[17617];
assign g[50384] = b[14] & g[17617];
assign g[34002] = a[14] & g[17618];
assign g[50385] = b[14] & g[17618];
assign g[34003] = a[14] & g[17619];
assign g[50386] = b[14] & g[17619];
assign g[34004] = a[14] & g[17620];
assign g[50387] = b[14] & g[17620];
assign g[34005] = a[14] & g[17621];
assign g[50388] = b[14] & g[17621];
assign g[34006] = a[14] & g[17622];
assign g[50389] = b[14] & g[17622];
assign g[34007] = a[14] & g[17623];
assign g[50390] = b[14] & g[17623];
assign g[34008] = a[14] & g[17624];
assign g[50391] = b[14] & g[17624];
assign g[34009] = a[14] & g[17625];
assign g[50392] = b[14] & g[17625];
assign g[34010] = a[14] & g[17626];
assign g[50393] = b[14] & g[17626];
assign g[34011] = a[14] & g[17627];
assign g[50394] = b[14] & g[17627];
assign g[34012] = a[14] & g[17628];
assign g[50395] = b[14] & g[17628];
assign g[34013] = a[14] & g[17629];
assign g[50396] = b[14] & g[17629];
assign g[34014] = a[14] & g[17630];
assign g[50397] = b[14] & g[17630];
assign g[34015] = a[14] & g[17631];
assign g[50398] = b[14] & g[17631];
assign g[34016] = a[14] & g[17632];
assign g[50399] = b[14] & g[17632];
assign g[34017] = a[14] & g[17633];
assign g[50400] = b[14] & g[17633];
assign g[34018] = a[14] & g[17634];
assign g[50401] = b[14] & g[17634];
assign g[34019] = a[14] & g[17635];
assign g[50402] = b[14] & g[17635];
assign g[34020] = a[14] & g[17636];
assign g[50403] = b[14] & g[17636];
assign g[34021] = a[14] & g[17637];
assign g[50404] = b[14] & g[17637];
assign g[34022] = a[14] & g[17638];
assign g[50405] = b[14] & g[17638];
assign g[34023] = a[14] & g[17639];
assign g[50406] = b[14] & g[17639];
assign g[34024] = a[14] & g[17640];
assign g[50407] = b[14] & g[17640];
assign g[34025] = a[14] & g[17641];
assign g[50408] = b[14] & g[17641];
assign g[34026] = a[14] & g[17642];
assign g[50409] = b[14] & g[17642];
assign g[34027] = a[14] & g[17643];
assign g[50410] = b[14] & g[17643];
assign g[34028] = a[14] & g[17644];
assign g[50411] = b[14] & g[17644];
assign g[34029] = a[14] & g[17645];
assign g[50412] = b[14] & g[17645];
assign g[34030] = a[14] & g[17646];
assign g[50413] = b[14] & g[17646];
assign g[34031] = a[14] & g[17647];
assign g[50414] = b[14] & g[17647];
assign g[34032] = a[14] & g[17648];
assign g[50415] = b[14] & g[17648];
assign g[34033] = a[14] & g[17649];
assign g[50416] = b[14] & g[17649];
assign g[34034] = a[14] & g[17650];
assign g[50417] = b[14] & g[17650];
assign g[34035] = a[14] & g[17651];
assign g[50418] = b[14] & g[17651];
assign g[34036] = a[14] & g[17652];
assign g[50419] = b[14] & g[17652];
assign g[34037] = a[14] & g[17653];
assign g[50420] = b[14] & g[17653];
assign g[34038] = a[14] & g[17654];
assign g[50421] = b[14] & g[17654];
assign g[34039] = a[14] & g[17655];
assign g[50422] = b[14] & g[17655];
assign g[34040] = a[14] & g[17656];
assign g[50423] = b[14] & g[17656];
assign g[34041] = a[14] & g[17657];
assign g[50424] = b[14] & g[17657];
assign g[34042] = a[14] & g[17658];
assign g[50425] = b[14] & g[17658];
assign g[34043] = a[14] & g[17659];
assign g[50426] = b[14] & g[17659];
assign g[34044] = a[14] & g[17660];
assign g[50427] = b[14] & g[17660];
assign g[34045] = a[14] & g[17661];
assign g[50428] = b[14] & g[17661];
assign g[34046] = a[14] & g[17662];
assign g[50429] = b[14] & g[17662];
assign g[34047] = a[14] & g[17663];
assign g[50430] = b[14] & g[17663];
assign g[34048] = a[14] & g[17664];
assign g[50431] = b[14] & g[17664];
assign g[34049] = a[14] & g[17665];
assign g[50432] = b[14] & g[17665];
assign g[34050] = a[14] & g[17666];
assign g[50433] = b[14] & g[17666];
assign g[34051] = a[14] & g[17667];
assign g[50434] = b[14] & g[17667];
assign g[34052] = a[14] & g[17668];
assign g[50435] = b[14] & g[17668];
assign g[34053] = a[14] & g[17669];
assign g[50436] = b[14] & g[17669];
assign g[34054] = a[14] & g[17670];
assign g[50437] = b[14] & g[17670];
assign g[34055] = a[14] & g[17671];
assign g[50438] = b[14] & g[17671];
assign g[34056] = a[14] & g[17672];
assign g[50439] = b[14] & g[17672];
assign g[34057] = a[14] & g[17673];
assign g[50440] = b[14] & g[17673];
assign g[34058] = a[14] & g[17674];
assign g[50441] = b[14] & g[17674];
assign g[34059] = a[14] & g[17675];
assign g[50442] = b[14] & g[17675];
assign g[34060] = a[14] & g[17676];
assign g[50443] = b[14] & g[17676];
assign g[34061] = a[14] & g[17677];
assign g[50444] = b[14] & g[17677];
assign g[34062] = a[14] & g[17678];
assign g[50445] = b[14] & g[17678];
assign g[34063] = a[14] & g[17679];
assign g[50446] = b[14] & g[17679];
assign g[34064] = a[14] & g[17680];
assign g[50447] = b[14] & g[17680];
assign g[34065] = a[14] & g[17681];
assign g[50448] = b[14] & g[17681];
assign g[34066] = a[14] & g[17682];
assign g[50449] = b[14] & g[17682];
assign g[34067] = a[14] & g[17683];
assign g[50450] = b[14] & g[17683];
assign g[34068] = a[14] & g[17684];
assign g[50451] = b[14] & g[17684];
assign g[34069] = a[14] & g[17685];
assign g[50452] = b[14] & g[17685];
assign g[34070] = a[14] & g[17686];
assign g[50453] = b[14] & g[17686];
assign g[34071] = a[14] & g[17687];
assign g[50454] = b[14] & g[17687];
assign g[34072] = a[14] & g[17688];
assign g[50455] = b[14] & g[17688];
assign g[34073] = a[14] & g[17689];
assign g[50456] = b[14] & g[17689];
assign g[34074] = a[14] & g[17690];
assign g[50457] = b[14] & g[17690];
assign g[34075] = a[14] & g[17691];
assign g[50458] = b[14] & g[17691];
assign g[34076] = a[14] & g[17692];
assign g[50459] = b[14] & g[17692];
assign g[34077] = a[14] & g[17693];
assign g[50460] = b[14] & g[17693];
assign g[34078] = a[14] & g[17694];
assign g[50461] = b[14] & g[17694];
assign g[34079] = a[14] & g[17695];
assign g[50462] = b[14] & g[17695];
assign g[34080] = a[14] & g[17696];
assign g[50463] = b[14] & g[17696];
assign g[34081] = a[14] & g[17697];
assign g[50464] = b[14] & g[17697];
assign g[34082] = a[14] & g[17698];
assign g[50465] = b[14] & g[17698];
assign g[34083] = a[14] & g[17699];
assign g[50466] = b[14] & g[17699];
assign g[34084] = a[14] & g[17700];
assign g[50467] = b[14] & g[17700];
assign g[34085] = a[14] & g[17701];
assign g[50468] = b[14] & g[17701];
assign g[34086] = a[14] & g[17702];
assign g[50469] = b[14] & g[17702];
assign g[34087] = a[14] & g[17703];
assign g[50470] = b[14] & g[17703];
assign g[34088] = a[14] & g[17704];
assign g[50471] = b[14] & g[17704];
assign g[34089] = a[14] & g[17705];
assign g[50472] = b[14] & g[17705];
assign g[34090] = a[14] & g[17706];
assign g[50473] = b[14] & g[17706];
assign g[34091] = a[14] & g[17707];
assign g[50474] = b[14] & g[17707];
assign g[34092] = a[14] & g[17708];
assign g[50475] = b[14] & g[17708];
assign g[34093] = a[14] & g[17709];
assign g[50476] = b[14] & g[17709];
assign g[34094] = a[14] & g[17710];
assign g[50477] = b[14] & g[17710];
assign g[34095] = a[14] & g[17711];
assign g[50478] = b[14] & g[17711];
assign g[34096] = a[14] & g[17712];
assign g[50479] = b[14] & g[17712];
assign g[34097] = a[14] & g[17713];
assign g[50480] = b[14] & g[17713];
assign g[34098] = a[14] & g[17714];
assign g[50481] = b[14] & g[17714];
assign g[34099] = a[14] & g[17715];
assign g[50482] = b[14] & g[17715];
assign g[34100] = a[14] & g[17716];
assign g[50483] = b[14] & g[17716];
assign g[34101] = a[14] & g[17717];
assign g[50484] = b[14] & g[17717];
assign g[34102] = a[14] & g[17718];
assign g[50485] = b[14] & g[17718];
assign g[34103] = a[14] & g[17719];
assign g[50486] = b[14] & g[17719];
assign g[34104] = a[14] & g[17720];
assign g[50487] = b[14] & g[17720];
assign g[34105] = a[14] & g[17721];
assign g[50488] = b[14] & g[17721];
assign g[34106] = a[14] & g[17722];
assign g[50489] = b[14] & g[17722];
assign g[34107] = a[14] & g[17723];
assign g[50490] = b[14] & g[17723];
assign g[34108] = a[14] & g[17724];
assign g[50491] = b[14] & g[17724];
assign g[34109] = a[14] & g[17725];
assign g[50492] = b[14] & g[17725];
assign g[34110] = a[14] & g[17726];
assign g[50493] = b[14] & g[17726];
assign g[34111] = a[14] & g[17727];
assign g[50494] = b[14] & g[17727];
assign g[34112] = a[14] & g[17728];
assign g[50495] = b[14] & g[17728];
assign g[34113] = a[14] & g[17729];
assign g[50496] = b[14] & g[17729];
assign g[34114] = a[14] & g[17730];
assign g[50497] = b[14] & g[17730];
assign g[34115] = a[14] & g[17731];
assign g[50498] = b[14] & g[17731];
assign g[34116] = a[14] & g[17732];
assign g[50499] = b[14] & g[17732];
assign g[34117] = a[14] & g[17733];
assign g[50500] = b[14] & g[17733];
assign g[34118] = a[14] & g[17734];
assign g[50501] = b[14] & g[17734];
assign g[34119] = a[14] & g[17735];
assign g[50502] = b[14] & g[17735];
assign g[34120] = a[14] & g[17736];
assign g[50503] = b[14] & g[17736];
assign g[34121] = a[14] & g[17737];
assign g[50504] = b[14] & g[17737];
assign g[34122] = a[14] & g[17738];
assign g[50505] = b[14] & g[17738];
assign g[34123] = a[14] & g[17739];
assign g[50506] = b[14] & g[17739];
assign g[34124] = a[14] & g[17740];
assign g[50507] = b[14] & g[17740];
assign g[34125] = a[14] & g[17741];
assign g[50508] = b[14] & g[17741];
assign g[34126] = a[14] & g[17742];
assign g[50509] = b[14] & g[17742];
assign g[34127] = a[14] & g[17743];
assign g[50510] = b[14] & g[17743];
assign g[34128] = a[14] & g[17744];
assign g[50511] = b[14] & g[17744];
assign g[34129] = a[14] & g[17745];
assign g[50512] = b[14] & g[17745];
assign g[34130] = a[14] & g[17746];
assign g[50513] = b[14] & g[17746];
assign g[34131] = a[14] & g[17747];
assign g[50514] = b[14] & g[17747];
assign g[34132] = a[14] & g[17748];
assign g[50515] = b[14] & g[17748];
assign g[34133] = a[14] & g[17749];
assign g[50516] = b[14] & g[17749];
assign g[34134] = a[14] & g[17750];
assign g[50517] = b[14] & g[17750];
assign g[34135] = a[14] & g[17751];
assign g[50518] = b[14] & g[17751];
assign g[34136] = a[14] & g[17752];
assign g[50519] = b[14] & g[17752];
assign g[34137] = a[14] & g[17753];
assign g[50520] = b[14] & g[17753];
assign g[34138] = a[14] & g[17754];
assign g[50521] = b[14] & g[17754];
assign g[34139] = a[14] & g[17755];
assign g[50522] = b[14] & g[17755];
assign g[34140] = a[14] & g[17756];
assign g[50523] = b[14] & g[17756];
assign g[34141] = a[14] & g[17757];
assign g[50524] = b[14] & g[17757];
assign g[34142] = a[14] & g[17758];
assign g[50525] = b[14] & g[17758];
assign g[34143] = a[14] & g[17759];
assign g[50526] = b[14] & g[17759];
assign g[34144] = a[14] & g[17760];
assign g[50527] = b[14] & g[17760];
assign g[34145] = a[14] & g[17761];
assign g[50528] = b[14] & g[17761];
assign g[34146] = a[14] & g[17762];
assign g[50529] = b[14] & g[17762];
assign g[34147] = a[14] & g[17763];
assign g[50530] = b[14] & g[17763];
assign g[34148] = a[14] & g[17764];
assign g[50531] = b[14] & g[17764];
assign g[34149] = a[14] & g[17765];
assign g[50532] = b[14] & g[17765];
assign g[34150] = a[14] & g[17766];
assign g[50533] = b[14] & g[17766];
assign g[34151] = a[14] & g[17767];
assign g[50534] = b[14] & g[17767];
assign g[34152] = a[14] & g[17768];
assign g[50535] = b[14] & g[17768];
assign g[34153] = a[14] & g[17769];
assign g[50536] = b[14] & g[17769];
assign g[34154] = a[14] & g[17770];
assign g[50537] = b[14] & g[17770];
assign g[34155] = a[14] & g[17771];
assign g[50538] = b[14] & g[17771];
assign g[34156] = a[14] & g[17772];
assign g[50539] = b[14] & g[17772];
assign g[34157] = a[14] & g[17773];
assign g[50540] = b[14] & g[17773];
assign g[34158] = a[14] & g[17774];
assign g[50541] = b[14] & g[17774];
assign g[34159] = a[14] & g[17775];
assign g[50542] = b[14] & g[17775];
assign g[34160] = a[14] & g[17776];
assign g[50543] = b[14] & g[17776];
assign g[34161] = a[14] & g[17777];
assign g[50544] = b[14] & g[17777];
assign g[34162] = a[14] & g[17778];
assign g[50545] = b[14] & g[17778];
assign g[34163] = a[14] & g[17779];
assign g[50546] = b[14] & g[17779];
assign g[34164] = a[14] & g[17780];
assign g[50547] = b[14] & g[17780];
assign g[34165] = a[14] & g[17781];
assign g[50548] = b[14] & g[17781];
assign g[34166] = a[14] & g[17782];
assign g[50549] = b[14] & g[17782];
assign g[34167] = a[14] & g[17783];
assign g[50550] = b[14] & g[17783];
assign g[34168] = a[14] & g[17784];
assign g[50551] = b[14] & g[17784];
assign g[34169] = a[14] & g[17785];
assign g[50552] = b[14] & g[17785];
assign g[34170] = a[14] & g[17786];
assign g[50553] = b[14] & g[17786];
assign g[34171] = a[14] & g[17787];
assign g[50554] = b[14] & g[17787];
assign g[34172] = a[14] & g[17788];
assign g[50555] = b[14] & g[17788];
assign g[34173] = a[14] & g[17789];
assign g[50556] = b[14] & g[17789];
assign g[34174] = a[14] & g[17790];
assign g[50557] = b[14] & g[17790];
assign g[34175] = a[14] & g[17791];
assign g[50558] = b[14] & g[17791];
assign g[34176] = a[14] & g[17792];
assign g[50559] = b[14] & g[17792];
assign g[34177] = a[14] & g[17793];
assign g[50560] = b[14] & g[17793];
assign g[34178] = a[14] & g[17794];
assign g[50561] = b[14] & g[17794];
assign g[34179] = a[14] & g[17795];
assign g[50562] = b[14] & g[17795];
assign g[34180] = a[14] & g[17796];
assign g[50563] = b[14] & g[17796];
assign g[34181] = a[14] & g[17797];
assign g[50564] = b[14] & g[17797];
assign g[34182] = a[14] & g[17798];
assign g[50565] = b[14] & g[17798];
assign g[34183] = a[14] & g[17799];
assign g[50566] = b[14] & g[17799];
assign g[34184] = a[14] & g[17800];
assign g[50567] = b[14] & g[17800];
assign g[34185] = a[14] & g[17801];
assign g[50568] = b[14] & g[17801];
assign g[34186] = a[14] & g[17802];
assign g[50569] = b[14] & g[17802];
assign g[34187] = a[14] & g[17803];
assign g[50570] = b[14] & g[17803];
assign g[34188] = a[14] & g[17804];
assign g[50571] = b[14] & g[17804];
assign g[34189] = a[14] & g[17805];
assign g[50572] = b[14] & g[17805];
assign g[34190] = a[14] & g[17806];
assign g[50573] = b[14] & g[17806];
assign g[34191] = a[14] & g[17807];
assign g[50574] = b[14] & g[17807];
assign g[34192] = a[14] & g[17808];
assign g[50575] = b[14] & g[17808];
assign g[34193] = a[14] & g[17809];
assign g[50576] = b[14] & g[17809];
assign g[34194] = a[14] & g[17810];
assign g[50577] = b[14] & g[17810];
assign g[34195] = a[14] & g[17811];
assign g[50578] = b[14] & g[17811];
assign g[34196] = a[14] & g[17812];
assign g[50579] = b[14] & g[17812];
assign g[34197] = a[14] & g[17813];
assign g[50580] = b[14] & g[17813];
assign g[34198] = a[14] & g[17814];
assign g[50581] = b[14] & g[17814];
assign g[34199] = a[14] & g[17815];
assign g[50582] = b[14] & g[17815];
assign g[34200] = a[14] & g[17816];
assign g[50583] = b[14] & g[17816];
assign g[34201] = a[14] & g[17817];
assign g[50584] = b[14] & g[17817];
assign g[34202] = a[14] & g[17818];
assign g[50585] = b[14] & g[17818];
assign g[34203] = a[14] & g[17819];
assign g[50586] = b[14] & g[17819];
assign g[34204] = a[14] & g[17820];
assign g[50587] = b[14] & g[17820];
assign g[34205] = a[14] & g[17821];
assign g[50588] = b[14] & g[17821];
assign g[34206] = a[14] & g[17822];
assign g[50589] = b[14] & g[17822];
assign g[34207] = a[14] & g[17823];
assign g[50590] = b[14] & g[17823];
assign g[34208] = a[14] & g[17824];
assign g[50591] = b[14] & g[17824];
assign g[34209] = a[14] & g[17825];
assign g[50592] = b[14] & g[17825];
assign g[34210] = a[14] & g[17826];
assign g[50593] = b[14] & g[17826];
assign g[34211] = a[14] & g[17827];
assign g[50594] = b[14] & g[17827];
assign g[34212] = a[14] & g[17828];
assign g[50595] = b[14] & g[17828];
assign g[34213] = a[14] & g[17829];
assign g[50596] = b[14] & g[17829];
assign g[34214] = a[14] & g[17830];
assign g[50597] = b[14] & g[17830];
assign g[34215] = a[14] & g[17831];
assign g[50598] = b[14] & g[17831];
assign g[34216] = a[14] & g[17832];
assign g[50599] = b[14] & g[17832];
assign g[34217] = a[14] & g[17833];
assign g[50600] = b[14] & g[17833];
assign g[34218] = a[14] & g[17834];
assign g[50601] = b[14] & g[17834];
assign g[34219] = a[14] & g[17835];
assign g[50602] = b[14] & g[17835];
assign g[34220] = a[14] & g[17836];
assign g[50603] = b[14] & g[17836];
assign g[34221] = a[14] & g[17837];
assign g[50604] = b[14] & g[17837];
assign g[34222] = a[14] & g[17838];
assign g[50605] = b[14] & g[17838];
assign g[34223] = a[14] & g[17839];
assign g[50606] = b[14] & g[17839];
assign g[34224] = a[14] & g[17840];
assign g[50607] = b[14] & g[17840];
assign g[34225] = a[14] & g[17841];
assign g[50608] = b[14] & g[17841];
assign g[34226] = a[14] & g[17842];
assign g[50609] = b[14] & g[17842];
assign g[34227] = a[14] & g[17843];
assign g[50610] = b[14] & g[17843];
assign g[34228] = a[14] & g[17844];
assign g[50611] = b[14] & g[17844];
assign g[34229] = a[14] & g[17845];
assign g[50612] = b[14] & g[17845];
assign g[34230] = a[14] & g[17846];
assign g[50613] = b[14] & g[17846];
assign g[34231] = a[14] & g[17847];
assign g[50614] = b[14] & g[17847];
assign g[34232] = a[14] & g[17848];
assign g[50615] = b[14] & g[17848];
assign g[34233] = a[14] & g[17849];
assign g[50616] = b[14] & g[17849];
assign g[34234] = a[14] & g[17850];
assign g[50617] = b[14] & g[17850];
assign g[34235] = a[14] & g[17851];
assign g[50618] = b[14] & g[17851];
assign g[34236] = a[14] & g[17852];
assign g[50619] = b[14] & g[17852];
assign g[34237] = a[14] & g[17853];
assign g[50620] = b[14] & g[17853];
assign g[34238] = a[14] & g[17854];
assign g[50621] = b[14] & g[17854];
assign g[34239] = a[14] & g[17855];
assign g[50622] = b[14] & g[17855];
assign g[34240] = a[14] & g[17856];
assign g[50623] = b[14] & g[17856];
assign g[34241] = a[14] & g[17857];
assign g[50624] = b[14] & g[17857];
assign g[34242] = a[14] & g[17858];
assign g[50625] = b[14] & g[17858];
assign g[34243] = a[14] & g[17859];
assign g[50626] = b[14] & g[17859];
assign g[34244] = a[14] & g[17860];
assign g[50627] = b[14] & g[17860];
assign g[34245] = a[14] & g[17861];
assign g[50628] = b[14] & g[17861];
assign g[34246] = a[14] & g[17862];
assign g[50629] = b[14] & g[17862];
assign g[34247] = a[14] & g[17863];
assign g[50630] = b[14] & g[17863];
assign g[34248] = a[14] & g[17864];
assign g[50631] = b[14] & g[17864];
assign g[34249] = a[14] & g[17865];
assign g[50632] = b[14] & g[17865];
assign g[34250] = a[14] & g[17866];
assign g[50633] = b[14] & g[17866];
assign g[34251] = a[14] & g[17867];
assign g[50634] = b[14] & g[17867];
assign g[34252] = a[14] & g[17868];
assign g[50635] = b[14] & g[17868];
assign g[34253] = a[14] & g[17869];
assign g[50636] = b[14] & g[17869];
assign g[34254] = a[14] & g[17870];
assign g[50637] = b[14] & g[17870];
assign g[34255] = a[14] & g[17871];
assign g[50638] = b[14] & g[17871];
assign g[34256] = a[14] & g[17872];
assign g[50639] = b[14] & g[17872];
assign g[34257] = a[14] & g[17873];
assign g[50640] = b[14] & g[17873];
assign g[34258] = a[14] & g[17874];
assign g[50641] = b[14] & g[17874];
assign g[34259] = a[14] & g[17875];
assign g[50642] = b[14] & g[17875];
assign g[34260] = a[14] & g[17876];
assign g[50643] = b[14] & g[17876];
assign g[34261] = a[14] & g[17877];
assign g[50644] = b[14] & g[17877];
assign g[34262] = a[14] & g[17878];
assign g[50645] = b[14] & g[17878];
assign g[34263] = a[14] & g[17879];
assign g[50646] = b[14] & g[17879];
assign g[34264] = a[14] & g[17880];
assign g[50647] = b[14] & g[17880];
assign g[34265] = a[14] & g[17881];
assign g[50648] = b[14] & g[17881];
assign g[34266] = a[14] & g[17882];
assign g[50649] = b[14] & g[17882];
assign g[34267] = a[14] & g[17883];
assign g[50650] = b[14] & g[17883];
assign g[34268] = a[14] & g[17884];
assign g[50651] = b[14] & g[17884];
assign g[34269] = a[14] & g[17885];
assign g[50652] = b[14] & g[17885];
assign g[34270] = a[14] & g[17886];
assign g[50653] = b[14] & g[17886];
assign g[34271] = a[14] & g[17887];
assign g[50654] = b[14] & g[17887];
assign g[34272] = a[14] & g[17888];
assign g[50655] = b[14] & g[17888];
assign g[34273] = a[14] & g[17889];
assign g[50656] = b[14] & g[17889];
assign g[34274] = a[14] & g[17890];
assign g[50657] = b[14] & g[17890];
assign g[34275] = a[14] & g[17891];
assign g[50658] = b[14] & g[17891];
assign g[34276] = a[14] & g[17892];
assign g[50659] = b[14] & g[17892];
assign g[34277] = a[14] & g[17893];
assign g[50660] = b[14] & g[17893];
assign g[34278] = a[14] & g[17894];
assign g[50661] = b[14] & g[17894];
assign g[34279] = a[14] & g[17895];
assign g[50662] = b[14] & g[17895];
assign g[34280] = a[14] & g[17896];
assign g[50663] = b[14] & g[17896];
assign g[34281] = a[14] & g[17897];
assign g[50664] = b[14] & g[17897];
assign g[34282] = a[14] & g[17898];
assign g[50665] = b[14] & g[17898];
assign g[34283] = a[14] & g[17899];
assign g[50666] = b[14] & g[17899];
assign g[34284] = a[14] & g[17900];
assign g[50667] = b[14] & g[17900];
assign g[34285] = a[14] & g[17901];
assign g[50668] = b[14] & g[17901];
assign g[34286] = a[14] & g[17902];
assign g[50669] = b[14] & g[17902];
assign g[34287] = a[14] & g[17903];
assign g[50670] = b[14] & g[17903];
assign g[34288] = a[14] & g[17904];
assign g[50671] = b[14] & g[17904];
assign g[34289] = a[14] & g[17905];
assign g[50672] = b[14] & g[17905];
assign g[34290] = a[14] & g[17906];
assign g[50673] = b[14] & g[17906];
assign g[34291] = a[14] & g[17907];
assign g[50674] = b[14] & g[17907];
assign g[34292] = a[14] & g[17908];
assign g[50675] = b[14] & g[17908];
assign g[34293] = a[14] & g[17909];
assign g[50676] = b[14] & g[17909];
assign g[34294] = a[14] & g[17910];
assign g[50677] = b[14] & g[17910];
assign g[34295] = a[14] & g[17911];
assign g[50678] = b[14] & g[17911];
assign g[34296] = a[14] & g[17912];
assign g[50679] = b[14] & g[17912];
assign g[34297] = a[14] & g[17913];
assign g[50680] = b[14] & g[17913];
assign g[34298] = a[14] & g[17914];
assign g[50681] = b[14] & g[17914];
assign g[34299] = a[14] & g[17915];
assign g[50682] = b[14] & g[17915];
assign g[34300] = a[14] & g[17916];
assign g[50683] = b[14] & g[17916];
assign g[34301] = a[14] & g[17917];
assign g[50684] = b[14] & g[17917];
assign g[34302] = a[14] & g[17918];
assign g[50685] = b[14] & g[17918];
assign g[34303] = a[14] & g[17919];
assign g[50686] = b[14] & g[17919];
assign g[34304] = a[14] & g[17920];
assign g[50687] = b[14] & g[17920];
assign g[34305] = a[14] & g[17921];
assign g[50688] = b[14] & g[17921];
assign g[34306] = a[14] & g[17922];
assign g[50689] = b[14] & g[17922];
assign g[34307] = a[14] & g[17923];
assign g[50690] = b[14] & g[17923];
assign g[34308] = a[14] & g[17924];
assign g[50691] = b[14] & g[17924];
assign g[34309] = a[14] & g[17925];
assign g[50692] = b[14] & g[17925];
assign g[34310] = a[14] & g[17926];
assign g[50693] = b[14] & g[17926];
assign g[34311] = a[14] & g[17927];
assign g[50694] = b[14] & g[17927];
assign g[34312] = a[14] & g[17928];
assign g[50695] = b[14] & g[17928];
assign g[34313] = a[14] & g[17929];
assign g[50696] = b[14] & g[17929];
assign g[34314] = a[14] & g[17930];
assign g[50697] = b[14] & g[17930];
assign g[34315] = a[14] & g[17931];
assign g[50698] = b[14] & g[17931];
assign g[34316] = a[14] & g[17932];
assign g[50699] = b[14] & g[17932];
assign g[34317] = a[14] & g[17933];
assign g[50700] = b[14] & g[17933];
assign g[34318] = a[14] & g[17934];
assign g[50701] = b[14] & g[17934];
assign g[34319] = a[14] & g[17935];
assign g[50702] = b[14] & g[17935];
assign g[34320] = a[14] & g[17936];
assign g[50703] = b[14] & g[17936];
assign g[34321] = a[14] & g[17937];
assign g[50704] = b[14] & g[17937];
assign g[34322] = a[14] & g[17938];
assign g[50705] = b[14] & g[17938];
assign g[34323] = a[14] & g[17939];
assign g[50706] = b[14] & g[17939];
assign g[34324] = a[14] & g[17940];
assign g[50707] = b[14] & g[17940];
assign g[34325] = a[14] & g[17941];
assign g[50708] = b[14] & g[17941];
assign g[34326] = a[14] & g[17942];
assign g[50709] = b[14] & g[17942];
assign g[34327] = a[14] & g[17943];
assign g[50710] = b[14] & g[17943];
assign g[34328] = a[14] & g[17944];
assign g[50711] = b[14] & g[17944];
assign g[34329] = a[14] & g[17945];
assign g[50712] = b[14] & g[17945];
assign g[34330] = a[14] & g[17946];
assign g[50713] = b[14] & g[17946];
assign g[34331] = a[14] & g[17947];
assign g[50714] = b[14] & g[17947];
assign g[34332] = a[14] & g[17948];
assign g[50715] = b[14] & g[17948];
assign g[34333] = a[14] & g[17949];
assign g[50716] = b[14] & g[17949];
assign g[34334] = a[14] & g[17950];
assign g[50717] = b[14] & g[17950];
assign g[34335] = a[14] & g[17951];
assign g[50718] = b[14] & g[17951];
assign g[34336] = a[14] & g[17952];
assign g[50719] = b[14] & g[17952];
assign g[34337] = a[14] & g[17953];
assign g[50720] = b[14] & g[17953];
assign g[34338] = a[14] & g[17954];
assign g[50721] = b[14] & g[17954];
assign g[34339] = a[14] & g[17955];
assign g[50722] = b[14] & g[17955];
assign g[34340] = a[14] & g[17956];
assign g[50723] = b[14] & g[17956];
assign g[34341] = a[14] & g[17957];
assign g[50724] = b[14] & g[17957];
assign g[34342] = a[14] & g[17958];
assign g[50725] = b[14] & g[17958];
assign g[34343] = a[14] & g[17959];
assign g[50726] = b[14] & g[17959];
assign g[34344] = a[14] & g[17960];
assign g[50727] = b[14] & g[17960];
assign g[34345] = a[14] & g[17961];
assign g[50728] = b[14] & g[17961];
assign g[34346] = a[14] & g[17962];
assign g[50729] = b[14] & g[17962];
assign g[34347] = a[14] & g[17963];
assign g[50730] = b[14] & g[17963];
assign g[34348] = a[14] & g[17964];
assign g[50731] = b[14] & g[17964];
assign g[34349] = a[14] & g[17965];
assign g[50732] = b[14] & g[17965];
assign g[34350] = a[14] & g[17966];
assign g[50733] = b[14] & g[17966];
assign g[34351] = a[14] & g[17967];
assign g[50734] = b[14] & g[17967];
assign g[34352] = a[14] & g[17968];
assign g[50735] = b[14] & g[17968];
assign g[34353] = a[14] & g[17969];
assign g[50736] = b[14] & g[17969];
assign g[34354] = a[14] & g[17970];
assign g[50737] = b[14] & g[17970];
assign g[34355] = a[14] & g[17971];
assign g[50738] = b[14] & g[17971];
assign g[34356] = a[14] & g[17972];
assign g[50739] = b[14] & g[17972];
assign g[34357] = a[14] & g[17973];
assign g[50740] = b[14] & g[17973];
assign g[34358] = a[14] & g[17974];
assign g[50741] = b[14] & g[17974];
assign g[34359] = a[14] & g[17975];
assign g[50742] = b[14] & g[17975];
assign g[34360] = a[14] & g[17976];
assign g[50743] = b[14] & g[17976];
assign g[34361] = a[14] & g[17977];
assign g[50744] = b[14] & g[17977];
assign g[34362] = a[14] & g[17978];
assign g[50745] = b[14] & g[17978];
assign g[34363] = a[14] & g[17979];
assign g[50746] = b[14] & g[17979];
assign g[34364] = a[14] & g[17980];
assign g[50747] = b[14] & g[17980];
assign g[34365] = a[14] & g[17981];
assign g[50748] = b[14] & g[17981];
assign g[34366] = a[14] & g[17982];
assign g[50749] = b[14] & g[17982];
assign g[34367] = a[14] & g[17983];
assign g[50750] = b[14] & g[17983];
assign g[34368] = a[14] & g[17984];
assign g[50751] = b[14] & g[17984];
assign g[34369] = a[14] & g[17985];
assign g[50752] = b[14] & g[17985];
assign g[34370] = a[14] & g[17986];
assign g[50753] = b[14] & g[17986];
assign g[34371] = a[14] & g[17987];
assign g[50754] = b[14] & g[17987];
assign g[34372] = a[14] & g[17988];
assign g[50755] = b[14] & g[17988];
assign g[34373] = a[14] & g[17989];
assign g[50756] = b[14] & g[17989];
assign g[34374] = a[14] & g[17990];
assign g[50757] = b[14] & g[17990];
assign g[34375] = a[14] & g[17991];
assign g[50758] = b[14] & g[17991];
assign g[34376] = a[14] & g[17992];
assign g[50759] = b[14] & g[17992];
assign g[34377] = a[14] & g[17993];
assign g[50760] = b[14] & g[17993];
assign g[34378] = a[14] & g[17994];
assign g[50761] = b[14] & g[17994];
assign g[34379] = a[14] & g[17995];
assign g[50762] = b[14] & g[17995];
assign g[34380] = a[14] & g[17996];
assign g[50763] = b[14] & g[17996];
assign g[34381] = a[14] & g[17997];
assign g[50764] = b[14] & g[17997];
assign g[34382] = a[14] & g[17998];
assign g[50765] = b[14] & g[17998];
assign g[34383] = a[14] & g[17999];
assign g[50766] = b[14] & g[17999];
assign g[34384] = a[14] & g[18000];
assign g[50767] = b[14] & g[18000];
assign g[34385] = a[14] & g[18001];
assign g[50768] = b[14] & g[18001];
assign g[34386] = a[14] & g[18002];
assign g[50769] = b[14] & g[18002];
assign g[34387] = a[14] & g[18003];
assign g[50770] = b[14] & g[18003];
assign g[34388] = a[14] & g[18004];
assign g[50771] = b[14] & g[18004];
assign g[34389] = a[14] & g[18005];
assign g[50772] = b[14] & g[18005];
assign g[34390] = a[14] & g[18006];
assign g[50773] = b[14] & g[18006];
assign g[34391] = a[14] & g[18007];
assign g[50774] = b[14] & g[18007];
assign g[34392] = a[14] & g[18008];
assign g[50775] = b[14] & g[18008];
assign g[34393] = a[14] & g[18009];
assign g[50776] = b[14] & g[18009];
assign g[34394] = a[14] & g[18010];
assign g[50777] = b[14] & g[18010];
assign g[34395] = a[14] & g[18011];
assign g[50778] = b[14] & g[18011];
assign g[34396] = a[14] & g[18012];
assign g[50779] = b[14] & g[18012];
assign g[34397] = a[14] & g[18013];
assign g[50780] = b[14] & g[18013];
assign g[34398] = a[14] & g[18014];
assign g[50781] = b[14] & g[18014];
assign g[34399] = a[14] & g[18015];
assign g[50782] = b[14] & g[18015];
assign g[34400] = a[14] & g[18016];
assign g[50783] = b[14] & g[18016];
assign g[34401] = a[14] & g[18017];
assign g[50784] = b[14] & g[18017];
assign g[34402] = a[14] & g[18018];
assign g[50785] = b[14] & g[18018];
assign g[34403] = a[14] & g[18019];
assign g[50786] = b[14] & g[18019];
assign g[34404] = a[14] & g[18020];
assign g[50787] = b[14] & g[18020];
assign g[34405] = a[14] & g[18021];
assign g[50788] = b[14] & g[18021];
assign g[34406] = a[14] & g[18022];
assign g[50789] = b[14] & g[18022];
assign g[34407] = a[14] & g[18023];
assign g[50790] = b[14] & g[18023];
assign g[34408] = a[14] & g[18024];
assign g[50791] = b[14] & g[18024];
assign g[34409] = a[14] & g[18025];
assign g[50792] = b[14] & g[18025];
assign g[34410] = a[14] & g[18026];
assign g[50793] = b[14] & g[18026];
assign g[34411] = a[14] & g[18027];
assign g[50794] = b[14] & g[18027];
assign g[34412] = a[14] & g[18028];
assign g[50795] = b[14] & g[18028];
assign g[34413] = a[14] & g[18029];
assign g[50796] = b[14] & g[18029];
assign g[34414] = a[14] & g[18030];
assign g[50797] = b[14] & g[18030];
assign g[34415] = a[14] & g[18031];
assign g[50798] = b[14] & g[18031];
assign g[34416] = a[14] & g[18032];
assign g[50799] = b[14] & g[18032];
assign g[34417] = a[14] & g[18033];
assign g[50800] = b[14] & g[18033];
assign g[34418] = a[14] & g[18034];
assign g[50801] = b[14] & g[18034];
assign g[34419] = a[14] & g[18035];
assign g[50802] = b[14] & g[18035];
assign g[34420] = a[14] & g[18036];
assign g[50803] = b[14] & g[18036];
assign g[34421] = a[14] & g[18037];
assign g[50804] = b[14] & g[18037];
assign g[34422] = a[14] & g[18038];
assign g[50805] = b[14] & g[18038];
assign g[34423] = a[14] & g[18039];
assign g[50806] = b[14] & g[18039];
assign g[34424] = a[14] & g[18040];
assign g[50807] = b[14] & g[18040];
assign g[34425] = a[14] & g[18041];
assign g[50808] = b[14] & g[18041];
assign g[34426] = a[14] & g[18042];
assign g[50809] = b[14] & g[18042];
assign g[34427] = a[14] & g[18043];
assign g[50810] = b[14] & g[18043];
assign g[34428] = a[14] & g[18044];
assign g[50811] = b[14] & g[18044];
assign g[34429] = a[14] & g[18045];
assign g[50812] = b[14] & g[18045];
assign g[34430] = a[14] & g[18046];
assign g[50813] = b[14] & g[18046];
assign g[34431] = a[14] & g[18047];
assign g[50814] = b[14] & g[18047];
assign g[34432] = a[14] & g[18048];
assign g[50815] = b[14] & g[18048];
assign g[34433] = a[14] & g[18049];
assign g[50816] = b[14] & g[18049];
assign g[34434] = a[14] & g[18050];
assign g[50817] = b[14] & g[18050];
assign g[34435] = a[14] & g[18051];
assign g[50818] = b[14] & g[18051];
assign g[34436] = a[14] & g[18052];
assign g[50819] = b[14] & g[18052];
assign g[34437] = a[14] & g[18053];
assign g[50820] = b[14] & g[18053];
assign g[34438] = a[14] & g[18054];
assign g[50821] = b[14] & g[18054];
assign g[34439] = a[14] & g[18055];
assign g[50822] = b[14] & g[18055];
assign g[34440] = a[14] & g[18056];
assign g[50823] = b[14] & g[18056];
assign g[34441] = a[14] & g[18057];
assign g[50824] = b[14] & g[18057];
assign g[34442] = a[14] & g[18058];
assign g[50825] = b[14] & g[18058];
assign g[34443] = a[14] & g[18059];
assign g[50826] = b[14] & g[18059];
assign g[34444] = a[14] & g[18060];
assign g[50827] = b[14] & g[18060];
assign g[34445] = a[14] & g[18061];
assign g[50828] = b[14] & g[18061];
assign g[34446] = a[14] & g[18062];
assign g[50829] = b[14] & g[18062];
assign g[34447] = a[14] & g[18063];
assign g[50830] = b[14] & g[18063];
assign g[34448] = a[14] & g[18064];
assign g[50831] = b[14] & g[18064];
assign g[34449] = a[14] & g[18065];
assign g[50832] = b[14] & g[18065];
assign g[34450] = a[14] & g[18066];
assign g[50833] = b[14] & g[18066];
assign g[34451] = a[14] & g[18067];
assign g[50834] = b[14] & g[18067];
assign g[34452] = a[14] & g[18068];
assign g[50835] = b[14] & g[18068];
assign g[34453] = a[14] & g[18069];
assign g[50836] = b[14] & g[18069];
assign g[34454] = a[14] & g[18070];
assign g[50837] = b[14] & g[18070];
assign g[34455] = a[14] & g[18071];
assign g[50838] = b[14] & g[18071];
assign g[34456] = a[14] & g[18072];
assign g[50839] = b[14] & g[18072];
assign g[34457] = a[14] & g[18073];
assign g[50840] = b[14] & g[18073];
assign g[34458] = a[14] & g[18074];
assign g[50841] = b[14] & g[18074];
assign g[34459] = a[14] & g[18075];
assign g[50842] = b[14] & g[18075];
assign g[34460] = a[14] & g[18076];
assign g[50843] = b[14] & g[18076];
assign g[34461] = a[14] & g[18077];
assign g[50844] = b[14] & g[18077];
assign g[34462] = a[14] & g[18078];
assign g[50845] = b[14] & g[18078];
assign g[34463] = a[14] & g[18079];
assign g[50846] = b[14] & g[18079];
assign g[34464] = a[14] & g[18080];
assign g[50847] = b[14] & g[18080];
assign g[34465] = a[14] & g[18081];
assign g[50848] = b[14] & g[18081];
assign g[34466] = a[14] & g[18082];
assign g[50849] = b[14] & g[18082];
assign g[34467] = a[14] & g[18083];
assign g[50850] = b[14] & g[18083];
assign g[34468] = a[14] & g[18084];
assign g[50851] = b[14] & g[18084];
assign g[34469] = a[14] & g[18085];
assign g[50852] = b[14] & g[18085];
assign g[34470] = a[14] & g[18086];
assign g[50853] = b[14] & g[18086];
assign g[34471] = a[14] & g[18087];
assign g[50854] = b[14] & g[18087];
assign g[34472] = a[14] & g[18088];
assign g[50855] = b[14] & g[18088];
assign g[34473] = a[14] & g[18089];
assign g[50856] = b[14] & g[18089];
assign g[34474] = a[14] & g[18090];
assign g[50857] = b[14] & g[18090];
assign g[34475] = a[14] & g[18091];
assign g[50858] = b[14] & g[18091];
assign g[34476] = a[14] & g[18092];
assign g[50859] = b[14] & g[18092];
assign g[34477] = a[14] & g[18093];
assign g[50860] = b[14] & g[18093];
assign g[34478] = a[14] & g[18094];
assign g[50861] = b[14] & g[18094];
assign g[34479] = a[14] & g[18095];
assign g[50862] = b[14] & g[18095];
assign g[34480] = a[14] & g[18096];
assign g[50863] = b[14] & g[18096];
assign g[34481] = a[14] & g[18097];
assign g[50864] = b[14] & g[18097];
assign g[34482] = a[14] & g[18098];
assign g[50865] = b[14] & g[18098];
assign g[34483] = a[14] & g[18099];
assign g[50866] = b[14] & g[18099];
assign g[34484] = a[14] & g[18100];
assign g[50867] = b[14] & g[18100];
assign g[34485] = a[14] & g[18101];
assign g[50868] = b[14] & g[18101];
assign g[34486] = a[14] & g[18102];
assign g[50869] = b[14] & g[18102];
assign g[34487] = a[14] & g[18103];
assign g[50870] = b[14] & g[18103];
assign g[34488] = a[14] & g[18104];
assign g[50871] = b[14] & g[18104];
assign g[34489] = a[14] & g[18105];
assign g[50872] = b[14] & g[18105];
assign g[34490] = a[14] & g[18106];
assign g[50873] = b[14] & g[18106];
assign g[34491] = a[14] & g[18107];
assign g[50874] = b[14] & g[18107];
assign g[34492] = a[14] & g[18108];
assign g[50875] = b[14] & g[18108];
assign g[34493] = a[14] & g[18109];
assign g[50876] = b[14] & g[18109];
assign g[34494] = a[14] & g[18110];
assign g[50877] = b[14] & g[18110];
assign g[34495] = a[14] & g[18111];
assign g[50878] = b[14] & g[18111];
assign g[34496] = a[14] & g[18112];
assign g[50879] = b[14] & g[18112];
assign g[34497] = a[14] & g[18113];
assign g[50880] = b[14] & g[18113];
assign g[34498] = a[14] & g[18114];
assign g[50881] = b[14] & g[18114];
assign g[34499] = a[14] & g[18115];
assign g[50882] = b[14] & g[18115];
assign g[34500] = a[14] & g[18116];
assign g[50883] = b[14] & g[18116];
assign g[34501] = a[14] & g[18117];
assign g[50884] = b[14] & g[18117];
assign g[34502] = a[14] & g[18118];
assign g[50885] = b[14] & g[18118];
assign g[34503] = a[14] & g[18119];
assign g[50886] = b[14] & g[18119];
assign g[34504] = a[14] & g[18120];
assign g[50887] = b[14] & g[18120];
assign g[34505] = a[14] & g[18121];
assign g[50888] = b[14] & g[18121];
assign g[34506] = a[14] & g[18122];
assign g[50889] = b[14] & g[18122];
assign g[34507] = a[14] & g[18123];
assign g[50890] = b[14] & g[18123];
assign g[34508] = a[14] & g[18124];
assign g[50891] = b[14] & g[18124];
assign g[34509] = a[14] & g[18125];
assign g[50892] = b[14] & g[18125];
assign g[34510] = a[14] & g[18126];
assign g[50893] = b[14] & g[18126];
assign g[34511] = a[14] & g[18127];
assign g[50894] = b[14] & g[18127];
assign g[34512] = a[14] & g[18128];
assign g[50895] = b[14] & g[18128];
assign g[34513] = a[14] & g[18129];
assign g[50896] = b[14] & g[18129];
assign g[34514] = a[14] & g[18130];
assign g[50897] = b[14] & g[18130];
assign g[34515] = a[14] & g[18131];
assign g[50898] = b[14] & g[18131];
assign g[34516] = a[14] & g[18132];
assign g[50899] = b[14] & g[18132];
assign g[34517] = a[14] & g[18133];
assign g[50900] = b[14] & g[18133];
assign g[34518] = a[14] & g[18134];
assign g[50901] = b[14] & g[18134];
assign g[34519] = a[14] & g[18135];
assign g[50902] = b[14] & g[18135];
assign g[34520] = a[14] & g[18136];
assign g[50903] = b[14] & g[18136];
assign g[34521] = a[14] & g[18137];
assign g[50904] = b[14] & g[18137];
assign g[34522] = a[14] & g[18138];
assign g[50905] = b[14] & g[18138];
assign g[34523] = a[14] & g[18139];
assign g[50906] = b[14] & g[18139];
assign g[34524] = a[14] & g[18140];
assign g[50907] = b[14] & g[18140];
assign g[34525] = a[14] & g[18141];
assign g[50908] = b[14] & g[18141];
assign g[34526] = a[14] & g[18142];
assign g[50909] = b[14] & g[18142];
assign g[34527] = a[14] & g[18143];
assign g[50910] = b[14] & g[18143];
assign g[34528] = a[14] & g[18144];
assign g[50911] = b[14] & g[18144];
assign g[34529] = a[14] & g[18145];
assign g[50912] = b[14] & g[18145];
assign g[34530] = a[14] & g[18146];
assign g[50913] = b[14] & g[18146];
assign g[34531] = a[14] & g[18147];
assign g[50914] = b[14] & g[18147];
assign g[34532] = a[14] & g[18148];
assign g[50915] = b[14] & g[18148];
assign g[34533] = a[14] & g[18149];
assign g[50916] = b[14] & g[18149];
assign g[34534] = a[14] & g[18150];
assign g[50917] = b[14] & g[18150];
assign g[34535] = a[14] & g[18151];
assign g[50918] = b[14] & g[18151];
assign g[34536] = a[14] & g[18152];
assign g[50919] = b[14] & g[18152];
assign g[34537] = a[14] & g[18153];
assign g[50920] = b[14] & g[18153];
assign g[34538] = a[14] & g[18154];
assign g[50921] = b[14] & g[18154];
assign g[34539] = a[14] & g[18155];
assign g[50922] = b[14] & g[18155];
assign g[34540] = a[14] & g[18156];
assign g[50923] = b[14] & g[18156];
assign g[34541] = a[14] & g[18157];
assign g[50924] = b[14] & g[18157];
assign g[34542] = a[14] & g[18158];
assign g[50925] = b[14] & g[18158];
assign g[34543] = a[14] & g[18159];
assign g[50926] = b[14] & g[18159];
assign g[34544] = a[14] & g[18160];
assign g[50927] = b[14] & g[18160];
assign g[34545] = a[14] & g[18161];
assign g[50928] = b[14] & g[18161];
assign g[34546] = a[14] & g[18162];
assign g[50929] = b[14] & g[18162];
assign g[34547] = a[14] & g[18163];
assign g[50930] = b[14] & g[18163];
assign g[34548] = a[14] & g[18164];
assign g[50931] = b[14] & g[18164];
assign g[34549] = a[14] & g[18165];
assign g[50932] = b[14] & g[18165];
assign g[34550] = a[14] & g[18166];
assign g[50933] = b[14] & g[18166];
assign g[34551] = a[14] & g[18167];
assign g[50934] = b[14] & g[18167];
assign g[34552] = a[14] & g[18168];
assign g[50935] = b[14] & g[18168];
assign g[34553] = a[14] & g[18169];
assign g[50936] = b[14] & g[18169];
assign g[34554] = a[14] & g[18170];
assign g[50937] = b[14] & g[18170];
assign g[34555] = a[14] & g[18171];
assign g[50938] = b[14] & g[18171];
assign g[34556] = a[14] & g[18172];
assign g[50939] = b[14] & g[18172];
assign g[34557] = a[14] & g[18173];
assign g[50940] = b[14] & g[18173];
assign g[34558] = a[14] & g[18174];
assign g[50941] = b[14] & g[18174];
assign g[34559] = a[14] & g[18175];
assign g[50942] = b[14] & g[18175];
assign g[34560] = a[14] & g[18176];
assign g[50943] = b[14] & g[18176];
assign g[34561] = a[14] & g[18177];
assign g[50944] = b[14] & g[18177];
assign g[34562] = a[14] & g[18178];
assign g[50945] = b[14] & g[18178];
assign g[34563] = a[14] & g[18179];
assign g[50946] = b[14] & g[18179];
assign g[34564] = a[14] & g[18180];
assign g[50947] = b[14] & g[18180];
assign g[34565] = a[14] & g[18181];
assign g[50948] = b[14] & g[18181];
assign g[34566] = a[14] & g[18182];
assign g[50949] = b[14] & g[18182];
assign g[34567] = a[14] & g[18183];
assign g[50950] = b[14] & g[18183];
assign g[34568] = a[14] & g[18184];
assign g[50951] = b[14] & g[18184];
assign g[34569] = a[14] & g[18185];
assign g[50952] = b[14] & g[18185];
assign g[34570] = a[14] & g[18186];
assign g[50953] = b[14] & g[18186];
assign g[34571] = a[14] & g[18187];
assign g[50954] = b[14] & g[18187];
assign g[34572] = a[14] & g[18188];
assign g[50955] = b[14] & g[18188];
assign g[34573] = a[14] & g[18189];
assign g[50956] = b[14] & g[18189];
assign g[34574] = a[14] & g[18190];
assign g[50957] = b[14] & g[18190];
assign g[34575] = a[14] & g[18191];
assign g[50958] = b[14] & g[18191];
assign g[34576] = a[14] & g[18192];
assign g[50959] = b[14] & g[18192];
assign g[34577] = a[14] & g[18193];
assign g[50960] = b[14] & g[18193];
assign g[34578] = a[14] & g[18194];
assign g[50961] = b[14] & g[18194];
assign g[34579] = a[14] & g[18195];
assign g[50962] = b[14] & g[18195];
assign g[34580] = a[14] & g[18196];
assign g[50963] = b[14] & g[18196];
assign g[34581] = a[14] & g[18197];
assign g[50964] = b[14] & g[18197];
assign g[34582] = a[14] & g[18198];
assign g[50965] = b[14] & g[18198];
assign g[34583] = a[14] & g[18199];
assign g[50966] = b[14] & g[18199];
assign g[34584] = a[14] & g[18200];
assign g[50967] = b[14] & g[18200];
assign g[34585] = a[14] & g[18201];
assign g[50968] = b[14] & g[18201];
assign g[34586] = a[14] & g[18202];
assign g[50969] = b[14] & g[18202];
assign g[34587] = a[14] & g[18203];
assign g[50970] = b[14] & g[18203];
assign g[34588] = a[14] & g[18204];
assign g[50971] = b[14] & g[18204];
assign g[34589] = a[14] & g[18205];
assign g[50972] = b[14] & g[18205];
assign g[34590] = a[14] & g[18206];
assign g[50973] = b[14] & g[18206];
assign g[34591] = a[14] & g[18207];
assign g[50974] = b[14] & g[18207];
assign g[34592] = a[14] & g[18208];
assign g[50975] = b[14] & g[18208];
assign g[34593] = a[14] & g[18209];
assign g[50976] = b[14] & g[18209];
assign g[34594] = a[14] & g[18210];
assign g[50977] = b[14] & g[18210];
assign g[34595] = a[14] & g[18211];
assign g[50978] = b[14] & g[18211];
assign g[34596] = a[14] & g[18212];
assign g[50979] = b[14] & g[18212];
assign g[34597] = a[14] & g[18213];
assign g[50980] = b[14] & g[18213];
assign g[34598] = a[14] & g[18214];
assign g[50981] = b[14] & g[18214];
assign g[34599] = a[14] & g[18215];
assign g[50982] = b[14] & g[18215];
assign g[34600] = a[14] & g[18216];
assign g[50983] = b[14] & g[18216];
assign g[34601] = a[14] & g[18217];
assign g[50984] = b[14] & g[18217];
assign g[34602] = a[14] & g[18218];
assign g[50985] = b[14] & g[18218];
assign g[34603] = a[14] & g[18219];
assign g[50986] = b[14] & g[18219];
assign g[34604] = a[14] & g[18220];
assign g[50987] = b[14] & g[18220];
assign g[34605] = a[14] & g[18221];
assign g[50988] = b[14] & g[18221];
assign g[34606] = a[14] & g[18222];
assign g[50989] = b[14] & g[18222];
assign g[34607] = a[14] & g[18223];
assign g[50990] = b[14] & g[18223];
assign g[34608] = a[14] & g[18224];
assign g[50991] = b[14] & g[18224];
assign g[34609] = a[14] & g[18225];
assign g[50992] = b[14] & g[18225];
assign g[34610] = a[14] & g[18226];
assign g[50993] = b[14] & g[18226];
assign g[34611] = a[14] & g[18227];
assign g[50994] = b[14] & g[18227];
assign g[34612] = a[14] & g[18228];
assign g[50995] = b[14] & g[18228];
assign g[34613] = a[14] & g[18229];
assign g[50996] = b[14] & g[18229];
assign g[34614] = a[14] & g[18230];
assign g[50997] = b[14] & g[18230];
assign g[34615] = a[14] & g[18231];
assign g[50998] = b[14] & g[18231];
assign g[34616] = a[14] & g[18232];
assign g[50999] = b[14] & g[18232];
assign g[34617] = a[14] & g[18233];
assign g[51000] = b[14] & g[18233];
assign g[34618] = a[14] & g[18234];
assign g[51001] = b[14] & g[18234];
assign g[34619] = a[14] & g[18235];
assign g[51002] = b[14] & g[18235];
assign g[34620] = a[14] & g[18236];
assign g[51003] = b[14] & g[18236];
assign g[34621] = a[14] & g[18237];
assign g[51004] = b[14] & g[18237];
assign g[34622] = a[14] & g[18238];
assign g[51005] = b[14] & g[18238];
assign g[34623] = a[14] & g[18239];
assign g[51006] = b[14] & g[18239];
assign g[34624] = a[14] & g[18240];
assign g[51007] = b[14] & g[18240];
assign g[34625] = a[14] & g[18241];
assign g[51008] = b[14] & g[18241];
assign g[34626] = a[14] & g[18242];
assign g[51009] = b[14] & g[18242];
assign g[34627] = a[14] & g[18243];
assign g[51010] = b[14] & g[18243];
assign g[34628] = a[14] & g[18244];
assign g[51011] = b[14] & g[18244];
assign g[34629] = a[14] & g[18245];
assign g[51012] = b[14] & g[18245];
assign g[34630] = a[14] & g[18246];
assign g[51013] = b[14] & g[18246];
assign g[34631] = a[14] & g[18247];
assign g[51014] = b[14] & g[18247];
assign g[34632] = a[14] & g[18248];
assign g[51015] = b[14] & g[18248];
assign g[34633] = a[14] & g[18249];
assign g[51016] = b[14] & g[18249];
assign g[34634] = a[14] & g[18250];
assign g[51017] = b[14] & g[18250];
assign g[34635] = a[14] & g[18251];
assign g[51018] = b[14] & g[18251];
assign g[34636] = a[14] & g[18252];
assign g[51019] = b[14] & g[18252];
assign g[34637] = a[14] & g[18253];
assign g[51020] = b[14] & g[18253];
assign g[34638] = a[14] & g[18254];
assign g[51021] = b[14] & g[18254];
assign g[34639] = a[14] & g[18255];
assign g[51022] = b[14] & g[18255];
assign g[34640] = a[14] & g[18256];
assign g[51023] = b[14] & g[18256];
assign g[34641] = a[14] & g[18257];
assign g[51024] = b[14] & g[18257];
assign g[34642] = a[14] & g[18258];
assign g[51025] = b[14] & g[18258];
assign g[34643] = a[14] & g[18259];
assign g[51026] = b[14] & g[18259];
assign g[34644] = a[14] & g[18260];
assign g[51027] = b[14] & g[18260];
assign g[34645] = a[14] & g[18261];
assign g[51028] = b[14] & g[18261];
assign g[34646] = a[14] & g[18262];
assign g[51029] = b[14] & g[18262];
assign g[34647] = a[14] & g[18263];
assign g[51030] = b[14] & g[18263];
assign g[34648] = a[14] & g[18264];
assign g[51031] = b[14] & g[18264];
assign g[34649] = a[14] & g[18265];
assign g[51032] = b[14] & g[18265];
assign g[34650] = a[14] & g[18266];
assign g[51033] = b[14] & g[18266];
assign g[34651] = a[14] & g[18267];
assign g[51034] = b[14] & g[18267];
assign g[34652] = a[14] & g[18268];
assign g[51035] = b[14] & g[18268];
assign g[34653] = a[14] & g[18269];
assign g[51036] = b[14] & g[18269];
assign g[34654] = a[14] & g[18270];
assign g[51037] = b[14] & g[18270];
assign g[34655] = a[14] & g[18271];
assign g[51038] = b[14] & g[18271];
assign g[34656] = a[14] & g[18272];
assign g[51039] = b[14] & g[18272];
assign g[34657] = a[14] & g[18273];
assign g[51040] = b[14] & g[18273];
assign g[34658] = a[14] & g[18274];
assign g[51041] = b[14] & g[18274];
assign g[34659] = a[14] & g[18275];
assign g[51042] = b[14] & g[18275];
assign g[34660] = a[14] & g[18276];
assign g[51043] = b[14] & g[18276];
assign g[34661] = a[14] & g[18277];
assign g[51044] = b[14] & g[18277];
assign g[34662] = a[14] & g[18278];
assign g[51045] = b[14] & g[18278];
assign g[34663] = a[14] & g[18279];
assign g[51046] = b[14] & g[18279];
assign g[34664] = a[14] & g[18280];
assign g[51047] = b[14] & g[18280];
assign g[34665] = a[14] & g[18281];
assign g[51048] = b[14] & g[18281];
assign g[34666] = a[14] & g[18282];
assign g[51049] = b[14] & g[18282];
assign g[34667] = a[14] & g[18283];
assign g[51050] = b[14] & g[18283];
assign g[34668] = a[14] & g[18284];
assign g[51051] = b[14] & g[18284];
assign g[34669] = a[14] & g[18285];
assign g[51052] = b[14] & g[18285];
assign g[34670] = a[14] & g[18286];
assign g[51053] = b[14] & g[18286];
assign g[34671] = a[14] & g[18287];
assign g[51054] = b[14] & g[18287];
assign g[34672] = a[14] & g[18288];
assign g[51055] = b[14] & g[18288];
assign g[34673] = a[14] & g[18289];
assign g[51056] = b[14] & g[18289];
assign g[34674] = a[14] & g[18290];
assign g[51057] = b[14] & g[18290];
assign g[34675] = a[14] & g[18291];
assign g[51058] = b[14] & g[18291];
assign g[34676] = a[14] & g[18292];
assign g[51059] = b[14] & g[18292];
assign g[34677] = a[14] & g[18293];
assign g[51060] = b[14] & g[18293];
assign g[34678] = a[14] & g[18294];
assign g[51061] = b[14] & g[18294];
assign g[34679] = a[14] & g[18295];
assign g[51062] = b[14] & g[18295];
assign g[34680] = a[14] & g[18296];
assign g[51063] = b[14] & g[18296];
assign g[34681] = a[14] & g[18297];
assign g[51064] = b[14] & g[18297];
assign g[34682] = a[14] & g[18298];
assign g[51065] = b[14] & g[18298];
assign g[34683] = a[14] & g[18299];
assign g[51066] = b[14] & g[18299];
assign g[34684] = a[14] & g[18300];
assign g[51067] = b[14] & g[18300];
assign g[34685] = a[14] & g[18301];
assign g[51068] = b[14] & g[18301];
assign g[34686] = a[14] & g[18302];
assign g[51069] = b[14] & g[18302];
assign g[34687] = a[14] & g[18303];
assign g[51070] = b[14] & g[18303];
assign g[34688] = a[14] & g[18304];
assign g[51071] = b[14] & g[18304];
assign g[34689] = a[14] & g[18305];
assign g[51072] = b[14] & g[18305];
assign g[34690] = a[14] & g[18306];
assign g[51073] = b[14] & g[18306];
assign g[34691] = a[14] & g[18307];
assign g[51074] = b[14] & g[18307];
assign g[34692] = a[14] & g[18308];
assign g[51075] = b[14] & g[18308];
assign g[34693] = a[14] & g[18309];
assign g[51076] = b[14] & g[18309];
assign g[34694] = a[14] & g[18310];
assign g[51077] = b[14] & g[18310];
assign g[34695] = a[14] & g[18311];
assign g[51078] = b[14] & g[18311];
assign g[34696] = a[14] & g[18312];
assign g[51079] = b[14] & g[18312];
assign g[34697] = a[14] & g[18313];
assign g[51080] = b[14] & g[18313];
assign g[34698] = a[14] & g[18314];
assign g[51081] = b[14] & g[18314];
assign g[34699] = a[14] & g[18315];
assign g[51082] = b[14] & g[18315];
assign g[34700] = a[14] & g[18316];
assign g[51083] = b[14] & g[18316];
assign g[34701] = a[14] & g[18317];
assign g[51084] = b[14] & g[18317];
assign g[34702] = a[14] & g[18318];
assign g[51085] = b[14] & g[18318];
assign g[34703] = a[14] & g[18319];
assign g[51086] = b[14] & g[18319];
assign g[34704] = a[14] & g[18320];
assign g[51087] = b[14] & g[18320];
assign g[34705] = a[14] & g[18321];
assign g[51088] = b[14] & g[18321];
assign g[34706] = a[14] & g[18322];
assign g[51089] = b[14] & g[18322];
assign g[34707] = a[14] & g[18323];
assign g[51090] = b[14] & g[18323];
assign g[34708] = a[14] & g[18324];
assign g[51091] = b[14] & g[18324];
assign g[34709] = a[14] & g[18325];
assign g[51092] = b[14] & g[18325];
assign g[34710] = a[14] & g[18326];
assign g[51093] = b[14] & g[18326];
assign g[34711] = a[14] & g[18327];
assign g[51094] = b[14] & g[18327];
assign g[34712] = a[14] & g[18328];
assign g[51095] = b[14] & g[18328];
assign g[34713] = a[14] & g[18329];
assign g[51096] = b[14] & g[18329];
assign g[34714] = a[14] & g[18330];
assign g[51097] = b[14] & g[18330];
assign g[34715] = a[14] & g[18331];
assign g[51098] = b[14] & g[18331];
assign g[34716] = a[14] & g[18332];
assign g[51099] = b[14] & g[18332];
assign g[34717] = a[14] & g[18333];
assign g[51100] = b[14] & g[18333];
assign g[34718] = a[14] & g[18334];
assign g[51101] = b[14] & g[18334];
assign g[34719] = a[14] & g[18335];
assign g[51102] = b[14] & g[18335];
assign g[34720] = a[14] & g[18336];
assign g[51103] = b[14] & g[18336];
assign g[34721] = a[14] & g[18337];
assign g[51104] = b[14] & g[18337];
assign g[34722] = a[14] & g[18338];
assign g[51105] = b[14] & g[18338];
assign g[34723] = a[14] & g[18339];
assign g[51106] = b[14] & g[18339];
assign g[34724] = a[14] & g[18340];
assign g[51107] = b[14] & g[18340];
assign g[34725] = a[14] & g[18341];
assign g[51108] = b[14] & g[18341];
assign g[34726] = a[14] & g[18342];
assign g[51109] = b[14] & g[18342];
assign g[34727] = a[14] & g[18343];
assign g[51110] = b[14] & g[18343];
assign g[34728] = a[14] & g[18344];
assign g[51111] = b[14] & g[18344];
assign g[34729] = a[14] & g[18345];
assign g[51112] = b[14] & g[18345];
assign g[34730] = a[14] & g[18346];
assign g[51113] = b[14] & g[18346];
assign g[34731] = a[14] & g[18347];
assign g[51114] = b[14] & g[18347];
assign g[34732] = a[14] & g[18348];
assign g[51115] = b[14] & g[18348];
assign g[34733] = a[14] & g[18349];
assign g[51116] = b[14] & g[18349];
assign g[34734] = a[14] & g[18350];
assign g[51117] = b[14] & g[18350];
assign g[34735] = a[14] & g[18351];
assign g[51118] = b[14] & g[18351];
assign g[34736] = a[14] & g[18352];
assign g[51119] = b[14] & g[18352];
assign g[34737] = a[14] & g[18353];
assign g[51120] = b[14] & g[18353];
assign g[34738] = a[14] & g[18354];
assign g[51121] = b[14] & g[18354];
assign g[34739] = a[14] & g[18355];
assign g[51122] = b[14] & g[18355];
assign g[34740] = a[14] & g[18356];
assign g[51123] = b[14] & g[18356];
assign g[34741] = a[14] & g[18357];
assign g[51124] = b[14] & g[18357];
assign g[34742] = a[14] & g[18358];
assign g[51125] = b[14] & g[18358];
assign g[34743] = a[14] & g[18359];
assign g[51126] = b[14] & g[18359];
assign g[34744] = a[14] & g[18360];
assign g[51127] = b[14] & g[18360];
assign g[34745] = a[14] & g[18361];
assign g[51128] = b[14] & g[18361];
assign g[34746] = a[14] & g[18362];
assign g[51129] = b[14] & g[18362];
assign g[34747] = a[14] & g[18363];
assign g[51130] = b[14] & g[18363];
assign g[34748] = a[14] & g[18364];
assign g[51131] = b[14] & g[18364];
assign g[34749] = a[14] & g[18365];
assign g[51132] = b[14] & g[18365];
assign g[34750] = a[14] & g[18366];
assign g[51133] = b[14] & g[18366];
assign g[34751] = a[14] & g[18367];
assign g[51134] = b[14] & g[18367];
assign g[34752] = a[14] & g[18368];
assign g[51135] = b[14] & g[18368];
assign g[34753] = a[14] & g[18369];
assign g[51136] = b[14] & g[18369];
assign g[34754] = a[14] & g[18370];
assign g[51137] = b[14] & g[18370];
assign g[34755] = a[14] & g[18371];
assign g[51138] = b[14] & g[18371];
assign g[34756] = a[14] & g[18372];
assign g[51139] = b[14] & g[18372];
assign g[34757] = a[14] & g[18373];
assign g[51140] = b[14] & g[18373];
assign g[34758] = a[14] & g[18374];
assign g[51141] = b[14] & g[18374];
assign g[34759] = a[14] & g[18375];
assign g[51142] = b[14] & g[18375];
assign g[34760] = a[14] & g[18376];
assign g[51143] = b[14] & g[18376];
assign g[34761] = a[14] & g[18377];
assign g[51144] = b[14] & g[18377];
assign g[34762] = a[14] & g[18378];
assign g[51145] = b[14] & g[18378];
assign g[34763] = a[14] & g[18379];
assign g[51146] = b[14] & g[18379];
assign g[34764] = a[14] & g[18380];
assign g[51147] = b[14] & g[18380];
assign g[34765] = a[14] & g[18381];
assign g[51148] = b[14] & g[18381];
assign g[34766] = a[14] & g[18382];
assign g[51149] = b[14] & g[18382];
assign g[34767] = a[14] & g[18383];
assign g[51150] = b[14] & g[18383];
assign g[34768] = a[14] & g[18384];
assign g[51151] = b[14] & g[18384];
assign g[34769] = a[14] & g[18385];
assign g[51152] = b[14] & g[18385];
assign g[34770] = a[14] & g[18386];
assign g[51153] = b[14] & g[18386];
assign g[34771] = a[14] & g[18387];
assign g[51154] = b[14] & g[18387];
assign g[34772] = a[14] & g[18388];
assign g[51155] = b[14] & g[18388];
assign g[34773] = a[14] & g[18389];
assign g[51156] = b[14] & g[18389];
assign g[34774] = a[14] & g[18390];
assign g[51157] = b[14] & g[18390];
assign g[34775] = a[14] & g[18391];
assign g[51158] = b[14] & g[18391];
assign g[34776] = a[14] & g[18392];
assign g[51159] = b[14] & g[18392];
assign g[34777] = a[14] & g[18393];
assign g[51160] = b[14] & g[18393];
assign g[34778] = a[14] & g[18394];
assign g[51161] = b[14] & g[18394];
assign g[34779] = a[14] & g[18395];
assign g[51162] = b[14] & g[18395];
assign g[34780] = a[14] & g[18396];
assign g[51163] = b[14] & g[18396];
assign g[34781] = a[14] & g[18397];
assign g[51164] = b[14] & g[18397];
assign g[34782] = a[14] & g[18398];
assign g[51165] = b[14] & g[18398];
assign g[34783] = a[14] & g[18399];
assign g[51166] = b[14] & g[18399];
assign g[34784] = a[14] & g[18400];
assign g[51167] = b[14] & g[18400];
assign g[34785] = a[14] & g[18401];
assign g[51168] = b[14] & g[18401];
assign g[34786] = a[14] & g[18402];
assign g[51169] = b[14] & g[18402];
assign g[34787] = a[14] & g[18403];
assign g[51170] = b[14] & g[18403];
assign g[34788] = a[14] & g[18404];
assign g[51171] = b[14] & g[18404];
assign g[34789] = a[14] & g[18405];
assign g[51172] = b[14] & g[18405];
assign g[34790] = a[14] & g[18406];
assign g[51173] = b[14] & g[18406];
assign g[34791] = a[14] & g[18407];
assign g[51174] = b[14] & g[18407];
assign g[34792] = a[14] & g[18408];
assign g[51175] = b[14] & g[18408];
assign g[34793] = a[14] & g[18409];
assign g[51176] = b[14] & g[18409];
assign g[34794] = a[14] & g[18410];
assign g[51177] = b[14] & g[18410];
assign g[34795] = a[14] & g[18411];
assign g[51178] = b[14] & g[18411];
assign g[34796] = a[14] & g[18412];
assign g[51179] = b[14] & g[18412];
assign g[34797] = a[14] & g[18413];
assign g[51180] = b[14] & g[18413];
assign g[34798] = a[14] & g[18414];
assign g[51181] = b[14] & g[18414];
assign g[34799] = a[14] & g[18415];
assign g[51182] = b[14] & g[18415];
assign g[34800] = a[14] & g[18416];
assign g[51183] = b[14] & g[18416];
assign g[34801] = a[14] & g[18417];
assign g[51184] = b[14] & g[18417];
assign g[34802] = a[14] & g[18418];
assign g[51185] = b[14] & g[18418];
assign g[34803] = a[14] & g[18419];
assign g[51186] = b[14] & g[18419];
assign g[34804] = a[14] & g[18420];
assign g[51187] = b[14] & g[18420];
assign g[34805] = a[14] & g[18421];
assign g[51188] = b[14] & g[18421];
assign g[34806] = a[14] & g[18422];
assign g[51189] = b[14] & g[18422];
assign g[34807] = a[14] & g[18423];
assign g[51190] = b[14] & g[18423];
assign g[34808] = a[14] & g[18424];
assign g[51191] = b[14] & g[18424];
assign g[34809] = a[14] & g[18425];
assign g[51192] = b[14] & g[18425];
assign g[34810] = a[14] & g[18426];
assign g[51193] = b[14] & g[18426];
assign g[34811] = a[14] & g[18427];
assign g[51194] = b[14] & g[18427];
assign g[34812] = a[14] & g[18428];
assign g[51195] = b[14] & g[18428];
assign g[34813] = a[14] & g[18429];
assign g[51196] = b[14] & g[18429];
assign g[34814] = a[14] & g[18430];
assign g[51197] = b[14] & g[18430];
assign g[34815] = a[14] & g[18431];
assign g[51198] = b[14] & g[18431];
assign g[34816] = a[14] & g[18432];
assign g[51199] = b[14] & g[18432];
assign g[34817] = a[14] & g[18433];
assign g[51200] = b[14] & g[18433];
assign g[34818] = a[14] & g[18434];
assign g[51201] = b[14] & g[18434];
assign g[34819] = a[14] & g[18435];
assign g[51202] = b[14] & g[18435];
assign g[34820] = a[14] & g[18436];
assign g[51203] = b[14] & g[18436];
assign g[34821] = a[14] & g[18437];
assign g[51204] = b[14] & g[18437];
assign g[34822] = a[14] & g[18438];
assign g[51205] = b[14] & g[18438];
assign g[34823] = a[14] & g[18439];
assign g[51206] = b[14] & g[18439];
assign g[34824] = a[14] & g[18440];
assign g[51207] = b[14] & g[18440];
assign g[34825] = a[14] & g[18441];
assign g[51208] = b[14] & g[18441];
assign g[34826] = a[14] & g[18442];
assign g[51209] = b[14] & g[18442];
assign g[34827] = a[14] & g[18443];
assign g[51210] = b[14] & g[18443];
assign g[34828] = a[14] & g[18444];
assign g[51211] = b[14] & g[18444];
assign g[34829] = a[14] & g[18445];
assign g[51212] = b[14] & g[18445];
assign g[34830] = a[14] & g[18446];
assign g[51213] = b[14] & g[18446];
assign g[34831] = a[14] & g[18447];
assign g[51214] = b[14] & g[18447];
assign g[34832] = a[14] & g[18448];
assign g[51215] = b[14] & g[18448];
assign g[34833] = a[14] & g[18449];
assign g[51216] = b[14] & g[18449];
assign g[34834] = a[14] & g[18450];
assign g[51217] = b[14] & g[18450];
assign g[34835] = a[14] & g[18451];
assign g[51218] = b[14] & g[18451];
assign g[34836] = a[14] & g[18452];
assign g[51219] = b[14] & g[18452];
assign g[34837] = a[14] & g[18453];
assign g[51220] = b[14] & g[18453];
assign g[34838] = a[14] & g[18454];
assign g[51221] = b[14] & g[18454];
assign g[34839] = a[14] & g[18455];
assign g[51222] = b[14] & g[18455];
assign g[34840] = a[14] & g[18456];
assign g[51223] = b[14] & g[18456];
assign g[34841] = a[14] & g[18457];
assign g[51224] = b[14] & g[18457];
assign g[34842] = a[14] & g[18458];
assign g[51225] = b[14] & g[18458];
assign g[34843] = a[14] & g[18459];
assign g[51226] = b[14] & g[18459];
assign g[34844] = a[14] & g[18460];
assign g[51227] = b[14] & g[18460];
assign g[34845] = a[14] & g[18461];
assign g[51228] = b[14] & g[18461];
assign g[34846] = a[14] & g[18462];
assign g[51229] = b[14] & g[18462];
assign g[34847] = a[14] & g[18463];
assign g[51230] = b[14] & g[18463];
assign g[34848] = a[14] & g[18464];
assign g[51231] = b[14] & g[18464];
assign g[34849] = a[14] & g[18465];
assign g[51232] = b[14] & g[18465];
assign g[34850] = a[14] & g[18466];
assign g[51233] = b[14] & g[18466];
assign g[34851] = a[14] & g[18467];
assign g[51234] = b[14] & g[18467];
assign g[34852] = a[14] & g[18468];
assign g[51235] = b[14] & g[18468];
assign g[34853] = a[14] & g[18469];
assign g[51236] = b[14] & g[18469];
assign g[34854] = a[14] & g[18470];
assign g[51237] = b[14] & g[18470];
assign g[34855] = a[14] & g[18471];
assign g[51238] = b[14] & g[18471];
assign g[34856] = a[14] & g[18472];
assign g[51239] = b[14] & g[18472];
assign g[34857] = a[14] & g[18473];
assign g[51240] = b[14] & g[18473];
assign g[34858] = a[14] & g[18474];
assign g[51241] = b[14] & g[18474];
assign g[34859] = a[14] & g[18475];
assign g[51242] = b[14] & g[18475];
assign g[34860] = a[14] & g[18476];
assign g[51243] = b[14] & g[18476];
assign g[34861] = a[14] & g[18477];
assign g[51244] = b[14] & g[18477];
assign g[34862] = a[14] & g[18478];
assign g[51245] = b[14] & g[18478];
assign g[34863] = a[14] & g[18479];
assign g[51246] = b[14] & g[18479];
assign g[34864] = a[14] & g[18480];
assign g[51247] = b[14] & g[18480];
assign g[34865] = a[14] & g[18481];
assign g[51248] = b[14] & g[18481];
assign g[34866] = a[14] & g[18482];
assign g[51249] = b[14] & g[18482];
assign g[34867] = a[14] & g[18483];
assign g[51250] = b[14] & g[18483];
assign g[34868] = a[14] & g[18484];
assign g[51251] = b[14] & g[18484];
assign g[34869] = a[14] & g[18485];
assign g[51252] = b[14] & g[18485];
assign g[34870] = a[14] & g[18486];
assign g[51253] = b[14] & g[18486];
assign g[34871] = a[14] & g[18487];
assign g[51254] = b[14] & g[18487];
assign g[34872] = a[14] & g[18488];
assign g[51255] = b[14] & g[18488];
assign g[34873] = a[14] & g[18489];
assign g[51256] = b[14] & g[18489];
assign g[34874] = a[14] & g[18490];
assign g[51257] = b[14] & g[18490];
assign g[34875] = a[14] & g[18491];
assign g[51258] = b[14] & g[18491];
assign g[34876] = a[14] & g[18492];
assign g[51259] = b[14] & g[18492];
assign g[34877] = a[14] & g[18493];
assign g[51260] = b[14] & g[18493];
assign g[34878] = a[14] & g[18494];
assign g[51261] = b[14] & g[18494];
assign g[34879] = a[14] & g[18495];
assign g[51262] = b[14] & g[18495];
assign g[34880] = a[14] & g[18496];
assign g[51263] = b[14] & g[18496];
assign g[34881] = a[14] & g[18497];
assign g[51264] = b[14] & g[18497];
assign g[34882] = a[14] & g[18498];
assign g[51265] = b[14] & g[18498];
assign g[34883] = a[14] & g[18499];
assign g[51266] = b[14] & g[18499];
assign g[34884] = a[14] & g[18500];
assign g[51267] = b[14] & g[18500];
assign g[34885] = a[14] & g[18501];
assign g[51268] = b[14] & g[18501];
assign g[34886] = a[14] & g[18502];
assign g[51269] = b[14] & g[18502];
assign g[34887] = a[14] & g[18503];
assign g[51270] = b[14] & g[18503];
assign g[34888] = a[14] & g[18504];
assign g[51271] = b[14] & g[18504];
assign g[34889] = a[14] & g[18505];
assign g[51272] = b[14] & g[18505];
assign g[34890] = a[14] & g[18506];
assign g[51273] = b[14] & g[18506];
assign g[34891] = a[14] & g[18507];
assign g[51274] = b[14] & g[18507];
assign g[34892] = a[14] & g[18508];
assign g[51275] = b[14] & g[18508];
assign g[34893] = a[14] & g[18509];
assign g[51276] = b[14] & g[18509];
assign g[34894] = a[14] & g[18510];
assign g[51277] = b[14] & g[18510];
assign g[34895] = a[14] & g[18511];
assign g[51278] = b[14] & g[18511];
assign g[34896] = a[14] & g[18512];
assign g[51279] = b[14] & g[18512];
assign g[34897] = a[14] & g[18513];
assign g[51280] = b[14] & g[18513];
assign g[34898] = a[14] & g[18514];
assign g[51281] = b[14] & g[18514];
assign g[34899] = a[14] & g[18515];
assign g[51282] = b[14] & g[18515];
assign g[34900] = a[14] & g[18516];
assign g[51283] = b[14] & g[18516];
assign g[34901] = a[14] & g[18517];
assign g[51284] = b[14] & g[18517];
assign g[34902] = a[14] & g[18518];
assign g[51285] = b[14] & g[18518];
assign g[34903] = a[14] & g[18519];
assign g[51286] = b[14] & g[18519];
assign g[34904] = a[14] & g[18520];
assign g[51287] = b[14] & g[18520];
assign g[34905] = a[14] & g[18521];
assign g[51288] = b[14] & g[18521];
assign g[34906] = a[14] & g[18522];
assign g[51289] = b[14] & g[18522];
assign g[34907] = a[14] & g[18523];
assign g[51290] = b[14] & g[18523];
assign g[34908] = a[14] & g[18524];
assign g[51291] = b[14] & g[18524];
assign g[34909] = a[14] & g[18525];
assign g[51292] = b[14] & g[18525];
assign g[34910] = a[14] & g[18526];
assign g[51293] = b[14] & g[18526];
assign g[34911] = a[14] & g[18527];
assign g[51294] = b[14] & g[18527];
assign g[34912] = a[14] & g[18528];
assign g[51295] = b[14] & g[18528];
assign g[34913] = a[14] & g[18529];
assign g[51296] = b[14] & g[18529];
assign g[34914] = a[14] & g[18530];
assign g[51297] = b[14] & g[18530];
assign g[34915] = a[14] & g[18531];
assign g[51298] = b[14] & g[18531];
assign g[34916] = a[14] & g[18532];
assign g[51299] = b[14] & g[18532];
assign g[34917] = a[14] & g[18533];
assign g[51300] = b[14] & g[18533];
assign g[34918] = a[14] & g[18534];
assign g[51301] = b[14] & g[18534];
assign g[34919] = a[14] & g[18535];
assign g[51302] = b[14] & g[18535];
assign g[34920] = a[14] & g[18536];
assign g[51303] = b[14] & g[18536];
assign g[34921] = a[14] & g[18537];
assign g[51304] = b[14] & g[18537];
assign g[34922] = a[14] & g[18538];
assign g[51305] = b[14] & g[18538];
assign g[34923] = a[14] & g[18539];
assign g[51306] = b[14] & g[18539];
assign g[34924] = a[14] & g[18540];
assign g[51307] = b[14] & g[18540];
assign g[34925] = a[14] & g[18541];
assign g[51308] = b[14] & g[18541];
assign g[34926] = a[14] & g[18542];
assign g[51309] = b[14] & g[18542];
assign g[34927] = a[14] & g[18543];
assign g[51310] = b[14] & g[18543];
assign g[34928] = a[14] & g[18544];
assign g[51311] = b[14] & g[18544];
assign g[34929] = a[14] & g[18545];
assign g[51312] = b[14] & g[18545];
assign g[34930] = a[14] & g[18546];
assign g[51313] = b[14] & g[18546];
assign g[34931] = a[14] & g[18547];
assign g[51314] = b[14] & g[18547];
assign g[34932] = a[14] & g[18548];
assign g[51315] = b[14] & g[18548];
assign g[34933] = a[14] & g[18549];
assign g[51316] = b[14] & g[18549];
assign g[34934] = a[14] & g[18550];
assign g[51317] = b[14] & g[18550];
assign g[34935] = a[14] & g[18551];
assign g[51318] = b[14] & g[18551];
assign g[34936] = a[14] & g[18552];
assign g[51319] = b[14] & g[18552];
assign g[34937] = a[14] & g[18553];
assign g[51320] = b[14] & g[18553];
assign g[34938] = a[14] & g[18554];
assign g[51321] = b[14] & g[18554];
assign g[34939] = a[14] & g[18555];
assign g[51322] = b[14] & g[18555];
assign g[34940] = a[14] & g[18556];
assign g[51323] = b[14] & g[18556];
assign g[34941] = a[14] & g[18557];
assign g[51324] = b[14] & g[18557];
assign g[34942] = a[14] & g[18558];
assign g[51325] = b[14] & g[18558];
assign g[34943] = a[14] & g[18559];
assign g[51326] = b[14] & g[18559];
assign g[34944] = a[14] & g[18560];
assign g[51327] = b[14] & g[18560];
assign g[34945] = a[14] & g[18561];
assign g[51328] = b[14] & g[18561];
assign g[34946] = a[14] & g[18562];
assign g[51329] = b[14] & g[18562];
assign g[34947] = a[14] & g[18563];
assign g[51330] = b[14] & g[18563];
assign g[34948] = a[14] & g[18564];
assign g[51331] = b[14] & g[18564];
assign g[34949] = a[14] & g[18565];
assign g[51332] = b[14] & g[18565];
assign g[34950] = a[14] & g[18566];
assign g[51333] = b[14] & g[18566];
assign g[34951] = a[14] & g[18567];
assign g[51334] = b[14] & g[18567];
assign g[34952] = a[14] & g[18568];
assign g[51335] = b[14] & g[18568];
assign g[34953] = a[14] & g[18569];
assign g[51336] = b[14] & g[18569];
assign g[34954] = a[14] & g[18570];
assign g[51337] = b[14] & g[18570];
assign g[34955] = a[14] & g[18571];
assign g[51338] = b[14] & g[18571];
assign g[34956] = a[14] & g[18572];
assign g[51339] = b[14] & g[18572];
assign g[34957] = a[14] & g[18573];
assign g[51340] = b[14] & g[18573];
assign g[34958] = a[14] & g[18574];
assign g[51341] = b[14] & g[18574];
assign g[34959] = a[14] & g[18575];
assign g[51342] = b[14] & g[18575];
assign g[34960] = a[14] & g[18576];
assign g[51343] = b[14] & g[18576];
assign g[34961] = a[14] & g[18577];
assign g[51344] = b[14] & g[18577];
assign g[34962] = a[14] & g[18578];
assign g[51345] = b[14] & g[18578];
assign g[34963] = a[14] & g[18579];
assign g[51346] = b[14] & g[18579];
assign g[34964] = a[14] & g[18580];
assign g[51347] = b[14] & g[18580];
assign g[34965] = a[14] & g[18581];
assign g[51348] = b[14] & g[18581];
assign g[34966] = a[14] & g[18582];
assign g[51349] = b[14] & g[18582];
assign g[34967] = a[14] & g[18583];
assign g[51350] = b[14] & g[18583];
assign g[34968] = a[14] & g[18584];
assign g[51351] = b[14] & g[18584];
assign g[34969] = a[14] & g[18585];
assign g[51352] = b[14] & g[18585];
assign g[34970] = a[14] & g[18586];
assign g[51353] = b[14] & g[18586];
assign g[34971] = a[14] & g[18587];
assign g[51354] = b[14] & g[18587];
assign g[34972] = a[14] & g[18588];
assign g[51355] = b[14] & g[18588];
assign g[34973] = a[14] & g[18589];
assign g[51356] = b[14] & g[18589];
assign g[34974] = a[14] & g[18590];
assign g[51357] = b[14] & g[18590];
assign g[34975] = a[14] & g[18591];
assign g[51358] = b[14] & g[18591];
assign g[34976] = a[14] & g[18592];
assign g[51359] = b[14] & g[18592];
assign g[34977] = a[14] & g[18593];
assign g[51360] = b[14] & g[18593];
assign g[34978] = a[14] & g[18594];
assign g[51361] = b[14] & g[18594];
assign g[34979] = a[14] & g[18595];
assign g[51362] = b[14] & g[18595];
assign g[34980] = a[14] & g[18596];
assign g[51363] = b[14] & g[18596];
assign g[34981] = a[14] & g[18597];
assign g[51364] = b[14] & g[18597];
assign g[34982] = a[14] & g[18598];
assign g[51365] = b[14] & g[18598];
assign g[34983] = a[14] & g[18599];
assign g[51366] = b[14] & g[18599];
assign g[34984] = a[14] & g[18600];
assign g[51367] = b[14] & g[18600];
assign g[34985] = a[14] & g[18601];
assign g[51368] = b[14] & g[18601];
assign g[34986] = a[14] & g[18602];
assign g[51369] = b[14] & g[18602];
assign g[34987] = a[14] & g[18603];
assign g[51370] = b[14] & g[18603];
assign g[34988] = a[14] & g[18604];
assign g[51371] = b[14] & g[18604];
assign g[34989] = a[14] & g[18605];
assign g[51372] = b[14] & g[18605];
assign g[34990] = a[14] & g[18606];
assign g[51373] = b[14] & g[18606];
assign g[34991] = a[14] & g[18607];
assign g[51374] = b[14] & g[18607];
assign g[34992] = a[14] & g[18608];
assign g[51375] = b[14] & g[18608];
assign g[34993] = a[14] & g[18609];
assign g[51376] = b[14] & g[18609];
assign g[34994] = a[14] & g[18610];
assign g[51377] = b[14] & g[18610];
assign g[34995] = a[14] & g[18611];
assign g[51378] = b[14] & g[18611];
assign g[34996] = a[14] & g[18612];
assign g[51379] = b[14] & g[18612];
assign g[34997] = a[14] & g[18613];
assign g[51380] = b[14] & g[18613];
assign g[34998] = a[14] & g[18614];
assign g[51381] = b[14] & g[18614];
assign g[34999] = a[14] & g[18615];
assign g[51382] = b[14] & g[18615];
assign g[35000] = a[14] & g[18616];
assign g[51383] = b[14] & g[18616];
assign g[35001] = a[14] & g[18617];
assign g[51384] = b[14] & g[18617];
assign g[35002] = a[14] & g[18618];
assign g[51385] = b[14] & g[18618];
assign g[35003] = a[14] & g[18619];
assign g[51386] = b[14] & g[18619];
assign g[35004] = a[14] & g[18620];
assign g[51387] = b[14] & g[18620];
assign g[35005] = a[14] & g[18621];
assign g[51388] = b[14] & g[18621];
assign g[35006] = a[14] & g[18622];
assign g[51389] = b[14] & g[18622];
assign g[35007] = a[14] & g[18623];
assign g[51390] = b[14] & g[18623];
assign g[35008] = a[14] & g[18624];
assign g[51391] = b[14] & g[18624];
assign g[35009] = a[14] & g[18625];
assign g[51392] = b[14] & g[18625];
assign g[35010] = a[14] & g[18626];
assign g[51393] = b[14] & g[18626];
assign g[35011] = a[14] & g[18627];
assign g[51394] = b[14] & g[18627];
assign g[35012] = a[14] & g[18628];
assign g[51395] = b[14] & g[18628];
assign g[35013] = a[14] & g[18629];
assign g[51396] = b[14] & g[18629];
assign g[35014] = a[14] & g[18630];
assign g[51397] = b[14] & g[18630];
assign g[35015] = a[14] & g[18631];
assign g[51398] = b[14] & g[18631];
assign g[35016] = a[14] & g[18632];
assign g[51399] = b[14] & g[18632];
assign g[35017] = a[14] & g[18633];
assign g[51400] = b[14] & g[18633];
assign g[35018] = a[14] & g[18634];
assign g[51401] = b[14] & g[18634];
assign g[35019] = a[14] & g[18635];
assign g[51402] = b[14] & g[18635];
assign g[35020] = a[14] & g[18636];
assign g[51403] = b[14] & g[18636];
assign g[35021] = a[14] & g[18637];
assign g[51404] = b[14] & g[18637];
assign g[35022] = a[14] & g[18638];
assign g[51405] = b[14] & g[18638];
assign g[35023] = a[14] & g[18639];
assign g[51406] = b[14] & g[18639];
assign g[35024] = a[14] & g[18640];
assign g[51407] = b[14] & g[18640];
assign g[35025] = a[14] & g[18641];
assign g[51408] = b[14] & g[18641];
assign g[35026] = a[14] & g[18642];
assign g[51409] = b[14] & g[18642];
assign g[35027] = a[14] & g[18643];
assign g[51410] = b[14] & g[18643];
assign g[35028] = a[14] & g[18644];
assign g[51411] = b[14] & g[18644];
assign g[35029] = a[14] & g[18645];
assign g[51412] = b[14] & g[18645];
assign g[35030] = a[14] & g[18646];
assign g[51413] = b[14] & g[18646];
assign g[35031] = a[14] & g[18647];
assign g[51414] = b[14] & g[18647];
assign g[35032] = a[14] & g[18648];
assign g[51415] = b[14] & g[18648];
assign g[35033] = a[14] & g[18649];
assign g[51416] = b[14] & g[18649];
assign g[35034] = a[14] & g[18650];
assign g[51417] = b[14] & g[18650];
assign g[35035] = a[14] & g[18651];
assign g[51418] = b[14] & g[18651];
assign g[35036] = a[14] & g[18652];
assign g[51419] = b[14] & g[18652];
assign g[35037] = a[14] & g[18653];
assign g[51420] = b[14] & g[18653];
assign g[35038] = a[14] & g[18654];
assign g[51421] = b[14] & g[18654];
assign g[35039] = a[14] & g[18655];
assign g[51422] = b[14] & g[18655];
assign g[35040] = a[14] & g[18656];
assign g[51423] = b[14] & g[18656];
assign g[35041] = a[14] & g[18657];
assign g[51424] = b[14] & g[18657];
assign g[35042] = a[14] & g[18658];
assign g[51425] = b[14] & g[18658];
assign g[35043] = a[14] & g[18659];
assign g[51426] = b[14] & g[18659];
assign g[35044] = a[14] & g[18660];
assign g[51427] = b[14] & g[18660];
assign g[35045] = a[14] & g[18661];
assign g[51428] = b[14] & g[18661];
assign g[35046] = a[14] & g[18662];
assign g[51429] = b[14] & g[18662];
assign g[35047] = a[14] & g[18663];
assign g[51430] = b[14] & g[18663];
assign g[35048] = a[14] & g[18664];
assign g[51431] = b[14] & g[18664];
assign g[35049] = a[14] & g[18665];
assign g[51432] = b[14] & g[18665];
assign g[35050] = a[14] & g[18666];
assign g[51433] = b[14] & g[18666];
assign g[35051] = a[14] & g[18667];
assign g[51434] = b[14] & g[18667];
assign g[35052] = a[14] & g[18668];
assign g[51435] = b[14] & g[18668];
assign g[35053] = a[14] & g[18669];
assign g[51436] = b[14] & g[18669];
assign g[35054] = a[14] & g[18670];
assign g[51437] = b[14] & g[18670];
assign g[35055] = a[14] & g[18671];
assign g[51438] = b[14] & g[18671];
assign g[35056] = a[14] & g[18672];
assign g[51439] = b[14] & g[18672];
assign g[35057] = a[14] & g[18673];
assign g[51440] = b[14] & g[18673];
assign g[35058] = a[14] & g[18674];
assign g[51441] = b[14] & g[18674];
assign g[35059] = a[14] & g[18675];
assign g[51442] = b[14] & g[18675];
assign g[35060] = a[14] & g[18676];
assign g[51443] = b[14] & g[18676];
assign g[35061] = a[14] & g[18677];
assign g[51444] = b[14] & g[18677];
assign g[35062] = a[14] & g[18678];
assign g[51445] = b[14] & g[18678];
assign g[35063] = a[14] & g[18679];
assign g[51446] = b[14] & g[18679];
assign g[35064] = a[14] & g[18680];
assign g[51447] = b[14] & g[18680];
assign g[35065] = a[14] & g[18681];
assign g[51448] = b[14] & g[18681];
assign g[35066] = a[14] & g[18682];
assign g[51449] = b[14] & g[18682];
assign g[35067] = a[14] & g[18683];
assign g[51450] = b[14] & g[18683];
assign g[35068] = a[14] & g[18684];
assign g[51451] = b[14] & g[18684];
assign g[35069] = a[14] & g[18685];
assign g[51452] = b[14] & g[18685];
assign g[35070] = a[14] & g[18686];
assign g[51453] = b[14] & g[18686];
assign g[35071] = a[14] & g[18687];
assign g[51454] = b[14] & g[18687];
assign g[35072] = a[14] & g[18688];
assign g[51455] = b[14] & g[18688];
assign g[35073] = a[14] & g[18689];
assign g[51456] = b[14] & g[18689];
assign g[35074] = a[14] & g[18690];
assign g[51457] = b[14] & g[18690];
assign g[35075] = a[14] & g[18691];
assign g[51458] = b[14] & g[18691];
assign g[35076] = a[14] & g[18692];
assign g[51459] = b[14] & g[18692];
assign g[35077] = a[14] & g[18693];
assign g[51460] = b[14] & g[18693];
assign g[35078] = a[14] & g[18694];
assign g[51461] = b[14] & g[18694];
assign g[35079] = a[14] & g[18695];
assign g[51462] = b[14] & g[18695];
assign g[35080] = a[14] & g[18696];
assign g[51463] = b[14] & g[18696];
assign g[35081] = a[14] & g[18697];
assign g[51464] = b[14] & g[18697];
assign g[35082] = a[14] & g[18698];
assign g[51465] = b[14] & g[18698];
assign g[35083] = a[14] & g[18699];
assign g[51466] = b[14] & g[18699];
assign g[35084] = a[14] & g[18700];
assign g[51467] = b[14] & g[18700];
assign g[35085] = a[14] & g[18701];
assign g[51468] = b[14] & g[18701];
assign g[35086] = a[14] & g[18702];
assign g[51469] = b[14] & g[18702];
assign g[35087] = a[14] & g[18703];
assign g[51470] = b[14] & g[18703];
assign g[35088] = a[14] & g[18704];
assign g[51471] = b[14] & g[18704];
assign g[35089] = a[14] & g[18705];
assign g[51472] = b[14] & g[18705];
assign g[35090] = a[14] & g[18706];
assign g[51473] = b[14] & g[18706];
assign g[35091] = a[14] & g[18707];
assign g[51474] = b[14] & g[18707];
assign g[35092] = a[14] & g[18708];
assign g[51475] = b[14] & g[18708];
assign g[35093] = a[14] & g[18709];
assign g[51476] = b[14] & g[18709];
assign g[35094] = a[14] & g[18710];
assign g[51477] = b[14] & g[18710];
assign g[35095] = a[14] & g[18711];
assign g[51478] = b[14] & g[18711];
assign g[35096] = a[14] & g[18712];
assign g[51479] = b[14] & g[18712];
assign g[35097] = a[14] & g[18713];
assign g[51480] = b[14] & g[18713];
assign g[35098] = a[14] & g[18714];
assign g[51481] = b[14] & g[18714];
assign g[35099] = a[14] & g[18715];
assign g[51482] = b[14] & g[18715];
assign g[35100] = a[14] & g[18716];
assign g[51483] = b[14] & g[18716];
assign g[35101] = a[14] & g[18717];
assign g[51484] = b[14] & g[18717];
assign g[35102] = a[14] & g[18718];
assign g[51485] = b[14] & g[18718];
assign g[35103] = a[14] & g[18719];
assign g[51486] = b[14] & g[18719];
assign g[35104] = a[14] & g[18720];
assign g[51487] = b[14] & g[18720];
assign g[35105] = a[14] & g[18721];
assign g[51488] = b[14] & g[18721];
assign g[35106] = a[14] & g[18722];
assign g[51489] = b[14] & g[18722];
assign g[35107] = a[14] & g[18723];
assign g[51490] = b[14] & g[18723];
assign g[35108] = a[14] & g[18724];
assign g[51491] = b[14] & g[18724];
assign g[35109] = a[14] & g[18725];
assign g[51492] = b[14] & g[18725];
assign g[35110] = a[14] & g[18726];
assign g[51493] = b[14] & g[18726];
assign g[35111] = a[14] & g[18727];
assign g[51494] = b[14] & g[18727];
assign g[35112] = a[14] & g[18728];
assign g[51495] = b[14] & g[18728];
assign g[35113] = a[14] & g[18729];
assign g[51496] = b[14] & g[18729];
assign g[35114] = a[14] & g[18730];
assign g[51497] = b[14] & g[18730];
assign g[35115] = a[14] & g[18731];
assign g[51498] = b[14] & g[18731];
assign g[35116] = a[14] & g[18732];
assign g[51499] = b[14] & g[18732];
assign g[35117] = a[14] & g[18733];
assign g[51500] = b[14] & g[18733];
assign g[35118] = a[14] & g[18734];
assign g[51501] = b[14] & g[18734];
assign g[35119] = a[14] & g[18735];
assign g[51502] = b[14] & g[18735];
assign g[35120] = a[14] & g[18736];
assign g[51503] = b[14] & g[18736];
assign g[35121] = a[14] & g[18737];
assign g[51504] = b[14] & g[18737];
assign g[35122] = a[14] & g[18738];
assign g[51505] = b[14] & g[18738];
assign g[35123] = a[14] & g[18739];
assign g[51506] = b[14] & g[18739];
assign g[35124] = a[14] & g[18740];
assign g[51507] = b[14] & g[18740];
assign g[35125] = a[14] & g[18741];
assign g[51508] = b[14] & g[18741];
assign g[35126] = a[14] & g[18742];
assign g[51509] = b[14] & g[18742];
assign g[35127] = a[14] & g[18743];
assign g[51510] = b[14] & g[18743];
assign g[35128] = a[14] & g[18744];
assign g[51511] = b[14] & g[18744];
assign g[35129] = a[14] & g[18745];
assign g[51512] = b[14] & g[18745];
assign g[35130] = a[14] & g[18746];
assign g[51513] = b[14] & g[18746];
assign g[35131] = a[14] & g[18747];
assign g[51514] = b[14] & g[18747];
assign g[35132] = a[14] & g[18748];
assign g[51515] = b[14] & g[18748];
assign g[35133] = a[14] & g[18749];
assign g[51516] = b[14] & g[18749];
assign g[35134] = a[14] & g[18750];
assign g[51517] = b[14] & g[18750];
assign g[35135] = a[14] & g[18751];
assign g[51518] = b[14] & g[18751];
assign g[35136] = a[14] & g[18752];
assign g[51519] = b[14] & g[18752];
assign g[35137] = a[14] & g[18753];
assign g[51520] = b[14] & g[18753];
assign g[35138] = a[14] & g[18754];
assign g[51521] = b[14] & g[18754];
assign g[35139] = a[14] & g[18755];
assign g[51522] = b[14] & g[18755];
assign g[35140] = a[14] & g[18756];
assign g[51523] = b[14] & g[18756];
assign g[35141] = a[14] & g[18757];
assign g[51524] = b[14] & g[18757];
assign g[35142] = a[14] & g[18758];
assign g[51525] = b[14] & g[18758];
assign g[35143] = a[14] & g[18759];
assign g[51526] = b[14] & g[18759];
assign g[35144] = a[14] & g[18760];
assign g[51527] = b[14] & g[18760];
assign g[35145] = a[14] & g[18761];
assign g[51528] = b[14] & g[18761];
assign g[35146] = a[14] & g[18762];
assign g[51529] = b[14] & g[18762];
assign g[35147] = a[14] & g[18763];
assign g[51530] = b[14] & g[18763];
assign g[35148] = a[14] & g[18764];
assign g[51531] = b[14] & g[18764];
assign g[35149] = a[14] & g[18765];
assign g[51532] = b[14] & g[18765];
assign g[35150] = a[14] & g[18766];
assign g[51533] = b[14] & g[18766];
assign g[35151] = a[14] & g[18767];
assign g[51534] = b[14] & g[18767];
assign g[35152] = a[14] & g[18768];
assign g[51535] = b[14] & g[18768];
assign g[35153] = a[14] & g[18769];
assign g[51536] = b[14] & g[18769];
assign g[35154] = a[14] & g[18770];
assign g[51537] = b[14] & g[18770];
assign g[35155] = a[14] & g[18771];
assign g[51538] = b[14] & g[18771];
assign g[35156] = a[14] & g[18772];
assign g[51539] = b[14] & g[18772];
assign g[35157] = a[14] & g[18773];
assign g[51540] = b[14] & g[18773];
assign g[35158] = a[14] & g[18774];
assign g[51541] = b[14] & g[18774];
assign g[35159] = a[14] & g[18775];
assign g[51542] = b[14] & g[18775];
assign g[35160] = a[14] & g[18776];
assign g[51543] = b[14] & g[18776];
assign g[35161] = a[14] & g[18777];
assign g[51544] = b[14] & g[18777];
assign g[35162] = a[14] & g[18778];
assign g[51545] = b[14] & g[18778];
assign g[35163] = a[14] & g[18779];
assign g[51546] = b[14] & g[18779];
assign g[35164] = a[14] & g[18780];
assign g[51547] = b[14] & g[18780];
assign g[35165] = a[14] & g[18781];
assign g[51548] = b[14] & g[18781];
assign g[35166] = a[14] & g[18782];
assign g[51549] = b[14] & g[18782];
assign g[35167] = a[14] & g[18783];
assign g[51550] = b[14] & g[18783];
assign g[35168] = a[14] & g[18784];
assign g[51551] = b[14] & g[18784];
assign g[35169] = a[14] & g[18785];
assign g[51552] = b[14] & g[18785];
assign g[35170] = a[14] & g[18786];
assign g[51553] = b[14] & g[18786];
assign g[35171] = a[14] & g[18787];
assign g[51554] = b[14] & g[18787];
assign g[35172] = a[14] & g[18788];
assign g[51555] = b[14] & g[18788];
assign g[35173] = a[14] & g[18789];
assign g[51556] = b[14] & g[18789];
assign g[35174] = a[14] & g[18790];
assign g[51557] = b[14] & g[18790];
assign g[35175] = a[14] & g[18791];
assign g[51558] = b[14] & g[18791];
assign g[35176] = a[14] & g[18792];
assign g[51559] = b[14] & g[18792];
assign g[35177] = a[14] & g[18793];
assign g[51560] = b[14] & g[18793];
assign g[35178] = a[14] & g[18794];
assign g[51561] = b[14] & g[18794];
assign g[35179] = a[14] & g[18795];
assign g[51562] = b[14] & g[18795];
assign g[35180] = a[14] & g[18796];
assign g[51563] = b[14] & g[18796];
assign g[35181] = a[14] & g[18797];
assign g[51564] = b[14] & g[18797];
assign g[35182] = a[14] & g[18798];
assign g[51565] = b[14] & g[18798];
assign g[35183] = a[14] & g[18799];
assign g[51566] = b[14] & g[18799];
assign g[35184] = a[14] & g[18800];
assign g[51567] = b[14] & g[18800];
assign g[35185] = a[14] & g[18801];
assign g[51568] = b[14] & g[18801];
assign g[35186] = a[14] & g[18802];
assign g[51569] = b[14] & g[18802];
assign g[35187] = a[14] & g[18803];
assign g[51570] = b[14] & g[18803];
assign g[35188] = a[14] & g[18804];
assign g[51571] = b[14] & g[18804];
assign g[35189] = a[14] & g[18805];
assign g[51572] = b[14] & g[18805];
assign g[35190] = a[14] & g[18806];
assign g[51573] = b[14] & g[18806];
assign g[35191] = a[14] & g[18807];
assign g[51574] = b[14] & g[18807];
assign g[35192] = a[14] & g[18808];
assign g[51575] = b[14] & g[18808];
assign g[35193] = a[14] & g[18809];
assign g[51576] = b[14] & g[18809];
assign g[35194] = a[14] & g[18810];
assign g[51577] = b[14] & g[18810];
assign g[35195] = a[14] & g[18811];
assign g[51578] = b[14] & g[18811];
assign g[35196] = a[14] & g[18812];
assign g[51579] = b[14] & g[18812];
assign g[35197] = a[14] & g[18813];
assign g[51580] = b[14] & g[18813];
assign g[35198] = a[14] & g[18814];
assign g[51581] = b[14] & g[18814];
assign g[35199] = a[14] & g[18815];
assign g[51582] = b[14] & g[18815];
assign g[35200] = a[14] & g[18816];
assign g[51583] = b[14] & g[18816];
assign g[35201] = a[14] & g[18817];
assign g[51584] = b[14] & g[18817];
assign g[35202] = a[14] & g[18818];
assign g[51585] = b[14] & g[18818];
assign g[35203] = a[14] & g[18819];
assign g[51586] = b[14] & g[18819];
assign g[35204] = a[14] & g[18820];
assign g[51587] = b[14] & g[18820];
assign g[35205] = a[14] & g[18821];
assign g[51588] = b[14] & g[18821];
assign g[35206] = a[14] & g[18822];
assign g[51589] = b[14] & g[18822];
assign g[35207] = a[14] & g[18823];
assign g[51590] = b[14] & g[18823];
assign g[35208] = a[14] & g[18824];
assign g[51591] = b[14] & g[18824];
assign g[35209] = a[14] & g[18825];
assign g[51592] = b[14] & g[18825];
assign g[35210] = a[14] & g[18826];
assign g[51593] = b[14] & g[18826];
assign g[35211] = a[14] & g[18827];
assign g[51594] = b[14] & g[18827];
assign g[35212] = a[14] & g[18828];
assign g[51595] = b[14] & g[18828];
assign g[35213] = a[14] & g[18829];
assign g[51596] = b[14] & g[18829];
assign g[35214] = a[14] & g[18830];
assign g[51597] = b[14] & g[18830];
assign g[35215] = a[14] & g[18831];
assign g[51598] = b[14] & g[18831];
assign g[35216] = a[14] & g[18832];
assign g[51599] = b[14] & g[18832];
assign g[35217] = a[14] & g[18833];
assign g[51600] = b[14] & g[18833];
assign g[35218] = a[14] & g[18834];
assign g[51601] = b[14] & g[18834];
assign g[35219] = a[14] & g[18835];
assign g[51602] = b[14] & g[18835];
assign g[35220] = a[14] & g[18836];
assign g[51603] = b[14] & g[18836];
assign g[35221] = a[14] & g[18837];
assign g[51604] = b[14] & g[18837];
assign g[35222] = a[14] & g[18838];
assign g[51605] = b[14] & g[18838];
assign g[35223] = a[14] & g[18839];
assign g[51606] = b[14] & g[18839];
assign g[35224] = a[14] & g[18840];
assign g[51607] = b[14] & g[18840];
assign g[35225] = a[14] & g[18841];
assign g[51608] = b[14] & g[18841];
assign g[35226] = a[14] & g[18842];
assign g[51609] = b[14] & g[18842];
assign g[35227] = a[14] & g[18843];
assign g[51610] = b[14] & g[18843];
assign g[35228] = a[14] & g[18844];
assign g[51611] = b[14] & g[18844];
assign g[35229] = a[14] & g[18845];
assign g[51612] = b[14] & g[18845];
assign g[35230] = a[14] & g[18846];
assign g[51613] = b[14] & g[18846];
assign g[35231] = a[14] & g[18847];
assign g[51614] = b[14] & g[18847];
assign g[35232] = a[14] & g[18848];
assign g[51615] = b[14] & g[18848];
assign g[35233] = a[14] & g[18849];
assign g[51616] = b[14] & g[18849];
assign g[35234] = a[14] & g[18850];
assign g[51617] = b[14] & g[18850];
assign g[35235] = a[14] & g[18851];
assign g[51618] = b[14] & g[18851];
assign g[35236] = a[14] & g[18852];
assign g[51619] = b[14] & g[18852];
assign g[35237] = a[14] & g[18853];
assign g[51620] = b[14] & g[18853];
assign g[35238] = a[14] & g[18854];
assign g[51621] = b[14] & g[18854];
assign g[35239] = a[14] & g[18855];
assign g[51622] = b[14] & g[18855];
assign g[35240] = a[14] & g[18856];
assign g[51623] = b[14] & g[18856];
assign g[35241] = a[14] & g[18857];
assign g[51624] = b[14] & g[18857];
assign g[35242] = a[14] & g[18858];
assign g[51625] = b[14] & g[18858];
assign g[35243] = a[14] & g[18859];
assign g[51626] = b[14] & g[18859];
assign g[35244] = a[14] & g[18860];
assign g[51627] = b[14] & g[18860];
assign g[35245] = a[14] & g[18861];
assign g[51628] = b[14] & g[18861];
assign g[35246] = a[14] & g[18862];
assign g[51629] = b[14] & g[18862];
assign g[35247] = a[14] & g[18863];
assign g[51630] = b[14] & g[18863];
assign g[35248] = a[14] & g[18864];
assign g[51631] = b[14] & g[18864];
assign g[35249] = a[14] & g[18865];
assign g[51632] = b[14] & g[18865];
assign g[35250] = a[14] & g[18866];
assign g[51633] = b[14] & g[18866];
assign g[35251] = a[14] & g[18867];
assign g[51634] = b[14] & g[18867];
assign g[35252] = a[14] & g[18868];
assign g[51635] = b[14] & g[18868];
assign g[35253] = a[14] & g[18869];
assign g[51636] = b[14] & g[18869];
assign g[35254] = a[14] & g[18870];
assign g[51637] = b[14] & g[18870];
assign g[35255] = a[14] & g[18871];
assign g[51638] = b[14] & g[18871];
assign g[35256] = a[14] & g[18872];
assign g[51639] = b[14] & g[18872];
assign g[35257] = a[14] & g[18873];
assign g[51640] = b[14] & g[18873];
assign g[35258] = a[14] & g[18874];
assign g[51641] = b[14] & g[18874];
assign g[35259] = a[14] & g[18875];
assign g[51642] = b[14] & g[18875];
assign g[35260] = a[14] & g[18876];
assign g[51643] = b[14] & g[18876];
assign g[35261] = a[14] & g[18877];
assign g[51644] = b[14] & g[18877];
assign g[35262] = a[14] & g[18878];
assign g[51645] = b[14] & g[18878];
assign g[35263] = a[14] & g[18879];
assign g[51646] = b[14] & g[18879];
assign g[35264] = a[14] & g[18880];
assign g[51647] = b[14] & g[18880];
assign g[35265] = a[14] & g[18881];
assign g[51648] = b[14] & g[18881];
assign g[35266] = a[14] & g[18882];
assign g[51649] = b[14] & g[18882];
assign g[35267] = a[14] & g[18883];
assign g[51650] = b[14] & g[18883];
assign g[35268] = a[14] & g[18884];
assign g[51651] = b[14] & g[18884];
assign g[35269] = a[14] & g[18885];
assign g[51652] = b[14] & g[18885];
assign g[35270] = a[14] & g[18886];
assign g[51653] = b[14] & g[18886];
assign g[35271] = a[14] & g[18887];
assign g[51654] = b[14] & g[18887];
assign g[35272] = a[14] & g[18888];
assign g[51655] = b[14] & g[18888];
assign g[35273] = a[14] & g[18889];
assign g[51656] = b[14] & g[18889];
assign g[35274] = a[14] & g[18890];
assign g[51657] = b[14] & g[18890];
assign g[35275] = a[14] & g[18891];
assign g[51658] = b[14] & g[18891];
assign g[35276] = a[14] & g[18892];
assign g[51659] = b[14] & g[18892];
assign g[35277] = a[14] & g[18893];
assign g[51660] = b[14] & g[18893];
assign g[35278] = a[14] & g[18894];
assign g[51661] = b[14] & g[18894];
assign g[35279] = a[14] & g[18895];
assign g[51662] = b[14] & g[18895];
assign g[35280] = a[14] & g[18896];
assign g[51663] = b[14] & g[18896];
assign g[35281] = a[14] & g[18897];
assign g[51664] = b[14] & g[18897];
assign g[35282] = a[14] & g[18898];
assign g[51665] = b[14] & g[18898];
assign g[35283] = a[14] & g[18899];
assign g[51666] = b[14] & g[18899];
assign g[35284] = a[14] & g[18900];
assign g[51667] = b[14] & g[18900];
assign g[35285] = a[14] & g[18901];
assign g[51668] = b[14] & g[18901];
assign g[35286] = a[14] & g[18902];
assign g[51669] = b[14] & g[18902];
assign g[35287] = a[14] & g[18903];
assign g[51670] = b[14] & g[18903];
assign g[35288] = a[14] & g[18904];
assign g[51671] = b[14] & g[18904];
assign g[35289] = a[14] & g[18905];
assign g[51672] = b[14] & g[18905];
assign g[35290] = a[14] & g[18906];
assign g[51673] = b[14] & g[18906];
assign g[35291] = a[14] & g[18907];
assign g[51674] = b[14] & g[18907];
assign g[35292] = a[14] & g[18908];
assign g[51675] = b[14] & g[18908];
assign g[35293] = a[14] & g[18909];
assign g[51676] = b[14] & g[18909];
assign g[35294] = a[14] & g[18910];
assign g[51677] = b[14] & g[18910];
assign g[35295] = a[14] & g[18911];
assign g[51678] = b[14] & g[18911];
assign g[35296] = a[14] & g[18912];
assign g[51679] = b[14] & g[18912];
assign g[35297] = a[14] & g[18913];
assign g[51680] = b[14] & g[18913];
assign g[35298] = a[14] & g[18914];
assign g[51681] = b[14] & g[18914];
assign g[35299] = a[14] & g[18915];
assign g[51682] = b[14] & g[18915];
assign g[35300] = a[14] & g[18916];
assign g[51683] = b[14] & g[18916];
assign g[35301] = a[14] & g[18917];
assign g[51684] = b[14] & g[18917];
assign g[35302] = a[14] & g[18918];
assign g[51685] = b[14] & g[18918];
assign g[35303] = a[14] & g[18919];
assign g[51686] = b[14] & g[18919];
assign g[35304] = a[14] & g[18920];
assign g[51687] = b[14] & g[18920];
assign g[35305] = a[14] & g[18921];
assign g[51688] = b[14] & g[18921];
assign g[35306] = a[14] & g[18922];
assign g[51689] = b[14] & g[18922];
assign g[35307] = a[14] & g[18923];
assign g[51690] = b[14] & g[18923];
assign g[35308] = a[14] & g[18924];
assign g[51691] = b[14] & g[18924];
assign g[35309] = a[14] & g[18925];
assign g[51692] = b[14] & g[18925];
assign g[35310] = a[14] & g[18926];
assign g[51693] = b[14] & g[18926];
assign g[35311] = a[14] & g[18927];
assign g[51694] = b[14] & g[18927];
assign g[35312] = a[14] & g[18928];
assign g[51695] = b[14] & g[18928];
assign g[35313] = a[14] & g[18929];
assign g[51696] = b[14] & g[18929];
assign g[35314] = a[14] & g[18930];
assign g[51697] = b[14] & g[18930];
assign g[35315] = a[14] & g[18931];
assign g[51698] = b[14] & g[18931];
assign g[35316] = a[14] & g[18932];
assign g[51699] = b[14] & g[18932];
assign g[35317] = a[14] & g[18933];
assign g[51700] = b[14] & g[18933];
assign g[35318] = a[14] & g[18934];
assign g[51701] = b[14] & g[18934];
assign g[35319] = a[14] & g[18935];
assign g[51702] = b[14] & g[18935];
assign g[35320] = a[14] & g[18936];
assign g[51703] = b[14] & g[18936];
assign g[35321] = a[14] & g[18937];
assign g[51704] = b[14] & g[18937];
assign g[35322] = a[14] & g[18938];
assign g[51705] = b[14] & g[18938];
assign g[35323] = a[14] & g[18939];
assign g[51706] = b[14] & g[18939];
assign g[35324] = a[14] & g[18940];
assign g[51707] = b[14] & g[18940];
assign g[35325] = a[14] & g[18941];
assign g[51708] = b[14] & g[18941];
assign g[35326] = a[14] & g[18942];
assign g[51709] = b[14] & g[18942];
assign g[35327] = a[14] & g[18943];
assign g[51710] = b[14] & g[18943];
assign g[35328] = a[14] & g[18944];
assign g[51711] = b[14] & g[18944];
assign g[35329] = a[14] & g[18945];
assign g[51712] = b[14] & g[18945];
assign g[35330] = a[14] & g[18946];
assign g[51713] = b[14] & g[18946];
assign g[35331] = a[14] & g[18947];
assign g[51714] = b[14] & g[18947];
assign g[35332] = a[14] & g[18948];
assign g[51715] = b[14] & g[18948];
assign g[35333] = a[14] & g[18949];
assign g[51716] = b[14] & g[18949];
assign g[35334] = a[14] & g[18950];
assign g[51717] = b[14] & g[18950];
assign g[35335] = a[14] & g[18951];
assign g[51718] = b[14] & g[18951];
assign g[35336] = a[14] & g[18952];
assign g[51719] = b[14] & g[18952];
assign g[35337] = a[14] & g[18953];
assign g[51720] = b[14] & g[18953];
assign g[35338] = a[14] & g[18954];
assign g[51721] = b[14] & g[18954];
assign g[35339] = a[14] & g[18955];
assign g[51722] = b[14] & g[18955];
assign g[35340] = a[14] & g[18956];
assign g[51723] = b[14] & g[18956];
assign g[35341] = a[14] & g[18957];
assign g[51724] = b[14] & g[18957];
assign g[35342] = a[14] & g[18958];
assign g[51725] = b[14] & g[18958];
assign g[35343] = a[14] & g[18959];
assign g[51726] = b[14] & g[18959];
assign g[35344] = a[14] & g[18960];
assign g[51727] = b[14] & g[18960];
assign g[35345] = a[14] & g[18961];
assign g[51728] = b[14] & g[18961];
assign g[35346] = a[14] & g[18962];
assign g[51729] = b[14] & g[18962];
assign g[35347] = a[14] & g[18963];
assign g[51730] = b[14] & g[18963];
assign g[35348] = a[14] & g[18964];
assign g[51731] = b[14] & g[18964];
assign g[35349] = a[14] & g[18965];
assign g[51732] = b[14] & g[18965];
assign g[35350] = a[14] & g[18966];
assign g[51733] = b[14] & g[18966];
assign g[35351] = a[14] & g[18967];
assign g[51734] = b[14] & g[18967];
assign g[35352] = a[14] & g[18968];
assign g[51735] = b[14] & g[18968];
assign g[35353] = a[14] & g[18969];
assign g[51736] = b[14] & g[18969];
assign g[35354] = a[14] & g[18970];
assign g[51737] = b[14] & g[18970];
assign g[35355] = a[14] & g[18971];
assign g[51738] = b[14] & g[18971];
assign g[35356] = a[14] & g[18972];
assign g[51739] = b[14] & g[18972];
assign g[35357] = a[14] & g[18973];
assign g[51740] = b[14] & g[18973];
assign g[35358] = a[14] & g[18974];
assign g[51741] = b[14] & g[18974];
assign g[35359] = a[14] & g[18975];
assign g[51742] = b[14] & g[18975];
assign g[35360] = a[14] & g[18976];
assign g[51743] = b[14] & g[18976];
assign g[35361] = a[14] & g[18977];
assign g[51744] = b[14] & g[18977];
assign g[35362] = a[14] & g[18978];
assign g[51745] = b[14] & g[18978];
assign g[35363] = a[14] & g[18979];
assign g[51746] = b[14] & g[18979];
assign g[35364] = a[14] & g[18980];
assign g[51747] = b[14] & g[18980];
assign g[35365] = a[14] & g[18981];
assign g[51748] = b[14] & g[18981];
assign g[35366] = a[14] & g[18982];
assign g[51749] = b[14] & g[18982];
assign g[35367] = a[14] & g[18983];
assign g[51750] = b[14] & g[18983];
assign g[35368] = a[14] & g[18984];
assign g[51751] = b[14] & g[18984];
assign g[35369] = a[14] & g[18985];
assign g[51752] = b[14] & g[18985];
assign g[35370] = a[14] & g[18986];
assign g[51753] = b[14] & g[18986];
assign g[35371] = a[14] & g[18987];
assign g[51754] = b[14] & g[18987];
assign g[35372] = a[14] & g[18988];
assign g[51755] = b[14] & g[18988];
assign g[35373] = a[14] & g[18989];
assign g[51756] = b[14] & g[18989];
assign g[35374] = a[14] & g[18990];
assign g[51757] = b[14] & g[18990];
assign g[35375] = a[14] & g[18991];
assign g[51758] = b[14] & g[18991];
assign g[35376] = a[14] & g[18992];
assign g[51759] = b[14] & g[18992];
assign g[35377] = a[14] & g[18993];
assign g[51760] = b[14] & g[18993];
assign g[35378] = a[14] & g[18994];
assign g[51761] = b[14] & g[18994];
assign g[35379] = a[14] & g[18995];
assign g[51762] = b[14] & g[18995];
assign g[35380] = a[14] & g[18996];
assign g[51763] = b[14] & g[18996];
assign g[35381] = a[14] & g[18997];
assign g[51764] = b[14] & g[18997];
assign g[35382] = a[14] & g[18998];
assign g[51765] = b[14] & g[18998];
assign g[35383] = a[14] & g[18999];
assign g[51766] = b[14] & g[18999];
assign g[35384] = a[14] & g[19000];
assign g[51767] = b[14] & g[19000];
assign g[35385] = a[14] & g[19001];
assign g[51768] = b[14] & g[19001];
assign g[35386] = a[14] & g[19002];
assign g[51769] = b[14] & g[19002];
assign g[35387] = a[14] & g[19003];
assign g[51770] = b[14] & g[19003];
assign g[35388] = a[14] & g[19004];
assign g[51771] = b[14] & g[19004];
assign g[35389] = a[14] & g[19005];
assign g[51772] = b[14] & g[19005];
assign g[35390] = a[14] & g[19006];
assign g[51773] = b[14] & g[19006];
assign g[35391] = a[14] & g[19007];
assign g[51774] = b[14] & g[19007];
assign g[35392] = a[14] & g[19008];
assign g[51775] = b[14] & g[19008];
assign g[35393] = a[14] & g[19009];
assign g[51776] = b[14] & g[19009];
assign g[35394] = a[14] & g[19010];
assign g[51777] = b[14] & g[19010];
assign g[35395] = a[14] & g[19011];
assign g[51778] = b[14] & g[19011];
assign g[35396] = a[14] & g[19012];
assign g[51779] = b[14] & g[19012];
assign g[35397] = a[14] & g[19013];
assign g[51780] = b[14] & g[19013];
assign g[35398] = a[14] & g[19014];
assign g[51781] = b[14] & g[19014];
assign g[35399] = a[14] & g[19015];
assign g[51782] = b[14] & g[19015];
assign g[35400] = a[14] & g[19016];
assign g[51783] = b[14] & g[19016];
assign g[35401] = a[14] & g[19017];
assign g[51784] = b[14] & g[19017];
assign g[35402] = a[14] & g[19018];
assign g[51785] = b[14] & g[19018];
assign g[35403] = a[14] & g[19019];
assign g[51786] = b[14] & g[19019];
assign g[35404] = a[14] & g[19020];
assign g[51787] = b[14] & g[19020];
assign g[35405] = a[14] & g[19021];
assign g[51788] = b[14] & g[19021];
assign g[35406] = a[14] & g[19022];
assign g[51789] = b[14] & g[19022];
assign g[35407] = a[14] & g[19023];
assign g[51790] = b[14] & g[19023];
assign g[35408] = a[14] & g[19024];
assign g[51791] = b[14] & g[19024];
assign g[35409] = a[14] & g[19025];
assign g[51792] = b[14] & g[19025];
assign g[35410] = a[14] & g[19026];
assign g[51793] = b[14] & g[19026];
assign g[35411] = a[14] & g[19027];
assign g[51794] = b[14] & g[19027];
assign g[35412] = a[14] & g[19028];
assign g[51795] = b[14] & g[19028];
assign g[35413] = a[14] & g[19029];
assign g[51796] = b[14] & g[19029];
assign g[35414] = a[14] & g[19030];
assign g[51797] = b[14] & g[19030];
assign g[35415] = a[14] & g[19031];
assign g[51798] = b[14] & g[19031];
assign g[35416] = a[14] & g[19032];
assign g[51799] = b[14] & g[19032];
assign g[35417] = a[14] & g[19033];
assign g[51800] = b[14] & g[19033];
assign g[35418] = a[14] & g[19034];
assign g[51801] = b[14] & g[19034];
assign g[35419] = a[14] & g[19035];
assign g[51802] = b[14] & g[19035];
assign g[35420] = a[14] & g[19036];
assign g[51803] = b[14] & g[19036];
assign g[35421] = a[14] & g[19037];
assign g[51804] = b[14] & g[19037];
assign g[35422] = a[14] & g[19038];
assign g[51805] = b[14] & g[19038];
assign g[35423] = a[14] & g[19039];
assign g[51806] = b[14] & g[19039];
assign g[35424] = a[14] & g[19040];
assign g[51807] = b[14] & g[19040];
assign g[35425] = a[14] & g[19041];
assign g[51808] = b[14] & g[19041];
assign g[35426] = a[14] & g[19042];
assign g[51809] = b[14] & g[19042];
assign g[35427] = a[14] & g[19043];
assign g[51810] = b[14] & g[19043];
assign g[35428] = a[14] & g[19044];
assign g[51811] = b[14] & g[19044];
assign g[35429] = a[14] & g[19045];
assign g[51812] = b[14] & g[19045];
assign g[35430] = a[14] & g[19046];
assign g[51813] = b[14] & g[19046];
assign g[35431] = a[14] & g[19047];
assign g[51814] = b[14] & g[19047];
assign g[35432] = a[14] & g[19048];
assign g[51815] = b[14] & g[19048];
assign g[35433] = a[14] & g[19049];
assign g[51816] = b[14] & g[19049];
assign g[35434] = a[14] & g[19050];
assign g[51817] = b[14] & g[19050];
assign g[35435] = a[14] & g[19051];
assign g[51818] = b[14] & g[19051];
assign g[35436] = a[14] & g[19052];
assign g[51819] = b[14] & g[19052];
assign g[35437] = a[14] & g[19053];
assign g[51820] = b[14] & g[19053];
assign g[35438] = a[14] & g[19054];
assign g[51821] = b[14] & g[19054];
assign g[35439] = a[14] & g[19055];
assign g[51822] = b[14] & g[19055];
assign g[35440] = a[14] & g[19056];
assign g[51823] = b[14] & g[19056];
assign g[35441] = a[14] & g[19057];
assign g[51824] = b[14] & g[19057];
assign g[35442] = a[14] & g[19058];
assign g[51825] = b[14] & g[19058];
assign g[35443] = a[14] & g[19059];
assign g[51826] = b[14] & g[19059];
assign g[35444] = a[14] & g[19060];
assign g[51827] = b[14] & g[19060];
assign g[35445] = a[14] & g[19061];
assign g[51828] = b[14] & g[19061];
assign g[35446] = a[14] & g[19062];
assign g[51829] = b[14] & g[19062];
assign g[35447] = a[14] & g[19063];
assign g[51830] = b[14] & g[19063];
assign g[35448] = a[14] & g[19064];
assign g[51831] = b[14] & g[19064];
assign g[35449] = a[14] & g[19065];
assign g[51832] = b[14] & g[19065];
assign g[35450] = a[14] & g[19066];
assign g[51833] = b[14] & g[19066];
assign g[35451] = a[14] & g[19067];
assign g[51834] = b[14] & g[19067];
assign g[35452] = a[14] & g[19068];
assign g[51835] = b[14] & g[19068];
assign g[35453] = a[14] & g[19069];
assign g[51836] = b[14] & g[19069];
assign g[35454] = a[14] & g[19070];
assign g[51837] = b[14] & g[19070];
assign g[35455] = a[14] & g[19071];
assign g[51838] = b[14] & g[19071];
assign g[35456] = a[14] & g[19072];
assign g[51839] = b[14] & g[19072];
assign g[35457] = a[14] & g[19073];
assign g[51840] = b[14] & g[19073];
assign g[35458] = a[14] & g[19074];
assign g[51841] = b[14] & g[19074];
assign g[35459] = a[14] & g[19075];
assign g[51842] = b[14] & g[19075];
assign g[35460] = a[14] & g[19076];
assign g[51843] = b[14] & g[19076];
assign g[35461] = a[14] & g[19077];
assign g[51844] = b[14] & g[19077];
assign g[35462] = a[14] & g[19078];
assign g[51845] = b[14] & g[19078];
assign g[35463] = a[14] & g[19079];
assign g[51846] = b[14] & g[19079];
assign g[35464] = a[14] & g[19080];
assign g[51847] = b[14] & g[19080];
assign g[35465] = a[14] & g[19081];
assign g[51848] = b[14] & g[19081];
assign g[35466] = a[14] & g[19082];
assign g[51849] = b[14] & g[19082];
assign g[35467] = a[14] & g[19083];
assign g[51850] = b[14] & g[19083];
assign g[35468] = a[14] & g[19084];
assign g[51851] = b[14] & g[19084];
assign g[35469] = a[14] & g[19085];
assign g[51852] = b[14] & g[19085];
assign g[35470] = a[14] & g[19086];
assign g[51853] = b[14] & g[19086];
assign g[35471] = a[14] & g[19087];
assign g[51854] = b[14] & g[19087];
assign g[35472] = a[14] & g[19088];
assign g[51855] = b[14] & g[19088];
assign g[35473] = a[14] & g[19089];
assign g[51856] = b[14] & g[19089];
assign g[35474] = a[14] & g[19090];
assign g[51857] = b[14] & g[19090];
assign g[35475] = a[14] & g[19091];
assign g[51858] = b[14] & g[19091];
assign g[35476] = a[14] & g[19092];
assign g[51859] = b[14] & g[19092];
assign g[35477] = a[14] & g[19093];
assign g[51860] = b[14] & g[19093];
assign g[35478] = a[14] & g[19094];
assign g[51861] = b[14] & g[19094];
assign g[35479] = a[14] & g[19095];
assign g[51862] = b[14] & g[19095];
assign g[35480] = a[14] & g[19096];
assign g[51863] = b[14] & g[19096];
assign g[35481] = a[14] & g[19097];
assign g[51864] = b[14] & g[19097];
assign g[35482] = a[14] & g[19098];
assign g[51865] = b[14] & g[19098];
assign g[35483] = a[14] & g[19099];
assign g[51866] = b[14] & g[19099];
assign g[35484] = a[14] & g[19100];
assign g[51867] = b[14] & g[19100];
assign g[35485] = a[14] & g[19101];
assign g[51868] = b[14] & g[19101];
assign g[35486] = a[14] & g[19102];
assign g[51869] = b[14] & g[19102];
assign g[35487] = a[14] & g[19103];
assign g[51870] = b[14] & g[19103];
assign g[35488] = a[14] & g[19104];
assign g[51871] = b[14] & g[19104];
assign g[35489] = a[14] & g[19105];
assign g[51872] = b[14] & g[19105];
assign g[35490] = a[14] & g[19106];
assign g[51873] = b[14] & g[19106];
assign g[35491] = a[14] & g[19107];
assign g[51874] = b[14] & g[19107];
assign g[35492] = a[14] & g[19108];
assign g[51875] = b[14] & g[19108];
assign g[35493] = a[14] & g[19109];
assign g[51876] = b[14] & g[19109];
assign g[35494] = a[14] & g[19110];
assign g[51877] = b[14] & g[19110];
assign g[35495] = a[14] & g[19111];
assign g[51878] = b[14] & g[19111];
assign g[35496] = a[14] & g[19112];
assign g[51879] = b[14] & g[19112];
assign g[35497] = a[14] & g[19113];
assign g[51880] = b[14] & g[19113];
assign g[35498] = a[14] & g[19114];
assign g[51881] = b[14] & g[19114];
assign g[35499] = a[14] & g[19115];
assign g[51882] = b[14] & g[19115];
assign g[35500] = a[14] & g[19116];
assign g[51883] = b[14] & g[19116];
assign g[35501] = a[14] & g[19117];
assign g[51884] = b[14] & g[19117];
assign g[35502] = a[14] & g[19118];
assign g[51885] = b[14] & g[19118];
assign g[35503] = a[14] & g[19119];
assign g[51886] = b[14] & g[19119];
assign g[35504] = a[14] & g[19120];
assign g[51887] = b[14] & g[19120];
assign g[35505] = a[14] & g[19121];
assign g[51888] = b[14] & g[19121];
assign g[35506] = a[14] & g[19122];
assign g[51889] = b[14] & g[19122];
assign g[35507] = a[14] & g[19123];
assign g[51890] = b[14] & g[19123];
assign g[35508] = a[14] & g[19124];
assign g[51891] = b[14] & g[19124];
assign g[35509] = a[14] & g[19125];
assign g[51892] = b[14] & g[19125];
assign g[35510] = a[14] & g[19126];
assign g[51893] = b[14] & g[19126];
assign g[35511] = a[14] & g[19127];
assign g[51894] = b[14] & g[19127];
assign g[35512] = a[14] & g[19128];
assign g[51895] = b[14] & g[19128];
assign g[35513] = a[14] & g[19129];
assign g[51896] = b[14] & g[19129];
assign g[35514] = a[14] & g[19130];
assign g[51897] = b[14] & g[19130];
assign g[35515] = a[14] & g[19131];
assign g[51898] = b[14] & g[19131];
assign g[35516] = a[14] & g[19132];
assign g[51899] = b[14] & g[19132];
assign g[35517] = a[14] & g[19133];
assign g[51900] = b[14] & g[19133];
assign g[35518] = a[14] & g[19134];
assign g[51901] = b[14] & g[19134];
assign g[35519] = a[14] & g[19135];
assign g[51902] = b[14] & g[19135];
assign g[35520] = a[14] & g[19136];
assign g[51903] = b[14] & g[19136];
assign g[35521] = a[14] & g[19137];
assign g[51904] = b[14] & g[19137];
assign g[35522] = a[14] & g[19138];
assign g[51905] = b[14] & g[19138];
assign g[35523] = a[14] & g[19139];
assign g[51906] = b[14] & g[19139];
assign g[35524] = a[14] & g[19140];
assign g[51907] = b[14] & g[19140];
assign g[35525] = a[14] & g[19141];
assign g[51908] = b[14] & g[19141];
assign g[35526] = a[14] & g[19142];
assign g[51909] = b[14] & g[19142];
assign g[35527] = a[14] & g[19143];
assign g[51910] = b[14] & g[19143];
assign g[35528] = a[14] & g[19144];
assign g[51911] = b[14] & g[19144];
assign g[35529] = a[14] & g[19145];
assign g[51912] = b[14] & g[19145];
assign g[35530] = a[14] & g[19146];
assign g[51913] = b[14] & g[19146];
assign g[35531] = a[14] & g[19147];
assign g[51914] = b[14] & g[19147];
assign g[35532] = a[14] & g[19148];
assign g[51915] = b[14] & g[19148];
assign g[35533] = a[14] & g[19149];
assign g[51916] = b[14] & g[19149];
assign g[35534] = a[14] & g[19150];
assign g[51917] = b[14] & g[19150];
assign g[35535] = a[14] & g[19151];
assign g[51918] = b[14] & g[19151];
assign g[35536] = a[14] & g[19152];
assign g[51919] = b[14] & g[19152];
assign g[35537] = a[14] & g[19153];
assign g[51920] = b[14] & g[19153];
assign g[35538] = a[14] & g[19154];
assign g[51921] = b[14] & g[19154];
assign g[35539] = a[14] & g[19155];
assign g[51922] = b[14] & g[19155];
assign g[35540] = a[14] & g[19156];
assign g[51923] = b[14] & g[19156];
assign g[35541] = a[14] & g[19157];
assign g[51924] = b[14] & g[19157];
assign g[35542] = a[14] & g[19158];
assign g[51925] = b[14] & g[19158];
assign g[35543] = a[14] & g[19159];
assign g[51926] = b[14] & g[19159];
assign g[35544] = a[14] & g[19160];
assign g[51927] = b[14] & g[19160];
assign g[35545] = a[14] & g[19161];
assign g[51928] = b[14] & g[19161];
assign g[35546] = a[14] & g[19162];
assign g[51929] = b[14] & g[19162];
assign g[35547] = a[14] & g[19163];
assign g[51930] = b[14] & g[19163];
assign g[35548] = a[14] & g[19164];
assign g[51931] = b[14] & g[19164];
assign g[35549] = a[14] & g[19165];
assign g[51932] = b[14] & g[19165];
assign g[35550] = a[14] & g[19166];
assign g[51933] = b[14] & g[19166];
assign g[35551] = a[14] & g[19167];
assign g[51934] = b[14] & g[19167];
assign g[35552] = a[14] & g[19168];
assign g[51935] = b[14] & g[19168];
assign g[35553] = a[14] & g[19169];
assign g[51936] = b[14] & g[19169];
assign g[35554] = a[14] & g[19170];
assign g[51937] = b[14] & g[19170];
assign g[35555] = a[14] & g[19171];
assign g[51938] = b[14] & g[19171];
assign g[35556] = a[14] & g[19172];
assign g[51939] = b[14] & g[19172];
assign g[35557] = a[14] & g[19173];
assign g[51940] = b[14] & g[19173];
assign g[35558] = a[14] & g[19174];
assign g[51941] = b[14] & g[19174];
assign g[35559] = a[14] & g[19175];
assign g[51942] = b[14] & g[19175];
assign g[35560] = a[14] & g[19176];
assign g[51943] = b[14] & g[19176];
assign g[35561] = a[14] & g[19177];
assign g[51944] = b[14] & g[19177];
assign g[35562] = a[14] & g[19178];
assign g[51945] = b[14] & g[19178];
assign g[35563] = a[14] & g[19179];
assign g[51946] = b[14] & g[19179];
assign g[35564] = a[14] & g[19180];
assign g[51947] = b[14] & g[19180];
assign g[35565] = a[14] & g[19181];
assign g[51948] = b[14] & g[19181];
assign g[35566] = a[14] & g[19182];
assign g[51949] = b[14] & g[19182];
assign g[35567] = a[14] & g[19183];
assign g[51950] = b[14] & g[19183];
assign g[35568] = a[14] & g[19184];
assign g[51951] = b[14] & g[19184];
assign g[35569] = a[14] & g[19185];
assign g[51952] = b[14] & g[19185];
assign g[35570] = a[14] & g[19186];
assign g[51953] = b[14] & g[19186];
assign g[35571] = a[14] & g[19187];
assign g[51954] = b[14] & g[19187];
assign g[35572] = a[14] & g[19188];
assign g[51955] = b[14] & g[19188];
assign g[35573] = a[14] & g[19189];
assign g[51956] = b[14] & g[19189];
assign g[35574] = a[14] & g[19190];
assign g[51957] = b[14] & g[19190];
assign g[35575] = a[14] & g[19191];
assign g[51958] = b[14] & g[19191];
assign g[35576] = a[14] & g[19192];
assign g[51959] = b[14] & g[19192];
assign g[35577] = a[14] & g[19193];
assign g[51960] = b[14] & g[19193];
assign g[35578] = a[14] & g[19194];
assign g[51961] = b[14] & g[19194];
assign g[35579] = a[14] & g[19195];
assign g[51962] = b[14] & g[19195];
assign g[35580] = a[14] & g[19196];
assign g[51963] = b[14] & g[19196];
assign g[35581] = a[14] & g[19197];
assign g[51964] = b[14] & g[19197];
assign g[35582] = a[14] & g[19198];
assign g[51965] = b[14] & g[19198];
assign g[35583] = a[14] & g[19199];
assign g[51966] = b[14] & g[19199];
assign g[35584] = a[14] & g[19200];
assign g[51967] = b[14] & g[19200];
assign g[35585] = a[14] & g[19201];
assign g[51968] = b[14] & g[19201];
assign g[35586] = a[14] & g[19202];
assign g[51969] = b[14] & g[19202];
assign g[35587] = a[14] & g[19203];
assign g[51970] = b[14] & g[19203];
assign g[35588] = a[14] & g[19204];
assign g[51971] = b[14] & g[19204];
assign g[35589] = a[14] & g[19205];
assign g[51972] = b[14] & g[19205];
assign g[35590] = a[14] & g[19206];
assign g[51973] = b[14] & g[19206];
assign g[35591] = a[14] & g[19207];
assign g[51974] = b[14] & g[19207];
assign g[35592] = a[14] & g[19208];
assign g[51975] = b[14] & g[19208];
assign g[35593] = a[14] & g[19209];
assign g[51976] = b[14] & g[19209];
assign g[35594] = a[14] & g[19210];
assign g[51977] = b[14] & g[19210];
assign g[35595] = a[14] & g[19211];
assign g[51978] = b[14] & g[19211];
assign g[35596] = a[14] & g[19212];
assign g[51979] = b[14] & g[19212];
assign g[35597] = a[14] & g[19213];
assign g[51980] = b[14] & g[19213];
assign g[35598] = a[14] & g[19214];
assign g[51981] = b[14] & g[19214];
assign g[35599] = a[14] & g[19215];
assign g[51982] = b[14] & g[19215];
assign g[35600] = a[14] & g[19216];
assign g[51983] = b[14] & g[19216];
assign g[35601] = a[14] & g[19217];
assign g[51984] = b[14] & g[19217];
assign g[35602] = a[14] & g[19218];
assign g[51985] = b[14] & g[19218];
assign g[35603] = a[14] & g[19219];
assign g[51986] = b[14] & g[19219];
assign g[35604] = a[14] & g[19220];
assign g[51987] = b[14] & g[19220];
assign g[35605] = a[14] & g[19221];
assign g[51988] = b[14] & g[19221];
assign g[35606] = a[14] & g[19222];
assign g[51989] = b[14] & g[19222];
assign g[35607] = a[14] & g[19223];
assign g[51990] = b[14] & g[19223];
assign g[35608] = a[14] & g[19224];
assign g[51991] = b[14] & g[19224];
assign g[35609] = a[14] & g[19225];
assign g[51992] = b[14] & g[19225];
assign g[35610] = a[14] & g[19226];
assign g[51993] = b[14] & g[19226];
assign g[35611] = a[14] & g[19227];
assign g[51994] = b[14] & g[19227];
assign g[35612] = a[14] & g[19228];
assign g[51995] = b[14] & g[19228];
assign g[35613] = a[14] & g[19229];
assign g[51996] = b[14] & g[19229];
assign g[35614] = a[14] & g[19230];
assign g[51997] = b[14] & g[19230];
assign g[35615] = a[14] & g[19231];
assign g[51998] = b[14] & g[19231];
assign g[35616] = a[14] & g[19232];
assign g[51999] = b[14] & g[19232];
assign g[35617] = a[14] & g[19233];
assign g[52000] = b[14] & g[19233];
assign g[35618] = a[14] & g[19234];
assign g[52001] = b[14] & g[19234];
assign g[35619] = a[14] & g[19235];
assign g[52002] = b[14] & g[19235];
assign g[35620] = a[14] & g[19236];
assign g[52003] = b[14] & g[19236];
assign g[35621] = a[14] & g[19237];
assign g[52004] = b[14] & g[19237];
assign g[35622] = a[14] & g[19238];
assign g[52005] = b[14] & g[19238];
assign g[35623] = a[14] & g[19239];
assign g[52006] = b[14] & g[19239];
assign g[35624] = a[14] & g[19240];
assign g[52007] = b[14] & g[19240];
assign g[35625] = a[14] & g[19241];
assign g[52008] = b[14] & g[19241];
assign g[35626] = a[14] & g[19242];
assign g[52009] = b[14] & g[19242];
assign g[35627] = a[14] & g[19243];
assign g[52010] = b[14] & g[19243];
assign g[35628] = a[14] & g[19244];
assign g[52011] = b[14] & g[19244];
assign g[35629] = a[14] & g[19245];
assign g[52012] = b[14] & g[19245];
assign g[35630] = a[14] & g[19246];
assign g[52013] = b[14] & g[19246];
assign g[35631] = a[14] & g[19247];
assign g[52014] = b[14] & g[19247];
assign g[35632] = a[14] & g[19248];
assign g[52015] = b[14] & g[19248];
assign g[35633] = a[14] & g[19249];
assign g[52016] = b[14] & g[19249];
assign g[35634] = a[14] & g[19250];
assign g[52017] = b[14] & g[19250];
assign g[35635] = a[14] & g[19251];
assign g[52018] = b[14] & g[19251];
assign g[35636] = a[14] & g[19252];
assign g[52019] = b[14] & g[19252];
assign g[35637] = a[14] & g[19253];
assign g[52020] = b[14] & g[19253];
assign g[35638] = a[14] & g[19254];
assign g[52021] = b[14] & g[19254];
assign g[35639] = a[14] & g[19255];
assign g[52022] = b[14] & g[19255];
assign g[35640] = a[14] & g[19256];
assign g[52023] = b[14] & g[19256];
assign g[35641] = a[14] & g[19257];
assign g[52024] = b[14] & g[19257];
assign g[35642] = a[14] & g[19258];
assign g[52025] = b[14] & g[19258];
assign g[35643] = a[14] & g[19259];
assign g[52026] = b[14] & g[19259];
assign g[35644] = a[14] & g[19260];
assign g[52027] = b[14] & g[19260];
assign g[35645] = a[14] & g[19261];
assign g[52028] = b[14] & g[19261];
assign g[35646] = a[14] & g[19262];
assign g[52029] = b[14] & g[19262];
assign g[35647] = a[14] & g[19263];
assign g[52030] = b[14] & g[19263];
assign g[35648] = a[14] & g[19264];
assign g[52031] = b[14] & g[19264];
assign g[35649] = a[14] & g[19265];
assign g[52032] = b[14] & g[19265];
assign g[35650] = a[14] & g[19266];
assign g[52033] = b[14] & g[19266];
assign g[35651] = a[14] & g[19267];
assign g[52034] = b[14] & g[19267];
assign g[35652] = a[14] & g[19268];
assign g[52035] = b[14] & g[19268];
assign g[35653] = a[14] & g[19269];
assign g[52036] = b[14] & g[19269];
assign g[35654] = a[14] & g[19270];
assign g[52037] = b[14] & g[19270];
assign g[35655] = a[14] & g[19271];
assign g[52038] = b[14] & g[19271];
assign g[35656] = a[14] & g[19272];
assign g[52039] = b[14] & g[19272];
assign g[35657] = a[14] & g[19273];
assign g[52040] = b[14] & g[19273];
assign g[35658] = a[14] & g[19274];
assign g[52041] = b[14] & g[19274];
assign g[35659] = a[14] & g[19275];
assign g[52042] = b[14] & g[19275];
assign g[35660] = a[14] & g[19276];
assign g[52043] = b[14] & g[19276];
assign g[35661] = a[14] & g[19277];
assign g[52044] = b[14] & g[19277];
assign g[35662] = a[14] & g[19278];
assign g[52045] = b[14] & g[19278];
assign g[35663] = a[14] & g[19279];
assign g[52046] = b[14] & g[19279];
assign g[35664] = a[14] & g[19280];
assign g[52047] = b[14] & g[19280];
assign g[35665] = a[14] & g[19281];
assign g[52048] = b[14] & g[19281];
assign g[35666] = a[14] & g[19282];
assign g[52049] = b[14] & g[19282];
assign g[35667] = a[14] & g[19283];
assign g[52050] = b[14] & g[19283];
assign g[35668] = a[14] & g[19284];
assign g[52051] = b[14] & g[19284];
assign g[35669] = a[14] & g[19285];
assign g[52052] = b[14] & g[19285];
assign g[35670] = a[14] & g[19286];
assign g[52053] = b[14] & g[19286];
assign g[35671] = a[14] & g[19287];
assign g[52054] = b[14] & g[19287];
assign g[35672] = a[14] & g[19288];
assign g[52055] = b[14] & g[19288];
assign g[35673] = a[14] & g[19289];
assign g[52056] = b[14] & g[19289];
assign g[35674] = a[14] & g[19290];
assign g[52057] = b[14] & g[19290];
assign g[35675] = a[14] & g[19291];
assign g[52058] = b[14] & g[19291];
assign g[35676] = a[14] & g[19292];
assign g[52059] = b[14] & g[19292];
assign g[35677] = a[14] & g[19293];
assign g[52060] = b[14] & g[19293];
assign g[35678] = a[14] & g[19294];
assign g[52061] = b[14] & g[19294];
assign g[35679] = a[14] & g[19295];
assign g[52062] = b[14] & g[19295];
assign g[35680] = a[14] & g[19296];
assign g[52063] = b[14] & g[19296];
assign g[35681] = a[14] & g[19297];
assign g[52064] = b[14] & g[19297];
assign g[35682] = a[14] & g[19298];
assign g[52065] = b[14] & g[19298];
assign g[35683] = a[14] & g[19299];
assign g[52066] = b[14] & g[19299];
assign g[35684] = a[14] & g[19300];
assign g[52067] = b[14] & g[19300];
assign g[35685] = a[14] & g[19301];
assign g[52068] = b[14] & g[19301];
assign g[35686] = a[14] & g[19302];
assign g[52069] = b[14] & g[19302];
assign g[35687] = a[14] & g[19303];
assign g[52070] = b[14] & g[19303];
assign g[35688] = a[14] & g[19304];
assign g[52071] = b[14] & g[19304];
assign g[35689] = a[14] & g[19305];
assign g[52072] = b[14] & g[19305];
assign g[35690] = a[14] & g[19306];
assign g[52073] = b[14] & g[19306];
assign g[35691] = a[14] & g[19307];
assign g[52074] = b[14] & g[19307];
assign g[35692] = a[14] & g[19308];
assign g[52075] = b[14] & g[19308];
assign g[35693] = a[14] & g[19309];
assign g[52076] = b[14] & g[19309];
assign g[35694] = a[14] & g[19310];
assign g[52077] = b[14] & g[19310];
assign g[35695] = a[14] & g[19311];
assign g[52078] = b[14] & g[19311];
assign g[35696] = a[14] & g[19312];
assign g[52079] = b[14] & g[19312];
assign g[35697] = a[14] & g[19313];
assign g[52080] = b[14] & g[19313];
assign g[35698] = a[14] & g[19314];
assign g[52081] = b[14] & g[19314];
assign g[35699] = a[14] & g[19315];
assign g[52082] = b[14] & g[19315];
assign g[35700] = a[14] & g[19316];
assign g[52083] = b[14] & g[19316];
assign g[35701] = a[14] & g[19317];
assign g[52084] = b[14] & g[19317];
assign g[35702] = a[14] & g[19318];
assign g[52085] = b[14] & g[19318];
assign g[35703] = a[14] & g[19319];
assign g[52086] = b[14] & g[19319];
assign g[35704] = a[14] & g[19320];
assign g[52087] = b[14] & g[19320];
assign g[35705] = a[14] & g[19321];
assign g[52088] = b[14] & g[19321];
assign g[35706] = a[14] & g[19322];
assign g[52089] = b[14] & g[19322];
assign g[35707] = a[14] & g[19323];
assign g[52090] = b[14] & g[19323];
assign g[35708] = a[14] & g[19324];
assign g[52091] = b[14] & g[19324];
assign g[35709] = a[14] & g[19325];
assign g[52092] = b[14] & g[19325];
assign g[35710] = a[14] & g[19326];
assign g[52093] = b[14] & g[19326];
assign g[35711] = a[14] & g[19327];
assign g[52094] = b[14] & g[19327];
assign g[35712] = a[14] & g[19328];
assign g[52095] = b[14] & g[19328];
assign g[35713] = a[14] & g[19329];
assign g[52096] = b[14] & g[19329];
assign g[35714] = a[14] & g[19330];
assign g[52097] = b[14] & g[19330];
assign g[35715] = a[14] & g[19331];
assign g[52098] = b[14] & g[19331];
assign g[35716] = a[14] & g[19332];
assign g[52099] = b[14] & g[19332];
assign g[35717] = a[14] & g[19333];
assign g[52100] = b[14] & g[19333];
assign g[35718] = a[14] & g[19334];
assign g[52101] = b[14] & g[19334];
assign g[35719] = a[14] & g[19335];
assign g[52102] = b[14] & g[19335];
assign g[35720] = a[14] & g[19336];
assign g[52103] = b[14] & g[19336];
assign g[35721] = a[14] & g[19337];
assign g[52104] = b[14] & g[19337];
assign g[35722] = a[14] & g[19338];
assign g[52105] = b[14] & g[19338];
assign g[35723] = a[14] & g[19339];
assign g[52106] = b[14] & g[19339];
assign g[35724] = a[14] & g[19340];
assign g[52107] = b[14] & g[19340];
assign g[35725] = a[14] & g[19341];
assign g[52108] = b[14] & g[19341];
assign g[35726] = a[14] & g[19342];
assign g[52109] = b[14] & g[19342];
assign g[35727] = a[14] & g[19343];
assign g[52110] = b[14] & g[19343];
assign g[35728] = a[14] & g[19344];
assign g[52111] = b[14] & g[19344];
assign g[35729] = a[14] & g[19345];
assign g[52112] = b[14] & g[19345];
assign g[35730] = a[14] & g[19346];
assign g[52113] = b[14] & g[19346];
assign g[35731] = a[14] & g[19347];
assign g[52114] = b[14] & g[19347];
assign g[35732] = a[14] & g[19348];
assign g[52115] = b[14] & g[19348];
assign g[35733] = a[14] & g[19349];
assign g[52116] = b[14] & g[19349];
assign g[35734] = a[14] & g[19350];
assign g[52117] = b[14] & g[19350];
assign g[35735] = a[14] & g[19351];
assign g[52118] = b[14] & g[19351];
assign g[35736] = a[14] & g[19352];
assign g[52119] = b[14] & g[19352];
assign g[35737] = a[14] & g[19353];
assign g[52120] = b[14] & g[19353];
assign g[35738] = a[14] & g[19354];
assign g[52121] = b[14] & g[19354];
assign g[35739] = a[14] & g[19355];
assign g[52122] = b[14] & g[19355];
assign g[35740] = a[14] & g[19356];
assign g[52123] = b[14] & g[19356];
assign g[35741] = a[14] & g[19357];
assign g[52124] = b[14] & g[19357];
assign g[35742] = a[14] & g[19358];
assign g[52125] = b[14] & g[19358];
assign g[35743] = a[14] & g[19359];
assign g[52126] = b[14] & g[19359];
assign g[35744] = a[14] & g[19360];
assign g[52127] = b[14] & g[19360];
assign g[35745] = a[14] & g[19361];
assign g[52128] = b[14] & g[19361];
assign g[35746] = a[14] & g[19362];
assign g[52129] = b[14] & g[19362];
assign g[35747] = a[14] & g[19363];
assign g[52130] = b[14] & g[19363];
assign g[35748] = a[14] & g[19364];
assign g[52131] = b[14] & g[19364];
assign g[35749] = a[14] & g[19365];
assign g[52132] = b[14] & g[19365];
assign g[35750] = a[14] & g[19366];
assign g[52133] = b[14] & g[19366];
assign g[35751] = a[14] & g[19367];
assign g[52134] = b[14] & g[19367];
assign g[35752] = a[14] & g[19368];
assign g[52135] = b[14] & g[19368];
assign g[35753] = a[14] & g[19369];
assign g[52136] = b[14] & g[19369];
assign g[35754] = a[14] & g[19370];
assign g[52137] = b[14] & g[19370];
assign g[35755] = a[14] & g[19371];
assign g[52138] = b[14] & g[19371];
assign g[35756] = a[14] & g[19372];
assign g[52139] = b[14] & g[19372];
assign g[35757] = a[14] & g[19373];
assign g[52140] = b[14] & g[19373];
assign g[35758] = a[14] & g[19374];
assign g[52141] = b[14] & g[19374];
assign g[35759] = a[14] & g[19375];
assign g[52142] = b[14] & g[19375];
assign g[35760] = a[14] & g[19376];
assign g[52143] = b[14] & g[19376];
assign g[35761] = a[14] & g[19377];
assign g[52144] = b[14] & g[19377];
assign g[35762] = a[14] & g[19378];
assign g[52145] = b[14] & g[19378];
assign g[35763] = a[14] & g[19379];
assign g[52146] = b[14] & g[19379];
assign g[35764] = a[14] & g[19380];
assign g[52147] = b[14] & g[19380];
assign g[35765] = a[14] & g[19381];
assign g[52148] = b[14] & g[19381];
assign g[35766] = a[14] & g[19382];
assign g[52149] = b[14] & g[19382];
assign g[35767] = a[14] & g[19383];
assign g[52150] = b[14] & g[19383];
assign g[35768] = a[14] & g[19384];
assign g[52151] = b[14] & g[19384];
assign g[35769] = a[14] & g[19385];
assign g[52152] = b[14] & g[19385];
assign g[35770] = a[14] & g[19386];
assign g[52153] = b[14] & g[19386];
assign g[35771] = a[14] & g[19387];
assign g[52154] = b[14] & g[19387];
assign g[35772] = a[14] & g[19388];
assign g[52155] = b[14] & g[19388];
assign g[35773] = a[14] & g[19389];
assign g[52156] = b[14] & g[19389];
assign g[35774] = a[14] & g[19390];
assign g[52157] = b[14] & g[19390];
assign g[35775] = a[14] & g[19391];
assign g[52158] = b[14] & g[19391];
assign g[35776] = a[14] & g[19392];
assign g[52159] = b[14] & g[19392];
assign g[35777] = a[14] & g[19393];
assign g[52160] = b[14] & g[19393];
assign g[35778] = a[14] & g[19394];
assign g[52161] = b[14] & g[19394];
assign g[35779] = a[14] & g[19395];
assign g[52162] = b[14] & g[19395];
assign g[35780] = a[14] & g[19396];
assign g[52163] = b[14] & g[19396];
assign g[35781] = a[14] & g[19397];
assign g[52164] = b[14] & g[19397];
assign g[35782] = a[14] & g[19398];
assign g[52165] = b[14] & g[19398];
assign g[35783] = a[14] & g[19399];
assign g[52166] = b[14] & g[19399];
assign g[35784] = a[14] & g[19400];
assign g[52167] = b[14] & g[19400];
assign g[35785] = a[14] & g[19401];
assign g[52168] = b[14] & g[19401];
assign g[35786] = a[14] & g[19402];
assign g[52169] = b[14] & g[19402];
assign g[35787] = a[14] & g[19403];
assign g[52170] = b[14] & g[19403];
assign g[35788] = a[14] & g[19404];
assign g[52171] = b[14] & g[19404];
assign g[35789] = a[14] & g[19405];
assign g[52172] = b[14] & g[19405];
assign g[35790] = a[14] & g[19406];
assign g[52173] = b[14] & g[19406];
assign g[35791] = a[14] & g[19407];
assign g[52174] = b[14] & g[19407];
assign g[35792] = a[14] & g[19408];
assign g[52175] = b[14] & g[19408];
assign g[35793] = a[14] & g[19409];
assign g[52176] = b[14] & g[19409];
assign g[35794] = a[14] & g[19410];
assign g[52177] = b[14] & g[19410];
assign g[35795] = a[14] & g[19411];
assign g[52178] = b[14] & g[19411];
assign g[35796] = a[14] & g[19412];
assign g[52179] = b[14] & g[19412];
assign g[35797] = a[14] & g[19413];
assign g[52180] = b[14] & g[19413];
assign g[35798] = a[14] & g[19414];
assign g[52181] = b[14] & g[19414];
assign g[35799] = a[14] & g[19415];
assign g[52182] = b[14] & g[19415];
assign g[35800] = a[14] & g[19416];
assign g[52183] = b[14] & g[19416];
assign g[35801] = a[14] & g[19417];
assign g[52184] = b[14] & g[19417];
assign g[35802] = a[14] & g[19418];
assign g[52185] = b[14] & g[19418];
assign g[35803] = a[14] & g[19419];
assign g[52186] = b[14] & g[19419];
assign g[35804] = a[14] & g[19420];
assign g[52187] = b[14] & g[19420];
assign g[35805] = a[14] & g[19421];
assign g[52188] = b[14] & g[19421];
assign g[35806] = a[14] & g[19422];
assign g[52189] = b[14] & g[19422];
assign g[35807] = a[14] & g[19423];
assign g[52190] = b[14] & g[19423];
assign g[35808] = a[14] & g[19424];
assign g[52191] = b[14] & g[19424];
assign g[35809] = a[14] & g[19425];
assign g[52192] = b[14] & g[19425];
assign g[35810] = a[14] & g[19426];
assign g[52193] = b[14] & g[19426];
assign g[35811] = a[14] & g[19427];
assign g[52194] = b[14] & g[19427];
assign g[35812] = a[14] & g[19428];
assign g[52195] = b[14] & g[19428];
assign g[35813] = a[14] & g[19429];
assign g[52196] = b[14] & g[19429];
assign g[35814] = a[14] & g[19430];
assign g[52197] = b[14] & g[19430];
assign g[35815] = a[14] & g[19431];
assign g[52198] = b[14] & g[19431];
assign g[35816] = a[14] & g[19432];
assign g[52199] = b[14] & g[19432];
assign g[35817] = a[14] & g[19433];
assign g[52200] = b[14] & g[19433];
assign g[35818] = a[14] & g[19434];
assign g[52201] = b[14] & g[19434];
assign g[35819] = a[14] & g[19435];
assign g[52202] = b[14] & g[19435];
assign g[35820] = a[14] & g[19436];
assign g[52203] = b[14] & g[19436];
assign g[35821] = a[14] & g[19437];
assign g[52204] = b[14] & g[19437];
assign g[35822] = a[14] & g[19438];
assign g[52205] = b[14] & g[19438];
assign g[35823] = a[14] & g[19439];
assign g[52206] = b[14] & g[19439];
assign g[35824] = a[14] & g[19440];
assign g[52207] = b[14] & g[19440];
assign g[35825] = a[14] & g[19441];
assign g[52208] = b[14] & g[19441];
assign g[35826] = a[14] & g[19442];
assign g[52209] = b[14] & g[19442];
assign g[35827] = a[14] & g[19443];
assign g[52210] = b[14] & g[19443];
assign g[35828] = a[14] & g[19444];
assign g[52211] = b[14] & g[19444];
assign g[35829] = a[14] & g[19445];
assign g[52212] = b[14] & g[19445];
assign g[35830] = a[14] & g[19446];
assign g[52213] = b[14] & g[19446];
assign g[35831] = a[14] & g[19447];
assign g[52214] = b[14] & g[19447];
assign g[35832] = a[14] & g[19448];
assign g[52215] = b[14] & g[19448];
assign g[35833] = a[14] & g[19449];
assign g[52216] = b[14] & g[19449];
assign g[35834] = a[14] & g[19450];
assign g[52217] = b[14] & g[19450];
assign g[35835] = a[14] & g[19451];
assign g[52218] = b[14] & g[19451];
assign g[35836] = a[14] & g[19452];
assign g[52219] = b[14] & g[19452];
assign g[35837] = a[14] & g[19453];
assign g[52220] = b[14] & g[19453];
assign g[35838] = a[14] & g[19454];
assign g[52221] = b[14] & g[19454];
assign g[35839] = a[14] & g[19455];
assign g[52222] = b[14] & g[19455];
assign g[35840] = a[14] & g[19456];
assign g[52223] = b[14] & g[19456];
assign g[35841] = a[14] & g[19457];
assign g[52224] = b[14] & g[19457];
assign g[35842] = a[14] & g[19458];
assign g[52225] = b[14] & g[19458];
assign g[35843] = a[14] & g[19459];
assign g[52226] = b[14] & g[19459];
assign g[35844] = a[14] & g[19460];
assign g[52227] = b[14] & g[19460];
assign g[35845] = a[14] & g[19461];
assign g[52228] = b[14] & g[19461];
assign g[35846] = a[14] & g[19462];
assign g[52229] = b[14] & g[19462];
assign g[35847] = a[14] & g[19463];
assign g[52230] = b[14] & g[19463];
assign g[35848] = a[14] & g[19464];
assign g[52231] = b[14] & g[19464];
assign g[35849] = a[14] & g[19465];
assign g[52232] = b[14] & g[19465];
assign g[35850] = a[14] & g[19466];
assign g[52233] = b[14] & g[19466];
assign g[35851] = a[14] & g[19467];
assign g[52234] = b[14] & g[19467];
assign g[35852] = a[14] & g[19468];
assign g[52235] = b[14] & g[19468];
assign g[35853] = a[14] & g[19469];
assign g[52236] = b[14] & g[19469];
assign g[35854] = a[14] & g[19470];
assign g[52237] = b[14] & g[19470];
assign g[35855] = a[14] & g[19471];
assign g[52238] = b[14] & g[19471];
assign g[35856] = a[14] & g[19472];
assign g[52239] = b[14] & g[19472];
assign g[35857] = a[14] & g[19473];
assign g[52240] = b[14] & g[19473];
assign g[35858] = a[14] & g[19474];
assign g[52241] = b[14] & g[19474];
assign g[35859] = a[14] & g[19475];
assign g[52242] = b[14] & g[19475];
assign g[35860] = a[14] & g[19476];
assign g[52243] = b[14] & g[19476];
assign g[35861] = a[14] & g[19477];
assign g[52244] = b[14] & g[19477];
assign g[35862] = a[14] & g[19478];
assign g[52245] = b[14] & g[19478];
assign g[35863] = a[14] & g[19479];
assign g[52246] = b[14] & g[19479];
assign g[35864] = a[14] & g[19480];
assign g[52247] = b[14] & g[19480];
assign g[35865] = a[14] & g[19481];
assign g[52248] = b[14] & g[19481];
assign g[35866] = a[14] & g[19482];
assign g[52249] = b[14] & g[19482];
assign g[35867] = a[14] & g[19483];
assign g[52250] = b[14] & g[19483];
assign g[35868] = a[14] & g[19484];
assign g[52251] = b[14] & g[19484];
assign g[35869] = a[14] & g[19485];
assign g[52252] = b[14] & g[19485];
assign g[35870] = a[14] & g[19486];
assign g[52253] = b[14] & g[19486];
assign g[35871] = a[14] & g[19487];
assign g[52254] = b[14] & g[19487];
assign g[35872] = a[14] & g[19488];
assign g[52255] = b[14] & g[19488];
assign g[35873] = a[14] & g[19489];
assign g[52256] = b[14] & g[19489];
assign g[35874] = a[14] & g[19490];
assign g[52257] = b[14] & g[19490];
assign g[35875] = a[14] & g[19491];
assign g[52258] = b[14] & g[19491];
assign g[35876] = a[14] & g[19492];
assign g[52259] = b[14] & g[19492];
assign g[35877] = a[14] & g[19493];
assign g[52260] = b[14] & g[19493];
assign g[35878] = a[14] & g[19494];
assign g[52261] = b[14] & g[19494];
assign g[35879] = a[14] & g[19495];
assign g[52262] = b[14] & g[19495];
assign g[35880] = a[14] & g[19496];
assign g[52263] = b[14] & g[19496];
assign g[35881] = a[14] & g[19497];
assign g[52264] = b[14] & g[19497];
assign g[35882] = a[14] & g[19498];
assign g[52265] = b[14] & g[19498];
assign g[35883] = a[14] & g[19499];
assign g[52266] = b[14] & g[19499];
assign g[35884] = a[14] & g[19500];
assign g[52267] = b[14] & g[19500];
assign g[35885] = a[14] & g[19501];
assign g[52268] = b[14] & g[19501];
assign g[35886] = a[14] & g[19502];
assign g[52269] = b[14] & g[19502];
assign g[35887] = a[14] & g[19503];
assign g[52270] = b[14] & g[19503];
assign g[35888] = a[14] & g[19504];
assign g[52271] = b[14] & g[19504];
assign g[35889] = a[14] & g[19505];
assign g[52272] = b[14] & g[19505];
assign g[35890] = a[14] & g[19506];
assign g[52273] = b[14] & g[19506];
assign g[35891] = a[14] & g[19507];
assign g[52274] = b[14] & g[19507];
assign g[35892] = a[14] & g[19508];
assign g[52275] = b[14] & g[19508];
assign g[35893] = a[14] & g[19509];
assign g[52276] = b[14] & g[19509];
assign g[35894] = a[14] & g[19510];
assign g[52277] = b[14] & g[19510];
assign g[35895] = a[14] & g[19511];
assign g[52278] = b[14] & g[19511];
assign g[35896] = a[14] & g[19512];
assign g[52279] = b[14] & g[19512];
assign g[35897] = a[14] & g[19513];
assign g[52280] = b[14] & g[19513];
assign g[35898] = a[14] & g[19514];
assign g[52281] = b[14] & g[19514];
assign g[35899] = a[14] & g[19515];
assign g[52282] = b[14] & g[19515];
assign g[35900] = a[14] & g[19516];
assign g[52283] = b[14] & g[19516];
assign g[35901] = a[14] & g[19517];
assign g[52284] = b[14] & g[19517];
assign g[35902] = a[14] & g[19518];
assign g[52285] = b[14] & g[19518];
assign g[35903] = a[14] & g[19519];
assign g[52286] = b[14] & g[19519];
assign g[35904] = a[14] & g[19520];
assign g[52287] = b[14] & g[19520];
assign g[35905] = a[14] & g[19521];
assign g[52288] = b[14] & g[19521];
assign g[35906] = a[14] & g[19522];
assign g[52289] = b[14] & g[19522];
assign g[35907] = a[14] & g[19523];
assign g[52290] = b[14] & g[19523];
assign g[35908] = a[14] & g[19524];
assign g[52291] = b[14] & g[19524];
assign g[35909] = a[14] & g[19525];
assign g[52292] = b[14] & g[19525];
assign g[35910] = a[14] & g[19526];
assign g[52293] = b[14] & g[19526];
assign g[35911] = a[14] & g[19527];
assign g[52294] = b[14] & g[19527];
assign g[35912] = a[14] & g[19528];
assign g[52295] = b[14] & g[19528];
assign g[35913] = a[14] & g[19529];
assign g[52296] = b[14] & g[19529];
assign g[35914] = a[14] & g[19530];
assign g[52297] = b[14] & g[19530];
assign g[35915] = a[14] & g[19531];
assign g[52298] = b[14] & g[19531];
assign g[35916] = a[14] & g[19532];
assign g[52299] = b[14] & g[19532];
assign g[35917] = a[14] & g[19533];
assign g[52300] = b[14] & g[19533];
assign g[35918] = a[14] & g[19534];
assign g[52301] = b[14] & g[19534];
assign g[35919] = a[14] & g[19535];
assign g[52302] = b[14] & g[19535];
assign g[35920] = a[14] & g[19536];
assign g[52303] = b[14] & g[19536];
assign g[35921] = a[14] & g[19537];
assign g[52304] = b[14] & g[19537];
assign g[35922] = a[14] & g[19538];
assign g[52305] = b[14] & g[19538];
assign g[35923] = a[14] & g[19539];
assign g[52306] = b[14] & g[19539];
assign g[35924] = a[14] & g[19540];
assign g[52307] = b[14] & g[19540];
assign g[35925] = a[14] & g[19541];
assign g[52308] = b[14] & g[19541];
assign g[35926] = a[14] & g[19542];
assign g[52309] = b[14] & g[19542];
assign g[35927] = a[14] & g[19543];
assign g[52310] = b[14] & g[19543];
assign g[35928] = a[14] & g[19544];
assign g[52311] = b[14] & g[19544];
assign g[35929] = a[14] & g[19545];
assign g[52312] = b[14] & g[19545];
assign g[35930] = a[14] & g[19546];
assign g[52313] = b[14] & g[19546];
assign g[35931] = a[14] & g[19547];
assign g[52314] = b[14] & g[19547];
assign g[35932] = a[14] & g[19548];
assign g[52315] = b[14] & g[19548];
assign g[35933] = a[14] & g[19549];
assign g[52316] = b[14] & g[19549];
assign g[35934] = a[14] & g[19550];
assign g[52317] = b[14] & g[19550];
assign g[35935] = a[14] & g[19551];
assign g[52318] = b[14] & g[19551];
assign g[35936] = a[14] & g[19552];
assign g[52319] = b[14] & g[19552];
assign g[35937] = a[14] & g[19553];
assign g[52320] = b[14] & g[19553];
assign g[35938] = a[14] & g[19554];
assign g[52321] = b[14] & g[19554];
assign g[35939] = a[14] & g[19555];
assign g[52322] = b[14] & g[19555];
assign g[35940] = a[14] & g[19556];
assign g[52323] = b[14] & g[19556];
assign g[35941] = a[14] & g[19557];
assign g[52324] = b[14] & g[19557];
assign g[35942] = a[14] & g[19558];
assign g[52325] = b[14] & g[19558];
assign g[35943] = a[14] & g[19559];
assign g[52326] = b[14] & g[19559];
assign g[35944] = a[14] & g[19560];
assign g[52327] = b[14] & g[19560];
assign g[35945] = a[14] & g[19561];
assign g[52328] = b[14] & g[19561];
assign g[35946] = a[14] & g[19562];
assign g[52329] = b[14] & g[19562];
assign g[35947] = a[14] & g[19563];
assign g[52330] = b[14] & g[19563];
assign g[35948] = a[14] & g[19564];
assign g[52331] = b[14] & g[19564];
assign g[35949] = a[14] & g[19565];
assign g[52332] = b[14] & g[19565];
assign g[35950] = a[14] & g[19566];
assign g[52333] = b[14] & g[19566];
assign g[35951] = a[14] & g[19567];
assign g[52334] = b[14] & g[19567];
assign g[35952] = a[14] & g[19568];
assign g[52335] = b[14] & g[19568];
assign g[35953] = a[14] & g[19569];
assign g[52336] = b[14] & g[19569];
assign g[35954] = a[14] & g[19570];
assign g[52337] = b[14] & g[19570];
assign g[35955] = a[14] & g[19571];
assign g[52338] = b[14] & g[19571];
assign g[35956] = a[14] & g[19572];
assign g[52339] = b[14] & g[19572];
assign g[35957] = a[14] & g[19573];
assign g[52340] = b[14] & g[19573];
assign g[35958] = a[14] & g[19574];
assign g[52341] = b[14] & g[19574];
assign g[35959] = a[14] & g[19575];
assign g[52342] = b[14] & g[19575];
assign g[35960] = a[14] & g[19576];
assign g[52343] = b[14] & g[19576];
assign g[35961] = a[14] & g[19577];
assign g[52344] = b[14] & g[19577];
assign g[35962] = a[14] & g[19578];
assign g[52345] = b[14] & g[19578];
assign g[35963] = a[14] & g[19579];
assign g[52346] = b[14] & g[19579];
assign g[35964] = a[14] & g[19580];
assign g[52347] = b[14] & g[19580];
assign g[35965] = a[14] & g[19581];
assign g[52348] = b[14] & g[19581];
assign g[35966] = a[14] & g[19582];
assign g[52349] = b[14] & g[19582];
assign g[35967] = a[14] & g[19583];
assign g[52350] = b[14] & g[19583];
assign g[35968] = a[14] & g[19584];
assign g[52351] = b[14] & g[19584];
assign g[35969] = a[14] & g[19585];
assign g[52352] = b[14] & g[19585];
assign g[35970] = a[14] & g[19586];
assign g[52353] = b[14] & g[19586];
assign g[35971] = a[14] & g[19587];
assign g[52354] = b[14] & g[19587];
assign g[35972] = a[14] & g[19588];
assign g[52355] = b[14] & g[19588];
assign g[35973] = a[14] & g[19589];
assign g[52356] = b[14] & g[19589];
assign g[35974] = a[14] & g[19590];
assign g[52357] = b[14] & g[19590];
assign g[35975] = a[14] & g[19591];
assign g[52358] = b[14] & g[19591];
assign g[35976] = a[14] & g[19592];
assign g[52359] = b[14] & g[19592];
assign g[35977] = a[14] & g[19593];
assign g[52360] = b[14] & g[19593];
assign g[35978] = a[14] & g[19594];
assign g[52361] = b[14] & g[19594];
assign g[35979] = a[14] & g[19595];
assign g[52362] = b[14] & g[19595];
assign g[35980] = a[14] & g[19596];
assign g[52363] = b[14] & g[19596];
assign g[35981] = a[14] & g[19597];
assign g[52364] = b[14] & g[19597];
assign g[35982] = a[14] & g[19598];
assign g[52365] = b[14] & g[19598];
assign g[35983] = a[14] & g[19599];
assign g[52366] = b[14] & g[19599];
assign g[35984] = a[14] & g[19600];
assign g[52367] = b[14] & g[19600];
assign g[35985] = a[14] & g[19601];
assign g[52368] = b[14] & g[19601];
assign g[35986] = a[14] & g[19602];
assign g[52369] = b[14] & g[19602];
assign g[35987] = a[14] & g[19603];
assign g[52370] = b[14] & g[19603];
assign g[35988] = a[14] & g[19604];
assign g[52371] = b[14] & g[19604];
assign g[35989] = a[14] & g[19605];
assign g[52372] = b[14] & g[19605];
assign g[35990] = a[14] & g[19606];
assign g[52373] = b[14] & g[19606];
assign g[35991] = a[14] & g[19607];
assign g[52374] = b[14] & g[19607];
assign g[35992] = a[14] & g[19608];
assign g[52375] = b[14] & g[19608];
assign g[35993] = a[14] & g[19609];
assign g[52376] = b[14] & g[19609];
assign g[35994] = a[14] & g[19610];
assign g[52377] = b[14] & g[19610];
assign g[35995] = a[14] & g[19611];
assign g[52378] = b[14] & g[19611];
assign g[35996] = a[14] & g[19612];
assign g[52379] = b[14] & g[19612];
assign g[35997] = a[14] & g[19613];
assign g[52380] = b[14] & g[19613];
assign g[35998] = a[14] & g[19614];
assign g[52381] = b[14] & g[19614];
assign g[35999] = a[14] & g[19615];
assign g[52382] = b[14] & g[19615];
assign g[36000] = a[14] & g[19616];
assign g[52383] = b[14] & g[19616];
assign g[36001] = a[14] & g[19617];
assign g[52384] = b[14] & g[19617];
assign g[36002] = a[14] & g[19618];
assign g[52385] = b[14] & g[19618];
assign g[36003] = a[14] & g[19619];
assign g[52386] = b[14] & g[19619];
assign g[36004] = a[14] & g[19620];
assign g[52387] = b[14] & g[19620];
assign g[36005] = a[14] & g[19621];
assign g[52388] = b[14] & g[19621];
assign g[36006] = a[14] & g[19622];
assign g[52389] = b[14] & g[19622];
assign g[36007] = a[14] & g[19623];
assign g[52390] = b[14] & g[19623];
assign g[36008] = a[14] & g[19624];
assign g[52391] = b[14] & g[19624];
assign g[36009] = a[14] & g[19625];
assign g[52392] = b[14] & g[19625];
assign g[36010] = a[14] & g[19626];
assign g[52393] = b[14] & g[19626];
assign g[36011] = a[14] & g[19627];
assign g[52394] = b[14] & g[19627];
assign g[36012] = a[14] & g[19628];
assign g[52395] = b[14] & g[19628];
assign g[36013] = a[14] & g[19629];
assign g[52396] = b[14] & g[19629];
assign g[36014] = a[14] & g[19630];
assign g[52397] = b[14] & g[19630];
assign g[36015] = a[14] & g[19631];
assign g[52398] = b[14] & g[19631];
assign g[36016] = a[14] & g[19632];
assign g[52399] = b[14] & g[19632];
assign g[36017] = a[14] & g[19633];
assign g[52400] = b[14] & g[19633];
assign g[36018] = a[14] & g[19634];
assign g[52401] = b[14] & g[19634];
assign g[36019] = a[14] & g[19635];
assign g[52402] = b[14] & g[19635];
assign g[36020] = a[14] & g[19636];
assign g[52403] = b[14] & g[19636];
assign g[36021] = a[14] & g[19637];
assign g[52404] = b[14] & g[19637];
assign g[36022] = a[14] & g[19638];
assign g[52405] = b[14] & g[19638];
assign g[36023] = a[14] & g[19639];
assign g[52406] = b[14] & g[19639];
assign g[36024] = a[14] & g[19640];
assign g[52407] = b[14] & g[19640];
assign g[36025] = a[14] & g[19641];
assign g[52408] = b[14] & g[19641];
assign g[36026] = a[14] & g[19642];
assign g[52409] = b[14] & g[19642];
assign g[36027] = a[14] & g[19643];
assign g[52410] = b[14] & g[19643];
assign g[36028] = a[14] & g[19644];
assign g[52411] = b[14] & g[19644];
assign g[36029] = a[14] & g[19645];
assign g[52412] = b[14] & g[19645];
assign g[36030] = a[14] & g[19646];
assign g[52413] = b[14] & g[19646];
assign g[36031] = a[14] & g[19647];
assign g[52414] = b[14] & g[19647];
assign g[36032] = a[14] & g[19648];
assign g[52415] = b[14] & g[19648];
assign g[36033] = a[14] & g[19649];
assign g[52416] = b[14] & g[19649];
assign g[36034] = a[14] & g[19650];
assign g[52417] = b[14] & g[19650];
assign g[36035] = a[14] & g[19651];
assign g[52418] = b[14] & g[19651];
assign g[36036] = a[14] & g[19652];
assign g[52419] = b[14] & g[19652];
assign g[36037] = a[14] & g[19653];
assign g[52420] = b[14] & g[19653];
assign g[36038] = a[14] & g[19654];
assign g[52421] = b[14] & g[19654];
assign g[36039] = a[14] & g[19655];
assign g[52422] = b[14] & g[19655];
assign g[36040] = a[14] & g[19656];
assign g[52423] = b[14] & g[19656];
assign g[36041] = a[14] & g[19657];
assign g[52424] = b[14] & g[19657];
assign g[36042] = a[14] & g[19658];
assign g[52425] = b[14] & g[19658];
assign g[36043] = a[14] & g[19659];
assign g[52426] = b[14] & g[19659];
assign g[36044] = a[14] & g[19660];
assign g[52427] = b[14] & g[19660];
assign g[36045] = a[14] & g[19661];
assign g[52428] = b[14] & g[19661];
assign g[36046] = a[14] & g[19662];
assign g[52429] = b[14] & g[19662];
assign g[36047] = a[14] & g[19663];
assign g[52430] = b[14] & g[19663];
assign g[36048] = a[14] & g[19664];
assign g[52431] = b[14] & g[19664];
assign g[36049] = a[14] & g[19665];
assign g[52432] = b[14] & g[19665];
assign g[36050] = a[14] & g[19666];
assign g[52433] = b[14] & g[19666];
assign g[36051] = a[14] & g[19667];
assign g[52434] = b[14] & g[19667];
assign g[36052] = a[14] & g[19668];
assign g[52435] = b[14] & g[19668];
assign g[36053] = a[14] & g[19669];
assign g[52436] = b[14] & g[19669];
assign g[36054] = a[14] & g[19670];
assign g[52437] = b[14] & g[19670];
assign g[36055] = a[14] & g[19671];
assign g[52438] = b[14] & g[19671];
assign g[36056] = a[14] & g[19672];
assign g[52439] = b[14] & g[19672];
assign g[36057] = a[14] & g[19673];
assign g[52440] = b[14] & g[19673];
assign g[36058] = a[14] & g[19674];
assign g[52441] = b[14] & g[19674];
assign g[36059] = a[14] & g[19675];
assign g[52442] = b[14] & g[19675];
assign g[36060] = a[14] & g[19676];
assign g[52443] = b[14] & g[19676];
assign g[36061] = a[14] & g[19677];
assign g[52444] = b[14] & g[19677];
assign g[36062] = a[14] & g[19678];
assign g[52445] = b[14] & g[19678];
assign g[36063] = a[14] & g[19679];
assign g[52446] = b[14] & g[19679];
assign g[36064] = a[14] & g[19680];
assign g[52447] = b[14] & g[19680];
assign g[36065] = a[14] & g[19681];
assign g[52448] = b[14] & g[19681];
assign g[36066] = a[14] & g[19682];
assign g[52449] = b[14] & g[19682];
assign g[36067] = a[14] & g[19683];
assign g[52450] = b[14] & g[19683];
assign g[36068] = a[14] & g[19684];
assign g[52451] = b[14] & g[19684];
assign g[36069] = a[14] & g[19685];
assign g[52452] = b[14] & g[19685];
assign g[36070] = a[14] & g[19686];
assign g[52453] = b[14] & g[19686];
assign g[36071] = a[14] & g[19687];
assign g[52454] = b[14] & g[19687];
assign g[36072] = a[14] & g[19688];
assign g[52455] = b[14] & g[19688];
assign g[36073] = a[14] & g[19689];
assign g[52456] = b[14] & g[19689];
assign g[36074] = a[14] & g[19690];
assign g[52457] = b[14] & g[19690];
assign g[36075] = a[14] & g[19691];
assign g[52458] = b[14] & g[19691];
assign g[36076] = a[14] & g[19692];
assign g[52459] = b[14] & g[19692];
assign g[36077] = a[14] & g[19693];
assign g[52460] = b[14] & g[19693];
assign g[36078] = a[14] & g[19694];
assign g[52461] = b[14] & g[19694];
assign g[36079] = a[14] & g[19695];
assign g[52462] = b[14] & g[19695];
assign g[36080] = a[14] & g[19696];
assign g[52463] = b[14] & g[19696];
assign g[36081] = a[14] & g[19697];
assign g[52464] = b[14] & g[19697];
assign g[36082] = a[14] & g[19698];
assign g[52465] = b[14] & g[19698];
assign g[36083] = a[14] & g[19699];
assign g[52466] = b[14] & g[19699];
assign g[36084] = a[14] & g[19700];
assign g[52467] = b[14] & g[19700];
assign g[36085] = a[14] & g[19701];
assign g[52468] = b[14] & g[19701];
assign g[36086] = a[14] & g[19702];
assign g[52469] = b[14] & g[19702];
assign g[36087] = a[14] & g[19703];
assign g[52470] = b[14] & g[19703];
assign g[36088] = a[14] & g[19704];
assign g[52471] = b[14] & g[19704];
assign g[36089] = a[14] & g[19705];
assign g[52472] = b[14] & g[19705];
assign g[36090] = a[14] & g[19706];
assign g[52473] = b[14] & g[19706];
assign g[36091] = a[14] & g[19707];
assign g[52474] = b[14] & g[19707];
assign g[36092] = a[14] & g[19708];
assign g[52475] = b[14] & g[19708];
assign g[36093] = a[14] & g[19709];
assign g[52476] = b[14] & g[19709];
assign g[36094] = a[14] & g[19710];
assign g[52477] = b[14] & g[19710];
assign g[36095] = a[14] & g[19711];
assign g[52478] = b[14] & g[19711];
assign g[36096] = a[14] & g[19712];
assign g[52479] = b[14] & g[19712];
assign g[36097] = a[14] & g[19713];
assign g[52480] = b[14] & g[19713];
assign g[36098] = a[14] & g[19714];
assign g[52481] = b[14] & g[19714];
assign g[36099] = a[14] & g[19715];
assign g[52482] = b[14] & g[19715];
assign g[36100] = a[14] & g[19716];
assign g[52483] = b[14] & g[19716];
assign g[36101] = a[14] & g[19717];
assign g[52484] = b[14] & g[19717];
assign g[36102] = a[14] & g[19718];
assign g[52485] = b[14] & g[19718];
assign g[36103] = a[14] & g[19719];
assign g[52486] = b[14] & g[19719];
assign g[36104] = a[14] & g[19720];
assign g[52487] = b[14] & g[19720];
assign g[36105] = a[14] & g[19721];
assign g[52488] = b[14] & g[19721];
assign g[36106] = a[14] & g[19722];
assign g[52489] = b[14] & g[19722];
assign g[36107] = a[14] & g[19723];
assign g[52490] = b[14] & g[19723];
assign g[36108] = a[14] & g[19724];
assign g[52491] = b[14] & g[19724];
assign g[36109] = a[14] & g[19725];
assign g[52492] = b[14] & g[19725];
assign g[36110] = a[14] & g[19726];
assign g[52493] = b[14] & g[19726];
assign g[36111] = a[14] & g[19727];
assign g[52494] = b[14] & g[19727];
assign g[36112] = a[14] & g[19728];
assign g[52495] = b[14] & g[19728];
assign g[36113] = a[14] & g[19729];
assign g[52496] = b[14] & g[19729];
assign g[36114] = a[14] & g[19730];
assign g[52497] = b[14] & g[19730];
assign g[36115] = a[14] & g[19731];
assign g[52498] = b[14] & g[19731];
assign g[36116] = a[14] & g[19732];
assign g[52499] = b[14] & g[19732];
assign g[36117] = a[14] & g[19733];
assign g[52500] = b[14] & g[19733];
assign g[36118] = a[14] & g[19734];
assign g[52501] = b[14] & g[19734];
assign g[36119] = a[14] & g[19735];
assign g[52502] = b[14] & g[19735];
assign g[36120] = a[14] & g[19736];
assign g[52503] = b[14] & g[19736];
assign g[36121] = a[14] & g[19737];
assign g[52504] = b[14] & g[19737];
assign g[36122] = a[14] & g[19738];
assign g[52505] = b[14] & g[19738];
assign g[36123] = a[14] & g[19739];
assign g[52506] = b[14] & g[19739];
assign g[36124] = a[14] & g[19740];
assign g[52507] = b[14] & g[19740];
assign g[36125] = a[14] & g[19741];
assign g[52508] = b[14] & g[19741];
assign g[36126] = a[14] & g[19742];
assign g[52509] = b[14] & g[19742];
assign g[36127] = a[14] & g[19743];
assign g[52510] = b[14] & g[19743];
assign g[36128] = a[14] & g[19744];
assign g[52511] = b[14] & g[19744];
assign g[36129] = a[14] & g[19745];
assign g[52512] = b[14] & g[19745];
assign g[36130] = a[14] & g[19746];
assign g[52513] = b[14] & g[19746];
assign g[36131] = a[14] & g[19747];
assign g[52514] = b[14] & g[19747];
assign g[36132] = a[14] & g[19748];
assign g[52515] = b[14] & g[19748];
assign g[36133] = a[14] & g[19749];
assign g[52516] = b[14] & g[19749];
assign g[36134] = a[14] & g[19750];
assign g[52517] = b[14] & g[19750];
assign g[36135] = a[14] & g[19751];
assign g[52518] = b[14] & g[19751];
assign g[36136] = a[14] & g[19752];
assign g[52519] = b[14] & g[19752];
assign g[36137] = a[14] & g[19753];
assign g[52520] = b[14] & g[19753];
assign g[36138] = a[14] & g[19754];
assign g[52521] = b[14] & g[19754];
assign g[36139] = a[14] & g[19755];
assign g[52522] = b[14] & g[19755];
assign g[36140] = a[14] & g[19756];
assign g[52523] = b[14] & g[19756];
assign g[36141] = a[14] & g[19757];
assign g[52524] = b[14] & g[19757];
assign g[36142] = a[14] & g[19758];
assign g[52525] = b[14] & g[19758];
assign g[36143] = a[14] & g[19759];
assign g[52526] = b[14] & g[19759];
assign g[36144] = a[14] & g[19760];
assign g[52527] = b[14] & g[19760];
assign g[36145] = a[14] & g[19761];
assign g[52528] = b[14] & g[19761];
assign g[36146] = a[14] & g[19762];
assign g[52529] = b[14] & g[19762];
assign g[36147] = a[14] & g[19763];
assign g[52530] = b[14] & g[19763];
assign g[36148] = a[14] & g[19764];
assign g[52531] = b[14] & g[19764];
assign g[36149] = a[14] & g[19765];
assign g[52532] = b[14] & g[19765];
assign g[36150] = a[14] & g[19766];
assign g[52533] = b[14] & g[19766];
assign g[36151] = a[14] & g[19767];
assign g[52534] = b[14] & g[19767];
assign g[36152] = a[14] & g[19768];
assign g[52535] = b[14] & g[19768];
assign g[36153] = a[14] & g[19769];
assign g[52536] = b[14] & g[19769];
assign g[36154] = a[14] & g[19770];
assign g[52537] = b[14] & g[19770];
assign g[36155] = a[14] & g[19771];
assign g[52538] = b[14] & g[19771];
assign g[36156] = a[14] & g[19772];
assign g[52539] = b[14] & g[19772];
assign g[36157] = a[14] & g[19773];
assign g[52540] = b[14] & g[19773];
assign g[36158] = a[14] & g[19774];
assign g[52541] = b[14] & g[19774];
assign g[36159] = a[14] & g[19775];
assign g[52542] = b[14] & g[19775];
assign g[36160] = a[14] & g[19776];
assign g[52543] = b[14] & g[19776];
assign g[36161] = a[14] & g[19777];
assign g[52544] = b[14] & g[19777];
assign g[36162] = a[14] & g[19778];
assign g[52545] = b[14] & g[19778];
assign g[36163] = a[14] & g[19779];
assign g[52546] = b[14] & g[19779];
assign g[36164] = a[14] & g[19780];
assign g[52547] = b[14] & g[19780];
assign g[36165] = a[14] & g[19781];
assign g[52548] = b[14] & g[19781];
assign g[36166] = a[14] & g[19782];
assign g[52549] = b[14] & g[19782];
assign g[36167] = a[14] & g[19783];
assign g[52550] = b[14] & g[19783];
assign g[36168] = a[14] & g[19784];
assign g[52551] = b[14] & g[19784];
assign g[36169] = a[14] & g[19785];
assign g[52552] = b[14] & g[19785];
assign g[36170] = a[14] & g[19786];
assign g[52553] = b[14] & g[19786];
assign g[36171] = a[14] & g[19787];
assign g[52554] = b[14] & g[19787];
assign g[36172] = a[14] & g[19788];
assign g[52555] = b[14] & g[19788];
assign g[36173] = a[14] & g[19789];
assign g[52556] = b[14] & g[19789];
assign g[36174] = a[14] & g[19790];
assign g[52557] = b[14] & g[19790];
assign g[36175] = a[14] & g[19791];
assign g[52558] = b[14] & g[19791];
assign g[36176] = a[14] & g[19792];
assign g[52559] = b[14] & g[19792];
assign g[36177] = a[14] & g[19793];
assign g[52560] = b[14] & g[19793];
assign g[36178] = a[14] & g[19794];
assign g[52561] = b[14] & g[19794];
assign g[36179] = a[14] & g[19795];
assign g[52562] = b[14] & g[19795];
assign g[36180] = a[14] & g[19796];
assign g[52563] = b[14] & g[19796];
assign g[36181] = a[14] & g[19797];
assign g[52564] = b[14] & g[19797];
assign g[36182] = a[14] & g[19798];
assign g[52565] = b[14] & g[19798];
assign g[36183] = a[14] & g[19799];
assign g[52566] = b[14] & g[19799];
assign g[36184] = a[14] & g[19800];
assign g[52567] = b[14] & g[19800];
assign g[36185] = a[14] & g[19801];
assign g[52568] = b[14] & g[19801];
assign g[36186] = a[14] & g[19802];
assign g[52569] = b[14] & g[19802];
assign g[36187] = a[14] & g[19803];
assign g[52570] = b[14] & g[19803];
assign g[36188] = a[14] & g[19804];
assign g[52571] = b[14] & g[19804];
assign g[36189] = a[14] & g[19805];
assign g[52572] = b[14] & g[19805];
assign g[36190] = a[14] & g[19806];
assign g[52573] = b[14] & g[19806];
assign g[36191] = a[14] & g[19807];
assign g[52574] = b[14] & g[19807];
assign g[36192] = a[14] & g[19808];
assign g[52575] = b[14] & g[19808];
assign g[36193] = a[14] & g[19809];
assign g[52576] = b[14] & g[19809];
assign g[36194] = a[14] & g[19810];
assign g[52577] = b[14] & g[19810];
assign g[36195] = a[14] & g[19811];
assign g[52578] = b[14] & g[19811];
assign g[36196] = a[14] & g[19812];
assign g[52579] = b[14] & g[19812];
assign g[36197] = a[14] & g[19813];
assign g[52580] = b[14] & g[19813];
assign g[36198] = a[14] & g[19814];
assign g[52581] = b[14] & g[19814];
assign g[36199] = a[14] & g[19815];
assign g[52582] = b[14] & g[19815];
assign g[36200] = a[14] & g[19816];
assign g[52583] = b[14] & g[19816];
assign g[36201] = a[14] & g[19817];
assign g[52584] = b[14] & g[19817];
assign g[36202] = a[14] & g[19818];
assign g[52585] = b[14] & g[19818];
assign g[36203] = a[14] & g[19819];
assign g[52586] = b[14] & g[19819];
assign g[36204] = a[14] & g[19820];
assign g[52587] = b[14] & g[19820];
assign g[36205] = a[14] & g[19821];
assign g[52588] = b[14] & g[19821];
assign g[36206] = a[14] & g[19822];
assign g[52589] = b[14] & g[19822];
assign g[36207] = a[14] & g[19823];
assign g[52590] = b[14] & g[19823];
assign g[36208] = a[14] & g[19824];
assign g[52591] = b[14] & g[19824];
assign g[36209] = a[14] & g[19825];
assign g[52592] = b[14] & g[19825];
assign g[36210] = a[14] & g[19826];
assign g[52593] = b[14] & g[19826];
assign g[36211] = a[14] & g[19827];
assign g[52594] = b[14] & g[19827];
assign g[36212] = a[14] & g[19828];
assign g[52595] = b[14] & g[19828];
assign g[36213] = a[14] & g[19829];
assign g[52596] = b[14] & g[19829];
assign g[36214] = a[14] & g[19830];
assign g[52597] = b[14] & g[19830];
assign g[36215] = a[14] & g[19831];
assign g[52598] = b[14] & g[19831];
assign g[36216] = a[14] & g[19832];
assign g[52599] = b[14] & g[19832];
assign g[36217] = a[14] & g[19833];
assign g[52600] = b[14] & g[19833];
assign g[36218] = a[14] & g[19834];
assign g[52601] = b[14] & g[19834];
assign g[36219] = a[14] & g[19835];
assign g[52602] = b[14] & g[19835];
assign g[36220] = a[14] & g[19836];
assign g[52603] = b[14] & g[19836];
assign g[36221] = a[14] & g[19837];
assign g[52604] = b[14] & g[19837];
assign g[36222] = a[14] & g[19838];
assign g[52605] = b[14] & g[19838];
assign g[36223] = a[14] & g[19839];
assign g[52606] = b[14] & g[19839];
assign g[36224] = a[14] & g[19840];
assign g[52607] = b[14] & g[19840];
assign g[36225] = a[14] & g[19841];
assign g[52608] = b[14] & g[19841];
assign g[36226] = a[14] & g[19842];
assign g[52609] = b[14] & g[19842];
assign g[36227] = a[14] & g[19843];
assign g[52610] = b[14] & g[19843];
assign g[36228] = a[14] & g[19844];
assign g[52611] = b[14] & g[19844];
assign g[36229] = a[14] & g[19845];
assign g[52612] = b[14] & g[19845];
assign g[36230] = a[14] & g[19846];
assign g[52613] = b[14] & g[19846];
assign g[36231] = a[14] & g[19847];
assign g[52614] = b[14] & g[19847];
assign g[36232] = a[14] & g[19848];
assign g[52615] = b[14] & g[19848];
assign g[36233] = a[14] & g[19849];
assign g[52616] = b[14] & g[19849];
assign g[36234] = a[14] & g[19850];
assign g[52617] = b[14] & g[19850];
assign g[36235] = a[14] & g[19851];
assign g[52618] = b[14] & g[19851];
assign g[36236] = a[14] & g[19852];
assign g[52619] = b[14] & g[19852];
assign g[36237] = a[14] & g[19853];
assign g[52620] = b[14] & g[19853];
assign g[36238] = a[14] & g[19854];
assign g[52621] = b[14] & g[19854];
assign g[36239] = a[14] & g[19855];
assign g[52622] = b[14] & g[19855];
assign g[36240] = a[14] & g[19856];
assign g[52623] = b[14] & g[19856];
assign g[36241] = a[14] & g[19857];
assign g[52624] = b[14] & g[19857];
assign g[36242] = a[14] & g[19858];
assign g[52625] = b[14] & g[19858];
assign g[36243] = a[14] & g[19859];
assign g[52626] = b[14] & g[19859];
assign g[36244] = a[14] & g[19860];
assign g[52627] = b[14] & g[19860];
assign g[36245] = a[14] & g[19861];
assign g[52628] = b[14] & g[19861];
assign g[36246] = a[14] & g[19862];
assign g[52629] = b[14] & g[19862];
assign g[36247] = a[14] & g[19863];
assign g[52630] = b[14] & g[19863];
assign g[36248] = a[14] & g[19864];
assign g[52631] = b[14] & g[19864];
assign g[36249] = a[14] & g[19865];
assign g[52632] = b[14] & g[19865];
assign g[36250] = a[14] & g[19866];
assign g[52633] = b[14] & g[19866];
assign g[36251] = a[14] & g[19867];
assign g[52634] = b[14] & g[19867];
assign g[36252] = a[14] & g[19868];
assign g[52635] = b[14] & g[19868];
assign g[36253] = a[14] & g[19869];
assign g[52636] = b[14] & g[19869];
assign g[36254] = a[14] & g[19870];
assign g[52637] = b[14] & g[19870];
assign g[36255] = a[14] & g[19871];
assign g[52638] = b[14] & g[19871];
assign g[36256] = a[14] & g[19872];
assign g[52639] = b[14] & g[19872];
assign g[36257] = a[14] & g[19873];
assign g[52640] = b[14] & g[19873];
assign g[36258] = a[14] & g[19874];
assign g[52641] = b[14] & g[19874];
assign g[36259] = a[14] & g[19875];
assign g[52642] = b[14] & g[19875];
assign g[36260] = a[14] & g[19876];
assign g[52643] = b[14] & g[19876];
assign g[36261] = a[14] & g[19877];
assign g[52644] = b[14] & g[19877];
assign g[36262] = a[14] & g[19878];
assign g[52645] = b[14] & g[19878];
assign g[36263] = a[14] & g[19879];
assign g[52646] = b[14] & g[19879];
assign g[36264] = a[14] & g[19880];
assign g[52647] = b[14] & g[19880];
assign g[36265] = a[14] & g[19881];
assign g[52648] = b[14] & g[19881];
assign g[36266] = a[14] & g[19882];
assign g[52649] = b[14] & g[19882];
assign g[36267] = a[14] & g[19883];
assign g[52650] = b[14] & g[19883];
assign g[36268] = a[14] & g[19884];
assign g[52651] = b[14] & g[19884];
assign g[36269] = a[14] & g[19885];
assign g[52652] = b[14] & g[19885];
assign g[36270] = a[14] & g[19886];
assign g[52653] = b[14] & g[19886];
assign g[36271] = a[14] & g[19887];
assign g[52654] = b[14] & g[19887];
assign g[36272] = a[14] & g[19888];
assign g[52655] = b[14] & g[19888];
assign g[36273] = a[14] & g[19889];
assign g[52656] = b[14] & g[19889];
assign g[36274] = a[14] & g[19890];
assign g[52657] = b[14] & g[19890];
assign g[36275] = a[14] & g[19891];
assign g[52658] = b[14] & g[19891];
assign g[36276] = a[14] & g[19892];
assign g[52659] = b[14] & g[19892];
assign g[36277] = a[14] & g[19893];
assign g[52660] = b[14] & g[19893];
assign g[36278] = a[14] & g[19894];
assign g[52661] = b[14] & g[19894];
assign g[36279] = a[14] & g[19895];
assign g[52662] = b[14] & g[19895];
assign g[36280] = a[14] & g[19896];
assign g[52663] = b[14] & g[19896];
assign g[36281] = a[14] & g[19897];
assign g[52664] = b[14] & g[19897];
assign g[36282] = a[14] & g[19898];
assign g[52665] = b[14] & g[19898];
assign g[36283] = a[14] & g[19899];
assign g[52666] = b[14] & g[19899];
assign g[36284] = a[14] & g[19900];
assign g[52667] = b[14] & g[19900];
assign g[36285] = a[14] & g[19901];
assign g[52668] = b[14] & g[19901];
assign g[36286] = a[14] & g[19902];
assign g[52669] = b[14] & g[19902];
assign g[36287] = a[14] & g[19903];
assign g[52670] = b[14] & g[19903];
assign g[36288] = a[14] & g[19904];
assign g[52671] = b[14] & g[19904];
assign g[36289] = a[14] & g[19905];
assign g[52672] = b[14] & g[19905];
assign g[36290] = a[14] & g[19906];
assign g[52673] = b[14] & g[19906];
assign g[36291] = a[14] & g[19907];
assign g[52674] = b[14] & g[19907];
assign g[36292] = a[14] & g[19908];
assign g[52675] = b[14] & g[19908];
assign g[36293] = a[14] & g[19909];
assign g[52676] = b[14] & g[19909];
assign g[36294] = a[14] & g[19910];
assign g[52677] = b[14] & g[19910];
assign g[36295] = a[14] & g[19911];
assign g[52678] = b[14] & g[19911];
assign g[36296] = a[14] & g[19912];
assign g[52679] = b[14] & g[19912];
assign g[36297] = a[14] & g[19913];
assign g[52680] = b[14] & g[19913];
assign g[36298] = a[14] & g[19914];
assign g[52681] = b[14] & g[19914];
assign g[36299] = a[14] & g[19915];
assign g[52682] = b[14] & g[19915];
assign g[36300] = a[14] & g[19916];
assign g[52683] = b[14] & g[19916];
assign g[36301] = a[14] & g[19917];
assign g[52684] = b[14] & g[19917];
assign g[36302] = a[14] & g[19918];
assign g[52685] = b[14] & g[19918];
assign g[36303] = a[14] & g[19919];
assign g[52686] = b[14] & g[19919];
assign g[36304] = a[14] & g[19920];
assign g[52687] = b[14] & g[19920];
assign g[36305] = a[14] & g[19921];
assign g[52688] = b[14] & g[19921];
assign g[36306] = a[14] & g[19922];
assign g[52689] = b[14] & g[19922];
assign g[36307] = a[14] & g[19923];
assign g[52690] = b[14] & g[19923];
assign g[36308] = a[14] & g[19924];
assign g[52691] = b[14] & g[19924];
assign g[36309] = a[14] & g[19925];
assign g[52692] = b[14] & g[19925];
assign g[36310] = a[14] & g[19926];
assign g[52693] = b[14] & g[19926];
assign g[36311] = a[14] & g[19927];
assign g[52694] = b[14] & g[19927];
assign g[36312] = a[14] & g[19928];
assign g[52695] = b[14] & g[19928];
assign g[36313] = a[14] & g[19929];
assign g[52696] = b[14] & g[19929];
assign g[36314] = a[14] & g[19930];
assign g[52697] = b[14] & g[19930];
assign g[36315] = a[14] & g[19931];
assign g[52698] = b[14] & g[19931];
assign g[36316] = a[14] & g[19932];
assign g[52699] = b[14] & g[19932];
assign g[36317] = a[14] & g[19933];
assign g[52700] = b[14] & g[19933];
assign g[36318] = a[14] & g[19934];
assign g[52701] = b[14] & g[19934];
assign g[36319] = a[14] & g[19935];
assign g[52702] = b[14] & g[19935];
assign g[36320] = a[14] & g[19936];
assign g[52703] = b[14] & g[19936];
assign g[36321] = a[14] & g[19937];
assign g[52704] = b[14] & g[19937];
assign g[36322] = a[14] & g[19938];
assign g[52705] = b[14] & g[19938];
assign g[36323] = a[14] & g[19939];
assign g[52706] = b[14] & g[19939];
assign g[36324] = a[14] & g[19940];
assign g[52707] = b[14] & g[19940];
assign g[36325] = a[14] & g[19941];
assign g[52708] = b[14] & g[19941];
assign g[36326] = a[14] & g[19942];
assign g[52709] = b[14] & g[19942];
assign g[36327] = a[14] & g[19943];
assign g[52710] = b[14] & g[19943];
assign g[36328] = a[14] & g[19944];
assign g[52711] = b[14] & g[19944];
assign g[36329] = a[14] & g[19945];
assign g[52712] = b[14] & g[19945];
assign g[36330] = a[14] & g[19946];
assign g[52713] = b[14] & g[19946];
assign g[36331] = a[14] & g[19947];
assign g[52714] = b[14] & g[19947];
assign g[36332] = a[14] & g[19948];
assign g[52715] = b[14] & g[19948];
assign g[36333] = a[14] & g[19949];
assign g[52716] = b[14] & g[19949];
assign g[36334] = a[14] & g[19950];
assign g[52717] = b[14] & g[19950];
assign g[36335] = a[14] & g[19951];
assign g[52718] = b[14] & g[19951];
assign g[36336] = a[14] & g[19952];
assign g[52719] = b[14] & g[19952];
assign g[36337] = a[14] & g[19953];
assign g[52720] = b[14] & g[19953];
assign g[36338] = a[14] & g[19954];
assign g[52721] = b[14] & g[19954];
assign g[36339] = a[14] & g[19955];
assign g[52722] = b[14] & g[19955];
assign g[36340] = a[14] & g[19956];
assign g[52723] = b[14] & g[19956];
assign g[36341] = a[14] & g[19957];
assign g[52724] = b[14] & g[19957];
assign g[36342] = a[14] & g[19958];
assign g[52725] = b[14] & g[19958];
assign g[36343] = a[14] & g[19959];
assign g[52726] = b[14] & g[19959];
assign g[36344] = a[14] & g[19960];
assign g[52727] = b[14] & g[19960];
assign g[36345] = a[14] & g[19961];
assign g[52728] = b[14] & g[19961];
assign g[36346] = a[14] & g[19962];
assign g[52729] = b[14] & g[19962];
assign g[36347] = a[14] & g[19963];
assign g[52730] = b[14] & g[19963];
assign g[36348] = a[14] & g[19964];
assign g[52731] = b[14] & g[19964];
assign g[36349] = a[14] & g[19965];
assign g[52732] = b[14] & g[19965];
assign g[36350] = a[14] & g[19966];
assign g[52733] = b[14] & g[19966];
assign g[36351] = a[14] & g[19967];
assign g[52734] = b[14] & g[19967];
assign g[36352] = a[14] & g[19968];
assign g[52735] = b[14] & g[19968];
assign g[36353] = a[14] & g[19969];
assign g[52736] = b[14] & g[19969];
assign g[36354] = a[14] & g[19970];
assign g[52737] = b[14] & g[19970];
assign g[36355] = a[14] & g[19971];
assign g[52738] = b[14] & g[19971];
assign g[36356] = a[14] & g[19972];
assign g[52739] = b[14] & g[19972];
assign g[36357] = a[14] & g[19973];
assign g[52740] = b[14] & g[19973];
assign g[36358] = a[14] & g[19974];
assign g[52741] = b[14] & g[19974];
assign g[36359] = a[14] & g[19975];
assign g[52742] = b[14] & g[19975];
assign g[36360] = a[14] & g[19976];
assign g[52743] = b[14] & g[19976];
assign g[36361] = a[14] & g[19977];
assign g[52744] = b[14] & g[19977];
assign g[36362] = a[14] & g[19978];
assign g[52745] = b[14] & g[19978];
assign g[36363] = a[14] & g[19979];
assign g[52746] = b[14] & g[19979];
assign g[36364] = a[14] & g[19980];
assign g[52747] = b[14] & g[19980];
assign g[36365] = a[14] & g[19981];
assign g[52748] = b[14] & g[19981];
assign g[36366] = a[14] & g[19982];
assign g[52749] = b[14] & g[19982];
assign g[36367] = a[14] & g[19983];
assign g[52750] = b[14] & g[19983];
assign g[36368] = a[14] & g[19984];
assign g[52751] = b[14] & g[19984];
assign g[36369] = a[14] & g[19985];
assign g[52752] = b[14] & g[19985];
assign g[36370] = a[14] & g[19986];
assign g[52753] = b[14] & g[19986];
assign g[36371] = a[14] & g[19987];
assign g[52754] = b[14] & g[19987];
assign g[36372] = a[14] & g[19988];
assign g[52755] = b[14] & g[19988];
assign g[36373] = a[14] & g[19989];
assign g[52756] = b[14] & g[19989];
assign g[36374] = a[14] & g[19990];
assign g[52757] = b[14] & g[19990];
assign g[36375] = a[14] & g[19991];
assign g[52758] = b[14] & g[19991];
assign g[36376] = a[14] & g[19992];
assign g[52759] = b[14] & g[19992];
assign g[36377] = a[14] & g[19993];
assign g[52760] = b[14] & g[19993];
assign g[36378] = a[14] & g[19994];
assign g[52761] = b[14] & g[19994];
assign g[36379] = a[14] & g[19995];
assign g[52762] = b[14] & g[19995];
assign g[36380] = a[14] & g[19996];
assign g[52763] = b[14] & g[19996];
assign g[36381] = a[14] & g[19997];
assign g[52764] = b[14] & g[19997];
assign g[36382] = a[14] & g[19998];
assign g[52765] = b[14] & g[19998];
assign g[36383] = a[14] & g[19999];
assign g[52766] = b[14] & g[19999];
assign g[36384] = a[14] & g[20000];
assign g[52767] = b[14] & g[20000];
assign g[36385] = a[14] & g[20001];
assign g[52768] = b[14] & g[20001];
assign g[36386] = a[14] & g[20002];
assign g[52769] = b[14] & g[20002];
assign g[36387] = a[14] & g[20003];
assign g[52770] = b[14] & g[20003];
assign g[36388] = a[14] & g[20004];
assign g[52771] = b[14] & g[20004];
assign g[36389] = a[14] & g[20005];
assign g[52772] = b[14] & g[20005];
assign g[36390] = a[14] & g[20006];
assign g[52773] = b[14] & g[20006];
assign g[36391] = a[14] & g[20007];
assign g[52774] = b[14] & g[20007];
assign g[36392] = a[14] & g[20008];
assign g[52775] = b[14] & g[20008];
assign g[36393] = a[14] & g[20009];
assign g[52776] = b[14] & g[20009];
assign g[36394] = a[14] & g[20010];
assign g[52777] = b[14] & g[20010];
assign g[36395] = a[14] & g[20011];
assign g[52778] = b[14] & g[20011];
assign g[36396] = a[14] & g[20012];
assign g[52779] = b[14] & g[20012];
assign g[36397] = a[14] & g[20013];
assign g[52780] = b[14] & g[20013];
assign g[36398] = a[14] & g[20014];
assign g[52781] = b[14] & g[20014];
assign g[36399] = a[14] & g[20015];
assign g[52782] = b[14] & g[20015];
assign g[36400] = a[14] & g[20016];
assign g[52783] = b[14] & g[20016];
assign g[36401] = a[14] & g[20017];
assign g[52784] = b[14] & g[20017];
assign g[36402] = a[14] & g[20018];
assign g[52785] = b[14] & g[20018];
assign g[36403] = a[14] & g[20019];
assign g[52786] = b[14] & g[20019];
assign g[36404] = a[14] & g[20020];
assign g[52787] = b[14] & g[20020];
assign g[36405] = a[14] & g[20021];
assign g[52788] = b[14] & g[20021];
assign g[36406] = a[14] & g[20022];
assign g[52789] = b[14] & g[20022];
assign g[36407] = a[14] & g[20023];
assign g[52790] = b[14] & g[20023];
assign g[36408] = a[14] & g[20024];
assign g[52791] = b[14] & g[20024];
assign g[36409] = a[14] & g[20025];
assign g[52792] = b[14] & g[20025];
assign g[36410] = a[14] & g[20026];
assign g[52793] = b[14] & g[20026];
assign g[36411] = a[14] & g[20027];
assign g[52794] = b[14] & g[20027];
assign g[36412] = a[14] & g[20028];
assign g[52795] = b[14] & g[20028];
assign g[36413] = a[14] & g[20029];
assign g[52796] = b[14] & g[20029];
assign g[36414] = a[14] & g[20030];
assign g[52797] = b[14] & g[20030];
assign g[36415] = a[14] & g[20031];
assign g[52798] = b[14] & g[20031];
assign g[36416] = a[14] & g[20032];
assign g[52799] = b[14] & g[20032];
assign g[36417] = a[14] & g[20033];
assign g[52800] = b[14] & g[20033];
assign g[36418] = a[14] & g[20034];
assign g[52801] = b[14] & g[20034];
assign g[36419] = a[14] & g[20035];
assign g[52802] = b[14] & g[20035];
assign g[36420] = a[14] & g[20036];
assign g[52803] = b[14] & g[20036];
assign g[36421] = a[14] & g[20037];
assign g[52804] = b[14] & g[20037];
assign g[36422] = a[14] & g[20038];
assign g[52805] = b[14] & g[20038];
assign g[36423] = a[14] & g[20039];
assign g[52806] = b[14] & g[20039];
assign g[36424] = a[14] & g[20040];
assign g[52807] = b[14] & g[20040];
assign g[36425] = a[14] & g[20041];
assign g[52808] = b[14] & g[20041];
assign g[36426] = a[14] & g[20042];
assign g[52809] = b[14] & g[20042];
assign g[36427] = a[14] & g[20043];
assign g[52810] = b[14] & g[20043];
assign g[36428] = a[14] & g[20044];
assign g[52811] = b[14] & g[20044];
assign g[36429] = a[14] & g[20045];
assign g[52812] = b[14] & g[20045];
assign g[36430] = a[14] & g[20046];
assign g[52813] = b[14] & g[20046];
assign g[36431] = a[14] & g[20047];
assign g[52814] = b[14] & g[20047];
assign g[36432] = a[14] & g[20048];
assign g[52815] = b[14] & g[20048];
assign g[36433] = a[14] & g[20049];
assign g[52816] = b[14] & g[20049];
assign g[36434] = a[14] & g[20050];
assign g[52817] = b[14] & g[20050];
assign g[36435] = a[14] & g[20051];
assign g[52818] = b[14] & g[20051];
assign g[36436] = a[14] & g[20052];
assign g[52819] = b[14] & g[20052];
assign g[36437] = a[14] & g[20053];
assign g[52820] = b[14] & g[20053];
assign g[36438] = a[14] & g[20054];
assign g[52821] = b[14] & g[20054];
assign g[36439] = a[14] & g[20055];
assign g[52822] = b[14] & g[20055];
assign g[36440] = a[14] & g[20056];
assign g[52823] = b[14] & g[20056];
assign g[36441] = a[14] & g[20057];
assign g[52824] = b[14] & g[20057];
assign g[36442] = a[14] & g[20058];
assign g[52825] = b[14] & g[20058];
assign g[36443] = a[14] & g[20059];
assign g[52826] = b[14] & g[20059];
assign g[36444] = a[14] & g[20060];
assign g[52827] = b[14] & g[20060];
assign g[36445] = a[14] & g[20061];
assign g[52828] = b[14] & g[20061];
assign g[36446] = a[14] & g[20062];
assign g[52829] = b[14] & g[20062];
assign g[36447] = a[14] & g[20063];
assign g[52830] = b[14] & g[20063];
assign g[36448] = a[14] & g[20064];
assign g[52831] = b[14] & g[20064];
assign g[36449] = a[14] & g[20065];
assign g[52832] = b[14] & g[20065];
assign g[36450] = a[14] & g[20066];
assign g[52833] = b[14] & g[20066];
assign g[36451] = a[14] & g[20067];
assign g[52834] = b[14] & g[20067];
assign g[36452] = a[14] & g[20068];
assign g[52835] = b[14] & g[20068];
assign g[36453] = a[14] & g[20069];
assign g[52836] = b[14] & g[20069];
assign g[36454] = a[14] & g[20070];
assign g[52837] = b[14] & g[20070];
assign g[36455] = a[14] & g[20071];
assign g[52838] = b[14] & g[20071];
assign g[36456] = a[14] & g[20072];
assign g[52839] = b[14] & g[20072];
assign g[36457] = a[14] & g[20073];
assign g[52840] = b[14] & g[20073];
assign g[36458] = a[14] & g[20074];
assign g[52841] = b[14] & g[20074];
assign g[36459] = a[14] & g[20075];
assign g[52842] = b[14] & g[20075];
assign g[36460] = a[14] & g[20076];
assign g[52843] = b[14] & g[20076];
assign g[36461] = a[14] & g[20077];
assign g[52844] = b[14] & g[20077];
assign g[36462] = a[14] & g[20078];
assign g[52845] = b[14] & g[20078];
assign g[36463] = a[14] & g[20079];
assign g[52846] = b[14] & g[20079];
assign g[36464] = a[14] & g[20080];
assign g[52847] = b[14] & g[20080];
assign g[36465] = a[14] & g[20081];
assign g[52848] = b[14] & g[20081];
assign g[36466] = a[14] & g[20082];
assign g[52849] = b[14] & g[20082];
assign g[36467] = a[14] & g[20083];
assign g[52850] = b[14] & g[20083];
assign g[36468] = a[14] & g[20084];
assign g[52851] = b[14] & g[20084];
assign g[36469] = a[14] & g[20085];
assign g[52852] = b[14] & g[20085];
assign g[36470] = a[14] & g[20086];
assign g[52853] = b[14] & g[20086];
assign g[36471] = a[14] & g[20087];
assign g[52854] = b[14] & g[20087];
assign g[36472] = a[14] & g[20088];
assign g[52855] = b[14] & g[20088];
assign g[36473] = a[14] & g[20089];
assign g[52856] = b[14] & g[20089];
assign g[36474] = a[14] & g[20090];
assign g[52857] = b[14] & g[20090];
assign g[36475] = a[14] & g[20091];
assign g[52858] = b[14] & g[20091];
assign g[36476] = a[14] & g[20092];
assign g[52859] = b[14] & g[20092];
assign g[36477] = a[14] & g[20093];
assign g[52860] = b[14] & g[20093];
assign g[36478] = a[14] & g[20094];
assign g[52861] = b[14] & g[20094];
assign g[36479] = a[14] & g[20095];
assign g[52862] = b[14] & g[20095];
assign g[36480] = a[14] & g[20096];
assign g[52863] = b[14] & g[20096];
assign g[36481] = a[14] & g[20097];
assign g[52864] = b[14] & g[20097];
assign g[36482] = a[14] & g[20098];
assign g[52865] = b[14] & g[20098];
assign g[36483] = a[14] & g[20099];
assign g[52866] = b[14] & g[20099];
assign g[36484] = a[14] & g[20100];
assign g[52867] = b[14] & g[20100];
assign g[36485] = a[14] & g[20101];
assign g[52868] = b[14] & g[20101];
assign g[36486] = a[14] & g[20102];
assign g[52869] = b[14] & g[20102];
assign g[36487] = a[14] & g[20103];
assign g[52870] = b[14] & g[20103];
assign g[36488] = a[14] & g[20104];
assign g[52871] = b[14] & g[20104];
assign g[36489] = a[14] & g[20105];
assign g[52872] = b[14] & g[20105];
assign g[36490] = a[14] & g[20106];
assign g[52873] = b[14] & g[20106];
assign g[36491] = a[14] & g[20107];
assign g[52874] = b[14] & g[20107];
assign g[36492] = a[14] & g[20108];
assign g[52875] = b[14] & g[20108];
assign g[36493] = a[14] & g[20109];
assign g[52876] = b[14] & g[20109];
assign g[36494] = a[14] & g[20110];
assign g[52877] = b[14] & g[20110];
assign g[36495] = a[14] & g[20111];
assign g[52878] = b[14] & g[20111];
assign g[36496] = a[14] & g[20112];
assign g[52879] = b[14] & g[20112];
assign g[36497] = a[14] & g[20113];
assign g[52880] = b[14] & g[20113];
assign g[36498] = a[14] & g[20114];
assign g[52881] = b[14] & g[20114];
assign g[36499] = a[14] & g[20115];
assign g[52882] = b[14] & g[20115];
assign g[36500] = a[14] & g[20116];
assign g[52883] = b[14] & g[20116];
assign g[36501] = a[14] & g[20117];
assign g[52884] = b[14] & g[20117];
assign g[36502] = a[14] & g[20118];
assign g[52885] = b[14] & g[20118];
assign g[36503] = a[14] & g[20119];
assign g[52886] = b[14] & g[20119];
assign g[36504] = a[14] & g[20120];
assign g[52887] = b[14] & g[20120];
assign g[36505] = a[14] & g[20121];
assign g[52888] = b[14] & g[20121];
assign g[36506] = a[14] & g[20122];
assign g[52889] = b[14] & g[20122];
assign g[36507] = a[14] & g[20123];
assign g[52890] = b[14] & g[20123];
assign g[36508] = a[14] & g[20124];
assign g[52891] = b[14] & g[20124];
assign g[36509] = a[14] & g[20125];
assign g[52892] = b[14] & g[20125];
assign g[36510] = a[14] & g[20126];
assign g[52893] = b[14] & g[20126];
assign g[36511] = a[14] & g[20127];
assign g[52894] = b[14] & g[20127];
assign g[36512] = a[14] & g[20128];
assign g[52895] = b[14] & g[20128];
assign g[36513] = a[14] & g[20129];
assign g[52896] = b[14] & g[20129];
assign g[36514] = a[14] & g[20130];
assign g[52897] = b[14] & g[20130];
assign g[36515] = a[14] & g[20131];
assign g[52898] = b[14] & g[20131];
assign g[36516] = a[14] & g[20132];
assign g[52899] = b[14] & g[20132];
assign g[36517] = a[14] & g[20133];
assign g[52900] = b[14] & g[20133];
assign g[36518] = a[14] & g[20134];
assign g[52901] = b[14] & g[20134];
assign g[36519] = a[14] & g[20135];
assign g[52902] = b[14] & g[20135];
assign g[36520] = a[14] & g[20136];
assign g[52903] = b[14] & g[20136];
assign g[36521] = a[14] & g[20137];
assign g[52904] = b[14] & g[20137];
assign g[36522] = a[14] & g[20138];
assign g[52905] = b[14] & g[20138];
assign g[36523] = a[14] & g[20139];
assign g[52906] = b[14] & g[20139];
assign g[36524] = a[14] & g[20140];
assign g[52907] = b[14] & g[20140];
assign g[36525] = a[14] & g[20141];
assign g[52908] = b[14] & g[20141];
assign g[36526] = a[14] & g[20142];
assign g[52909] = b[14] & g[20142];
assign g[36527] = a[14] & g[20143];
assign g[52910] = b[14] & g[20143];
assign g[36528] = a[14] & g[20144];
assign g[52911] = b[14] & g[20144];
assign g[36529] = a[14] & g[20145];
assign g[52912] = b[14] & g[20145];
assign g[36530] = a[14] & g[20146];
assign g[52913] = b[14] & g[20146];
assign g[36531] = a[14] & g[20147];
assign g[52914] = b[14] & g[20147];
assign g[36532] = a[14] & g[20148];
assign g[52915] = b[14] & g[20148];
assign g[36533] = a[14] & g[20149];
assign g[52916] = b[14] & g[20149];
assign g[36534] = a[14] & g[20150];
assign g[52917] = b[14] & g[20150];
assign g[36535] = a[14] & g[20151];
assign g[52918] = b[14] & g[20151];
assign g[36536] = a[14] & g[20152];
assign g[52919] = b[14] & g[20152];
assign g[36537] = a[14] & g[20153];
assign g[52920] = b[14] & g[20153];
assign g[36538] = a[14] & g[20154];
assign g[52921] = b[14] & g[20154];
assign g[36539] = a[14] & g[20155];
assign g[52922] = b[14] & g[20155];
assign g[36540] = a[14] & g[20156];
assign g[52923] = b[14] & g[20156];
assign g[36541] = a[14] & g[20157];
assign g[52924] = b[14] & g[20157];
assign g[36542] = a[14] & g[20158];
assign g[52925] = b[14] & g[20158];
assign g[36543] = a[14] & g[20159];
assign g[52926] = b[14] & g[20159];
assign g[36544] = a[14] & g[20160];
assign g[52927] = b[14] & g[20160];
assign g[36545] = a[14] & g[20161];
assign g[52928] = b[14] & g[20161];
assign g[36546] = a[14] & g[20162];
assign g[52929] = b[14] & g[20162];
assign g[36547] = a[14] & g[20163];
assign g[52930] = b[14] & g[20163];
assign g[36548] = a[14] & g[20164];
assign g[52931] = b[14] & g[20164];
assign g[36549] = a[14] & g[20165];
assign g[52932] = b[14] & g[20165];
assign g[36550] = a[14] & g[20166];
assign g[52933] = b[14] & g[20166];
assign g[36551] = a[14] & g[20167];
assign g[52934] = b[14] & g[20167];
assign g[36552] = a[14] & g[20168];
assign g[52935] = b[14] & g[20168];
assign g[36553] = a[14] & g[20169];
assign g[52936] = b[14] & g[20169];
assign g[36554] = a[14] & g[20170];
assign g[52937] = b[14] & g[20170];
assign g[36555] = a[14] & g[20171];
assign g[52938] = b[14] & g[20171];
assign g[36556] = a[14] & g[20172];
assign g[52939] = b[14] & g[20172];
assign g[36557] = a[14] & g[20173];
assign g[52940] = b[14] & g[20173];
assign g[36558] = a[14] & g[20174];
assign g[52941] = b[14] & g[20174];
assign g[36559] = a[14] & g[20175];
assign g[52942] = b[14] & g[20175];
assign g[36560] = a[14] & g[20176];
assign g[52943] = b[14] & g[20176];
assign g[36561] = a[14] & g[20177];
assign g[52944] = b[14] & g[20177];
assign g[36562] = a[14] & g[20178];
assign g[52945] = b[14] & g[20178];
assign g[36563] = a[14] & g[20179];
assign g[52946] = b[14] & g[20179];
assign g[36564] = a[14] & g[20180];
assign g[52947] = b[14] & g[20180];
assign g[36565] = a[14] & g[20181];
assign g[52948] = b[14] & g[20181];
assign g[36566] = a[14] & g[20182];
assign g[52949] = b[14] & g[20182];
assign g[36567] = a[14] & g[20183];
assign g[52950] = b[14] & g[20183];
assign g[36568] = a[14] & g[20184];
assign g[52951] = b[14] & g[20184];
assign g[36569] = a[14] & g[20185];
assign g[52952] = b[14] & g[20185];
assign g[36570] = a[14] & g[20186];
assign g[52953] = b[14] & g[20186];
assign g[36571] = a[14] & g[20187];
assign g[52954] = b[14] & g[20187];
assign g[36572] = a[14] & g[20188];
assign g[52955] = b[14] & g[20188];
assign g[36573] = a[14] & g[20189];
assign g[52956] = b[14] & g[20189];
assign g[36574] = a[14] & g[20190];
assign g[52957] = b[14] & g[20190];
assign g[36575] = a[14] & g[20191];
assign g[52958] = b[14] & g[20191];
assign g[36576] = a[14] & g[20192];
assign g[52959] = b[14] & g[20192];
assign g[36577] = a[14] & g[20193];
assign g[52960] = b[14] & g[20193];
assign g[36578] = a[14] & g[20194];
assign g[52961] = b[14] & g[20194];
assign g[36579] = a[14] & g[20195];
assign g[52962] = b[14] & g[20195];
assign g[36580] = a[14] & g[20196];
assign g[52963] = b[14] & g[20196];
assign g[36581] = a[14] & g[20197];
assign g[52964] = b[14] & g[20197];
assign g[36582] = a[14] & g[20198];
assign g[52965] = b[14] & g[20198];
assign g[36583] = a[14] & g[20199];
assign g[52966] = b[14] & g[20199];
assign g[36584] = a[14] & g[20200];
assign g[52967] = b[14] & g[20200];
assign g[36585] = a[14] & g[20201];
assign g[52968] = b[14] & g[20201];
assign g[36586] = a[14] & g[20202];
assign g[52969] = b[14] & g[20202];
assign g[36587] = a[14] & g[20203];
assign g[52970] = b[14] & g[20203];
assign g[36588] = a[14] & g[20204];
assign g[52971] = b[14] & g[20204];
assign g[36589] = a[14] & g[20205];
assign g[52972] = b[14] & g[20205];
assign g[36590] = a[14] & g[20206];
assign g[52973] = b[14] & g[20206];
assign g[36591] = a[14] & g[20207];
assign g[52974] = b[14] & g[20207];
assign g[36592] = a[14] & g[20208];
assign g[52975] = b[14] & g[20208];
assign g[36593] = a[14] & g[20209];
assign g[52976] = b[14] & g[20209];
assign g[36594] = a[14] & g[20210];
assign g[52977] = b[14] & g[20210];
assign g[36595] = a[14] & g[20211];
assign g[52978] = b[14] & g[20211];
assign g[36596] = a[14] & g[20212];
assign g[52979] = b[14] & g[20212];
assign g[36597] = a[14] & g[20213];
assign g[52980] = b[14] & g[20213];
assign g[36598] = a[14] & g[20214];
assign g[52981] = b[14] & g[20214];
assign g[36599] = a[14] & g[20215];
assign g[52982] = b[14] & g[20215];
assign g[36600] = a[14] & g[20216];
assign g[52983] = b[14] & g[20216];
assign g[36601] = a[14] & g[20217];
assign g[52984] = b[14] & g[20217];
assign g[36602] = a[14] & g[20218];
assign g[52985] = b[14] & g[20218];
assign g[36603] = a[14] & g[20219];
assign g[52986] = b[14] & g[20219];
assign g[36604] = a[14] & g[20220];
assign g[52987] = b[14] & g[20220];
assign g[36605] = a[14] & g[20221];
assign g[52988] = b[14] & g[20221];
assign g[36606] = a[14] & g[20222];
assign g[52989] = b[14] & g[20222];
assign g[36607] = a[14] & g[20223];
assign g[52990] = b[14] & g[20223];
assign g[36608] = a[14] & g[20224];
assign g[52991] = b[14] & g[20224];
assign g[36609] = a[14] & g[20225];
assign g[52992] = b[14] & g[20225];
assign g[36610] = a[14] & g[20226];
assign g[52993] = b[14] & g[20226];
assign g[36611] = a[14] & g[20227];
assign g[52994] = b[14] & g[20227];
assign g[36612] = a[14] & g[20228];
assign g[52995] = b[14] & g[20228];
assign g[36613] = a[14] & g[20229];
assign g[52996] = b[14] & g[20229];
assign g[36614] = a[14] & g[20230];
assign g[52997] = b[14] & g[20230];
assign g[36615] = a[14] & g[20231];
assign g[52998] = b[14] & g[20231];
assign g[36616] = a[14] & g[20232];
assign g[52999] = b[14] & g[20232];
assign g[36617] = a[14] & g[20233];
assign g[53000] = b[14] & g[20233];
assign g[36618] = a[14] & g[20234];
assign g[53001] = b[14] & g[20234];
assign g[36619] = a[14] & g[20235];
assign g[53002] = b[14] & g[20235];
assign g[36620] = a[14] & g[20236];
assign g[53003] = b[14] & g[20236];
assign g[36621] = a[14] & g[20237];
assign g[53004] = b[14] & g[20237];
assign g[36622] = a[14] & g[20238];
assign g[53005] = b[14] & g[20238];
assign g[36623] = a[14] & g[20239];
assign g[53006] = b[14] & g[20239];
assign g[36624] = a[14] & g[20240];
assign g[53007] = b[14] & g[20240];
assign g[36625] = a[14] & g[20241];
assign g[53008] = b[14] & g[20241];
assign g[36626] = a[14] & g[20242];
assign g[53009] = b[14] & g[20242];
assign g[36627] = a[14] & g[20243];
assign g[53010] = b[14] & g[20243];
assign g[36628] = a[14] & g[20244];
assign g[53011] = b[14] & g[20244];
assign g[36629] = a[14] & g[20245];
assign g[53012] = b[14] & g[20245];
assign g[36630] = a[14] & g[20246];
assign g[53013] = b[14] & g[20246];
assign g[36631] = a[14] & g[20247];
assign g[53014] = b[14] & g[20247];
assign g[36632] = a[14] & g[20248];
assign g[53015] = b[14] & g[20248];
assign g[36633] = a[14] & g[20249];
assign g[53016] = b[14] & g[20249];
assign g[36634] = a[14] & g[20250];
assign g[53017] = b[14] & g[20250];
assign g[36635] = a[14] & g[20251];
assign g[53018] = b[14] & g[20251];
assign g[36636] = a[14] & g[20252];
assign g[53019] = b[14] & g[20252];
assign g[36637] = a[14] & g[20253];
assign g[53020] = b[14] & g[20253];
assign g[36638] = a[14] & g[20254];
assign g[53021] = b[14] & g[20254];
assign g[36639] = a[14] & g[20255];
assign g[53022] = b[14] & g[20255];
assign g[36640] = a[14] & g[20256];
assign g[53023] = b[14] & g[20256];
assign g[36641] = a[14] & g[20257];
assign g[53024] = b[14] & g[20257];
assign g[36642] = a[14] & g[20258];
assign g[53025] = b[14] & g[20258];
assign g[36643] = a[14] & g[20259];
assign g[53026] = b[14] & g[20259];
assign g[36644] = a[14] & g[20260];
assign g[53027] = b[14] & g[20260];
assign g[36645] = a[14] & g[20261];
assign g[53028] = b[14] & g[20261];
assign g[36646] = a[14] & g[20262];
assign g[53029] = b[14] & g[20262];
assign g[36647] = a[14] & g[20263];
assign g[53030] = b[14] & g[20263];
assign g[36648] = a[14] & g[20264];
assign g[53031] = b[14] & g[20264];
assign g[36649] = a[14] & g[20265];
assign g[53032] = b[14] & g[20265];
assign g[36650] = a[14] & g[20266];
assign g[53033] = b[14] & g[20266];
assign g[36651] = a[14] & g[20267];
assign g[53034] = b[14] & g[20267];
assign g[36652] = a[14] & g[20268];
assign g[53035] = b[14] & g[20268];
assign g[36653] = a[14] & g[20269];
assign g[53036] = b[14] & g[20269];
assign g[36654] = a[14] & g[20270];
assign g[53037] = b[14] & g[20270];
assign g[36655] = a[14] & g[20271];
assign g[53038] = b[14] & g[20271];
assign g[36656] = a[14] & g[20272];
assign g[53039] = b[14] & g[20272];
assign g[36657] = a[14] & g[20273];
assign g[53040] = b[14] & g[20273];
assign g[36658] = a[14] & g[20274];
assign g[53041] = b[14] & g[20274];
assign g[36659] = a[14] & g[20275];
assign g[53042] = b[14] & g[20275];
assign g[36660] = a[14] & g[20276];
assign g[53043] = b[14] & g[20276];
assign g[36661] = a[14] & g[20277];
assign g[53044] = b[14] & g[20277];
assign g[36662] = a[14] & g[20278];
assign g[53045] = b[14] & g[20278];
assign g[36663] = a[14] & g[20279];
assign g[53046] = b[14] & g[20279];
assign g[36664] = a[14] & g[20280];
assign g[53047] = b[14] & g[20280];
assign g[36665] = a[14] & g[20281];
assign g[53048] = b[14] & g[20281];
assign g[36666] = a[14] & g[20282];
assign g[53049] = b[14] & g[20282];
assign g[36667] = a[14] & g[20283];
assign g[53050] = b[14] & g[20283];
assign g[36668] = a[14] & g[20284];
assign g[53051] = b[14] & g[20284];
assign g[36669] = a[14] & g[20285];
assign g[53052] = b[14] & g[20285];
assign g[36670] = a[14] & g[20286];
assign g[53053] = b[14] & g[20286];
assign g[36671] = a[14] & g[20287];
assign g[53054] = b[14] & g[20287];
assign g[36672] = a[14] & g[20288];
assign g[53055] = b[14] & g[20288];
assign g[36673] = a[14] & g[20289];
assign g[53056] = b[14] & g[20289];
assign g[36674] = a[14] & g[20290];
assign g[53057] = b[14] & g[20290];
assign g[36675] = a[14] & g[20291];
assign g[53058] = b[14] & g[20291];
assign g[36676] = a[14] & g[20292];
assign g[53059] = b[14] & g[20292];
assign g[36677] = a[14] & g[20293];
assign g[53060] = b[14] & g[20293];
assign g[36678] = a[14] & g[20294];
assign g[53061] = b[14] & g[20294];
assign g[36679] = a[14] & g[20295];
assign g[53062] = b[14] & g[20295];
assign g[36680] = a[14] & g[20296];
assign g[53063] = b[14] & g[20296];
assign g[36681] = a[14] & g[20297];
assign g[53064] = b[14] & g[20297];
assign g[36682] = a[14] & g[20298];
assign g[53065] = b[14] & g[20298];
assign g[36683] = a[14] & g[20299];
assign g[53066] = b[14] & g[20299];
assign g[36684] = a[14] & g[20300];
assign g[53067] = b[14] & g[20300];
assign g[36685] = a[14] & g[20301];
assign g[53068] = b[14] & g[20301];
assign g[36686] = a[14] & g[20302];
assign g[53069] = b[14] & g[20302];
assign g[36687] = a[14] & g[20303];
assign g[53070] = b[14] & g[20303];
assign g[36688] = a[14] & g[20304];
assign g[53071] = b[14] & g[20304];
assign g[36689] = a[14] & g[20305];
assign g[53072] = b[14] & g[20305];
assign g[36690] = a[14] & g[20306];
assign g[53073] = b[14] & g[20306];
assign g[36691] = a[14] & g[20307];
assign g[53074] = b[14] & g[20307];
assign g[36692] = a[14] & g[20308];
assign g[53075] = b[14] & g[20308];
assign g[36693] = a[14] & g[20309];
assign g[53076] = b[14] & g[20309];
assign g[36694] = a[14] & g[20310];
assign g[53077] = b[14] & g[20310];
assign g[36695] = a[14] & g[20311];
assign g[53078] = b[14] & g[20311];
assign g[36696] = a[14] & g[20312];
assign g[53079] = b[14] & g[20312];
assign g[36697] = a[14] & g[20313];
assign g[53080] = b[14] & g[20313];
assign g[36698] = a[14] & g[20314];
assign g[53081] = b[14] & g[20314];
assign g[36699] = a[14] & g[20315];
assign g[53082] = b[14] & g[20315];
assign g[36700] = a[14] & g[20316];
assign g[53083] = b[14] & g[20316];
assign g[36701] = a[14] & g[20317];
assign g[53084] = b[14] & g[20317];
assign g[36702] = a[14] & g[20318];
assign g[53085] = b[14] & g[20318];
assign g[36703] = a[14] & g[20319];
assign g[53086] = b[14] & g[20319];
assign g[36704] = a[14] & g[20320];
assign g[53087] = b[14] & g[20320];
assign g[36705] = a[14] & g[20321];
assign g[53088] = b[14] & g[20321];
assign g[36706] = a[14] & g[20322];
assign g[53089] = b[14] & g[20322];
assign g[36707] = a[14] & g[20323];
assign g[53090] = b[14] & g[20323];
assign g[36708] = a[14] & g[20324];
assign g[53091] = b[14] & g[20324];
assign g[36709] = a[14] & g[20325];
assign g[53092] = b[14] & g[20325];
assign g[36710] = a[14] & g[20326];
assign g[53093] = b[14] & g[20326];
assign g[36711] = a[14] & g[20327];
assign g[53094] = b[14] & g[20327];
assign g[36712] = a[14] & g[20328];
assign g[53095] = b[14] & g[20328];
assign g[36713] = a[14] & g[20329];
assign g[53096] = b[14] & g[20329];
assign g[36714] = a[14] & g[20330];
assign g[53097] = b[14] & g[20330];
assign g[36715] = a[14] & g[20331];
assign g[53098] = b[14] & g[20331];
assign g[36716] = a[14] & g[20332];
assign g[53099] = b[14] & g[20332];
assign g[36717] = a[14] & g[20333];
assign g[53100] = b[14] & g[20333];
assign g[36718] = a[14] & g[20334];
assign g[53101] = b[14] & g[20334];
assign g[36719] = a[14] & g[20335];
assign g[53102] = b[14] & g[20335];
assign g[36720] = a[14] & g[20336];
assign g[53103] = b[14] & g[20336];
assign g[36721] = a[14] & g[20337];
assign g[53104] = b[14] & g[20337];
assign g[36722] = a[14] & g[20338];
assign g[53105] = b[14] & g[20338];
assign g[36723] = a[14] & g[20339];
assign g[53106] = b[14] & g[20339];
assign g[36724] = a[14] & g[20340];
assign g[53107] = b[14] & g[20340];
assign g[36725] = a[14] & g[20341];
assign g[53108] = b[14] & g[20341];
assign g[36726] = a[14] & g[20342];
assign g[53109] = b[14] & g[20342];
assign g[36727] = a[14] & g[20343];
assign g[53110] = b[14] & g[20343];
assign g[36728] = a[14] & g[20344];
assign g[53111] = b[14] & g[20344];
assign g[36729] = a[14] & g[20345];
assign g[53112] = b[14] & g[20345];
assign g[36730] = a[14] & g[20346];
assign g[53113] = b[14] & g[20346];
assign g[36731] = a[14] & g[20347];
assign g[53114] = b[14] & g[20347];
assign g[36732] = a[14] & g[20348];
assign g[53115] = b[14] & g[20348];
assign g[36733] = a[14] & g[20349];
assign g[53116] = b[14] & g[20349];
assign g[36734] = a[14] & g[20350];
assign g[53117] = b[14] & g[20350];
assign g[36735] = a[14] & g[20351];
assign g[53118] = b[14] & g[20351];
assign g[36736] = a[14] & g[20352];
assign g[53119] = b[14] & g[20352];
assign g[36737] = a[14] & g[20353];
assign g[53120] = b[14] & g[20353];
assign g[36738] = a[14] & g[20354];
assign g[53121] = b[14] & g[20354];
assign g[36739] = a[14] & g[20355];
assign g[53122] = b[14] & g[20355];
assign g[36740] = a[14] & g[20356];
assign g[53123] = b[14] & g[20356];
assign g[36741] = a[14] & g[20357];
assign g[53124] = b[14] & g[20357];
assign g[36742] = a[14] & g[20358];
assign g[53125] = b[14] & g[20358];
assign g[36743] = a[14] & g[20359];
assign g[53126] = b[14] & g[20359];
assign g[36744] = a[14] & g[20360];
assign g[53127] = b[14] & g[20360];
assign g[36745] = a[14] & g[20361];
assign g[53128] = b[14] & g[20361];
assign g[36746] = a[14] & g[20362];
assign g[53129] = b[14] & g[20362];
assign g[36747] = a[14] & g[20363];
assign g[53130] = b[14] & g[20363];
assign g[36748] = a[14] & g[20364];
assign g[53131] = b[14] & g[20364];
assign g[36749] = a[14] & g[20365];
assign g[53132] = b[14] & g[20365];
assign g[36750] = a[14] & g[20366];
assign g[53133] = b[14] & g[20366];
assign g[36751] = a[14] & g[20367];
assign g[53134] = b[14] & g[20367];
assign g[36752] = a[14] & g[20368];
assign g[53135] = b[14] & g[20368];
assign g[36753] = a[14] & g[20369];
assign g[53136] = b[14] & g[20369];
assign g[36754] = a[14] & g[20370];
assign g[53137] = b[14] & g[20370];
assign g[36755] = a[14] & g[20371];
assign g[53138] = b[14] & g[20371];
assign g[36756] = a[14] & g[20372];
assign g[53139] = b[14] & g[20372];
assign g[36757] = a[14] & g[20373];
assign g[53140] = b[14] & g[20373];
assign g[36758] = a[14] & g[20374];
assign g[53141] = b[14] & g[20374];
assign g[36759] = a[14] & g[20375];
assign g[53142] = b[14] & g[20375];
assign g[36760] = a[14] & g[20376];
assign g[53143] = b[14] & g[20376];
assign g[36761] = a[14] & g[20377];
assign g[53144] = b[14] & g[20377];
assign g[36762] = a[14] & g[20378];
assign g[53145] = b[14] & g[20378];
assign g[36763] = a[14] & g[20379];
assign g[53146] = b[14] & g[20379];
assign g[36764] = a[14] & g[20380];
assign g[53147] = b[14] & g[20380];
assign g[36765] = a[14] & g[20381];
assign g[53148] = b[14] & g[20381];
assign g[36766] = a[14] & g[20382];
assign g[53149] = b[14] & g[20382];
assign g[36767] = a[14] & g[20383];
assign g[53150] = b[14] & g[20383];
assign g[36768] = a[14] & g[20384];
assign g[53151] = b[14] & g[20384];
assign g[36769] = a[14] & g[20385];
assign g[53152] = b[14] & g[20385];
assign g[36770] = a[14] & g[20386];
assign g[53153] = b[14] & g[20386];
assign g[36771] = a[14] & g[20387];
assign g[53154] = b[14] & g[20387];
assign g[36772] = a[14] & g[20388];
assign g[53155] = b[14] & g[20388];
assign g[36773] = a[14] & g[20389];
assign g[53156] = b[14] & g[20389];
assign g[36774] = a[14] & g[20390];
assign g[53157] = b[14] & g[20390];
assign g[36775] = a[14] & g[20391];
assign g[53158] = b[14] & g[20391];
assign g[36776] = a[14] & g[20392];
assign g[53159] = b[14] & g[20392];
assign g[36777] = a[14] & g[20393];
assign g[53160] = b[14] & g[20393];
assign g[36778] = a[14] & g[20394];
assign g[53161] = b[14] & g[20394];
assign g[36779] = a[14] & g[20395];
assign g[53162] = b[14] & g[20395];
assign g[36780] = a[14] & g[20396];
assign g[53163] = b[14] & g[20396];
assign g[36781] = a[14] & g[20397];
assign g[53164] = b[14] & g[20397];
assign g[36782] = a[14] & g[20398];
assign g[53165] = b[14] & g[20398];
assign g[36783] = a[14] & g[20399];
assign g[53166] = b[14] & g[20399];
assign g[36784] = a[14] & g[20400];
assign g[53167] = b[14] & g[20400];
assign g[36785] = a[14] & g[20401];
assign g[53168] = b[14] & g[20401];
assign g[36786] = a[14] & g[20402];
assign g[53169] = b[14] & g[20402];
assign g[36787] = a[14] & g[20403];
assign g[53170] = b[14] & g[20403];
assign g[36788] = a[14] & g[20404];
assign g[53171] = b[14] & g[20404];
assign g[36789] = a[14] & g[20405];
assign g[53172] = b[14] & g[20405];
assign g[36790] = a[14] & g[20406];
assign g[53173] = b[14] & g[20406];
assign g[36791] = a[14] & g[20407];
assign g[53174] = b[14] & g[20407];
assign g[36792] = a[14] & g[20408];
assign g[53175] = b[14] & g[20408];
assign g[36793] = a[14] & g[20409];
assign g[53176] = b[14] & g[20409];
assign g[36794] = a[14] & g[20410];
assign g[53177] = b[14] & g[20410];
assign g[36795] = a[14] & g[20411];
assign g[53178] = b[14] & g[20411];
assign g[36796] = a[14] & g[20412];
assign g[53179] = b[14] & g[20412];
assign g[36797] = a[14] & g[20413];
assign g[53180] = b[14] & g[20413];
assign g[36798] = a[14] & g[20414];
assign g[53181] = b[14] & g[20414];
assign g[36799] = a[14] & g[20415];
assign g[53182] = b[14] & g[20415];
assign g[36800] = a[14] & g[20416];
assign g[53183] = b[14] & g[20416];
assign g[36801] = a[14] & g[20417];
assign g[53184] = b[14] & g[20417];
assign g[36802] = a[14] & g[20418];
assign g[53185] = b[14] & g[20418];
assign g[36803] = a[14] & g[20419];
assign g[53186] = b[14] & g[20419];
assign g[36804] = a[14] & g[20420];
assign g[53187] = b[14] & g[20420];
assign g[36805] = a[14] & g[20421];
assign g[53188] = b[14] & g[20421];
assign g[36806] = a[14] & g[20422];
assign g[53189] = b[14] & g[20422];
assign g[36807] = a[14] & g[20423];
assign g[53190] = b[14] & g[20423];
assign g[36808] = a[14] & g[20424];
assign g[53191] = b[14] & g[20424];
assign g[36809] = a[14] & g[20425];
assign g[53192] = b[14] & g[20425];
assign g[36810] = a[14] & g[20426];
assign g[53193] = b[14] & g[20426];
assign g[36811] = a[14] & g[20427];
assign g[53194] = b[14] & g[20427];
assign g[36812] = a[14] & g[20428];
assign g[53195] = b[14] & g[20428];
assign g[36813] = a[14] & g[20429];
assign g[53196] = b[14] & g[20429];
assign g[36814] = a[14] & g[20430];
assign g[53197] = b[14] & g[20430];
assign g[36815] = a[14] & g[20431];
assign g[53198] = b[14] & g[20431];
assign g[36816] = a[14] & g[20432];
assign g[53199] = b[14] & g[20432];
assign g[36817] = a[14] & g[20433];
assign g[53200] = b[14] & g[20433];
assign g[36818] = a[14] & g[20434];
assign g[53201] = b[14] & g[20434];
assign g[36819] = a[14] & g[20435];
assign g[53202] = b[14] & g[20435];
assign g[36820] = a[14] & g[20436];
assign g[53203] = b[14] & g[20436];
assign g[36821] = a[14] & g[20437];
assign g[53204] = b[14] & g[20437];
assign g[36822] = a[14] & g[20438];
assign g[53205] = b[14] & g[20438];
assign g[36823] = a[14] & g[20439];
assign g[53206] = b[14] & g[20439];
assign g[36824] = a[14] & g[20440];
assign g[53207] = b[14] & g[20440];
assign g[36825] = a[14] & g[20441];
assign g[53208] = b[14] & g[20441];
assign g[36826] = a[14] & g[20442];
assign g[53209] = b[14] & g[20442];
assign g[36827] = a[14] & g[20443];
assign g[53210] = b[14] & g[20443];
assign g[36828] = a[14] & g[20444];
assign g[53211] = b[14] & g[20444];
assign g[36829] = a[14] & g[20445];
assign g[53212] = b[14] & g[20445];
assign g[36830] = a[14] & g[20446];
assign g[53213] = b[14] & g[20446];
assign g[36831] = a[14] & g[20447];
assign g[53214] = b[14] & g[20447];
assign g[36832] = a[14] & g[20448];
assign g[53215] = b[14] & g[20448];
assign g[36833] = a[14] & g[20449];
assign g[53216] = b[14] & g[20449];
assign g[36834] = a[14] & g[20450];
assign g[53217] = b[14] & g[20450];
assign g[36835] = a[14] & g[20451];
assign g[53218] = b[14] & g[20451];
assign g[36836] = a[14] & g[20452];
assign g[53219] = b[14] & g[20452];
assign g[36837] = a[14] & g[20453];
assign g[53220] = b[14] & g[20453];
assign g[36838] = a[14] & g[20454];
assign g[53221] = b[14] & g[20454];
assign g[36839] = a[14] & g[20455];
assign g[53222] = b[14] & g[20455];
assign g[36840] = a[14] & g[20456];
assign g[53223] = b[14] & g[20456];
assign g[36841] = a[14] & g[20457];
assign g[53224] = b[14] & g[20457];
assign g[36842] = a[14] & g[20458];
assign g[53225] = b[14] & g[20458];
assign g[36843] = a[14] & g[20459];
assign g[53226] = b[14] & g[20459];
assign g[36844] = a[14] & g[20460];
assign g[53227] = b[14] & g[20460];
assign g[36845] = a[14] & g[20461];
assign g[53228] = b[14] & g[20461];
assign g[36846] = a[14] & g[20462];
assign g[53229] = b[14] & g[20462];
assign g[36847] = a[14] & g[20463];
assign g[53230] = b[14] & g[20463];
assign g[36848] = a[14] & g[20464];
assign g[53231] = b[14] & g[20464];
assign g[36849] = a[14] & g[20465];
assign g[53232] = b[14] & g[20465];
assign g[36850] = a[14] & g[20466];
assign g[53233] = b[14] & g[20466];
assign g[36851] = a[14] & g[20467];
assign g[53234] = b[14] & g[20467];
assign g[36852] = a[14] & g[20468];
assign g[53235] = b[14] & g[20468];
assign g[36853] = a[14] & g[20469];
assign g[53236] = b[14] & g[20469];
assign g[36854] = a[14] & g[20470];
assign g[53237] = b[14] & g[20470];
assign g[36855] = a[14] & g[20471];
assign g[53238] = b[14] & g[20471];
assign g[36856] = a[14] & g[20472];
assign g[53239] = b[14] & g[20472];
assign g[36857] = a[14] & g[20473];
assign g[53240] = b[14] & g[20473];
assign g[36858] = a[14] & g[20474];
assign g[53241] = b[14] & g[20474];
assign g[36859] = a[14] & g[20475];
assign g[53242] = b[14] & g[20475];
assign g[36860] = a[14] & g[20476];
assign g[53243] = b[14] & g[20476];
assign g[36861] = a[14] & g[20477];
assign g[53244] = b[14] & g[20477];
assign g[36862] = a[14] & g[20478];
assign g[53245] = b[14] & g[20478];
assign g[36863] = a[14] & g[20479];
assign g[53246] = b[14] & g[20479];
assign g[36864] = a[14] & g[20480];
assign g[53247] = b[14] & g[20480];
assign g[36865] = a[14] & g[20481];
assign g[53248] = b[14] & g[20481];
assign g[36866] = a[14] & g[20482];
assign g[53249] = b[14] & g[20482];
assign g[36867] = a[14] & g[20483];
assign g[53250] = b[14] & g[20483];
assign g[36868] = a[14] & g[20484];
assign g[53251] = b[14] & g[20484];
assign g[36869] = a[14] & g[20485];
assign g[53252] = b[14] & g[20485];
assign g[36870] = a[14] & g[20486];
assign g[53253] = b[14] & g[20486];
assign g[36871] = a[14] & g[20487];
assign g[53254] = b[14] & g[20487];
assign g[36872] = a[14] & g[20488];
assign g[53255] = b[14] & g[20488];
assign g[36873] = a[14] & g[20489];
assign g[53256] = b[14] & g[20489];
assign g[36874] = a[14] & g[20490];
assign g[53257] = b[14] & g[20490];
assign g[36875] = a[14] & g[20491];
assign g[53258] = b[14] & g[20491];
assign g[36876] = a[14] & g[20492];
assign g[53259] = b[14] & g[20492];
assign g[36877] = a[14] & g[20493];
assign g[53260] = b[14] & g[20493];
assign g[36878] = a[14] & g[20494];
assign g[53261] = b[14] & g[20494];
assign g[36879] = a[14] & g[20495];
assign g[53262] = b[14] & g[20495];
assign g[36880] = a[14] & g[20496];
assign g[53263] = b[14] & g[20496];
assign g[36881] = a[14] & g[20497];
assign g[53264] = b[14] & g[20497];
assign g[36882] = a[14] & g[20498];
assign g[53265] = b[14] & g[20498];
assign g[36883] = a[14] & g[20499];
assign g[53266] = b[14] & g[20499];
assign g[36884] = a[14] & g[20500];
assign g[53267] = b[14] & g[20500];
assign g[36885] = a[14] & g[20501];
assign g[53268] = b[14] & g[20501];
assign g[36886] = a[14] & g[20502];
assign g[53269] = b[14] & g[20502];
assign g[36887] = a[14] & g[20503];
assign g[53270] = b[14] & g[20503];
assign g[36888] = a[14] & g[20504];
assign g[53271] = b[14] & g[20504];
assign g[36889] = a[14] & g[20505];
assign g[53272] = b[14] & g[20505];
assign g[36890] = a[14] & g[20506];
assign g[53273] = b[14] & g[20506];
assign g[36891] = a[14] & g[20507];
assign g[53274] = b[14] & g[20507];
assign g[36892] = a[14] & g[20508];
assign g[53275] = b[14] & g[20508];
assign g[36893] = a[14] & g[20509];
assign g[53276] = b[14] & g[20509];
assign g[36894] = a[14] & g[20510];
assign g[53277] = b[14] & g[20510];
assign g[36895] = a[14] & g[20511];
assign g[53278] = b[14] & g[20511];
assign g[36896] = a[14] & g[20512];
assign g[53279] = b[14] & g[20512];
assign g[36897] = a[14] & g[20513];
assign g[53280] = b[14] & g[20513];
assign g[36898] = a[14] & g[20514];
assign g[53281] = b[14] & g[20514];
assign g[36899] = a[14] & g[20515];
assign g[53282] = b[14] & g[20515];
assign g[36900] = a[14] & g[20516];
assign g[53283] = b[14] & g[20516];
assign g[36901] = a[14] & g[20517];
assign g[53284] = b[14] & g[20517];
assign g[36902] = a[14] & g[20518];
assign g[53285] = b[14] & g[20518];
assign g[36903] = a[14] & g[20519];
assign g[53286] = b[14] & g[20519];
assign g[36904] = a[14] & g[20520];
assign g[53287] = b[14] & g[20520];
assign g[36905] = a[14] & g[20521];
assign g[53288] = b[14] & g[20521];
assign g[36906] = a[14] & g[20522];
assign g[53289] = b[14] & g[20522];
assign g[36907] = a[14] & g[20523];
assign g[53290] = b[14] & g[20523];
assign g[36908] = a[14] & g[20524];
assign g[53291] = b[14] & g[20524];
assign g[36909] = a[14] & g[20525];
assign g[53292] = b[14] & g[20525];
assign g[36910] = a[14] & g[20526];
assign g[53293] = b[14] & g[20526];
assign g[36911] = a[14] & g[20527];
assign g[53294] = b[14] & g[20527];
assign g[36912] = a[14] & g[20528];
assign g[53295] = b[14] & g[20528];
assign g[36913] = a[14] & g[20529];
assign g[53296] = b[14] & g[20529];
assign g[36914] = a[14] & g[20530];
assign g[53297] = b[14] & g[20530];
assign g[36915] = a[14] & g[20531];
assign g[53298] = b[14] & g[20531];
assign g[36916] = a[14] & g[20532];
assign g[53299] = b[14] & g[20532];
assign g[36917] = a[14] & g[20533];
assign g[53300] = b[14] & g[20533];
assign g[36918] = a[14] & g[20534];
assign g[53301] = b[14] & g[20534];
assign g[36919] = a[14] & g[20535];
assign g[53302] = b[14] & g[20535];
assign g[36920] = a[14] & g[20536];
assign g[53303] = b[14] & g[20536];
assign g[36921] = a[14] & g[20537];
assign g[53304] = b[14] & g[20537];
assign g[36922] = a[14] & g[20538];
assign g[53305] = b[14] & g[20538];
assign g[36923] = a[14] & g[20539];
assign g[53306] = b[14] & g[20539];
assign g[36924] = a[14] & g[20540];
assign g[53307] = b[14] & g[20540];
assign g[36925] = a[14] & g[20541];
assign g[53308] = b[14] & g[20541];
assign g[36926] = a[14] & g[20542];
assign g[53309] = b[14] & g[20542];
assign g[36927] = a[14] & g[20543];
assign g[53310] = b[14] & g[20543];
assign g[36928] = a[14] & g[20544];
assign g[53311] = b[14] & g[20544];
assign g[36929] = a[14] & g[20545];
assign g[53312] = b[14] & g[20545];
assign g[36930] = a[14] & g[20546];
assign g[53313] = b[14] & g[20546];
assign g[36931] = a[14] & g[20547];
assign g[53314] = b[14] & g[20547];
assign g[36932] = a[14] & g[20548];
assign g[53315] = b[14] & g[20548];
assign g[36933] = a[14] & g[20549];
assign g[53316] = b[14] & g[20549];
assign g[36934] = a[14] & g[20550];
assign g[53317] = b[14] & g[20550];
assign g[36935] = a[14] & g[20551];
assign g[53318] = b[14] & g[20551];
assign g[36936] = a[14] & g[20552];
assign g[53319] = b[14] & g[20552];
assign g[36937] = a[14] & g[20553];
assign g[53320] = b[14] & g[20553];
assign g[36938] = a[14] & g[20554];
assign g[53321] = b[14] & g[20554];
assign g[36939] = a[14] & g[20555];
assign g[53322] = b[14] & g[20555];
assign g[36940] = a[14] & g[20556];
assign g[53323] = b[14] & g[20556];
assign g[36941] = a[14] & g[20557];
assign g[53324] = b[14] & g[20557];
assign g[36942] = a[14] & g[20558];
assign g[53325] = b[14] & g[20558];
assign g[36943] = a[14] & g[20559];
assign g[53326] = b[14] & g[20559];
assign g[36944] = a[14] & g[20560];
assign g[53327] = b[14] & g[20560];
assign g[36945] = a[14] & g[20561];
assign g[53328] = b[14] & g[20561];
assign g[36946] = a[14] & g[20562];
assign g[53329] = b[14] & g[20562];
assign g[36947] = a[14] & g[20563];
assign g[53330] = b[14] & g[20563];
assign g[36948] = a[14] & g[20564];
assign g[53331] = b[14] & g[20564];
assign g[36949] = a[14] & g[20565];
assign g[53332] = b[14] & g[20565];
assign g[36950] = a[14] & g[20566];
assign g[53333] = b[14] & g[20566];
assign g[36951] = a[14] & g[20567];
assign g[53334] = b[14] & g[20567];
assign g[36952] = a[14] & g[20568];
assign g[53335] = b[14] & g[20568];
assign g[36953] = a[14] & g[20569];
assign g[53336] = b[14] & g[20569];
assign g[36954] = a[14] & g[20570];
assign g[53337] = b[14] & g[20570];
assign g[36955] = a[14] & g[20571];
assign g[53338] = b[14] & g[20571];
assign g[36956] = a[14] & g[20572];
assign g[53339] = b[14] & g[20572];
assign g[36957] = a[14] & g[20573];
assign g[53340] = b[14] & g[20573];
assign g[36958] = a[14] & g[20574];
assign g[53341] = b[14] & g[20574];
assign g[36959] = a[14] & g[20575];
assign g[53342] = b[14] & g[20575];
assign g[36960] = a[14] & g[20576];
assign g[53343] = b[14] & g[20576];
assign g[36961] = a[14] & g[20577];
assign g[53344] = b[14] & g[20577];
assign g[36962] = a[14] & g[20578];
assign g[53345] = b[14] & g[20578];
assign g[36963] = a[14] & g[20579];
assign g[53346] = b[14] & g[20579];
assign g[36964] = a[14] & g[20580];
assign g[53347] = b[14] & g[20580];
assign g[36965] = a[14] & g[20581];
assign g[53348] = b[14] & g[20581];
assign g[36966] = a[14] & g[20582];
assign g[53349] = b[14] & g[20582];
assign g[36967] = a[14] & g[20583];
assign g[53350] = b[14] & g[20583];
assign g[36968] = a[14] & g[20584];
assign g[53351] = b[14] & g[20584];
assign g[36969] = a[14] & g[20585];
assign g[53352] = b[14] & g[20585];
assign g[36970] = a[14] & g[20586];
assign g[53353] = b[14] & g[20586];
assign g[36971] = a[14] & g[20587];
assign g[53354] = b[14] & g[20587];
assign g[36972] = a[14] & g[20588];
assign g[53355] = b[14] & g[20588];
assign g[36973] = a[14] & g[20589];
assign g[53356] = b[14] & g[20589];
assign g[36974] = a[14] & g[20590];
assign g[53357] = b[14] & g[20590];
assign g[36975] = a[14] & g[20591];
assign g[53358] = b[14] & g[20591];
assign g[36976] = a[14] & g[20592];
assign g[53359] = b[14] & g[20592];
assign g[36977] = a[14] & g[20593];
assign g[53360] = b[14] & g[20593];
assign g[36978] = a[14] & g[20594];
assign g[53361] = b[14] & g[20594];
assign g[36979] = a[14] & g[20595];
assign g[53362] = b[14] & g[20595];
assign g[36980] = a[14] & g[20596];
assign g[53363] = b[14] & g[20596];
assign g[36981] = a[14] & g[20597];
assign g[53364] = b[14] & g[20597];
assign g[36982] = a[14] & g[20598];
assign g[53365] = b[14] & g[20598];
assign g[36983] = a[14] & g[20599];
assign g[53366] = b[14] & g[20599];
assign g[36984] = a[14] & g[20600];
assign g[53367] = b[14] & g[20600];
assign g[36985] = a[14] & g[20601];
assign g[53368] = b[14] & g[20601];
assign g[36986] = a[14] & g[20602];
assign g[53369] = b[14] & g[20602];
assign g[36987] = a[14] & g[20603];
assign g[53370] = b[14] & g[20603];
assign g[36988] = a[14] & g[20604];
assign g[53371] = b[14] & g[20604];
assign g[36989] = a[14] & g[20605];
assign g[53372] = b[14] & g[20605];
assign g[36990] = a[14] & g[20606];
assign g[53373] = b[14] & g[20606];
assign g[36991] = a[14] & g[20607];
assign g[53374] = b[14] & g[20607];
assign g[36992] = a[14] & g[20608];
assign g[53375] = b[14] & g[20608];
assign g[36993] = a[14] & g[20609];
assign g[53376] = b[14] & g[20609];
assign g[36994] = a[14] & g[20610];
assign g[53377] = b[14] & g[20610];
assign g[36995] = a[14] & g[20611];
assign g[53378] = b[14] & g[20611];
assign g[36996] = a[14] & g[20612];
assign g[53379] = b[14] & g[20612];
assign g[36997] = a[14] & g[20613];
assign g[53380] = b[14] & g[20613];
assign g[36998] = a[14] & g[20614];
assign g[53381] = b[14] & g[20614];
assign g[36999] = a[14] & g[20615];
assign g[53382] = b[14] & g[20615];
assign g[37000] = a[14] & g[20616];
assign g[53383] = b[14] & g[20616];
assign g[37001] = a[14] & g[20617];
assign g[53384] = b[14] & g[20617];
assign g[37002] = a[14] & g[20618];
assign g[53385] = b[14] & g[20618];
assign g[37003] = a[14] & g[20619];
assign g[53386] = b[14] & g[20619];
assign g[37004] = a[14] & g[20620];
assign g[53387] = b[14] & g[20620];
assign g[37005] = a[14] & g[20621];
assign g[53388] = b[14] & g[20621];
assign g[37006] = a[14] & g[20622];
assign g[53389] = b[14] & g[20622];
assign g[37007] = a[14] & g[20623];
assign g[53390] = b[14] & g[20623];
assign g[37008] = a[14] & g[20624];
assign g[53391] = b[14] & g[20624];
assign g[37009] = a[14] & g[20625];
assign g[53392] = b[14] & g[20625];
assign g[37010] = a[14] & g[20626];
assign g[53393] = b[14] & g[20626];
assign g[37011] = a[14] & g[20627];
assign g[53394] = b[14] & g[20627];
assign g[37012] = a[14] & g[20628];
assign g[53395] = b[14] & g[20628];
assign g[37013] = a[14] & g[20629];
assign g[53396] = b[14] & g[20629];
assign g[37014] = a[14] & g[20630];
assign g[53397] = b[14] & g[20630];
assign g[37015] = a[14] & g[20631];
assign g[53398] = b[14] & g[20631];
assign g[37016] = a[14] & g[20632];
assign g[53399] = b[14] & g[20632];
assign g[37017] = a[14] & g[20633];
assign g[53400] = b[14] & g[20633];
assign g[37018] = a[14] & g[20634];
assign g[53401] = b[14] & g[20634];
assign g[37019] = a[14] & g[20635];
assign g[53402] = b[14] & g[20635];
assign g[37020] = a[14] & g[20636];
assign g[53403] = b[14] & g[20636];
assign g[37021] = a[14] & g[20637];
assign g[53404] = b[14] & g[20637];
assign g[37022] = a[14] & g[20638];
assign g[53405] = b[14] & g[20638];
assign g[37023] = a[14] & g[20639];
assign g[53406] = b[14] & g[20639];
assign g[37024] = a[14] & g[20640];
assign g[53407] = b[14] & g[20640];
assign g[37025] = a[14] & g[20641];
assign g[53408] = b[14] & g[20641];
assign g[37026] = a[14] & g[20642];
assign g[53409] = b[14] & g[20642];
assign g[37027] = a[14] & g[20643];
assign g[53410] = b[14] & g[20643];
assign g[37028] = a[14] & g[20644];
assign g[53411] = b[14] & g[20644];
assign g[37029] = a[14] & g[20645];
assign g[53412] = b[14] & g[20645];
assign g[37030] = a[14] & g[20646];
assign g[53413] = b[14] & g[20646];
assign g[37031] = a[14] & g[20647];
assign g[53414] = b[14] & g[20647];
assign g[37032] = a[14] & g[20648];
assign g[53415] = b[14] & g[20648];
assign g[37033] = a[14] & g[20649];
assign g[53416] = b[14] & g[20649];
assign g[37034] = a[14] & g[20650];
assign g[53417] = b[14] & g[20650];
assign g[37035] = a[14] & g[20651];
assign g[53418] = b[14] & g[20651];
assign g[37036] = a[14] & g[20652];
assign g[53419] = b[14] & g[20652];
assign g[37037] = a[14] & g[20653];
assign g[53420] = b[14] & g[20653];
assign g[37038] = a[14] & g[20654];
assign g[53421] = b[14] & g[20654];
assign g[37039] = a[14] & g[20655];
assign g[53422] = b[14] & g[20655];
assign g[37040] = a[14] & g[20656];
assign g[53423] = b[14] & g[20656];
assign g[37041] = a[14] & g[20657];
assign g[53424] = b[14] & g[20657];
assign g[37042] = a[14] & g[20658];
assign g[53425] = b[14] & g[20658];
assign g[37043] = a[14] & g[20659];
assign g[53426] = b[14] & g[20659];
assign g[37044] = a[14] & g[20660];
assign g[53427] = b[14] & g[20660];
assign g[37045] = a[14] & g[20661];
assign g[53428] = b[14] & g[20661];
assign g[37046] = a[14] & g[20662];
assign g[53429] = b[14] & g[20662];
assign g[37047] = a[14] & g[20663];
assign g[53430] = b[14] & g[20663];
assign g[37048] = a[14] & g[20664];
assign g[53431] = b[14] & g[20664];
assign g[37049] = a[14] & g[20665];
assign g[53432] = b[14] & g[20665];
assign g[37050] = a[14] & g[20666];
assign g[53433] = b[14] & g[20666];
assign g[37051] = a[14] & g[20667];
assign g[53434] = b[14] & g[20667];
assign g[37052] = a[14] & g[20668];
assign g[53435] = b[14] & g[20668];
assign g[37053] = a[14] & g[20669];
assign g[53436] = b[14] & g[20669];
assign g[37054] = a[14] & g[20670];
assign g[53437] = b[14] & g[20670];
assign g[37055] = a[14] & g[20671];
assign g[53438] = b[14] & g[20671];
assign g[37056] = a[14] & g[20672];
assign g[53439] = b[14] & g[20672];
assign g[37057] = a[14] & g[20673];
assign g[53440] = b[14] & g[20673];
assign g[37058] = a[14] & g[20674];
assign g[53441] = b[14] & g[20674];
assign g[37059] = a[14] & g[20675];
assign g[53442] = b[14] & g[20675];
assign g[37060] = a[14] & g[20676];
assign g[53443] = b[14] & g[20676];
assign g[37061] = a[14] & g[20677];
assign g[53444] = b[14] & g[20677];
assign g[37062] = a[14] & g[20678];
assign g[53445] = b[14] & g[20678];
assign g[37063] = a[14] & g[20679];
assign g[53446] = b[14] & g[20679];
assign g[37064] = a[14] & g[20680];
assign g[53447] = b[14] & g[20680];
assign g[37065] = a[14] & g[20681];
assign g[53448] = b[14] & g[20681];
assign g[37066] = a[14] & g[20682];
assign g[53449] = b[14] & g[20682];
assign g[37067] = a[14] & g[20683];
assign g[53450] = b[14] & g[20683];
assign g[37068] = a[14] & g[20684];
assign g[53451] = b[14] & g[20684];
assign g[37069] = a[14] & g[20685];
assign g[53452] = b[14] & g[20685];
assign g[37070] = a[14] & g[20686];
assign g[53453] = b[14] & g[20686];
assign g[37071] = a[14] & g[20687];
assign g[53454] = b[14] & g[20687];
assign g[37072] = a[14] & g[20688];
assign g[53455] = b[14] & g[20688];
assign g[37073] = a[14] & g[20689];
assign g[53456] = b[14] & g[20689];
assign g[37074] = a[14] & g[20690];
assign g[53457] = b[14] & g[20690];
assign g[37075] = a[14] & g[20691];
assign g[53458] = b[14] & g[20691];
assign g[37076] = a[14] & g[20692];
assign g[53459] = b[14] & g[20692];
assign g[37077] = a[14] & g[20693];
assign g[53460] = b[14] & g[20693];
assign g[37078] = a[14] & g[20694];
assign g[53461] = b[14] & g[20694];
assign g[37079] = a[14] & g[20695];
assign g[53462] = b[14] & g[20695];
assign g[37080] = a[14] & g[20696];
assign g[53463] = b[14] & g[20696];
assign g[37081] = a[14] & g[20697];
assign g[53464] = b[14] & g[20697];
assign g[37082] = a[14] & g[20698];
assign g[53465] = b[14] & g[20698];
assign g[37083] = a[14] & g[20699];
assign g[53466] = b[14] & g[20699];
assign g[37084] = a[14] & g[20700];
assign g[53467] = b[14] & g[20700];
assign g[37085] = a[14] & g[20701];
assign g[53468] = b[14] & g[20701];
assign g[37086] = a[14] & g[20702];
assign g[53469] = b[14] & g[20702];
assign g[37087] = a[14] & g[20703];
assign g[53470] = b[14] & g[20703];
assign g[37088] = a[14] & g[20704];
assign g[53471] = b[14] & g[20704];
assign g[37089] = a[14] & g[20705];
assign g[53472] = b[14] & g[20705];
assign g[37090] = a[14] & g[20706];
assign g[53473] = b[14] & g[20706];
assign g[37091] = a[14] & g[20707];
assign g[53474] = b[14] & g[20707];
assign g[37092] = a[14] & g[20708];
assign g[53475] = b[14] & g[20708];
assign g[37093] = a[14] & g[20709];
assign g[53476] = b[14] & g[20709];
assign g[37094] = a[14] & g[20710];
assign g[53477] = b[14] & g[20710];
assign g[37095] = a[14] & g[20711];
assign g[53478] = b[14] & g[20711];
assign g[37096] = a[14] & g[20712];
assign g[53479] = b[14] & g[20712];
assign g[37097] = a[14] & g[20713];
assign g[53480] = b[14] & g[20713];
assign g[37098] = a[14] & g[20714];
assign g[53481] = b[14] & g[20714];
assign g[37099] = a[14] & g[20715];
assign g[53482] = b[14] & g[20715];
assign g[37100] = a[14] & g[20716];
assign g[53483] = b[14] & g[20716];
assign g[37101] = a[14] & g[20717];
assign g[53484] = b[14] & g[20717];
assign g[37102] = a[14] & g[20718];
assign g[53485] = b[14] & g[20718];
assign g[37103] = a[14] & g[20719];
assign g[53486] = b[14] & g[20719];
assign g[37104] = a[14] & g[20720];
assign g[53487] = b[14] & g[20720];
assign g[37105] = a[14] & g[20721];
assign g[53488] = b[14] & g[20721];
assign g[37106] = a[14] & g[20722];
assign g[53489] = b[14] & g[20722];
assign g[37107] = a[14] & g[20723];
assign g[53490] = b[14] & g[20723];
assign g[37108] = a[14] & g[20724];
assign g[53491] = b[14] & g[20724];
assign g[37109] = a[14] & g[20725];
assign g[53492] = b[14] & g[20725];
assign g[37110] = a[14] & g[20726];
assign g[53493] = b[14] & g[20726];
assign g[37111] = a[14] & g[20727];
assign g[53494] = b[14] & g[20727];
assign g[37112] = a[14] & g[20728];
assign g[53495] = b[14] & g[20728];
assign g[37113] = a[14] & g[20729];
assign g[53496] = b[14] & g[20729];
assign g[37114] = a[14] & g[20730];
assign g[53497] = b[14] & g[20730];
assign g[37115] = a[14] & g[20731];
assign g[53498] = b[14] & g[20731];
assign g[37116] = a[14] & g[20732];
assign g[53499] = b[14] & g[20732];
assign g[37117] = a[14] & g[20733];
assign g[53500] = b[14] & g[20733];
assign g[37118] = a[14] & g[20734];
assign g[53501] = b[14] & g[20734];
assign g[37119] = a[14] & g[20735];
assign g[53502] = b[14] & g[20735];
assign g[37120] = a[14] & g[20736];
assign g[53503] = b[14] & g[20736];
assign g[37121] = a[14] & g[20737];
assign g[53504] = b[14] & g[20737];
assign g[37122] = a[14] & g[20738];
assign g[53505] = b[14] & g[20738];
assign g[37123] = a[14] & g[20739];
assign g[53506] = b[14] & g[20739];
assign g[37124] = a[14] & g[20740];
assign g[53507] = b[14] & g[20740];
assign g[37125] = a[14] & g[20741];
assign g[53508] = b[14] & g[20741];
assign g[37126] = a[14] & g[20742];
assign g[53509] = b[14] & g[20742];
assign g[37127] = a[14] & g[20743];
assign g[53510] = b[14] & g[20743];
assign g[37128] = a[14] & g[20744];
assign g[53511] = b[14] & g[20744];
assign g[37129] = a[14] & g[20745];
assign g[53512] = b[14] & g[20745];
assign g[37130] = a[14] & g[20746];
assign g[53513] = b[14] & g[20746];
assign g[37131] = a[14] & g[20747];
assign g[53514] = b[14] & g[20747];
assign g[37132] = a[14] & g[20748];
assign g[53515] = b[14] & g[20748];
assign g[37133] = a[14] & g[20749];
assign g[53516] = b[14] & g[20749];
assign g[37134] = a[14] & g[20750];
assign g[53517] = b[14] & g[20750];
assign g[37135] = a[14] & g[20751];
assign g[53518] = b[14] & g[20751];
assign g[37136] = a[14] & g[20752];
assign g[53519] = b[14] & g[20752];
assign g[37137] = a[14] & g[20753];
assign g[53520] = b[14] & g[20753];
assign g[37138] = a[14] & g[20754];
assign g[53521] = b[14] & g[20754];
assign g[37139] = a[14] & g[20755];
assign g[53522] = b[14] & g[20755];
assign g[37140] = a[14] & g[20756];
assign g[53523] = b[14] & g[20756];
assign g[37141] = a[14] & g[20757];
assign g[53524] = b[14] & g[20757];
assign g[37142] = a[14] & g[20758];
assign g[53525] = b[14] & g[20758];
assign g[37143] = a[14] & g[20759];
assign g[53526] = b[14] & g[20759];
assign g[37144] = a[14] & g[20760];
assign g[53527] = b[14] & g[20760];
assign g[37145] = a[14] & g[20761];
assign g[53528] = b[14] & g[20761];
assign g[37146] = a[14] & g[20762];
assign g[53529] = b[14] & g[20762];
assign g[37147] = a[14] & g[20763];
assign g[53530] = b[14] & g[20763];
assign g[37148] = a[14] & g[20764];
assign g[53531] = b[14] & g[20764];
assign g[37149] = a[14] & g[20765];
assign g[53532] = b[14] & g[20765];
assign g[37150] = a[14] & g[20766];
assign g[53533] = b[14] & g[20766];
assign g[37151] = a[14] & g[20767];
assign g[53534] = b[14] & g[20767];
assign g[37152] = a[14] & g[20768];
assign g[53535] = b[14] & g[20768];
assign g[37153] = a[14] & g[20769];
assign g[53536] = b[14] & g[20769];
assign g[37154] = a[14] & g[20770];
assign g[53537] = b[14] & g[20770];
assign g[37155] = a[14] & g[20771];
assign g[53538] = b[14] & g[20771];
assign g[37156] = a[14] & g[20772];
assign g[53539] = b[14] & g[20772];
assign g[37157] = a[14] & g[20773];
assign g[53540] = b[14] & g[20773];
assign g[37158] = a[14] & g[20774];
assign g[53541] = b[14] & g[20774];
assign g[37159] = a[14] & g[20775];
assign g[53542] = b[14] & g[20775];
assign g[37160] = a[14] & g[20776];
assign g[53543] = b[14] & g[20776];
assign g[37161] = a[14] & g[20777];
assign g[53544] = b[14] & g[20777];
assign g[37162] = a[14] & g[20778];
assign g[53545] = b[14] & g[20778];
assign g[37163] = a[14] & g[20779];
assign g[53546] = b[14] & g[20779];
assign g[37164] = a[14] & g[20780];
assign g[53547] = b[14] & g[20780];
assign g[37165] = a[14] & g[20781];
assign g[53548] = b[14] & g[20781];
assign g[37166] = a[14] & g[20782];
assign g[53549] = b[14] & g[20782];
assign g[37167] = a[14] & g[20783];
assign g[53550] = b[14] & g[20783];
assign g[37168] = a[14] & g[20784];
assign g[53551] = b[14] & g[20784];
assign g[37169] = a[14] & g[20785];
assign g[53552] = b[14] & g[20785];
assign g[37170] = a[14] & g[20786];
assign g[53553] = b[14] & g[20786];
assign g[37171] = a[14] & g[20787];
assign g[53554] = b[14] & g[20787];
assign g[37172] = a[14] & g[20788];
assign g[53555] = b[14] & g[20788];
assign g[37173] = a[14] & g[20789];
assign g[53556] = b[14] & g[20789];
assign g[37174] = a[14] & g[20790];
assign g[53557] = b[14] & g[20790];
assign g[37175] = a[14] & g[20791];
assign g[53558] = b[14] & g[20791];
assign g[37176] = a[14] & g[20792];
assign g[53559] = b[14] & g[20792];
assign g[37177] = a[14] & g[20793];
assign g[53560] = b[14] & g[20793];
assign g[37178] = a[14] & g[20794];
assign g[53561] = b[14] & g[20794];
assign g[37179] = a[14] & g[20795];
assign g[53562] = b[14] & g[20795];
assign g[37180] = a[14] & g[20796];
assign g[53563] = b[14] & g[20796];
assign g[37181] = a[14] & g[20797];
assign g[53564] = b[14] & g[20797];
assign g[37182] = a[14] & g[20798];
assign g[53565] = b[14] & g[20798];
assign g[37183] = a[14] & g[20799];
assign g[53566] = b[14] & g[20799];
assign g[37184] = a[14] & g[20800];
assign g[53567] = b[14] & g[20800];
assign g[37185] = a[14] & g[20801];
assign g[53568] = b[14] & g[20801];
assign g[37186] = a[14] & g[20802];
assign g[53569] = b[14] & g[20802];
assign g[37187] = a[14] & g[20803];
assign g[53570] = b[14] & g[20803];
assign g[37188] = a[14] & g[20804];
assign g[53571] = b[14] & g[20804];
assign g[37189] = a[14] & g[20805];
assign g[53572] = b[14] & g[20805];
assign g[37190] = a[14] & g[20806];
assign g[53573] = b[14] & g[20806];
assign g[37191] = a[14] & g[20807];
assign g[53574] = b[14] & g[20807];
assign g[37192] = a[14] & g[20808];
assign g[53575] = b[14] & g[20808];
assign g[37193] = a[14] & g[20809];
assign g[53576] = b[14] & g[20809];
assign g[37194] = a[14] & g[20810];
assign g[53577] = b[14] & g[20810];
assign g[37195] = a[14] & g[20811];
assign g[53578] = b[14] & g[20811];
assign g[37196] = a[14] & g[20812];
assign g[53579] = b[14] & g[20812];
assign g[37197] = a[14] & g[20813];
assign g[53580] = b[14] & g[20813];
assign g[37198] = a[14] & g[20814];
assign g[53581] = b[14] & g[20814];
assign g[37199] = a[14] & g[20815];
assign g[53582] = b[14] & g[20815];
assign g[37200] = a[14] & g[20816];
assign g[53583] = b[14] & g[20816];
assign g[37201] = a[14] & g[20817];
assign g[53584] = b[14] & g[20817];
assign g[37202] = a[14] & g[20818];
assign g[53585] = b[14] & g[20818];
assign g[37203] = a[14] & g[20819];
assign g[53586] = b[14] & g[20819];
assign g[37204] = a[14] & g[20820];
assign g[53587] = b[14] & g[20820];
assign g[37205] = a[14] & g[20821];
assign g[53588] = b[14] & g[20821];
assign g[37206] = a[14] & g[20822];
assign g[53589] = b[14] & g[20822];
assign g[37207] = a[14] & g[20823];
assign g[53590] = b[14] & g[20823];
assign g[37208] = a[14] & g[20824];
assign g[53591] = b[14] & g[20824];
assign g[37209] = a[14] & g[20825];
assign g[53592] = b[14] & g[20825];
assign g[37210] = a[14] & g[20826];
assign g[53593] = b[14] & g[20826];
assign g[37211] = a[14] & g[20827];
assign g[53594] = b[14] & g[20827];
assign g[37212] = a[14] & g[20828];
assign g[53595] = b[14] & g[20828];
assign g[37213] = a[14] & g[20829];
assign g[53596] = b[14] & g[20829];
assign g[37214] = a[14] & g[20830];
assign g[53597] = b[14] & g[20830];
assign g[37215] = a[14] & g[20831];
assign g[53598] = b[14] & g[20831];
assign g[37216] = a[14] & g[20832];
assign g[53599] = b[14] & g[20832];
assign g[37217] = a[14] & g[20833];
assign g[53600] = b[14] & g[20833];
assign g[37218] = a[14] & g[20834];
assign g[53601] = b[14] & g[20834];
assign g[37219] = a[14] & g[20835];
assign g[53602] = b[14] & g[20835];
assign g[37220] = a[14] & g[20836];
assign g[53603] = b[14] & g[20836];
assign g[37221] = a[14] & g[20837];
assign g[53604] = b[14] & g[20837];
assign g[37222] = a[14] & g[20838];
assign g[53605] = b[14] & g[20838];
assign g[37223] = a[14] & g[20839];
assign g[53606] = b[14] & g[20839];
assign g[37224] = a[14] & g[20840];
assign g[53607] = b[14] & g[20840];
assign g[37225] = a[14] & g[20841];
assign g[53608] = b[14] & g[20841];
assign g[37226] = a[14] & g[20842];
assign g[53609] = b[14] & g[20842];
assign g[37227] = a[14] & g[20843];
assign g[53610] = b[14] & g[20843];
assign g[37228] = a[14] & g[20844];
assign g[53611] = b[14] & g[20844];
assign g[37229] = a[14] & g[20845];
assign g[53612] = b[14] & g[20845];
assign g[37230] = a[14] & g[20846];
assign g[53613] = b[14] & g[20846];
assign g[37231] = a[14] & g[20847];
assign g[53614] = b[14] & g[20847];
assign g[37232] = a[14] & g[20848];
assign g[53615] = b[14] & g[20848];
assign g[37233] = a[14] & g[20849];
assign g[53616] = b[14] & g[20849];
assign g[37234] = a[14] & g[20850];
assign g[53617] = b[14] & g[20850];
assign g[37235] = a[14] & g[20851];
assign g[53618] = b[14] & g[20851];
assign g[37236] = a[14] & g[20852];
assign g[53619] = b[14] & g[20852];
assign g[37237] = a[14] & g[20853];
assign g[53620] = b[14] & g[20853];
assign g[37238] = a[14] & g[20854];
assign g[53621] = b[14] & g[20854];
assign g[37239] = a[14] & g[20855];
assign g[53622] = b[14] & g[20855];
assign g[37240] = a[14] & g[20856];
assign g[53623] = b[14] & g[20856];
assign g[37241] = a[14] & g[20857];
assign g[53624] = b[14] & g[20857];
assign g[37242] = a[14] & g[20858];
assign g[53625] = b[14] & g[20858];
assign g[37243] = a[14] & g[20859];
assign g[53626] = b[14] & g[20859];
assign g[37244] = a[14] & g[20860];
assign g[53627] = b[14] & g[20860];
assign g[37245] = a[14] & g[20861];
assign g[53628] = b[14] & g[20861];
assign g[37246] = a[14] & g[20862];
assign g[53629] = b[14] & g[20862];
assign g[37247] = a[14] & g[20863];
assign g[53630] = b[14] & g[20863];
assign g[37248] = a[14] & g[20864];
assign g[53631] = b[14] & g[20864];
assign g[37249] = a[14] & g[20865];
assign g[53632] = b[14] & g[20865];
assign g[37250] = a[14] & g[20866];
assign g[53633] = b[14] & g[20866];
assign g[37251] = a[14] & g[20867];
assign g[53634] = b[14] & g[20867];
assign g[37252] = a[14] & g[20868];
assign g[53635] = b[14] & g[20868];
assign g[37253] = a[14] & g[20869];
assign g[53636] = b[14] & g[20869];
assign g[37254] = a[14] & g[20870];
assign g[53637] = b[14] & g[20870];
assign g[37255] = a[14] & g[20871];
assign g[53638] = b[14] & g[20871];
assign g[37256] = a[14] & g[20872];
assign g[53639] = b[14] & g[20872];
assign g[37257] = a[14] & g[20873];
assign g[53640] = b[14] & g[20873];
assign g[37258] = a[14] & g[20874];
assign g[53641] = b[14] & g[20874];
assign g[37259] = a[14] & g[20875];
assign g[53642] = b[14] & g[20875];
assign g[37260] = a[14] & g[20876];
assign g[53643] = b[14] & g[20876];
assign g[37261] = a[14] & g[20877];
assign g[53644] = b[14] & g[20877];
assign g[37262] = a[14] & g[20878];
assign g[53645] = b[14] & g[20878];
assign g[37263] = a[14] & g[20879];
assign g[53646] = b[14] & g[20879];
assign g[37264] = a[14] & g[20880];
assign g[53647] = b[14] & g[20880];
assign g[37265] = a[14] & g[20881];
assign g[53648] = b[14] & g[20881];
assign g[37266] = a[14] & g[20882];
assign g[53649] = b[14] & g[20882];
assign g[37267] = a[14] & g[20883];
assign g[53650] = b[14] & g[20883];
assign g[37268] = a[14] & g[20884];
assign g[53651] = b[14] & g[20884];
assign g[37269] = a[14] & g[20885];
assign g[53652] = b[14] & g[20885];
assign g[37270] = a[14] & g[20886];
assign g[53653] = b[14] & g[20886];
assign g[37271] = a[14] & g[20887];
assign g[53654] = b[14] & g[20887];
assign g[37272] = a[14] & g[20888];
assign g[53655] = b[14] & g[20888];
assign g[37273] = a[14] & g[20889];
assign g[53656] = b[14] & g[20889];
assign g[37274] = a[14] & g[20890];
assign g[53657] = b[14] & g[20890];
assign g[37275] = a[14] & g[20891];
assign g[53658] = b[14] & g[20891];
assign g[37276] = a[14] & g[20892];
assign g[53659] = b[14] & g[20892];
assign g[37277] = a[14] & g[20893];
assign g[53660] = b[14] & g[20893];
assign g[37278] = a[14] & g[20894];
assign g[53661] = b[14] & g[20894];
assign g[37279] = a[14] & g[20895];
assign g[53662] = b[14] & g[20895];
assign g[37280] = a[14] & g[20896];
assign g[53663] = b[14] & g[20896];
assign g[37281] = a[14] & g[20897];
assign g[53664] = b[14] & g[20897];
assign g[37282] = a[14] & g[20898];
assign g[53665] = b[14] & g[20898];
assign g[37283] = a[14] & g[20899];
assign g[53666] = b[14] & g[20899];
assign g[37284] = a[14] & g[20900];
assign g[53667] = b[14] & g[20900];
assign g[37285] = a[14] & g[20901];
assign g[53668] = b[14] & g[20901];
assign g[37286] = a[14] & g[20902];
assign g[53669] = b[14] & g[20902];
assign g[37287] = a[14] & g[20903];
assign g[53670] = b[14] & g[20903];
assign g[37288] = a[14] & g[20904];
assign g[53671] = b[14] & g[20904];
assign g[37289] = a[14] & g[20905];
assign g[53672] = b[14] & g[20905];
assign g[37290] = a[14] & g[20906];
assign g[53673] = b[14] & g[20906];
assign g[37291] = a[14] & g[20907];
assign g[53674] = b[14] & g[20907];
assign g[37292] = a[14] & g[20908];
assign g[53675] = b[14] & g[20908];
assign g[37293] = a[14] & g[20909];
assign g[53676] = b[14] & g[20909];
assign g[37294] = a[14] & g[20910];
assign g[53677] = b[14] & g[20910];
assign g[37295] = a[14] & g[20911];
assign g[53678] = b[14] & g[20911];
assign g[37296] = a[14] & g[20912];
assign g[53679] = b[14] & g[20912];
assign g[37297] = a[14] & g[20913];
assign g[53680] = b[14] & g[20913];
assign g[37298] = a[14] & g[20914];
assign g[53681] = b[14] & g[20914];
assign g[37299] = a[14] & g[20915];
assign g[53682] = b[14] & g[20915];
assign g[37300] = a[14] & g[20916];
assign g[53683] = b[14] & g[20916];
assign g[37301] = a[14] & g[20917];
assign g[53684] = b[14] & g[20917];
assign g[37302] = a[14] & g[20918];
assign g[53685] = b[14] & g[20918];
assign g[37303] = a[14] & g[20919];
assign g[53686] = b[14] & g[20919];
assign g[37304] = a[14] & g[20920];
assign g[53687] = b[14] & g[20920];
assign g[37305] = a[14] & g[20921];
assign g[53688] = b[14] & g[20921];
assign g[37306] = a[14] & g[20922];
assign g[53689] = b[14] & g[20922];
assign g[37307] = a[14] & g[20923];
assign g[53690] = b[14] & g[20923];
assign g[37308] = a[14] & g[20924];
assign g[53691] = b[14] & g[20924];
assign g[37309] = a[14] & g[20925];
assign g[53692] = b[14] & g[20925];
assign g[37310] = a[14] & g[20926];
assign g[53693] = b[14] & g[20926];
assign g[37311] = a[14] & g[20927];
assign g[53694] = b[14] & g[20927];
assign g[37312] = a[14] & g[20928];
assign g[53695] = b[14] & g[20928];
assign g[37313] = a[14] & g[20929];
assign g[53696] = b[14] & g[20929];
assign g[37314] = a[14] & g[20930];
assign g[53697] = b[14] & g[20930];
assign g[37315] = a[14] & g[20931];
assign g[53698] = b[14] & g[20931];
assign g[37316] = a[14] & g[20932];
assign g[53699] = b[14] & g[20932];
assign g[37317] = a[14] & g[20933];
assign g[53700] = b[14] & g[20933];
assign g[37318] = a[14] & g[20934];
assign g[53701] = b[14] & g[20934];
assign g[37319] = a[14] & g[20935];
assign g[53702] = b[14] & g[20935];
assign g[37320] = a[14] & g[20936];
assign g[53703] = b[14] & g[20936];
assign g[37321] = a[14] & g[20937];
assign g[53704] = b[14] & g[20937];
assign g[37322] = a[14] & g[20938];
assign g[53705] = b[14] & g[20938];
assign g[37323] = a[14] & g[20939];
assign g[53706] = b[14] & g[20939];
assign g[37324] = a[14] & g[20940];
assign g[53707] = b[14] & g[20940];
assign g[37325] = a[14] & g[20941];
assign g[53708] = b[14] & g[20941];
assign g[37326] = a[14] & g[20942];
assign g[53709] = b[14] & g[20942];
assign g[37327] = a[14] & g[20943];
assign g[53710] = b[14] & g[20943];
assign g[37328] = a[14] & g[20944];
assign g[53711] = b[14] & g[20944];
assign g[37329] = a[14] & g[20945];
assign g[53712] = b[14] & g[20945];
assign g[37330] = a[14] & g[20946];
assign g[53713] = b[14] & g[20946];
assign g[37331] = a[14] & g[20947];
assign g[53714] = b[14] & g[20947];
assign g[37332] = a[14] & g[20948];
assign g[53715] = b[14] & g[20948];
assign g[37333] = a[14] & g[20949];
assign g[53716] = b[14] & g[20949];
assign g[37334] = a[14] & g[20950];
assign g[53717] = b[14] & g[20950];
assign g[37335] = a[14] & g[20951];
assign g[53718] = b[14] & g[20951];
assign g[37336] = a[14] & g[20952];
assign g[53719] = b[14] & g[20952];
assign g[37337] = a[14] & g[20953];
assign g[53720] = b[14] & g[20953];
assign g[37338] = a[14] & g[20954];
assign g[53721] = b[14] & g[20954];
assign g[37339] = a[14] & g[20955];
assign g[53722] = b[14] & g[20955];
assign g[37340] = a[14] & g[20956];
assign g[53723] = b[14] & g[20956];
assign g[37341] = a[14] & g[20957];
assign g[53724] = b[14] & g[20957];
assign g[37342] = a[14] & g[20958];
assign g[53725] = b[14] & g[20958];
assign g[37343] = a[14] & g[20959];
assign g[53726] = b[14] & g[20959];
assign g[37344] = a[14] & g[20960];
assign g[53727] = b[14] & g[20960];
assign g[37345] = a[14] & g[20961];
assign g[53728] = b[14] & g[20961];
assign g[37346] = a[14] & g[20962];
assign g[53729] = b[14] & g[20962];
assign g[37347] = a[14] & g[20963];
assign g[53730] = b[14] & g[20963];
assign g[37348] = a[14] & g[20964];
assign g[53731] = b[14] & g[20964];
assign g[37349] = a[14] & g[20965];
assign g[53732] = b[14] & g[20965];
assign g[37350] = a[14] & g[20966];
assign g[53733] = b[14] & g[20966];
assign g[37351] = a[14] & g[20967];
assign g[53734] = b[14] & g[20967];
assign g[37352] = a[14] & g[20968];
assign g[53735] = b[14] & g[20968];
assign g[37353] = a[14] & g[20969];
assign g[53736] = b[14] & g[20969];
assign g[37354] = a[14] & g[20970];
assign g[53737] = b[14] & g[20970];
assign g[37355] = a[14] & g[20971];
assign g[53738] = b[14] & g[20971];
assign g[37356] = a[14] & g[20972];
assign g[53739] = b[14] & g[20972];
assign g[37357] = a[14] & g[20973];
assign g[53740] = b[14] & g[20973];
assign g[37358] = a[14] & g[20974];
assign g[53741] = b[14] & g[20974];
assign g[37359] = a[14] & g[20975];
assign g[53742] = b[14] & g[20975];
assign g[37360] = a[14] & g[20976];
assign g[53743] = b[14] & g[20976];
assign g[37361] = a[14] & g[20977];
assign g[53744] = b[14] & g[20977];
assign g[37362] = a[14] & g[20978];
assign g[53745] = b[14] & g[20978];
assign g[37363] = a[14] & g[20979];
assign g[53746] = b[14] & g[20979];
assign g[37364] = a[14] & g[20980];
assign g[53747] = b[14] & g[20980];
assign g[37365] = a[14] & g[20981];
assign g[53748] = b[14] & g[20981];
assign g[37366] = a[14] & g[20982];
assign g[53749] = b[14] & g[20982];
assign g[37367] = a[14] & g[20983];
assign g[53750] = b[14] & g[20983];
assign g[37368] = a[14] & g[20984];
assign g[53751] = b[14] & g[20984];
assign g[37369] = a[14] & g[20985];
assign g[53752] = b[14] & g[20985];
assign g[37370] = a[14] & g[20986];
assign g[53753] = b[14] & g[20986];
assign g[37371] = a[14] & g[20987];
assign g[53754] = b[14] & g[20987];
assign g[37372] = a[14] & g[20988];
assign g[53755] = b[14] & g[20988];
assign g[37373] = a[14] & g[20989];
assign g[53756] = b[14] & g[20989];
assign g[37374] = a[14] & g[20990];
assign g[53757] = b[14] & g[20990];
assign g[37375] = a[14] & g[20991];
assign g[53758] = b[14] & g[20991];
assign g[37376] = a[14] & g[20992];
assign g[53759] = b[14] & g[20992];
assign g[37377] = a[14] & g[20993];
assign g[53760] = b[14] & g[20993];
assign g[37378] = a[14] & g[20994];
assign g[53761] = b[14] & g[20994];
assign g[37379] = a[14] & g[20995];
assign g[53762] = b[14] & g[20995];
assign g[37380] = a[14] & g[20996];
assign g[53763] = b[14] & g[20996];
assign g[37381] = a[14] & g[20997];
assign g[53764] = b[14] & g[20997];
assign g[37382] = a[14] & g[20998];
assign g[53765] = b[14] & g[20998];
assign g[37383] = a[14] & g[20999];
assign g[53766] = b[14] & g[20999];
assign g[37384] = a[14] & g[21000];
assign g[53767] = b[14] & g[21000];
assign g[37385] = a[14] & g[21001];
assign g[53768] = b[14] & g[21001];
assign g[37386] = a[14] & g[21002];
assign g[53769] = b[14] & g[21002];
assign g[37387] = a[14] & g[21003];
assign g[53770] = b[14] & g[21003];
assign g[37388] = a[14] & g[21004];
assign g[53771] = b[14] & g[21004];
assign g[37389] = a[14] & g[21005];
assign g[53772] = b[14] & g[21005];
assign g[37390] = a[14] & g[21006];
assign g[53773] = b[14] & g[21006];
assign g[37391] = a[14] & g[21007];
assign g[53774] = b[14] & g[21007];
assign g[37392] = a[14] & g[21008];
assign g[53775] = b[14] & g[21008];
assign g[37393] = a[14] & g[21009];
assign g[53776] = b[14] & g[21009];
assign g[37394] = a[14] & g[21010];
assign g[53777] = b[14] & g[21010];
assign g[37395] = a[14] & g[21011];
assign g[53778] = b[14] & g[21011];
assign g[37396] = a[14] & g[21012];
assign g[53779] = b[14] & g[21012];
assign g[37397] = a[14] & g[21013];
assign g[53780] = b[14] & g[21013];
assign g[37398] = a[14] & g[21014];
assign g[53781] = b[14] & g[21014];
assign g[37399] = a[14] & g[21015];
assign g[53782] = b[14] & g[21015];
assign g[37400] = a[14] & g[21016];
assign g[53783] = b[14] & g[21016];
assign g[37401] = a[14] & g[21017];
assign g[53784] = b[14] & g[21017];
assign g[37402] = a[14] & g[21018];
assign g[53785] = b[14] & g[21018];
assign g[37403] = a[14] & g[21019];
assign g[53786] = b[14] & g[21019];
assign g[37404] = a[14] & g[21020];
assign g[53787] = b[14] & g[21020];
assign g[37405] = a[14] & g[21021];
assign g[53788] = b[14] & g[21021];
assign g[37406] = a[14] & g[21022];
assign g[53789] = b[14] & g[21022];
assign g[37407] = a[14] & g[21023];
assign g[53790] = b[14] & g[21023];
assign g[37408] = a[14] & g[21024];
assign g[53791] = b[14] & g[21024];
assign g[37409] = a[14] & g[21025];
assign g[53792] = b[14] & g[21025];
assign g[37410] = a[14] & g[21026];
assign g[53793] = b[14] & g[21026];
assign g[37411] = a[14] & g[21027];
assign g[53794] = b[14] & g[21027];
assign g[37412] = a[14] & g[21028];
assign g[53795] = b[14] & g[21028];
assign g[37413] = a[14] & g[21029];
assign g[53796] = b[14] & g[21029];
assign g[37414] = a[14] & g[21030];
assign g[53797] = b[14] & g[21030];
assign g[37415] = a[14] & g[21031];
assign g[53798] = b[14] & g[21031];
assign g[37416] = a[14] & g[21032];
assign g[53799] = b[14] & g[21032];
assign g[37417] = a[14] & g[21033];
assign g[53800] = b[14] & g[21033];
assign g[37418] = a[14] & g[21034];
assign g[53801] = b[14] & g[21034];
assign g[37419] = a[14] & g[21035];
assign g[53802] = b[14] & g[21035];
assign g[37420] = a[14] & g[21036];
assign g[53803] = b[14] & g[21036];
assign g[37421] = a[14] & g[21037];
assign g[53804] = b[14] & g[21037];
assign g[37422] = a[14] & g[21038];
assign g[53805] = b[14] & g[21038];
assign g[37423] = a[14] & g[21039];
assign g[53806] = b[14] & g[21039];
assign g[37424] = a[14] & g[21040];
assign g[53807] = b[14] & g[21040];
assign g[37425] = a[14] & g[21041];
assign g[53808] = b[14] & g[21041];
assign g[37426] = a[14] & g[21042];
assign g[53809] = b[14] & g[21042];
assign g[37427] = a[14] & g[21043];
assign g[53810] = b[14] & g[21043];
assign g[37428] = a[14] & g[21044];
assign g[53811] = b[14] & g[21044];
assign g[37429] = a[14] & g[21045];
assign g[53812] = b[14] & g[21045];
assign g[37430] = a[14] & g[21046];
assign g[53813] = b[14] & g[21046];
assign g[37431] = a[14] & g[21047];
assign g[53814] = b[14] & g[21047];
assign g[37432] = a[14] & g[21048];
assign g[53815] = b[14] & g[21048];
assign g[37433] = a[14] & g[21049];
assign g[53816] = b[14] & g[21049];
assign g[37434] = a[14] & g[21050];
assign g[53817] = b[14] & g[21050];
assign g[37435] = a[14] & g[21051];
assign g[53818] = b[14] & g[21051];
assign g[37436] = a[14] & g[21052];
assign g[53819] = b[14] & g[21052];
assign g[37437] = a[14] & g[21053];
assign g[53820] = b[14] & g[21053];
assign g[37438] = a[14] & g[21054];
assign g[53821] = b[14] & g[21054];
assign g[37439] = a[14] & g[21055];
assign g[53822] = b[14] & g[21055];
assign g[37440] = a[14] & g[21056];
assign g[53823] = b[14] & g[21056];
assign g[37441] = a[14] & g[21057];
assign g[53824] = b[14] & g[21057];
assign g[37442] = a[14] & g[21058];
assign g[53825] = b[14] & g[21058];
assign g[37443] = a[14] & g[21059];
assign g[53826] = b[14] & g[21059];
assign g[37444] = a[14] & g[21060];
assign g[53827] = b[14] & g[21060];
assign g[37445] = a[14] & g[21061];
assign g[53828] = b[14] & g[21061];
assign g[37446] = a[14] & g[21062];
assign g[53829] = b[14] & g[21062];
assign g[37447] = a[14] & g[21063];
assign g[53830] = b[14] & g[21063];
assign g[37448] = a[14] & g[21064];
assign g[53831] = b[14] & g[21064];
assign g[37449] = a[14] & g[21065];
assign g[53832] = b[14] & g[21065];
assign g[37450] = a[14] & g[21066];
assign g[53833] = b[14] & g[21066];
assign g[37451] = a[14] & g[21067];
assign g[53834] = b[14] & g[21067];
assign g[37452] = a[14] & g[21068];
assign g[53835] = b[14] & g[21068];
assign g[37453] = a[14] & g[21069];
assign g[53836] = b[14] & g[21069];
assign g[37454] = a[14] & g[21070];
assign g[53837] = b[14] & g[21070];
assign g[37455] = a[14] & g[21071];
assign g[53838] = b[14] & g[21071];
assign g[37456] = a[14] & g[21072];
assign g[53839] = b[14] & g[21072];
assign g[37457] = a[14] & g[21073];
assign g[53840] = b[14] & g[21073];
assign g[37458] = a[14] & g[21074];
assign g[53841] = b[14] & g[21074];
assign g[37459] = a[14] & g[21075];
assign g[53842] = b[14] & g[21075];
assign g[37460] = a[14] & g[21076];
assign g[53843] = b[14] & g[21076];
assign g[37461] = a[14] & g[21077];
assign g[53844] = b[14] & g[21077];
assign g[37462] = a[14] & g[21078];
assign g[53845] = b[14] & g[21078];
assign g[37463] = a[14] & g[21079];
assign g[53846] = b[14] & g[21079];
assign g[37464] = a[14] & g[21080];
assign g[53847] = b[14] & g[21080];
assign g[37465] = a[14] & g[21081];
assign g[53848] = b[14] & g[21081];
assign g[37466] = a[14] & g[21082];
assign g[53849] = b[14] & g[21082];
assign g[37467] = a[14] & g[21083];
assign g[53850] = b[14] & g[21083];
assign g[37468] = a[14] & g[21084];
assign g[53851] = b[14] & g[21084];
assign g[37469] = a[14] & g[21085];
assign g[53852] = b[14] & g[21085];
assign g[37470] = a[14] & g[21086];
assign g[53853] = b[14] & g[21086];
assign g[37471] = a[14] & g[21087];
assign g[53854] = b[14] & g[21087];
assign g[37472] = a[14] & g[21088];
assign g[53855] = b[14] & g[21088];
assign g[37473] = a[14] & g[21089];
assign g[53856] = b[14] & g[21089];
assign g[37474] = a[14] & g[21090];
assign g[53857] = b[14] & g[21090];
assign g[37475] = a[14] & g[21091];
assign g[53858] = b[14] & g[21091];
assign g[37476] = a[14] & g[21092];
assign g[53859] = b[14] & g[21092];
assign g[37477] = a[14] & g[21093];
assign g[53860] = b[14] & g[21093];
assign g[37478] = a[14] & g[21094];
assign g[53861] = b[14] & g[21094];
assign g[37479] = a[14] & g[21095];
assign g[53862] = b[14] & g[21095];
assign g[37480] = a[14] & g[21096];
assign g[53863] = b[14] & g[21096];
assign g[37481] = a[14] & g[21097];
assign g[53864] = b[14] & g[21097];
assign g[37482] = a[14] & g[21098];
assign g[53865] = b[14] & g[21098];
assign g[37483] = a[14] & g[21099];
assign g[53866] = b[14] & g[21099];
assign g[37484] = a[14] & g[21100];
assign g[53867] = b[14] & g[21100];
assign g[37485] = a[14] & g[21101];
assign g[53868] = b[14] & g[21101];
assign g[37486] = a[14] & g[21102];
assign g[53869] = b[14] & g[21102];
assign g[37487] = a[14] & g[21103];
assign g[53870] = b[14] & g[21103];
assign g[37488] = a[14] & g[21104];
assign g[53871] = b[14] & g[21104];
assign g[37489] = a[14] & g[21105];
assign g[53872] = b[14] & g[21105];
assign g[37490] = a[14] & g[21106];
assign g[53873] = b[14] & g[21106];
assign g[37491] = a[14] & g[21107];
assign g[53874] = b[14] & g[21107];
assign g[37492] = a[14] & g[21108];
assign g[53875] = b[14] & g[21108];
assign g[37493] = a[14] & g[21109];
assign g[53876] = b[14] & g[21109];
assign g[37494] = a[14] & g[21110];
assign g[53877] = b[14] & g[21110];
assign g[37495] = a[14] & g[21111];
assign g[53878] = b[14] & g[21111];
assign g[37496] = a[14] & g[21112];
assign g[53879] = b[14] & g[21112];
assign g[37497] = a[14] & g[21113];
assign g[53880] = b[14] & g[21113];
assign g[37498] = a[14] & g[21114];
assign g[53881] = b[14] & g[21114];
assign g[37499] = a[14] & g[21115];
assign g[53882] = b[14] & g[21115];
assign g[37500] = a[14] & g[21116];
assign g[53883] = b[14] & g[21116];
assign g[37501] = a[14] & g[21117];
assign g[53884] = b[14] & g[21117];
assign g[37502] = a[14] & g[21118];
assign g[53885] = b[14] & g[21118];
assign g[37503] = a[14] & g[21119];
assign g[53886] = b[14] & g[21119];
assign g[37504] = a[14] & g[21120];
assign g[53887] = b[14] & g[21120];
assign g[37505] = a[14] & g[21121];
assign g[53888] = b[14] & g[21121];
assign g[37506] = a[14] & g[21122];
assign g[53889] = b[14] & g[21122];
assign g[37507] = a[14] & g[21123];
assign g[53890] = b[14] & g[21123];
assign g[37508] = a[14] & g[21124];
assign g[53891] = b[14] & g[21124];
assign g[37509] = a[14] & g[21125];
assign g[53892] = b[14] & g[21125];
assign g[37510] = a[14] & g[21126];
assign g[53893] = b[14] & g[21126];
assign g[37511] = a[14] & g[21127];
assign g[53894] = b[14] & g[21127];
assign g[37512] = a[14] & g[21128];
assign g[53895] = b[14] & g[21128];
assign g[37513] = a[14] & g[21129];
assign g[53896] = b[14] & g[21129];
assign g[37514] = a[14] & g[21130];
assign g[53897] = b[14] & g[21130];
assign g[37515] = a[14] & g[21131];
assign g[53898] = b[14] & g[21131];
assign g[37516] = a[14] & g[21132];
assign g[53899] = b[14] & g[21132];
assign g[37517] = a[14] & g[21133];
assign g[53900] = b[14] & g[21133];
assign g[37518] = a[14] & g[21134];
assign g[53901] = b[14] & g[21134];
assign g[37519] = a[14] & g[21135];
assign g[53902] = b[14] & g[21135];
assign g[37520] = a[14] & g[21136];
assign g[53903] = b[14] & g[21136];
assign g[37521] = a[14] & g[21137];
assign g[53904] = b[14] & g[21137];
assign g[37522] = a[14] & g[21138];
assign g[53905] = b[14] & g[21138];
assign g[37523] = a[14] & g[21139];
assign g[53906] = b[14] & g[21139];
assign g[37524] = a[14] & g[21140];
assign g[53907] = b[14] & g[21140];
assign g[37525] = a[14] & g[21141];
assign g[53908] = b[14] & g[21141];
assign g[37526] = a[14] & g[21142];
assign g[53909] = b[14] & g[21142];
assign g[37527] = a[14] & g[21143];
assign g[53910] = b[14] & g[21143];
assign g[37528] = a[14] & g[21144];
assign g[53911] = b[14] & g[21144];
assign g[37529] = a[14] & g[21145];
assign g[53912] = b[14] & g[21145];
assign g[37530] = a[14] & g[21146];
assign g[53913] = b[14] & g[21146];
assign g[37531] = a[14] & g[21147];
assign g[53914] = b[14] & g[21147];
assign g[37532] = a[14] & g[21148];
assign g[53915] = b[14] & g[21148];
assign g[37533] = a[14] & g[21149];
assign g[53916] = b[14] & g[21149];
assign g[37534] = a[14] & g[21150];
assign g[53917] = b[14] & g[21150];
assign g[37535] = a[14] & g[21151];
assign g[53918] = b[14] & g[21151];
assign g[37536] = a[14] & g[21152];
assign g[53919] = b[14] & g[21152];
assign g[37537] = a[14] & g[21153];
assign g[53920] = b[14] & g[21153];
assign g[37538] = a[14] & g[21154];
assign g[53921] = b[14] & g[21154];
assign g[37539] = a[14] & g[21155];
assign g[53922] = b[14] & g[21155];
assign g[37540] = a[14] & g[21156];
assign g[53923] = b[14] & g[21156];
assign g[37541] = a[14] & g[21157];
assign g[53924] = b[14] & g[21157];
assign g[37542] = a[14] & g[21158];
assign g[53925] = b[14] & g[21158];
assign g[37543] = a[14] & g[21159];
assign g[53926] = b[14] & g[21159];
assign g[37544] = a[14] & g[21160];
assign g[53927] = b[14] & g[21160];
assign g[37545] = a[14] & g[21161];
assign g[53928] = b[14] & g[21161];
assign g[37546] = a[14] & g[21162];
assign g[53929] = b[14] & g[21162];
assign g[37547] = a[14] & g[21163];
assign g[53930] = b[14] & g[21163];
assign g[37548] = a[14] & g[21164];
assign g[53931] = b[14] & g[21164];
assign g[37549] = a[14] & g[21165];
assign g[53932] = b[14] & g[21165];
assign g[37550] = a[14] & g[21166];
assign g[53933] = b[14] & g[21166];
assign g[37551] = a[14] & g[21167];
assign g[53934] = b[14] & g[21167];
assign g[37552] = a[14] & g[21168];
assign g[53935] = b[14] & g[21168];
assign g[37553] = a[14] & g[21169];
assign g[53936] = b[14] & g[21169];
assign g[37554] = a[14] & g[21170];
assign g[53937] = b[14] & g[21170];
assign g[37555] = a[14] & g[21171];
assign g[53938] = b[14] & g[21171];
assign g[37556] = a[14] & g[21172];
assign g[53939] = b[14] & g[21172];
assign g[37557] = a[14] & g[21173];
assign g[53940] = b[14] & g[21173];
assign g[37558] = a[14] & g[21174];
assign g[53941] = b[14] & g[21174];
assign g[37559] = a[14] & g[21175];
assign g[53942] = b[14] & g[21175];
assign g[37560] = a[14] & g[21176];
assign g[53943] = b[14] & g[21176];
assign g[37561] = a[14] & g[21177];
assign g[53944] = b[14] & g[21177];
assign g[37562] = a[14] & g[21178];
assign g[53945] = b[14] & g[21178];
assign g[37563] = a[14] & g[21179];
assign g[53946] = b[14] & g[21179];
assign g[37564] = a[14] & g[21180];
assign g[53947] = b[14] & g[21180];
assign g[37565] = a[14] & g[21181];
assign g[53948] = b[14] & g[21181];
assign g[37566] = a[14] & g[21182];
assign g[53949] = b[14] & g[21182];
assign g[37567] = a[14] & g[21183];
assign g[53950] = b[14] & g[21183];
assign g[37568] = a[14] & g[21184];
assign g[53951] = b[14] & g[21184];
assign g[37569] = a[14] & g[21185];
assign g[53952] = b[14] & g[21185];
assign g[37570] = a[14] & g[21186];
assign g[53953] = b[14] & g[21186];
assign g[37571] = a[14] & g[21187];
assign g[53954] = b[14] & g[21187];
assign g[37572] = a[14] & g[21188];
assign g[53955] = b[14] & g[21188];
assign g[37573] = a[14] & g[21189];
assign g[53956] = b[14] & g[21189];
assign g[37574] = a[14] & g[21190];
assign g[53957] = b[14] & g[21190];
assign g[37575] = a[14] & g[21191];
assign g[53958] = b[14] & g[21191];
assign g[37576] = a[14] & g[21192];
assign g[53959] = b[14] & g[21192];
assign g[37577] = a[14] & g[21193];
assign g[53960] = b[14] & g[21193];
assign g[37578] = a[14] & g[21194];
assign g[53961] = b[14] & g[21194];
assign g[37579] = a[14] & g[21195];
assign g[53962] = b[14] & g[21195];
assign g[37580] = a[14] & g[21196];
assign g[53963] = b[14] & g[21196];
assign g[37581] = a[14] & g[21197];
assign g[53964] = b[14] & g[21197];
assign g[37582] = a[14] & g[21198];
assign g[53965] = b[14] & g[21198];
assign g[37583] = a[14] & g[21199];
assign g[53966] = b[14] & g[21199];
assign g[37584] = a[14] & g[21200];
assign g[53967] = b[14] & g[21200];
assign g[37585] = a[14] & g[21201];
assign g[53968] = b[14] & g[21201];
assign g[37586] = a[14] & g[21202];
assign g[53969] = b[14] & g[21202];
assign g[37587] = a[14] & g[21203];
assign g[53970] = b[14] & g[21203];
assign g[37588] = a[14] & g[21204];
assign g[53971] = b[14] & g[21204];
assign g[37589] = a[14] & g[21205];
assign g[53972] = b[14] & g[21205];
assign g[37590] = a[14] & g[21206];
assign g[53973] = b[14] & g[21206];
assign g[37591] = a[14] & g[21207];
assign g[53974] = b[14] & g[21207];
assign g[37592] = a[14] & g[21208];
assign g[53975] = b[14] & g[21208];
assign g[37593] = a[14] & g[21209];
assign g[53976] = b[14] & g[21209];
assign g[37594] = a[14] & g[21210];
assign g[53977] = b[14] & g[21210];
assign g[37595] = a[14] & g[21211];
assign g[53978] = b[14] & g[21211];
assign g[37596] = a[14] & g[21212];
assign g[53979] = b[14] & g[21212];
assign g[37597] = a[14] & g[21213];
assign g[53980] = b[14] & g[21213];
assign g[37598] = a[14] & g[21214];
assign g[53981] = b[14] & g[21214];
assign g[37599] = a[14] & g[21215];
assign g[53982] = b[14] & g[21215];
assign g[37600] = a[14] & g[21216];
assign g[53983] = b[14] & g[21216];
assign g[37601] = a[14] & g[21217];
assign g[53984] = b[14] & g[21217];
assign g[37602] = a[14] & g[21218];
assign g[53985] = b[14] & g[21218];
assign g[37603] = a[14] & g[21219];
assign g[53986] = b[14] & g[21219];
assign g[37604] = a[14] & g[21220];
assign g[53987] = b[14] & g[21220];
assign g[37605] = a[14] & g[21221];
assign g[53988] = b[14] & g[21221];
assign g[37606] = a[14] & g[21222];
assign g[53989] = b[14] & g[21222];
assign g[37607] = a[14] & g[21223];
assign g[53990] = b[14] & g[21223];
assign g[37608] = a[14] & g[21224];
assign g[53991] = b[14] & g[21224];
assign g[37609] = a[14] & g[21225];
assign g[53992] = b[14] & g[21225];
assign g[37610] = a[14] & g[21226];
assign g[53993] = b[14] & g[21226];
assign g[37611] = a[14] & g[21227];
assign g[53994] = b[14] & g[21227];
assign g[37612] = a[14] & g[21228];
assign g[53995] = b[14] & g[21228];
assign g[37613] = a[14] & g[21229];
assign g[53996] = b[14] & g[21229];
assign g[37614] = a[14] & g[21230];
assign g[53997] = b[14] & g[21230];
assign g[37615] = a[14] & g[21231];
assign g[53998] = b[14] & g[21231];
assign g[37616] = a[14] & g[21232];
assign g[53999] = b[14] & g[21232];
assign g[37617] = a[14] & g[21233];
assign g[54000] = b[14] & g[21233];
assign g[37618] = a[14] & g[21234];
assign g[54001] = b[14] & g[21234];
assign g[37619] = a[14] & g[21235];
assign g[54002] = b[14] & g[21235];
assign g[37620] = a[14] & g[21236];
assign g[54003] = b[14] & g[21236];
assign g[37621] = a[14] & g[21237];
assign g[54004] = b[14] & g[21237];
assign g[37622] = a[14] & g[21238];
assign g[54005] = b[14] & g[21238];
assign g[37623] = a[14] & g[21239];
assign g[54006] = b[14] & g[21239];
assign g[37624] = a[14] & g[21240];
assign g[54007] = b[14] & g[21240];
assign g[37625] = a[14] & g[21241];
assign g[54008] = b[14] & g[21241];
assign g[37626] = a[14] & g[21242];
assign g[54009] = b[14] & g[21242];
assign g[37627] = a[14] & g[21243];
assign g[54010] = b[14] & g[21243];
assign g[37628] = a[14] & g[21244];
assign g[54011] = b[14] & g[21244];
assign g[37629] = a[14] & g[21245];
assign g[54012] = b[14] & g[21245];
assign g[37630] = a[14] & g[21246];
assign g[54013] = b[14] & g[21246];
assign g[37631] = a[14] & g[21247];
assign g[54014] = b[14] & g[21247];
assign g[37632] = a[14] & g[21248];
assign g[54015] = b[14] & g[21248];
assign g[37633] = a[14] & g[21249];
assign g[54016] = b[14] & g[21249];
assign g[37634] = a[14] & g[21250];
assign g[54017] = b[14] & g[21250];
assign g[37635] = a[14] & g[21251];
assign g[54018] = b[14] & g[21251];
assign g[37636] = a[14] & g[21252];
assign g[54019] = b[14] & g[21252];
assign g[37637] = a[14] & g[21253];
assign g[54020] = b[14] & g[21253];
assign g[37638] = a[14] & g[21254];
assign g[54021] = b[14] & g[21254];
assign g[37639] = a[14] & g[21255];
assign g[54022] = b[14] & g[21255];
assign g[37640] = a[14] & g[21256];
assign g[54023] = b[14] & g[21256];
assign g[37641] = a[14] & g[21257];
assign g[54024] = b[14] & g[21257];
assign g[37642] = a[14] & g[21258];
assign g[54025] = b[14] & g[21258];
assign g[37643] = a[14] & g[21259];
assign g[54026] = b[14] & g[21259];
assign g[37644] = a[14] & g[21260];
assign g[54027] = b[14] & g[21260];
assign g[37645] = a[14] & g[21261];
assign g[54028] = b[14] & g[21261];
assign g[37646] = a[14] & g[21262];
assign g[54029] = b[14] & g[21262];
assign g[37647] = a[14] & g[21263];
assign g[54030] = b[14] & g[21263];
assign g[37648] = a[14] & g[21264];
assign g[54031] = b[14] & g[21264];
assign g[37649] = a[14] & g[21265];
assign g[54032] = b[14] & g[21265];
assign g[37650] = a[14] & g[21266];
assign g[54033] = b[14] & g[21266];
assign g[37651] = a[14] & g[21267];
assign g[54034] = b[14] & g[21267];
assign g[37652] = a[14] & g[21268];
assign g[54035] = b[14] & g[21268];
assign g[37653] = a[14] & g[21269];
assign g[54036] = b[14] & g[21269];
assign g[37654] = a[14] & g[21270];
assign g[54037] = b[14] & g[21270];
assign g[37655] = a[14] & g[21271];
assign g[54038] = b[14] & g[21271];
assign g[37656] = a[14] & g[21272];
assign g[54039] = b[14] & g[21272];
assign g[37657] = a[14] & g[21273];
assign g[54040] = b[14] & g[21273];
assign g[37658] = a[14] & g[21274];
assign g[54041] = b[14] & g[21274];
assign g[37659] = a[14] & g[21275];
assign g[54042] = b[14] & g[21275];
assign g[37660] = a[14] & g[21276];
assign g[54043] = b[14] & g[21276];
assign g[37661] = a[14] & g[21277];
assign g[54044] = b[14] & g[21277];
assign g[37662] = a[14] & g[21278];
assign g[54045] = b[14] & g[21278];
assign g[37663] = a[14] & g[21279];
assign g[54046] = b[14] & g[21279];
assign g[37664] = a[14] & g[21280];
assign g[54047] = b[14] & g[21280];
assign g[37665] = a[14] & g[21281];
assign g[54048] = b[14] & g[21281];
assign g[37666] = a[14] & g[21282];
assign g[54049] = b[14] & g[21282];
assign g[37667] = a[14] & g[21283];
assign g[54050] = b[14] & g[21283];
assign g[37668] = a[14] & g[21284];
assign g[54051] = b[14] & g[21284];
assign g[37669] = a[14] & g[21285];
assign g[54052] = b[14] & g[21285];
assign g[37670] = a[14] & g[21286];
assign g[54053] = b[14] & g[21286];
assign g[37671] = a[14] & g[21287];
assign g[54054] = b[14] & g[21287];
assign g[37672] = a[14] & g[21288];
assign g[54055] = b[14] & g[21288];
assign g[37673] = a[14] & g[21289];
assign g[54056] = b[14] & g[21289];
assign g[37674] = a[14] & g[21290];
assign g[54057] = b[14] & g[21290];
assign g[37675] = a[14] & g[21291];
assign g[54058] = b[14] & g[21291];
assign g[37676] = a[14] & g[21292];
assign g[54059] = b[14] & g[21292];
assign g[37677] = a[14] & g[21293];
assign g[54060] = b[14] & g[21293];
assign g[37678] = a[14] & g[21294];
assign g[54061] = b[14] & g[21294];
assign g[37679] = a[14] & g[21295];
assign g[54062] = b[14] & g[21295];
assign g[37680] = a[14] & g[21296];
assign g[54063] = b[14] & g[21296];
assign g[37681] = a[14] & g[21297];
assign g[54064] = b[14] & g[21297];
assign g[37682] = a[14] & g[21298];
assign g[54065] = b[14] & g[21298];
assign g[37683] = a[14] & g[21299];
assign g[54066] = b[14] & g[21299];
assign g[37684] = a[14] & g[21300];
assign g[54067] = b[14] & g[21300];
assign g[37685] = a[14] & g[21301];
assign g[54068] = b[14] & g[21301];
assign g[37686] = a[14] & g[21302];
assign g[54069] = b[14] & g[21302];
assign g[37687] = a[14] & g[21303];
assign g[54070] = b[14] & g[21303];
assign g[37688] = a[14] & g[21304];
assign g[54071] = b[14] & g[21304];
assign g[37689] = a[14] & g[21305];
assign g[54072] = b[14] & g[21305];
assign g[37690] = a[14] & g[21306];
assign g[54073] = b[14] & g[21306];
assign g[37691] = a[14] & g[21307];
assign g[54074] = b[14] & g[21307];
assign g[37692] = a[14] & g[21308];
assign g[54075] = b[14] & g[21308];
assign g[37693] = a[14] & g[21309];
assign g[54076] = b[14] & g[21309];
assign g[37694] = a[14] & g[21310];
assign g[54077] = b[14] & g[21310];
assign g[37695] = a[14] & g[21311];
assign g[54078] = b[14] & g[21311];
assign g[37696] = a[14] & g[21312];
assign g[54079] = b[14] & g[21312];
assign g[37697] = a[14] & g[21313];
assign g[54080] = b[14] & g[21313];
assign g[37698] = a[14] & g[21314];
assign g[54081] = b[14] & g[21314];
assign g[37699] = a[14] & g[21315];
assign g[54082] = b[14] & g[21315];
assign g[37700] = a[14] & g[21316];
assign g[54083] = b[14] & g[21316];
assign g[37701] = a[14] & g[21317];
assign g[54084] = b[14] & g[21317];
assign g[37702] = a[14] & g[21318];
assign g[54085] = b[14] & g[21318];
assign g[37703] = a[14] & g[21319];
assign g[54086] = b[14] & g[21319];
assign g[37704] = a[14] & g[21320];
assign g[54087] = b[14] & g[21320];
assign g[37705] = a[14] & g[21321];
assign g[54088] = b[14] & g[21321];
assign g[37706] = a[14] & g[21322];
assign g[54089] = b[14] & g[21322];
assign g[37707] = a[14] & g[21323];
assign g[54090] = b[14] & g[21323];
assign g[37708] = a[14] & g[21324];
assign g[54091] = b[14] & g[21324];
assign g[37709] = a[14] & g[21325];
assign g[54092] = b[14] & g[21325];
assign g[37710] = a[14] & g[21326];
assign g[54093] = b[14] & g[21326];
assign g[37711] = a[14] & g[21327];
assign g[54094] = b[14] & g[21327];
assign g[37712] = a[14] & g[21328];
assign g[54095] = b[14] & g[21328];
assign g[37713] = a[14] & g[21329];
assign g[54096] = b[14] & g[21329];
assign g[37714] = a[14] & g[21330];
assign g[54097] = b[14] & g[21330];
assign g[37715] = a[14] & g[21331];
assign g[54098] = b[14] & g[21331];
assign g[37716] = a[14] & g[21332];
assign g[54099] = b[14] & g[21332];
assign g[37717] = a[14] & g[21333];
assign g[54100] = b[14] & g[21333];
assign g[37718] = a[14] & g[21334];
assign g[54101] = b[14] & g[21334];
assign g[37719] = a[14] & g[21335];
assign g[54102] = b[14] & g[21335];
assign g[37720] = a[14] & g[21336];
assign g[54103] = b[14] & g[21336];
assign g[37721] = a[14] & g[21337];
assign g[54104] = b[14] & g[21337];
assign g[37722] = a[14] & g[21338];
assign g[54105] = b[14] & g[21338];
assign g[37723] = a[14] & g[21339];
assign g[54106] = b[14] & g[21339];
assign g[37724] = a[14] & g[21340];
assign g[54107] = b[14] & g[21340];
assign g[37725] = a[14] & g[21341];
assign g[54108] = b[14] & g[21341];
assign g[37726] = a[14] & g[21342];
assign g[54109] = b[14] & g[21342];
assign g[37727] = a[14] & g[21343];
assign g[54110] = b[14] & g[21343];
assign g[37728] = a[14] & g[21344];
assign g[54111] = b[14] & g[21344];
assign g[37729] = a[14] & g[21345];
assign g[54112] = b[14] & g[21345];
assign g[37730] = a[14] & g[21346];
assign g[54113] = b[14] & g[21346];
assign g[37731] = a[14] & g[21347];
assign g[54114] = b[14] & g[21347];
assign g[37732] = a[14] & g[21348];
assign g[54115] = b[14] & g[21348];
assign g[37733] = a[14] & g[21349];
assign g[54116] = b[14] & g[21349];
assign g[37734] = a[14] & g[21350];
assign g[54117] = b[14] & g[21350];
assign g[37735] = a[14] & g[21351];
assign g[54118] = b[14] & g[21351];
assign g[37736] = a[14] & g[21352];
assign g[54119] = b[14] & g[21352];
assign g[37737] = a[14] & g[21353];
assign g[54120] = b[14] & g[21353];
assign g[37738] = a[14] & g[21354];
assign g[54121] = b[14] & g[21354];
assign g[37739] = a[14] & g[21355];
assign g[54122] = b[14] & g[21355];
assign g[37740] = a[14] & g[21356];
assign g[54123] = b[14] & g[21356];
assign g[37741] = a[14] & g[21357];
assign g[54124] = b[14] & g[21357];
assign g[37742] = a[14] & g[21358];
assign g[54125] = b[14] & g[21358];
assign g[37743] = a[14] & g[21359];
assign g[54126] = b[14] & g[21359];
assign g[37744] = a[14] & g[21360];
assign g[54127] = b[14] & g[21360];
assign g[37745] = a[14] & g[21361];
assign g[54128] = b[14] & g[21361];
assign g[37746] = a[14] & g[21362];
assign g[54129] = b[14] & g[21362];
assign g[37747] = a[14] & g[21363];
assign g[54130] = b[14] & g[21363];
assign g[37748] = a[14] & g[21364];
assign g[54131] = b[14] & g[21364];
assign g[37749] = a[14] & g[21365];
assign g[54132] = b[14] & g[21365];
assign g[37750] = a[14] & g[21366];
assign g[54133] = b[14] & g[21366];
assign g[37751] = a[14] & g[21367];
assign g[54134] = b[14] & g[21367];
assign g[37752] = a[14] & g[21368];
assign g[54135] = b[14] & g[21368];
assign g[37753] = a[14] & g[21369];
assign g[54136] = b[14] & g[21369];
assign g[37754] = a[14] & g[21370];
assign g[54137] = b[14] & g[21370];
assign g[37755] = a[14] & g[21371];
assign g[54138] = b[14] & g[21371];
assign g[37756] = a[14] & g[21372];
assign g[54139] = b[14] & g[21372];
assign g[37757] = a[14] & g[21373];
assign g[54140] = b[14] & g[21373];
assign g[37758] = a[14] & g[21374];
assign g[54141] = b[14] & g[21374];
assign g[37759] = a[14] & g[21375];
assign g[54142] = b[14] & g[21375];
assign g[37760] = a[14] & g[21376];
assign g[54143] = b[14] & g[21376];
assign g[37761] = a[14] & g[21377];
assign g[54144] = b[14] & g[21377];
assign g[37762] = a[14] & g[21378];
assign g[54145] = b[14] & g[21378];
assign g[37763] = a[14] & g[21379];
assign g[54146] = b[14] & g[21379];
assign g[37764] = a[14] & g[21380];
assign g[54147] = b[14] & g[21380];
assign g[37765] = a[14] & g[21381];
assign g[54148] = b[14] & g[21381];
assign g[37766] = a[14] & g[21382];
assign g[54149] = b[14] & g[21382];
assign g[37767] = a[14] & g[21383];
assign g[54150] = b[14] & g[21383];
assign g[37768] = a[14] & g[21384];
assign g[54151] = b[14] & g[21384];
assign g[37769] = a[14] & g[21385];
assign g[54152] = b[14] & g[21385];
assign g[37770] = a[14] & g[21386];
assign g[54153] = b[14] & g[21386];
assign g[37771] = a[14] & g[21387];
assign g[54154] = b[14] & g[21387];
assign g[37772] = a[14] & g[21388];
assign g[54155] = b[14] & g[21388];
assign g[37773] = a[14] & g[21389];
assign g[54156] = b[14] & g[21389];
assign g[37774] = a[14] & g[21390];
assign g[54157] = b[14] & g[21390];
assign g[37775] = a[14] & g[21391];
assign g[54158] = b[14] & g[21391];
assign g[37776] = a[14] & g[21392];
assign g[54159] = b[14] & g[21392];
assign g[37777] = a[14] & g[21393];
assign g[54160] = b[14] & g[21393];
assign g[37778] = a[14] & g[21394];
assign g[54161] = b[14] & g[21394];
assign g[37779] = a[14] & g[21395];
assign g[54162] = b[14] & g[21395];
assign g[37780] = a[14] & g[21396];
assign g[54163] = b[14] & g[21396];
assign g[37781] = a[14] & g[21397];
assign g[54164] = b[14] & g[21397];
assign g[37782] = a[14] & g[21398];
assign g[54165] = b[14] & g[21398];
assign g[37783] = a[14] & g[21399];
assign g[54166] = b[14] & g[21399];
assign g[37784] = a[14] & g[21400];
assign g[54167] = b[14] & g[21400];
assign g[37785] = a[14] & g[21401];
assign g[54168] = b[14] & g[21401];
assign g[37786] = a[14] & g[21402];
assign g[54169] = b[14] & g[21402];
assign g[37787] = a[14] & g[21403];
assign g[54170] = b[14] & g[21403];
assign g[37788] = a[14] & g[21404];
assign g[54171] = b[14] & g[21404];
assign g[37789] = a[14] & g[21405];
assign g[54172] = b[14] & g[21405];
assign g[37790] = a[14] & g[21406];
assign g[54173] = b[14] & g[21406];
assign g[37791] = a[14] & g[21407];
assign g[54174] = b[14] & g[21407];
assign g[37792] = a[14] & g[21408];
assign g[54175] = b[14] & g[21408];
assign g[37793] = a[14] & g[21409];
assign g[54176] = b[14] & g[21409];
assign g[37794] = a[14] & g[21410];
assign g[54177] = b[14] & g[21410];
assign g[37795] = a[14] & g[21411];
assign g[54178] = b[14] & g[21411];
assign g[37796] = a[14] & g[21412];
assign g[54179] = b[14] & g[21412];
assign g[37797] = a[14] & g[21413];
assign g[54180] = b[14] & g[21413];
assign g[37798] = a[14] & g[21414];
assign g[54181] = b[14] & g[21414];
assign g[37799] = a[14] & g[21415];
assign g[54182] = b[14] & g[21415];
assign g[37800] = a[14] & g[21416];
assign g[54183] = b[14] & g[21416];
assign g[37801] = a[14] & g[21417];
assign g[54184] = b[14] & g[21417];
assign g[37802] = a[14] & g[21418];
assign g[54185] = b[14] & g[21418];
assign g[37803] = a[14] & g[21419];
assign g[54186] = b[14] & g[21419];
assign g[37804] = a[14] & g[21420];
assign g[54187] = b[14] & g[21420];
assign g[37805] = a[14] & g[21421];
assign g[54188] = b[14] & g[21421];
assign g[37806] = a[14] & g[21422];
assign g[54189] = b[14] & g[21422];
assign g[37807] = a[14] & g[21423];
assign g[54190] = b[14] & g[21423];
assign g[37808] = a[14] & g[21424];
assign g[54191] = b[14] & g[21424];
assign g[37809] = a[14] & g[21425];
assign g[54192] = b[14] & g[21425];
assign g[37810] = a[14] & g[21426];
assign g[54193] = b[14] & g[21426];
assign g[37811] = a[14] & g[21427];
assign g[54194] = b[14] & g[21427];
assign g[37812] = a[14] & g[21428];
assign g[54195] = b[14] & g[21428];
assign g[37813] = a[14] & g[21429];
assign g[54196] = b[14] & g[21429];
assign g[37814] = a[14] & g[21430];
assign g[54197] = b[14] & g[21430];
assign g[37815] = a[14] & g[21431];
assign g[54198] = b[14] & g[21431];
assign g[37816] = a[14] & g[21432];
assign g[54199] = b[14] & g[21432];
assign g[37817] = a[14] & g[21433];
assign g[54200] = b[14] & g[21433];
assign g[37818] = a[14] & g[21434];
assign g[54201] = b[14] & g[21434];
assign g[37819] = a[14] & g[21435];
assign g[54202] = b[14] & g[21435];
assign g[37820] = a[14] & g[21436];
assign g[54203] = b[14] & g[21436];
assign g[37821] = a[14] & g[21437];
assign g[54204] = b[14] & g[21437];
assign g[37822] = a[14] & g[21438];
assign g[54205] = b[14] & g[21438];
assign g[37823] = a[14] & g[21439];
assign g[54206] = b[14] & g[21439];
assign g[37824] = a[14] & g[21440];
assign g[54207] = b[14] & g[21440];
assign g[37825] = a[14] & g[21441];
assign g[54208] = b[14] & g[21441];
assign g[37826] = a[14] & g[21442];
assign g[54209] = b[14] & g[21442];
assign g[37827] = a[14] & g[21443];
assign g[54210] = b[14] & g[21443];
assign g[37828] = a[14] & g[21444];
assign g[54211] = b[14] & g[21444];
assign g[37829] = a[14] & g[21445];
assign g[54212] = b[14] & g[21445];
assign g[37830] = a[14] & g[21446];
assign g[54213] = b[14] & g[21446];
assign g[37831] = a[14] & g[21447];
assign g[54214] = b[14] & g[21447];
assign g[37832] = a[14] & g[21448];
assign g[54215] = b[14] & g[21448];
assign g[37833] = a[14] & g[21449];
assign g[54216] = b[14] & g[21449];
assign g[37834] = a[14] & g[21450];
assign g[54217] = b[14] & g[21450];
assign g[37835] = a[14] & g[21451];
assign g[54218] = b[14] & g[21451];
assign g[37836] = a[14] & g[21452];
assign g[54219] = b[14] & g[21452];
assign g[37837] = a[14] & g[21453];
assign g[54220] = b[14] & g[21453];
assign g[37838] = a[14] & g[21454];
assign g[54221] = b[14] & g[21454];
assign g[37839] = a[14] & g[21455];
assign g[54222] = b[14] & g[21455];
assign g[37840] = a[14] & g[21456];
assign g[54223] = b[14] & g[21456];
assign g[37841] = a[14] & g[21457];
assign g[54224] = b[14] & g[21457];
assign g[37842] = a[14] & g[21458];
assign g[54225] = b[14] & g[21458];
assign g[37843] = a[14] & g[21459];
assign g[54226] = b[14] & g[21459];
assign g[37844] = a[14] & g[21460];
assign g[54227] = b[14] & g[21460];
assign g[37845] = a[14] & g[21461];
assign g[54228] = b[14] & g[21461];
assign g[37846] = a[14] & g[21462];
assign g[54229] = b[14] & g[21462];
assign g[37847] = a[14] & g[21463];
assign g[54230] = b[14] & g[21463];
assign g[37848] = a[14] & g[21464];
assign g[54231] = b[14] & g[21464];
assign g[37849] = a[14] & g[21465];
assign g[54232] = b[14] & g[21465];
assign g[37850] = a[14] & g[21466];
assign g[54233] = b[14] & g[21466];
assign g[37851] = a[14] & g[21467];
assign g[54234] = b[14] & g[21467];
assign g[37852] = a[14] & g[21468];
assign g[54235] = b[14] & g[21468];
assign g[37853] = a[14] & g[21469];
assign g[54236] = b[14] & g[21469];
assign g[37854] = a[14] & g[21470];
assign g[54237] = b[14] & g[21470];
assign g[37855] = a[14] & g[21471];
assign g[54238] = b[14] & g[21471];
assign g[37856] = a[14] & g[21472];
assign g[54239] = b[14] & g[21472];
assign g[37857] = a[14] & g[21473];
assign g[54240] = b[14] & g[21473];
assign g[37858] = a[14] & g[21474];
assign g[54241] = b[14] & g[21474];
assign g[37859] = a[14] & g[21475];
assign g[54242] = b[14] & g[21475];
assign g[37860] = a[14] & g[21476];
assign g[54243] = b[14] & g[21476];
assign g[37861] = a[14] & g[21477];
assign g[54244] = b[14] & g[21477];
assign g[37862] = a[14] & g[21478];
assign g[54245] = b[14] & g[21478];
assign g[37863] = a[14] & g[21479];
assign g[54246] = b[14] & g[21479];
assign g[37864] = a[14] & g[21480];
assign g[54247] = b[14] & g[21480];
assign g[37865] = a[14] & g[21481];
assign g[54248] = b[14] & g[21481];
assign g[37866] = a[14] & g[21482];
assign g[54249] = b[14] & g[21482];
assign g[37867] = a[14] & g[21483];
assign g[54250] = b[14] & g[21483];
assign g[37868] = a[14] & g[21484];
assign g[54251] = b[14] & g[21484];
assign g[37869] = a[14] & g[21485];
assign g[54252] = b[14] & g[21485];
assign g[37870] = a[14] & g[21486];
assign g[54253] = b[14] & g[21486];
assign g[37871] = a[14] & g[21487];
assign g[54254] = b[14] & g[21487];
assign g[37872] = a[14] & g[21488];
assign g[54255] = b[14] & g[21488];
assign g[37873] = a[14] & g[21489];
assign g[54256] = b[14] & g[21489];
assign g[37874] = a[14] & g[21490];
assign g[54257] = b[14] & g[21490];
assign g[37875] = a[14] & g[21491];
assign g[54258] = b[14] & g[21491];
assign g[37876] = a[14] & g[21492];
assign g[54259] = b[14] & g[21492];
assign g[37877] = a[14] & g[21493];
assign g[54260] = b[14] & g[21493];
assign g[37878] = a[14] & g[21494];
assign g[54261] = b[14] & g[21494];
assign g[37879] = a[14] & g[21495];
assign g[54262] = b[14] & g[21495];
assign g[37880] = a[14] & g[21496];
assign g[54263] = b[14] & g[21496];
assign g[37881] = a[14] & g[21497];
assign g[54264] = b[14] & g[21497];
assign g[37882] = a[14] & g[21498];
assign g[54265] = b[14] & g[21498];
assign g[37883] = a[14] & g[21499];
assign g[54266] = b[14] & g[21499];
assign g[37884] = a[14] & g[21500];
assign g[54267] = b[14] & g[21500];
assign g[37885] = a[14] & g[21501];
assign g[54268] = b[14] & g[21501];
assign g[37886] = a[14] & g[21502];
assign g[54269] = b[14] & g[21502];
assign g[37887] = a[14] & g[21503];
assign g[54270] = b[14] & g[21503];
assign g[37888] = a[14] & g[21504];
assign g[54271] = b[14] & g[21504];
assign g[37889] = a[14] & g[21505];
assign g[54272] = b[14] & g[21505];
assign g[37890] = a[14] & g[21506];
assign g[54273] = b[14] & g[21506];
assign g[37891] = a[14] & g[21507];
assign g[54274] = b[14] & g[21507];
assign g[37892] = a[14] & g[21508];
assign g[54275] = b[14] & g[21508];
assign g[37893] = a[14] & g[21509];
assign g[54276] = b[14] & g[21509];
assign g[37894] = a[14] & g[21510];
assign g[54277] = b[14] & g[21510];
assign g[37895] = a[14] & g[21511];
assign g[54278] = b[14] & g[21511];
assign g[37896] = a[14] & g[21512];
assign g[54279] = b[14] & g[21512];
assign g[37897] = a[14] & g[21513];
assign g[54280] = b[14] & g[21513];
assign g[37898] = a[14] & g[21514];
assign g[54281] = b[14] & g[21514];
assign g[37899] = a[14] & g[21515];
assign g[54282] = b[14] & g[21515];
assign g[37900] = a[14] & g[21516];
assign g[54283] = b[14] & g[21516];
assign g[37901] = a[14] & g[21517];
assign g[54284] = b[14] & g[21517];
assign g[37902] = a[14] & g[21518];
assign g[54285] = b[14] & g[21518];
assign g[37903] = a[14] & g[21519];
assign g[54286] = b[14] & g[21519];
assign g[37904] = a[14] & g[21520];
assign g[54287] = b[14] & g[21520];
assign g[37905] = a[14] & g[21521];
assign g[54288] = b[14] & g[21521];
assign g[37906] = a[14] & g[21522];
assign g[54289] = b[14] & g[21522];
assign g[37907] = a[14] & g[21523];
assign g[54290] = b[14] & g[21523];
assign g[37908] = a[14] & g[21524];
assign g[54291] = b[14] & g[21524];
assign g[37909] = a[14] & g[21525];
assign g[54292] = b[14] & g[21525];
assign g[37910] = a[14] & g[21526];
assign g[54293] = b[14] & g[21526];
assign g[37911] = a[14] & g[21527];
assign g[54294] = b[14] & g[21527];
assign g[37912] = a[14] & g[21528];
assign g[54295] = b[14] & g[21528];
assign g[37913] = a[14] & g[21529];
assign g[54296] = b[14] & g[21529];
assign g[37914] = a[14] & g[21530];
assign g[54297] = b[14] & g[21530];
assign g[37915] = a[14] & g[21531];
assign g[54298] = b[14] & g[21531];
assign g[37916] = a[14] & g[21532];
assign g[54299] = b[14] & g[21532];
assign g[37917] = a[14] & g[21533];
assign g[54300] = b[14] & g[21533];
assign g[37918] = a[14] & g[21534];
assign g[54301] = b[14] & g[21534];
assign g[37919] = a[14] & g[21535];
assign g[54302] = b[14] & g[21535];
assign g[37920] = a[14] & g[21536];
assign g[54303] = b[14] & g[21536];
assign g[37921] = a[14] & g[21537];
assign g[54304] = b[14] & g[21537];
assign g[37922] = a[14] & g[21538];
assign g[54305] = b[14] & g[21538];
assign g[37923] = a[14] & g[21539];
assign g[54306] = b[14] & g[21539];
assign g[37924] = a[14] & g[21540];
assign g[54307] = b[14] & g[21540];
assign g[37925] = a[14] & g[21541];
assign g[54308] = b[14] & g[21541];
assign g[37926] = a[14] & g[21542];
assign g[54309] = b[14] & g[21542];
assign g[37927] = a[14] & g[21543];
assign g[54310] = b[14] & g[21543];
assign g[37928] = a[14] & g[21544];
assign g[54311] = b[14] & g[21544];
assign g[37929] = a[14] & g[21545];
assign g[54312] = b[14] & g[21545];
assign g[37930] = a[14] & g[21546];
assign g[54313] = b[14] & g[21546];
assign g[37931] = a[14] & g[21547];
assign g[54314] = b[14] & g[21547];
assign g[37932] = a[14] & g[21548];
assign g[54315] = b[14] & g[21548];
assign g[37933] = a[14] & g[21549];
assign g[54316] = b[14] & g[21549];
assign g[37934] = a[14] & g[21550];
assign g[54317] = b[14] & g[21550];
assign g[37935] = a[14] & g[21551];
assign g[54318] = b[14] & g[21551];
assign g[37936] = a[14] & g[21552];
assign g[54319] = b[14] & g[21552];
assign g[37937] = a[14] & g[21553];
assign g[54320] = b[14] & g[21553];
assign g[37938] = a[14] & g[21554];
assign g[54321] = b[14] & g[21554];
assign g[37939] = a[14] & g[21555];
assign g[54322] = b[14] & g[21555];
assign g[37940] = a[14] & g[21556];
assign g[54323] = b[14] & g[21556];
assign g[37941] = a[14] & g[21557];
assign g[54324] = b[14] & g[21557];
assign g[37942] = a[14] & g[21558];
assign g[54325] = b[14] & g[21558];
assign g[37943] = a[14] & g[21559];
assign g[54326] = b[14] & g[21559];
assign g[37944] = a[14] & g[21560];
assign g[54327] = b[14] & g[21560];
assign g[37945] = a[14] & g[21561];
assign g[54328] = b[14] & g[21561];
assign g[37946] = a[14] & g[21562];
assign g[54329] = b[14] & g[21562];
assign g[37947] = a[14] & g[21563];
assign g[54330] = b[14] & g[21563];
assign g[37948] = a[14] & g[21564];
assign g[54331] = b[14] & g[21564];
assign g[37949] = a[14] & g[21565];
assign g[54332] = b[14] & g[21565];
assign g[37950] = a[14] & g[21566];
assign g[54333] = b[14] & g[21566];
assign g[37951] = a[14] & g[21567];
assign g[54334] = b[14] & g[21567];
assign g[37952] = a[14] & g[21568];
assign g[54335] = b[14] & g[21568];
assign g[37953] = a[14] & g[21569];
assign g[54336] = b[14] & g[21569];
assign g[37954] = a[14] & g[21570];
assign g[54337] = b[14] & g[21570];
assign g[37955] = a[14] & g[21571];
assign g[54338] = b[14] & g[21571];
assign g[37956] = a[14] & g[21572];
assign g[54339] = b[14] & g[21572];
assign g[37957] = a[14] & g[21573];
assign g[54340] = b[14] & g[21573];
assign g[37958] = a[14] & g[21574];
assign g[54341] = b[14] & g[21574];
assign g[37959] = a[14] & g[21575];
assign g[54342] = b[14] & g[21575];
assign g[37960] = a[14] & g[21576];
assign g[54343] = b[14] & g[21576];
assign g[37961] = a[14] & g[21577];
assign g[54344] = b[14] & g[21577];
assign g[37962] = a[14] & g[21578];
assign g[54345] = b[14] & g[21578];
assign g[37963] = a[14] & g[21579];
assign g[54346] = b[14] & g[21579];
assign g[37964] = a[14] & g[21580];
assign g[54347] = b[14] & g[21580];
assign g[37965] = a[14] & g[21581];
assign g[54348] = b[14] & g[21581];
assign g[37966] = a[14] & g[21582];
assign g[54349] = b[14] & g[21582];
assign g[37967] = a[14] & g[21583];
assign g[54350] = b[14] & g[21583];
assign g[37968] = a[14] & g[21584];
assign g[54351] = b[14] & g[21584];
assign g[37969] = a[14] & g[21585];
assign g[54352] = b[14] & g[21585];
assign g[37970] = a[14] & g[21586];
assign g[54353] = b[14] & g[21586];
assign g[37971] = a[14] & g[21587];
assign g[54354] = b[14] & g[21587];
assign g[37972] = a[14] & g[21588];
assign g[54355] = b[14] & g[21588];
assign g[37973] = a[14] & g[21589];
assign g[54356] = b[14] & g[21589];
assign g[37974] = a[14] & g[21590];
assign g[54357] = b[14] & g[21590];
assign g[37975] = a[14] & g[21591];
assign g[54358] = b[14] & g[21591];
assign g[37976] = a[14] & g[21592];
assign g[54359] = b[14] & g[21592];
assign g[37977] = a[14] & g[21593];
assign g[54360] = b[14] & g[21593];
assign g[37978] = a[14] & g[21594];
assign g[54361] = b[14] & g[21594];
assign g[37979] = a[14] & g[21595];
assign g[54362] = b[14] & g[21595];
assign g[37980] = a[14] & g[21596];
assign g[54363] = b[14] & g[21596];
assign g[37981] = a[14] & g[21597];
assign g[54364] = b[14] & g[21597];
assign g[37982] = a[14] & g[21598];
assign g[54365] = b[14] & g[21598];
assign g[37983] = a[14] & g[21599];
assign g[54366] = b[14] & g[21599];
assign g[37984] = a[14] & g[21600];
assign g[54367] = b[14] & g[21600];
assign g[37985] = a[14] & g[21601];
assign g[54368] = b[14] & g[21601];
assign g[37986] = a[14] & g[21602];
assign g[54369] = b[14] & g[21602];
assign g[37987] = a[14] & g[21603];
assign g[54370] = b[14] & g[21603];
assign g[37988] = a[14] & g[21604];
assign g[54371] = b[14] & g[21604];
assign g[37989] = a[14] & g[21605];
assign g[54372] = b[14] & g[21605];
assign g[37990] = a[14] & g[21606];
assign g[54373] = b[14] & g[21606];
assign g[37991] = a[14] & g[21607];
assign g[54374] = b[14] & g[21607];
assign g[37992] = a[14] & g[21608];
assign g[54375] = b[14] & g[21608];
assign g[37993] = a[14] & g[21609];
assign g[54376] = b[14] & g[21609];
assign g[37994] = a[14] & g[21610];
assign g[54377] = b[14] & g[21610];
assign g[37995] = a[14] & g[21611];
assign g[54378] = b[14] & g[21611];
assign g[37996] = a[14] & g[21612];
assign g[54379] = b[14] & g[21612];
assign g[37997] = a[14] & g[21613];
assign g[54380] = b[14] & g[21613];
assign g[37998] = a[14] & g[21614];
assign g[54381] = b[14] & g[21614];
assign g[37999] = a[14] & g[21615];
assign g[54382] = b[14] & g[21615];
assign g[38000] = a[14] & g[21616];
assign g[54383] = b[14] & g[21616];
assign g[38001] = a[14] & g[21617];
assign g[54384] = b[14] & g[21617];
assign g[38002] = a[14] & g[21618];
assign g[54385] = b[14] & g[21618];
assign g[38003] = a[14] & g[21619];
assign g[54386] = b[14] & g[21619];
assign g[38004] = a[14] & g[21620];
assign g[54387] = b[14] & g[21620];
assign g[38005] = a[14] & g[21621];
assign g[54388] = b[14] & g[21621];
assign g[38006] = a[14] & g[21622];
assign g[54389] = b[14] & g[21622];
assign g[38007] = a[14] & g[21623];
assign g[54390] = b[14] & g[21623];
assign g[38008] = a[14] & g[21624];
assign g[54391] = b[14] & g[21624];
assign g[38009] = a[14] & g[21625];
assign g[54392] = b[14] & g[21625];
assign g[38010] = a[14] & g[21626];
assign g[54393] = b[14] & g[21626];
assign g[38011] = a[14] & g[21627];
assign g[54394] = b[14] & g[21627];
assign g[38012] = a[14] & g[21628];
assign g[54395] = b[14] & g[21628];
assign g[38013] = a[14] & g[21629];
assign g[54396] = b[14] & g[21629];
assign g[38014] = a[14] & g[21630];
assign g[54397] = b[14] & g[21630];
assign g[38015] = a[14] & g[21631];
assign g[54398] = b[14] & g[21631];
assign g[38016] = a[14] & g[21632];
assign g[54399] = b[14] & g[21632];
assign g[38017] = a[14] & g[21633];
assign g[54400] = b[14] & g[21633];
assign g[38018] = a[14] & g[21634];
assign g[54401] = b[14] & g[21634];
assign g[38019] = a[14] & g[21635];
assign g[54402] = b[14] & g[21635];
assign g[38020] = a[14] & g[21636];
assign g[54403] = b[14] & g[21636];
assign g[38021] = a[14] & g[21637];
assign g[54404] = b[14] & g[21637];
assign g[38022] = a[14] & g[21638];
assign g[54405] = b[14] & g[21638];
assign g[38023] = a[14] & g[21639];
assign g[54406] = b[14] & g[21639];
assign g[38024] = a[14] & g[21640];
assign g[54407] = b[14] & g[21640];
assign g[38025] = a[14] & g[21641];
assign g[54408] = b[14] & g[21641];
assign g[38026] = a[14] & g[21642];
assign g[54409] = b[14] & g[21642];
assign g[38027] = a[14] & g[21643];
assign g[54410] = b[14] & g[21643];
assign g[38028] = a[14] & g[21644];
assign g[54411] = b[14] & g[21644];
assign g[38029] = a[14] & g[21645];
assign g[54412] = b[14] & g[21645];
assign g[38030] = a[14] & g[21646];
assign g[54413] = b[14] & g[21646];
assign g[38031] = a[14] & g[21647];
assign g[54414] = b[14] & g[21647];
assign g[38032] = a[14] & g[21648];
assign g[54415] = b[14] & g[21648];
assign g[38033] = a[14] & g[21649];
assign g[54416] = b[14] & g[21649];
assign g[38034] = a[14] & g[21650];
assign g[54417] = b[14] & g[21650];
assign g[38035] = a[14] & g[21651];
assign g[54418] = b[14] & g[21651];
assign g[38036] = a[14] & g[21652];
assign g[54419] = b[14] & g[21652];
assign g[38037] = a[14] & g[21653];
assign g[54420] = b[14] & g[21653];
assign g[38038] = a[14] & g[21654];
assign g[54421] = b[14] & g[21654];
assign g[38039] = a[14] & g[21655];
assign g[54422] = b[14] & g[21655];
assign g[38040] = a[14] & g[21656];
assign g[54423] = b[14] & g[21656];
assign g[38041] = a[14] & g[21657];
assign g[54424] = b[14] & g[21657];
assign g[38042] = a[14] & g[21658];
assign g[54425] = b[14] & g[21658];
assign g[38043] = a[14] & g[21659];
assign g[54426] = b[14] & g[21659];
assign g[38044] = a[14] & g[21660];
assign g[54427] = b[14] & g[21660];
assign g[38045] = a[14] & g[21661];
assign g[54428] = b[14] & g[21661];
assign g[38046] = a[14] & g[21662];
assign g[54429] = b[14] & g[21662];
assign g[38047] = a[14] & g[21663];
assign g[54430] = b[14] & g[21663];
assign g[38048] = a[14] & g[21664];
assign g[54431] = b[14] & g[21664];
assign g[38049] = a[14] & g[21665];
assign g[54432] = b[14] & g[21665];
assign g[38050] = a[14] & g[21666];
assign g[54433] = b[14] & g[21666];
assign g[38051] = a[14] & g[21667];
assign g[54434] = b[14] & g[21667];
assign g[38052] = a[14] & g[21668];
assign g[54435] = b[14] & g[21668];
assign g[38053] = a[14] & g[21669];
assign g[54436] = b[14] & g[21669];
assign g[38054] = a[14] & g[21670];
assign g[54437] = b[14] & g[21670];
assign g[38055] = a[14] & g[21671];
assign g[54438] = b[14] & g[21671];
assign g[38056] = a[14] & g[21672];
assign g[54439] = b[14] & g[21672];
assign g[38057] = a[14] & g[21673];
assign g[54440] = b[14] & g[21673];
assign g[38058] = a[14] & g[21674];
assign g[54441] = b[14] & g[21674];
assign g[38059] = a[14] & g[21675];
assign g[54442] = b[14] & g[21675];
assign g[38060] = a[14] & g[21676];
assign g[54443] = b[14] & g[21676];
assign g[38061] = a[14] & g[21677];
assign g[54444] = b[14] & g[21677];
assign g[38062] = a[14] & g[21678];
assign g[54445] = b[14] & g[21678];
assign g[38063] = a[14] & g[21679];
assign g[54446] = b[14] & g[21679];
assign g[38064] = a[14] & g[21680];
assign g[54447] = b[14] & g[21680];
assign g[38065] = a[14] & g[21681];
assign g[54448] = b[14] & g[21681];
assign g[38066] = a[14] & g[21682];
assign g[54449] = b[14] & g[21682];
assign g[38067] = a[14] & g[21683];
assign g[54450] = b[14] & g[21683];
assign g[38068] = a[14] & g[21684];
assign g[54451] = b[14] & g[21684];
assign g[38069] = a[14] & g[21685];
assign g[54452] = b[14] & g[21685];
assign g[38070] = a[14] & g[21686];
assign g[54453] = b[14] & g[21686];
assign g[38071] = a[14] & g[21687];
assign g[54454] = b[14] & g[21687];
assign g[38072] = a[14] & g[21688];
assign g[54455] = b[14] & g[21688];
assign g[38073] = a[14] & g[21689];
assign g[54456] = b[14] & g[21689];
assign g[38074] = a[14] & g[21690];
assign g[54457] = b[14] & g[21690];
assign g[38075] = a[14] & g[21691];
assign g[54458] = b[14] & g[21691];
assign g[38076] = a[14] & g[21692];
assign g[54459] = b[14] & g[21692];
assign g[38077] = a[14] & g[21693];
assign g[54460] = b[14] & g[21693];
assign g[38078] = a[14] & g[21694];
assign g[54461] = b[14] & g[21694];
assign g[38079] = a[14] & g[21695];
assign g[54462] = b[14] & g[21695];
assign g[38080] = a[14] & g[21696];
assign g[54463] = b[14] & g[21696];
assign g[38081] = a[14] & g[21697];
assign g[54464] = b[14] & g[21697];
assign g[38082] = a[14] & g[21698];
assign g[54465] = b[14] & g[21698];
assign g[38083] = a[14] & g[21699];
assign g[54466] = b[14] & g[21699];
assign g[38084] = a[14] & g[21700];
assign g[54467] = b[14] & g[21700];
assign g[38085] = a[14] & g[21701];
assign g[54468] = b[14] & g[21701];
assign g[38086] = a[14] & g[21702];
assign g[54469] = b[14] & g[21702];
assign g[38087] = a[14] & g[21703];
assign g[54470] = b[14] & g[21703];
assign g[38088] = a[14] & g[21704];
assign g[54471] = b[14] & g[21704];
assign g[38089] = a[14] & g[21705];
assign g[54472] = b[14] & g[21705];
assign g[38090] = a[14] & g[21706];
assign g[54473] = b[14] & g[21706];
assign g[38091] = a[14] & g[21707];
assign g[54474] = b[14] & g[21707];
assign g[38092] = a[14] & g[21708];
assign g[54475] = b[14] & g[21708];
assign g[38093] = a[14] & g[21709];
assign g[54476] = b[14] & g[21709];
assign g[38094] = a[14] & g[21710];
assign g[54477] = b[14] & g[21710];
assign g[38095] = a[14] & g[21711];
assign g[54478] = b[14] & g[21711];
assign g[38096] = a[14] & g[21712];
assign g[54479] = b[14] & g[21712];
assign g[38097] = a[14] & g[21713];
assign g[54480] = b[14] & g[21713];
assign g[38098] = a[14] & g[21714];
assign g[54481] = b[14] & g[21714];
assign g[38099] = a[14] & g[21715];
assign g[54482] = b[14] & g[21715];
assign g[38100] = a[14] & g[21716];
assign g[54483] = b[14] & g[21716];
assign g[38101] = a[14] & g[21717];
assign g[54484] = b[14] & g[21717];
assign g[38102] = a[14] & g[21718];
assign g[54485] = b[14] & g[21718];
assign g[38103] = a[14] & g[21719];
assign g[54486] = b[14] & g[21719];
assign g[38104] = a[14] & g[21720];
assign g[54487] = b[14] & g[21720];
assign g[38105] = a[14] & g[21721];
assign g[54488] = b[14] & g[21721];
assign g[38106] = a[14] & g[21722];
assign g[54489] = b[14] & g[21722];
assign g[38107] = a[14] & g[21723];
assign g[54490] = b[14] & g[21723];
assign g[38108] = a[14] & g[21724];
assign g[54491] = b[14] & g[21724];
assign g[38109] = a[14] & g[21725];
assign g[54492] = b[14] & g[21725];
assign g[38110] = a[14] & g[21726];
assign g[54493] = b[14] & g[21726];
assign g[38111] = a[14] & g[21727];
assign g[54494] = b[14] & g[21727];
assign g[38112] = a[14] & g[21728];
assign g[54495] = b[14] & g[21728];
assign g[38113] = a[14] & g[21729];
assign g[54496] = b[14] & g[21729];
assign g[38114] = a[14] & g[21730];
assign g[54497] = b[14] & g[21730];
assign g[38115] = a[14] & g[21731];
assign g[54498] = b[14] & g[21731];
assign g[38116] = a[14] & g[21732];
assign g[54499] = b[14] & g[21732];
assign g[38117] = a[14] & g[21733];
assign g[54500] = b[14] & g[21733];
assign g[38118] = a[14] & g[21734];
assign g[54501] = b[14] & g[21734];
assign g[38119] = a[14] & g[21735];
assign g[54502] = b[14] & g[21735];
assign g[38120] = a[14] & g[21736];
assign g[54503] = b[14] & g[21736];
assign g[38121] = a[14] & g[21737];
assign g[54504] = b[14] & g[21737];
assign g[38122] = a[14] & g[21738];
assign g[54505] = b[14] & g[21738];
assign g[38123] = a[14] & g[21739];
assign g[54506] = b[14] & g[21739];
assign g[38124] = a[14] & g[21740];
assign g[54507] = b[14] & g[21740];
assign g[38125] = a[14] & g[21741];
assign g[54508] = b[14] & g[21741];
assign g[38126] = a[14] & g[21742];
assign g[54509] = b[14] & g[21742];
assign g[38127] = a[14] & g[21743];
assign g[54510] = b[14] & g[21743];
assign g[38128] = a[14] & g[21744];
assign g[54511] = b[14] & g[21744];
assign g[38129] = a[14] & g[21745];
assign g[54512] = b[14] & g[21745];
assign g[38130] = a[14] & g[21746];
assign g[54513] = b[14] & g[21746];
assign g[38131] = a[14] & g[21747];
assign g[54514] = b[14] & g[21747];
assign g[38132] = a[14] & g[21748];
assign g[54515] = b[14] & g[21748];
assign g[38133] = a[14] & g[21749];
assign g[54516] = b[14] & g[21749];
assign g[38134] = a[14] & g[21750];
assign g[54517] = b[14] & g[21750];
assign g[38135] = a[14] & g[21751];
assign g[54518] = b[14] & g[21751];
assign g[38136] = a[14] & g[21752];
assign g[54519] = b[14] & g[21752];
assign g[38137] = a[14] & g[21753];
assign g[54520] = b[14] & g[21753];
assign g[38138] = a[14] & g[21754];
assign g[54521] = b[14] & g[21754];
assign g[38139] = a[14] & g[21755];
assign g[54522] = b[14] & g[21755];
assign g[38140] = a[14] & g[21756];
assign g[54523] = b[14] & g[21756];
assign g[38141] = a[14] & g[21757];
assign g[54524] = b[14] & g[21757];
assign g[38142] = a[14] & g[21758];
assign g[54525] = b[14] & g[21758];
assign g[38143] = a[14] & g[21759];
assign g[54526] = b[14] & g[21759];
assign g[38144] = a[14] & g[21760];
assign g[54527] = b[14] & g[21760];
assign g[38145] = a[14] & g[21761];
assign g[54528] = b[14] & g[21761];
assign g[38146] = a[14] & g[21762];
assign g[54529] = b[14] & g[21762];
assign g[38147] = a[14] & g[21763];
assign g[54530] = b[14] & g[21763];
assign g[38148] = a[14] & g[21764];
assign g[54531] = b[14] & g[21764];
assign g[38149] = a[14] & g[21765];
assign g[54532] = b[14] & g[21765];
assign g[38150] = a[14] & g[21766];
assign g[54533] = b[14] & g[21766];
assign g[38151] = a[14] & g[21767];
assign g[54534] = b[14] & g[21767];
assign g[38152] = a[14] & g[21768];
assign g[54535] = b[14] & g[21768];
assign g[38153] = a[14] & g[21769];
assign g[54536] = b[14] & g[21769];
assign g[38154] = a[14] & g[21770];
assign g[54537] = b[14] & g[21770];
assign g[38155] = a[14] & g[21771];
assign g[54538] = b[14] & g[21771];
assign g[38156] = a[14] & g[21772];
assign g[54539] = b[14] & g[21772];
assign g[38157] = a[14] & g[21773];
assign g[54540] = b[14] & g[21773];
assign g[38158] = a[14] & g[21774];
assign g[54541] = b[14] & g[21774];
assign g[38159] = a[14] & g[21775];
assign g[54542] = b[14] & g[21775];
assign g[38160] = a[14] & g[21776];
assign g[54543] = b[14] & g[21776];
assign g[38161] = a[14] & g[21777];
assign g[54544] = b[14] & g[21777];
assign g[38162] = a[14] & g[21778];
assign g[54545] = b[14] & g[21778];
assign g[38163] = a[14] & g[21779];
assign g[54546] = b[14] & g[21779];
assign g[38164] = a[14] & g[21780];
assign g[54547] = b[14] & g[21780];
assign g[38165] = a[14] & g[21781];
assign g[54548] = b[14] & g[21781];
assign g[38166] = a[14] & g[21782];
assign g[54549] = b[14] & g[21782];
assign g[38167] = a[14] & g[21783];
assign g[54550] = b[14] & g[21783];
assign g[38168] = a[14] & g[21784];
assign g[54551] = b[14] & g[21784];
assign g[38169] = a[14] & g[21785];
assign g[54552] = b[14] & g[21785];
assign g[38170] = a[14] & g[21786];
assign g[54553] = b[14] & g[21786];
assign g[38171] = a[14] & g[21787];
assign g[54554] = b[14] & g[21787];
assign g[38172] = a[14] & g[21788];
assign g[54555] = b[14] & g[21788];
assign g[38173] = a[14] & g[21789];
assign g[54556] = b[14] & g[21789];
assign g[38174] = a[14] & g[21790];
assign g[54557] = b[14] & g[21790];
assign g[38175] = a[14] & g[21791];
assign g[54558] = b[14] & g[21791];
assign g[38176] = a[14] & g[21792];
assign g[54559] = b[14] & g[21792];
assign g[38177] = a[14] & g[21793];
assign g[54560] = b[14] & g[21793];
assign g[38178] = a[14] & g[21794];
assign g[54561] = b[14] & g[21794];
assign g[38179] = a[14] & g[21795];
assign g[54562] = b[14] & g[21795];
assign g[38180] = a[14] & g[21796];
assign g[54563] = b[14] & g[21796];
assign g[38181] = a[14] & g[21797];
assign g[54564] = b[14] & g[21797];
assign g[38182] = a[14] & g[21798];
assign g[54565] = b[14] & g[21798];
assign g[38183] = a[14] & g[21799];
assign g[54566] = b[14] & g[21799];
assign g[38184] = a[14] & g[21800];
assign g[54567] = b[14] & g[21800];
assign g[38185] = a[14] & g[21801];
assign g[54568] = b[14] & g[21801];
assign g[38186] = a[14] & g[21802];
assign g[54569] = b[14] & g[21802];
assign g[38187] = a[14] & g[21803];
assign g[54570] = b[14] & g[21803];
assign g[38188] = a[14] & g[21804];
assign g[54571] = b[14] & g[21804];
assign g[38189] = a[14] & g[21805];
assign g[54572] = b[14] & g[21805];
assign g[38190] = a[14] & g[21806];
assign g[54573] = b[14] & g[21806];
assign g[38191] = a[14] & g[21807];
assign g[54574] = b[14] & g[21807];
assign g[38192] = a[14] & g[21808];
assign g[54575] = b[14] & g[21808];
assign g[38193] = a[14] & g[21809];
assign g[54576] = b[14] & g[21809];
assign g[38194] = a[14] & g[21810];
assign g[54577] = b[14] & g[21810];
assign g[38195] = a[14] & g[21811];
assign g[54578] = b[14] & g[21811];
assign g[38196] = a[14] & g[21812];
assign g[54579] = b[14] & g[21812];
assign g[38197] = a[14] & g[21813];
assign g[54580] = b[14] & g[21813];
assign g[38198] = a[14] & g[21814];
assign g[54581] = b[14] & g[21814];
assign g[38199] = a[14] & g[21815];
assign g[54582] = b[14] & g[21815];
assign g[38200] = a[14] & g[21816];
assign g[54583] = b[14] & g[21816];
assign g[38201] = a[14] & g[21817];
assign g[54584] = b[14] & g[21817];
assign g[38202] = a[14] & g[21818];
assign g[54585] = b[14] & g[21818];
assign g[38203] = a[14] & g[21819];
assign g[54586] = b[14] & g[21819];
assign g[38204] = a[14] & g[21820];
assign g[54587] = b[14] & g[21820];
assign g[38205] = a[14] & g[21821];
assign g[54588] = b[14] & g[21821];
assign g[38206] = a[14] & g[21822];
assign g[54589] = b[14] & g[21822];
assign g[38207] = a[14] & g[21823];
assign g[54590] = b[14] & g[21823];
assign g[38208] = a[14] & g[21824];
assign g[54591] = b[14] & g[21824];
assign g[38209] = a[14] & g[21825];
assign g[54592] = b[14] & g[21825];
assign g[38210] = a[14] & g[21826];
assign g[54593] = b[14] & g[21826];
assign g[38211] = a[14] & g[21827];
assign g[54594] = b[14] & g[21827];
assign g[38212] = a[14] & g[21828];
assign g[54595] = b[14] & g[21828];
assign g[38213] = a[14] & g[21829];
assign g[54596] = b[14] & g[21829];
assign g[38214] = a[14] & g[21830];
assign g[54597] = b[14] & g[21830];
assign g[38215] = a[14] & g[21831];
assign g[54598] = b[14] & g[21831];
assign g[38216] = a[14] & g[21832];
assign g[54599] = b[14] & g[21832];
assign g[38217] = a[14] & g[21833];
assign g[54600] = b[14] & g[21833];
assign g[38218] = a[14] & g[21834];
assign g[54601] = b[14] & g[21834];
assign g[38219] = a[14] & g[21835];
assign g[54602] = b[14] & g[21835];
assign g[38220] = a[14] & g[21836];
assign g[54603] = b[14] & g[21836];
assign g[38221] = a[14] & g[21837];
assign g[54604] = b[14] & g[21837];
assign g[38222] = a[14] & g[21838];
assign g[54605] = b[14] & g[21838];
assign g[38223] = a[14] & g[21839];
assign g[54606] = b[14] & g[21839];
assign g[38224] = a[14] & g[21840];
assign g[54607] = b[14] & g[21840];
assign g[38225] = a[14] & g[21841];
assign g[54608] = b[14] & g[21841];
assign g[38226] = a[14] & g[21842];
assign g[54609] = b[14] & g[21842];
assign g[38227] = a[14] & g[21843];
assign g[54610] = b[14] & g[21843];
assign g[38228] = a[14] & g[21844];
assign g[54611] = b[14] & g[21844];
assign g[38229] = a[14] & g[21845];
assign g[54612] = b[14] & g[21845];
assign g[38230] = a[14] & g[21846];
assign g[54613] = b[14] & g[21846];
assign g[38231] = a[14] & g[21847];
assign g[54614] = b[14] & g[21847];
assign g[38232] = a[14] & g[21848];
assign g[54615] = b[14] & g[21848];
assign g[38233] = a[14] & g[21849];
assign g[54616] = b[14] & g[21849];
assign g[38234] = a[14] & g[21850];
assign g[54617] = b[14] & g[21850];
assign g[38235] = a[14] & g[21851];
assign g[54618] = b[14] & g[21851];
assign g[38236] = a[14] & g[21852];
assign g[54619] = b[14] & g[21852];
assign g[38237] = a[14] & g[21853];
assign g[54620] = b[14] & g[21853];
assign g[38238] = a[14] & g[21854];
assign g[54621] = b[14] & g[21854];
assign g[38239] = a[14] & g[21855];
assign g[54622] = b[14] & g[21855];
assign g[38240] = a[14] & g[21856];
assign g[54623] = b[14] & g[21856];
assign g[38241] = a[14] & g[21857];
assign g[54624] = b[14] & g[21857];
assign g[38242] = a[14] & g[21858];
assign g[54625] = b[14] & g[21858];
assign g[38243] = a[14] & g[21859];
assign g[54626] = b[14] & g[21859];
assign g[38244] = a[14] & g[21860];
assign g[54627] = b[14] & g[21860];
assign g[38245] = a[14] & g[21861];
assign g[54628] = b[14] & g[21861];
assign g[38246] = a[14] & g[21862];
assign g[54629] = b[14] & g[21862];
assign g[38247] = a[14] & g[21863];
assign g[54630] = b[14] & g[21863];
assign g[38248] = a[14] & g[21864];
assign g[54631] = b[14] & g[21864];
assign g[38249] = a[14] & g[21865];
assign g[54632] = b[14] & g[21865];
assign g[38250] = a[14] & g[21866];
assign g[54633] = b[14] & g[21866];
assign g[38251] = a[14] & g[21867];
assign g[54634] = b[14] & g[21867];
assign g[38252] = a[14] & g[21868];
assign g[54635] = b[14] & g[21868];
assign g[38253] = a[14] & g[21869];
assign g[54636] = b[14] & g[21869];
assign g[38254] = a[14] & g[21870];
assign g[54637] = b[14] & g[21870];
assign g[38255] = a[14] & g[21871];
assign g[54638] = b[14] & g[21871];
assign g[38256] = a[14] & g[21872];
assign g[54639] = b[14] & g[21872];
assign g[38257] = a[14] & g[21873];
assign g[54640] = b[14] & g[21873];
assign g[38258] = a[14] & g[21874];
assign g[54641] = b[14] & g[21874];
assign g[38259] = a[14] & g[21875];
assign g[54642] = b[14] & g[21875];
assign g[38260] = a[14] & g[21876];
assign g[54643] = b[14] & g[21876];
assign g[38261] = a[14] & g[21877];
assign g[54644] = b[14] & g[21877];
assign g[38262] = a[14] & g[21878];
assign g[54645] = b[14] & g[21878];
assign g[38263] = a[14] & g[21879];
assign g[54646] = b[14] & g[21879];
assign g[38264] = a[14] & g[21880];
assign g[54647] = b[14] & g[21880];
assign g[38265] = a[14] & g[21881];
assign g[54648] = b[14] & g[21881];
assign g[38266] = a[14] & g[21882];
assign g[54649] = b[14] & g[21882];
assign g[38267] = a[14] & g[21883];
assign g[54650] = b[14] & g[21883];
assign g[38268] = a[14] & g[21884];
assign g[54651] = b[14] & g[21884];
assign g[38269] = a[14] & g[21885];
assign g[54652] = b[14] & g[21885];
assign g[38270] = a[14] & g[21886];
assign g[54653] = b[14] & g[21886];
assign g[38271] = a[14] & g[21887];
assign g[54654] = b[14] & g[21887];
assign g[38272] = a[14] & g[21888];
assign g[54655] = b[14] & g[21888];
assign g[38273] = a[14] & g[21889];
assign g[54656] = b[14] & g[21889];
assign g[38274] = a[14] & g[21890];
assign g[54657] = b[14] & g[21890];
assign g[38275] = a[14] & g[21891];
assign g[54658] = b[14] & g[21891];
assign g[38276] = a[14] & g[21892];
assign g[54659] = b[14] & g[21892];
assign g[38277] = a[14] & g[21893];
assign g[54660] = b[14] & g[21893];
assign g[38278] = a[14] & g[21894];
assign g[54661] = b[14] & g[21894];
assign g[38279] = a[14] & g[21895];
assign g[54662] = b[14] & g[21895];
assign g[38280] = a[14] & g[21896];
assign g[54663] = b[14] & g[21896];
assign g[38281] = a[14] & g[21897];
assign g[54664] = b[14] & g[21897];
assign g[38282] = a[14] & g[21898];
assign g[54665] = b[14] & g[21898];
assign g[38283] = a[14] & g[21899];
assign g[54666] = b[14] & g[21899];
assign g[38284] = a[14] & g[21900];
assign g[54667] = b[14] & g[21900];
assign g[38285] = a[14] & g[21901];
assign g[54668] = b[14] & g[21901];
assign g[38286] = a[14] & g[21902];
assign g[54669] = b[14] & g[21902];
assign g[38287] = a[14] & g[21903];
assign g[54670] = b[14] & g[21903];
assign g[38288] = a[14] & g[21904];
assign g[54671] = b[14] & g[21904];
assign g[38289] = a[14] & g[21905];
assign g[54672] = b[14] & g[21905];
assign g[38290] = a[14] & g[21906];
assign g[54673] = b[14] & g[21906];
assign g[38291] = a[14] & g[21907];
assign g[54674] = b[14] & g[21907];
assign g[38292] = a[14] & g[21908];
assign g[54675] = b[14] & g[21908];
assign g[38293] = a[14] & g[21909];
assign g[54676] = b[14] & g[21909];
assign g[38294] = a[14] & g[21910];
assign g[54677] = b[14] & g[21910];
assign g[38295] = a[14] & g[21911];
assign g[54678] = b[14] & g[21911];
assign g[38296] = a[14] & g[21912];
assign g[54679] = b[14] & g[21912];
assign g[38297] = a[14] & g[21913];
assign g[54680] = b[14] & g[21913];
assign g[38298] = a[14] & g[21914];
assign g[54681] = b[14] & g[21914];
assign g[38299] = a[14] & g[21915];
assign g[54682] = b[14] & g[21915];
assign g[38300] = a[14] & g[21916];
assign g[54683] = b[14] & g[21916];
assign g[38301] = a[14] & g[21917];
assign g[54684] = b[14] & g[21917];
assign g[38302] = a[14] & g[21918];
assign g[54685] = b[14] & g[21918];
assign g[38303] = a[14] & g[21919];
assign g[54686] = b[14] & g[21919];
assign g[38304] = a[14] & g[21920];
assign g[54687] = b[14] & g[21920];
assign g[38305] = a[14] & g[21921];
assign g[54688] = b[14] & g[21921];
assign g[38306] = a[14] & g[21922];
assign g[54689] = b[14] & g[21922];
assign g[38307] = a[14] & g[21923];
assign g[54690] = b[14] & g[21923];
assign g[38308] = a[14] & g[21924];
assign g[54691] = b[14] & g[21924];
assign g[38309] = a[14] & g[21925];
assign g[54692] = b[14] & g[21925];
assign g[38310] = a[14] & g[21926];
assign g[54693] = b[14] & g[21926];
assign g[38311] = a[14] & g[21927];
assign g[54694] = b[14] & g[21927];
assign g[38312] = a[14] & g[21928];
assign g[54695] = b[14] & g[21928];
assign g[38313] = a[14] & g[21929];
assign g[54696] = b[14] & g[21929];
assign g[38314] = a[14] & g[21930];
assign g[54697] = b[14] & g[21930];
assign g[38315] = a[14] & g[21931];
assign g[54698] = b[14] & g[21931];
assign g[38316] = a[14] & g[21932];
assign g[54699] = b[14] & g[21932];
assign g[38317] = a[14] & g[21933];
assign g[54700] = b[14] & g[21933];
assign g[38318] = a[14] & g[21934];
assign g[54701] = b[14] & g[21934];
assign g[38319] = a[14] & g[21935];
assign g[54702] = b[14] & g[21935];
assign g[38320] = a[14] & g[21936];
assign g[54703] = b[14] & g[21936];
assign g[38321] = a[14] & g[21937];
assign g[54704] = b[14] & g[21937];
assign g[38322] = a[14] & g[21938];
assign g[54705] = b[14] & g[21938];
assign g[38323] = a[14] & g[21939];
assign g[54706] = b[14] & g[21939];
assign g[38324] = a[14] & g[21940];
assign g[54707] = b[14] & g[21940];
assign g[38325] = a[14] & g[21941];
assign g[54708] = b[14] & g[21941];
assign g[38326] = a[14] & g[21942];
assign g[54709] = b[14] & g[21942];
assign g[38327] = a[14] & g[21943];
assign g[54710] = b[14] & g[21943];
assign g[38328] = a[14] & g[21944];
assign g[54711] = b[14] & g[21944];
assign g[38329] = a[14] & g[21945];
assign g[54712] = b[14] & g[21945];
assign g[38330] = a[14] & g[21946];
assign g[54713] = b[14] & g[21946];
assign g[38331] = a[14] & g[21947];
assign g[54714] = b[14] & g[21947];
assign g[38332] = a[14] & g[21948];
assign g[54715] = b[14] & g[21948];
assign g[38333] = a[14] & g[21949];
assign g[54716] = b[14] & g[21949];
assign g[38334] = a[14] & g[21950];
assign g[54717] = b[14] & g[21950];
assign g[38335] = a[14] & g[21951];
assign g[54718] = b[14] & g[21951];
assign g[38336] = a[14] & g[21952];
assign g[54719] = b[14] & g[21952];
assign g[38337] = a[14] & g[21953];
assign g[54720] = b[14] & g[21953];
assign g[38338] = a[14] & g[21954];
assign g[54721] = b[14] & g[21954];
assign g[38339] = a[14] & g[21955];
assign g[54722] = b[14] & g[21955];
assign g[38340] = a[14] & g[21956];
assign g[54723] = b[14] & g[21956];
assign g[38341] = a[14] & g[21957];
assign g[54724] = b[14] & g[21957];
assign g[38342] = a[14] & g[21958];
assign g[54725] = b[14] & g[21958];
assign g[38343] = a[14] & g[21959];
assign g[54726] = b[14] & g[21959];
assign g[38344] = a[14] & g[21960];
assign g[54727] = b[14] & g[21960];
assign g[38345] = a[14] & g[21961];
assign g[54728] = b[14] & g[21961];
assign g[38346] = a[14] & g[21962];
assign g[54729] = b[14] & g[21962];
assign g[38347] = a[14] & g[21963];
assign g[54730] = b[14] & g[21963];
assign g[38348] = a[14] & g[21964];
assign g[54731] = b[14] & g[21964];
assign g[38349] = a[14] & g[21965];
assign g[54732] = b[14] & g[21965];
assign g[38350] = a[14] & g[21966];
assign g[54733] = b[14] & g[21966];
assign g[38351] = a[14] & g[21967];
assign g[54734] = b[14] & g[21967];
assign g[38352] = a[14] & g[21968];
assign g[54735] = b[14] & g[21968];
assign g[38353] = a[14] & g[21969];
assign g[54736] = b[14] & g[21969];
assign g[38354] = a[14] & g[21970];
assign g[54737] = b[14] & g[21970];
assign g[38355] = a[14] & g[21971];
assign g[54738] = b[14] & g[21971];
assign g[38356] = a[14] & g[21972];
assign g[54739] = b[14] & g[21972];
assign g[38357] = a[14] & g[21973];
assign g[54740] = b[14] & g[21973];
assign g[38358] = a[14] & g[21974];
assign g[54741] = b[14] & g[21974];
assign g[38359] = a[14] & g[21975];
assign g[54742] = b[14] & g[21975];
assign g[38360] = a[14] & g[21976];
assign g[54743] = b[14] & g[21976];
assign g[38361] = a[14] & g[21977];
assign g[54744] = b[14] & g[21977];
assign g[38362] = a[14] & g[21978];
assign g[54745] = b[14] & g[21978];
assign g[38363] = a[14] & g[21979];
assign g[54746] = b[14] & g[21979];
assign g[38364] = a[14] & g[21980];
assign g[54747] = b[14] & g[21980];
assign g[38365] = a[14] & g[21981];
assign g[54748] = b[14] & g[21981];
assign g[38366] = a[14] & g[21982];
assign g[54749] = b[14] & g[21982];
assign g[38367] = a[14] & g[21983];
assign g[54750] = b[14] & g[21983];
assign g[38368] = a[14] & g[21984];
assign g[54751] = b[14] & g[21984];
assign g[38369] = a[14] & g[21985];
assign g[54752] = b[14] & g[21985];
assign g[38370] = a[14] & g[21986];
assign g[54753] = b[14] & g[21986];
assign g[38371] = a[14] & g[21987];
assign g[54754] = b[14] & g[21987];
assign g[38372] = a[14] & g[21988];
assign g[54755] = b[14] & g[21988];
assign g[38373] = a[14] & g[21989];
assign g[54756] = b[14] & g[21989];
assign g[38374] = a[14] & g[21990];
assign g[54757] = b[14] & g[21990];
assign g[38375] = a[14] & g[21991];
assign g[54758] = b[14] & g[21991];
assign g[38376] = a[14] & g[21992];
assign g[54759] = b[14] & g[21992];
assign g[38377] = a[14] & g[21993];
assign g[54760] = b[14] & g[21993];
assign g[38378] = a[14] & g[21994];
assign g[54761] = b[14] & g[21994];
assign g[38379] = a[14] & g[21995];
assign g[54762] = b[14] & g[21995];
assign g[38380] = a[14] & g[21996];
assign g[54763] = b[14] & g[21996];
assign g[38381] = a[14] & g[21997];
assign g[54764] = b[14] & g[21997];
assign g[38382] = a[14] & g[21998];
assign g[54765] = b[14] & g[21998];
assign g[38383] = a[14] & g[21999];
assign g[54766] = b[14] & g[21999];
assign g[38384] = a[14] & g[22000];
assign g[54767] = b[14] & g[22000];
assign g[38385] = a[14] & g[22001];
assign g[54768] = b[14] & g[22001];
assign g[38386] = a[14] & g[22002];
assign g[54769] = b[14] & g[22002];
assign g[38387] = a[14] & g[22003];
assign g[54770] = b[14] & g[22003];
assign g[38388] = a[14] & g[22004];
assign g[54771] = b[14] & g[22004];
assign g[38389] = a[14] & g[22005];
assign g[54772] = b[14] & g[22005];
assign g[38390] = a[14] & g[22006];
assign g[54773] = b[14] & g[22006];
assign g[38391] = a[14] & g[22007];
assign g[54774] = b[14] & g[22007];
assign g[38392] = a[14] & g[22008];
assign g[54775] = b[14] & g[22008];
assign g[38393] = a[14] & g[22009];
assign g[54776] = b[14] & g[22009];
assign g[38394] = a[14] & g[22010];
assign g[54777] = b[14] & g[22010];
assign g[38395] = a[14] & g[22011];
assign g[54778] = b[14] & g[22011];
assign g[38396] = a[14] & g[22012];
assign g[54779] = b[14] & g[22012];
assign g[38397] = a[14] & g[22013];
assign g[54780] = b[14] & g[22013];
assign g[38398] = a[14] & g[22014];
assign g[54781] = b[14] & g[22014];
assign g[38399] = a[14] & g[22015];
assign g[54782] = b[14] & g[22015];
assign g[38400] = a[14] & g[22016];
assign g[54783] = b[14] & g[22016];
assign g[38401] = a[14] & g[22017];
assign g[54784] = b[14] & g[22017];
assign g[38402] = a[14] & g[22018];
assign g[54785] = b[14] & g[22018];
assign g[38403] = a[14] & g[22019];
assign g[54786] = b[14] & g[22019];
assign g[38404] = a[14] & g[22020];
assign g[54787] = b[14] & g[22020];
assign g[38405] = a[14] & g[22021];
assign g[54788] = b[14] & g[22021];
assign g[38406] = a[14] & g[22022];
assign g[54789] = b[14] & g[22022];
assign g[38407] = a[14] & g[22023];
assign g[54790] = b[14] & g[22023];
assign g[38408] = a[14] & g[22024];
assign g[54791] = b[14] & g[22024];
assign g[38409] = a[14] & g[22025];
assign g[54792] = b[14] & g[22025];
assign g[38410] = a[14] & g[22026];
assign g[54793] = b[14] & g[22026];
assign g[38411] = a[14] & g[22027];
assign g[54794] = b[14] & g[22027];
assign g[38412] = a[14] & g[22028];
assign g[54795] = b[14] & g[22028];
assign g[38413] = a[14] & g[22029];
assign g[54796] = b[14] & g[22029];
assign g[38414] = a[14] & g[22030];
assign g[54797] = b[14] & g[22030];
assign g[38415] = a[14] & g[22031];
assign g[54798] = b[14] & g[22031];
assign g[38416] = a[14] & g[22032];
assign g[54799] = b[14] & g[22032];
assign g[38417] = a[14] & g[22033];
assign g[54800] = b[14] & g[22033];
assign g[38418] = a[14] & g[22034];
assign g[54801] = b[14] & g[22034];
assign g[38419] = a[14] & g[22035];
assign g[54802] = b[14] & g[22035];
assign g[38420] = a[14] & g[22036];
assign g[54803] = b[14] & g[22036];
assign g[38421] = a[14] & g[22037];
assign g[54804] = b[14] & g[22037];
assign g[38422] = a[14] & g[22038];
assign g[54805] = b[14] & g[22038];
assign g[38423] = a[14] & g[22039];
assign g[54806] = b[14] & g[22039];
assign g[38424] = a[14] & g[22040];
assign g[54807] = b[14] & g[22040];
assign g[38425] = a[14] & g[22041];
assign g[54808] = b[14] & g[22041];
assign g[38426] = a[14] & g[22042];
assign g[54809] = b[14] & g[22042];
assign g[38427] = a[14] & g[22043];
assign g[54810] = b[14] & g[22043];
assign g[38428] = a[14] & g[22044];
assign g[54811] = b[14] & g[22044];
assign g[38429] = a[14] & g[22045];
assign g[54812] = b[14] & g[22045];
assign g[38430] = a[14] & g[22046];
assign g[54813] = b[14] & g[22046];
assign g[38431] = a[14] & g[22047];
assign g[54814] = b[14] & g[22047];
assign g[38432] = a[14] & g[22048];
assign g[54815] = b[14] & g[22048];
assign g[38433] = a[14] & g[22049];
assign g[54816] = b[14] & g[22049];
assign g[38434] = a[14] & g[22050];
assign g[54817] = b[14] & g[22050];
assign g[38435] = a[14] & g[22051];
assign g[54818] = b[14] & g[22051];
assign g[38436] = a[14] & g[22052];
assign g[54819] = b[14] & g[22052];
assign g[38437] = a[14] & g[22053];
assign g[54820] = b[14] & g[22053];
assign g[38438] = a[14] & g[22054];
assign g[54821] = b[14] & g[22054];
assign g[38439] = a[14] & g[22055];
assign g[54822] = b[14] & g[22055];
assign g[38440] = a[14] & g[22056];
assign g[54823] = b[14] & g[22056];
assign g[38441] = a[14] & g[22057];
assign g[54824] = b[14] & g[22057];
assign g[38442] = a[14] & g[22058];
assign g[54825] = b[14] & g[22058];
assign g[38443] = a[14] & g[22059];
assign g[54826] = b[14] & g[22059];
assign g[38444] = a[14] & g[22060];
assign g[54827] = b[14] & g[22060];
assign g[38445] = a[14] & g[22061];
assign g[54828] = b[14] & g[22061];
assign g[38446] = a[14] & g[22062];
assign g[54829] = b[14] & g[22062];
assign g[38447] = a[14] & g[22063];
assign g[54830] = b[14] & g[22063];
assign g[38448] = a[14] & g[22064];
assign g[54831] = b[14] & g[22064];
assign g[38449] = a[14] & g[22065];
assign g[54832] = b[14] & g[22065];
assign g[38450] = a[14] & g[22066];
assign g[54833] = b[14] & g[22066];
assign g[38451] = a[14] & g[22067];
assign g[54834] = b[14] & g[22067];
assign g[38452] = a[14] & g[22068];
assign g[54835] = b[14] & g[22068];
assign g[38453] = a[14] & g[22069];
assign g[54836] = b[14] & g[22069];
assign g[38454] = a[14] & g[22070];
assign g[54837] = b[14] & g[22070];
assign g[38455] = a[14] & g[22071];
assign g[54838] = b[14] & g[22071];
assign g[38456] = a[14] & g[22072];
assign g[54839] = b[14] & g[22072];
assign g[38457] = a[14] & g[22073];
assign g[54840] = b[14] & g[22073];
assign g[38458] = a[14] & g[22074];
assign g[54841] = b[14] & g[22074];
assign g[38459] = a[14] & g[22075];
assign g[54842] = b[14] & g[22075];
assign g[38460] = a[14] & g[22076];
assign g[54843] = b[14] & g[22076];
assign g[38461] = a[14] & g[22077];
assign g[54844] = b[14] & g[22077];
assign g[38462] = a[14] & g[22078];
assign g[54845] = b[14] & g[22078];
assign g[38463] = a[14] & g[22079];
assign g[54846] = b[14] & g[22079];
assign g[38464] = a[14] & g[22080];
assign g[54847] = b[14] & g[22080];
assign g[38465] = a[14] & g[22081];
assign g[54848] = b[14] & g[22081];
assign g[38466] = a[14] & g[22082];
assign g[54849] = b[14] & g[22082];
assign g[38467] = a[14] & g[22083];
assign g[54850] = b[14] & g[22083];
assign g[38468] = a[14] & g[22084];
assign g[54851] = b[14] & g[22084];
assign g[38469] = a[14] & g[22085];
assign g[54852] = b[14] & g[22085];
assign g[38470] = a[14] & g[22086];
assign g[54853] = b[14] & g[22086];
assign g[38471] = a[14] & g[22087];
assign g[54854] = b[14] & g[22087];
assign g[38472] = a[14] & g[22088];
assign g[54855] = b[14] & g[22088];
assign g[38473] = a[14] & g[22089];
assign g[54856] = b[14] & g[22089];
assign g[38474] = a[14] & g[22090];
assign g[54857] = b[14] & g[22090];
assign g[38475] = a[14] & g[22091];
assign g[54858] = b[14] & g[22091];
assign g[38476] = a[14] & g[22092];
assign g[54859] = b[14] & g[22092];
assign g[38477] = a[14] & g[22093];
assign g[54860] = b[14] & g[22093];
assign g[38478] = a[14] & g[22094];
assign g[54861] = b[14] & g[22094];
assign g[38479] = a[14] & g[22095];
assign g[54862] = b[14] & g[22095];
assign g[38480] = a[14] & g[22096];
assign g[54863] = b[14] & g[22096];
assign g[38481] = a[14] & g[22097];
assign g[54864] = b[14] & g[22097];
assign g[38482] = a[14] & g[22098];
assign g[54865] = b[14] & g[22098];
assign g[38483] = a[14] & g[22099];
assign g[54866] = b[14] & g[22099];
assign g[38484] = a[14] & g[22100];
assign g[54867] = b[14] & g[22100];
assign g[38485] = a[14] & g[22101];
assign g[54868] = b[14] & g[22101];
assign g[38486] = a[14] & g[22102];
assign g[54869] = b[14] & g[22102];
assign g[38487] = a[14] & g[22103];
assign g[54870] = b[14] & g[22103];
assign g[38488] = a[14] & g[22104];
assign g[54871] = b[14] & g[22104];
assign g[38489] = a[14] & g[22105];
assign g[54872] = b[14] & g[22105];
assign g[38490] = a[14] & g[22106];
assign g[54873] = b[14] & g[22106];
assign g[38491] = a[14] & g[22107];
assign g[54874] = b[14] & g[22107];
assign g[38492] = a[14] & g[22108];
assign g[54875] = b[14] & g[22108];
assign g[38493] = a[14] & g[22109];
assign g[54876] = b[14] & g[22109];
assign g[38494] = a[14] & g[22110];
assign g[54877] = b[14] & g[22110];
assign g[38495] = a[14] & g[22111];
assign g[54878] = b[14] & g[22111];
assign g[38496] = a[14] & g[22112];
assign g[54879] = b[14] & g[22112];
assign g[38497] = a[14] & g[22113];
assign g[54880] = b[14] & g[22113];
assign g[38498] = a[14] & g[22114];
assign g[54881] = b[14] & g[22114];
assign g[38499] = a[14] & g[22115];
assign g[54882] = b[14] & g[22115];
assign g[38500] = a[14] & g[22116];
assign g[54883] = b[14] & g[22116];
assign g[38501] = a[14] & g[22117];
assign g[54884] = b[14] & g[22117];
assign g[38502] = a[14] & g[22118];
assign g[54885] = b[14] & g[22118];
assign g[38503] = a[14] & g[22119];
assign g[54886] = b[14] & g[22119];
assign g[38504] = a[14] & g[22120];
assign g[54887] = b[14] & g[22120];
assign g[38505] = a[14] & g[22121];
assign g[54888] = b[14] & g[22121];
assign g[38506] = a[14] & g[22122];
assign g[54889] = b[14] & g[22122];
assign g[38507] = a[14] & g[22123];
assign g[54890] = b[14] & g[22123];
assign g[38508] = a[14] & g[22124];
assign g[54891] = b[14] & g[22124];
assign g[38509] = a[14] & g[22125];
assign g[54892] = b[14] & g[22125];
assign g[38510] = a[14] & g[22126];
assign g[54893] = b[14] & g[22126];
assign g[38511] = a[14] & g[22127];
assign g[54894] = b[14] & g[22127];
assign g[38512] = a[14] & g[22128];
assign g[54895] = b[14] & g[22128];
assign g[38513] = a[14] & g[22129];
assign g[54896] = b[14] & g[22129];
assign g[38514] = a[14] & g[22130];
assign g[54897] = b[14] & g[22130];
assign g[38515] = a[14] & g[22131];
assign g[54898] = b[14] & g[22131];
assign g[38516] = a[14] & g[22132];
assign g[54899] = b[14] & g[22132];
assign g[38517] = a[14] & g[22133];
assign g[54900] = b[14] & g[22133];
assign g[38518] = a[14] & g[22134];
assign g[54901] = b[14] & g[22134];
assign g[38519] = a[14] & g[22135];
assign g[54902] = b[14] & g[22135];
assign g[38520] = a[14] & g[22136];
assign g[54903] = b[14] & g[22136];
assign g[38521] = a[14] & g[22137];
assign g[54904] = b[14] & g[22137];
assign g[38522] = a[14] & g[22138];
assign g[54905] = b[14] & g[22138];
assign g[38523] = a[14] & g[22139];
assign g[54906] = b[14] & g[22139];
assign g[38524] = a[14] & g[22140];
assign g[54907] = b[14] & g[22140];
assign g[38525] = a[14] & g[22141];
assign g[54908] = b[14] & g[22141];
assign g[38526] = a[14] & g[22142];
assign g[54909] = b[14] & g[22142];
assign g[38527] = a[14] & g[22143];
assign g[54910] = b[14] & g[22143];
assign g[38528] = a[14] & g[22144];
assign g[54911] = b[14] & g[22144];
assign g[38529] = a[14] & g[22145];
assign g[54912] = b[14] & g[22145];
assign g[38530] = a[14] & g[22146];
assign g[54913] = b[14] & g[22146];
assign g[38531] = a[14] & g[22147];
assign g[54914] = b[14] & g[22147];
assign g[38532] = a[14] & g[22148];
assign g[54915] = b[14] & g[22148];
assign g[38533] = a[14] & g[22149];
assign g[54916] = b[14] & g[22149];
assign g[38534] = a[14] & g[22150];
assign g[54917] = b[14] & g[22150];
assign g[38535] = a[14] & g[22151];
assign g[54918] = b[14] & g[22151];
assign g[38536] = a[14] & g[22152];
assign g[54919] = b[14] & g[22152];
assign g[38537] = a[14] & g[22153];
assign g[54920] = b[14] & g[22153];
assign g[38538] = a[14] & g[22154];
assign g[54921] = b[14] & g[22154];
assign g[38539] = a[14] & g[22155];
assign g[54922] = b[14] & g[22155];
assign g[38540] = a[14] & g[22156];
assign g[54923] = b[14] & g[22156];
assign g[38541] = a[14] & g[22157];
assign g[54924] = b[14] & g[22157];
assign g[38542] = a[14] & g[22158];
assign g[54925] = b[14] & g[22158];
assign g[38543] = a[14] & g[22159];
assign g[54926] = b[14] & g[22159];
assign g[38544] = a[14] & g[22160];
assign g[54927] = b[14] & g[22160];
assign g[38545] = a[14] & g[22161];
assign g[54928] = b[14] & g[22161];
assign g[38546] = a[14] & g[22162];
assign g[54929] = b[14] & g[22162];
assign g[38547] = a[14] & g[22163];
assign g[54930] = b[14] & g[22163];
assign g[38548] = a[14] & g[22164];
assign g[54931] = b[14] & g[22164];
assign g[38549] = a[14] & g[22165];
assign g[54932] = b[14] & g[22165];
assign g[38550] = a[14] & g[22166];
assign g[54933] = b[14] & g[22166];
assign g[38551] = a[14] & g[22167];
assign g[54934] = b[14] & g[22167];
assign g[38552] = a[14] & g[22168];
assign g[54935] = b[14] & g[22168];
assign g[38553] = a[14] & g[22169];
assign g[54936] = b[14] & g[22169];
assign g[38554] = a[14] & g[22170];
assign g[54937] = b[14] & g[22170];
assign g[38555] = a[14] & g[22171];
assign g[54938] = b[14] & g[22171];
assign g[38556] = a[14] & g[22172];
assign g[54939] = b[14] & g[22172];
assign g[38557] = a[14] & g[22173];
assign g[54940] = b[14] & g[22173];
assign g[38558] = a[14] & g[22174];
assign g[54941] = b[14] & g[22174];
assign g[38559] = a[14] & g[22175];
assign g[54942] = b[14] & g[22175];
assign g[38560] = a[14] & g[22176];
assign g[54943] = b[14] & g[22176];
assign g[38561] = a[14] & g[22177];
assign g[54944] = b[14] & g[22177];
assign g[38562] = a[14] & g[22178];
assign g[54945] = b[14] & g[22178];
assign g[38563] = a[14] & g[22179];
assign g[54946] = b[14] & g[22179];
assign g[38564] = a[14] & g[22180];
assign g[54947] = b[14] & g[22180];
assign g[38565] = a[14] & g[22181];
assign g[54948] = b[14] & g[22181];
assign g[38566] = a[14] & g[22182];
assign g[54949] = b[14] & g[22182];
assign g[38567] = a[14] & g[22183];
assign g[54950] = b[14] & g[22183];
assign g[38568] = a[14] & g[22184];
assign g[54951] = b[14] & g[22184];
assign g[38569] = a[14] & g[22185];
assign g[54952] = b[14] & g[22185];
assign g[38570] = a[14] & g[22186];
assign g[54953] = b[14] & g[22186];
assign g[38571] = a[14] & g[22187];
assign g[54954] = b[14] & g[22187];
assign g[38572] = a[14] & g[22188];
assign g[54955] = b[14] & g[22188];
assign g[38573] = a[14] & g[22189];
assign g[54956] = b[14] & g[22189];
assign g[38574] = a[14] & g[22190];
assign g[54957] = b[14] & g[22190];
assign g[38575] = a[14] & g[22191];
assign g[54958] = b[14] & g[22191];
assign g[38576] = a[14] & g[22192];
assign g[54959] = b[14] & g[22192];
assign g[38577] = a[14] & g[22193];
assign g[54960] = b[14] & g[22193];
assign g[38578] = a[14] & g[22194];
assign g[54961] = b[14] & g[22194];
assign g[38579] = a[14] & g[22195];
assign g[54962] = b[14] & g[22195];
assign g[38580] = a[14] & g[22196];
assign g[54963] = b[14] & g[22196];
assign g[38581] = a[14] & g[22197];
assign g[54964] = b[14] & g[22197];
assign g[38582] = a[14] & g[22198];
assign g[54965] = b[14] & g[22198];
assign g[38583] = a[14] & g[22199];
assign g[54966] = b[14] & g[22199];
assign g[38584] = a[14] & g[22200];
assign g[54967] = b[14] & g[22200];
assign g[38585] = a[14] & g[22201];
assign g[54968] = b[14] & g[22201];
assign g[38586] = a[14] & g[22202];
assign g[54969] = b[14] & g[22202];
assign g[38587] = a[14] & g[22203];
assign g[54970] = b[14] & g[22203];
assign g[38588] = a[14] & g[22204];
assign g[54971] = b[14] & g[22204];
assign g[38589] = a[14] & g[22205];
assign g[54972] = b[14] & g[22205];
assign g[38590] = a[14] & g[22206];
assign g[54973] = b[14] & g[22206];
assign g[38591] = a[14] & g[22207];
assign g[54974] = b[14] & g[22207];
assign g[38592] = a[14] & g[22208];
assign g[54975] = b[14] & g[22208];
assign g[38593] = a[14] & g[22209];
assign g[54976] = b[14] & g[22209];
assign g[38594] = a[14] & g[22210];
assign g[54977] = b[14] & g[22210];
assign g[38595] = a[14] & g[22211];
assign g[54978] = b[14] & g[22211];
assign g[38596] = a[14] & g[22212];
assign g[54979] = b[14] & g[22212];
assign g[38597] = a[14] & g[22213];
assign g[54980] = b[14] & g[22213];
assign g[38598] = a[14] & g[22214];
assign g[54981] = b[14] & g[22214];
assign g[38599] = a[14] & g[22215];
assign g[54982] = b[14] & g[22215];
assign g[38600] = a[14] & g[22216];
assign g[54983] = b[14] & g[22216];
assign g[38601] = a[14] & g[22217];
assign g[54984] = b[14] & g[22217];
assign g[38602] = a[14] & g[22218];
assign g[54985] = b[14] & g[22218];
assign g[38603] = a[14] & g[22219];
assign g[54986] = b[14] & g[22219];
assign g[38604] = a[14] & g[22220];
assign g[54987] = b[14] & g[22220];
assign g[38605] = a[14] & g[22221];
assign g[54988] = b[14] & g[22221];
assign g[38606] = a[14] & g[22222];
assign g[54989] = b[14] & g[22222];
assign g[38607] = a[14] & g[22223];
assign g[54990] = b[14] & g[22223];
assign g[38608] = a[14] & g[22224];
assign g[54991] = b[14] & g[22224];
assign g[38609] = a[14] & g[22225];
assign g[54992] = b[14] & g[22225];
assign g[38610] = a[14] & g[22226];
assign g[54993] = b[14] & g[22226];
assign g[38611] = a[14] & g[22227];
assign g[54994] = b[14] & g[22227];
assign g[38612] = a[14] & g[22228];
assign g[54995] = b[14] & g[22228];
assign g[38613] = a[14] & g[22229];
assign g[54996] = b[14] & g[22229];
assign g[38614] = a[14] & g[22230];
assign g[54997] = b[14] & g[22230];
assign g[38615] = a[14] & g[22231];
assign g[54998] = b[14] & g[22231];
assign g[38616] = a[14] & g[22232];
assign g[54999] = b[14] & g[22232];
assign g[38617] = a[14] & g[22233];
assign g[55000] = b[14] & g[22233];
assign g[38618] = a[14] & g[22234];
assign g[55001] = b[14] & g[22234];
assign g[38619] = a[14] & g[22235];
assign g[55002] = b[14] & g[22235];
assign g[38620] = a[14] & g[22236];
assign g[55003] = b[14] & g[22236];
assign g[38621] = a[14] & g[22237];
assign g[55004] = b[14] & g[22237];
assign g[38622] = a[14] & g[22238];
assign g[55005] = b[14] & g[22238];
assign g[38623] = a[14] & g[22239];
assign g[55006] = b[14] & g[22239];
assign g[38624] = a[14] & g[22240];
assign g[55007] = b[14] & g[22240];
assign g[38625] = a[14] & g[22241];
assign g[55008] = b[14] & g[22241];
assign g[38626] = a[14] & g[22242];
assign g[55009] = b[14] & g[22242];
assign g[38627] = a[14] & g[22243];
assign g[55010] = b[14] & g[22243];
assign g[38628] = a[14] & g[22244];
assign g[55011] = b[14] & g[22244];
assign g[38629] = a[14] & g[22245];
assign g[55012] = b[14] & g[22245];
assign g[38630] = a[14] & g[22246];
assign g[55013] = b[14] & g[22246];
assign g[38631] = a[14] & g[22247];
assign g[55014] = b[14] & g[22247];
assign g[38632] = a[14] & g[22248];
assign g[55015] = b[14] & g[22248];
assign g[38633] = a[14] & g[22249];
assign g[55016] = b[14] & g[22249];
assign g[38634] = a[14] & g[22250];
assign g[55017] = b[14] & g[22250];
assign g[38635] = a[14] & g[22251];
assign g[55018] = b[14] & g[22251];
assign g[38636] = a[14] & g[22252];
assign g[55019] = b[14] & g[22252];
assign g[38637] = a[14] & g[22253];
assign g[55020] = b[14] & g[22253];
assign g[38638] = a[14] & g[22254];
assign g[55021] = b[14] & g[22254];
assign g[38639] = a[14] & g[22255];
assign g[55022] = b[14] & g[22255];
assign g[38640] = a[14] & g[22256];
assign g[55023] = b[14] & g[22256];
assign g[38641] = a[14] & g[22257];
assign g[55024] = b[14] & g[22257];
assign g[38642] = a[14] & g[22258];
assign g[55025] = b[14] & g[22258];
assign g[38643] = a[14] & g[22259];
assign g[55026] = b[14] & g[22259];
assign g[38644] = a[14] & g[22260];
assign g[55027] = b[14] & g[22260];
assign g[38645] = a[14] & g[22261];
assign g[55028] = b[14] & g[22261];
assign g[38646] = a[14] & g[22262];
assign g[55029] = b[14] & g[22262];
assign g[38647] = a[14] & g[22263];
assign g[55030] = b[14] & g[22263];
assign g[38648] = a[14] & g[22264];
assign g[55031] = b[14] & g[22264];
assign g[38649] = a[14] & g[22265];
assign g[55032] = b[14] & g[22265];
assign g[38650] = a[14] & g[22266];
assign g[55033] = b[14] & g[22266];
assign g[38651] = a[14] & g[22267];
assign g[55034] = b[14] & g[22267];
assign g[38652] = a[14] & g[22268];
assign g[55035] = b[14] & g[22268];
assign g[38653] = a[14] & g[22269];
assign g[55036] = b[14] & g[22269];
assign g[38654] = a[14] & g[22270];
assign g[55037] = b[14] & g[22270];
assign g[38655] = a[14] & g[22271];
assign g[55038] = b[14] & g[22271];
assign g[38656] = a[14] & g[22272];
assign g[55039] = b[14] & g[22272];
assign g[38657] = a[14] & g[22273];
assign g[55040] = b[14] & g[22273];
assign g[38658] = a[14] & g[22274];
assign g[55041] = b[14] & g[22274];
assign g[38659] = a[14] & g[22275];
assign g[55042] = b[14] & g[22275];
assign g[38660] = a[14] & g[22276];
assign g[55043] = b[14] & g[22276];
assign g[38661] = a[14] & g[22277];
assign g[55044] = b[14] & g[22277];
assign g[38662] = a[14] & g[22278];
assign g[55045] = b[14] & g[22278];
assign g[38663] = a[14] & g[22279];
assign g[55046] = b[14] & g[22279];
assign g[38664] = a[14] & g[22280];
assign g[55047] = b[14] & g[22280];
assign g[38665] = a[14] & g[22281];
assign g[55048] = b[14] & g[22281];
assign g[38666] = a[14] & g[22282];
assign g[55049] = b[14] & g[22282];
assign g[38667] = a[14] & g[22283];
assign g[55050] = b[14] & g[22283];
assign g[38668] = a[14] & g[22284];
assign g[55051] = b[14] & g[22284];
assign g[38669] = a[14] & g[22285];
assign g[55052] = b[14] & g[22285];
assign g[38670] = a[14] & g[22286];
assign g[55053] = b[14] & g[22286];
assign g[38671] = a[14] & g[22287];
assign g[55054] = b[14] & g[22287];
assign g[38672] = a[14] & g[22288];
assign g[55055] = b[14] & g[22288];
assign g[38673] = a[14] & g[22289];
assign g[55056] = b[14] & g[22289];
assign g[38674] = a[14] & g[22290];
assign g[55057] = b[14] & g[22290];
assign g[38675] = a[14] & g[22291];
assign g[55058] = b[14] & g[22291];
assign g[38676] = a[14] & g[22292];
assign g[55059] = b[14] & g[22292];
assign g[38677] = a[14] & g[22293];
assign g[55060] = b[14] & g[22293];
assign g[38678] = a[14] & g[22294];
assign g[55061] = b[14] & g[22294];
assign g[38679] = a[14] & g[22295];
assign g[55062] = b[14] & g[22295];
assign g[38680] = a[14] & g[22296];
assign g[55063] = b[14] & g[22296];
assign g[38681] = a[14] & g[22297];
assign g[55064] = b[14] & g[22297];
assign g[38682] = a[14] & g[22298];
assign g[55065] = b[14] & g[22298];
assign g[38683] = a[14] & g[22299];
assign g[55066] = b[14] & g[22299];
assign g[38684] = a[14] & g[22300];
assign g[55067] = b[14] & g[22300];
assign g[38685] = a[14] & g[22301];
assign g[55068] = b[14] & g[22301];
assign g[38686] = a[14] & g[22302];
assign g[55069] = b[14] & g[22302];
assign g[38687] = a[14] & g[22303];
assign g[55070] = b[14] & g[22303];
assign g[38688] = a[14] & g[22304];
assign g[55071] = b[14] & g[22304];
assign g[38689] = a[14] & g[22305];
assign g[55072] = b[14] & g[22305];
assign g[38690] = a[14] & g[22306];
assign g[55073] = b[14] & g[22306];
assign g[38691] = a[14] & g[22307];
assign g[55074] = b[14] & g[22307];
assign g[38692] = a[14] & g[22308];
assign g[55075] = b[14] & g[22308];
assign g[38693] = a[14] & g[22309];
assign g[55076] = b[14] & g[22309];
assign g[38694] = a[14] & g[22310];
assign g[55077] = b[14] & g[22310];
assign g[38695] = a[14] & g[22311];
assign g[55078] = b[14] & g[22311];
assign g[38696] = a[14] & g[22312];
assign g[55079] = b[14] & g[22312];
assign g[38697] = a[14] & g[22313];
assign g[55080] = b[14] & g[22313];
assign g[38698] = a[14] & g[22314];
assign g[55081] = b[14] & g[22314];
assign g[38699] = a[14] & g[22315];
assign g[55082] = b[14] & g[22315];
assign g[38700] = a[14] & g[22316];
assign g[55083] = b[14] & g[22316];
assign g[38701] = a[14] & g[22317];
assign g[55084] = b[14] & g[22317];
assign g[38702] = a[14] & g[22318];
assign g[55085] = b[14] & g[22318];
assign g[38703] = a[14] & g[22319];
assign g[55086] = b[14] & g[22319];
assign g[38704] = a[14] & g[22320];
assign g[55087] = b[14] & g[22320];
assign g[38705] = a[14] & g[22321];
assign g[55088] = b[14] & g[22321];
assign g[38706] = a[14] & g[22322];
assign g[55089] = b[14] & g[22322];
assign g[38707] = a[14] & g[22323];
assign g[55090] = b[14] & g[22323];
assign g[38708] = a[14] & g[22324];
assign g[55091] = b[14] & g[22324];
assign g[38709] = a[14] & g[22325];
assign g[55092] = b[14] & g[22325];
assign g[38710] = a[14] & g[22326];
assign g[55093] = b[14] & g[22326];
assign g[38711] = a[14] & g[22327];
assign g[55094] = b[14] & g[22327];
assign g[38712] = a[14] & g[22328];
assign g[55095] = b[14] & g[22328];
assign g[38713] = a[14] & g[22329];
assign g[55096] = b[14] & g[22329];
assign g[38714] = a[14] & g[22330];
assign g[55097] = b[14] & g[22330];
assign g[38715] = a[14] & g[22331];
assign g[55098] = b[14] & g[22331];
assign g[38716] = a[14] & g[22332];
assign g[55099] = b[14] & g[22332];
assign g[38717] = a[14] & g[22333];
assign g[55100] = b[14] & g[22333];
assign g[38718] = a[14] & g[22334];
assign g[55101] = b[14] & g[22334];
assign g[38719] = a[14] & g[22335];
assign g[55102] = b[14] & g[22335];
assign g[38720] = a[14] & g[22336];
assign g[55103] = b[14] & g[22336];
assign g[38721] = a[14] & g[22337];
assign g[55104] = b[14] & g[22337];
assign g[38722] = a[14] & g[22338];
assign g[55105] = b[14] & g[22338];
assign g[38723] = a[14] & g[22339];
assign g[55106] = b[14] & g[22339];
assign g[38724] = a[14] & g[22340];
assign g[55107] = b[14] & g[22340];
assign g[38725] = a[14] & g[22341];
assign g[55108] = b[14] & g[22341];
assign g[38726] = a[14] & g[22342];
assign g[55109] = b[14] & g[22342];
assign g[38727] = a[14] & g[22343];
assign g[55110] = b[14] & g[22343];
assign g[38728] = a[14] & g[22344];
assign g[55111] = b[14] & g[22344];
assign g[38729] = a[14] & g[22345];
assign g[55112] = b[14] & g[22345];
assign g[38730] = a[14] & g[22346];
assign g[55113] = b[14] & g[22346];
assign g[38731] = a[14] & g[22347];
assign g[55114] = b[14] & g[22347];
assign g[38732] = a[14] & g[22348];
assign g[55115] = b[14] & g[22348];
assign g[38733] = a[14] & g[22349];
assign g[55116] = b[14] & g[22349];
assign g[38734] = a[14] & g[22350];
assign g[55117] = b[14] & g[22350];
assign g[38735] = a[14] & g[22351];
assign g[55118] = b[14] & g[22351];
assign g[38736] = a[14] & g[22352];
assign g[55119] = b[14] & g[22352];
assign g[38737] = a[14] & g[22353];
assign g[55120] = b[14] & g[22353];
assign g[38738] = a[14] & g[22354];
assign g[55121] = b[14] & g[22354];
assign g[38739] = a[14] & g[22355];
assign g[55122] = b[14] & g[22355];
assign g[38740] = a[14] & g[22356];
assign g[55123] = b[14] & g[22356];
assign g[38741] = a[14] & g[22357];
assign g[55124] = b[14] & g[22357];
assign g[38742] = a[14] & g[22358];
assign g[55125] = b[14] & g[22358];
assign g[38743] = a[14] & g[22359];
assign g[55126] = b[14] & g[22359];
assign g[38744] = a[14] & g[22360];
assign g[55127] = b[14] & g[22360];
assign g[38745] = a[14] & g[22361];
assign g[55128] = b[14] & g[22361];
assign g[38746] = a[14] & g[22362];
assign g[55129] = b[14] & g[22362];
assign g[38747] = a[14] & g[22363];
assign g[55130] = b[14] & g[22363];
assign g[38748] = a[14] & g[22364];
assign g[55131] = b[14] & g[22364];
assign g[38749] = a[14] & g[22365];
assign g[55132] = b[14] & g[22365];
assign g[38750] = a[14] & g[22366];
assign g[55133] = b[14] & g[22366];
assign g[38751] = a[14] & g[22367];
assign g[55134] = b[14] & g[22367];
assign g[38752] = a[14] & g[22368];
assign g[55135] = b[14] & g[22368];
assign g[38753] = a[14] & g[22369];
assign g[55136] = b[14] & g[22369];
assign g[38754] = a[14] & g[22370];
assign g[55137] = b[14] & g[22370];
assign g[38755] = a[14] & g[22371];
assign g[55138] = b[14] & g[22371];
assign g[38756] = a[14] & g[22372];
assign g[55139] = b[14] & g[22372];
assign g[38757] = a[14] & g[22373];
assign g[55140] = b[14] & g[22373];
assign g[38758] = a[14] & g[22374];
assign g[55141] = b[14] & g[22374];
assign g[38759] = a[14] & g[22375];
assign g[55142] = b[14] & g[22375];
assign g[38760] = a[14] & g[22376];
assign g[55143] = b[14] & g[22376];
assign g[38761] = a[14] & g[22377];
assign g[55144] = b[14] & g[22377];
assign g[38762] = a[14] & g[22378];
assign g[55145] = b[14] & g[22378];
assign g[38763] = a[14] & g[22379];
assign g[55146] = b[14] & g[22379];
assign g[38764] = a[14] & g[22380];
assign g[55147] = b[14] & g[22380];
assign g[38765] = a[14] & g[22381];
assign g[55148] = b[14] & g[22381];
assign g[38766] = a[14] & g[22382];
assign g[55149] = b[14] & g[22382];
assign g[38767] = a[14] & g[22383];
assign g[55150] = b[14] & g[22383];
assign g[38768] = a[14] & g[22384];
assign g[55151] = b[14] & g[22384];
assign g[38769] = a[14] & g[22385];
assign g[55152] = b[14] & g[22385];
assign g[38770] = a[14] & g[22386];
assign g[55153] = b[14] & g[22386];
assign g[38771] = a[14] & g[22387];
assign g[55154] = b[14] & g[22387];
assign g[38772] = a[14] & g[22388];
assign g[55155] = b[14] & g[22388];
assign g[38773] = a[14] & g[22389];
assign g[55156] = b[14] & g[22389];
assign g[38774] = a[14] & g[22390];
assign g[55157] = b[14] & g[22390];
assign g[38775] = a[14] & g[22391];
assign g[55158] = b[14] & g[22391];
assign g[38776] = a[14] & g[22392];
assign g[55159] = b[14] & g[22392];
assign g[38777] = a[14] & g[22393];
assign g[55160] = b[14] & g[22393];
assign g[38778] = a[14] & g[22394];
assign g[55161] = b[14] & g[22394];
assign g[38779] = a[14] & g[22395];
assign g[55162] = b[14] & g[22395];
assign g[38780] = a[14] & g[22396];
assign g[55163] = b[14] & g[22396];
assign g[38781] = a[14] & g[22397];
assign g[55164] = b[14] & g[22397];
assign g[38782] = a[14] & g[22398];
assign g[55165] = b[14] & g[22398];
assign g[38783] = a[14] & g[22399];
assign g[55166] = b[14] & g[22399];
assign g[38784] = a[14] & g[22400];
assign g[55167] = b[14] & g[22400];
assign g[38785] = a[14] & g[22401];
assign g[55168] = b[14] & g[22401];
assign g[38786] = a[14] & g[22402];
assign g[55169] = b[14] & g[22402];
assign g[38787] = a[14] & g[22403];
assign g[55170] = b[14] & g[22403];
assign g[38788] = a[14] & g[22404];
assign g[55171] = b[14] & g[22404];
assign g[38789] = a[14] & g[22405];
assign g[55172] = b[14] & g[22405];
assign g[38790] = a[14] & g[22406];
assign g[55173] = b[14] & g[22406];
assign g[38791] = a[14] & g[22407];
assign g[55174] = b[14] & g[22407];
assign g[38792] = a[14] & g[22408];
assign g[55175] = b[14] & g[22408];
assign g[38793] = a[14] & g[22409];
assign g[55176] = b[14] & g[22409];
assign g[38794] = a[14] & g[22410];
assign g[55177] = b[14] & g[22410];
assign g[38795] = a[14] & g[22411];
assign g[55178] = b[14] & g[22411];
assign g[38796] = a[14] & g[22412];
assign g[55179] = b[14] & g[22412];
assign g[38797] = a[14] & g[22413];
assign g[55180] = b[14] & g[22413];
assign g[38798] = a[14] & g[22414];
assign g[55181] = b[14] & g[22414];
assign g[38799] = a[14] & g[22415];
assign g[55182] = b[14] & g[22415];
assign g[38800] = a[14] & g[22416];
assign g[55183] = b[14] & g[22416];
assign g[38801] = a[14] & g[22417];
assign g[55184] = b[14] & g[22417];
assign g[38802] = a[14] & g[22418];
assign g[55185] = b[14] & g[22418];
assign g[38803] = a[14] & g[22419];
assign g[55186] = b[14] & g[22419];
assign g[38804] = a[14] & g[22420];
assign g[55187] = b[14] & g[22420];
assign g[38805] = a[14] & g[22421];
assign g[55188] = b[14] & g[22421];
assign g[38806] = a[14] & g[22422];
assign g[55189] = b[14] & g[22422];
assign g[38807] = a[14] & g[22423];
assign g[55190] = b[14] & g[22423];
assign g[38808] = a[14] & g[22424];
assign g[55191] = b[14] & g[22424];
assign g[38809] = a[14] & g[22425];
assign g[55192] = b[14] & g[22425];
assign g[38810] = a[14] & g[22426];
assign g[55193] = b[14] & g[22426];
assign g[38811] = a[14] & g[22427];
assign g[55194] = b[14] & g[22427];
assign g[38812] = a[14] & g[22428];
assign g[55195] = b[14] & g[22428];
assign g[38813] = a[14] & g[22429];
assign g[55196] = b[14] & g[22429];
assign g[38814] = a[14] & g[22430];
assign g[55197] = b[14] & g[22430];
assign g[38815] = a[14] & g[22431];
assign g[55198] = b[14] & g[22431];
assign g[38816] = a[14] & g[22432];
assign g[55199] = b[14] & g[22432];
assign g[38817] = a[14] & g[22433];
assign g[55200] = b[14] & g[22433];
assign g[38818] = a[14] & g[22434];
assign g[55201] = b[14] & g[22434];
assign g[38819] = a[14] & g[22435];
assign g[55202] = b[14] & g[22435];
assign g[38820] = a[14] & g[22436];
assign g[55203] = b[14] & g[22436];
assign g[38821] = a[14] & g[22437];
assign g[55204] = b[14] & g[22437];
assign g[38822] = a[14] & g[22438];
assign g[55205] = b[14] & g[22438];
assign g[38823] = a[14] & g[22439];
assign g[55206] = b[14] & g[22439];
assign g[38824] = a[14] & g[22440];
assign g[55207] = b[14] & g[22440];
assign g[38825] = a[14] & g[22441];
assign g[55208] = b[14] & g[22441];
assign g[38826] = a[14] & g[22442];
assign g[55209] = b[14] & g[22442];
assign g[38827] = a[14] & g[22443];
assign g[55210] = b[14] & g[22443];
assign g[38828] = a[14] & g[22444];
assign g[55211] = b[14] & g[22444];
assign g[38829] = a[14] & g[22445];
assign g[55212] = b[14] & g[22445];
assign g[38830] = a[14] & g[22446];
assign g[55213] = b[14] & g[22446];
assign g[38831] = a[14] & g[22447];
assign g[55214] = b[14] & g[22447];
assign g[38832] = a[14] & g[22448];
assign g[55215] = b[14] & g[22448];
assign g[38833] = a[14] & g[22449];
assign g[55216] = b[14] & g[22449];
assign g[38834] = a[14] & g[22450];
assign g[55217] = b[14] & g[22450];
assign g[38835] = a[14] & g[22451];
assign g[55218] = b[14] & g[22451];
assign g[38836] = a[14] & g[22452];
assign g[55219] = b[14] & g[22452];
assign g[38837] = a[14] & g[22453];
assign g[55220] = b[14] & g[22453];
assign g[38838] = a[14] & g[22454];
assign g[55221] = b[14] & g[22454];
assign g[38839] = a[14] & g[22455];
assign g[55222] = b[14] & g[22455];
assign g[38840] = a[14] & g[22456];
assign g[55223] = b[14] & g[22456];
assign g[38841] = a[14] & g[22457];
assign g[55224] = b[14] & g[22457];
assign g[38842] = a[14] & g[22458];
assign g[55225] = b[14] & g[22458];
assign g[38843] = a[14] & g[22459];
assign g[55226] = b[14] & g[22459];
assign g[38844] = a[14] & g[22460];
assign g[55227] = b[14] & g[22460];
assign g[38845] = a[14] & g[22461];
assign g[55228] = b[14] & g[22461];
assign g[38846] = a[14] & g[22462];
assign g[55229] = b[14] & g[22462];
assign g[38847] = a[14] & g[22463];
assign g[55230] = b[14] & g[22463];
assign g[38848] = a[14] & g[22464];
assign g[55231] = b[14] & g[22464];
assign g[38849] = a[14] & g[22465];
assign g[55232] = b[14] & g[22465];
assign g[38850] = a[14] & g[22466];
assign g[55233] = b[14] & g[22466];
assign g[38851] = a[14] & g[22467];
assign g[55234] = b[14] & g[22467];
assign g[38852] = a[14] & g[22468];
assign g[55235] = b[14] & g[22468];
assign g[38853] = a[14] & g[22469];
assign g[55236] = b[14] & g[22469];
assign g[38854] = a[14] & g[22470];
assign g[55237] = b[14] & g[22470];
assign g[38855] = a[14] & g[22471];
assign g[55238] = b[14] & g[22471];
assign g[38856] = a[14] & g[22472];
assign g[55239] = b[14] & g[22472];
assign g[38857] = a[14] & g[22473];
assign g[55240] = b[14] & g[22473];
assign g[38858] = a[14] & g[22474];
assign g[55241] = b[14] & g[22474];
assign g[38859] = a[14] & g[22475];
assign g[55242] = b[14] & g[22475];
assign g[38860] = a[14] & g[22476];
assign g[55243] = b[14] & g[22476];
assign g[38861] = a[14] & g[22477];
assign g[55244] = b[14] & g[22477];
assign g[38862] = a[14] & g[22478];
assign g[55245] = b[14] & g[22478];
assign g[38863] = a[14] & g[22479];
assign g[55246] = b[14] & g[22479];
assign g[38864] = a[14] & g[22480];
assign g[55247] = b[14] & g[22480];
assign g[38865] = a[14] & g[22481];
assign g[55248] = b[14] & g[22481];
assign g[38866] = a[14] & g[22482];
assign g[55249] = b[14] & g[22482];
assign g[38867] = a[14] & g[22483];
assign g[55250] = b[14] & g[22483];
assign g[38868] = a[14] & g[22484];
assign g[55251] = b[14] & g[22484];
assign g[38869] = a[14] & g[22485];
assign g[55252] = b[14] & g[22485];
assign g[38870] = a[14] & g[22486];
assign g[55253] = b[14] & g[22486];
assign g[38871] = a[14] & g[22487];
assign g[55254] = b[14] & g[22487];
assign g[38872] = a[14] & g[22488];
assign g[55255] = b[14] & g[22488];
assign g[38873] = a[14] & g[22489];
assign g[55256] = b[14] & g[22489];
assign g[38874] = a[14] & g[22490];
assign g[55257] = b[14] & g[22490];
assign g[38875] = a[14] & g[22491];
assign g[55258] = b[14] & g[22491];
assign g[38876] = a[14] & g[22492];
assign g[55259] = b[14] & g[22492];
assign g[38877] = a[14] & g[22493];
assign g[55260] = b[14] & g[22493];
assign g[38878] = a[14] & g[22494];
assign g[55261] = b[14] & g[22494];
assign g[38879] = a[14] & g[22495];
assign g[55262] = b[14] & g[22495];
assign g[38880] = a[14] & g[22496];
assign g[55263] = b[14] & g[22496];
assign g[38881] = a[14] & g[22497];
assign g[55264] = b[14] & g[22497];
assign g[38882] = a[14] & g[22498];
assign g[55265] = b[14] & g[22498];
assign g[38883] = a[14] & g[22499];
assign g[55266] = b[14] & g[22499];
assign g[38884] = a[14] & g[22500];
assign g[55267] = b[14] & g[22500];
assign g[38885] = a[14] & g[22501];
assign g[55268] = b[14] & g[22501];
assign g[38886] = a[14] & g[22502];
assign g[55269] = b[14] & g[22502];
assign g[38887] = a[14] & g[22503];
assign g[55270] = b[14] & g[22503];
assign g[38888] = a[14] & g[22504];
assign g[55271] = b[14] & g[22504];
assign g[38889] = a[14] & g[22505];
assign g[55272] = b[14] & g[22505];
assign g[38890] = a[14] & g[22506];
assign g[55273] = b[14] & g[22506];
assign g[38891] = a[14] & g[22507];
assign g[55274] = b[14] & g[22507];
assign g[38892] = a[14] & g[22508];
assign g[55275] = b[14] & g[22508];
assign g[38893] = a[14] & g[22509];
assign g[55276] = b[14] & g[22509];
assign g[38894] = a[14] & g[22510];
assign g[55277] = b[14] & g[22510];
assign g[38895] = a[14] & g[22511];
assign g[55278] = b[14] & g[22511];
assign g[38896] = a[14] & g[22512];
assign g[55279] = b[14] & g[22512];
assign g[38897] = a[14] & g[22513];
assign g[55280] = b[14] & g[22513];
assign g[38898] = a[14] & g[22514];
assign g[55281] = b[14] & g[22514];
assign g[38899] = a[14] & g[22515];
assign g[55282] = b[14] & g[22515];
assign g[38900] = a[14] & g[22516];
assign g[55283] = b[14] & g[22516];
assign g[38901] = a[14] & g[22517];
assign g[55284] = b[14] & g[22517];
assign g[38902] = a[14] & g[22518];
assign g[55285] = b[14] & g[22518];
assign g[38903] = a[14] & g[22519];
assign g[55286] = b[14] & g[22519];
assign g[38904] = a[14] & g[22520];
assign g[55287] = b[14] & g[22520];
assign g[38905] = a[14] & g[22521];
assign g[55288] = b[14] & g[22521];
assign g[38906] = a[14] & g[22522];
assign g[55289] = b[14] & g[22522];
assign g[38907] = a[14] & g[22523];
assign g[55290] = b[14] & g[22523];
assign g[38908] = a[14] & g[22524];
assign g[55291] = b[14] & g[22524];
assign g[38909] = a[14] & g[22525];
assign g[55292] = b[14] & g[22525];
assign g[38910] = a[14] & g[22526];
assign g[55293] = b[14] & g[22526];
assign g[38911] = a[14] & g[22527];
assign g[55294] = b[14] & g[22527];
assign g[38912] = a[14] & g[22528];
assign g[55295] = b[14] & g[22528];
assign g[38913] = a[14] & g[22529];
assign g[55296] = b[14] & g[22529];
assign g[38914] = a[14] & g[22530];
assign g[55297] = b[14] & g[22530];
assign g[38915] = a[14] & g[22531];
assign g[55298] = b[14] & g[22531];
assign g[38916] = a[14] & g[22532];
assign g[55299] = b[14] & g[22532];
assign g[38917] = a[14] & g[22533];
assign g[55300] = b[14] & g[22533];
assign g[38918] = a[14] & g[22534];
assign g[55301] = b[14] & g[22534];
assign g[38919] = a[14] & g[22535];
assign g[55302] = b[14] & g[22535];
assign g[38920] = a[14] & g[22536];
assign g[55303] = b[14] & g[22536];
assign g[38921] = a[14] & g[22537];
assign g[55304] = b[14] & g[22537];
assign g[38922] = a[14] & g[22538];
assign g[55305] = b[14] & g[22538];
assign g[38923] = a[14] & g[22539];
assign g[55306] = b[14] & g[22539];
assign g[38924] = a[14] & g[22540];
assign g[55307] = b[14] & g[22540];
assign g[38925] = a[14] & g[22541];
assign g[55308] = b[14] & g[22541];
assign g[38926] = a[14] & g[22542];
assign g[55309] = b[14] & g[22542];
assign g[38927] = a[14] & g[22543];
assign g[55310] = b[14] & g[22543];
assign g[38928] = a[14] & g[22544];
assign g[55311] = b[14] & g[22544];
assign g[38929] = a[14] & g[22545];
assign g[55312] = b[14] & g[22545];
assign g[38930] = a[14] & g[22546];
assign g[55313] = b[14] & g[22546];
assign g[38931] = a[14] & g[22547];
assign g[55314] = b[14] & g[22547];
assign g[38932] = a[14] & g[22548];
assign g[55315] = b[14] & g[22548];
assign g[38933] = a[14] & g[22549];
assign g[55316] = b[14] & g[22549];
assign g[38934] = a[14] & g[22550];
assign g[55317] = b[14] & g[22550];
assign g[38935] = a[14] & g[22551];
assign g[55318] = b[14] & g[22551];
assign g[38936] = a[14] & g[22552];
assign g[55319] = b[14] & g[22552];
assign g[38937] = a[14] & g[22553];
assign g[55320] = b[14] & g[22553];
assign g[38938] = a[14] & g[22554];
assign g[55321] = b[14] & g[22554];
assign g[38939] = a[14] & g[22555];
assign g[55322] = b[14] & g[22555];
assign g[38940] = a[14] & g[22556];
assign g[55323] = b[14] & g[22556];
assign g[38941] = a[14] & g[22557];
assign g[55324] = b[14] & g[22557];
assign g[38942] = a[14] & g[22558];
assign g[55325] = b[14] & g[22558];
assign g[38943] = a[14] & g[22559];
assign g[55326] = b[14] & g[22559];
assign g[38944] = a[14] & g[22560];
assign g[55327] = b[14] & g[22560];
assign g[38945] = a[14] & g[22561];
assign g[55328] = b[14] & g[22561];
assign g[38946] = a[14] & g[22562];
assign g[55329] = b[14] & g[22562];
assign g[38947] = a[14] & g[22563];
assign g[55330] = b[14] & g[22563];
assign g[38948] = a[14] & g[22564];
assign g[55331] = b[14] & g[22564];
assign g[38949] = a[14] & g[22565];
assign g[55332] = b[14] & g[22565];
assign g[38950] = a[14] & g[22566];
assign g[55333] = b[14] & g[22566];
assign g[38951] = a[14] & g[22567];
assign g[55334] = b[14] & g[22567];
assign g[38952] = a[14] & g[22568];
assign g[55335] = b[14] & g[22568];
assign g[38953] = a[14] & g[22569];
assign g[55336] = b[14] & g[22569];
assign g[38954] = a[14] & g[22570];
assign g[55337] = b[14] & g[22570];
assign g[38955] = a[14] & g[22571];
assign g[55338] = b[14] & g[22571];
assign g[38956] = a[14] & g[22572];
assign g[55339] = b[14] & g[22572];
assign g[38957] = a[14] & g[22573];
assign g[55340] = b[14] & g[22573];
assign g[38958] = a[14] & g[22574];
assign g[55341] = b[14] & g[22574];
assign g[38959] = a[14] & g[22575];
assign g[55342] = b[14] & g[22575];
assign g[38960] = a[14] & g[22576];
assign g[55343] = b[14] & g[22576];
assign g[38961] = a[14] & g[22577];
assign g[55344] = b[14] & g[22577];
assign g[38962] = a[14] & g[22578];
assign g[55345] = b[14] & g[22578];
assign g[38963] = a[14] & g[22579];
assign g[55346] = b[14] & g[22579];
assign g[38964] = a[14] & g[22580];
assign g[55347] = b[14] & g[22580];
assign g[38965] = a[14] & g[22581];
assign g[55348] = b[14] & g[22581];
assign g[38966] = a[14] & g[22582];
assign g[55349] = b[14] & g[22582];
assign g[38967] = a[14] & g[22583];
assign g[55350] = b[14] & g[22583];
assign g[38968] = a[14] & g[22584];
assign g[55351] = b[14] & g[22584];
assign g[38969] = a[14] & g[22585];
assign g[55352] = b[14] & g[22585];
assign g[38970] = a[14] & g[22586];
assign g[55353] = b[14] & g[22586];
assign g[38971] = a[14] & g[22587];
assign g[55354] = b[14] & g[22587];
assign g[38972] = a[14] & g[22588];
assign g[55355] = b[14] & g[22588];
assign g[38973] = a[14] & g[22589];
assign g[55356] = b[14] & g[22589];
assign g[38974] = a[14] & g[22590];
assign g[55357] = b[14] & g[22590];
assign g[38975] = a[14] & g[22591];
assign g[55358] = b[14] & g[22591];
assign g[38976] = a[14] & g[22592];
assign g[55359] = b[14] & g[22592];
assign g[38977] = a[14] & g[22593];
assign g[55360] = b[14] & g[22593];
assign g[38978] = a[14] & g[22594];
assign g[55361] = b[14] & g[22594];
assign g[38979] = a[14] & g[22595];
assign g[55362] = b[14] & g[22595];
assign g[38980] = a[14] & g[22596];
assign g[55363] = b[14] & g[22596];
assign g[38981] = a[14] & g[22597];
assign g[55364] = b[14] & g[22597];
assign g[38982] = a[14] & g[22598];
assign g[55365] = b[14] & g[22598];
assign g[38983] = a[14] & g[22599];
assign g[55366] = b[14] & g[22599];
assign g[38984] = a[14] & g[22600];
assign g[55367] = b[14] & g[22600];
assign g[38985] = a[14] & g[22601];
assign g[55368] = b[14] & g[22601];
assign g[38986] = a[14] & g[22602];
assign g[55369] = b[14] & g[22602];
assign g[38987] = a[14] & g[22603];
assign g[55370] = b[14] & g[22603];
assign g[38988] = a[14] & g[22604];
assign g[55371] = b[14] & g[22604];
assign g[38989] = a[14] & g[22605];
assign g[55372] = b[14] & g[22605];
assign g[38990] = a[14] & g[22606];
assign g[55373] = b[14] & g[22606];
assign g[38991] = a[14] & g[22607];
assign g[55374] = b[14] & g[22607];
assign g[38992] = a[14] & g[22608];
assign g[55375] = b[14] & g[22608];
assign g[38993] = a[14] & g[22609];
assign g[55376] = b[14] & g[22609];
assign g[38994] = a[14] & g[22610];
assign g[55377] = b[14] & g[22610];
assign g[38995] = a[14] & g[22611];
assign g[55378] = b[14] & g[22611];
assign g[38996] = a[14] & g[22612];
assign g[55379] = b[14] & g[22612];
assign g[38997] = a[14] & g[22613];
assign g[55380] = b[14] & g[22613];
assign g[38998] = a[14] & g[22614];
assign g[55381] = b[14] & g[22614];
assign g[38999] = a[14] & g[22615];
assign g[55382] = b[14] & g[22615];
assign g[39000] = a[14] & g[22616];
assign g[55383] = b[14] & g[22616];
assign g[39001] = a[14] & g[22617];
assign g[55384] = b[14] & g[22617];
assign g[39002] = a[14] & g[22618];
assign g[55385] = b[14] & g[22618];
assign g[39003] = a[14] & g[22619];
assign g[55386] = b[14] & g[22619];
assign g[39004] = a[14] & g[22620];
assign g[55387] = b[14] & g[22620];
assign g[39005] = a[14] & g[22621];
assign g[55388] = b[14] & g[22621];
assign g[39006] = a[14] & g[22622];
assign g[55389] = b[14] & g[22622];
assign g[39007] = a[14] & g[22623];
assign g[55390] = b[14] & g[22623];
assign g[39008] = a[14] & g[22624];
assign g[55391] = b[14] & g[22624];
assign g[39009] = a[14] & g[22625];
assign g[55392] = b[14] & g[22625];
assign g[39010] = a[14] & g[22626];
assign g[55393] = b[14] & g[22626];
assign g[39011] = a[14] & g[22627];
assign g[55394] = b[14] & g[22627];
assign g[39012] = a[14] & g[22628];
assign g[55395] = b[14] & g[22628];
assign g[39013] = a[14] & g[22629];
assign g[55396] = b[14] & g[22629];
assign g[39014] = a[14] & g[22630];
assign g[55397] = b[14] & g[22630];
assign g[39015] = a[14] & g[22631];
assign g[55398] = b[14] & g[22631];
assign g[39016] = a[14] & g[22632];
assign g[55399] = b[14] & g[22632];
assign g[39017] = a[14] & g[22633];
assign g[55400] = b[14] & g[22633];
assign g[39018] = a[14] & g[22634];
assign g[55401] = b[14] & g[22634];
assign g[39019] = a[14] & g[22635];
assign g[55402] = b[14] & g[22635];
assign g[39020] = a[14] & g[22636];
assign g[55403] = b[14] & g[22636];
assign g[39021] = a[14] & g[22637];
assign g[55404] = b[14] & g[22637];
assign g[39022] = a[14] & g[22638];
assign g[55405] = b[14] & g[22638];
assign g[39023] = a[14] & g[22639];
assign g[55406] = b[14] & g[22639];
assign g[39024] = a[14] & g[22640];
assign g[55407] = b[14] & g[22640];
assign g[39025] = a[14] & g[22641];
assign g[55408] = b[14] & g[22641];
assign g[39026] = a[14] & g[22642];
assign g[55409] = b[14] & g[22642];
assign g[39027] = a[14] & g[22643];
assign g[55410] = b[14] & g[22643];
assign g[39028] = a[14] & g[22644];
assign g[55411] = b[14] & g[22644];
assign g[39029] = a[14] & g[22645];
assign g[55412] = b[14] & g[22645];
assign g[39030] = a[14] & g[22646];
assign g[55413] = b[14] & g[22646];
assign g[39031] = a[14] & g[22647];
assign g[55414] = b[14] & g[22647];
assign g[39032] = a[14] & g[22648];
assign g[55415] = b[14] & g[22648];
assign g[39033] = a[14] & g[22649];
assign g[55416] = b[14] & g[22649];
assign g[39034] = a[14] & g[22650];
assign g[55417] = b[14] & g[22650];
assign g[39035] = a[14] & g[22651];
assign g[55418] = b[14] & g[22651];
assign g[39036] = a[14] & g[22652];
assign g[55419] = b[14] & g[22652];
assign g[39037] = a[14] & g[22653];
assign g[55420] = b[14] & g[22653];
assign g[39038] = a[14] & g[22654];
assign g[55421] = b[14] & g[22654];
assign g[39039] = a[14] & g[22655];
assign g[55422] = b[14] & g[22655];
assign g[39040] = a[14] & g[22656];
assign g[55423] = b[14] & g[22656];
assign g[39041] = a[14] & g[22657];
assign g[55424] = b[14] & g[22657];
assign g[39042] = a[14] & g[22658];
assign g[55425] = b[14] & g[22658];
assign g[39043] = a[14] & g[22659];
assign g[55426] = b[14] & g[22659];
assign g[39044] = a[14] & g[22660];
assign g[55427] = b[14] & g[22660];
assign g[39045] = a[14] & g[22661];
assign g[55428] = b[14] & g[22661];
assign g[39046] = a[14] & g[22662];
assign g[55429] = b[14] & g[22662];
assign g[39047] = a[14] & g[22663];
assign g[55430] = b[14] & g[22663];
assign g[39048] = a[14] & g[22664];
assign g[55431] = b[14] & g[22664];
assign g[39049] = a[14] & g[22665];
assign g[55432] = b[14] & g[22665];
assign g[39050] = a[14] & g[22666];
assign g[55433] = b[14] & g[22666];
assign g[39051] = a[14] & g[22667];
assign g[55434] = b[14] & g[22667];
assign g[39052] = a[14] & g[22668];
assign g[55435] = b[14] & g[22668];
assign g[39053] = a[14] & g[22669];
assign g[55436] = b[14] & g[22669];
assign g[39054] = a[14] & g[22670];
assign g[55437] = b[14] & g[22670];
assign g[39055] = a[14] & g[22671];
assign g[55438] = b[14] & g[22671];
assign g[39056] = a[14] & g[22672];
assign g[55439] = b[14] & g[22672];
assign g[39057] = a[14] & g[22673];
assign g[55440] = b[14] & g[22673];
assign g[39058] = a[14] & g[22674];
assign g[55441] = b[14] & g[22674];
assign g[39059] = a[14] & g[22675];
assign g[55442] = b[14] & g[22675];
assign g[39060] = a[14] & g[22676];
assign g[55443] = b[14] & g[22676];
assign g[39061] = a[14] & g[22677];
assign g[55444] = b[14] & g[22677];
assign g[39062] = a[14] & g[22678];
assign g[55445] = b[14] & g[22678];
assign g[39063] = a[14] & g[22679];
assign g[55446] = b[14] & g[22679];
assign g[39064] = a[14] & g[22680];
assign g[55447] = b[14] & g[22680];
assign g[39065] = a[14] & g[22681];
assign g[55448] = b[14] & g[22681];
assign g[39066] = a[14] & g[22682];
assign g[55449] = b[14] & g[22682];
assign g[39067] = a[14] & g[22683];
assign g[55450] = b[14] & g[22683];
assign g[39068] = a[14] & g[22684];
assign g[55451] = b[14] & g[22684];
assign g[39069] = a[14] & g[22685];
assign g[55452] = b[14] & g[22685];
assign g[39070] = a[14] & g[22686];
assign g[55453] = b[14] & g[22686];
assign g[39071] = a[14] & g[22687];
assign g[55454] = b[14] & g[22687];
assign g[39072] = a[14] & g[22688];
assign g[55455] = b[14] & g[22688];
assign g[39073] = a[14] & g[22689];
assign g[55456] = b[14] & g[22689];
assign g[39074] = a[14] & g[22690];
assign g[55457] = b[14] & g[22690];
assign g[39075] = a[14] & g[22691];
assign g[55458] = b[14] & g[22691];
assign g[39076] = a[14] & g[22692];
assign g[55459] = b[14] & g[22692];
assign g[39077] = a[14] & g[22693];
assign g[55460] = b[14] & g[22693];
assign g[39078] = a[14] & g[22694];
assign g[55461] = b[14] & g[22694];
assign g[39079] = a[14] & g[22695];
assign g[55462] = b[14] & g[22695];
assign g[39080] = a[14] & g[22696];
assign g[55463] = b[14] & g[22696];
assign g[39081] = a[14] & g[22697];
assign g[55464] = b[14] & g[22697];
assign g[39082] = a[14] & g[22698];
assign g[55465] = b[14] & g[22698];
assign g[39083] = a[14] & g[22699];
assign g[55466] = b[14] & g[22699];
assign g[39084] = a[14] & g[22700];
assign g[55467] = b[14] & g[22700];
assign g[39085] = a[14] & g[22701];
assign g[55468] = b[14] & g[22701];
assign g[39086] = a[14] & g[22702];
assign g[55469] = b[14] & g[22702];
assign g[39087] = a[14] & g[22703];
assign g[55470] = b[14] & g[22703];
assign g[39088] = a[14] & g[22704];
assign g[55471] = b[14] & g[22704];
assign g[39089] = a[14] & g[22705];
assign g[55472] = b[14] & g[22705];
assign g[39090] = a[14] & g[22706];
assign g[55473] = b[14] & g[22706];
assign g[39091] = a[14] & g[22707];
assign g[55474] = b[14] & g[22707];
assign g[39092] = a[14] & g[22708];
assign g[55475] = b[14] & g[22708];
assign g[39093] = a[14] & g[22709];
assign g[55476] = b[14] & g[22709];
assign g[39094] = a[14] & g[22710];
assign g[55477] = b[14] & g[22710];
assign g[39095] = a[14] & g[22711];
assign g[55478] = b[14] & g[22711];
assign g[39096] = a[14] & g[22712];
assign g[55479] = b[14] & g[22712];
assign g[39097] = a[14] & g[22713];
assign g[55480] = b[14] & g[22713];
assign g[39098] = a[14] & g[22714];
assign g[55481] = b[14] & g[22714];
assign g[39099] = a[14] & g[22715];
assign g[55482] = b[14] & g[22715];
assign g[39100] = a[14] & g[22716];
assign g[55483] = b[14] & g[22716];
assign g[39101] = a[14] & g[22717];
assign g[55484] = b[14] & g[22717];
assign g[39102] = a[14] & g[22718];
assign g[55485] = b[14] & g[22718];
assign g[39103] = a[14] & g[22719];
assign g[55486] = b[14] & g[22719];
assign g[39104] = a[14] & g[22720];
assign g[55487] = b[14] & g[22720];
assign g[39105] = a[14] & g[22721];
assign g[55488] = b[14] & g[22721];
assign g[39106] = a[14] & g[22722];
assign g[55489] = b[14] & g[22722];
assign g[39107] = a[14] & g[22723];
assign g[55490] = b[14] & g[22723];
assign g[39108] = a[14] & g[22724];
assign g[55491] = b[14] & g[22724];
assign g[39109] = a[14] & g[22725];
assign g[55492] = b[14] & g[22725];
assign g[39110] = a[14] & g[22726];
assign g[55493] = b[14] & g[22726];
assign g[39111] = a[14] & g[22727];
assign g[55494] = b[14] & g[22727];
assign g[39112] = a[14] & g[22728];
assign g[55495] = b[14] & g[22728];
assign g[39113] = a[14] & g[22729];
assign g[55496] = b[14] & g[22729];
assign g[39114] = a[14] & g[22730];
assign g[55497] = b[14] & g[22730];
assign g[39115] = a[14] & g[22731];
assign g[55498] = b[14] & g[22731];
assign g[39116] = a[14] & g[22732];
assign g[55499] = b[14] & g[22732];
assign g[39117] = a[14] & g[22733];
assign g[55500] = b[14] & g[22733];
assign g[39118] = a[14] & g[22734];
assign g[55501] = b[14] & g[22734];
assign g[39119] = a[14] & g[22735];
assign g[55502] = b[14] & g[22735];
assign g[39120] = a[14] & g[22736];
assign g[55503] = b[14] & g[22736];
assign g[39121] = a[14] & g[22737];
assign g[55504] = b[14] & g[22737];
assign g[39122] = a[14] & g[22738];
assign g[55505] = b[14] & g[22738];
assign g[39123] = a[14] & g[22739];
assign g[55506] = b[14] & g[22739];
assign g[39124] = a[14] & g[22740];
assign g[55507] = b[14] & g[22740];
assign g[39125] = a[14] & g[22741];
assign g[55508] = b[14] & g[22741];
assign g[39126] = a[14] & g[22742];
assign g[55509] = b[14] & g[22742];
assign g[39127] = a[14] & g[22743];
assign g[55510] = b[14] & g[22743];
assign g[39128] = a[14] & g[22744];
assign g[55511] = b[14] & g[22744];
assign g[39129] = a[14] & g[22745];
assign g[55512] = b[14] & g[22745];
assign g[39130] = a[14] & g[22746];
assign g[55513] = b[14] & g[22746];
assign g[39131] = a[14] & g[22747];
assign g[55514] = b[14] & g[22747];
assign g[39132] = a[14] & g[22748];
assign g[55515] = b[14] & g[22748];
assign g[39133] = a[14] & g[22749];
assign g[55516] = b[14] & g[22749];
assign g[39134] = a[14] & g[22750];
assign g[55517] = b[14] & g[22750];
assign g[39135] = a[14] & g[22751];
assign g[55518] = b[14] & g[22751];
assign g[39136] = a[14] & g[22752];
assign g[55519] = b[14] & g[22752];
assign g[39137] = a[14] & g[22753];
assign g[55520] = b[14] & g[22753];
assign g[39138] = a[14] & g[22754];
assign g[55521] = b[14] & g[22754];
assign g[39139] = a[14] & g[22755];
assign g[55522] = b[14] & g[22755];
assign g[39140] = a[14] & g[22756];
assign g[55523] = b[14] & g[22756];
assign g[39141] = a[14] & g[22757];
assign g[55524] = b[14] & g[22757];
assign g[39142] = a[14] & g[22758];
assign g[55525] = b[14] & g[22758];
assign g[39143] = a[14] & g[22759];
assign g[55526] = b[14] & g[22759];
assign g[39144] = a[14] & g[22760];
assign g[55527] = b[14] & g[22760];
assign g[39145] = a[14] & g[22761];
assign g[55528] = b[14] & g[22761];
assign g[39146] = a[14] & g[22762];
assign g[55529] = b[14] & g[22762];
assign g[39147] = a[14] & g[22763];
assign g[55530] = b[14] & g[22763];
assign g[39148] = a[14] & g[22764];
assign g[55531] = b[14] & g[22764];
assign g[39149] = a[14] & g[22765];
assign g[55532] = b[14] & g[22765];
assign g[39150] = a[14] & g[22766];
assign g[55533] = b[14] & g[22766];
assign g[39151] = a[14] & g[22767];
assign g[55534] = b[14] & g[22767];
assign g[39152] = a[14] & g[22768];
assign g[55535] = b[14] & g[22768];
assign g[39153] = a[14] & g[22769];
assign g[55536] = b[14] & g[22769];
assign g[39154] = a[14] & g[22770];
assign g[55537] = b[14] & g[22770];
assign g[39155] = a[14] & g[22771];
assign g[55538] = b[14] & g[22771];
assign g[39156] = a[14] & g[22772];
assign g[55539] = b[14] & g[22772];
assign g[39157] = a[14] & g[22773];
assign g[55540] = b[14] & g[22773];
assign g[39158] = a[14] & g[22774];
assign g[55541] = b[14] & g[22774];
assign g[39159] = a[14] & g[22775];
assign g[55542] = b[14] & g[22775];
assign g[39160] = a[14] & g[22776];
assign g[55543] = b[14] & g[22776];
assign g[39161] = a[14] & g[22777];
assign g[55544] = b[14] & g[22777];
assign g[39162] = a[14] & g[22778];
assign g[55545] = b[14] & g[22778];
assign g[39163] = a[14] & g[22779];
assign g[55546] = b[14] & g[22779];
assign g[39164] = a[14] & g[22780];
assign g[55547] = b[14] & g[22780];
assign g[39165] = a[14] & g[22781];
assign g[55548] = b[14] & g[22781];
assign g[39166] = a[14] & g[22782];
assign g[55549] = b[14] & g[22782];
assign g[39167] = a[14] & g[22783];
assign g[55550] = b[14] & g[22783];
assign g[39168] = a[14] & g[22784];
assign g[55551] = b[14] & g[22784];
assign g[39169] = a[14] & g[22785];
assign g[55552] = b[14] & g[22785];
assign g[39170] = a[14] & g[22786];
assign g[55553] = b[14] & g[22786];
assign g[39171] = a[14] & g[22787];
assign g[55554] = b[14] & g[22787];
assign g[39172] = a[14] & g[22788];
assign g[55555] = b[14] & g[22788];
assign g[39173] = a[14] & g[22789];
assign g[55556] = b[14] & g[22789];
assign g[39174] = a[14] & g[22790];
assign g[55557] = b[14] & g[22790];
assign g[39175] = a[14] & g[22791];
assign g[55558] = b[14] & g[22791];
assign g[39176] = a[14] & g[22792];
assign g[55559] = b[14] & g[22792];
assign g[39177] = a[14] & g[22793];
assign g[55560] = b[14] & g[22793];
assign g[39178] = a[14] & g[22794];
assign g[55561] = b[14] & g[22794];
assign g[39179] = a[14] & g[22795];
assign g[55562] = b[14] & g[22795];
assign g[39180] = a[14] & g[22796];
assign g[55563] = b[14] & g[22796];
assign g[39181] = a[14] & g[22797];
assign g[55564] = b[14] & g[22797];
assign g[39182] = a[14] & g[22798];
assign g[55565] = b[14] & g[22798];
assign g[39183] = a[14] & g[22799];
assign g[55566] = b[14] & g[22799];
assign g[39184] = a[14] & g[22800];
assign g[55567] = b[14] & g[22800];
assign g[39185] = a[14] & g[22801];
assign g[55568] = b[14] & g[22801];
assign g[39186] = a[14] & g[22802];
assign g[55569] = b[14] & g[22802];
assign g[39187] = a[14] & g[22803];
assign g[55570] = b[14] & g[22803];
assign g[39188] = a[14] & g[22804];
assign g[55571] = b[14] & g[22804];
assign g[39189] = a[14] & g[22805];
assign g[55572] = b[14] & g[22805];
assign g[39190] = a[14] & g[22806];
assign g[55573] = b[14] & g[22806];
assign g[39191] = a[14] & g[22807];
assign g[55574] = b[14] & g[22807];
assign g[39192] = a[14] & g[22808];
assign g[55575] = b[14] & g[22808];
assign g[39193] = a[14] & g[22809];
assign g[55576] = b[14] & g[22809];
assign g[39194] = a[14] & g[22810];
assign g[55577] = b[14] & g[22810];
assign g[39195] = a[14] & g[22811];
assign g[55578] = b[14] & g[22811];
assign g[39196] = a[14] & g[22812];
assign g[55579] = b[14] & g[22812];
assign g[39197] = a[14] & g[22813];
assign g[55580] = b[14] & g[22813];
assign g[39198] = a[14] & g[22814];
assign g[55581] = b[14] & g[22814];
assign g[39199] = a[14] & g[22815];
assign g[55582] = b[14] & g[22815];
assign g[39200] = a[14] & g[22816];
assign g[55583] = b[14] & g[22816];
assign g[39201] = a[14] & g[22817];
assign g[55584] = b[14] & g[22817];
assign g[39202] = a[14] & g[22818];
assign g[55585] = b[14] & g[22818];
assign g[39203] = a[14] & g[22819];
assign g[55586] = b[14] & g[22819];
assign g[39204] = a[14] & g[22820];
assign g[55587] = b[14] & g[22820];
assign g[39205] = a[14] & g[22821];
assign g[55588] = b[14] & g[22821];
assign g[39206] = a[14] & g[22822];
assign g[55589] = b[14] & g[22822];
assign g[39207] = a[14] & g[22823];
assign g[55590] = b[14] & g[22823];
assign g[39208] = a[14] & g[22824];
assign g[55591] = b[14] & g[22824];
assign g[39209] = a[14] & g[22825];
assign g[55592] = b[14] & g[22825];
assign g[39210] = a[14] & g[22826];
assign g[55593] = b[14] & g[22826];
assign g[39211] = a[14] & g[22827];
assign g[55594] = b[14] & g[22827];
assign g[39212] = a[14] & g[22828];
assign g[55595] = b[14] & g[22828];
assign g[39213] = a[14] & g[22829];
assign g[55596] = b[14] & g[22829];
assign g[39214] = a[14] & g[22830];
assign g[55597] = b[14] & g[22830];
assign g[39215] = a[14] & g[22831];
assign g[55598] = b[14] & g[22831];
assign g[39216] = a[14] & g[22832];
assign g[55599] = b[14] & g[22832];
assign g[39217] = a[14] & g[22833];
assign g[55600] = b[14] & g[22833];
assign g[39218] = a[14] & g[22834];
assign g[55601] = b[14] & g[22834];
assign g[39219] = a[14] & g[22835];
assign g[55602] = b[14] & g[22835];
assign g[39220] = a[14] & g[22836];
assign g[55603] = b[14] & g[22836];
assign g[39221] = a[14] & g[22837];
assign g[55604] = b[14] & g[22837];
assign g[39222] = a[14] & g[22838];
assign g[55605] = b[14] & g[22838];
assign g[39223] = a[14] & g[22839];
assign g[55606] = b[14] & g[22839];
assign g[39224] = a[14] & g[22840];
assign g[55607] = b[14] & g[22840];
assign g[39225] = a[14] & g[22841];
assign g[55608] = b[14] & g[22841];
assign g[39226] = a[14] & g[22842];
assign g[55609] = b[14] & g[22842];
assign g[39227] = a[14] & g[22843];
assign g[55610] = b[14] & g[22843];
assign g[39228] = a[14] & g[22844];
assign g[55611] = b[14] & g[22844];
assign g[39229] = a[14] & g[22845];
assign g[55612] = b[14] & g[22845];
assign g[39230] = a[14] & g[22846];
assign g[55613] = b[14] & g[22846];
assign g[39231] = a[14] & g[22847];
assign g[55614] = b[14] & g[22847];
assign g[39232] = a[14] & g[22848];
assign g[55615] = b[14] & g[22848];
assign g[39233] = a[14] & g[22849];
assign g[55616] = b[14] & g[22849];
assign g[39234] = a[14] & g[22850];
assign g[55617] = b[14] & g[22850];
assign g[39235] = a[14] & g[22851];
assign g[55618] = b[14] & g[22851];
assign g[39236] = a[14] & g[22852];
assign g[55619] = b[14] & g[22852];
assign g[39237] = a[14] & g[22853];
assign g[55620] = b[14] & g[22853];
assign g[39238] = a[14] & g[22854];
assign g[55621] = b[14] & g[22854];
assign g[39239] = a[14] & g[22855];
assign g[55622] = b[14] & g[22855];
assign g[39240] = a[14] & g[22856];
assign g[55623] = b[14] & g[22856];
assign g[39241] = a[14] & g[22857];
assign g[55624] = b[14] & g[22857];
assign g[39242] = a[14] & g[22858];
assign g[55625] = b[14] & g[22858];
assign g[39243] = a[14] & g[22859];
assign g[55626] = b[14] & g[22859];
assign g[39244] = a[14] & g[22860];
assign g[55627] = b[14] & g[22860];
assign g[39245] = a[14] & g[22861];
assign g[55628] = b[14] & g[22861];
assign g[39246] = a[14] & g[22862];
assign g[55629] = b[14] & g[22862];
assign g[39247] = a[14] & g[22863];
assign g[55630] = b[14] & g[22863];
assign g[39248] = a[14] & g[22864];
assign g[55631] = b[14] & g[22864];
assign g[39249] = a[14] & g[22865];
assign g[55632] = b[14] & g[22865];
assign g[39250] = a[14] & g[22866];
assign g[55633] = b[14] & g[22866];
assign g[39251] = a[14] & g[22867];
assign g[55634] = b[14] & g[22867];
assign g[39252] = a[14] & g[22868];
assign g[55635] = b[14] & g[22868];
assign g[39253] = a[14] & g[22869];
assign g[55636] = b[14] & g[22869];
assign g[39254] = a[14] & g[22870];
assign g[55637] = b[14] & g[22870];
assign g[39255] = a[14] & g[22871];
assign g[55638] = b[14] & g[22871];
assign g[39256] = a[14] & g[22872];
assign g[55639] = b[14] & g[22872];
assign g[39257] = a[14] & g[22873];
assign g[55640] = b[14] & g[22873];
assign g[39258] = a[14] & g[22874];
assign g[55641] = b[14] & g[22874];
assign g[39259] = a[14] & g[22875];
assign g[55642] = b[14] & g[22875];
assign g[39260] = a[14] & g[22876];
assign g[55643] = b[14] & g[22876];
assign g[39261] = a[14] & g[22877];
assign g[55644] = b[14] & g[22877];
assign g[39262] = a[14] & g[22878];
assign g[55645] = b[14] & g[22878];
assign g[39263] = a[14] & g[22879];
assign g[55646] = b[14] & g[22879];
assign g[39264] = a[14] & g[22880];
assign g[55647] = b[14] & g[22880];
assign g[39265] = a[14] & g[22881];
assign g[55648] = b[14] & g[22881];
assign g[39266] = a[14] & g[22882];
assign g[55649] = b[14] & g[22882];
assign g[39267] = a[14] & g[22883];
assign g[55650] = b[14] & g[22883];
assign g[39268] = a[14] & g[22884];
assign g[55651] = b[14] & g[22884];
assign g[39269] = a[14] & g[22885];
assign g[55652] = b[14] & g[22885];
assign g[39270] = a[14] & g[22886];
assign g[55653] = b[14] & g[22886];
assign g[39271] = a[14] & g[22887];
assign g[55654] = b[14] & g[22887];
assign g[39272] = a[14] & g[22888];
assign g[55655] = b[14] & g[22888];
assign g[39273] = a[14] & g[22889];
assign g[55656] = b[14] & g[22889];
assign g[39274] = a[14] & g[22890];
assign g[55657] = b[14] & g[22890];
assign g[39275] = a[14] & g[22891];
assign g[55658] = b[14] & g[22891];
assign g[39276] = a[14] & g[22892];
assign g[55659] = b[14] & g[22892];
assign g[39277] = a[14] & g[22893];
assign g[55660] = b[14] & g[22893];
assign g[39278] = a[14] & g[22894];
assign g[55661] = b[14] & g[22894];
assign g[39279] = a[14] & g[22895];
assign g[55662] = b[14] & g[22895];
assign g[39280] = a[14] & g[22896];
assign g[55663] = b[14] & g[22896];
assign g[39281] = a[14] & g[22897];
assign g[55664] = b[14] & g[22897];
assign g[39282] = a[14] & g[22898];
assign g[55665] = b[14] & g[22898];
assign g[39283] = a[14] & g[22899];
assign g[55666] = b[14] & g[22899];
assign g[39284] = a[14] & g[22900];
assign g[55667] = b[14] & g[22900];
assign g[39285] = a[14] & g[22901];
assign g[55668] = b[14] & g[22901];
assign g[39286] = a[14] & g[22902];
assign g[55669] = b[14] & g[22902];
assign g[39287] = a[14] & g[22903];
assign g[55670] = b[14] & g[22903];
assign g[39288] = a[14] & g[22904];
assign g[55671] = b[14] & g[22904];
assign g[39289] = a[14] & g[22905];
assign g[55672] = b[14] & g[22905];
assign g[39290] = a[14] & g[22906];
assign g[55673] = b[14] & g[22906];
assign g[39291] = a[14] & g[22907];
assign g[55674] = b[14] & g[22907];
assign g[39292] = a[14] & g[22908];
assign g[55675] = b[14] & g[22908];
assign g[39293] = a[14] & g[22909];
assign g[55676] = b[14] & g[22909];
assign g[39294] = a[14] & g[22910];
assign g[55677] = b[14] & g[22910];
assign g[39295] = a[14] & g[22911];
assign g[55678] = b[14] & g[22911];
assign g[39296] = a[14] & g[22912];
assign g[55679] = b[14] & g[22912];
assign g[39297] = a[14] & g[22913];
assign g[55680] = b[14] & g[22913];
assign g[39298] = a[14] & g[22914];
assign g[55681] = b[14] & g[22914];
assign g[39299] = a[14] & g[22915];
assign g[55682] = b[14] & g[22915];
assign g[39300] = a[14] & g[22916];
assign g[55683] = b[14] & g[22916];
assign g[39301] = a[14] & g[22917];
assign g[55684] = b[14] & g[22917];
assign g[39302] = a[14] & g[22918];
assign g[55685] = b[14] & g[22918];
assign g[39303] = a[14] & g[22919];
assign g[55686] = b[14] & g[22919];
assign g[39304] = a[14] & g[22920];
assign g[55687] = b[14] & g[22920];
assign g[39305] = a[14] & g[22921];
assign g[55688] = b[14] & g[22921];
assign g[39306] = a[14] & g[22922];
assign g[55689] = b[14] & g[22922];
assign g[39307] = a[14] & g[22923];
assign g[55690] = b[14] & g[22923];
assign g[39308] = a[14] & g[22924];
assign g[55691] = b[14] & g[22924];
assign g[39309] = a[14] & g[22925];
assign g[55692] = b[14] & g[22925];
assign g[39310] = a[14] & g[22926];
assign g[55693] = b[14] & g[22926];
assign g[39311] = a[14] & g[22927];
assign g[55694] = b[14] & g[22927];
assign g[39312] = a[14] & g[22928];
assign g[55695] = b[14] & g[22928];
assign g[39313] = a[14] & g[22929];
assign g[55696] = b[14] & g[22929];
assign g[39314] = a[14] & g[22930];
assign g[55697] = b[14] & g[22930];
assign g[39315] = a[14] & g[22931];
assign g[55698] = b[14] & g[22931];
assign g[39316] = a[14] & g[22932];
assign g[55699] = b[14] & g[22932];
assign g[39317] = a[14] & g[22933];
assign g[55700] = b[14] & g[22933];
assign g[39318] = a[14] & g[22934];
assign g[55701] = b[14] & g[22934];
assign g[39319] = a[14] & g[22935];
assign g[55702] = b[14] & g[22935];
assign g[39320] = a[14] & g[22936];
assign g[55703] = b[14] & g[22936];
assign g[39321] = a[14] & g[22937];
assign g[55704] = b[14] & g[22937];
assign g[39322] = a[14] & g[22938];
assign g[55705] = b[14] & g[22938];
assign g[39323] = a[14] & g[22939];
assign g[55706] = b[14] & g[22939];
assign g[39324] = a[14] & g[22940];
assign g[55707] = b[14] & g[22940];
assign g[39325] = a[14] & g[22941];
assign g[55708] = b[14] & g[22941];
assign g[39326] = a[14] & g[22942];
assign g[55709] = b[14] & g[22942];
assign g[39327] = a[14] & g[22943];
assign g[55710] = b[14] & g[22943];
assign g[39328] = a[14] & g[22944];
assign g[55711] = b[14] & g[22944];
assign g[39329] = a[14] & g[22945];
assign g[55712] = b[14] & g[22945];
assign g[39330] = a[14] & g[22946];
assign g[55713] = b[14] & g[22946];
assign g[39331] = a[14] & g[22947];
assign g[55714] = b[14] & g[22947];
assign g[39332] = a[14] & g[22948];
assign g[55715] = b[14] & g[22948];
assign g[39333] = a[14] & g[22949];
assign g[55716] = b[14] & g[22949];
assign g[39334] = a[14] & g[22950];
assign g[55717] = b[14] & g[22950];
assign g[39335] = a[14] & g[22951];
assign g[55718] = b[14] & g[22951];
assign g[39336] = a[14] & g[22952];
assign g[55719] = b[14] & g[22952];
assign g[39337] = a[14] & g[22953];
assign g[55720] = b[14] & g[22953];
assign g[39338] = a[14] & g[22954];
assign g[55721] = b[14] & g[22954];
assign g[39339] = a[14] & g[22955];
assign g[55722] = b[14] & g[22955];
assign g[39340] = a[14] & g[22956];
assign g[55723] = b[14] & g[22956];
assign g[39341] = a[14] & g[22957];
assign g[55724] = b[14] & g[22957];
assign g[39342] = a[14] & g[22958];
assign g[55725] = b[14] & g[22958];
assign g[39343] = a[14] & g[22959];
assign g[55726] = b[14] & g[22959];
assign g[39344] = a[14] & g[22960];
assign g[55727] = b[14] & g[22960];
assign g[39345] = a[14] & g[22961];
assign g[55728] = b[14] & g[22961];
assign g[39346] = a[14] & g[22962];
assign g[55729] = b[14] & g[22962];
assign g[39347] = a[14] & g[22963];
assign g[55730] = b[14] & g[22963];
assign g[39348] = a[14] & g[22964];
assign g[55731] = b[14] & g[22964];
assign g[39349] = a[14] & g[22965];
assign g[55732] = b[14] & g[22965];
assign g[39350] = a[14] & g[22966];
assign g[55733] = b[14] & g[22966];
assign g[39351] = a[14] & g[22967];
assign g[55734] = b[14] & g[22967];
assign g[39352] = a[14] & g[22968];
assign g[55735] = b[14] & g[22968];
assign g[39353] = a[14] & g[22969];
assign g[55736] = b[14] & g[22969];
assign g[39354] = a[14] & g[22970];
assign g[55737] = b[14] & g[22970];
assign g[39355] = a[14] & g[22971];
assign g[55738] = b[14] & g[22971];
assign g[39356] = a[14] & g[22972];
assign g[55739] = b[14] & g[22972];
assign g[39357] = a[14] & g[22973];
assign g[55740] = b[14] & g[22973];
assign g[39358] = a[14] & g[22974];
assign g[55741] = b[14] & g[22974];
assign g[39359] = a[14] & g[22975];
assign g[55742] = b[14] & g[22975];
assign g[39360] = a[14] & g[22976];
assign g[55743] = b[14] & g[22976];
assign g[39361] = a[14] & g[22977];
assign g[55744] = b[14] & g[22977];
assign g[39362] = a[14] & g[22978];
assign g[55745] = b[14] & g[22978];
assign g[39363] = a[14] & g[22979];
assign g[55746] = b[14] & g[22979];
assign g[39364] = a[14] & g[22980];
assign g[55747] = b[14] & g[22980];
assign g[39365] = a[14] & g[22981];
assign g[55748] = b[14] & g[22981];
assign g[39366] = a[14] & g[22982];
assign g[55749] = b[14] & g[22982];
assign g[39367] = a[14] & g[22983];
assign g[55750] = b[14] & g[22983];
assign g[39368] = a[14] & g[22984];
assign g[55751] = b[14] & g[22984];
assign g[39369] = a[14] & g[22985];
assign g[55752] = b[14] & g[22985];
assign g[39370] = a[14] & g[22986];
assign g[55753] = b[14] & g[22986];
assign g[39371] = a[14] & g[22987];
assign g[55754] = b[14] & g[22987];
assign g[39372] = a[14] & g[22988];
assign g[55755] = b[14] & g[22988];
assign g[39373] = a[14] & g[22989];
assign g[55756] = b[14] & g[22989];
assign g[39374] = a[14] & g[22990];
assign g[55757] = b[14] & g[22990];
assign g[39375] = a[14] & g[22991];
assign g[55758] = b[14] & g[22991];
assign g[39376] = a[14] & g[22992];
assign g[55759] = b[14] & g[22992];
assign g[39377] = a[14] & g[22993];
assign g[55760] = b[14] & g[22993];
assign g[39378] = a[14] & g[22994];
assign g[55761] = b[14] & g[22994];
assign g[39379] = a[14] & g[22995];
assign g[55762] = b[14] & g[22995];
assign g[39380] = a[14] & g[22996];
assign g[55763] = b[14] & g[22996];
assign g[39381] = a[14] & g[22997];
assign g[55764] = b[14] & g[22997];
assign g[39382] = a[14] & g[22998];
assign g[55765] = b[14] & g[22998];
assign g[39383] = a[14] & g[22999];
assign g[55766] = b[14] & g[22999];
assign g[39384] = a[14] & g[23000];
assign g[55767] = b[14] & g[23000];
assign g[39385] = a[14] & g[23001];
assign g[55768] = b[14] & g[23001];
assign g[39386] = a[14] & g[23002];
assign g[55769] = b[14] & g[23002];
assign g[39387] = a[14] & g[23003];
assign g[55770] = b[14] & g[23003];
assign g[39388] = a[14] & g[23004];
assign g[55771] = b[14] & g[23004];
assign g[39389] = a[14] & g[23005];
assign g[55772] = b[14] & g[23005];
assign g[39390] = a[14] & g[23006];
assign g[55773] = b[14] & g[23006];
assign g[39391] = a[14] & g[23007];
assign g[55774] = b[14] & g[23007];
assign g[39392] = a[14] & g[23008];
assign g[55775] = b[14] & g[23008];
assign g[39393] = a[14] & g[23009];
assign g[55776] = b[14] & g[23009];
assign g[39394] = a[14] & g[23010];
assign g[55777] = b[14] & g[23010];
assign g[39395] = a[14] & g[23011];
assign g[55778] = b[14] & g[23011];
assign g[39396] = a[14] & g[23012];
assign g[55779] = b[14] & g[23012];
assign g[39397] = a[14] & g[23013];
assign g[55780] = b[14] & g[23013];
assign g[39398] = a[14] & g[23014];
assign g[55781] = b[14] & g[23014];
assign g[39399] = a[14] & g[23015];
assign g[55782] = b[14] & g[23015];
assign g[39400] = a[14] & g[23016];
assign g[55783] = b[14] & g[23016];
assign g[39401] = a[14] & g[23017];
assign g[55784] = b[14] & g[23017];
assign g[39402] = a[14] & g[23018];
assign g[55785] = b[14] & g[23018];
assign g[39403] = a[14] & g[23019];
assign g[55786] = b[14] & g[23019];
assign g[39404] = a[14] & g[23020];
assign g[55787] = b[14] & g[23020];
assign g[39405] = a[14] & g[23021];
assign g[55788] = b[14] & g[23021];
assign g[39406] = a[14] & g[23022];
assign g[55789] = b[14] & g[23022];
assign g[39407] = a[14] & g[23023];
assign g[55790] = b[14] & g[23023];
assign g[39408] = a[14] & g[23024];
assign g[55791] = b[14] & g[23024];
assign g[39409] = a[14] & g[23025];
assign g[55792] = b[14] & g[23025];
assign g[39410] = a[14] & g[23026];
assign g[55793] = b[14] & g[23026];
assign g[39411] = a[14] & g[23027];
assign g[55794] = b[14] & g[23027];
assign g[39412] = a[14] & g[23028];
assign g[55795] = b[14] & g[23028];
assign g[39413] = a[14] & g[23029];
assign g[55796] = b[14] & g[23029];
assign g[39414] = a[14] & g[23030];
assign g[55797] = b[14] & g[23030];
assign g[39415] = a[14] & g[23031];
assign g[55798] = b[14] & g[23031];
assign g[39416] = a[14] & g[23032];
assign g[55799] = b[14] & g[23032];
assign g[39417] = a[14] & g[23033];
assign g[55800] = b[14] & g[23033];
assign g[39418] = a[14] & g[23034];
assign g[55801] = b[14] & g[23034];
assign g[39419] = a[14] & g[23035];
assign g[55802] = b[14] & g[23035];
assign g[39420] = a[14] & g[23036];
assign g[55803] = b[14] & g[23036];
assign g[39421] = a[14] & g[23037];
assign g[55804] = b[14] & g[23037];
assign g[39422] = a[14] & g[23038];
assign g[55805] = b[14] & g[23038];
assign g[39423] = a[14] & g[23039];
assign g[55806] = b[14] & g[23039];
assign g[39424] = a[14] & g[23040];
assign g[55807] = b[14] & g[23040];
assign g[39425] = a[14] & g[23041];
assign g[55808] = b[14] & g[23041];
assign g[39426] = a[14] & g[23042];
assign g[55809] = b[14] & g[23042];
assign g[39427] = a[14] & g[23043];
assign g[55810] = b[14] & g[23043];
assign g[39428] = a[14] & g[23044];
assign g[55811] = b[14] & g[23044];
assign g[39429] = a[14] & g[23045];
assign g[55812] = b[14] & g[23045];
assign g[39430] = a[14] & g[23046];
assign g[55813] = b[14] & g[23046];
assign g[39431] = a[14] & g[23047];
assign g[55814] = b[14] & g[23047];
assign g[39432] = a[14] & g[23048];
assign g[55815] = b[14] & g[23048];
assign g[39433] = a[14] & g[23049];
assign g[55816] = b[14] & g[23049];
assign g[39434] = a[14] & g[23050];
assign g[55817] = b[14] & g[23050];
assign g[39435] = a[14] & g[23051];
assign g[55818] = b[14] & g[23051];
assign g[39436] = a[14] & g[23052];
assign g[55819] = b[14] & g[23052];
assign g[39437] = a[14] & g[23053];
assign g[55820] = b[14] & g[23053];
assign g[39438] = a[14] & g[23054];
assign g[55821] = b[14] & g[23054];
assign g[39439] = a[14] & g[23055];
assign g[55822] = b[14] & g[23055];
assign g[39440] = a[14] & g[23056];
assign g[55823] = b[14] & g[23056];
assign g[39441] = a[14] & g[23057];
assign g[55824] = b[14] & g[23057];
assign g[39442] = a[14] & g[23058];
assign g[55825] = b[14] & g[23058];
assign g[39443] = a[14] & g[23059];
assign g[55826] = b[14] & g[23059];
assign g[39444] = a[14] & g[23060];
assign g[55827] = b[14] & g[23060];
assign g[39445] = a[14] & g[23061];
assign g[55828] = b[14] & g[23061];
assign g[39446] = a[14] & g[23062];
assign g[55829] = b[14] & g[23062];
assign g[39447] = a[14] & g[23063];
assign g[55830] = b[14] & g[23063];
assign g[39448] = a[14] & g[23064];
assign g[55831] = b[14] & g[23064];
assign g[39449] = a[14] & g[23065];
assign g[55832] = b[14] & g[23065];
assign g[39450] = a[14] & g[23066];
assign g[55833] = b[14] & g[23066];
assign g[39451] = a[14] & g[23067];
assign g[55834] = b[14] & g[23067];
assign g[39452] = a[14] & g[23068];
assign g[55835] = b[14] & g[23068];
assign g[39453] = a[14] & g[23069];
assign g[55836] = b[14] & g[23069];
assign g[39454] = a[14] & g[23070];
assign g[55837] = b[14] & g[23070];
assign g[39455] = a[14] & g[23071];
assign g[55838] = b[14] & g[23071];
assign g[39456] = a[14] & g[23072];
assign g[55839] = b[14] & g[23072];
assign g[39457] = a[14] & g[23073];
assign g[55840] = b[14] & g[23073];
assign g[39458] = a[14] & g[23074];
assign g[55841] = b[14] & g[23074];
assign g[39459] = a[14] & g[23075];
assign g[55842] = b[14] & g[23075];
assign g[39460] = a[14] & g[23076];
assign g[55843] = b[14] & g[23076];
assign g[39461] = a[14] & g[23077];
assign g[55844] = b[14] & g[23077];
assign g[39462] = a[14] & g[23078];
assign g[55845] = b[14] & g[23078];
assign g[39463] = a[14] & g[23079];
assign g[55846] = b[14] & g[23079];
assign g[39464] = a[14] & g[23080];
assign g[55847] = b[14] & g[23080];
assign g[39465] = a[14] & g[23081];
assign g[55848] = b[14] & g[23081];
assign g[39466] = a[14] & g[23082];
assign g[55849] = b[14] & g[23082];
assign g[39467] = a[14] & g[23083];
assign g[55850] = b[14] & g[23083];
assign g[39468] = a[14] & g[23084];
assign g[55851] = b[14] & g[23084];
assign g[39469] = a[14] & g[23085];
assign g[55852] = b[14] & g[23085];
assign g[39470] = a[14] & g[23086];
assign g[55853] = b[14] & g[23086];
assign g[39471] = a[14] & g[23087];
assign g[55854] = b[14] & g[23087];
assign g[39472] = a[14] & g[23088];
assign g[55855] = b[14] & g[23088];
assign g[39473] = a[14] & g[23089];
assign g[55856] = b[14] & g[23089];
assign g[39474] = a[14] & g[23090];
assign g[55857] = b[14] & g[23090];
assign g[39475] = a[14] & g[23091];
assign g[55858] = b[14] & g[23091];
assign g[39476] = a[14] & g[23092];
assign g[55859] = b[14] & g[23092];
assign g[39477] = a[14] & g[23093];
assign g[55860] = b[14] & g[23093];
assign g[39478] = a[14] & g[23094];
assign g[55861] = b[14] & g[23094];
assign g[39479] = a[14] & g[23095];
assign g[55862] = b[14] & g[23095];
assign g[39480] = a[14] & g[23096];
assign g[55863] = b[14] & g[23096];
assign g[39481] = a[14] & g[23097];
assign g[55864] = b[14] & g[23097];
assign g[39482] = a[14] & g[23098];
assign g[55865] = b[14] & g[23098];
assign g[39483] = a[14] & g[23099];
assign g[55866] = b[14] & g[23099];
assign g[39484] = a[14] & g[23100];
assign g[55867] = b[14] & g[23100];
assign g[39485] = a[14] & g[23101];
assign g[55868] = b[14] & g[23101];
assign g[39486] = a[14] & g[23102];
assign g[55869] = b[14] & g[23102];
assign g[39487] = a[14] & g[23103];
assign g[55870] = b[14] & g[23103];
assign g[39488] = a[14] & g[23104];
assign g[55871] = b[14] & g[23104];
assign g[39489] = a[14] & g[23105];
assign g[55872] = b[14] & g[23105];
assign g[39490] = a[14] & g[23106];
assign g[55873] = b[14] & g[23106];
assign g[39491] = a[14] & g[23107];
assign g[55874] = b[14] & g[23107];
assign g[39492] = a[14] & g[23108];
assign g[55875] = b[14] & g[23108];
assign g[39493] = a[14] & g[23109];
assign g[55876] = b[14] & g[23109];
assign g[39494] = a[14] & g[23110];
assign g[55877] = b[14] & g[23110];
assign g[39495] = a[14] & g[23111];
assign g[55878] = b[14] & g[23111];
assign g[39496] = a[14] & g[23112];
assign g[55879] = b[14] & g[23112];
assign g[39497] = a[14] & g[23113];
assign g[55880] = b[14] & g[23113];
assign g[39498] = a[14] & g[23114];
assign g[55881] = b[14] & g[23114];
assign g[39499] = a[14] & g[23115];
assign g[55882] = b[14] & g[23115];
assign g[39500] = a[14] & g[23116];
assign g[55883] = b[14] & g[23116];
assign g[39501] = a[14] & g[23117];
assign g[55884] = b[14] & g[23117];
assign g[39502] = a[14] & g[23118];
assign g[55885] = b[14] & g[23118];
assign g[39503] = a[14] & g[23119];
assign g[55886] = b[14] & g[23119];
assign g[39504] = a[14] & g[23120];
assign g[55887] = b[14] & g[23120];
assign g[39505] = a[14] & g[23121];
assign g[55888] = b[14] & g[23121];
assign g[39506] = a[14] & g[23122];
assign g[55889] = b[14] & g[23122];
assign g[39507] = a[14] & g[23123];
assign g[55890] = b[14] & g[23123];
assign g[39508] = a[14] & g[23124];
assign g[55891] = b[14] & g[23124];
assign g[39509] = a[14] & g[23125];
assign g[55892] = b[14] & g[23125];
assign g[39510] = a[14] & g[23126];
assign g[55893] = b[14] & g[23126];
assign g[39511] = a[14] & g[23127];
assign g[55894] = b[14] & g[23127];
assign g[39512] = a[14] & g[23128];
assign g[55895] = b[14] & g[23128];
assign g[39513] = a[14] & g[23129];
assign g[55896] = b[14] & g[23129];
assign g[39514] = a[14] & g[23130];
assign g[55897] = b[14] & g[23130];
assign g[39515] = a[14] & g[23131];
assign g[55898] = b[14] & g[23131];
assign g[39516] = a[14] & g[23132];
assign g[55899] = b[14] & g[23132];
assign g[39517] = a[14] & g[23133];
assign g[55900] = b[14] & g[23133];
assign g[39518] = a[14] & g[23134];
assign g[55901] = b[14] & g[23134];
assign g[39519] = a[14] & g[23135];
assign g[55902] = b[14] & g[23135];
assign g[39520] = a[14] & g[23136];
assign g[55903] = b[14] & g[23136];
assign g[39521] = a[14] & g[23137];
assign g[55904] = b[14] & g[23137];
assign g[39522] = a[14] & g[23138];
assign g[55905] = b[14] & g[23138];
assign g[39523] = a[14] & g[23139];
assign g[55906] = b[14] & g[23139];
assign g[39524] = a[14] & g[23140];
assign g[55907] = b[14] & g[23140];
assign g[39525] = a[14] & g[23141];
assign g[55908] = b[14] & g[23141];
assign g[39526] = a[14] & g[23142];
assign g[55909] = b[14] & g[23142];
assign g[39527] = a[14] & g[23143];
assign g[55910] = b[14] & g[23143];
assign g[39528] = a[14] & g[23144];
assign g[55911] = b[14] & g[23144];
assign g[39529] = a[14] & g[23145];
assign g[55912] = b[14] & g[23145];
assign g[39530] = a[14] & g[23146];
assign g[55913] = b[14] & g[23146];
assign g[39531] = a[14] & g[23147];
assign g[55914] = b[14] & g[23147];
assign g[39532] = a[14] & g[23148];
assign g[55915] = b[14] & g[23148];
assign g[39533] = a[14] & g[23149];
assign g[55916] = b[14] & g[23149];
assign g[39534] = a[14] & g[23150];
assign g[55917] = b[14] & g[23150];
assign g[39535] = a[14] & g[23151];
assign g[55918] = b[14] & g[23151];
assign g[39536] = a[14] & g[23152];
assign g[55919] = b[14] & g[23152];
assign g[39537] = a[14] & g[23153];
assign g[55920] = b[14] & g[23153];
assign g[39538] = a[14] & g[23154];
assign g[55921] = b[14] & g[23154];
assign g[39539] = a[14] & g[23155];
assign g[55922] = b[14] & g[23155];
assign g[39540] = a[14] & g[23156];
assign g[55923] = b[14] & g[23156];
assign g[39541] = a[14] & g[23157];
assign g[55924] = b[14] & g[23157];
assign g[39542] = a[14] & g[23158];
assign g[55925] = b[14] & g[23158];
assign g[39543] = a[14] & g[23159];
assign g[55926] = b[14] & g[23159];
assign g[39544] = a[14] & g[23160];
assign g[55927] = b[14] & g[23160];
assign g[39545] = a[14] & g[23161];
assign g[55928] = b[14] & g[23161];
assign g[39546] = a[14] & g[23162];
assign g[55929] = b[14] & g[23162];
assign g[39547] = a[14] & g[23163];
assign g[55930] = b[14] & g[23163];
assign g[39548] = a[14] & g[23164];
assign g[55931] = b[14] & g[23164];
assign g[39549] = a[14] & g[23165];
assign g[55932] = b[14] & g[23165];
assign g[39550] = a[14] & g[23166];
assign g[55933] = b[14] & g[23166];
assign g[39551] = a[14] & g[23167];
assign g[55934] = b[14] & g[23167];
assign g[39552] = a[14] & g[23168];
assign g[55935] = b[14] & g[23168];
assign g[39553] = a[14] & g[23169];
assign g[55936] = b[14] & g[23169];
assign g[39554] = a[14] & g[23170];
assign g[55937] = b[14] & g[23170];
assign g[39555] = a[14] & g[23171];
assign g[55938] = b[14] & g[23171];
assign g[39556] = a[14] & g[23172];
assign g[55939] = b[14] & g[23172];
assign g[39557] = a[14] & g[23173];
assign g[55940] = b[14] & g[23173];
assign g[39558] = a[14] & g[23174];
assign g[55941] = b[14] & g[23174];
assign g[39559] = a[14] & g[23175];
assign g[55942] = b[14] & g[23175];
assign g[39560] = a[14] & g[23176];
assign g[55943] = b[14] & g[23176];
assign g[39561] = a[14] & g[23177];
assign g[55944] = b[14] & g[23177];
assign g[39562] = a[14] & g[23178];
assign g[55945] = b[14] & g[23178];
assign g[39563] = a[14] & g[23179];
assign g[55946] = b[14] & g[23179];
assign g[39564] = a[14] & g[23180];
assign g[55947] = b[14] & g[23180];
assign g[39565] = a[14] & g[23181];
assign g[55948] = b[14] & g[23181];
assign g[39566] = a[14] & g[23182];
assign g[55949] = b[14] & g[23182];
assign g[39567] = a[14] & g[23183];
assign g[55950] = b[14] & g[23183];
assign g[39568] = a[14] & g[23184];
assign g[55951] = b[14] & g[23184];
assign g[39569] = a[14] & g[23185];
assign g[55952] = b[14] & g[23185];
assign g[39570] = a[14] & g[23186];
assign g[55953] = b[14] & g[23186];
assign g[39571] = a[14] & g[23187];
assign g[55954] = b[14] & g[23187];
assign g[39572] = a[14] & g[23188];
assign g[55955] = b[14] & g[23188];
assign g[39573] = a[14] & g[23189];
assign g[55956] = b[14] & g[23189];
assign g[39574] = a[14] & g[23190];
assign g[55957] = b[14] & g[23190];
assign g[39575] = a[14] & g[23191];
assign g[55958] = b[14] & g[23191];
assign g[39576] = a[14] & g[23192];
assign g[55959] = b[14] & g[23192];
assign g[39577] = a[14] & g[23193];
assign g[55960] = b[14] & g[23193];
assign g[39578] = a[14] & g[23194];
assign g[55961] = b[14] & g[23194];
assign g[39579] = a[14] & g[23195];
assign g[55962] = b[14] & g[23195];
assign g[39580] = a[14] & g[23196];
assign g[55963] = b[14] & g[23196];
assign g[39581] = a[14] & g[23197];
assign g[55964] = b[14] & g[23197];
assign g[39582] = a[14] & g[23198];
assign g[55965] = b[14] & g[23198];
assign g[39583] = a[14] & g[23199];
assign g[55966] = b[14] & g[23199];
assign g[39584] = a[14] & g[23200];
assign g[55967] = b[14] & g[23200];
assign g[39585] = a[14] & g[23201];
assign g[55968] = b[14] & g[23201];
assign g[39586] = a[14] & g[23202];
assign g[55969] = b[14] & g[23202];
assign g[39587] = a[14] & g[23203];
assign g[55970] = b[14] & g[23203];
assign g[39588] = a[14] & g[23204];
assign g[55971] = b[14] & g[23204];
assign g[39589] = a[14] & g[23205];
assign g[55972] = b[14] & g[23205];
assign g[39590] = a[14] & g[23206];
assign g[55973] = b[14] & g[23206];
assign g[39591] = a[14] & g[23207];
assign g[55974] = b[14] & g[23207];
assign g[39592] = a[14] & g[23208];
assign g[55975] = b[14] & g[23208];
assign g[39593] = a[14] & g[23209];
assign g[55976] = b[14] & g[23209];
assign g[39594] = a[14] & g[23210];
assign g[55977] = b[14] & g[23210];
assign g[39595] = a[14] & g[23211];
assign g[55978] = b[14] & g[23211];
assign g[39596] = a[14] & g[23212];
assign g[55979] = b[14] & g[23212];
assign g[39597] = a[14] & g[23213];
assign g[55980] = b[14] & g[23213];
assign g[39598] = a[14] & g[23214];
assign g[55981] = b[14] & g[23214];
assign g[39599] = a[14] & g[23215];
assign g[55982] = b[14] & g[23215];
assign g[39600] = a[14] & g[23216];
assign g[55983] = b[14] & g[23216];
assign g[39601] = a[14] & g[23217];
assign g[55984] = b[14] & g[23217];
assign g[39602] = a[14] & g[23218];
assign g[55985] = b[14] & g[23218];
assign g[39603] = a[14] & g[23219];
assign g[55986] = b[14] & g[23219];
assign g[39604] = a[14] & g[23220];
assign g[55987] = b[14] & g[23220];
assign g[39605] = a[14] & g[23221];
assign g[55988] = b[14] & g[23221];
assign g[39606] = a[14] & g[23222];
assign g[55989] = b[14] & g[23222];
assign g[39607] = a[14] & g[23223];
assign g[55990] = b[14] & g[23223];
assign g[39608] = a[14] & g[23224];
assign g[55991] = b[14] & g[23224];
assign g[39609] = a[14] & g[23225];
assign g[55992] = b[14] & g[23225];
assign g[39610] = a[14] & g[23226];
assign g[55993] = b[14] & g[23226];
assign g[39611] = a[14] & g[23227];
assign g[55994] = b[14] & g[23227];
assign g[39612] = a[14] & g[23228];
assign g[55995] = b[14] & g[23228];
assign g[39613] = a[14] & g[23229];
assign g[55996] = b[14] & g[23229];
assign g[39614] = a[14] & g[23230];
assign g[55997] = b[14] & g[23230];
assign g[39615] = a[14] & g[23231];
assign g[55998] = b[14] & g[23231];
assign g[39616] = a[14] & g[23232];
assign g[55999] = b[14] & g[23232];
assign g[39617] = a[14] & g[23233];
assign g[56000] = b[14] & g[23233];
assign g[39618] = a[14] & g[23234];
assign g[56001] = b[14] & g[23234];
assign g[39619] = a[14] & g[23235];
assign g[56002] = b[14] & g[23235];
assign g[39620] = a[14] & g[23236];
assign g[56003] = b[14] & g[23236];
assign g[39621] = a[14] & g[23237];
assign g[56004] = b[14] & g[23237];
assign g[39622] = a[14] & g[23238];
assign g[56005] = b[14] & g[23238];
assign g[39623] = a[14] & g[23239];
assign g[56006] = b[14] & g[23239];
assign g[39624] = a[14] & g[23240];
assign g[56007] = b[14] & g[23240];
assign g[39625] = a[14] & g[23241];
assign g[56008] = b[14] & g[23241];
assign g[39626] = a[14] & g[23242];
assign g[56009] = b[14] & g[23242];
assign g[39627] = a[14] & g[23243];
assign g[56010] = b[14] & g[23243];
assign g[39628] = a[14] & g[23244];
assign g[56011] = b[14] & g[23244];
assign g[39629] = a[14] & g[23245];
assign g[56012] = b[14] & g[23245];
assign g[39630] = a[14] & g[23246];
assign g[56013] = b[14] & g[23246];
assign g[39631] = a[14] & g[23247];
assign g[56014] = b[14] & g[23247];
assign g[39632] = a[14] & g[23248];
assign g[56015] = b[14] & g[23248];
assign g[39633] = a[14] & g[23249];
assign g[56016] = b[14] & g[23249];
assign g[39634] = a[14] & g[23250];
assign g[56017] = b[14] & g[23250];
assign g[39635] = a[14] & g[23251];
assign g[56018] = b[14] & g[23251];
assign g[39636] = a[14] & g[23252];
assign g[56019] = b[14] & g[23252];
assign g[39637] = a[14] & g[23253];
assign g[56020] = b[14] & g[23253];
assign g[39638] = a[14] & g[23254];
assign g[56021] = b[14] & g[23254];
assign g[39639] = a[14] & g[23255];
assign g[56022] = b[14] & g[23255];
assign g[39640] = a[14] & g[23256];
assign g[56023] = b[14] & g[23256];
assign g[39641] = a[14] & g[23257];
assign g[56024] = b[14] & g[23257];
assign g[39642] = a[14] & g[23258];
assign g[56025] = b[14] & g[23258];
assign g[39643] = a[14] & g[23259];
assign g[56026] = b[14] & g[23259];
assign g[39644] = a[14] & g[23260];
assign g[56027] = b[14] & g[23260];
assign g[39645] = a[14] & g[23261];
assign g[56028] = b[14] & g[23261];
assign g[39646] = a[14] & g[23262];
assign g[56029] = b[14] & g[23262];
assign g[39647] = a[14] & g[23263];
assign g[56030] = b[14] & g[23263];
assign g[39648] = a[14] & g[23264];
assign g[56031] = b[14] & g[23264];
assign g[39649] = a[14] & g[23265];
assign g[56032] = b[14] & g[23265];
assign g[39650] = a[14] & g[23266];
assign g[56033] = b[14] & g[23266];
assign g[39651] = a[14] & g[23267];
assign g[56034] = b[14] & g[23267];
assign g[39652] = a[14] & g[23268];
assign g[56035] = b[14] & g[23268];
assign g[39653] = a[14] & g[23269];
assign g[56036] = b[14] & g[23269];
assign g[39654] = a[14] & g[23270];
assign g[56037] = b[14] & g[23270];
assign g[39655] = a[14] & g[23271];
assign g[56038] = b[14] & g[23271];
assign g[39656] = a[14] & g[23272];
assign g[56039] = b[14] & g[23272];
assign g[39657] = a[14] & g[23273];
assign g[56040] = b[14] & g[23273];
assign g[39658] = a[14] & g[23274];
assign g[56041] = b[14] & g[23274];
assign g[39659] = a[14] & g[23275];
assign g[56042] = b[14] & g[23275];
assign g[39660] = a[14] & g[23276];
assign g[56043] = b[14] & g[23276];
assign g[39661] = a[14] & g[23277];
assign g[56044] = b[14] & g[23277];
assign g[39662] = a[14] & g[23278];
assign g[56045] = b[14] & g[23278];
assign g[39663] = a[14] & g[23279];
assign g[56046] = b[14] & g[23279];
assign g[39664] = a[14] & g[23280];
assign g[56047] = b[14] & g[23280];
assign g[39665] = a[14] & g[23281];
assign g[56048] = b[14] & g[23281];
assign g[39666] = a[14] & g[23282];
assign g[56049] = b[14] & g[23282];
assign g[39667] = a[14] & g[23283];
assign g[56050] = b[14] & g[23283];
assign g[39668] = a[14] & g[23284];
assign g[56051] = b[14] & g[23284];
assign g[39669] = a[14] & g[23285];
assign g[56052] = b[14] & g[23285];
assign g[39670] = a[14] & g[23286];
assign g[56053] = b[14] & g[23286];
assign g[39671] = a[14] & g[23287];
assign g[56054] = b[14] & g[23287];
assign g[39672] = a[14] & g[23288];
assign g[56055] = b[14] & g[23288];
assign g[39673] = a[14] & g[23289];
assign g[56056] = b[14] & g[23289];
assign g[39674] = a[14] & g[23290];
assign g[56057] = b[14] & g[23290];
assign g[39675] = a[14] & g[23291];
assign g[56058] = b[14] & g[23291];
assign g[39676] = a[14] & g[23292];
assign g[56059] = b[14] & g[23292];
assign g[39677] = a[14] & g[23293];
assign g[56060] = b[14] & g[23293];
assign g[39678] = a[14] & g[23294];
assign g[56061] = b[14] & g[23294];
assign g[39679] = a[14] & g[23295];
assign g[56062] = b[14] & g[23295];
assign g[39680] = a[14] & g[23296];
assign g[56063] = b[14] & g[23296];
assign g[39681] = a[14] & g[23297];
assign g[56064] = b[14] & g[23297];
assign g[39682] = a[14] & g[23298];
assign g[56065] = b[14] & g[23298];
assign g[39683] = a[14] & g[23299];
assign g[56066] = b[14] & g[23299];
assign g[39684] = a[14] & g[23300];
assign g[56067] = b[14] & g[23300];
assign g[39685] = a[14] & g[23301];
assign g[56068] = b[14] & g[23301];
assign g[39686] = a[14] & g[23302];
assign g[56069] = b[14] & g[23302];
assign g[39687] = a[14] & g[23303];
assign g[56070] = b[14] & g[23303];
assign g[39688] = a[14] & g[23304];
assign g[56071] = b[14] & g[23304];
assign g[39689] = a[14] & g[23305];
assign g[56072] = b[14] & g[23305];
assign g[39690] = a[14] & g[23306];
assign g[56073] = b[14] & g[23306];
assign g[39691] = a[14] & g[23307];
assign g[56074] = b[14] & g[23307];
assign g[39692] = a[14] & g[23308];
assign g[56075] = b[14] & g[23308];
assign g[39693] = a[14] & g[23309];
assign g[56076] = b[14] & g[23309];
assign g[39694] = a[14] & g[23310];
assign g[56077] = b[14] & g[23310];
assign g[39695] = a[14] & g[23311];
assign g[56078] = b[14] & g[23311];
assign g[39696] = a[14] & g[23312];
assign g[56079] = b[14] & g[23312];
assign g[39697] = a[14] & g[23313];
assign g[56080] = b[14] & g[23313];
assign g[39698] = a[14] & g[23314];
assign g[56081] = b[14] & g[23314];
assign g[39699] = a[14] & g[23315];
assign g[56082] = b[14] & g[23315];
assign g[39700] = a[14] & g[23316];
assign g[56083] = b[14] & g[23316];
assign g[39701] = a[14] & g[23317];
assign g[56084] = b[14] & g[23317];
assign g[39702] = a[14] & g[23318];
assign g[56085] = b[14] & g[23318];
assign g[39703] = a[14] & g[23319];
assign g[56086] = b[14] & g[23319];
assign g[39704] = a[14] & g[23320];
assign g[56087] = b[14] & g[23320];
assign g[39705] = a[14] & g[23321];
assign g[56088] = b[14] & g[23321];
assign g[39706] = a[14] & g[23322];
assign g[56089] = b[14] & g[23322];
assign g[39707] = a[14] & g[23323];
assign g[56090] = b[14] & g[23323];
assign g[39708] = a[14] & g[23324];
assign g[56091] = b[14] & g[23324];
assign g[39709] = a[14] & g[23325];
assign g[56092] = b[14] & g[23325];
assign g[39710] = a[14] & g[23326];
assign g[56093] = b[14] & g[23326];
assign g[39711] = a[14] & g[23327];
assign g[56094] = b[14] & g[23327];
assign g[39712] = a[14] & g[23328];
assign g[56095] = b[14] & g[23328];
assign g[39713] = a[14] & g[23329];
assign g[56096] = b[14] & g[23329];
assign g[39714] = a[14] & g[23330];
assign g[56097] = b[14] & g[23330];
assign g[39715] = a[14] & g[23331];
assign g[56098] = b[14] & g[23331];
assign g[39716] = a[14] & g[23332];
assign g[56099] = b[14] & g[23332];
assign g[39717] = a[14] & g[23333];
assign g[56100] = b[14] & g[23333];
assign g[39718] = a[14] & g[23334];
assign g[56101] = b[14] & g[23334];
assign g[39719] = a[14] & g[23335];
assign g[56102] = b[14] & g[23335];
assign g[39720] = a[14] & g[23336];
assign g[56103] = b[14] & g[23336];
assign g[39721] = a[14] & g[23337];
assign g[56104] = b[14] & g[23337];
assign g[39722] = a[14] & g[23338];
assign g[56105] = b[14] & g[23338];
assign g[39723] = a[14] & g[23339];
assign g[56106] = b[14] & g[23339];
assign g[39724] = a[14] & g[23340];
assign g[56107] = b[14] & g[23340];
assign g[39725] = a[14] & g[23341];
assign g[56108] = b[14] & g[23341];
assign g[39726] = a[14] & g[23342];
assign g[56109] = b[14] & g[23342];
assign g[39727] = a[14] & g[23343];
assign g[56110] = b[14] & g[23343];
assign g[39728] = a[14] & g[23344];
assign g[56111] = b[14] & g[23344];
assign g[39729] = a[14] & g[23345];
assign g[56112] = b[14] & g[23345];
assign g[39730] = a[14] & g[23346];
assign g[56113] = b[14] & g[23346];
assign g[39731] = a[14] & g[23347];
assign g[56114] = b[14] & g[23347];
assign g[39732] = a[14] & g[23348];
assign g[56115] = b[14] & g[23348];
assign g[39733] = a[14] & g[23349];
assign g[56116] = b[14] & g[23349];
assign g[39734] = a[14] & g[23350];
assign g[56117] = b[14] & g[23350];
assign g[39735] = a[14] & g[23351];
assign g[56118] = b[14] & g[23351];
assign g[39736] = a[14] & g[23352];
assign g[56119] = b[14] & g[23352];
assign g[39737] = a[14] & g[23353];
assign g[56120] = b[14] & g[23353];
assign g[39738] = a[14] & g[23354];
assign g[56121] = b[14] & g[23354];
assign g[39739] = a[14] & g[23355];
assign g[56122] = b[14] & g[23355];
assign g[39740] = a[14] & g[23356];
assign g[56123] = b[14] & g[23356];
assign g[39741] = a[14] & g[23357];
assign g[56124] = b[14] & g[23357];
assign g[39742] = a[14] & g[23358];
assign g[56125] = b[14] & g[23358];
assign g[39743] = a[14] & g[23359];
assign g[56126] = b[14] & g[23359];
assign g[39744] = a[14] & g[23360];
assign g[56127] = b[14] & g[23360];
assign g[39745] = a[14] & g[23361];
assign g[56128] = b[14] & g[23361];
assign g[39746] = a[14] & g[23362];
assign g[56129] = b[14] & g[23362];
assign g[39747] = a[14] & g[23363];
assign g[56130] = b[14] & g[23363];
assign g[39748] = a[14] & g[23364];
assign g[56131] = b[14] & g[23364];
assign g[39749] = a[14] & g[23365];
assign g[56132] = b[14] & g[23365];
assign g[39750] = a[14] & g[23366];
assign g[56133] = b[14] & g[23366];
assign g[39751] = a[14] & g[23367];
assign g[56134] = b[14] & g[23367];
assign g[39752] = a[14] & g[23368];
assign g[56135] = b[14] & g[23368];
assign g[39753] = a[14] & g[23369];
assign g[56136] = b[14] & g[23369];
assign g[39754] = a[14] & g[23370];
assign g[56137] = b[14] & g[23370];
assign g[39755] = a[14] & g[23371];
assign g[56138] = b[14] & g[23371];
assign g[39756] = a[14] & g[23372];
assign g[56139] = b[14] & g[23372];
assign g[39757] = a[14] & g[23373];
assign g[56140] = b[14] & g[23373];
assign g[39758] = a[14] & g[23374];
assign g[56141] = b[14] & g[23374];
assign g[39759] = a[14] & g[23375];
assign g[56142] = b[14] & g[23375];
assign g[39760] = a[14] & g[23376];
assign g[56143] = b[14] & g[23376];
assign g[39761] = a[14] & g[23377];
assign g[56144] = b[14] & g[23377];
assign g[39762] = a[14] & g[23378];
assign g[56145] = b[14] & g[23378];
assign g[39763] = a[14] & g[23379];
assign g[56146] = b[14] & g[23379];
assign g[39764] = a[14] & g[23380];
assign g[56147] = b[14] & g[23380];
assign g[39765] = a[14] & g[23381];
assign g[56148] = b[14] & g[23381];
assign g[39766] = a[14] & g[23382];
assign g[56149] = b[14] & g[23382];
assign g[39767] = a[14] & g[23383];
assign g[56150] = b[14] & g[23383];
assign g[39768] = a[14] & g[23384];
assign g[56151] = b[14] & g[23384];
assign g[39769] = a[14] & g[23385];
assign g[56152] = b[14] & g[23385];
assign g[39770] = a[14] & g[23386];
assign g[56153] = b[14] & g[23386];
assign g[39771] = a[14] & g[23387];
assign g[56154] = b[14] & g[23387];
assign g[39772] = a[14] & g[23388];
assign g[56155] = b[14] & g[23388];
assign g[39773] = a[14] & g[23389];
assign g[56156] = b[14] & g[23389];
assign g[39774] = a[14] & g[23390];
assign g[56157] = b[14] & g[23390];
assign g[39775] = a[14] & g[23391];
assign g[56158] = b[14] & g[23391];
assign g[39776] = a[14] & g[23392];
assign g[56159] = b[14] & g[23392];
assign g[39777] = a[14] & g[23393];
assign g[56160] = b[14] & g[23393];
assign g[39778] = a[14] & g[23394];
assign g[56161] = b[14] & g[23394];
assign g[39779] = a[14] & g[23395];
assign g[56162] = b[14] & g[23395];
assign g[39780] = a[14] & g[23396];
assign g[56163] = b[14] & g[23396];
assign g[39781] = a[14] & g[23397];
assign g[56164] = b[14] & g[23397];
assign g[39782] = a[14] & g[23398];
assign g[56165] = b[14] & g[23398];
assign g[39783] = a[14] & g[23399];
assign g[56166] = b[14] & g[23399];
assign g[39784] = a[14] & g[23400];
assign g[56167] = b[14] & g[23400];
assign g[39785] = a[14] & g[23401];
assign g[56168] = b[14] & g[23401];
assign g[39786] = a[14] & g[23402];
assign g[56169] = b[14] & g[23402];
assign g[39787] = a[14] & g[23403];
assign g[56170] = b[14] & g[23403];
assign g[39788] = a[14] & g[23404];
assign g[56171] = b[14] & g[23404];
assign g[39789] = a[14] & g[23405];
assign g[56172] = b[14] & g[23405];
assign g[39790] = a[14] & g[23406];
assign g[56173] = b[14] & g[23406];
assign g[39791] = a[14] & g[23407];
assign g[56174] = b[14] & g[23407];
assign g[39792] = a[14] & g[23408];
assign g[56175] = b[14] & g[23408];
assign g[39793] = a[14] & g[23409];
assign g[56176] = b[14] & g[23409];
assign g[39794] = a[14] & g[23410];
assign g[56177] = b[14] & g[23410];
assign g[39795] = a[14] & g[23411];
assign g[56178] = b[14] & g[23411];
assign g[39796] = a[14] & g[23412];
assign g[56179] = b[14] & g[23412];
assign g[39797] = a[14] & g[23413];
assign g[56180] = b[14] & g[23413];
assign g[39798] = a[14] & g[23414];
assign g[56181] = b[14] & g[23414];
assign g[39799] = a[14] & g[23415];
assign g[56182] = b[14] & g[23415];
assign g[39800] = a[14] & g[23416];
assign g[56183] = b[14] & g[23416];
assign g[39801] = a[14] & g[23417];
assign g[56184] = b[14] & g[23417];
assign g[39802] = a[14] & g[23418];
assign g[56185] = b[14] & g[23418];
assign g[39803] = a[14] & g[23419];
assign g[56186] = b[14] & g[23419];
assign g[39804] = a[14] & g[23420];
assign g[56187] = b[14] & g[23420];
assign g[39805] = a[14] & g[23421];
assign g[56188] = b[14] & g[23421];
assign g[39806] = a[14] & g[23422];
assign g[56189] = b[14] & g[23422];
assign g[39807] = a[14] & g[23423];
assign g[56190] = b[14] & g[23423];
assign g[39808] = a[14] & g[23424];
assign g[56191] = b[14] & g[23424];
assign g[39809] = a[14] & g[23425];
assign g[56192] = b[14] & g[23425];
assign g[39810] = a[14] & g[23426];
assign g[56193] = b[14] & g[23426];
assign g[39811] = a[14] & g[23427];
assign g[56194] = b[14] & g[23427];
assign g[39812] = a[14] & g[23428];
assign g[56195] = b[14] & g[23428];
assign g[39813] = a[14] & g[23429];
assign g[56196] = b[14] & g[23429];
assign g[39814] = a[14] & g[23430];
assign g[56197] = b[14] & g[23430];
assign g[39815] = a[14] & g[23431];
assign g[56198] = b[14] & g[23431];
assign g[39816] = a[14] & g[23432];
assign g[56199] = b[14] & g[23432];
assign g[39817] = a[14] & g[23433];
assign g[56200] = b[14] & g[23433];
assign g[39818] = a[14] & g[23434];
assign g[56201] = b[14] & g[23434];
assign g[39819] = a[14] & g[23435];
assign g[56202] = b[14] & g[23435];
assign g[39820] = a[14] & g[23436];
assign g[56203] = b[14] & g[23436];
assign g[39821] = a[14] & g[23437];
assign g[56204] = b[14] & g[23437];
assign g[39822] = a[14] & g[23438];
assign g[56205] = b[14] & g[23438];
assign g[39823] = a[14] & g[23439];
assign g[56206] = b[14] & g[23439];
assign g[39824] = a[14] & g[23440];
assign g[56207] = b[14] & g[23440];
assign g[39825] = a[14] & g[23441];
assign g[56208] = b[14] & g[23441];
assign g[39826] = a[14] & g[23442];
assign g[56209] = b[14] & g[23442];
assign g[39827] = a[14] & g[23443];
assign g[56210] = b[14] & g[23443];
assign g[39828] = a[14] & g[23444];
assign g[56211] = b[14] & g[23444];
assign g[39829] = a[14] & g[23445];
assign g[56212] = b[14] & g[23445];
assign g[39830] = a[14] & g[23446];
assign g[56213] = b[14] & g[23446];
assign g[39831] = a[14] & g[23447];
assign g[56214] = b[14] & g[23447];
assign g[39832] = a[14] & g[23448];
assign g[56215] = b[14] & g[23448];
assign g[39833] = a[14] & g[23449];
assign g[56216] = b[14] & g[23449];
assign g[39834] = a[14] & g[23450];
assign g[56217] = b[14] & g[23450];
assign g[39835] = a[14] & g[23451];
assign g[56218] = b[14] & g[23451];
assign g[39836] = a[14] & g[23452];
assign g[56219] = b[14] & g[23452];
assign g[39837] = a[14] & g[23453];
assign g[56220] = b[14] & g[23453];
assign g[39838] = a[14] & g[23454];
assign g[56221] = b[14] & g[23454];
assign g[39839] = a[14] & g[23455];
assign g[56222] = b[14] & g[23455];
assign g[39840] = a[14] & g[23456];
assign g[56223] = b[14] & g[23456];
assign g[39841] = a[14] & g[23457];
assign g[56224] = b[14] & g[23457];
assign g[39842] = a[14] & g[23458];
assign g[56225] = b[14] & g[23458];
assign g[39843] = a[14] & g[23459];
assign g[56226] = b[14] & g[23459];
assign g[39844] = a[14] & g[23460];
assign g[56227] = b[14] & g[23460];
assign g[39845] = a[14] & g[23461];
assign g[56228] = b[14] & g[23461];
assign g[39846] = a[14] & g[23462];
assign g[56229] = b[14] & g[23462];
assign g[39847] = a[14] & g[23463];
assign g[56230] = b[14] & g[23463];
assign g[39848] = a[14] & g[23464];
assign g[56231] = b[14] & g[23464];
assign g[39849] = a[14] & g[23465];
assign g[56232] = b[14] & g[23465];
assign g[39850] = a[14] & g[23466];
assign g[56233] = b[14] & g[23466];
assign g[39851] = a[14] & g[23467];
assign g[56234] = b[14] & g[23467];
assign g[39852] = a[14] & g[23468];
assign g[56235] = b[14] & g[23468];
assign g[39853] = a[14] & g[23469];
assign g[56236] = b[14] & g[23469];
assign g[39854] = a[14] & g[23470];
assign g[56237] = b[14] & g[23470];
assign g[39855] = a[14] & g[23471];
assign g[56238] = b[14] & g[23471];
assign g[39856] = a[14] & g[23472];
assign g[56239] = b[14] & g[23472];
assign g[39857] = a[14] & g[23473];
assign g[56240] = b[14] & g[23473];
assign g[39858] = a[14] & g[23474];
assign g[56241] = b[14] & g[23474];
assign g[39859] = a[14] & g[23475];
assign g[56242] = b[14] & g[23475];
assign g[39860] = a[14] & g[23476];
assign g[56243] = b[14] & g[23476];
assign g[39861] = a[14] & g[23477];
assign g[56244] = b[14] & g[23477];
assign g[39862] = a[14] & g[23478];
assign g[56245] = b[14] & g[23478];
assign g[39863] = a[14] & g[23479];
assign g[56246] = b[14] & g[23479];
assign g[39864] = a[14] & g[23480];
assign g[56247] = b[14] & g[23480];
assign g[39865] = a[14] & g[23481];
assign g[56248] = b[14] & g[23481];
assign g[39866] = a[14] & g[23482];
assign g[56249] = b[14] & g[23482];
assign g[39867] = a[14] & g[23483];
assign g[56250] = b[14] & g[23483];
assign g[39868] = a[14] & g[23484];
assign g[56251] = b[14] & g[23484];
assign g[39869] = a[14] & g[23485];
assign g[56252] = b[14] & g[23485];
assign g[39870] = a[14] & g[23486];
assign g[56253] = b[14] & g[23486];
assign g[39871] = a[14] & g[23487];
assign g[56254] = b[14] & g[23487];
assign g[39872] = a[14] & g[23488];
assign g[56255] = b[14] & g[23488];
assign g[39873] = a[14] & g[23489];
assign g[56256] = b[14] & g[23489];
assign g[39874] = a[14] & g[23490];
assign g[56257] = b[14] & g[23490];
assign g[39875] = a[14] & g[23491];
assign g[56258] = b[14] & g[23491];
assign g[39876] = a[14] & g[23492];
assign g[56259] = b[14] & g[23492];
assign g[39877] = a[14] & g[23493];
assign g[56260] = b[14] & g[23493];
assign g[39878] = a[14] & g[23494];
assign g[56261] = b[14] & g[23494];
assign g[39879] = a[14] & g[23495];
assign g[56262] = b[14] & g[23495];
assign g[39880] = a[14] & g[23496];
assign g[56263] = b[14] & g[23496];
assign g[39881] = a[14] & g[23497];
assign g[56264] = b[14] & g[23497];
assign g[39882] = a[14] & g[23498];
assign g[56265] = b[14] & g[23498];
assign g[39883] = a[14] & g[23499];
assign g[56266] = b[14] & g[23499];
assign g[39884] = a[14] & g[23500];
assign g[56267] = b[14] & g[23500];
assign g[39885] = a[14] & g[23501];
assign g[56268] = b[14] & g[23501];
assign g[39886] = a[14] & g[23502];
assign g[56269] = b[14] & g[23502];
assign g[39887] = a[14] & g[23503];
assign g[56270] = b[14] & g[23503];
assign g[39888] = a[14] & g[23504];
assign g[56271] = b[14] & g[23504];
assign g[39889] = a[14] & g[23505];
assign g[56272] = b[14] & g[23505];
assign g[39890] = a[14] & g[23506];
assign g[56273] = b[14] & g[23506];
assign g[39891] = a[14] & g[23507];
assign g[56274] = b[14] & g[23507];
assign g[39892] = a[14] & g[23508];
assign g[56275] = b[14] & g[23508];
assign g[39893] = a[14] & g[23509];
assign g[56276] = b[14] & g[23509];
assign g[39894] = a[14] & g[23510];
assign g[56277] = b[14] & g[23510];
assign g[39895] = a[14] & g[23511];
assign g[56278] = b[14] & g[23511];
assign g[39896] = a[14] & g[23512];
assign g[56279] = b[14] & g[23512];
assign g[39897] = a[14] & g[23513];
assign g[56280] = b[14] & g[23513];
assign g[39898] = a[14] & g[23514];
assign g[56281] = b[14] & g[23514];
assign g[39899] = a[14] & g[23515];
assign g[56282] = b[14] & g[23515];
assign g[39900] = a[14] & g[23516];
assign g[56283] = b[14] & g[23516];
assign g[39901] = a[14] & g[23517];
assign g[56284] = b[14] & g[23517];
assign g[39902] = a[14] & g[23518];
assign g[56285] = b[14] & g[23518];
assign g[39903] = a[14] & g[23519];
assign g[56286] = b[14] & g[23519];
assign g[39904] = a[14] & g[23520];
assign g[56287] = b[14] & g[23520];
assign g[39905] = a[14] & g[23521];
assign g[56288] = b[14] & g[23521];
assign g[39906] = a[14] & g[23522];
assign g[56289] = b[14] & g[23522];
assign g[39907] = a[14] & g[23523];
assign g[56290] = b[14] & g[23523];
assign g[39908] = a[14] & g[23524];
assign g[56291] = b[14] & g[23524];
assign g[39909] = a[14] & g[23525];
assign g[56292] = b[14] & g[23525];
assign g[39910] = a[14] & g[23526];
assign g[56293] = b[14] & g[23526];
assign g[39911] = a[14] & g[23527];
assign g[56294] = b[14] & g[23527];
assign g[39912] = a[14] & g[23528];
assign g[56295] = b[14] & g[23528];
assign g[39913] = a[14] & g[23529];
assign g[56296] = b[14] & g[23529];
assign g[39914] = a[14] & g[23530];
assign g[56297] = b[14] & g[23530];
assign g[39915] = a[14] & g[23531];
assign g[56298] = b[14] & g[23531];
assign g[39916] = a[14] & g[23532];
assign g[56299] = b[14] & g[23532];
assign g[39917] = a[14] & g[23533];
assign g[56300] = b[14] & g[23533];
assign g[39918] = a[14] & g[23534];
assign g[56301] = b[14] & g[23534];
assign g[39919] = a[14] & g[23535];
assign g[56302] = b[14] & g[23535];
assign g[39920] = a[14] & g[23536];
assign g[56303] = b[14] & g[23536];
assign g[39921] = a[14] & g[23537];
assign g[56304] = b[14] & g[23537];
assign g[39922] = a[14] & g[23538];
assign g[56305] = b[14] & g[23538];
assign g[39923] = a[14] & g[23539];
assign g[56306] = b[14] & g[23539];
assign g[39924] = a[14] & g[23540];
assign g[56307] = b[14] & g[23540];
assign g[39925] = a[14] & g[23541];
assign g[56308] = b[14] & g[23541];
assign g[39926] = a[14] & g[23542];
assign g[56309] = b[14] & g[23542];
assign g[39927] = a[14] & g[23543];
assign g[56310] = b[14] & g[23543];
assign g[39928] = a[14] & g[23544];
assign g[56311] = b[14] & g[23544];
assign g[39929] = a[14] & g[23545];
assign g[56312] = b[14] & g[23545];
assign g[39930] = a[14] & g[23546];
assign g[56313] = b[14] & g[23546];
assign g[39931] = a[14] & g[23547];
assign g[56314] = b[14] & g[23547];
assign g[39932] = a[14] & g[23548];
assign g[56315] = b[14] & g[23548];
assign g[39933] = a[14] & g[23549];
assign g[56316] = b[14] & g[23549];
assign g[39934] = a[14] & g[23550];
assign g[56317] = b[14] & g[23550];
assign g[39935] = a[14] & g[23551];
assign g[56318] = b[14] & g[23551];
assign g[39936] = a[14] & g[23552];
assign g[56319] = b[14] & g[23552];
assign g[39937] = a[14] & g[23553];
assign g[56320] = b[14] & g[23553];
assign g[39938] = a[14] & g[23554];
assign g[56321] = b[14] & g[23554];
assign g[39939] = a[14] & g[23555];
assign g[56322] = b[14] & g[23555];
assign g[39940] = a[14] & g[23556];
assign g[56323] = b[14] & g[23556];
assign g[39941] = a[14] & g[23557];
assign g[56324] = b[14] & g[23557];
assign g[39942] = a[14] & g[23558];
assign g[56325] = b[14] & g[23558];
assign g[39943] = a[14] & g[23559];
assign g[56326] = b[14] & g[23559];
assign g[39944] = a[14] & g[23560];
assign g[56327] = b[14] & g[23560];
assign g[39945] = a[14] & g[23561];
assign g[56328] = b[14] & g[23561];
assign g[39946] = a[14] & g[23562];
assign g[56329] = b[14] & g[23562];
assign g[39947] = a[14] & g[23563];
assign g[56330] = b[14] & g[23563];
assign g[39948] = a[14] & g[23564];
assign g[56331] = b[14] & g[23564];
assign g[39949] = a[14] & g[23565];
assign g[56332] = b[14] & g[23565];
assign g[39950] = a[14] & g[23566];
assign g[56333] = b[14] & g[23566];
assign g[39951] = a[14] & g[23567];
assign g[56334] = b[14] & g[23567];
assign g[39952] = a[14] & g[23568];
assign g[56335] = b[14] & g[23568];
assign g[39953] = a[14] & g[23569];
assign g[56336] = b[14] & g[23569];
assign g[39954] = a[14] & g[23570];
assign g[56337] = b[14] & g[23570];
assign g[39955] = a[14] & g[23571];
assign g[56338] = b[14] & g[23571];
assign g[39956] = a[14] & g[23572];
assign g[56339] = b[14] & g[23572];
assign g[39957] = a[14] & g[23573];
assign g[56340] = b[14] & g[23573];
assign g[39958] = a[14] & g[23574];
assign g[56341] = b[14] & g[23574];
assign g[39959] = a[14] & g[23575];
assign g[56342] = b[14] & g[23575];
assign g[39960] = a[14] & g[23576];
assign g[56343] = b[14] & g[23576];
assign g[39961] = a[14] & g[23577];
assign g[56344] = b[14] & g[23577];
assign g[39962] = a[14] & g[23578];
assign g[56345] = b[14] & g[23578];
assign g[39963] = a[14] & g[23579];
assign g[56346] = b[14] & g[23579];
assign g[39964] = a[14] & g[23580];
assign g[56347] = b[14] & g[23580];
assign g[39965] = a[14] & g[23581];
assign g[56348] = b[14] & g[23581];
assign g[39966] = a[14] & g[23582];
assign g[56349] = b[14] & g[23582];
assign g[39967] = a[14] & g[23583];
assign g[56350] = b[14] & g[23583];
assign g[39968] = a[14] & g[23584];
assign g[56351] = b[14] & g[23584];
assign g[39969] = a[14] & g[23585];
assign g[56352] = b[14] & g[23585];
assign g[39970] = a[14] & g[23586];
assign g[56353] = b[14] & g[23586];
assign g[39971] = a[14] & g[23587];
assign g[56354] = b[14] & g[23587];
assign g[39972] = a[14] & g[23588];
assign g[56355] = b[14] & g[23588];
assign g[39973] = a[14] & g[23589];
assign g[56356] = b[14] & g[23589];
assign g[39974] = a[14] & g[23590];
assign g[56357] = b[14] & g[23590];
assign g[39975] = a[14] & g[23591];
assign g[56358] = b[14] & g[23591];
assign g[39976] = a[14] & g[23592];
assign g[56359] = b[14] & g[23592];
assign g[39977] = a[14] & g[23593];
assign g[56360] = b[14] & g[23593];
assign g[39978] = a[14] & g[23594];
assign g[56361] = b[14] & g[23594];
assign g[39979] = a[14] & g[23595];
assign g[56362] = b[14] & g[23595];
assign g[39980] = a[14] & g[23596];
assign g[56363] = b[14] & g[23596];
assign g[39981] = a[14] & g[23597];
assign g[56364] = b[14] & g[23597];
assign g[39982] = a[14] & g[23598];
assign g[56365] = b[14] & g[23598];
assign g[39983] = a[14] & g[23599];
assign g[56366] = b[14] & g[23599];
assign g[39984] = a[14] & g[23600];
assign g[56367] = b[14] & g[23600];
assign g[39985] = a[14] & g[23601];
assign g[56368] = b[14] & g[23601];
assign g[39986] = a[14] & g[23602];
assign g[56369] = b[14] & g[23602];
assign g[39987] = a[14] & g[23603];
assign g[56370] = b[14] & g[23603];
assign g[39988] = a[14] & g[23604];
assign g[56371] = b[14] & g[23604];
assign g[39989] = a[14] & g[23605];
assign g[56372] = b[14] & g[23605];
assign g[39990] = a[14] & g[23606];
assign g[56373] = b[14] & g[23606];
assign g[39991] = a[14] & g[23607];
assign g[56374] = b[14] & g[23607];
assign g[39992] = a[14] & g[23608];
assign g[56375] = b[14] & g[23608];
assign g[39993] = a[14] & g[23609];
assign g[56376] = b[14] & g[23609];
assign g[39994] = a[14] & g[23610];
assign g[56377] = b[14] & g[23610];
assign g[39995] = a[14] & g[23611];
assign g[56378] = b[14] & g[23611];
assign g[39996] = a[14] & g[23612];
assign g[56379] = b[14] & g[23612];
assign g[39997] = a[14] & g[23613];
assign g[56380] = b[14] & g[23613];
assign g[39998] = a[14] & g[23614];
assign g[56381] = b[14] & g[23614];
assign g[39999] = a[14] & g[23615];
assign g[56382] = b[14] & g[23615];
assign g[40000] = a[14] & g[23616];
assign g[56383] = b[14] & g[23616];
assign g[40001] = a[14] & g[23617];
assign g[56384] = b[14] & g[23617];
assign g[40002] = a[14] & g[23618];
assign g[56385] = b[14] & g[23618];
assign g[40003] = a[14] & g[23619];
assign g[56386] = b[14] & g[23619];
assign g[40004] = a[14] & g[23620];
assign g[56387] = b[14] & g[23620];
assign g[40005] = a[14] & g[23621];
assign g[56388] = b[14] & g[23621];
assign g[40006] = a[14] & g[23622];
assign g[56389] = b[14] & g[23622];
assign g[40007] = a[14] & g[23623];
assign g[56390] = b[14] & g[23623];
assign g[40008] = a[14] & g[23624];
assign g[56391] = b[14] & g[23624];
assign g[40009] = a[14] & g[23625];
assign g[56392] = b[14] & g[23625];
assign g[40010] = a[14] & g[23626];
assign g[56393] = b[14] & g[23626];
assign g[40011] = a[14] & g[23627];
assign g[56394] = b[14] & g[23627];
assign g[40012] = a[14] & g[23628];
assign g[56395] = b[14] & g[23628];
assign g[40013] = a[14] & g[23629];
assign g[56396] = b[14] & g[23629];
assign g[40014] = a[14] & g[23630];
assign g[56397] = b[14] & g[23630];
assign g[40015] = a[14] & g[23631];
assign g[56398] = b[14] & g[23631];
assign g[40016] = a[14] & g[23632];
assign g[56399] = b[14] & g[23632];
assign g[40017] = a[14] & g[23633];
assign g[56400] = b[14] & g[23633];
assign g[40018] = a[14] & g[23634];
assign g[56401] = b[14] & g[23634];
assign g[40019] = a[14] & g[23635];
assign g[56402] = b[14] & g[23635];
assign g[40020] = a[14] & g[23636];
assign g[56403] = b[14] & g[23636];
assign g[40021] = a[14] & g[23637];
assign g[56404] = b[14] & g[23637];
assign g[40022] = a[14] & g[23638];
assign g[56405] = b[14] & g[23638];
assign g[40023] = a[14] & g[23639];
assign g[56406] = b[14] & g[23639];
assign g[40024] = a[14] & g[23640];
assign g[56407] = b[14] & g[23640];
assign g[40025] = a[14] & g[23641];
assign g[56408] = b[14] & g[23641];
assign g[40026] = a[14] & g[23642];
assign g[56409] = b[14] & g[23642];
assign g[40027] = a[14] & g[23643];
assign g[56410] = b[14] & g[23643];
assign g[40028] = a[14] & g[23644];
assign g[56411] = b[14] & g[23644];
assign g[40029] = a[14] & g[23645];
assign g[56412] = b[14] & g[23645];
assign g[40030] = a[14] & g[23646];
assign g[56413] = b[14] & g[23646];
assign g[40031] = a[14] & g[23647];
assign g[56414] = b[14] & g[23647];
assign g[40032] = a[14] & g[23648];
assign g[56415] = b[14] & g[23648];
assign g[40033] = a[14] & g[23649];
assign g[56416] = b[14] & g[23649];
assign g[40034] = a[14] & g[23650];
assign g[56417] = b[14] & g[23650];
assign g[40035] = a[14] & g[23651];
assign g[56418] = b[14] & g[23651];
assign g[40036] = a[14] & g[23652];
assign g[56419] = b[14] & g[23652];
assign g[40037] = a[14] & g[23653];
assign g[56420] = b[14] & g[23653];
assign g[40038] = a[14] & g[23654];
assign g[56421] = b[14] & g[23654];
assign g[40039] = a[14] & g[23655];
assign g[56422] = b[14] & g[23655];
assign g[40040] = a[14] & g[23656];
assign g[56423] = b[14] & g[23656];
assign g[40041] = a[14] & g[23657];
assign g[56424] = b[14] & g[23657];
assign g[40042] = a[14] & g[23658];
assign g[56425] = b[14] & g[23658];
assign g[40043] = a[14] & g[23659];
assign g[56426] = b[14] & g[23659];
assign g[40044] = a[14] & g[23660];
assign g[56427] = b[14] & g[23660];
assign g[40045] = a[14] & g[23661];
assign g[56428] = b[14] & g[23661];
assign g[40046] = a[14] & g[23662];
assign g[56429] = b[14] & g[23662];
assign g[40047] = a[14] & g[23663];
assign g[56430] = b[14] & g[23663];
assign g[40048] = a[14] & g[23664];
assign g[56431] = b[14] & g[23664];
assign g[40049] = a[14] & g[23665];
assign g[56432] = b[14] & g[23665];
assign g[40050] = a[14] & g[23666];
assign g[56433] = b[14] & g[23666];
assign g[40051] = a[14] & g[23667];
assign g[56434] = b[14] & g[23667];
assign g[40052] = a[14] & g[23668];
assign g[56435] = b[14] & g[23668];
assign g[40053] = a[14] & g[23669];
assign g[56436] = b[14] & g[23669];
assign g[40054] = a[14] & g[23670];
assign g[56437] = b[14] & g[23670];
assign g[40055] = a[14] & g[23671];
assign g[56438] = b[14] & g[23671];
assign g[40056] = a[14] & g[23672];
assign g[56439] = b[14] & g[23672];
assign g[40057] = a[14] & g[23673];
assign g[56440] = b[14] & g[23673];
assign g[40058] = a[14] & g[23674];
assign g[56441] = b[14] & g[23674];
assign g[40059] = a[14] & g[23675];
assign g[56442] = b[14] & g[23675];
assign g[40060] = a[14] & g[23676];
assign g[56443] = b[14] & g[23676];
assign g[40061] = a[14] & g[23677];
assign g[56444] = b[14] & g[23677];
assign g[40062] = a[14] & g[23678];
assign g[56445] = b[14] & g[23678];
assign g[40063] = a[14] & g[23679];
assign g[56446] = b[14] & g[23679];
assign g[40064] = a[14] & g[23680];
assign g[56447] = b[14] & g[23680];
assign g[40065] = a[14] & g[23681];
assign g[56448] = b[14] & g[23681];
assign g[40066] = a[14] & g[23682];
assign g[56449] = b[14] & g[23682];
assign g[40067] = a[14] & g[23683];
assign g[56450] = b[14] & g[23683];
assign g[40068] = a[14] & g[23684];
assign g[56451] = b[14] & g[23684];
assign g[40069] = a[14] & g[23685];
assign g[56452] = b[14] & g[23685];
assign g[40070] = a[14] & g[23686];
assign g[56453] = b[14] & g[23686];
assign g[40071] = a[14] & g[23687];
assign g[56454] = b[14] & g[23687];
assign g[40072] = a[14] & g[23688];
assign g[56455] = b[14] & g[23688];
assign g[40073] = a[14] & g[23689];
assign g[56456] = b[14] & g[23689];
assign g[40074] = a[14] & g[23690];
assign g[56457] = b[14] & g[23690];
assign g[40075] = a[14] & g[23691];
assign g[56458] = b[14] & g[23691];
assign g[40076] = a[14] & g[23692];
assign g[56459] = b[14] & g[23692];
assign g[40077] = a[14] & g[23693];
assign g[56460] = b[14] & g[23693];
assign g[40078] = a[14] & g[23694];
assign g[56461] = b[14] & g[23694];
assign g[40079] = a[14] & g[23695];
assign g[56462] = b[14] & g[23695];
assign g[40080] = a[14] & g[23696];
assign g[56463] = b[14] & g[23696];
assign g[40081] = a[14] & g[23697];
assign g[56464] = b[14] & g[23697];
assign g[40082] = a[14] & g[23698];
assign g[56465] = b[14] & g[23698];
assign g[40083] = a[14] & g[23699];
assign g[56466] = b[14] & g[23699];
assign g[40084] = a[14] & g[23700];
assign g[56467] = b[14] & g[23700];
assign g[40085] = a[14] & g[23701];
assign g[56468] = b[14] & g[23701];
assign g[40086] = a[14] & g[23702];
assign g[56469] = b[14] & g[23702];
assign g[40087] = a[14] & g[23703];
assign g[56470] = b[14] & g[23703];
assign g[40088] = a[14] & g[23704];
assign g[56471] = b[14] & g[23704];
assign g[40089] = a[14] & g[23705];
assign g[56472] = b[14] & g[23705];
assign g[40090] = a[14] & g[23706];
assign g[56473] = b[14] & g[23706];
assign g[40091] = a[14] & g[23707];
assign g[56474] = b[14] & g[23707];
assign g[40092] = a[14] & g[23708];
assign g[56475] = b[14] & g[23708];
assign g[40093] = a[14] & g[23709];
assign g[56476] = b[14] & g[23709];
assign g[40094] = a[14] & g[23710];
assign g[56477] = b[14] & g[23710];
assign g[40095] = a[14] & g[23711];
assign g[56478] = b[14] & g[23711];
assign g[40096] = a[14] & g[23712];
assign g[56479] = b[14] & g[23712];
assign g[40097] = a[14] & g[23713];
assign g[56480] = b[14] & g[23713];
assign g[40098] = a[14] & g[23714];
assign g[56481] = b[14] & g[23714];
assign g[40099] = a[14] & g[23715];
assign g[56482] = b[14] & g[23715];
assign g[40100] = a[14] & g[23716];
assign g[56483] = b[14] & g[23716];
assign g[40101] = a[14] & g[23717];
assign g[56484] = b[14] & g[23717];
assign g[40102] = a[14] & g[23718];
assign g[56485] = b[14] & g[23718];
assign g[40103] = a[14] & g[23719];
assign g[56486] = b[14] & g[23719];
assign g[40104] = a[14] & g[23720];
assign g[56487] = b[14] & g[23720];
assign g[40105] = a[14] & g[23721];
assign g[56488] = b[14] & g[23721];
assign g[40106] = a[14] & g[23722];
assign g[56489] = b[14] & g[23722];
assign g[40107] = a[14] & g[23723];
assign g[56490] = b[14] & g[23723];
assign g[40108] = a[14] & g[23724];
assign g[56491] = b[14] & g[23724];
assign g[40109] = a[14] & g[23725];
assign g[56492] = b[14] & g[23725];
assign g[40110] = a[14] & g[23726];
assign g[56493] = b[14] & g[23726];
assign g[40111] = a[14] & g[23727];
assign g[56494] = b[14] & g[23727];
assign g[40112] = a[14] & g[23728];
assign g[56495] = b[14] & g[23728];
assign g[40113] = a[14] & g[23729];
assign g[56496] = b[14] & g[23729];
assign g[40114] = a[14] & g[23730];
assign g[56497] = b[14] & g[23730];
assign g[40115] = a[14] & g[23731];
assign g[56498] = b[14] & g[23731];
assign g[40116] = a[14] & g[23732];
assign g[56499] = b[14] & g[23732];
assign g[40117] = a[14] & g[23733];
assign g[56500] = b[14] & g[23733];
assign g[40118] = a[14] & g[23734];
assign g[56501] = b[14] & g[23734];
assign g[40119] = a[14] & g[23735];
assign g[56502] = b[14] & g[23735];
assign g[40120] = a[14] & g[23736];
assign g[56503] = b[14] & g[23736];
assign g[40121] = a[14] & g[23737];
assign g[56504] = b[14] & g[23737];
assign g[40122] = a[14] & g[23738];
assign g[56505] = b[14] & g[23738];
assign g[40123] = a[14] & g[23739];
assign g[56506] = b[14] & g[23739];
assign g[40124] = a[14] & g[23740];
assign g[56507] = b[14] & g[23740];
assign g[40125] = a[14] & g[23741];
assign g[56508] = b[14] & g[23741];
assign g[40126] = a[14] & g[23742];
assign g[56509] = b[14] & g[23742];
assign g[40127] = a[14] & g[23743];
assign g[56510] = b[14] & g[23743];
assign g[40128] = a[14] & g[23744];
assign g[56511] = b[14] & g[23744];
assign g[40129] = a[14] & g[23745];
assign g[56512] = b[14] & g[23745];
assign g[40130] = a[14] & g[23746];
assign g[56513] = b[14] & g[23746];
assign g[40131] = a[14] & g[23747];
assign g[56514] = b[14] & g[23747];
assign g[40132] = a[14] & g[23748];
assign g[56515] = b[14] & g[23748];
assign g[40133] = a[14] & g[23749];
assign g[56516] = b[14] & g[23749];
assign g[40134] = a[14] & g[23750];
assign g[56517] = b[14] & g[23750];
assign g[40135] = a[14] & g[23751];
assign g[56518] = b[14] & g[23751];
assign g[40136] = a[14] & g[23752];
assign g[56519] = b[14] & g[23752];
assign g[40137] = a[14] & g[23753];
assign g[56520] = b[14] & g[23753];
assign g[40138] = a[14] & g[23754];
assign g[56521] = b[14] & g[23754];
assign g[40139] = a[14] & g[23755];
assign g[56522] = b[14] & g[23755];
assign g[40140] = a[14] & g[23756];
assign g[56523] = b[14] & g[23756];
assign g[40141] = a[14] & g[23757];
assign g[56524] = b[14] & g[23757];
assign g[40142] = a[14] & g[23758];
assign g[56525] = b[14] & g[23758];
assign g[40143] = a[14] & g[23759];
assign g[56526] = b[14] & g[23759];
assign g[40144] = a[14] & g[23760];
assign g[56527] = b[14] & g[23760];
assign g[40145] = a[14] & g[23761];
assign g[56528] = b[14] & g[23761];
assign g[40146] = a[14] & g[23762];
assign g[56529] = b[14] & g[23762];
assign g[40147] = a[14] & g[23763];
assign g[56530] = b[14] & g[23763];
assign g[40148] = a[14] & g[23764];
assign g[56531] = b[14] & g[23764];
assign g[40149] = a[14] & g[23765];
assign g[56532] = b[14] & g[23765];
assign g[40150] = a[14] & g[23766];
assign g[56533] = b[14] & g[23766];
assign g[40151] = a[14] & g[23767];
assign g[56534] = b[14] & g[23767];
assign g[40152] = a[14] & g[23768];
assign g[56535] = b[14] & g[23768];
assign g[40153] = a[14] & g[23769];
assign g[56536] = b[14] & g[23769];
assign g[40154] = a[14] & g[23770];
assign g[56537] = b[14] & g[23770];
assign g[40155] = a[14] & g[23771];
assign g[56538] = b[14] & g[23771];
assign g[40156] = a[14] & g[23772];
assign g[56539] = b[14] & g[23772];
assign g[40157] = a[14] & g[23773];
assign g[56540] = b[14] & g[23773];
assign g[40158] = a[14] & g[23774];
assign g[56541] = b[14] & g[23774];
assign g[40159] = a[14] & g[23775];
assign g[56542] = b[14] & g[23775];
assign g[40160] = a[14] & g[23776];
assign g[56543] = b[14] & g[23776];
assign g[40161] = a[14] & g[23777];
assign g[56544] = b[14] & g[23777];
assign g[40162] = a[14] & g[23778];
assign g[56545] = b[14] & g[23778];
assign g[40163] = a[14] & g[23779];
assign g[56546] = b[14] & g[23779];
assign g[40164] = a[14] & g[23780];
assign g[56547] = b[14] & g[23780];
assign g[40165] = a[14] & g[23781];
assign g[56548] = b[14] & g[23781];
assign g[40166] = a[14] & g[23782];
assign g[56549] = b[14] & g[23782];
assign g[40167] = a[14] & g[23783];
assign g[56550] = b[14] & g[23783];
assign g[40168] = a[14] & g[23784];
assign g[56551] = b[14] & g[23784];
assign g[40169] = a[14] & g[23785];
assign g[56552] = b[14] & g[23785];
assign g[40170] = a[14] & g[23786];
assign g[56553] = b[14] & g[23786];
assign g[40171] = a[14] & g[23787];
assign g[56554] = b[14] & g[23787];
assign g[40172] = a[14] & g[23788];
assign g[56555] = b[14] & g[23788];
assign g[40173] = a[14] & g[23789];
assign g[56556] = b[14] & g[23789];
assign g[40174] = a[14] & g[23790];
assign g[56557] = b[14] & g[23790];
assign g[40175] = a[14] & g[23791];
assign g[56558] = b[14] & g[23791];
assign g[40176] = a[14] & g[23792];
assign g[56559] = b[14] & g[23792];
assign g[40177] = a[14] & g[23793];
assign g[56560] = b[14] & g[23793];
assign g[40178] = a[14] & g[23794];
assign g[56561] = b[14] & g[23794];
assign g[40179] = a[14] & g[23795];
assign g[56562] = b[14] & g[23795];
assign g[40180] = a[14] & g[23796];
assign g[56563] = b[14] & g[23796];
assign g[40181] = a[14] & g[23797];
assign g[56564] = b[14] & g[23797];
assign g[40182] = a[14] & g[23798];
assign g[56565] = b[14] & g[23798];
assign g[40183] = a[14] & g[23799];
assign g[56566] = b[14] & g[23799];
assign g[40184] = a[14] & g[23800];
assign g[56567] = b[14] & g[23800];
assign g[40185] = a[14] & g[23801];
assign g[56568] = b[14] & g[23801];
assign g[40186] = a[14] & g[23802];
assign g[56569] = b[14] & g[23802];
assign g[40187] = a[14] & g[23803];
assign g[56570] = b[14] & g[23803];
assign g[40188] = a[14] & g[23804];
assign g[56571] = b[14] & g[23804];
assign g[40189] = a[14] & g[23805];
assign g[56572] = b[14] & g[23805];
assign g[40190] = a[14] & g[23806];
assign g[56573] = b[14] & g[23806];
assign g[40191] = a[14] & g[23807];
assign g[56574] = b[14] & g[23807];
assign g[40192] = a[14] & g[23808];
assign g[56575] = b[14] & g[23808];
assign g[40193] = a[14] & g[23809];
assign g[56576] = b[14] & g[23809];
assign g[40194] = a[14] & g[23810];
assign g[56577] = b[14] & g[23810];
assign g[40195] = a[14] & g[23811];
assign g[56578] = b[14] & g[23811];
assign g[40196] = a[14] & g[23812];
assign g[56579] = b[14] & g[23812];
assign g[40197] = a[14] & g[23813];
assign g[56580] = b[14] & g[23813];
assign g[40198] = a[14] & g[23814];
assign g[56581] = b[14] & g[23814];
assign g[40199] = a[14] & g[23815];
assign g[56582] = b[14] & g[23815];
assign g[40200] = a[14] & g[23816];
assign g[56583] = b[14] & g[23816];
assign g[40201] = a[14] & g[23817];
assign g[56584] = b[14] & g[23817];
assign g[40202] = a[14] & g[23818];
assign g[56585] = b[14] & g[23818];
assign g[40203] = a[14] & g[23819];
assign g[56586] = b[14] & g[23819];
assign g[40204] = a[14] & g[23820];
assign g[56587] = b[14] & g[23820];
assign g[40205] = a[14] & g[23821];
assign g[56588] = b[14] & g[23821];
assign g[40206] = a[14] & g[23822];
assign g[56589] = b[14] & g[23822];
assign g[40207] = a[14] & g[23823];
assign g[56590] = b[14] & g[23823];
assign g[40208] = a[14] & g[23824];
assign g[56591] = b[14] & g[23824];
assign g[40209] = a[14] & g[23825];
assign g[56592] = b[14] & g[23825];
assign g[40210] = a[14] & g[23826];
assign g[56593] = b[14] & g[23826];
assign g[40211] = a[14] & g[23827];
assign g[56594] = b[14] & g[23827];
assign g[40212] = a[14] & g[23828];
assign g[56595] = b[14] & g[23828];
assign g[40213] = a[14] & g[23829];
assign g[56596] = b[14] & g[23829];
assign g[40214] = a[14] & g[23830];
assign g[56597] = b[14] & g[23830];
assign g[40215] = a[14] & g[23831];
assign g[56598] = b[14] & g[23831];
assign g[40216] = a[14] & g[23832];
assign g[56599] = b[14] & g[23832];
assign g[40217] = a[14] & g[23833];
assign g[56600] = b[14] & g[23833];
assign g[40218] = a[14] & g[23834];
assign g[56601] = b[14] & g[23834];
assign g[40219] = a[14] & g[23835];
assign g[56602] = b[14] & g[23835];
assign g[40220] = a[14] & g[23836];
assign g[56603] = b[14] & g[23836];
assign g[40221] = a[14] & g[23837];
assign g[56604] = b[14] & g[23837];
assign g[40222] = a[14] & g[23838];
assign g[56605] = b[14] & g[23838];
assign g[40223] = a[14] & g[23839];
assign g[56606] = b[14] & g[23839];
assign g[40224] = a[14] & g[23840];
assign g[56607] = b[14] & g[23840];
assign g[40225] = a[14] & g[23841];
assign g[56608] = b[14] & g[23841];
assign g[40226] = a[14] & g[23842];
assign g[56609] = b[14] & g[23842];
assign g[40227] = a[14] & g[23843];
assign g[56610] = b[14] & g[23843];
assign g[40228] = a[14] & g[23844];
assign g[56611] = b[14] & g[23844];
assign g[40229] = a[14] & g[23845];
assign g[56612] = b[14] & g[23845];
assign g[40230] = a[14] & g[23846];
assign g[56613] = b[14] & g[23846];
assign g[40231] = a[14] & g[23847];
assign g[56614] = b[14] & g[23847];
assign g[40232] = a[14] & g[23848];
assign g[56615] = b[14] & g[23848];
assign g[40233] = a[14] & g[23849];
assign g[56616] = b[14] & g[23849];
assign g[40234] = a[14] & g[23850];
assign g[56617] = b[14] & g[23850];
assign g[40235] = a[14] & g[23851];
assign g[56618] = b[14] & g[23851];
assign g[40236] = a[14] & g[23852];
assign g[56619] = b[14] & g[23852];
assign g[40237] = a[14] & g[23853];
assign g[56620] = b[14] & g[23853];
assign g[40238] = a[14] & g[23854];
assign g[56621] = b[14] & g[23854];
assign g[40239] = a[14] & g[23855];
assign g[56622] = b[14] & g[23855];
assign g[40240] = a[14] & g[23856];
assign g[56623] = b[14] & g[23856];
assign g[40241] = a[14] & g[23857];
assign g[56624] = b[14] & g[23857];
assign g[40242] = a[14] & g[23858];
assign g[56625] = b[14] & g[23858];
assign g[40243] = a[14] & g[23859];
assign g[56626] = b[14] & g[23859];
assign g[40244] = a[14] & g[23860];
assign g[56627] = b[14] & g[23860];
assign g[40245] = a[14] & g[23861];
assign g[56628] = b[14] & g[23861];
assign g[40246] = a[14] & g[23862];
assign g[56629] = b[14] & g[23862];
assign g[40247] = a[14] & g[23863];
assign g[56630] = b[14] & g[23863];
assign g[40248] = a[14] & g[23864];
assign g[56631] = b[14] & g[23864];
assign g[40249] = a[14] & g[23865];
assign g[56632] = b[14] & g[23865];
assign g[40250] = a[14] & g[23866];
assign g[56633] = b[14] & g[23866];
assign g[40251] = a[14] & g[23867];
assign g[56634] = b[14] & g[23867];
assign g[40252] = a[14] & g[23868];
assign g[56635] = b[14] & g[23868];
assign g[40253] = a[14] & g[23869];
assign g[56636] = b[14] & g[23869];
assign g[40254] = a[14] & g[23870];
assign g[56637] = b[14] & g[23870];
assign g[40255] = a[14] & g[23871];
assign g[56638] = b[14] & g[23871];
assign g[40256] = a[14] & g[23872];
assign g[56639] = b[14] & g[23872];
assign g[40257] = a[14] & g[23873];
assign g[56640] = b[14] & g[23873];
assign g[40258] = a[14] & g[23874];
assign g[56641] = b[14] & g[23874];
assign g[40259] = a[14] & g[23875];
assign g[56642] = b[14] & g[23875];
assign g[40260] = a[14] & g[23876];
assign g[56643] = b[14] & g[23876];
assign g[40261] = a[14] & g[23877];
assign g[56644] = b[14] & g[23877];
assign g[40262] = a[14] & g[23878];
assign g[56645] = b[14] & g[23878];
assign g[40263] = a[14] & g[23879];
assign g[56646] = b[14] & g[23879];
assign g[40264] = a[14] & g[23880];
assign g[56647] = b[14] & g[23880];
assign g[40265] = a[14] & g[23881];
assign g[56648] = b[14] & g[23881];
assign g[40266] = a[14] & g[23882];
assign g[56649] = b[14] & g[23882];
assign g[40267] = a[14] & g[23883];
assign g[56650] = b[14] & g[23883];
assign g[40268] = a[14] & g[23884];
assign g[56651] = b[14] & g[23884];
assign g[40269] = a[14] & g[23885];
assign g[56652] = b[14] & g[23885];
assign g[40270] = a[14] & g[23886];
assign g[56653] = b[14] & g[23886];
assign g[40271] = a[14] & g[23887];
assign g[56654] = b[14] & g[23887];
assign g[40272] = a[14] & g[23888];
assign g[56655] = b[14] & g[23888];
assign g[40273] = a[14] & g[23889];
assign g[56656] = b[14] & g[23889];
assign g[40274] = a[14] & g[23890];
assign g[56657] = b[14] & g[23890];
assign g[40275] = a[14] & g[23891];
assign g[56658] = b[14] & g[23891];
assign g[40276] = a[14] & g[23892];
assign g[56659] = b[14] & g[23892];
assign g[40277] = a[14] & g[23893];
assign g[56660] = b[14] & g[23893];
assign g[40278] = a[14] & g[23894];
assign g[56661] = b[14] & g[23894];
assign g[40279] = a[14] & g[23895];
assign g[56662] = b[14] & g[23895];
assign g[40280] = a[14] & g[23896];
assign g[56663] = b[14] & g[23896];
assign g[40281] = a[14] & g[23897];
assign g[56664] = b[14] & g[23897];
assign g[40282] = a[14] & g[23898];
assign g[56665] = b[14] & g[23898];
assign g[40283] = a[14] & g[23899];
assign g[56666] = b[14] & g[23899];
assign g[40284] = a[14] & g[23900];
assign g[56667] = b[14] & g[23900];
assign g[40285] = a[14] & g[23901];
assign g[56668] = b[14] & g[23901];
assign g[40286] = a[14] & g[23902];
assign g[56669] = b[14] & g[23902];
assign g[40287] = a[14] & g[23903];
assign g[56670] = b[14] & g[23903];
assign g[40288] = a[14] & g[23904];
assign g[56671] = b[14] & g[23904];
assign g[40289] = a[14] & g[23905];
assign g[56672] = b[14] & g[23905];
assign g[40290] = a[14] & g[23906];
assign g[56673] = b[14] & g[23906];
assign g[40291] = a[14] & g[23907];
assign g[56674] = b[14] & g[23907];
assign g[40292] = a[14] & g[23908];
assign g[56675] = b[14] & g[23908];
assign g[40293] = a[14] & g[23909];
assign g[56676] = b[14] & g[23909];
assign g[40294] = a[14] & g[23910];
assign g[56677] = b[14] & g[23910];
assign g[40295] = a[14] & g[23911];
assign g[56678] = b[14] & g[23911];
assign g[40296] = a[14] & g[23912];
assign g[56679] = b[14] & g[23912];
assign g[40297] = a[14] & g[23913];
assign g[56680] = b[14] & g[23913];
assign g[40298] = a[14] & g[23914];
assign g[56681] = b[14] & g[23914];
assign g[40299] = a[14] & g[23915];
assign g[56682] = b[14] & g[23915];
assign g[40300] = a[14] & g[23916];
assign g[56683] = b[14] & g[23916];
assign g[40301] = a[14] & g[23917];
assign g[56684] = b[14] & g[23917];
assign g[40302] = a[14] & g[23918];
assign g[56685] = b[14] & g[23918];
assign g[40303] = a[14] & g[23919];
assign g[56686] = b[14] & g[23919];
assign g[40304] = a[14] & g[23920];
assign g[56687] = b[14] & g[23920];
assign g[40305] = a[14] & g[23921];
assign g[56688] = b[14] & g[23921];
assign g[40306] = a[14] & g[23922];
assign g[56689] = b[14] & g[23922];
assign g[40307] = a[14] & g[23923];
assign g[56690] = b[14] & g[23923];
assign g[40308] = a[14] & g[23924];
assign g[56691] = b[14] & g[23924];
assign g[40309] = a[14] & g[23925];
assign g[56692] = b[14] & g[23925];
assign g[40310] = a[14] & g[23926];
assign g[56693] = b[14] & g[23926];
assign g[40311] = a[14] & g[23927];
assign g[56694] = b[14] & g[23927];
assign g[40312] = a[14] & g[23928];
assign g[56695] = b[14] & g[23928];
assign g[40313] = a[14] & g[23929];
assign g[56696] = b[14] & g[23929];
assign g[40314] = a[14] & g[23930];
assign g[56697] = b[14] & g[23930];
assign g[40315] = a[14] & g[23931];
assign g[56698] = b[14] & g[23931];
assign g[40316] = a[14] & g[23932];
assign g[56699] = b[14] & g[23932];
assign g[40317] = a[14] & g[23933];
assign g[56700] = b[14] & g[23933];
assign g[40318] = a[14] & g[23934];
assign g[56701] = b[14] & g[23934];
assign g[40319] = a[14] & g[23935];
assign g[56702] = b[14] & g[23935];
assign g[40320] = a[14] & g[23936];
assign g[56703] = b[14] & g[23936];
assign g[40321] = a[14] & g[23937];
assign g[56704] = b[14] & g[23937];
assign g[40322] = a[14] & g[23938];
assign g[56705] = b[14] & g[23938];
assign g[40323] = a[14] & g[23939];
assign g[56706] = b[14] & g[23939];
assign g[40324] = a[14] & g[23940];
assign g[56707] = b[14] & g[23940];
assign g[40325] = a[14] & g[23941];
assign g[56708] = b[14] & g[23941];
assign g[40326] = a[14] & g[23942];
assign g[56709] = b[14] & g[23942];
assign g[40327] = a[14] & g[23943];
assign g[56710] = b[14] & g[23943];
assign g[40328] = a[14] & g[23944];
assign g[56711] = b[14] & g[23944];
assign g[40329] = a[14] & g[23945];
assign g[56712] = b[14] & g[23945];
assign g[40330] = a[14] & g[23946];
assign g[56713] = b[14] & g[23946];
assign g[40331] = a[14] & g[23947];
assign g[56714] = b[14] & g[23947];
assign g[40332] = a[14] & g[23948];
assign g[56715] = b[14] & g[23948];
assign g[40333] = a[14] & g[23949];
assign g[56716] = b[14] & g[23949];
assign g[40334] = a[14] & g[23950];
assign g[56717] = b[14] & g[23950];
assign g[40335] = a[14] & g[23951];
assign g[56718] = b[14] & g[23951];
assign g[40336] = a[14] & g[23952];
assign g[56719] = b[14] & g[23952];
assign g[40337] = a[14] & g[23953];
assign g[56720] = b[14] & g[23953];
assign g[40338] = a[14] & g[23954];
assign g[56721] = b[14] & g[23954];
assign g[40339] = a[14] & g[23955];
assign g[56722] = b[14] & g[23955];
assign g[40340] = a[14] & g[23956];
assign g[56723] = b[14] & g[23956];
assign g[40341] = a[14] & g[23957];
assign g[56724] = b[14] & g[23957];
assign g[40342] = a[14] & g[23958];
assign g[56725] = b[14] & g[23958];
assign g[40343] = a[14] & g[23959];
assign g[56726] = b[14] & g[23959];
assign g[40344] = a[14] & g[23960];
assign g[56727] = b[14] & g[23960];
assign g[40345] = a[14] & g[23961];
assign g[56728] = b[14] & g[23961];
assign g[40346] = a[14] & g[23962];
assign g[56729] = b[14] & g[23962];
assign g[40347] = a[14] & g[23963];
assign g[56730] = b[14] & g[23963];
assign g[40348] = a[14] & g[23964];
assign g[56731] = b[14] & g[23964];
assign g[40349] = a[14] & g[23965];
assign g[56732] = b[14] & g[23965];
assign g[40350] = a[14] & g[23966];
assign g[56733] = b[14] & g[23966];
assign g[40351] = a[14] & g[23967];
assign g[56734] = b[14] & g[23967];
assign g[40352] = a[14] & g[23968];
assign g[56735] = b[14] & g[23968];
assign g[40353] = a[14] & g[23969];
assign g[56736] = b[14] & g[23969];
assign g[40354] = a[14] & g[23970];
assign g[56737] = b[14] & g[23970];
assign g[40355] = a[14] & g[23971];
assign g[56738] = b[14] & g[23971];
assign g[40356] = a[14] & g[23972];
assign g[56739] = b[14] & g[23972];
assign g[40357] = a[14] & g[23973];
assign g[56740] = b[14] & g[23973];
assign g[40358] = a[14] & g[23974];
assign g[56741] = b[14] & g[23974];
assign g[40359] = a[14] & g[23975];
assign g[56742] = b[14] & g[23975];
assign g[40360] = a[14] & g[23976];
assign g[56743] = b[14] & g[23976];
assign g[40361] = a[14] & g[23977];
assign g[56744] = b[14] & g[23977];
assign g[40362] = a[14] & g[23978];
assign g[56745] = b[14] & g[23978];
assign g[40363] = a[14] & g[23979];
assign g[56746] = b[14] & g[23979];
assign g[40364] = a[14] & g[23980];
assign g[56747] = b[14] & g[23980];
assign g[40365] = a[14] & g[23981];
assign g[56748] = b[14] & g[23981];
assign g[40366] = a[14] & g[23982];
assign g[56749] = b[14] & g[23982];
assign g[40367] = a[14] & g[23983];
assign g[56750] = b[14] & g[23983];
assign g[40368] = a[14] & g[23984];
assign g[56751] = b[14] & g[23984];
assign g[40369] = a[14] & g[23985];
assign g[56752] = b[14] & g[23985];
assign g[40370] = a[14] & g[23986];
assign g[56753] = b[14] & g[23986];
assign g[40371] = a[14] & g[23987];
assign g[56754] = b[14] & g[23987];
assign g[40372] = a[14] & g[23988];
assign g[56755] = b[14] & g[23988];
assign g[40373] = a[14] & g[23989];
assign g[56756] = b[14] & g[23989];
assign g[40374] = a[14] & g[23990];
assign g[56757] = b[14] & g[23990];
assign g[40375] = a[14] & g[23991];
assign g[56758] = b[14] & g[23991];
assign g[40376] = a[14] & g[23992];
assign g[56759] = b[14] & g[23992];
assign g[40377] = a[14] & g[23993];
assign g[56760] = b[14] & g[23993];
assign g[40378] = a[14] & g[23994];
assign g[56761] = b[14] & g[23994];
assign g[40379] = a[14] & g[23995];
assign g[56762] = b[14] & g[23995];
assign g[40380] = a[14] & g[23996];
assign g[56763] = b[14] & g[23996];
assign g[40381] = a[14] & g[23997];
assign g[56764] = b[14] & g[23997];
assign g[40382] = a[14] & g[23998];
assign g[56765] = b[14] & g[23998];
assign g[40383] = a[14] & g[23999];
assign g[56766] = b[14] & g[23999];
assign g[40384] = a[14] & g[24000];
assign g[56767] = b[14] & g[24000];
assign g[40385] = a[14] & g[24001];
assign g[56768] = b[14] & g[24001];
assign g[40386] = a[14] & g[24002];
assign g[56769] = b[14] & g[24002];
assign g[40387] = a[14] & g[24003];
assign g[56770] = b[14] & g[24003];
assign g[40388] = a[14] & g[24004];
assign g[56771] = b[14] & g[24004];
assign g[40389] = a[14] & g[24005];
assign g[56772] = b[14] & g[24005];
assign g[40390] = a[14] & g[24006];
assign g[56773] = b[14] & g[24006];
assign g[40391] = a[14] & g[24007];
assign g[56774] = b[14] & g[24007];
assign g[40392] = a[14] & g[24008];
assign g[56775] = b[14] & g[24008];
assign g[40393] = a[14] & g[24009];
assign g[56776] = b[14] & g[24009];
assign g[40394] = a[14] & g[24010];
assign g[56777] = b[14] & g[24010];
assign g[40395] = a[14] & g[24011];
assign g[56778] = b[14] & g[24011];
assign g[40396] = a[14] & g[24012];
assign g[56779] = b[14] & g[24012];
assign g[40397] = a[14] & g[24013];
assign g[56780] = b[14] & g[24013];
assign g[40398] = a[14] & g[24014];
assign g[56781] = b[14] & g[24014];
assign g[40399] = a[14] & g[24015];
assign g[56782] = b[14] & g[24015];
assign g[40400] = a[14] & g[24016];
assign g[56783] = b[14] & g[24016];
assign g[40401] = a[14] & g[24017];
assign g[56784] = b[14] & g[24017];
assign g[40402] = a[14] & g[24018];
assign g[56785] = b[14] & g[24018];
assign g[40403] = a[14] & g[24019];
assign g[56786] = b[14] & g[24019];
assign g[40404] = a[14] & g[24020];
assign g[56787] = b[14] & g[24020];
assign g[40405] = a[14] & g[24021];
assign g[56788] = b[14] & g[24021];
assign g[40406] = a[14] & g[24022];
assign g[56789] = b[14] & g[24022];
assign g[40407] = a[14] & g[24023];
assign g[56790] = b[14] & g[24023];
assign g[40408] = a[14] & g[24024];
assign g[56791] = b[14] & g[24024];
assign g[40409] = a[14] & g[24025];
assign g[56792] = b[14] & g[24025];
assign g[40410] = a[14] & g[24026];
assign g[56793] = b[14] & g[24026];
assign g[40411] = a[14] & g[24027];
assign g[56794] = b[14] & g[24027];
assign g[40412] = a[14] & g[24028];
assign g[56795] = b[14] & g[24028];
assign g[40413] = a[14] & g[24029];
assign g[56796] = b[14] & g[24029];
assign g[40414] = a[14] & g[24030];
assign g[56797] = b[14] & g[24030];
assign g[40415] = a[14] & g[24031];
assign g[56798] = b[14] & g[24031];
assign g[40416] = a[14] & g[24032];
assign g[56799] = b[14] & g[24032];
assign g[40417] = a[14] & g[24033];
assign g[56800] = b[14] & g[24033];
assign g[40418] = a[14] & g[24034];
assign g[56801] = b[14] & g[24034];
assign g[40419] = a[14] & g[24035];
assign g[56802] = b[14] & g[24035];
assign g[40420] = a[14] & g[24036];
assign g[56803] = b[14] & g[24036];
assign g[40421] = a[14] & g[24037];
assign g[56804] = b[14] & g[24037];
assign g[40422] = a[14] & g[24038];
assign g[56805] = b[14] & g[24038];
assign g[40423] = a[14] & g[24039];
assign g[56806] = b[14] & g[24039];
assign g[40424] = a[14] & g[24040];
assign g[56807] = b[14] & g[24040];
assign g[40425] = a[14] & g[24041];
assign g[56808] = b[14] & g[24041];
assign g[40426] = a[14] & g[24042];
assign g[56809] = b[14] & g[24042];
assign g[40427] = a[14] & g[24043];
assign g[56810] = b[14] & g[24043];
assign g[40428] = a[14] & g[24044];
assign g[56811] = b[14] & g[24044];
assign g[40429] = a[14] & g[24045];
assign g[56812] = b[14] & g[24045];
assign g[40430] = a[14] & g[24046];
assign g[56813] = b[14] & g[24046];
assign g[40431] = a[14] & g[24047];
assign g[56814] = b[14] & g[24047];
assign g[40432] = a[14] & g[24048];
assign g[56815] = b[14] & g[24048];
assign g[40433] = a[14] & g[24049];
assign g[56816] = b[14] & g[24049];
assign g[40434] = a[14] & g[24050];
assign g[56817] = b[14] & g[24050];
assign g[40435] = a[14] & g[24051];
assign g[56818] = b[14] & g[24051];
assign g[40436] = a[14] & g[24052];
assign g[56819] = b[14] & g[24052];
assign g[40437] = a[14] & g[24053];
assign g[56820] = b[14] & g[24053];
assign g[40438] = a[14] & g[24054];
assign g[56821] = b[14] & g[24054];
assign g[40439] = a[14] & g[24055];
assign g[56822] = b[14] & g[24055];
assign g[40440] = a[14] & g[24056];
assign g[56823] = b[14] & g[24056];
assign g[40441] = a[14] & g[24057];
assign g[56824] = b[14] & g[24057];
assign g[40442] = a[14] & g[24058];
assign g[56825] = b[14] & g[24058];
assign g[40443] = a[14] & g[24059];
assign g[56826] = b[14] & g[24059];
assign g[40444] = a[14] & g[24060];
assign g[56827] = b[14] & g[24060];
assign g[40445] = a[14] & g[24061];
assign g[56828] = b[14] & g[24061];
assign g[40446] = a[14] & g[24062];
assign g[56829] = b[14] & g[24062];
assign g[40447] = a[14] & g[24063];
assign g[56830] = b[14] & g[24063];
assign g[40448] = a[14] & g[24064];
assign g[56831] = b[14] & g[24064];
assign g[40449] = a[14] & g[24065];
assign g[56832] = b[14] & g[24065];
assign g[40450] = a[14] & g[24066];
assign g[56833] = b[14] & g[24066];
assign g[40451] = a[14] & g[24067];
assign g[56834] = b[14] & g[24067];
assign g[40452] = a[14] & g[24068];
assign g[56835] = b[14] & g[24068];
assign g[40453] = a[14] & g[24069];
assign g[56836] = b[14] & g[24069];
assign g[40454] = a[14] & g[24070];
assign g[56837] = b[14] & g[24070];
assign g[40455] = a[14] & g[24071];
assign g[56838] = b[14] & g[24071];
assign g[40456] = a[14] & g[24072];
assign g[56839] = b[14] & g[24072];
assign g[40457] = a[14] & g[24073];
assign g[56840] = b[14] & g[24073];
assign g[40458] = a[14] & g[24074];
assign g[56841] = b[14] & g[24074];
assign g[40459] = a[14] & g[24075];
assign g[56842] = b[14] & g[24075];
assign g[40460] = a[14] & g[24076];
assign g[56843] = b[14] & g[24076];
assign g[40461] = a[14] & g[24077];
assign g[56844] = b[14] & g[24077];
assign g[40462] = a[14] & g[24078];
assign g[56845] = b[14] & g[24078];
assign g[40463] = a[14] & g[24079];
assign g[56846] = b[14] & g[24079];
assign g[40464] = a[14] & g[24080];
assign g[56847] = b[14] & g[24080];
assign g[40465] = a[14] & g[24081];
assign g[56848] = b[14] & g[24081];
assign g[40466] = a[14] & g[24082];
assign g[56849] = b[14] & g[24082];
assign g[40467] = a[14] & g[24083];
assign g[56850] = b[14] & g[24083];
assign g[40468] = a[14] & g[24084];
assign g[56851] = b[14] & g[24084];
assign g[40469] = a[14] & g[24085];
assign g[56852] = b[14] & g[24085];
assign g[40470] = a[14] & g[24086];
assign g[56853] = b[14] & g[24086];
assign g[40471] = a[14] & g[24087];
assign g[56854] = b[14] & g[24087];
assign g[40472] = a[14] & g[24088];
assign g[56855] = b[14] & g[24088];
assign g[40473] = a[14] & g[24089];
assign g[56856] = b[14] & g[24089];
assign g[40474] = a[14] & g[24090];
assign g[56857] = b[14] & g[24090];
assign g[40475] = a[14] & g[24091];
assign g[56858] = b[14] & g[24091];
assign g[40476] = a[14] & g[24092];
assign g[56859] = b[14] & g[24092];
assign g[40477] = a[14] & g[24093];
assign g[56860] = b[14] & g[24093];
assign g[40478] = a[14] & g[24094];
assign g[56861] = b[14] & g[24094];
assign g[40479] = a[14] & g[24095];
assign g[56862] = b[14] & g[24095];
assign g[40480] = a[14] & g[24096];
assign g[56863] = b[14] & g[24096];
assign g[40481] = a[14] & g[24097];
assign g[56864] = b[14] & g[24097];
assign g[40482] = a[14] & g[24098];
assign g[56865] = b[14] & g[24098];
assign g[40483] = a[14] & g[24099];
assign g[56866] = b[14] & g[24099];
assign g[40484] = a[14] & g[24100];
assign g[56867] = b[14] & g[24100];
assign g[40485] = a[14] & g[24101];
assign g[56868] = b[14] & g[24101];
assign g[40486] = a[14] & g[24102];
assign g[56869] = b[14] & g[24102];
assign g[40487] = a[14] & g[24103];
assign g[56870] = b[14] & g[24103];
assign g[40488] = a[14] & g[24104];
assign g[56871] = b[14] & g[24104];
assign g[40489] = a[14] & g[24105];
assign g[56872] = b[14] & g[24105];
assign g[40490] = a[14] & g[24106];
assign g[56873] = b[14] & g[24106];
assign g[40491] = a[14] & g[24107];
assign g[56874] = b[14] & g[24107];
assign g[40492] = a[14] & g[24108];
assign g[56875] = b[14] & g[24108];
assign g[40493] = a[14] & g[24109];
assign g[56876] = b[14] & g[24109];
assign g[40494] = a[14] & g[24110];
assign g[56877] = b[14] & g[24110];
assign g[40495] = a[14] & g[24111];
assign g[56878] = b[14] & g[24111];
assign g[40496] = a[14] & g[24112];
assign g[56879] = b[14] & g[24112];
assign g[40497] = a[14] & g[24113];
assign g[56880] = b[14] & g[24113];
assign g[40498] = a[14] & g[24114];
assign g[56881] = b[14] & g[24114];
assign g[40499] = a[14] & g[24115];
assign g[56882] = b[14] & g[24115];
assign g[40500] = a[14] & g[24116];
assign g[56883] = b[14] & g[24116];
assign g[40501] = a[14] & g[24117];
assign g[56884] = b[14] & g[24117];
assign g[40502] = a[14] & g[24118];
assign g[56885] = b[14] & g[24118];
assign g[40503] = a[14] & g[24119];
assign g[56886] = b[14] & g[24119];
assign g[40504] = a[14] & g[24120];
assign g[56887] = b[14] & g[24120];
assign g[40505] = a[14] & g[24121];
assign g[56888] = b[14] & g[24121];
assign g[40506] = a[14] & g[24122];
assign g[56889] = b[14] & g[24122];
assign g[40507] = a[14] & g[24123];
assign g[56890] = b[14] & g[24123];
assign g[40508] = a[14] & g[24124];
assign g[56891] = b[14] & g[24124];
assign g[40509] = a[14] & g[24125];
assign g[56892] = b[14] & g[24125];
assign g[40510] = a[14] & g[24126];
assign g[56893] = b[14] & g[24126];
assign g[40511] = a[14] & g[24127];
assign g[56894] = b[14] & g[24127];
assign g[40512] = a[14] & g[24128];
assign g[56895] = b[14] & g[24128];
assign g[40513] = a[14] & g[24129];
assign g[56896] = b[14] & g[24129];
assign g[40514] = a[14] & g[24130];
assign g[56897] = b[14] & g[24130];
assign g[40515] = a[14] & g[24131];
assign g[56898] = b[14] & g[24131];
assign g[40516] = a[14] & g[24132];
assign g[56899] = b[14] & g[24132];
assign g[40517] = a[14] & g[24133];
assign g[56900] = b[14] & g[24133];
assign g[40518] = a[14] & g[24134];
assign g[56901] = b[14] & g[24134];
assign g[40519] = a[14] & g[24135];
assign g[56902] = b[14] & g[24135];
assign g[40520] = a[14] & g[24136];
assign g[56903] = b[14] & g[24136];
assign g[40521] = a[14] & g[24137];
assign g[56904] = b[14] & g[24137];
assign g[40522] = a[14] & g[24138];
assign g[56905] = b[14] & g[24138];
assign g[40523] = a[14] & g[24139];
assign g[56906] = b[14] & g[24139];
assign g[40524] = a[14] & g[24140];
assign g[56907] = b[14] & g[24140];
assign g[40525] = a[14] & g[24141];
assign g[56908] = b[14] & g[24141];
assign g[40526] = a[14] & g[24142];
assign g[56909] = b[14] & g[24142];
assign g[40527] = a[14] & g[24143];
assign g[56910] = b[14] & g[24143];
assign g[40528] = a[14] & g[24144];
assign g[56911] = b[14] & g[24144];
assign g[40529] = a[14] & g[24145];
assign g[56912] = b[14] & g[24145];
assign g[40530] = a[14] & g[24146];
assign g[56913] = b[14] & g[24146];
assign g[40531] = a[14] & g[24147];
assign g[56914] = b[14] & g[24147];
assign g[40532] = a[14] & g[24148];
assign g[56915] = b[14] & g[24148];
assign g[40533] = a[14] & g[24149];
assign g[56916] = b[14] & g[24149];
assign g[40534] = a[14] & g[24150];
assign g[56917] = b[14] & g[24150];
assign g[40535] = a[14] & g[24151];
assign g[56918] = b[14] & g[24151];
assign g[40536] = a[14] & g[24152];
assign g[56919] = b[14] & g[24152];
assign g[40537] = a[14] & g[24153];
assign g[56920] = b[14] & g[24153];
assign g[40538] = a[14] & g[24154];
assign g[56921] = b[14] & g[24154];
assign g[40539] = a[14] & g[24155];
assign g[56922] = b[14] & g[24155];
assign g[40540] = a[14] & g[24156];
assign g[56923] = b[14] & g[24156];
assign g[40541] = a[14] & g[24157];
assign g[56924] = b[14] & g[24157];
assign g[40542] = a[14] & g[24158];
assign g[56925] = b[14] & g[24158];
assign g[40543] = a[14] & g[24159];
assign g[56926] = b[14] & g[24159];
assign g[40544] = a[14] & g[24160];
assign g[56927] = b[14] & g[24160];
assign g[40545] = a[14] & g[24161];
assign g[56928] = b[14] & g[24161];
assign g[40546] = a[14] & g[24162];
assign g[56929] = b[14] & g[24162];
assign g[40547] = a[14] & g[24163];
assign g[56930] = b[14] & g[24163];
assign g[40548] = a[14] & g[24164];
assign g[56931] = b[14] & g[24164];
assign g[40549] = a[14] & g[24165];
assign g[56932] = b[14] & g[24165];
assign g[40550] = a[14] & g[24166];
assign g[56933] = b[14] & g[24166];
assign g[40551] = a[14] & g[24167];
assign g[56934] = b[14] & g[24167];
assign g[40552] = a[14] & g[24168];
assign g[56935] = b[14] & g[24168];
assign g[40553] = a[14] & g[24169];
assign g[56936] = b[14] & g[24169];
assign g[40554] = a[14] & g[24170];
assign g[56937] = b[14] & g[24170];
assign g[40555] = a[14] & g[24171];
assign g[56938] = b[14] & g[24171];
assign g[40556] = a[14] & g[24172];
assign g[56939] = b[14] & g[24172];
assign g[40557] = a[14] & g[24173];
assign g[56940] = b[14] & g[24173];
assign g[40558] = a[14] & g[24174];
assign g[56941] = b[14] & g[24174];
assign g[40559] = a[14] & g[24175];
assign g[56942] = b[14] & g[24175];
assign g[40560] = a[14] & g[24176];
assign g[56943] = b[14] & g[24176];
assign g[40561] = a[14] & g[24177];
assign g[56944] = b[14] & g[24177];
assign g[40562] = a[14] & g[24178];
assign g[56945] = b[14] & g[24178];
assign g[40563] = a[14] & g[24179];
assign g[56946] = b[14] & g[24179];
assign g[40564] = a[14] & g[24180];
assign g[56947] = b[14] & g[24180];
assign g[40565] = a[14] & g[24181];
assign g[56948] = b[14] & g[24181];
assign g[40566] = a[14] & g[24182];
assign g[56949] = b[14] & g[24182];
assign g[40567] = a[14] & g[24183];
assign g[56950] = b[14] & g[24183];
assign g[40568] = a[14] & g[24184];
assign g[56951] = b[14] & g[24184];
assign g[40569] = a[14] & g[24185];
assign g[56952] = b[14] & g[24185];
assign g[40570] = a[14] & g[24186];
assign g[56953] = b[14] & g[24186];
assign g[40571] = a[14] & g[24187];
assign g[56954] = b[14] & g[24187];
assign g[40572] = a[14] & g[24188];
assign g[56955] = b[14] & g[24188];
assign g[40573] = a[14] & g[24189];
assign g[56956] = b[14] & g[24189];
assign g[40574] = a[14] & g[24190];
assign g[56957] = b[14] & g[24190];
assign g[40575] = a[14] & g[24191];
assign g[56958] = b[14] & g[24191];
assign g[40576] = a[14] & g[24192];
assign g[56959] = b[14] & g[24192];
assign g[40577] = a[14] & g[24193];
assign g[56960] = b[14] & g[24193];
assign g[40578] = a[14] & g[24194];
assign g[56961] = b[14] & g[24194];
assign g[40579] = a[14] & g[24195];
assign g[56962] = b[14] & g[24195];
assign g[40580] = a[14] & g[24196];
assign g[56963] = b[14] & g[24196];
assign g[40581] = a[14] & g[24197];
assign g[56964] = b[14] & g[24197];
assign g[40582] = a[14] & g[24198];
assign g[56965] = b[14] & g[24198];
assign g[40583] = a[14] & g[24199];
assign g[56966] = b[14] & g[24199];
assign g[40584] = a[14] & g[24200];
assign g[56967] = b[14] & g[24200];
assign g[40585] = a[14] & g[24201];
assign g[56968] = b[14] & g[24201];
assign g[40586] = a[14] & g[24202];
assign g[56969] = b[14] & g[24202];
assign g[40587] = a[14] & g[24203];
assign g[56970] = b[14] & g[24203];
assign g[40588] = a[14] & g[24204];
assign g[56971] = b[14] & g[24204];
assign g[40589] = a[14] & g[24205];
assign g[56972] = b[14] & g[24205];
assign g[40590] = a[14] & g[24206];
assign g[56973] = b[14] & g[24206];
assign g[40591] = a[14] & g[24207];
assign g[56974] = b[14] & g[24207];
assign g[40592] = a[14] & g[24208];
assign g[56975] = b[14] & g[24208];
assign g[40593] = a[14] & g[24209];
assign g[56976] = b[14] & g[24209];
assign g[40594] = a[14] & g[24210];
assign g[56977] = b[14] & g[24210];
assign g[40595] = a[14] & g[24211];
assign g[56978] = b[14] & g[24211];
assign g[40596] = a[14] & g[24212];
assign g[56979] = b[14] & g[24212];
assign g[40597] = a[14] & g[24213];
assign g[56980] = b[14] & g[24213];
assign g[40598] = a[14] & g[24214];
assign g[56981] = b[14] & g[24214];
assign g[40599] = a[14] & g[24215];
assign g[56982] = b[14] & g[24215];
assign g[40600] = a[14] & g[24216];
assign g[56983] = b[14] & g[24216];
assign g[40601] = a[14] & g[24217];
assign g[56984] = b[14] & g[24217];
assign g[40602] = a[14] & g[24218];
assign g[56985] = b[14] & g[24218];
assign g[40603] = a[14] & g[24219];
assign g[56986] = b[14] & g[24219];
assign g[40604] = a[14] & g[24220];
assign g[56987] = b[14] & g[24220];
assign g[40605] = a[14] & g[24221];
assign g[56988] = b[14] & g[24221];
assign g[40606] = a[14] & g[24222];
assign g[56989] = b[14] & g[24222];
assign g[40607] = a[14] & g[24223];
assign g[56990] = b[14] & g[24223];
assign g[40608] = a[14] & g[24224];
assign g[56991] = b[14] & g[24224];
assign g[40609] = a[14] & g[24225];
assign g[56992] = b[14] & g[24225];
assign g[40610] = a[14] & g[24226];
assign g[56993] = b[14] & g[24226];
assign g[40611] = a[14] & g[24227];
assign g[56994] = b[14] & g[24227];
assign g[40612] = a[14] & g[24228];
assign g[56995] = b[14] & g[24228];
assign g[40613] = a[14] & g[24229];
assign g[56996] = b[14] & g[24229];
assign g[40614] = a[14] & g[24230];
assign g[56997] = b[14] & g[24230];
assign g[40615] = a[14] & g[24231];
assign g[56998] = b[14] & g[24231];
assign g[40616] = a[14] & g[24232];
assign g[56999] = b[14] & g[24232];
assign g[40617] = a[14] & g[24233];
assign g[57000] = b[14] & g[24233];
assign g[40618] = a[14] & g[24234];
assign g[57001] = b[14] & g[24234];
assign g[40619] = a[14] & g[24235];
assign g[57002] = b[14] & g[24235];
assign g[40620] = a[14] & g[24236];
assign g[57003] = b[14] & g[24236];
assign g[40621] = a[14] & g[24237];
assign g[57004] = b[14] & g[24237];
assign g[40622] = a[14] & g[24238];
assign g[57005] = b[14] & g[24238];
assign g[40623] = a[14] & g[24239];
assign g[57006] = b[14] & g[24239];
assign g[40624] = a[14] & g[24240];
assign g[57007] = b[14] & g[24240];
assign g[40625] = a[14] & g[24241];
assign g[57008] = b[14] & g[24241];
assign g[40626] = a[14] & g[24242];
assign g[57009] = b[14] & g[24242];
assign g[40627] = a[14] & g[24243];
assign g[57010] = b[14] & g[24243];
assign g[40628] = a[14] & g[24244];
assign g[57011] = b[14] & g[24244];
assign g[40629] = a[14] & g[24245];
assign g[57012] = b[14] & g[24245];
assign g[40630] = a[14] & g[24246];
assign g[57013] = b[14] & g[24246];
assign g[40631] = a[14] & g[24247];
assign g[57014] = b[14] & g[24247];
assign g[40632] = a[14] & g[24248];
assign g[57015] = b[14] & g[24248];
assign g[40633] = a[14] & g[24249];
assign g[57016] = b[14] & g[24249];
assign g[40634] = a[14] & g[24250];
assign g[57017] = b[14] & g[24250];
assign g[40635] = a[14] & g[24251];
assign g[57018] = b[14] & g[24251];
assign g[40636] = a[14] & g[24252];
assign g[57019] = b[14] & g[24252];
assign g[40637] = a[14] & g[24253];
assign g[57020] = b[14] & g[24253];
assign g[40638] = a[14] & g[24254];
assign g[57021] = b[14] & g[24254];
assign g[40639] = a[14] & g[24255];
assign g[57022] = b[14] & g[24255];
assign g[40640] = a[14] & g[24256];
assign g[57023] = b[14] & g[24256];
assign g[40641] = a[14] & g[24257];
assign g[57024] = b[14] & g[24257];
assign g[40642] = a[14] & g[24258];
assign g[57025] = b[14] & g[24258];
assign g[40643] = a[14] & g[24259];
assign g[57026] = b[14] & g[24259];
assign g[40644] = a[14] & g[24260];
assign g[57027] = b[14] & g[24260];
assign g[40645] = a[14] & g[24261];
assign g[57028] = b[14] & g[24261];
assign g[40646] = a[14] & g[24262];
assign g[57029] = b[14] & g[24262];
assign g[40647] = a[14] & g[24263];
assign g[57030] = b[14] & g[24263];
assign g[40648] = a[14] & g[24264];
assign g[57031] = b[14] & g[24264];
assign g[40649] = a[14] & g[24265];
assign g[57032] = b[14] & g[24265];
assign g[40650] = a[14] & g[24266];
assign g[57033] = b[14] & g[24266];
assign g[40651] = a[14] & g[24267];
assign g[57034] = b[14] & g[24267];
assign g[40652] = a[14] & g[24268];
assign g[57035] = b[14] & g[24268];
assign g[40653] = a[14] & g[24269];
assign g[57036] = b[14] & g[24269];
assign g[40654] = a[14] & g[24270];
assign g[57037] = b[14] & g[24270];
assign g[40655] = a[14] & g[24271];
assign g[57038] = b[14] & g[24271];
assign g[40656] = a[14] & g[24272];
assign g[57039] = b[14] & g[24272];
assign g[40657] = a[14] & g[24273];
assign g[57040] = b[14] & g[24273];
assign g[40658] = a[14] & g[24274];
assign g[57041] = b[14] & g[24274];
assign g[40659] = a[14] & g[24275];
assign g[57042] = b[14] & g[24275];
assign g[40660] = a[14] & g[24276];
assign g[57043] = b[14] & g[24276];
assign g[40661] = a[14] & g[24277];
assign g[57044] = b[14] & g[24277];
assign g[40662] = a[14] & g[24278];
assign g[57045] = b[14] & g[24278];
assign g[40663] = a[14] & g[24279];
assign g[57046] = b[14] & g[24279];
assign g[40664] = a[14] & g[24280];
assign g[57047] = b[14] & g[24280];
assign g[40665] = a[14] & g[24281];
assign g[57048] = b[14] & g[24281];
assign g[40666] = a[14] & g[24282];
assign g[57049] = b[14] & g[24282];
assign g[40667] = a[14] & g[24283];
assign g[57050] = b[14] & g[24283];
assign g[40668] = a[14] & g[24284];
assign g[57051] = b[14] & g[24284];
assign g[40669] = a[14] & g[24285];
assign g[57052] = b[14] & g[24285];
assign g[40670] = a[14] & g[24286];
assign g[57053] = b[14] & g[24286];
assign g[40671] = a[14] & g[24287];
assign g[57054] = b[14] & g[24287];
assign g[40672] = a[14] & g[24288];
assign g[57055] = b[14] & g[24288];
assign g[40673] = a[14] & g[24289];
assign g[57056] = b[14] & g[24289];
assign g[40674] = a[14] & g[24290];
assign g[57057] = b[14] & g[24290];
assign g[40675] = a[14] & g[24291];
assign g[57058] = b[14] & g[24291];
assign g[40676] = a[14] & g[24292];
assign g[57059] = b[14] & g[24292];
assign g[40677] = a[14] & g[24293];
assign g[57060] = b[14] & g[24293];
assign g[40678] = a[14] & g[24294];
assign g[57061] = b[14] & g[24294];
assign g[40679] = a[14] & g[24295];
assign g[57062] = b[14] & g[24295];
assign g[40680] = a[14] & g[24296];
assign g[57063] = b[14] & g[24296];
assign g[40681] = a[14] & g[24297];
assign g[57064] = b[14] & g[24297];
assign g[40682] = a[14] & g[24298];
assign g[57065] = b[14] & g[24298];
assign g[40683] = a[14] & g[24299];
assign g[57066] = b[14] & g[24299];
assign g[40684] = a[14] & g[24300];
assign g[57067] = b[14] & g[24300];
assign g[40685] = a[14] & g[24301];
assign g[57068] = b[14] & g[24301];
assign g[40686] = a[14] & g[24302];
assign g[57069] = b[14] & g[24302];
assign g[40687] = a[14] & g[24303];
assign g[57070] = b[14] & g[24303];
assign g[40688] = a[14] & g[24304];
assign g[57071] = b[14] & g[24304];
assign g[40689] = a[14] & g[24305];
assign g[57072] = b[14] & g[24305];
assign g[40690] = a[14] & g[24306];
assign g[57073] = b[14] & g[24306];
assign g[40691] = a[14] & g[24307];
assign g[57074] = b[14] & g[24307];
assign g[40692] = a[14] & g[24308];
assign g[57075] = b[14] & g[24308];
assign g[40693] = a[14] & g[24309];
assign g[57076] = b[14] & g[24309];
assign g[40694] = a[14] & g[24310];
assign g[57077] = b[14] & g[24310];
assign g[40695] = a[14] & g[24311];
assign g[57078] = b[14] & g[24311];
assign g[40696] = a[14] & g[24312];
assign g[57079] = b[14] & g[24312];
assign g[40697] = a[14] & g[24313];
assign g[57080] = b[14] & g[24313];
assign g[40698] = a[14] & g[24314];
assign g[57081] = b[14] & g[24314];
assign g[40699] = a[14] & g[24315];
assign g[57082] = b[14] & g[24315];
assign g[40700] = a[14] & g[24316];
assign g[57083] = b[14] & g[24316];
assign g[40701] = a[14] & g[24317];
assign g[57084] = b[14] & g[24317];
assign g[40702] = a[14] & g[24318];
assign g[57085] = b[14] & g[24318];
assign g[40703] = a[14] & g[24319];
assign g[57086] = b[14] & g[24319];
assign g[40704] = a[14] & g[24320];
assign g[57087] = b[14] & g[24320];
assign g[40705] = a[14] & g[24321];
assign g[57088] = b[14] & g[24321];
assign g[40706] = a[14] & g[24322];
assign g[57089] = b[14] & g[24322];
assign g[40707] = a[14] & g[24323];
assign g[57090] = b[14] & g[24323];
assign g[40708] = a[14] & g[24324];
assign g[57091] = b[14] & g[24324];
assign g[40709] = a[14] & g[24325];
assign g[57092] = b[14] & g[24325];
assign g[40710] = a[14] & g[24326];
assign g[57093] = b[14] & g[24326];
assign g[40711] = a[14] & g[24327];
assign g[57094] = b[14] & g[24327];
assign g[40712] = a[14] & g[24328];
assign g[57095] = b[14] & g[24328];
assign g[40713] = a[14] & g[24329];
assign g[57096] = b[14] & g[24329];
assign g[40714] = a[14] & g[24330];
assign g[57097] = b[14] & g[24330];
assign g[40715] = a[14] & g[24331];
assign g[57098] = b[14] & g[24331];
assign g[40716] = a[14] & g[24332];
assign g[57099] = b[14] & g[24332];
assign g[40717] = a[14] & g[24333];
assign g[57100] = b[14] & g[24333];
assign g[40718] = a[14] & g[24334];
assign g[57101] = b[14] & g[24334];
assign g[40719] = a[14] & g[24335];
assign g[57102] = b[14] & g[24335];
assign g[40720] = a[14] & g[24336];
assign g[57103] = b[14] & g[24336];
assign g[40721] = a[14] & g[24337];
assign g[57104] = b[14] & g[24337];
assign g[40722] = a[14] & g[24338];
assign g[57105] = b[14] & g[24338];
assign g[40723] = a[14] & g[24339];
assign g[57106] = b[14] & g[24339];
assign g[40724] = a[14] & g[24340];
assign g[57107] = b[14] & g[24340];
assign g[40725] = a[14] & g[24341];
assign g[57108] = b[14] & g[24341];
assign g[40726] = a[14] & g[24342];
assign g[57109] = b[14] & g[24342];
assign g[40727] = a[14] & g[24343];
assign g[57110] = b[14] & g[24343];
assign g[40728] = a[14] & g[24344];
assign g[57111] = b[14] & g[24344];
assign g[40729] = a[14] & g[24345];
assign g[57112] = b[14] & g[24345];
assign g[40730] = a[14] & g[24346];
assign g[57113] = b[14] & g[24346];
assign g[40731] = a[14] & g[24347];
assign g[57114] = b[14] & g[24347];
assign g[40732] = a[14] & g[24348];
assign g[57115] = b[14] & g[24348];
assign g[40733] = a[14] & g[24349];
assign g[57116] = b[14] & g[24349];
assign g[40734] = a[14] & g[24350];
assign g[57117] = b[14] & g[24350];
assign g[40735] = a[14] & g[24351];
assign g[57118] = b[14] & g[24351];
assign g[40736] = a[14] & g[24352];
assign g[57119] = b[14] & g[24352];
assign g[40737] = a[14] & g[24353];
assign g[57120] = b[14] & g[24353];
assign g[40738] = a[14] & g[24354];
assign g[57121] = b[14] & g[24354];
assign g[40739] = a[14] & g[24355];
assign g[57122] = b[14] & g[24355];
assign g[40740] = a[14] & g[24356];
assign g[57123] = b[14] & g[24356];
assign g[40741] = a[14] & g[24357];
assign g[57124] = b[14] & g[24357];
assign g[40742] = a[14] & g[24358];
assign g[57125] = b[14] & g[24358];
assign g[40743] = a[14] & g[24359];
assign g[57126] = b[14] & g[24359];
assign g[40744] = a[14] & g[24360];
assign g[57127] = b[14] & g[24360];
assign g[40745] = a[14] & g[24361];
assign g[57128] = b[14] & g[24361];
assign g[40746] = a[14] & g[24362];
assign g[57129] = b[14] & g[24362];
assign g[40747] = a[14] & g[24363];
assign g[57130] = b[14] & g[24363];
assign g[40748] = a[14] & g[24364];
assign g[57131] = b[14] & g[24364];
assign g[40749] = a[14] & g[24365];
assign g[57132] = b[14] & g[24365];
assign g[40750] = a[14] & g[24366];
assign g[57133] = b[14] & g[24366];
assign g[40751] = a[14] & g[24367];
assign g[57134] = b[14] & g[24367];
assign g[40752] = a[14] & g[24368];
assign g[57135] = b[14] & g[24368];
assign g[40753] = a[14] & g[24369];
assign g[57136] = b[14] & g[24369];
assign g[40754] = a[14] & g[24370];
assign g[57137] = b[14] & g[24370];
assign g[40755] = a[14] & g[24371];
assign g[57138] = b[14] & g[24371];
assign g[40756] = a[14] & g[24372];
assign g[57139] = b[14] & g[24372];
assign g[40757] = a[14] & g[24373];
assign g[57140] = b[14] & g[24373];
assign g[40758] = a[14] & g[24374];
assign g[57141] = b[14] & g[24374];
assign g[40759] = a[14] & g[24375];
assign g[57142] = b[14] & g[24375];
assign g[40760] = a[14] & g[24376];
assign g[57143] = b[14] & g[24376];
assign g[40761] = a[14] & g[24377];
assign g[57144] = b[14] & g[24377];
assign g[40762] = a[14] & g[24378];
assign g[57145] = b[14] & g[24378];
assign g[40763] = a[14] & g[24379];
assign g[57146] = b[14] & g[24379];
assign g[40764] = a[14] & g[24380];
assign g[57147] = b[14] & g[24380];
assign g[40765] = a[14] & g[24381];
assign g[57148] = b[14] & g[24381];
assign g[40766] = a[14] & g[24382];
assign g[57149] = b[14] & g[24382];
assign g[40767] = a[14] & g[24383];
assign g[57150] = b[14] & g[24383];
assign g[40768] = a[14] & g[24384];
assign g[57151] = b[14] & g[24384];
assign g[40769] = a[14] & g[24385];
assign g[57152] = b[14] & g[24385];
assign g[40770] = a[14] & g[24386];
assign g[57153] = b[14] & g[24386];
assign g[40771] = a[14] & g[24387];
assign g[57154] = b[14] & g[24387];
assign g[40772] = a[14] & g[24388];
assign g[57155] = b[14] & g[24388];
assign g[40773] = a[14] & g[24389];
assign g[57156] = b[14] & g[24389];
assign g[40774] = a[14] & g[24390];
assign g[57157] = b[14] & g[24390];
assign g[40775] = a[14] & g[24391];
assign g[57158] = b[14] & g[24391];
assign g[40776] = a[14] & g[24392];
assign g[57159] = b[14] & g[24392];
assign g[40777] = a[14] & g[24393];
assign g[57160] = b[14] & g[24393];
assign g[40778] = a[14] & g[24394];
assign g[57161] = b[14] & g[24394];
assign g[40779] = a[14] & g[24395];
assign g[57162] = b[14] & g[24395];
assign g[40780] = a[14] & g[24396];
assign g[57163] = b[14] & g[24396];
assign g[40781] = a[14] & g[24397];
assign g[57164] = b[14] & g[24397];
assign g[40782] = a[14] & g[24398];
assign g[57165] = b[14] & g[24398];
assign g[40783] = a[14] & g[24399];
assign g[57166] = b[14] & g[24399];
assign g[40784] = a[14] & g[24400];
assign g[57167] = b[14] & g[24400];
assign g[40785] = a[14] & g[24401];
assign g[57168] = b[14] & g[24401];
assign g[40786] = a[14] & g[24402];
assign g[57169] = b[14] & g[24402];
assign g[40787] = a[14] & g[24403];
assign g[57170] = b[14] & g[24403];
assign g[40788] = a[14] & g[24404];
assign g[57171] = b[14] & g[24404];
assign g[40789] = a[14] & g[24405];
assign g[57172] = b[14] & g[24405];
assign g[40790] = a[14] & g[24406];
assign g[57173] = b[14] & g[24406];
assign g[40791] = a[14] & g[24407];
assign g[57174] = b[14] & g[24407];
assign g[40792] = a[14] & g[24408];
assign g[57175] = b[14] & g[24408];
assign g[40793] = a[14] & g[24409];
assign g[57176] = b[14] & g[24409];
assign g[40794] = a[14] & g[24410];
assign g[57177] = b[14] & g[24410];
assign g[40795] = a[14] & g[24411];
assign g[57178] = b[14] & g[24411];
assign g[40796] = a[14] & g[24412];
assign g[57179] = b[14] & g[24412];
assign g[40797] = a[14] & g[24413];
assign g[57180] = b[14] & g[24413];
assign g[40798] = a[14] & g[24414];
assign g[57181] = b[14] & g[24414];
assign g[40799] = a[14] & g[24415];
assign g[57182] = b[14] & g[24415];
assign g[40800] = a[14] & g[24416];
assign g[57183] = b[14] & g[24416];
assign g[40801] = a[14] & g[24417];
assign g[57184] = b[14] & g[24417];
assign g[40802] = a[14] & g[24418];
assign g[57185] = b[14] & g[24418];
assign g[40803] = a[14] & g[24419];
assign g[57186] = b[14] & g[24419];
assign g[40804] = a[14] & g[24420];
assign g[57187] = b[14] & g[24420];
assign g[40805] = a[14] & g[24421];
assign g[57188] = b[14] & g[24421];
assign g[40806] = a[14] & g[24422];
assign g[57189] = b[14] & g[24422];
assign g[40807] = a[14] & g[24423];
assign g[57190] = b[14] & g[24423];
assign g[40808] = a[14] & g[24424];
assign g[57191] = b[14] & g[24424];
assign g[40809] = a[14] & g[24425];
assign g[57192] = b[14] & g[24425];
assign g[40810] = a[14] & g[24426];
assign g[57193] = b[14] & g[24426];
assign g[40811] = a[14] & g[24427];
assign g[57194] = b[14] & g[24427];
assign g[40812] = a[14] & g[24428];
assign g[57195] = b[14] & g[24428];
assign g[40813] = a[14] & g[24429];
assign g[57196] = b[14] & g[24429];
assign g[40814] = a[14] & g[24430];
assign g[57197] = b[14] & g[24430];
assign g[40815] = a[14] & g[24431];
assign g[57198] = b[14] & g[24431];
assign g[40816] = a[14] & g[24432];
assign g[57199] = b[14] & g[24432];
assign g[40817] = a[14] & g[24433];
assign g[57200] = b[14] & g[24433];
assign g[40818] = a[14] & g[24434];
assign g[57201] = b[14] & g[24434];
assign g[40819] = a[14] & g[24435];
assign g[57202] = b[14] & g[24435];
assign g[40820] = a[14] & g[24436];
assign g[57203] = b[14] & g[24436];
assign g[40821] = a[14] & g[24437];
assign g[57204] = b[14] & g[24437];
assign g[40822] = a[14] & g[24438];
assign g[57205] = b[14] & g[24438];
assign g[40823] = a[14] & g[24439];
assign g[57206] = b[14] & g[24439];
assign g[40824] = a[14] & g[24440];
assign g[57207] = b[14] & g[24440];
assign g[40825] = a[14] & g[24441];
assign g[57208] = b[14] & g[24441];
assign g[40826] = a[14] & g[24442];
assign g[57209] = b[14] & g[24442];
assign g[40827] = a[14] & g[24443];
assign g[57210] = b[14] & g[24443];
assign g[40828] = a[14] & g[24444];
assign g[57211] = b[14] & g[24444];
assign g[40829] = a[14] & g[24445];
assign g[57212] = b[14] & g[24445];
assign g[40830] = a[14] & g[24446];
assign g[57213] = b[14] & g[24446];
assign g[40831] = a[14] & g[24447];
assign g[57214] = b[14] & g[24447];
assign g[40832] = a[14] & g[24448];
assign g[57215] = b[14] & g[24448];
assign g[40833] = a[14] & g[24449];
assign g[57216] = b[14] & g[24449];
assign g[40834] = a[14] & g[24450];
assign g[57217] = b[14] & g[24450];
assign g[40835] = a[14] & g[24451];
assign g[57218] = b[14] & g[24451];
assign g[40836] = a[14] & g[24452];
assign g[57219] = b[14] & g[24452];
assign g[40837] = a[14] & g[24453];
assign g[57220] = b[14] & g[24453];
assign g[40838] = a[14] & g[24454];
assign g[57221] = b[14] & g[24454];
assign g[40839] = a[14] & g[24455];
assign g[57222] = b[14] & g[24455];
assign g[40840] = a[14] & g[24456];
assign g[57223] = b[14] & g[24456];
assign g[40841] = a[14] & g[24457];
assign g[57224] = b[14] & g[24457];
assign g[40842] = a[14] & g[24458];
assign g[57225] = b[14] & g[24458];
assign g[40843] = a[14] & g[24459];
assign g[57226] = b[14] & g[24459];
assign g[40844] = a[14] & g[24460];
assign g[57227] = b[14] & g[24460];
assign g[40845] = a[14] & g[24461];
assign g[57228] = b[14] & g[24461];
assign g[40846] = a[14] & g[24462];
assign g[57229] = b[14] & g[24462];
assign g[40847] = a[14] & g[24463];
assign g[57230] = b[14] & g[24463];
assign g[40848] = a[14] & g[24464];
assign g[57231] = b[14] & g[24464];
assign g[40849] = a[14] & g[24465];
assign g[57232] = b[14] & g[24465];
assign g[40850] = a[14] & g[24466];
assign g[57233] = b[14] & g[24466];
assign g[40851] = a[14] & g[24467];
assign g[57234] = b[14] & g[24467];
assign g[40852] = a[14] & g[24468];
assign g[57235] = b[14] & g[24468];
assign g[40853] = a[14] & g[24469];
assign g[57236] = b[14] & g[24469];
assign g[40854] = a[14] & g[24470];
assign g[57237] = b[14] & g[24470];
assign g[40855] = a[14] & g[24471];
assign g[57238] = b[14] & g[24471];
assign g[40856] = a[14] & g[24472];
assign g[57239] = b[14] & g[24472];
assign g[40857] = a[14] & g[24473];
assign g[57240] = b[14] & g[24473];
assign g[40858] = a[14] & g[24474];
assign g[57241] = b[14] & g[24474];
assign g[40859] = a[14] & g[24475];
assign g[57242] = b[14] & g[24475];
assign g[40860] = a[14] & g[24476];
assign g[57243] = b[14] & g[24476];
assign g[40861] = a[14] & g[24477];
assign g[57244] = b[14] & g[24477];
assign g[40862] = a[14] & g[24478];
assign g[57245] = b[14] & g[24478];
assign g[40863] = a[14] & g[24479];
assign g[57246] = b[14] & g[24479];
assign g[40864] = a[14] & g[24480];
assign g[57247] = b[14] & g[24480];
assign g[40865] = a[14] & g[24481];
assign g[57248] = b[14] & g[24481];
assign g[40866] = a[14] & g[24482];
assign g[57249] = b[14] & g[24482];
assign g[40867] = a[14] & g[24483];
assign g[57250] = b[14] & g[24483];
assign g[40868] = a[14] & g[24484];
assign g[57251] = b[14] & g[24484];
assign g[40869] = a[14] & g[24485];
assign g[57252] = b[14] & g[24485];
assign g[40870] = a[14] & g[24486];
assign g[57253] = b[14] & g[24486];
assign g[40871] = a[14] & g[24487];
assign g[57254] = b[14] & g[24487];
assign g[40872] = a[14] & g[24488];
assign g[57255] = b[14] & g[24488];
assign g[40873] = a[14] & g[24489];
assign g[57256] = b[14] & g[24489];
assign g[40874] = a[14] & g[24490];
assign g[57257] = b[14] & g[24490];
assign g[40875] = a[14] & g[24491];
assign g[57258] = b[14] & g[24491];
assign g[40876] = a[14] & g[24492];
assign g[57259] = b[14] & g[24492];
assign g[40877] = a[14] & g[24493];
assign g[57260] = b[14] & g[24493];
assign g[40878] = a[14] & g[24494];
assign g[57261] = b[14] & g[24494];
assign g[40879] = a[14] & g[24495];
assign g[57262] = b[14] & g[24495];
assign g[40880] = a[14] & g[24496];
assign g[57263] = b[14] & g[24496];
assign g[40881] = a[14] & g[24497];
assign g[57264] = b[14] & g[24497];
assign g[40882] = a[14] & g[24498];
assign g[57265] = b[14] & g[24498];
assign g[40883] = a[14] & g[24499];
assign g[57266] = b[14] & g[24499];
assign g[40884] = a[14] & g[24500];
assign g[57267] = b[14] & g[24500];
assign g[40885] = a[14] & g[24501];
assign g[57268] = b[14] & g[24501];
assign g[40886] = a[14] & g[24502];
assign g[57269] = b[14] & g[24502];
assign g[40887] = a[14] & g[24503];
assign g[57270] = b[14] & g[24503];
assign g[40888] = a[14] & g[24504];
assign g[57271] = b[14] & g[24504];
assign g[40889] = a[14] & g[24505];
assign g[57272] = b[14] & g[24505];
assign g[40890] = a[14] & g[24506];
assign g[57273] = b[14] & g[24506];
assign g[40891] = a[14] & g[24507];
assign g[57274] = b[14] & g[24507];
assign g[40892] = a[14] & g[24508];
assign g[57275] = b[14] & g[24508];
assign g[40893] = a[14] & g[24509];
assign g[57276] = b[14] & g[24509];
assign g[40894] = a[14] & g[24510];
assign g[57277] = b[14] & g[24510];
assign g[40895] = a[14] & g[24511];
assign g[57278] = b[14] & g[24511];
assign g[40896] = a[14] & g[24512];
assign g[57279] = b[14] & g[24512];
assign g[40897] = a[14] & g[24513];
assign g[57280] = b[14] & g[24513];
assign g[40898] = a[14] & g[24514];
assign g[57281] = b[14] & g[24514];
assign g[40899] = a[14] & g[24515];
assign g[57282] = b[14] & g[24515];
assign g[40900] = a[14] & g[24516];
assign g[57283] = b[14] & g[24516];
assign g[40901] = a[14] & g[24517];
assign g[57284] = b[14] & g[24517];
assign g[40902] = a[14] & g[24518];
assign g[57285] = b[14] & g[24518];
assign g[40903] = a[14] & g[24519];
assign g[57286] = b[14] & g[24519];
assign g[40904] = a[14] & g[24520];
assign g[57287] = b[14] & g[24520];
assign g[40905] = a[14] & g[24521];
assign g[57288] = b[14] & g[24521];
assign g[40906] = a[14] & g[24522];
assign g[57289] = b[14] & g[24522];
assign g[40907] = a[14] & g[24523];
assign g[57290] = b[14] & g[24523];
assign g[40908] = a[14] & g[24524];
assign g[57291] = b[14] & g[24524];
assign g[40909] = a[14] & g[24525];
assign g[57292] = b[14] & g[24525];
assign g[40910] = a[14] & g[24526];
assign g[57293] = b[14] & g[24526];
assign g[40911] = a[14] & g[24527];
assign g[57294] = b[14] & g[24527];
assign g[40912] = a[14] & g[24528];
assign g[57295] = b[14] & g[24528];
assign g[40913] = a[14] & g[24529];
assign g[57296] = b[14] & g[24529];
assign g[40914] = a[14] & g[24530];
assign g[57297] = b[14] & g[24530];
assign g[40915] = a[14] & g[24531];
assign g[57298] = b[14] & g[24531];
assign g[40916] = a[14] & g[24532];
assign g[57299] = b[14] & g[24532];
assign g[40917] = a[14] & g[24533];
assign g[57300] = b[14] & g[24533];
assign g[40918] = a[14] & g[24534];
assign g[57301] = b[14] & g[24534];
assign g[40919] = a[14] & g[24535];
assign g[57302] = b[14] & g[24535];
assign g[40920] = a[14] & g[24536];
assign g[57303] = b[14] & g[24536];
assign g[40921] = a[14] & g[24537];
assign g[57304] = b[14] & g[24537];
assign g[40922] = a[14] & g[24538];
assign g[57305] = b[14] & g[24538];
assign g[40923] = a[14] & g[24539];
assign g[57306] = b[14] & g[24539];
assign g[40924] = a[14] & g[24540];
assign g[57307] = b[14] & g[24540];
assign g[40925] = a[14] & g[24541];
assign g[57308] = b[14] & g[24541];
assign g[40926] = a[14] & g[24542];
assign g[57309] = b[14] & g[24542];
assign g[40927] = a[14] & g[24543];
assign g[57310] = b[14] & g[24543];
assign g[40928] = a[14] & g[24544];
assign g[57311] = b[14] & g[24544];
assign g[40929] = a[14] & g[24545];
assign g[57312] = b[14] & g[24545];
assign g[40930] = a[14] & g[24546];
assign g[57313] = b[14] & g[24546];
assign g[40931] = a[14] & g[24547];
assign g[57314] = b[14] & g[24547];
assign g[40932] = a[14] & g[24548];
assign g[57315] = b[14] & g[24548];
assign g[40933] = a[14] & g[24549];
assign g[57316] = b[14] & g[24549];
assign g[40934] = a[14] & g[24550];
assign g[57317] = b[14] & g[24550];
assign g[40935] = a[14] & g[24551];
assign g[57318] = b[14] & g[24551];
assign g[40936] = a[14] & g[24552];
assign g[57319] = b[14] & g[24552];
assign g[40937] = a[14] & g[24553];
assign g[57320] = b[14] & g[24553];
assign g[40938] = a[14] & g[24554];
assign g[57321] = b[14] & g[24554];
assign g[40939] = a[14] & g[24555];
assign g[57322] = b[14] & g[24555];
assign g[40940] = a[14] & g[24556];
assign g[57323] = b[14] & g[24556];
assign g[40941] = a[14] & g[24557];
assign g[57324] = b[14] & g[24557];
assign g[40942] = a[14] & g[24558];
assign g[57325] = b[14] & g[24558];
assign g[40943] = a[14] & g[24559];
assign g[57326] = b[14] & g[24559];
assign g[40944] = a[14] & g[24560];
assign g[57327] = b[14] & g[24560];
assign g[40945] = a[14] & g[24561];
assign g[57328] = b[14] & g[24561];
assign g[40946] = a[14] & g[24562];
assign g[57329] = b[14] & g[24562];
assign g[40947] = a[14] & g[24563];
assign g[57330] = b[14] & g[24563];
assign g[40948] = a[14] & g[24564];
assign g[57331] = b[14] & g[24564];
assign g[40949] = a[14] & g[24565];
assign g[57332] = b[14] & g[24565];
assign g[40950] = a[14] & g[24566];
assign g[57333] = b[14] & g[24566];
assign g[40951] = a[14] & g[24567];
assign g[57334] = b[14] & g[24567];
assign g[40952] = a[14] & g[24568];
assign g[57335] = b[14] & g[24568];
assign g[40953] = a[14] & g[24569];
assign g[57336] = b[14] & g[24569];
assign g[40954] = a[14] & g[24570];
assign g[57337] = b[14] & g[24570];
assign g[40955] = a[14] & g[24571];
assign g[57338] = b[14] & g[24571];
assign g[40956] = a[14] & g[24572];
assign g[57339] = b[14] & g[24572];
assign g[40957] = a[14] & g[24573];
assign g[57340] = b[14] & g[24573];
assign g[40958] = a[14] & g[24574];
assign g[57341] = b[14] & g[24574];
assign g[40959] = a[14] & g[24575];
assign g[57342] = b[14] & g[24575];
assign g[40960] = a[14] & g[24576];
assign g[57343] = b[14] & g[24576];
assign g[40961] = a[14] & g[24577];
assign g[57344] = b[14] & g[24577];
assign g[40962] = a[14] & g[24578];
assign g[57345] = b[14] & g[24578];
assign g[40963] = a[14] & g[24579];
assign g[57346] = b[14] & g[24579];
assign g[40964] = a[14] & g[24580];
assign g[57347] = b[14] & g[24580];
assign g[40965] = a[14] & g[24581];
assign g[57348] = b[14] & g[24581];
assign g[40966] = a[14] & g[24582];
assign g[57349] = b[14] & g[24582];
assign g[40967] = a[14] & g[24583];
assign g[57350] = b[14] & g[24583];
assign g[40968] = a[14] & g[24584];
assign g[57351] = b[14] & g[24584];
assign g[40969] = a[14] & g[24585];
assign g[57352] = b[14] & g[24585];
assign g[40970] = a[14] & g[24586];
assign g[57353] = b[14] & g[24586];
assign g[40971] = a[14] & g[24587];
assign g[57354] = b[14] & g[24587];
assign g[40972] = a[14] & g[24588];
assign g[57355] = b[14] & g[24588];
assign g[40973] = a[14] & g[24589];
assign g[57356] = b[14] & g[24589];
assign g[40974] = a[14] & g[24590];
assign g[57357] = b[14] & g[24590];
assign g[40975] = a[14] & g[24591];
assign g[57358] = b[14] & g[24591];
assign g[40976] = a[14] & g[24592];
assign g[57359] = b[14] & g[24592];
assign g[40977] = a[14] & g[24593];
assign g[57360] = b[14] & g[24593];
assign g[40978] = a[14] & g[24594];
assign g[57361] = b[14] & g[24594];
assign g[40979] = a[14] & g[24595];
assign g[57362] = b[14] & g[24595];
assign g[40980] = a[14] & g[24596];
assign g[57363] = b[14] & g[24596];
assign g[40981] = a[14] & g[24597];
assign g[57364] = b[14] & g[24597];
assign g[40982] = a[14] & g[24598];
assign g[57365] = b[14] & g[24598];
assign g[40983] = a[14] & g[24599];
assign g[57366] = b[14] & g[24599];
assign g[40984] = a[14] & g[24600];
assign g[57367] = b[14] & g[24600];
assign g[40985] = a[14] & g[24601];
assign g[57368] = b[14] & g[24601];
assign g[40986] = a[14] & g[24602];
assign g[57369] = b[14] & g[24602];
assign g[40987] = a[14] & g[24603];
assign g[57370] = b[14] & g[24603];
assign g[40988] = a[14] & g[24604];
assign g[57371] = b[14] & g[24604];
assign g[40989] = a[14] & g[24605];
assign g[57372] = b[14] & g[24605];
assign g[40990] = a[14] & g[24606];
assign g[57373] = b[14] & g[24606];
assign g[40991] = a[14] & g[24607];
assign g[57374] = b[14] & g[24607];
assign g[40992] = a[14] & g[24608];
assign g[57375] = b[14] & g[24608];
assign g[40993] = a[14] & g[24609];
assign g[57376] = b[14] & g[24609];
assign g[40994] = a[14] & g[24610];
assign g[57377] = b[14] & g[24610];
assign g[40995] = a[14] & g[24611];
assign g[57378] = b[14] & g[24611];
assign g[40996] = a[14] & g[24612];
assign g[57379] = b[14] & g[24612];
assign g[40997] = a[14] & g[24613];
assign g[57380] = b[14] & g[24613];
assign g[40998] = a[14] & g[24614];
assign g[57381] = b[14] & g[24614];
assign g[40999] = a[14] & g[24615];
assign g[57382] = b[14] & g[24615];
assign g[41000] = a[14] & g[24616];
assign g[57383] = b[14] & g[24616];
assign g[41001] = a[14] & g[24617];
assign g[57384] = b[14] & g[24617];
assign g[41002] = a[14] & g[24618];
assign g[57385] = b[14] & g[24618];
assign g[41003] = a[14] & g[24619];
assign g[57386] = b[14] & g[24619];
assign g[41004] = a[14] & g[24620];
assign g[57387] = b[14] & g[24620];
assign g[41005] = a[14] & g[24621];
assign g[57388] = b[14] & g[24621];
assign g[41006] = a[14] & g[24622];
assign g[57389] = b[14] & g[24622];
assign g[41007] = a[14] & g[24623];
assign g[57390] = b[14] & g[24623];
assign g[41008] = a[14] & g[24624];
assign g[57391] = b[14] & g[24624];
assign g[41009] = a[14] & g[24625];
assign g[57392] = b[14] & g[24625];
assign g[41010] = a[14] & g[24626];
assign g[57393] = b[14] & g[24626];
assign g[41011] = a[14] & g[24627];
assign g[57394] = b[14] & g[24627];
assign g[41012] = a[14] & g[24628];
assign g[57395] = b[14] & g[24628];
assign g[41013] = a[14] & g[24629];
assign g[57396] = b[14] & g[24629];
assign g[41014] = a[14] & g[24630];
assign g[57397] = b[14] & g[24630];
assign g[41015] = a[14] & g[24631];
assign g[57398] = b[14] & g[24631];
assign g[41016] = a[14] & g[24632];
assign g[57399] = b[14] & g[24632];
assign g[41017] = a[14] & g[24633];
assign g[57400] = b[14] & g[24633];
assign g[41018] = a[14] & g[24634];
assign g[57401] = b[14] & g[24634];
assign g[41019] = a[14] & g[24635];
assign g[57402] = b[14] & g[24635];
assign g[41020] = a[14] & g[24636];
assign g[57403] = b[14] & g[24636];
assign g[41021] = a[14] & g[24637];
assign g[57404] = b[14] & g[24637];
assign g[41022] = a[14] & g[24638];
assign g[57405] = b[14] & g[24638];
assign g[41023] = a[14] & g[24639];
assign g[57406] = b[14] & g[24639];
assign g[41024] = a[14] & g[24640];
assign g[57407] = b[14] & g[24640];
assign g[41025] = a[14] & g[24641];
assign g[57408] = b[14] & g[24641];
assign g[41026] = a[14] & g[24642];
assign g[57409] = b[14] & g[24642];
assign g[41027] = a[14] & g[24643];
assign g[57410] = b[14] & g[24643];
assign g[41028] = a[14] & g[24644];
assign g[57411] = b[14] & g[24644];
assign g[41029] = a[14] & g[24645];
assign g[57412] = b[14] & g[24645];
assign g[41030] = a[14] & g[24646];
assign g[57413] = b[14] & g[24646];
assign g[41031] = a[14] & g[24647];
assign g[57414] = b[14] & g[24647];
assign g[41032] = a[14] & g[24648];
assign g[57415] = b[14] & g[24648];
assign g[41033] = a[14] & g[24649];
assign g[57416] = b[14] & g[24649];
assign g[41034] = a[14] & g[24650];
assign g[57417] = b[14] & g[24650];
assign g[41035] = a[14] & g[24651];
assign g[57418] = b[14] & g[24651];
assign g[41036] = a[14] & g[24652];
assign g[57419] = b[14] & g[24652];
assign g[41037] = a[14] & g[24653];
assign g[57420] = b[14] & g[24653];
assign g[41038] = a[14] & g[24654];
assign g[57421] = b[14] & g[24654];
assign g[41039] = a[14] & g[24655];
assign g[57422] = b[14] & g[24655];
assign g[41040] = a[14] & g[24656];
assign g[57423] = b[14] & g[24656];
assign g[41041] = a[14] & g[24657];
assign g[57424] = b[14] & g[24657];
assign g[41042] = a[14] & g[24658];
assign g[57425] = b[14] & g[24658];
assign g[41043] = a[14] & g[24659];
assign g[57426] = b[14] & g[24659];
assign g[41044] = a[14] & g[24660];
assign g[57427] = b[14] & g[24660];
assign g[41045] = a[14] & g[24661];
assign g[57428] = b[14] & g[24661];
assign g[41046] = a[14] & g[24662];
assign g[57429] = b[14] & g[24662];
assign g[41047] = a[14] & g[24663];
assign g[57430] = b[14] & g[24663];
assign g[41048] = a[14] & g[24664];
assign g[57431] = b[14] & g[24664];
assign g[41049] = a[14] & g[24665];
assign g[57432] = b[14] & g[24665];
assign g[41050] = a[14] & g[24666];
assign g[57433] = b[14] & g[24666];
assign g[41051] = a[14] & g[24667];
assign g[57434] = b[14] & g[24667];
assign g[41052] = a[14] & g[24668];
assign g[57435] = b[14] & g[24668];
assign g[41053] = a[14] & g[24669];
assign g[57436] = b[14] & g[24669];
assign g[41054] = a[14] & g[24670];
assign g[57437] = b[14] & g[24670];
assign g[41055] = a[14] & g[24671];
assign g[57438] = b[14] & g[24671];
assign g[41056] = a[14] & g[24672];
assign g[57439] = b[14] & g[24672];
assign g[41057] = a[14] & g[24673];
assign g[57440] = b[14] & g[24673];
assign g[41058] = a[14] & g[24674];
assign g[57441] = b[14] & g[24674];
assign g[41059] = a[14] & g[24675];
assign g[57442] = b[14] & g[24675];
assign g[41060] = a[14] & g[24676];
assign g[57443] = b[14] & g[24676];
assign g[41061] = a[14] & g[24677];
assign g[57444] = b[14] & g[24677];
assign g[41062] = a[14] & g[24678];
assign g[57445] = b[14] & g[24678];
assign g[41063] = a[14] & g[24679];
assign g[57446] = b[14] & g[24679];
assign g[41064] = a[14] & g[24680];
assign g[57447] = b[14] & g[24680];
assign g[41065] = a[14] & g[24681];
assign g[57448] = b[14] & g[24681];
assign g[41066] = a[14] & g[24682];
assign g[57449] = b[14] & g[24682];
assign g[41067] = a[14] & g[24683];
assign g[57450] = b[14] & g[24683];
assign g[41068] = a[14] & g[24684];
assign g[57451] = b[14] & g[24684];
assign g[41069] = a[14] & g[24685];
assign g[57452] = b[14] & g[24685];
assign g[41070] = a[14] & g[24686];
assign g[57453] = b[14] & g[24686];
assign g[41071] = a[14] & g[24687];
assign g[57454] = b[14] & g[24687];
assign g[41072] = a[14] & g[24688];
assign g[57455] = b[14] & g[24688];
assign g[41073] = a[14] & g[24689];
assign g[57456] = b[14] & g[24689];
assign g[41074] = a[14] & g[24690];
assign g[57457] = b[14] & g[24690];
assign g[41075] = a[14] & g[24691];
assign g[57458] = b[14] & g[24691];
assign g[41076] = a[14] & g[24692];
assign g[57459] = b[14] & g[24692];
assign g[41077] = a[14] & g[24693];
assign g[57460] = b[14] & g[24693];
assign g[41078] = a[14] & g[24694];
assign g[57461] = b[14] & g[24694];
assign g[41079] = a[14] & g[24695];
assign g[57462] = b[14] & g[24695];
assign g[41080] = a[14] & g[24696];
assign g[57463] = b[14] & g[24696];
assign g[41081] = a[14] & g[24697];
assign g[57464] = b[14] & g[24697];
assign g[41082] = a[14] & g[24698];
assign g[57465] = b[14] & g[24698];
assign g[41083] = a[14] & g[24699];
assign g[57466] = b[14] & g[24699];
assign g[41084] = a[14] & g[24700];
assign g[57467] = b[14] & g[24700];
assign g[41085] = a[14] & g[24701];
assign g[57468] = b[14] & g[24701];
assign g[41086] = a[14] & g[24702];
assign g[57469] = b[14] & g[24702];
assign g[41087] = a[14] & g[24703];
assign g[57470] = b[14] & g[24703];
assign g[41088] = a[14] & g[24704];
assign g[57471] = b[14] & g[24704];
assign g[41089] = a[14] & g[24705];
assign g[57472] = b[14] & g[24705];
assign g[41090] = a[14] & g[24706];
assign g[57473] = b[14] & g[24706];
assign g[41091] = a[14] & g[24707];
assign g[57474] = b[14] & g[24707];
assign g[41092] = a[14] & g[24708];
assign g[57475] = b[14] & g[24708];
assign g[41093] = a[14] & g[24709];
assign g[57476] = b[14] & g[24709];
assign g[41094] = a[14] & g[24710];
assign g[57477] = b[14] & g[24710];
assign g[41095] = a[14] & g[24711];
assign g[57478] = b[14] & g[24711];
assign g[41096] = a[14] & g[24712];
assign g[57479] = b[14] & g[24712];
assign g[41097] = a[14] & g[24713];
assign g[57480] = b[14] & g[24713];
assign g[41098] = a[14] & g[24714];
assign g[57481] = b[14] & g[24714];
assign g[41099] = a[14] & g[24715];
assign g[57482] = b[14] & g[24715];
assign g[41100] = a[14] & g[24716];
assign g[57483] = b[14] & g[24716];
assign g[41101] = a[14] & g[24717];
assign g[57484] = b[14] & g[24717];
assign g[41102] = a[14] & g[24718];
assign g[57485] = b[14] & g[24718];
assign g[41103] = a[14] & g[24719];
assign g[57486] = b[14] & g[24719];
assign g[41104] = a[14] & g[24720];
assign g[57487] = b[14] & g[24720];
assign g[41105] = a[14] & g[24721];
assign g[57488] = b[14] & g[24721];
assign g[41106] = a[14] & g[24722];
assign g[57489] = b[14] & g[24722];
assign g[41107] = a[14] & g[24723];
assign g[57490] = b[14] & g[24723];
assign g[41108] = a[14] & g[24724];
assign g[57491] = b[14] & g[24724];
assign g[41109] = a[14] & g[24725];
assign g[57492] = b[14] & g[24725];
assign g[41110] = a[14] & g[24726];
assign g[57493] = b[14] & g[24726];
assign g[41111] = a[14] & g[24727];
assign g[57494] = b[14] & g[24727];
assign g[41112] = a[14] & g[24728];
assign g[57495] = b[14] & g[24728];
assign g[41113] = a[14] & g[24729];
assign g[57496] = b[14] & g[24729];
assign g[41114] = a[14] & g[24730];
assign g[57497] = b[14] & g[24730];
assign g[41115] = a[14] & g[24731];
assign g[57498] = b[14] & g[24731];
assign g[41116] = a[14] & g[24732];
assign g[57499] = b[14] & g[24732];
assign g[41117] = a[14] & g[24733];
assign g[57500] = b[14] & g[24733];
assign g[41118] = a[14] & g[24734];
assign g[57501] = b[14] & g[24734];
assign g[41119] = a[14] & g[24735];
assign g[57502] = b[14] & g[24735];
assign g[41120] = a[14] & g[24736];
assign g[57503] = b[14] & g[24736];
assign g[41121] = a[14] & g[24737];
assign g[57504] = b[14] & g[24737];
assign g[41122] = a[14] & g[24738];
assign g[57505] = b[14] & g[24738];
assign g[41123] = a[14] & g[24739];
assign g[57506] = b[14] & g[24739];
assign g[41124] = a[14] & g[24740];
assign g[57507] = b[14] & g[24740];
assign g[41125] = a[14] & g[24741];
assign g[57508] = b[14] & g[24741];
assign g[41126] = a[14] & g[24742];
assign g[57509] = b[14] & g[24742];
assign g[41127] = a[14] & g[24743];
assign g[57510] = b[14] & g[24743];
assign g[41128] = a[14] & g[24744];
assign g[57511] = b[14] & g[24744];
assign g[41129] = a[14] & g[24745];
assign g[57512] = b[14] & g[24745];
assign g[41130] = a[14] & g[24746];
assign g[57513] = b[14] & g[24746];
assign g[41131] = a[14] & g[24747];
assign g[57514] = b[14] & g[24747];
assign g[41132] = a[14] & g[24748];
assign g[57515] = b[14] & g[24748];
assign g[41133] = a[14] & g[24749];
assign g[57516] = b[14] & g[24749];
assign g[41134] = a[14] & g[24750];
assign g[57517] = b[14] & g[24750];
assign g[41135] = a[14] & g[24751];
assign g[57518] = b[14] & g[24751];
assign g[41136] = a[14] & g[24752];
assign g[57519] = b[14] & g[24752];
assign g[41137] = a[14] & g[24753];
assign g[57520] = b[14] & g[24753];
assign g[41138] = a[14] & g[24754];
assign g[57521] = b[14] & g[24754];
assign g[41139] = a[14] & g[24755];
assign g[57522] = b[14] & g[24755];
assign g[41140] = a[14] & g[24756];
assign g[57523] = b[14] & g[24756];
assign g[41141] = a[14] & g[24757];
assign g[57524] = b[14] & g[24757];
assign g[41142] = a[14] & g[24758];
assign g[57525] = b[14] & g[24758];
assign g[41143] = a[14] & g[24759];
assign g[57526] = b[14] & g[24759];
assign g[41144] = a[14] & g[24760];
assign g[57527] = b[14] & g[24760];
assign g[41145] = a[14] & g[24761];
assign g[57528] = b[14] & g[24761];
assign g[41146] = a[14] & g[24762];
assign g[57529] = b[14] & g[24762];
assign g[41147] = a[14] & g[24763];
assign g[57530] = b[14] & g[24763];
assign g[41148] = a[14] & g[24764];
assign g[57531] = b[14] & g[24764];
assign g[41149] = a[14] & g[24765];
assign g[57532] = b[14] & g[24765];
assign g[41150] = a[14] & g[24766];
assign g[57533] = b[14] & g[24766];
assign g[41151] = a[14] & g[24767];
assign g[57534] = b[14] & g[24767];
assign g[41152] = a[14] & g[24768];
assign g[57535] = b[14] & g[24768];
assign g[41153] = a[14] & g[24769];
assign g[57536] = b[14] & g[24769];
assign g[41154] = a[14] & g[24770];
assign g[57537] = b[14] & g[24770];
assign g[41155] = a[14] & g[24771];
assign g[57538] = b[14] & g[24771];
assign g[41156] = a[14] & g[24772];
assign g[57539] = b[14] & g[24772];
assign g[41157] = a[14] & g[24773];
assign g[57540] = b[14] & g[24773];
assign g[41158] = a[14] & g[24774];
assign g[57541] = b[14] & g[24774];
assign g[41159] = a[14] & g[24775];
assign g[57542] = b[14] & g[24775];
assign g[41160] = a[14] & g[24776];
assign g[57543] = b[14] & g[24776];
assign g[41161] = a[14] & g[24777];
assign g[57544] = b[14] & g[24777];
assign g[41162] = a[14] & g[24778];
assign g[57545] = b[14] & g[24778];
assign g[41163] = a[14] & g[24779];
assign g[57546] = b[14] & g[24779];
assign g[41164] = a[14] & g[24780];
assign g[57547] = b[14] & g[24780];
assign g[41165] = a[14] & g[24781];
assign g[57548] = b[14] & g[24781];
assign g[41166] = a[14] & g[24782];
assign g[57549] = b[14] & g[24782];
assign g[41167] = a[14] & g[24783];
assign g[57550] = b[14] & g[24783];
assign g[41168] = a[14] & g[24784];
assign g[57551] = b[14] & g[24784];
assign g[41169] = a[14] & g[24785];
assign g[57552] = b[14] & g[24785];
assign g[41170] = a[14] & g[24786];
assign g[57553] = b[14] & g[24786];
assign g[41171] = a[14] & g[24787];
assign g[57554] = b[14] & g[24787];
assign g[41172] = a[14] & g[24788];
assign g[57555] = b[14] & g[24788];
assign g[41173] = a[14] & g[24789];
assign g[57556] = b[14] & g[24789];
assign g[41174] = a[14] & g[24790];
assign g[57557] = b[14] & g[24790];
assign g[41175] = a[14] & g[24791];
assign g[57558] = b[14] & g[24791];
assign g[41176] = a[14] & g[24792];
assign g[57559] = b[14] & g[24792];
assign g[41177] = a[14] & g[24793];
assign g[57560] = b[14] & g[24793];
assign g[41178] = a[14] & g[24794];
assign g[57561] = b[14] & g[24794];
assign g[41179] = a[14] & g[24795];
assign g[57562] = b[14] & g[24795];
assign g[41180] = a[14] & g[24796];
assign g[57563] = b[14] & g[24796];
assign g[41181] = a[14] & g[24797];
assign g[57564] = b[14] & g[24797];
assign g[41182] = a[14] & g[24798];
assign g[57565] = b[14] & g[24798];
assign g[41183] = a[14] & g[24799];
assign g[57566] = b[14] & g[24799];
assign g[41184] = a[14] & g[24800];
assign g[57567] = b[14] & g[24800];
assign g[41185] = a[14] & g[24801];
assign g[57568] = b[14] & g[24801];
assign g[41186] = a[14] & g[24802];
assign g[57569] = b[14] & g[24802];
assign g[41187] = a[14] & g[24803];
assign g[57570] = b[14] & g[24803];
assign g[41188] = a[14] & g[24804];
assign g[57571] = b[14] & g[24804];
assign g[41189] = a[14] & g[24805];
assign g[57572] = b[14] & g[24805];
assign g[41190] = a[14] & g[24806];
assign g[57573] = b[14] & g[24806];
assign g[41191] = a[14] & g[24807];
assign g[57574] = b[14] & g[24807];
assign g[41192] = a[14] & g[24808];
assign g[57575] = b[14] & g[24808];
assign g[41193] = a[14] & g[24809];
assign g[57576] = b[14] & g[24809];
assign g[41194] = a[14] & g[24810];
assign g[57577] = b[14] & g[24810];
assign g[41195] = a[14] & g[24811];
assign g[57578] = b[14] & g[24811];
assign g[41196] = a[14] & g[24812];
assign g[57579] = b[14] & g[24812];
assign g[41197] = a[14] & g[24813];
assign g[57580] = b[14] & g[24813];
assign g[41198] = a[14] & g[24814];
assign g[57581] = b[14] & g[24814];
assign g[41199] = a[14] & g[24815];
assign g[57582] = b[14] & g[24815];
assign g[41200] = a[14] & g[24816];
assign g[57583] = b[14] & g[24816];
assign g[41201] = a[14] & g[24817];
assign g[57584] = b[14] & g[24817];
assign g[41202] = a[14] & g[24818];
assign g[57585] = b[14] & g[24818];
assign g[41203] = a[14] & g[24819];
assign g[57586] = b[14] & g[24819];
assign g[41204] = a[14] & g[24820];
assign g[57587] = b[14] & g[24820];
assign g[41205] = a[14] & g[24821];
assign g[57588] = b[14] & g[24821];
assign g[41206] = a[14] & g[24822];
assign g[57589] = b[14] & g[24822];
assign g[41207] = a[14] & g[24823];
assign g[57590] = b[14] & g[24823];
assign g[41208] = a[14] & g[24824];
assign g[57591] = b[14] & g[24824];
assign g[41209] = a[14] & g[24825];
assign g[57592] = b[14] & g[24825];
assign g[41210] = a[14] & g[24826];
assign g[57593] = b[14] & g[24826];
assign g[41211] = a[14] & g[24827];
assign g[57594] = b[14] & g[24827];
assign g[41212] = a[14] & g[24828];
assign g[57595] = b[14] & g[24828];
assign g[41213] = a[14] & g[24829];
assign g[57596] = b[14] & g[24829];
assign g[41214] = a[14] & g[24830];
assign g[57597] = b[14] & g[24830];
assign g[41215] = a[14] & g[24831];
assign g[57598] = b[14] & g[24831];
assign g[41216] = a[14] & g[24832];
assign g[57599] = b[14] & g[24832];
assign g[41217] = a[14] & g[24833];
assign g[57600] = b[14] & g[24833];
assign g[41218] = a[14] & g[24834];
assign g[57601] = b[14] & g[24834];
assign g[41219] = a[14] & g[24835];
assign g[57602] = b[14] & g[24835];
assign g[41220] = a[14] & g[24836];
assign g[57603] = b[14] & g[24836];
assign g[41221] = a[14] & g[24837];
assign g[57604] = b[14] & g[24837];
assign g[41222] = a[14] & g[24838];
assign g[57605] = b[14] & g[24838];
assign g[41223] = a[14] & g[24839];
assign g[57606] = b[14] & g[24839];
assign g[41224] = a[14] & g[24840];
assign g[57607] = b[14] & g[24840];
assign g[41225] = a[14] & g[24841];
assign g[57608] = b[14] & g[24841];
assign g[41226] = a[14] & g[24842];
assign g[57609] = b[14] & g[24842];
assign g[41227] = a[14] & g[24843];
assign g[57610] = b[14] & g[24843];
assign g[41228] = a[14] & g[24844];
assign g[57611] = b[14] & g[24844];
assign g[41229] = a[14] & g[24845];
assign g[57612] = b[14] & g[24845];
assign g[41230] = a[14] & g[24846];
assign g[57613] = b[14] & g[24846];
assign g[41231] = a[14] & g[24847];
assign g[57614] = b[14] & g[24847];
assign g[41232] = a[14] & g[24848];
assign g[57615] = b[14] & g[24848];
assign g[41233] = a[14] & g[24849];
assign g[57616] = b[14] & g[24849];
assign g[41234] = a[14] & g[24850];
assign g[57617] = b[14] & g[24850];
assign g[41235] = a[14] & g[24851];
assign g[57618] = b[14] & g[24851];
assign g[41236] = a[14] & g[24852];
assign g[57619] = b[14] & g[24852];
assign g[41237] = a[14] & g[24853];
assign g[57620] = b[14] & g[24853];
assign g[41238] = a[14] & g[24854];
assign g[57621] = b[14] & g[24854];
assign g[41239] = a[14] & g[24855];
assign g[57622] = b[14] & g[24855];
assign g[41240] = a[14] & g[24856];
assign g[57623] = b[14] & g[24856];
assign g[41241] = a[14] & g[24857];
assign g[57624] = b[14] & g[24857];
assign g[41242] = a[14] & g[24858];
assign g[57625] = b[14] & g[24858];
assign g[41243] = a[14] & g[24859];
assign g[57626] = b[14] & g[24859];
assign g[41244] = a[14] & g[24860];
assign g[57627] = b[14] & g[24860];
assign g[41245] = a[14] & g[24861];
assign g[57628] = b[14] & g[24861];
assign g[41246] = a[14] & g[24862];
assign g[57629] = b[14] & g[24862];
assign g[41247] = a[14] & g[24863];
assign g[57630] = b[14] & g[24863];
assign g[41248] = a[14] & g[24864];
assign g[57631] = b[14] & g[24864];
assign g[41249] = a[14] & g[24865];
assign g[57632] = b[14] & g[24865];
assign g[41250] = a[14] & g[24866];
assign g[57633] = b[14] & g[24866];
assign g[41251] = a[14] & g[24867];
assign g[57634] = b[14] & g[24867];
assign g[41252] = a[14] & g[24868];
assign g[57635] = b[14] & g[24868];
assign g[41253] = a[14] & g[24869];
assign g[57636] = b[14] & g[24869];
assign g[41254] = a[14] & g[24870];
assign g[57637] = b[14] & g[24870];
assign g[41255] = a[14] & g[24871];
assign g[57638] = b[14] & g[24871];
assign g[41256] = a[14] & g[24872];
assign g[57639] = b[14] & g[24872];
assign g[41257] = a[14] & g[24873];
assign g[57640] = b[14] & g[24873];
assign g[41258] = a[14] & g[24874];
assign g[57641] = b[14] & g[24874];
assign g[41259] = a[14] & g[24875];
assign g[57642] = b[14] & g[24875];
assign g[41260] = a[14] & g[24876];
assign g[57643] = b[14] & g[24876];
assign g[41261] = a[14] & g[24877];
assign g[57644] = b[14] & g[24877];
assign g[41262] = a[14] & g[24878];
assign g[57645] = b[14] & g[24878];
assign g[41263] = a[14] & g[24879];
assign g[57646] = b[14] & g[24879];
assign g[41264] = a[14] & g[24880];
assign g[57647] = b[14] & g[24880];
assign g[41265] = a[14] & g[24881];
assign g[57648] = b[14] & g[24881];
assign g[41266] = a[14] & g[24882];
assign g[57649] = b[14] & g[24882];
assign g[41267] = a[14] & g[24883];
assign g[57650] = b[14] & g[24883];
assign g[41268] = a[14] & g[24884];
assign g[57651] = b[14] & g[24884];
assign g[41269] = a[14] & g[24885];
assign g[57652] = b[14] & g[24885];
assign g[41270] = a[14] & g[24886];
assign g[57653] = b[14] & g[24886];
assign g[41271] = a[14] & g[24887];
assign g[57654] = b[14] & g[24887];
assign g[41272] = a[14] & g[24888];
assign g[57655] = b[14] & g[24888];
assign g[41273] = a[14] & g[24889];
assign g[57656] = b[14] & g[24889];
assign g[41274] = a[14] & g[24890];
assign g[57657] = b[14] & g[24890];
assign g[41275] = a[14] & g[24891];
assign g[57658] = b[14] & g[24891];
assign g[41276] = a[14] & g[24892];
assign g[57659] = b[14] & g[24892];
assign g[41277] = a[14] & g[24893];
assign g[57660] = b[14] & g[24893];
assign g[41278] = a[14] & g[24894];
assign g[57661] = b[14] & g[24894];
assign g[41279] = a[14] & g[24895];
assign g[57662] = b[14] & g[24895];
assign g[41280] = a[14] & g[24896];
assign g[57663] = b[14] & g[24896];
assign g[41281] = a[14] & g[24897];
assign g[57664] = b[14] & g[24897];
assign g[41282] = a[14] & g[24898];
assign g[57665] = b[14] & g[24898];
assign g[41283] = a[14] & g[24899];
assign g[57666] = b[14] & g[24899];
assign g[41284] = a[14] & g[24900];
assign g[57667] = b[14] & g[24900];
assign g[41285] = a[14] & g[24901];
assign g[57668] = b[14] & g[24901];
assign g[41286] = a[14] & g[24902];
assign g[57669] = b[14] & g[24902];
assign g[41287] = a[14] & g[24903];
assign g[57670] = b[14] & g[24903];
assign g[41288] = a[14] & g[24904];
assign g[57671] = b[14] & g[24904];
assign g[41289] = a[14] & g[24905];
assign g[57672] = b[14] & g[24905];
assign g[41290] = a[14] & g[24906];
assign g[57673] = b[14] & g[24906];
assign g[41291] = a[14] & g[24907];
assign g[57674] = b[14] & g[24907];
assign g[41292] = a[14] & g[24908];
assign g[57675] = b[14] & g[24908];
assign g[41293] = a[14] & g[24909];
assign g[57676] = b[14] & g[24909];
assign g[41294] = a[14] & g[24910];
assign g[57677] = b[14] & g[24910];
assign g[41295] = a[14] & g[24911];
assign g[57678] = b[14] & g[24911];
assign g[41296] = a[14] & g[24912];
assign g[57679] = b[14] & g[24912];
assign g[41297] = a[14] & g[24913];
assign g[57680] = b[14] & g[24913];
assign g[41298] = a[14] & g[24914];
assign g[57681] = b[14] & g[24914];
assign g[41299] = a[14] & g[24915];
assign g[57682] = b[14] & g[24915];
assign g[41300] = a[14] & g[24916];
assign g[57683] = b[14] & g[24916];
assign g[41301] = a[14] & g[24917];
assign g[57684] = b[14] & g[24917];
assign g[41302] = a[14] & g[24918];
assign g[57685] = b[14] & g[24918];
assign g[41303] = a[14] & g[24919];
assign g[57686] = b[14] & g[24919];
assign g[41304] = a[14] & g[24920];
assign g[57687] = b[14] & g[24920];
assign g[41305] = a[14] & g[24921];
assign g[57688] = b[14] & g[24921];
assign g[41306] = a[14] & g[24922];
assign g[57689] = b[14] & g[24922];
assign g[41307] = a[14] & g[24923];
assign g[57690] = b[14] & g[24923];
assign g[41308] = a[14] & g[24924];
assign g[57691] = b[14] & g[24924];
assign g[41309] = a[14] & g[24925];
assign g[57692] = b[14] & g[24925];
assign g[41310] = a[14] & g[24926];
assign g[57693] = b[14] & g[24926];
assign g[41311] = a[14] & g[24927];
assign g[57694] = b[14] & g[24927];
assign g[41312] = a[14] & g[24928];
assign g[57695] = b[14] & g[24928];
assign g[41313] = a[14] & g[24929];
assign g[57696] = b[14] & g[24929];
assign g[41314] = a[14] & g[24930];
assign g[57697] = b[14] & g[24930];
assign g[41315] = a[14] & g[24931];
assign g[57698] = b[14] & g[24931];
assign g[41316] = a[14] & g[24932];
assign g[57699] = b[14] & g[24932];
assign g[41317] = a[14] & g[24933];
assign g[57700] = b[14] & g[24933];
assign g[41318] = a[14] & g[24934];
assign g[57701] = b[14] & g[24934];
assign g[41319] = a[14] & g[24935];
assign g[57702] = b[14] & g[24935];
assign g[41320] = a[14] & g[24936];
assign g[57703] = b[14] & g[24936];
assign g[41321] = a[14] & g[24937];
assign g[57704] = b[14] & g[24937];
assign g[41322] = a[14] & g[24938];
assign g[57705] = b[14] & g[24938];
assign g[41323] = a[14] & g[24939];
assign g[57706] = b[14] & g[24939];
assign g[41324] = a[14] & g[24940];
assign g[57707] = b[14] & g[24940];
assign g[41325] = a[14] & g[24941];
assign g[57708] = b[14] & g[24941];
assign g[41326] = a[14] & g[24942];
assign g[57709] = b[14] & g[24942];
assign g[41327] = a[14] & g[24943];
assign g[57710] = b[14] & g[24943];
assign g[41328] = a[14] & g[24944];
assign g[57711] = b[14] & g[24944];
assign g[41329] = a[14] & g[24945];
assign g[57712] = b[14] & g[24945];
assign g[41330] = a[14] & g[24946];
assign g[57713] = b[14] & g[24946];
assign g[41331] = a[14] & g[24947];
assign g[57714] = b[14] & g[24947];
assign g[41332] = a[14] & g[24948];
assign g[57715] = b[14] & g[24948];
assign g[41333] = a[14] & g[24949];
assign g[57716] = b[14] & g[24949];
assign g[41334] = a[14] & g[24950];
assign g[57717] = b[14] & g[24950];
assign g[41335] = a[14] & g[24951];
assign g[57718] = b[14] & g[24951];
assign g[41336] = a[14] & g[24952];
assign g[57719] = b[14] & g[24952];
assign g[41337] = a[14] & g[24953];
assign g[57720] = b[14] & g[24953];
assign g[41338] = a[14] & g[24954];
assign g[57721] = b[14] & g[24954];
assign g[41339] = a[14] & g[24955];
assign g[57722] = b[14] & g[24955];
assign g[41340] = a[14] & g[24956];
assign g[57723] = b[14] & g[24956];
assign g[41341] = a[14] & g[24957];
assign g[57724] = b[14] & g[24957];
assign g[41342] = a[14] & g[24958];
assign g[57725] = b[14] & g[24958];
assign g[41343] = a[14] & g[24959];
assign g[57726] = b[14] & g[24959];
assign g[41344] = a[14] & g[24960];
assign g[57727] = b[14] & g[24960];
assign g[41345] = a[14] & g[24961];
assign g[57728] = b[14] & g[24961];
assign g[41346] = a[14] & g[24962];
assign g[57729] = b[14] & g[24962];
assign g[41347] = a[14] & g[24963];
assign g[57730] = b[14] & g[24963];
assign g[41348] = a[14] & g[24964];
assign g[57731] = b[14] & g[24964];
assign g[41349] = a[14] & g[24965];
assign g[57732] = b[14] & g[24965];
assign g[41350] = a[14] & g[24966];
assign g[57733] = b[14] & g[24966];
assign g[41351] = a[14] & g[24967];
assign g[57734] = b[14] & g[24967];
assign g[41352] = a[14] & g[24968];
assign g[57735] = b[14] & g[24968];
assign g[41353] = a[14] & g[24969];
assign g[57736] = b[14] & g[24969];
assign g[41354] = a[14] & g[24970];
assign g[57737] = b[14] & g[24970];
assign g[41355] = a[14] & g[24971];
assign g[57738] = b[14] & g[24971];
assign g[41356] = a[14] & g[24972];
assign g[57739] = b[14] & g[24972];
assign g[41357] = a[14] & g[24973];
assign g[57740] = b[14] & g[24973];
assign g[41358] = a[14] & g[24974];
assign g[57741] = b[14] & g[24974];
assign g[41359] = a[14] & g[24975];
assign g[57742] = b[14] & g[24975];
assign g[41360] = a[14] & g[24976];
assign g[57743] = b[14] & g[24976];
assign g[41361] = a[14] & g[24977];
assign g[57744] = b[14] & g[24977];
assign g[41362] = a[14] & g[24978];
assign g[57745] = b[14] & g[24978];
assign g[41363] = a[14] & g[24979];
assign g[57746] = b[14] & g[24979];
assign g[41364] = a[14] & g[24980];
assign g[57747] = b[14] & g[24980];
assign g[41365] = a[14] & g[24981];
assign g[57748] = b[14] & g[24981];
assign g[41366] = a[14] & g[24982];
assign g[57749] = b[14] & g[24982];
assign g[41367] = a[14] & g[24983];
assign g[57750] = b[14] & g[24983];
assign g[41368] = a[14] & g[24984];
assign g[57751] = b[14] & g[24984];
assign g[41369] = a[14] & g[24985];
assign g[57752] = b[14] & g[24985];
assign g[41370] = a[14] & g[24986];
assign g[57753] = b[14] & g[24986];
assign g[41371] = a[14] & g[24987];
assign g[57754] = b[14] & g[24987];
assign g[41372] = a[14] & g[24988];
assign g[57755] = b[14] & g[24988];
assign g[41373] = a[14] & g[24989];
assign g[57756] = b[14] & g[24989];
assign g[41374] = a[14] & g[24990];
assign g[57757] = b[14] & g[24990];
assign g[41375] = a[14] & g[24991];
assign g[57758] = b[14] & g[24991];
assign g[41376] = a[14] & g[24992];
assign g[57759] = b[14] & g[24992];
assign g[41377] = a[14] & g[24993];
assign g[57760] = b[14] & g[24993];
assign g[41378] = a[14] & g[24994];
assign g[57761] = b[14] & g[24994];
assign g[41379] = a[14] & g[24995];
assign g[57762] = b[14] & g[24995];
assign g[41380] = a[14] & g[24996];
assign g[57763] = b[14] & g[24996];
assign g[41381] = a[14] & g[24997];
assign g[57764] = b[14] & g[24997];
assign g[41382] = a[14] & g[24998];
assign g[57765] = b[14] & g[24998];
assign g[41383] = a[14] & g[24999];
assign g[57766] = b[14] & g[24999];
assign g[41384] = a[14] & g[25000];
assign g[57767] = b[14] & g[25000];
assign g[41385] = a[14] & g[25001];
assign g[57768] = b[14] & g[25001];
assign g[41386] = a[14] & g[25002];
assign g[57769] = b[14] & g[25002];
assign g[41387] = a[14] & g[25003];
assign g[57770] = b[14] & g[25003];
assign g[41388] = a[14] & g[25004];
assign g[57771] = b[14] & g[25004];
assign g[41389] = a[14] & g[25005];
assign g[57772] = b[14] & g[25005];
assign g[41390] = a[14] & g[25006];
assign g[57773] = b[14] & g[25006];
assign g[41391] = a[14] & g[25007];
assign g[57774] = b[14] & g[25007];
assign g[41392] = a[14] & g[25008];
assign g[57775] = b[14] & g[25008];
assign g[41393] = a[14] & g[25009];
assign g[57776] = b[14] & g[25009];
assign g[41394] = a[14] & g[25010];
assign g[57777] = b[14] & g[25010];
assign g[41395] = a[14] & g[25011];
assign g[57778] = b[14] & g[25011];
assign g[41396] = a[14] & g[25012];
assign g[57779] = b[14] & g[25012];
assign g[41397] = a[14] & g[25013];
assign g[57780] = b[14] & g[25013];
assign g[41398] = a[14] & g[25014];
assign g[57781] = b[14] & g[25014];
assign g[41399] = a[14] & g[25015];
assign g[57782] = b[14] & g[25015];
assign g[41400] = a[14] & g[25016];
assign g[57783] = b[14] & g[25016];
assign g[41401] = a[14] & g[25017];
assign g[57784] = b[14] & g[25017];
assign g[41402] = a[14] & g[25018];
assign g[57785] = b[14] & g[25018];
assign g[41403] = a[14] & g[25019];
assign g[57786] = b[14] & g[25019];
assign g[41404] = a[14] & g[25020];
assign g[57787] = b[14] & g[25020];
assign g[41405] = a[14] & g[25021];
assign g[57788] = b[14] & g[25021];
assign g[41406] = a[14] & g[25022];
assign g[57789] = b[14] & g[25022];
assign g[41407] = a[14] & g[25023];
assign g[57790] = b[14] & g[25023];
assign g[41408] = a[14] & g[25024];
assign g[57791] = b[14] & g[25024];
assign g[41409] = a[14] & g[25025];
assign g[57792] = b[14] & g[25025];
assign g[41410] = a[14] & g[25026];
assign g[57793] = b[14] & g[25026];
assign g[41411] = a[14] & g[25027];
assign g[57794] = b[14] & g[25027];
assign g[41412] = a[14] & g[25028];
assign g[57795] = b[14] & g[25028];
assign g[41413] = a[14] & g[25029];
assign g[57796] = b[14] & g[25029];
assign g[41414] = a[14] & g[25030];
assign g[57797] = b[14] & g[25030];
assign g[41415] = a[14] & g[25031];
assign g[57798] = b[14] & g[25031];
assign g[41416] = a[14] & g[25032];
assign g[57799] = b[14] & g[25032];
assign g[41417] = a[14] & g[25033];
assign g[57800] = b[14] & g[25033];
assign g[41418] = a[14] & g[25034];
assign g[57801] = b[14] & g[25034];
assign g[41419] = a[14] & g[25035];
assign g[57802] = b[14] & g[25035];
assign g[41420] = a[14] & g[25036];
assign g[57803] = b[14] & g[25036];
assign g[41421] = a[14] & g[25037];
assign g[57804] = b[14] & g[25037];
assign g[41422] = a[14] & g[25038];
assign g[57805] = b[14] & g[25038];
assign g[41423] = a[14] & g[25039];
assign g[57806] = b[14] & g[25039];
assign g[41424] = a[14] & g[25040];
assign g[57807] = b[14] & g[25040];
assign g[41425] = a[14] & g[25041];
assign g[57808] = b[14] & g[25041];
assign g[41426] = a[14] & g[25042];
assign g[57809] = b[14] & g[25042];
assign g[41427] = a[14] & g[25043];
assign g[57810] = b[14] & g[25043];
assign g[41428] = a[14] & g[25044];
assign g[57811] = b[14] & g[25044];
assign g[41429] = a[14] & g[25045];
assign g[57812] = b[14] & g[25045];
assign g[41430] = a[14] & g[25046];
assign g[57813] = b[14] & g[25046];
assign g[41431] = a[14] & g[25047];
assign g[57814] = b[14] & g[25047];
assign g[41432] = a[14] & g[25048];
assign g[57815] = b[14] & g[25048];
assign g[41433] = a[14] & g[25049];
assign g[57816] = b[14] & g[25049];
assign g[41434] = a[14] & g[25050];
assign g[57817] = b[14] & g[25050];
assign g[41435] = a[14] & g[25051];
assign g[57818] = b[14] & g[25051];
assign g[41436] = a[14] & g[25052];
assign g[57819] = b[14] & g[25052];
assign g[41437] = a[14] & g[25053];
assign g[57820] = b[14] & g[25053];
assign g[41438] = a[14] & g[25054];
assign g[57821] = b[14] & g[25054];
assign g[41439] = a[14] & g[25055];
assign g[57822] = b[14] & g[25055];
assign g[41440] = a[14] & g[25056];
assign g[57823] = b[14] & g[25056];
assign g[41441] = a[14] & g[25057];
assign g[57824] = b[14] & g[25057];
assign g[41442] = a[14] & g[25058];
assign g[57825] = b[14] & g[25058];
assign g[41443] = a[14] & g[25059];
assign g[57826] = b[14] & g[25059];
assign g[41444] = a[14] & g[25060];
assign g[57827] = b[14] & g[25060];
assign g[41445] = a[14] & g[25061];
assign g[57828] = b[14] & g[25061];
assign g[41446] = a[14] & g[25062];
assign g[57829] = b[14] & g[25062];
assign g[41447] = a[14] & g[25063];
assign g[57830] = b[14] & g[25063];
assign g[41448] = a[14] & g[25064];
assign g[57831] = b[14] & g[25064];
assign g[41449] = a[14] & g[25065];
assign g[57832] = b[14] & g[25065];
assign g[41450] = a[14] & g[25066];
assign g[57833] = b[14] & g[25066];
assign g[41451] = a[14] & g[25067];
assign g[57834] = b[14] & g[25067];
assign g[41452] = a[14] & g[25068];
assign g[57835] = b[14] & g[25068];
assign g[41453] = a[14] & g[25069];
assign g[57836] = b[14] & g[25069];
assign g[41454] = a[14] & g[25070];
assign g[57837] = b[14] & g[25070];
assign g[41455] = a[14] & g[25071];
assign g[57838] = b[14] & g[25071];
assign g[41456] = a[14] & g[25072];
assign g[57839] = b[14] & g[25072];
assign g[41457] = a[14] & g[25073];
assign g[57840] = b[14] & g[25073];
assign g[41458] = a[14] & g[25074];
assign g[57841] = b[14] & g[25074];
assign g[41459] = a[14] & g[25075];
assign g[57842] = b[14] & g[25075];
assign g[41460] = a[14] & g[25076];
assign g[57843] = b[14] & g[25076];
assign g[41461] = a[14] & g[25077];
assign g[57844] = b[14] & g[25077];
assign g[41462] = a[14] & g[25078];
assign g[57845] = b[14] & g[25078];
assign g[41463] = a[14] & g[25079];
assign g[57846] = b[14] & g[25079];
assign g[41464] = a[14] & g[25080];
assign g[57847] = b[14] & g[25080];
assign g[41465] = a[14] & g[25081];
assign g[57848] = b[14] & g[25081];
assign g[41466] = a[14] & g[25082];
assign g[57849] = b[14] & g[25082];
assign g[41467] = a[14] & g[25083];
assign g[57850] = b[14] & g[25083];
assign g[41468] = a[14] & g[25084];
assign g[57851] = b[14] & g[25084];
assign g[41469] = a[14] & g[25085];
assign g[57852] = b[14] & g[25085];
assign g[41470] = a[14] & g[25086];
assign g[57853] = b[14] & g[25086];
assign g[41471] = a[14] & g[25087];
assign g[57854] = b[14] & g[25087];
assign g[41472] = a[14] & g[25088];
assign g[57855] = b[14] & g[25088];
assign g[41473] = a[14] & g[25089];
assign g[57856] = b[14] & g[25089];
assign g[41474] = a[14] & g[25090];
assign g[57857] = b[14] & g[25090];
assign g[41475] = a[14] & g[25091];
assign g[57858] = b[14] & g[25091];
assign g[41476] = a[14] & g[25092];
assign g[57859] = b[14] & g[25092];
assign g[41477] = a[14] & g[25093];
assign g[57860] = b[14] & g[25093];
assign g[41478] = a[14] & g[25094];
assign g[57861] = b[14] & g[25094];
assign g[41479] = a[14] & g[25095];
assign g[57862] = b[14] & g[25095];
assign g[41480] = a[14] & g[25096];
assign g[57863] = b[14] & g[25096];
assign g[41481] = a[14] & g[25097];
assign g[57864] = b[14] & g[25097];
assign g[41482] = a[14] & g[25098];
assign g[57865] = b[14] & g[25098];
assign g[41483] = a[14] & g[25099];
assign g[57866] = b[14] & g[25099];
assign g[41484] = a[14] & g[25100];
assign g[57867] = b[14] & g[25100];
assign g[41485] = a[14] & g[25101];
assign g[57868] = b[14] & g[25101];
assign g[41486] = a[14] & g[25102];
assign g[57869] = b[14] & g[25102];
assign g[41487] = a[14] & g[25103];
assign g[57870] = b[14] & g[25103];
assign g[41488] = a[14] & g[25104];
assign g[57871] = b[14] & g[25104];
assign g[41489] = a[14] & g[25105];
assign g[57872] = b[14] & g[25105];
assign g[41490] = a[14] & g[25106];
assign g[57873] = b[14] & g[25106];
assign g[41491] = a[14] & g[25107];
assign g[57874] = b[14] & g[25107];
assign g[41492] = a[14] & g[25108];
assign g[57875] = b[14] & g[25108];
assign g[41493] = a[14] & g[25109];
assign g[57876] = b[14] & g[25109];
assign g[41494] = a[14] & g[25110];
assign g[57877] = b[14] & g[25110];
assign g[41495] = a[14] & g[25111];
assign g[57878] = b[14] & g[25111];
assign g[41496] = a[14] & g[25112];
assign g[57879] = b[14] & g[25112];
assign g[41497] = a[14] & g[25113];
assign g[57880] = b[14] & g[25113];
assign g[41498] = a[14] & g[25114];
assign g[57881] = b[14] & g[25114];
assign g[41499] = a[14] & g[25115];
assign g[57882] = b[14] & g[25115];
assign g[41500] = a[14] & g[25116];
assign g[57883] = b[14] & g[25116];
assign g[41501] = a[14] & g[25117];
assign g[57884] = b[14] & g[25117];
assign g[41502] = a[14] & g[25118];
assign g[57885] = b[14] & g[25118];
assign g[41503] = a[14] & g[25119];
assign g[57886] = b[14] & g[25119];
assign g[41504] = a[14] & g[25120];
assign g[57887] = b[14] & g[25120];
assign g[41505] = a[14] & g[25121];
assign g[57888] = b[14] & g[25121];
assign g[41506] = a[14] & g[25122];
assign g[57889] = b[14] & g[25122];
assign g[41507] = a[14] & g[25123];
assign g[57890] = b[14] & g[25123];
assign g[41508] = a[14] & g[25124];
assign g[57891] = b[14] & g[25124];
assign g[41509] = a[14] & g[25125];
assign g[57892] = b[14] & g[25125];
assign g[41510] = a[14] & g[25126];
assign g[57893] = b[14] & g[25126];
assign g[41511] = a[14] & g[25127];
assign g[57894] = b[14] & g[25127];
assign g[41512] = a[14] & g[25128];
assign g[57895] = b[14] & g[25128];
assign g[41513] = a[14] & g[25129];
assign g[57896] = b[14] & g[25129];
assign g[41514] = a[14] & g[25130];
assign g[57897] = b[14] & g[25130];
assign g[41515] = a[14] & g[25131];
assign g[57898] = b[14] & g[25131];
assign g[41516] = a[14] & g[25132];
assign g[57899] = b[14] & g[25132];
assign g[41517] = a[14] & g[25133];
assign g[57900] = b[14] & g[25133];
assign g[41518] = a[14] & g[25134];
assign g[57901] = b[14] & g[25134];
assign g[41519] = a[14] & g[25135];
assign g[57902] = b[14] & g[25135];
assign g[41520] = a[14] & g[25136];
assign g[57903] = b[14] & g[25136];
assign g[41521] = a[14] & g[25137];
assign g[57904] = b[14] & g[25137];
assign g[41522] = a[14] & g[25138];
assign g[57905] = b[14] & g[25138];
assign g[41523] = a[14] & g[25139];
assign g[57906] = b[14] & g[25139];
assign g[41524] = a[14] & g[25140];
assign g[57907] = b[14] & g[25140];
assign g[41525] = a[14] & g[25141];
assign g[57908] = b[14] & g[25141];
assign g[41526] = a[14] & g[25142];
assign g[57909] = b[14] & g[25142];
assign g[41527] = a[14] & g[25143];
assign g[57910] = b[14] & g[25143];
assign g[41528] = a[14] & g[25144];
assign g[57911] = b[14] & g[25144];
assign g[41529] = a[14] & g[25145];
assign g[57912] = b[14] & g[25145];
assign g[41530] = a[14] & g[25146];
assign g[57913] = b[14] & g[25146];
assign g[41531] = a[14] & g[25147];
assign g[57914] = b[14] & g[25147];
assign g[41532] = a[14] & g[25148];
assign g[57915] = b[14] & g[25148];
assign g[41533] = a[14] & g[25149];
assign g[57916] = b[14] & g[25149];
assign g[41534] = a[14] & g[25150];
assign g[57917] = b[14] & g[25150];
assign g[41535] = a[14] & g[25151];
assign g[57918] = b[14] & g[25151];
assign g[41536] = a[14] & g[25152];
assign g[57919] = b[14] & g[25152];
assign g[41537] = a[14] & g[25153];
assign g[57920] = b[14] & g[25153];
assign g[41538] = a[14] & g[25154];
assign g[57921] = b[14] & g[25154];
assign g[41539] = a[14] & g[25155];
assign g[57922] = b[14] & g[25155];
assign g[41540] = a[14] & g[25156];
assign g[57923] = b[14] & g[25156];
assign g[41541] = a[14] & g[25157];
assign g[57924] = b[14] & g[25157];
assign g[41542] = a[14] & g[25158];
assign g[57925] = b[14] & g[25158];
assign g[41543] = a[14] & g[25159];
assign g[57926] = b[14] & g[25159];
assign g[41544] = a[14] & g[25160];
assign g[57927] = b[14] & g[25160];
assign g[41545] = a[14] & g[25161];
assign g[57928] = b[14] & g[25161];
assign g[41546] = a[14] & g[25162];
assign g[57929] = b[14] & g[25162];
assign g[41547] = a[14] & g[25163];
assign g[57930] = b[14] & g[25163];
assign g[41548] = a[14] & g[25164];
assign g[57931] = b[14] & g[25164];
assign g[41549] = a[14] & g[25165];
assign g[57932] = b[14] & g[25165];
assign g[41550] = a[14] & g[25166];
assign g[57933] = b[14] & g[25166];
assign g[41551] = a[14] & g[25167];
assign g[57934] = b[14] & g[25167];
assign g[41552] = a[14] & g[25168];
assign g[57935] = b[14] & g[25168];
assign g[41553] = a[14] & g[25169];
assign g[57936] = b[14] & g[25169];
assign g[41554] = a[14] & g[25170];
assign g[57937] = b[14] & g[25170];
assign g[41555] = a[14] & g[25171];
assign g[57938] = b[14] & g[25171];
assign g[41556] = a[14] & g[25172];
assign g[57939] = b[14] & g[25172];
assign g[41557] = a[14] & g[25173];
assign g[57940] = b[14] & g[25173];
assign g[41558] = a[14] & g[25174];
assign g[57941] = b[14] & g[25174];
assign g[41559] = a[14] & g[25175];
assign g[57942] = b[14] & g[25175];
assign g[41560] = a[14] & g[25176];
assign g[57943] = b[14] & g[25176];
assign g[41561] = a[14] & g[25177];
assign g[57944] = b[14] & g[25177];
assign g[41562] = a[14] & g[25178];
assign g[57945] = b[14] & g[25178];
assign g[41563] = a[14] & g[25179];
assign g[57946] = b[14] & g[25179];
assign g[41564] = a[14] & g[25180];
assign g[57947] = b[14] & g[25180];
assign g[41565] = a[14] & g[25181];
assign g[57948] = b[14] & g[25181];
assign g[41566] = a[14] & g[25182];
assign g[57949] = b[14] & g[25182];
assign g[41567] = a[14] & g[25183];
assign g[57950] = b[14] & g[25183];
assign g[41568] = a[14] & g[25184];
assign g[57951] = b[14] & g[25184];
assign g[41569] = a[14] & g[25185];
assign g[57952] = b[14] & g[25185];
assign g[41570] = a[14] & g[25186];
assign g[57953] = b[14] & g[25186];
assign g[41571] = a[14] & g[25187];
assign g[57954] = b[14] & g[25187];
assign g[41572] = a[14] & g[25188];
assign g[57955] = b[14] & g[25188];
assign g[41573] = a[14] & g[25189];
assign g[57956] = b[14] & g[25189];
assign g[41574] = a[14] & g[25190];
assign g[57957] = b[14] & g[25190];
assign g[41575] = a[14] & g[25191];
assign g[57958] = b[14] & g[25191];
assign g[41576] = a[14] & g[25192];
assign g[57959] = b[14] & g[25192];
assign g[41577] = a[14] & g[25193];
assign g[57960] = b[14] & g[25193];
assign g[41578] = a[14] & g[25194];
assign g[57961] = b[14] & g[25194];
assign g[41579] = a[14] & g[25195];
assign g[57962] = b[14] & g[25195];
assign g[41580] = a[14] & g[25196];
assign g[57963] = b[14] & g[25196];
assign g[41581] = a[14] & g[25197];
assign g[57964] = b[14] & g[25197];
assign g[41582] = a[14] & g[25198];
assign g[57965] = b[14] & g[25198];
assign g[41583] = a[14] & g[25199];
assign g[57966] = b[14] & g[25199];
assign g[41584] = a[14] & g[25200];
assign g[57967] = b[14] & g[25200];
assign g[41585] = a[14] & g[25201];
assign g[57968] = b[14] & g[25201];
assign g[41586] = a[14] & g[25202];
assign g[57969] = b[14] & g[25202];
assign g[41587] = a[14] & g[25203];
assign g[57970] = b[14] & g[25203];
assign g[41588] = a[14] & g[25204];
assign g[57971] = b[14] & g[25204];
assign g[41589] = a[14] & g[25205];
assign g[57972] = b[14] & g[25205];
assign g[41590] = a[14] & g[25206];
assign g[57973] = b[14] & g[25206];
assign g[41591] = a[14] & g[25207];
assign g[57974] = b[14] & g[25207];
assign g[41592] = a[14] & g[25208];
assign g[57975] = b[14] & g[25208];
assign g[41593] = a[14] & g[25209];
assign g[57976] = b[14] & g[25209];
assign g[41594] = a[14] & g[25210];
assign g[57977] = b[14] & g[25210];
assign g[41595] = a[14] & g[25211];
assign g[57978] = b[14] & g[25211];
assign g[41596] = a[14] & g[25212];
assign g[57979] = b[14] & g[25212];
assign g[41597] = a[14] & g[25213];
assign g[57980] = b[14] & g[25213];
assign g[41598] = a[14] & g[25214];
assign g[57981] = b[14] & g[25214];
assign g[41599] = a[14] & g[25215];
assign g[57982] = b[14] & g[25215];
assign g[41600] = a[14] & g[25216];
assign g[57983] = b[14] & g[25216];
assign g[41601] = a[14] & g[25217];
assign g[57984] = b[14] & g[25217];
assign g[41602] = a[14] & g[25218];
assign g[57985] = b[14] & g[25218];
assign g[41603] = a[14] & g[25219];
assign g[57986] = b[14] & g[25219];
assign g[41604] = a[14] & g[25220];
assign g[57987] = b[14] & g[25220];
assign g[41605] = a[14] & g[25221];
assign g[57988] = b[14] & g[25221];
assign g[41606] = a[14] & g[25222];
assign g[57989] = b[14] & g[25222];
assign g[41607] = a[14] & g[25223];
assign g[57990] = b[14] & g[25223];
assign g[41608] = a[14] & g[25224];
assign g[57991] = b[14] & g[25224];
assign g[41609] = a[14] & g[25225];
assign g[57992] = b[14] & g[25225];
assign g[41610] = a[14] & g[25226];
assign g[57993] = b[14] & g[25226];
assign g[41611] = a[14] & g[25227];
assign g[57994] = b[14] & g[25227];
assign g[41612] = a[14] & g[25228];
assign g[57995] = b[14] & g[25228];
assign g[41613] = a[14] & g[25229];
assign g[57996] = b[14] & g[25229];
assign g[41614] = a[14] & g[25230];
assign g[57997] = b[14] & g[25230];
assign g[41615] = a[14] & g[25231];
assign g[57998] = b[14] & g[25231];
assign g[41616] = a[14] & g[25232];
assign g[57999] = b[14] & g[25232];
assign g[41617] = a[14] & g[25233];
assign g[58000] = b[14] & g[25233];
assign g[41618] = a[14] & g[25234];
assign g[58001] = b[14] & g[25234];
assign g[41619] = a[14] & g[25235];
assign g[58002] = b[14] & g[25235];
assign g[41620] = a[14] & g[25236];
assign g[58003] = b[14] & g[25236];
assign g[41621] = a[14] & g[25237];
assign g[58004] = b[14] & g[25237];
assign g[41622] = a[14] & g[25238];
assign g[58005] = b[14] & g[25238];
assign g[41623] = a[14] & g[25239];
assign g[58006] = b[14] & g[25239];
assign g[41624] = a[14] & g[25240];
assign g[58007] = b[14] & g[25240];
assign g[41625] = a[14] & g[25241];
assign g[58008] = b[14] & g[25241];
assign g[41626] = a[14] & g[25242];
assign g[58009] = b[14] & g[25242];
assign g[41627] = a[14] & g[25243];
assign g[58010] = b[14] & g[25243];
assign g[41628] = a[14] & g[25244];
assign g[58011] = b[14] & g[25244];
assign g[41629] = a[14] & g[25245];
assign g[58012] = b[14] & g[25245];
assign g[41630] = a[14] & g[25246];
assign g[58013] = b[14] & g[25246];
assign g[41631] = a[14] & g[25247];
assign g[58014] = b[14] & g[25247];
assign g[41632] = a[14] & g[25248];
assign g[58015] = b[14] & g[25248];
assign g[41633] = a[14] & g[25249];
assign g[58016] = b[14] & g[25249];
assign g[41634] = a[14] & g[25250];
assign g[58017] = b[14] & g[25250];
assign g[41635] = a[14] & g[25251];
assign g[58018] = b[14] & g[25251];
assign g[41636] = a[14] & g[25252];
assign g[58019] = b[14] & g[25252];
assign g[41637] = a[14] & g[25253];
assign g[58020] = b[14] & g[25253];
assign g[41638] = a[14] & g[25254];
assign g[58021] = b[14] & g[25254];
assign g[41639] = a[14] & g[25255];
assign g[58022] = b[14] & g[25255];
assign g[41640] = a[14] & g[25256];
assign g[58023] = b[14] & g[25256];
assign g[41641] = a[14] & g[25257];
assign g[58024] = b[14] & g[25257];
assign g[41642] = a[14] & g[25258];
assign g[58025] = b[14] & g[25258];
assign g[41643] = a[14] & g[25259];
assign g[58026] = b[14] & g[25259];
assign g[41644] = a[14] & g[25260];
assign g[58027] = b[14] & g[25260];
assign g[41645] = a[14] & g[25261];
assign g[58028] = b[14] & g[25261];
assign g[41646] = a[14] & g[25262];
assign g[58029] = b[14] & g[25262];
assign g[41647] = a[14] & g[25263];
assign g[58030] = b[14] & g[25263];
assign g[41648] = a[14] & g[25264];
assign g[58031] = b[14] & g[25264];
assign g[41649] = a[14] & g[25265];
assign g[58032] = b[14] & g[25265];
assign g[41650] = a[14] & g[25266];
assign g[58033] = b[14] & g[25266];
assign g[41651] = a[14] & g[25267];
assign g[58034] = b[14] & g[25267];
assign g[41652] = a[14] & g[25268];
assign g[58035] = b[14] & g[25268];
assign g[41653] = a[14] & g[25269];
assign g[58036] = b[14] & g[25269];
assign g[41654] = a[14] & g[25270];
assign g[58037] = b[14] & g[25270];
assign g[41655] = a[14] & g[25271];
assign g[58038] = b[14] & g[25271];
assign g[41656] = a[14] & g[25272];
assign g[58039] = b[14] & g[25272];
assign g[41657] = a[14] & g[25273];
assign g[58040] = b[14] & g[25273];
assign g[41658] = a[14] & g[25274];
assign g[58041] = b[14] & g[25274];
assign g[41659] = a[14] & g[25275];
assign g[58042] = b[14] & g[25275];
assign g[41660] = a[14] & g[25276];
assign g[58043] = b[14] & g[25276];
assign g[41661] = a[14] & g[25277];
assign g[58044] = b[14] & g[25277];
assign g[41662] = a[14] & g[25278];
assign g[58045] = b[14] & g[25278];
assign g[41663] = a[14] & g[25279];
assign g[58046] = b[14] & g[25279];
assign g[41664] = a[14] & g[25280];
assign g[58047] = b[14] & g[25280];
assign g[41665] = a[14] & g[25281];
assign g[58048] = b[14] & g[25281];
assign g[41666] = a[14] & g[25282];
assign g[58049] = b[14] & g[25282];
assign g[41667] = a[14] & g[25283];
assign g[58050] = b[14] & g[25283];
assign g[41668] = a[14] & g[25284];
assign g[58051] = b[14] & g[25284];
assign g[41669] = a[14] & g[25285];
assign g[58052] = b[14] & g[25285];
assign g[41670] = a[14] & g[25286];
assign g[58053] = b[14] & g[25286];
assign g[41671] = a[14] & g[25287];
assign g[58054] = b[14] & g[25287];
assign g[41672] = a[14] & g[25288];
assign g[58055] = b[14] & g[25288];
assign g[41673] = a[14] & g[25289];
assign g[58056] = b[14] & g[25289];
assign g[41674] = a[14] & g[25290];
assign g[58057] = b[14] & g[25290];
assign g[41675] = a[14] & g[25291];
assign g[58058] = b[14] & g[25291];
assign g[41676] = a[14] & g[25292];
assign g[58059] = b[14] & g[25292];
assign g[41677] = a[14] & g[25293];
assign g[58060] = b[14] & g[25293];
assign g[41678] = a[14] & g[25294];
assign g[58061] = b[14] & g[25294];
assign g[41679] = a[14] & g[25295];
assign g[58062] = b[14] & g[25295];
assign g[41680] = a[14] & g[25296];
assign g[58063] = b[14] & g[25296];
assign g[41681] = a[14] & g[25297];
assign g[58064] = b[14] & g[25297];
assign g[41682] = a[14] & g[25298];
assign g[58065] = b[14] & g[25298];
assign g[41683] = a[14] & g[25299];
assign g[58066] = b[14] & g[25299];
assign g[41684] = a[14] & g[25300];
assign g[58067] = b[14] & g[25300];
assign g[41685] = a[14] & g[25301];
assign g[58068] = b[14] & g[25301];
assign g[41686] = a[14] & g[25302];
assign g[58069] = b[14] & g[25302];
assign g[41687] = a[14] & g[25303];
assign g[58070] = b[14] & g[25303];
assign g[41688] = a[14] & g[25304];
assign g[58071] = b[14] & g[25304];
assign g[41689] = a[14] & g[25305];
assign g[58072] = b[14] & g[25305];
assign g[41690] = a[14] & g[25306];
assign g[58073] = b[14] & g[25306];
assign g[41691] = a[14] & g[25307];
assign g[58074] = b[14] & g[25307];
assign g[41692] = a[14] & g[25308];
assign g[58075] = b[14] & g[25308];
assign g[41693] = a[14] & g[25309];
assign g[58076] = b[14] & g[25309];
assign g[41694] = a[14] & g[25310];
assign g[58077] = b[14] & g[25310];
assign g[41695] = a[14] & g[25311];
assign g[58078] = b[14] & g[25311];
assign g[41696] = a[14] & g[25312];
assign g[58079] = b[14] & g[25312];
assign g[41697] = a[14] & g[25313];
assign g[58080] = b[14] & g[25313];
assign g[41698] = a[14] & g[25314];
assign g[58081] = b[14] & g[25314];
assign g[41699] = a[14] & g[25315];
assign g[58082] = b[14] & g[25315];
assign g[41700] = a[14] & g[25316];
assign g[58083] = b[14] & g[25316];
assign g[41701] = a[14] & g[25317];
assign g[58084] = b[14] & g[25317];
assign g[41702] = a[14] & g[25318];
assign g[58085] = b[14] & g[25318];
assign g[41703] = a[14] & g[25319];
assign g[58086] = b[14] & g[25319];
assign g[41704] = a[14] & g[25320];
assign g[58087] = b[14] & g[25320];
assign g[41705] = a[14] & g[25321];
assign g[58088] = b[14] & g[25321];
assign g[41706] = a[14] & g[25322];
assign g[58089] = b[14] & g[25322];
assign g[41707] = a[14] & g[25323];
assign g[58090] = b[14] & g[25323];
assign g[41708] = a[14] & g[25324];
assign g[58091] = b[14] & g[25324];
assign g[41709] = a[14] & g[25325];
assign g[58092] = b[14] & g[25325];
assign g[41710] = a[14] & g[25326];
assign g[58093] = b[14] & g[25326];
assign g[41711] = a[14] & g[25327];
assign g[58094] = b[14] & g[25327];
assign g[41712] = a[14] & g[25328];
assign g[58095] = b[14] & g[25328];
assign g[41713] = a[14] & g[25329];
assign g[58096] = b[14] & g[25329];
assign g[41714] = a[14] & g[25330];
assign g[58097] = b[14] & g[25330];
assign g[41715] = a[14] & g[25331];
assign g[58098] = b[14] & g[25331];
assign g[41716] = a[14] & g[25332];
assign g[58099] = b[14] & g[25332];
assign g[41717] = a[14] & g[25333];
assign g[58100] = b[14] & g[25333];
assign g[41718] = a[14] & g[25334];
assign g[58101] = b[14] & g[25334];
assign g[41719] = a[14] & g[25335];
assign g[58102] = b[14] & g[25335];
assign g[41720] = a[14] & g[25336];
assign g[58103] = b[14] & g[25336];
assign g[41721] = a[14] & g[25337];
assign g[58104] = b[14] & g[25337];
assign g[41722] = a[14] & g[25338];
assign g[58105] = b[14] & g[25338];
assign g[41723] = a[14] & g[25339];
assign g[58106] = b[14] & g[25339];
assign g[41724] = a[14] & g[25340];
assign g[58107] = b[14] & g[25340];
assign g[41725] = a[14] & g[25341];
assign g[58108] = b[14] & g[25341];
assign g[41726] = a[14] & g[25342];
assign g[58109] = b[14] & g[25342];
assign g[41727] = a[14] & g[25343];
assign g[58110] = b[14] & g[25343];
assign g[41728] = a[14] & g[25344];
assign g[58111] = b[14] & g[25344];
assign g[41729] = a[14] & g[25345];
assign g[58112] = b[14] & g[25345];
assign g[41730] = a[14] & g[25346];
assign g[58113] = b[14] & g[25346];
assign g[41731] = a[14] & g[25347];
assign g[58114] = b[14] & g[25347];
assign g[41732] = a[14] & g[25348];
assign g[58115] = b[14] & g[25348];
assign g[41733] = a[14] & g[25349];
assign g[58116] = b[14] & g[25349];
assign g[41734] = a[14] & g[25350];
assign g[58117] = b[14] & g[25350];
assign g[41735] = a[14] & g[25351];
assign g[58118] = b[14] & g[25351];
assign g[41736] = a[14] & g[25352];
assign g[58119] = b[14] & g[25352];
assign g[41737] = a[14] & g[25353];
assign g[58120] = b[14] & g[25353];
assign g[41738] = a[14] & g[25354];
assign g[58121] = b[14] & g[25354];
assign g[41739] = a[14] & g[25355];
assign g[58122] = b[14] & g[25355];
assign g[41740] = a[14] & g[25356];
assign g[58123] = b[14] & g[25356];
assign g[41741] = a[14] & g[25357];
assign g[58124] = b[14] & g[25357];
assign g[41742] = a[14] & g[25358];
assign g[58125] = b[14] & g[25358];
assign g[41743] = a[14] & g[25359];
assign g[58126] = b[14] & g[25359];
assign g[41744] = a[14] & g[25360];
assign g[58127] = b[14] & g[25360];
assign g[41745] = a[14] & g[25361];
assign g[58128] = b[14] & g[25361];
assign g[41746] = a[14] & g[25362];
assign g[58129] = b[14] & g[25362];
assign g[41747] = a[14] & g[25363];
assign g[58130] = b[14] & g[25363];
assign g[41748] = a[14] & g[25364];
assign g[58131] = b[14] & g[25364];
assign g[41749] = a[14] & g[25365];
assign g[58132] = b[14] & g[25365];
assign g[41750] = a[14] & g[25366];
assign g[58133] = b[14] & g[25366];
assign g[41751] = a[14] & g[25367];
assign g[58134] = b[14] & g[25367];
assign g[41752] = a[14] & g[25368];
assign g[58135] = b[14] & g[25368];
assign g[41753] = a[14] & g[25369];
assign g[58136] = b[14] & g[25369];
assign g[41754] = a[14] & g[25370];
assign g[58137] = b[14] & g[25370];
assign g[41755] = a[14] & g[25371];
assign g[58138] = b[14] & g[25371];
assign g[41756] = a[14] & g[25372];
assign g[58139] = b[14] & g[25372];
assign g[41757] = a[14] & g[25373];
assign g[58140] = b[14] & g[25373];
assign g[41758] = a[14] & g[25374];
assign g[58141] = b[14] & g[25374];
assign g[41759] = a[14] & g[25375];
assign g[58142] = b[14] & g[25375];
assign g[41760] = a[14] & g[25376];
assign g[58143] = b[14] & g[25376];
assign g[41761] = a[14] & g[25377];
assign g[58144] = b[14] & g[25377];
assign g[41762] = a[14] & g[25378];
assign g[58145] = b[14] & g[25378];
assign g[41763] = a[14] & g[25379];
assign g[58146] = b[14] & g[25379];
assign g[41764] = a[14] & g[25380];
assign g[58147] = b[14] & g[25380];
assign g[41765] = a[14] & g[25381];
assign g[58148] = b[14] & g[25381];
assign g[41766] = a[14] & g[25382];
assign g[58149] = b[14] & g[25382];
assign g[41767] = a[14] & g[25383];
assign g[58150] = b[14] & g[25383];
assign g[41768] = a[14] & g[25384];
assign g[58151] = b[14] & g[25384];
assign g[41769] = a[14] & g[25385];
assign g[58152] = b[14] & g[25385];
assign g[41770] = a[14] & g[25386];
assign g[58153] = b[14] & g[25386];
assign g[41771] = a[14] & g[25387];
assign g[58154] = b[14] & g[25387];
assign g[41772] = a[14] & g[25388];
assign g[58155] = b[14] & g[25388];
assign g[41773] = a[14] & g[25389];
assign g[58156] = b[14] & g[25389];
assign g[41774] = a[14] & g[25390];
assign g[58157] = b[14] & g[25390];
assign g[41775] = a[14] & g[25391];
assign g[58158] = b[14] & g[25391];
assign g[41776] = a[14] & g[25392];
assign g[58159] = b[14] & g[25392];
assign g[41777] = a[14] & g[25393];
assign g[58160] = b[14] & g[25393];
assign g[41778] = a[14] & g[25394];
assign g[58161] = b[14] & g[25394];
assign g[41779] = a[14] & g[25395];
assign g[58162] = b[14] & g[25395];
assign g[41780] = a[14] & g[25396];
assign g[58163] = b[14] & g[25396];
assign g[41781] = a[14] & g[25397];
assign g[58164] = b[14] & g[25397];
assign g[41782] = a[14] & g[25398];
assign g[58165] = b[14] & g[25398];
assign g[41783] = a[14] & g[25399];
assign g[58166] = b[14] & g[25399];
assign g[41784] = a[14] & g[25400];
assign g[58167] = b[14] & g[25400];
assign g[41785] = a[14] & g[25401];
assign g[58168] = b[14] & g[25401];
assign g[41786] = a[14] & g[25402];
assign g[58169] = b[14] & g[25402];
assign g[41787] = a[14] & g[25403];
assign g[58170] = b[14] & g[25403];
assign g[41788] = a[14] & g[25404];
assign g[58171] = b[14] & g[25404];
assign g[41789] = a[14] & g[25405];
assign g[58172] = b[14] & g[25405];
assign g[41790] = a[14] & g[25406];
assign g[58173] = b[14] & g[25406];
assign g[41791] = a[14] & g[25407];
assign g[58174] = b[14] & g[25407];
assign g[41792] = a[14] & g[25408];
assign g[58175] = b[14] & g[25408];
assign g[41793] = a[14] & g[25409];
assign g[58176] = b[14] & g[25409];
assign g[41794] = a[14] & g[25410];
assign g[58177] = b[14] & g[25410];
assign g[41795] = a[14] & g[25411];
assign g[58178] = b[14] & g[25411];
assign g[41796] = a[14] & g[25412];
assign g[58179] = b[14] & g[25412];
assign g[41797] = a[14] & g[25413];
assign g[58180] = b[14] & g[25413];
assign g[41798] = a[14] & g[25414];
assign g[58181] = b[14] & g[25414];
assign g[41799] = a[14] & g[25415];
assign g[58182] = b[14] & g[25415];
assign g[41800] = a[14] & g[25416];
assign g[58183] = b[14] & g[25416];
assign g[41801] = a[14] & g[25417];
assign g[58184] = b[14] & g[25417];
assign g[41802] = a[14] & g[25418];
assign g[58185] = b[14] & g[25418];
assign g[41803] = a[14] & g[25419];
assign g[58186] = b[14] & g[25419];
assign g[41804] = a[14] & g[25420];
assign g[58187] = b[14] & g[25420];
assign g[41805] = a[14] & g[25421];
assign g[58188] = b[14] & g[25421];
assign g[41806] = a[14] & g[25422];
assign g[58189] = b[14] & g[25422];
assign g[41807] = a[14] & g[25423];
assign g[58190] = b[14] & g[25423];
assign g[41808] = a[14] & g[25424];
assign g[58191] = b[14] & g[25424];
assign g[41809] = a[14] & g[25425];
assign g[58192] = b[14] & g[25425];
assign g[41810] = a[14] & g[25426];
assign g[58193] = b[14] & g[25426];
assign g[41811] = a[14] & g[25427];
assign g[58194] = b[14] & g[25427];
assign g[41812] = a[14] & g[25428];
assign g[58195] = b[14] & g[25428];
assign g[41813] = a[14] & g[25429];
assign g[58196] = b[14] & g[25429];
assign g[41814] = a[14] & g[25430];
assign g[58197] = b[14] & g[25430];
assign g[41815] = a[14] & g[25431];
assign g[58198] = b[14] & g[25431];
assign g[41816] = a[14] & g[25432];
assign g[58199] = b[14] & g[25432];
assign g[41817] = a[14] & g[25433];
assign g[58200] = b[14] & g[25433];
assign g[41818] = a[14] & g[25434];
assign g[58201] = b[14] & g[25434];
assign g[41819] = a[14] & g[25435];
assign g[58202] = b[14] & g[25435];
assign g[41820] = a[14] & g[25436];
assign g[58203] = b[14] & g[25436];
assign g[41821] = a[14] & g[25437];
assign g[58204] = b[14] & g[25437];
assign g[41822] = a[14] & g[25438];
assign g[58205] = b[14] & g[25438];
assign g[41823] = a[14] & g[25439];
assign g[58206] = b[14] & g[25439];
assign g[41824] = a[14] & g[25440];
assign g[58207] = b[14] & g[25440];
assign g[41825] = a[14] & g[25441];
assign g[58208] = b[14] & g[25441];
assign g[41826] = a[14] & g[25442];
assign g[58209] = b[14] & g[25442];
assign g[41827] = a[14] & g[25443];
assign g[58210] = b[14] & g[25443];
assign g[41828] = a[14] & g[25444];
assign g[58211] = b[14] & g[25444];
assign g[41829] = a[14] & g[25445];
assign g[58212] = b[14] & g[25445];
assign g[41830] = a[14] & g[25446];
assign g[58213] = b[14] & g[25446];
assign g[41831] = a[14] & g[25447];
assign g[58214] = b[14] & g[25447];
assign g[41832] = a[14] & g[25448];
assign g[58215] = b[14] & g[25448];
assign g[41833] = a[14] & g[25449];
assign g[58216] = b[14] & g[25449];
assign g[41834] = a[14] & g[25450];
assign g[58217] = b[14] & g[25450];
assign g[41835] = a[14] & g[25451];
assign g[58218] = b[14] & g[25451];
assign g[41836] = a[14] & g[25452];
assign g[58219] = b[14] & g[25452];
assign g[41837] = a[14] & g[25453];
assign g[58220] = b[14] & g[25453];
assign g[41838] = a[14] & g[25454];
assign g[58221] = b[14] & g[25454];
assign g[41839] = a[14] & g[25455];
assign g[58222] = b[14] & g[25455];
assign g[41840] = a[14] & g[25456];
assign g[58223] = b[14] & g[25456];
assign g[41841] = a[14] & g[25457];
assign g[58224] = b[14] & g[25457];
assign g[41842] = a[14] & g[25458];
assign g[58225] = b[14] & g[25458];
assign g[41843] = a[14] & g[25459];
assign g[58226] = b[14] & g[25459];
assign g[41844] = a[14] & g[25460];
assign g[58227] = b[14] & g[25460];
assign g[41845] = a[14] & g[25461];
assign g[58228] = b[14] & g[25461];
assign g[41846] = a[14] & g[25462];
assign g[58229] = b[14] & g[25462];
assign g[41847] = a[14] & g[25463];
assign g[58230] = b[14] & g[25463];
assign g[41848] = a[14] & g[25464];
assign g[58231] = b[14] & g[25464];
assign g[41849] = a[14] & g[25465];
assign g[58232] = b[14] & g[25465];
assign g[41850] = a[14] & g[25466];
assign g[58233] = b[14] & g[25466];
assign g[41851] = a[14] & g[25467];
assign g[58234] = b[14] & g[25467];
assign g[41852] = a[14] & g[25468];
assign g[58235] = b[14] & g[25468];
assign g[41853] = a[14] & g[25469];
assign g[58236] = b[14] & g[25469];
assign g[41854] = a[14] & g[25470];
assign g[58237] = b[14] & g[25470];
assign g[41855] = a[14] & g[25471];
assign g[58238] = b[14] & g[25471];
assign g[41856] = a[14] & g[25472];
assign g[58239] = b[14] & g[25472];
assign g[41857] = a[14] & g[25473];
assign g[58240] = b[14] & g[25473];
assign g[41858] = a[14] & g[25474];
assign g[58241] = b[14] & g[25474];
assign g[41859] = a[14] & g[25475];
assign g[58242] = b[14] & g[25475];
assign g[41860] = a[14] & g[25476];
assign g[58243] = b[14] & g[25476];
assign g[41861] = a[14] & g[25477];
assign g[58244] = b[14] & g[25477];
assign g[41862] = a[14] & g[25478];
assign g[58245] = b[14] & g[25478];
assign g[41863] = a[14] & g[25479];
assign g[58246] = b[14] & g[25479];
assign g[41864] = a[14] & g[25480];
assign g[58247] = b[14] & g[25480];
assign g[41865] = a[14] & g[25481];
assign g[58248] = b[14] & g[25481];
assign g[41866] = a[14] & g[25482];
assign g[58249] = b[14] & g[25482];
assign g[41867] = a[14] & g[25483];
assign g[58250] = b[14] & g[25483];
assign g[41868] = a[14] & g[25484];
assign g[58251] = b[14] & g[25484];
assign g[41869] = a[14] & g[25485];
assign g[58252] = b[14] & g[25485];
assign g[41870] = a[14] & g[25486];
assign g[58253] = b[14] & g[25486];
assign g[41871] = a[14] & g[25487];
assign g[58254] = b[14] & g[25487];
assign g[41872] = a[14] & g[25488];
assign g[58255] = b[14] & g[25488];
assign g[41873] = a[14] & g[25489];
assign g[58256] = b[14] & g[25489];
assign g[41874] = a[14] & g[25490];
assign g[58257] = b[14] & g[25490];
assign g[41875] = a[14] & g[25491];
assign g[58258] = b[14] & g[25491];
assign g[41876] = a[14] & g[25492];
assign g[58259] = b[14] & g[25492];
assign g[41877] = a[14] & g[25493];
assign g[58260] = b[14] & g[25493];
assign g[41878] = a[14] & g[25494];
assign g[58261] = b[14] & g[25494];
assign g[41879] = a[14] & g[25495];
assign g[58262] = b[14] & g[25495];
assign g[41880] = a[14] & g[25496];
assign g[58263] = b[14] & g[25496];
assign g[41881] = a[14] & g[25497];
assign g[58264] = b[14] & g[25497];
assign g[41882] = a[14] & g[25498];
assign g[58265] = b[14] & g[25498];
assign g[41883] = a[14] & g[25499];
assign g[58266] = b[14] & g[25499];
assign g[41884] = a[14] & g[25500];
assign g[58267] = b[14] & g[25500];
assign g[41885] = a[14] & g[25501];
assign g[58268] = b[14] & g[25501];
assign g[41886] = a[14] & g[25502];
assign g[58269] = b[14] & g[25502];
assign g[41887] = a[14] & g[25503];
assign g[58270] = b[14] & g[25503];
assign g[41888] = a[14] & g[25504];
assign g[58271] = b[14] & g[25504];
assign g[41889] = a[14] & g[25505];
assign g[58272] = b[14] & g[25505];
assign g[41890] = a[14] & g[25506];
assign g[58273] = b[14] & g[25506];
assign g[41891] = a[14] & g[25507];
assign g[58274] = b[14] & g[25507];
assign g[41892] = a[14] & g[25508];
assign g[58275] = b[14] & g[25508];
assign g[41893] = a[14] & g[25509];
assign g[58276] = b[14] & g[25509];
assign g[41894] = a[14] & g[25510];
assign g[58277] = b[14] & g[25510];
assign g[41895] = a[14] & g[25511];
assign g[58278] = b[14] & g[25511];
assign g[41896] = a[14] & g[25512];
assign g[58279] = b[14] & g[25512];
assign g[41897] = a[14] & g[25513];
assign g[58280] = b[14] & g[25513];
assign g[41898] = a[14] & g[25514];
assign g[58281] = b[14] & g[25514];
assign g[41899] = a[14] & g[25515];
assign g[58282] = b[14] & g[25515];
assign g[41900] = a[14] & g[25516];
assign g[58283] = b[14] & g[25516];
assign g[41901] = a[14] & g[25517];
assign g[58284] = b[14] & g[25517];
assign g[41902] = a[14] & g[25518];
assign g[58285] = b[14] & g[25518];
assign g[41903] = a[14] & g[25519];
assign g[58286] = b[14] & g[25519];
assign g[41904] = a[14] & g[25520];
assign g[58287] = b[14] & g[25520];
assign g[41905] = a[14] & g[25521];
assign g[58288] = b[14] & g[25521];
assign g[41906] = a[14] & g[25522];
assign g[58289] = b[14] & g[25522];
assign g[41907] = a[14] & g[25523];
assign g[58290] = b[14] & g[25523];
assign g[41908] = a[14] & g[25524];
assign g[58291] = b[14] & g[25524];
assign g[41909] = a[14] & g[25525];
assign g[58292] = b[14] & g[25525];
assign g[41910] = a[14] & g[25526];
assign g[58293] = b[14] & g[25526];
assign g[41911] = a[14] & g[25527];
assign g[58294] = b[14] & g[25527];
assign g[41912] = a[14] & g[25528];
assign g[58295] = b[14] & g[25528];
assign g[41913] = a[14] & g[25529];
assign g[58296] = b[14] & g[25529];
assign g[41914] = a[14] & g[25530];
assign g[58297] = b[14] & g[25530];
assign g[41915] = a[14] & g[25531];
assign g[58298] = b[14] & g[25531];
assign g[41916] = a[14] & g[25532];
assign g[58299] = b[14] & g[25532];
assign g[41917] = a[14] & g[25533];
assign g[58300] = b[14] & g[25533];
assign g[41918] = a[14] & g[25534];
assign g[58301] = b[14] & g[25534];
assign g[41919] = a[14] & g[25535];
assign g[58302] = b[14] & g[25535];
assign g[41920] = a[14] & g[25536];
assign g[58303] = b[14] & g[25536];
assign g[41921] = a[14] & g[25537];
assign g[58304] = b[14] & g[25537];
assign g[41922] = a[14] & g[25538];
assign g[58305] = b[14] & g[25538];
assign g[41923] = a[14] & g[25539];
assign g[58306] = b[14] & g[25539];
assign g[41924] = a[14] & g[25540];
assign g[58307] = b[14] & g[25540];
assign g[41925] = a[14] & g[25541];
assign g[58308] = b[14] & g[25541];
assign g[41926] = a[14] & g[25542];
assign g[58309] = b[14] & g[25542];
assign g[41927] = a[14] & g[25543];
assign g[58310] = b[14] & g[25543];
assign g[41928] = a[14] & g[25544];
assign g[58311] = b[14] & g[25544];
assign g[41929] = a[14] & g[25545];
assign g[58312] = b[14] & g[25545];
assign g[41930] = a[14] & g[25546];
assign g[58313] = b[14] & g[25546];
assign g[41931] = a[14] & g[25547];
assign g[58314] = b[14] & g[25547];
assign g[41932] = a[14] & g[25548];
assign g[58315] = b[14] & g[25548];
assign g[41933] = a[14] & g[25549];
assign g[58316] = b[14] & g[25549];
assign g[41934] = a[14] & g[25550];
assign g[58317] = b[14] & g[25550];
assign g[41935] = a[14] & g[25551];
assign g[58318] = b[14] & g[25551];
assign g[41936] = a[14] & g[25552];
assign g[58319] = b[14] & g[25552];
assign g[41937] = a[14] & g[25553];
assign g[58320] = b[14] & g[25553];
assign g[41938] = a[14] & g[25554];
assign g[58321] = b[14] & g[25554];
assign g[41939] = a[14] & g[25555];
assign g[58322] = b[14] & g[25555];
assign g[41940] = a[14] & g[25556];
assign g[58323] = b[14] & g[25556];
assign g[41941] = a[14] & g[25557];
assign g[58324] = b[14] & g[25557];
assign g[41942] = a[14] & g[25558];
assign g[58325] = b[14] & g[25558];
assign g[41943] = a[14] & g[25559];
assign g[58326] = b[14] & g[25559];
assign g[41944] = a[14] & g[25560];
assign g[58327] = b[14] & g[25560];
assign g[41945] = a[14] & g[25561];
assign g[58328] = b[14] & g[25561];
assign g[41946] = a[14] & g[25562];
assign g[58329] = b[14] & g[25562];
assign g[41947] = a[14] & g[25563];
assign g[58330] = b[14] & g[25563];
assign g[41948] = a[14] & g[25564];
assign g[58331] = b[14] & g[25564];
assign g[41949] = a[14] & g[25565];
assign g[58332] = b[14] & g[25565];
assign g[41950] = a[14] & g[25566];
assign g[58333] = b[14] & g[25566];
assign g[41951] = a[14] & g[25567];
assign g[58334] = b[14] & g[25567];
assign g[41952] = a[14] & g[25568];
assign g[58335] = b[14] & g[25568];
assign g[41953] = a[14] & g[25569];
assign g[58336] = b[14] & g[25569];
assign g[41954] = a[14] & g[25570];
assign g[58337] = b[14] & g[25570];
assign g[41955] = a[14] & g[25571];
assign g[58338] = b[14] & g[25571];
assign g[41956] = a[14] & g[25572];
assign g[58339] = b[14] & g[25572];
assign g[41957] = a[14] & g[25573];
assign g[58340] = b[14] & g[25573];
assign g[41958] = a[14] & g[25574];
assign g[58341] = b[14] & g[25574];
assign g[41959] = a[14] & g[25575];
assign g[58342] = b[14] & g[25575];
assign g[41960] = a[14] & g[25576];
assign g[58343] = b[14] & g[25576];
assign g[41961] = a[14] & g[25577];
assign g[58344] = b[14] & g[25577];
assign g[41962] = a[14] & g[25578];
assign g[58345] = b[14] & g[25578];
assign g[41963] = a[14] & g[25579];
assign g[58346] = b[14] & g[25579];
assign g[41964] = a[14] & g[25580];
assign g[58347] = b[14] & g[25580];
assign g[41965] = a[14] & g[25581];
assign g[58348] = b[14] & g[25581];
assign g[41966] = a[14] & g[25582];
assign g[58349] = b[14] & g[25582];
assign g[41967] = a[14] & g[25583];
assign g[58350] = b[14] & g[25583];
assign g[41968] = a[14] & g[25584];
assign g[58351] = b[14] & g[25584];
assign g[41969] = a[14] & g[25585];
assign g[58352] = b[14] & g[25585];
assign g[41970] = a[14] & g[25586];
assign g[58353] = b[14] & g[25586];
assign g[41971] = a[14] & g[25587];
assign g[58354] = b[14] & g[25587];
assign g[41972] = a[14] & g[25588];
assign g[58355] = b[14] & g[25588];
assign g[41973] = a[14] & g[25589];
assign g[58356] = b[14] & g[25589];
assign g[41974] = a[14] & g[25590];
assign g[58357] = b[14] & g[25590];
assign g[41975] = a[14] & g[25591];
assign g[58358] = b[14] & g[25591];
assign g[41976] = a[14] & g[25592];
assign g[58359] = b[14] & g[25592];
assign g[41977] = a[14] & g[25593];
assign g[58360] = b[14] & g[25593];
assign g[41978] = a[14] & g[25594];
assign g[58361] = b[14] & g[25594];
assign g[41979] = a[14] & g[25595];
assign g[58362] = b[14] & g[25595];
assign g[41980] = a[14] & g[25596];
assign g[58363] = b[14] & g[25596];
assign g[41981] = a[14] & g[25597];
assign g[58364] = b[14] & g[25597];
assign g[41982] = a[14] & g[25598];
assign g[58365] = b[14] & g[25598];
assign g[41983] = a[14] & g[25599];
assign g[58366] = b[14] & g[25599];
assign g[41984] = a[14] & g[25600];
assign g[58367] = b[14] & g[25600];
assign g[41985] = a[14] & g[25601];
assign g[58368] = b[14] & g[25601];
assign g[41986] = a[14] & g[25602];
assign g[58369] = b[14] & g[25602];
assign g[41987] = a[14] & g[25603];
assign g[58370] = b[14] & g[25603];
assign g[41988] = a[14] & g[25604];
assign g[58371] = b[14] & g[25604];
assign g[41989] = a[14] & g[25605];
assign g[58372] = b[14] & g[25605];
assign g[41990] = a[14] & g[25606];
assign g[58373] = b[14] & g[25606];
assign g[41991] = a[14] & g[25607];
assign g[58374] = b[14] & g[25607];
assign g[41992] = a[14] & g[25608];
assign g[58375] = b[14] & g[25608];
assign g[41993] = a[14] & g[25609];
assign g[58376] = b[14] & g[25609];
assign g[41994] = a[14] & g[25610];
assign g[58377] = b[14] & g[25610];
assign g[41995] = a[14] & g[25611];
assign g[58378] = b[14] & g[25611];
assign g[41996] = a[14] & g[25612];
assign g[58379] = b[14] & g[25612];
assign g[41997] = a[14] & g[25613];
assign g[58380] = b[14] & g[25613];
assign g[41998] = a[14] & g[25614];
assign g[58381] = b[14] & g[25614];
assign g[41999] = a[14] & g[25615];
assign g[58382] = b[14] & g[25615];
assign g[42000] = a[14] & g[25616];
assign g[58383] = b[14] & g[25616];
assign g[42001] = a[14] & g[25617];
assign g[58384] = b[14] & g[25617];
assign g[42002] = a[14] & g[25618];
assign g[58385] = b[14] & g[25618];
assign g[42003] = a[14] & g[25619];
assign g[58386] = b[14] & g[25619];
assign g[42004] = a[14] & g[25620];
assign g[58387] = b[14] & g[25620];
assign g[42005] = a[14] & g[25621];
assign g[58388] = b[14] & g[25621];
assign g[42006] = a[14] & g[25622];
assign g[58389] = b[14] & g[25622];
assign g[42007] = a[14] & g[25623];
assign g[58390] = b[14] & g[25623];
assign g[42008] = a[14] & g[25624];
assign g[58391] = b[14] & g[25624];
assign g[42009] = a[14] & g[25625];
assign g[58392] = b[14] & g[25625];
assign g[42010] = a[14] & g[25626];
assign g[58393] = b[14] & g[25626];
assign g[42011] = a[14] & g[25627];
assign g[58394] = b[14] & g[25627];
assign g[42012] = a[14] & g[25628];
assign g[58395] = b[14] & g[25628];
assign g[42013] = a[14] & g[25629];
assign g[58396] = b[14] & g[25629];
assign g[42014] = a[14] & g[25630];
assign g[58397] = b[14] & g[25630];
assign g[42015] = a[14] & g[25631];
assign g[58398] = b[14] & g[25631];
assign g[42016] = a[14] & g[25632];
assign g[58399] = b[14] & g[25632];
assign g[42017] = a[14] & g[25633];
assign g[58400] = b[14] & g[25633];
assign g[42018] = a[14] & g[25634];
assign g[58401] = b[14] & g[25634];
assign g[42019] = a[14] & g[25635];
assign g[58402] = b[14] & g[25635];
assign g[42020] = a[14] & g[25636];
assign g[58403] = b[14] & g[25636];
assign g[42021] = a[14] & g[25637];
assign g[58404] = b[14] & g[25637];
assign g[42022] = a[14] & g[25638];
assign g[58405] = b[14] & g[25638];
assign g[42023] = a[14] & g[25639];
assign g[58406] = b[14] & g[25639];
assign g[42024] = a[14] & g[25640];
assign g[58407] = b[14] & g[25640];
assign g[42025] = a[14] & g[25641];
assign g[58408] = b[14] & g[25641];
assign g[42026] = a[14] & g[25642];
assign g[58409] = b[14] & g[25642];
assign g[42027] = a[14] & g[25643];
assign g[58410] = b[14] & g[25643];
assign g[42028] = a[14] & g[25644];
assign g[58411] = b[14] & g[25644];
assign g[42029] = a[14] & g[25645];
assign g[58412] = b[14] & g[25645];
assign g[42030] = a[14] & g[25646];
assign g[58413] = b[14] & g[25646];
assign g[42031] = a[14] & g[25647];
assign g[58414] = b[14] & g[25647];
assign g[42032] = a[14] & g[25648];
assign g[58415] = b[14] & g[25648];
assign g[42033] = a[14] & g[25649];
assign g[58416] = b[14] & g[25649];
assign g[42034] = a[14] & g[25650];
assign g[58417] = b[14] & g[25650];
assign g[42035] = a[14] & g[25651];
assign g[58418] = b[14] & g[25651];
assign g[42036] = a[14] & g[25652];
assign g[58419] = b[14] & g[25652];
assign g[42037] = a[14] & g[25653];
assign g[58420] = b[14] & g[25653];
assign g[42038] = a[14] & g[25654];
assign g[58421] = b[14] & g[25654];
assign g[42039] = a[14] & g[25655];
assign g[58422] = b[14] & g[25655];
assign g[42040] = a[14] & g[25656];
assign g[58423] = b[14] & g[25656];
assign g[42041] = a[14] & g[25657];
assign g[58424] = b[14] & g[25657];
assign g[42042] = a[14] & g[25658];
assign g[58425] = b[14] & g[25658];
assign g[42043] = a[14] & g[25659];
assign g[58426] = b[14] & g[25659];
assign g[42044] = a[14] & g[25660];
assign g[58427] = b[14] & g[25660];
assign g[42045] = a[14] & g[25661];
assign g[58428] = b[14] & g[25661];
assign g[42046] = a[14] & g[25662];
assign g[58429] = b[14] & g[25662];
assign g[42047] = a[14] & g[25663];
assign g[58430] = b[14] & g[25663];
assign g[42048] = a[14] & g[25664];
assign g[58431] = b[14] & g[25664];
assign g[42049] = a[14] & g[25665];
assign g[58432] = b[14] & g[25665];
assign g[42050] = a[14] & g[25666];
assign g[58433] = b[14] & g[25666];
assign g[42051] = a[14] & g[25667];
assign g[58434] = b[14] & g[25667];
assign g[42052] = a[14] & g[25668];
assign g[58435] = b[14] & g[25668];
assign g[42053] = a[14] & g[25669];
assign g[58436] = b[14] & g[25669];
assign g[42054] = a[14] & g[25670];
assign g[58437] = b[14] & g[25670];
assign g[42055] = a[14] & g[25671];
assign g[58438] = b[14] & g[25671];
assign g[42056] = a[14] & g[25672];
assign g[58439] = b[14] & g[25672];
assign g[42057] = a[14] & g[25673];
assign g[58440] = b[14] & g[25673];
assign g[42058] = a[14] & g[25674];
assign g[58441] = b[14] & g[25674];
assign g[42059] = a[14] & g[25675];
assign g[58442] = b[14] & g[25675];
assign g[42060] = a[14] & g[25676];
assign g[58443] = b[14] & g[25676];
assign g[42061] = a[14] & g[25677];
assign g[58444] = b[14] & g[25677];
assign g[42062] = a[14] & g[25678];
assign g[58445] = b[14] & g[25678];
assign g[42063] = a[14] & g[25679];
assign g[58446] = b[14] & g[25679];
assign g[42064] = a[14] & g[25680];
assign g[58447] = b[14] & g[25680];
assign g[42065] = a[14] & g[25681];
assign g[58448] = b[14] & g[25681];
assign g[42066] = a[14] & g[25682];
assign g[58449] = b[14] & g[25682];
assign g[42067] = a[14] & g[25683];
assign g[58450] = b[14] & g[25683];
assign g[42068] = a[14] & g[25684];
assign g[58451] = b[14] & g[25684];
assign g[42069] = a[14] & g[25685];
assign g[58452] = b[14] & g[25685];
assign g[42070] = a[14] & g[25686];
assign g[58453] = b[14] & g[25686];
assign g[42071] = a[14] & g[25687];
assign g[58454] = b[14] & g[25687];
assign g[42072] = a[14] & g[25688];
assign g[58455] = b[14] & g[25688];
assign g[42073] = a[14] & g[25689];
assign g[58456] = b[14] & g[25689];
assign g[42074] = a[14] & g[25690];
assign g[58457] = b[14] & g[25690];
assign g[42075] = a[14] & g[25691];
assign g[58458] = b[14] & g[25691];
assign g[42076] = a[14] & g[25692];
assign g[58459] = b[14] & g[25692];
assign g[42077] = a[14] & g[25693];
assign g[58460] = b[14] & g[25693];
assign g[42078] = a[14] & g[25694];
assign g[58461] = b[14] & g[25694];
assign g[42079] = a[14] & g[25695];
assign g[58462] = b[14] & g[25695];
assign g[42080] = a[14] & g[25696];
assign g[58463] = b[14] & g[25696];
assign g[42081] = a[14] & g[25697];
assign g[58464] = b[14] & g[25697];
assign g[42082] = a[14] & g[25698];
assign g[58465] = b[14] & g[25698];
assign g[42083] = a[14] & g[25699];
assign g[58466] = b[14] & g[25699];
assign g[42084] = a[14] & g[25700];
assign g[58467] = b[14] & g[25700];
assign g[42085] = a[14] & g[25701];
assign g[58468] = b[14] & g[25701];
assign g[42086] = a[14] & g[25702];
assign g[58469] = b[14] & g[25702];
assign g[42087] = a[14] & g[25703];
assign g[58470] = b[14] & g[25703];
assign g[42088] = a[14] & g[25704];
assign g[58471] = b[14] & g[25704];
assign g[42089] = a[14] & g[25705];
assign g[58472] = b[14] & g[25705];
assign g[42090] = a[14] & g[25706];
assign g[58473] = b[14] & g[25706];
assign g[42091] = a[14] & g[25707];
assign g[58474] = b[14] & g[25707];
assign g[42092] = a[14] & g[25708];
assign g[58475] = b[14] & g[25708];
assign g[42093] = a[14] & g[25709];
assign g[58476] = b[14] & g[25709];
assign g[42094] = a[14] & g[25710];
assign g[58477] = b[14] & g[25710];
assign g[42095] = a[14] & g[25711];
assign g[58478] = b[14] & g[25711];
assign g[42096] = a[14] & g[25712];
assign g[58479] = b[14] & g[25712];
assign g[42097] = a[14] & g[25713];
assign g[58480] = b[14] & g[25713];
assign g[42098] = a[14] & g[25714];
assign g[58481] = b[14] & g[25714];
assign g[42099] = a[14] & g[25715];
assign g[58482] = b[14] & g[25715];
assign g[42100] = a[14] & g[25716];
assign g[58483] = b[14] & g[25716];
assign g[42101] = a[14] & g[25717];
assign g[58484] = b[14] & g[25717];
assign g[42102] = a[14] & g[25718];
assign g[58485] = b[14] & g[25718];
assign g[42103] = a[14] & g[25719];
assign g[58486] = b[14] & g[25719];
assign g[42104] = a[14] & g[25720];
assign g[58487] = b[14] & g[25720];
assign g[42105] = a[14] & g[25721];
assign g[58488] = b[14] & g[25721];
assign g[42106] = a[14] & g[25722];
assign g[58489] = b[14] & g[25722];
assign g[42107] = a[14] & g[25723];
assign g[58490] = b[14] & g[25723];
assign g[42108] = a[14] & g[25724];
assign g[58491] = b[14] & g[25724];
assign g[42109] = a[14] & g[25725];
assign g[58492] = b[14] & g[25725];
assign g[42110] = a[14] & g[25726];
assign g[58493] = b[14] & g[25726];
assign g[42111] = a[14] & g[25727];
assign g[58494] = b[14] & g[25727];
assign g[42112] = a[14] & g[25728];
assign g[58495] = b[14] & g[25728];
assign g[42113] = a[14] & g[25729];
assign g[58496] = b[14] & g[25729];
assign g[42114] = a[14] & g[25730];
assign g[58497] = b[14] & g[25730];
assign g[42115] = a[14] & g[25731];
assign g[58498] = b[14] & g[25731];
assign g[42116] = a[14] & g[25732];
assign g[58499] = b[14] & g[25732];
assign g[42117] = a[14] & g[25733];
assign g[58500] = b[14] & g[25733];
assign g[42118] = a[14] & g[25734];
assign g[58501] = b[14] & g[25734];
assign g[42119] = a[14] & g[25735];
assign g[58502] = b[14] & g[25735];
assign g[42120] = a[14] & g[25736];
assign g[58503] = b[14] & g[25736];
assign g[42121] = a[14] & g[25737];
assign g[58504] = b[14] & g[25737];
assign g[42122] = a[14] & g[25738];
assign g[58505] = b[14] & g[25738];
assign g[42123] = a[14] & g[25739];
assign g[58506] = b[14] & g[25739];
assign g[42124] = a[14] & g[25740];
assign g[58507] = b[14] & g[25740];
assign g[42125] = a[14] & g[25741];
assign g[58508] = b[14] & g[25741];
assign g[42126] = a[14] & g[25742];
assign g[58509] = b[14] & g[25742];
assign g[42127] = a[14] & g[25743];
assign g[58510] = b[14] & g[25743];
assign g[42128] = a[14] & g[25744];
assign g[58511] = b[14] & g[25744];
assign g[42129] = a[14] & g[25745];
assign g[58512] = b[14] & g[25745];
assign g[42130] = a[14] & g[25746];
assign g[58513] = b[14] & g[25746];
assign g[42131] = a[14] & g[25747];
assign g[58514] = b[14] & g[25747];
assign g[42132] = a[14] & g[25748];
assign g[58515] = b[14] & g[25748];
assign g[42133] = a[14] & g[25749];
assign g[58516] = b[14] & g[25749];
assign g[42134] = a[14] & g[25750];
assign g[58517] = b[14] & g[25750];
assign g[42135] = a[14] & g[25751];
assign g[58518] = b[14] & g[25751];
assign g[42136] = a[14] & g[25752];
assign g[58519] = b[14] & g[25752];
assign g[42137] = a[14] & g[25753];
assign g[58520] = b[14] & g[25753];
assign g[42138] = a[14] & g[25754];
assign g[58521] = b[14] & g[25754];
assign g[42139] = a[14] & g[25755];
assign g[58522] = b[14] & g[25755];
assign g[42140] = a[14] & g[25756];
assign g[58523] = b[14] & g[25756];
assign g[42141] = a[14] & g[25757];
assign g[58524] = b[14] & g[25757];
assign g[42142] = a[14] & g[25758];
assign g[58525] = b[14] & g[25758];
assign g[42143] = a[14] & g[25759];
assign g[58526] = b[14] & g[25759];
assign g[42144] = a[14] & g[25760];
assign g[58527] = b[14] & g[25760];
assign g[42145] = a[14] & g[25761];
assign g[58528] = b[14] & g[25761];
assign g[42146] = a[14] & g[25762];
assign g[58529] = b[14] & g[25762];
assign g[42147] = a[14] & g[25763];
assign g[58530] = b[14] & g[25763];
assign g[42148] = a[14] & g[25764];
assign g[58531] = b[14] & g[25764];
assign g[42149] = a[14] & g[25765];
assign g[58532] = b[14] & g[25765];
assign g[42150] = a[14] & g[25766];
assign g[58533] = b[14] & g[25766];
assign g[42151] = a[14] & g[25767];
assign g[58534] = b[14] & g[25767];
assign g[42152] = a[14] & g[25768];
assign g[58535] = b[14] & g[25768];
assign g[42153] = a[14] & g[25769];
assign g[58536] = b[14] & g[25769];
assign g[42154] = a[14] & g[25770];
assign g[58537] = b[14] & g[25770];
assign g[42155] = a[14] & g[25771];
assign g[58538] = b[14] & g[25771];
assign g[42156] = a[14] & g[25772];
assign g[58539] = b[14] & g[25772];
assign g[42157] = a[14] & g[25773];
assign g[58540] = b[14] & g[25773];
assign g[42158] = a[14] & g[25774];
assign g[58541] = b[14] & g[25774];
assign g[42159] = a[14] & g[25775];
assign g[58542] = b[14] & g[25775];
assign g[42160] = a[14] & g[25776];
assign g[58543] = b[14] & g[25776];
assign g[42161] = a[14] & g[25777];
assign g[58544] = b[14] & g[25777];
assign g[42162] = a[14] & g[25778];
assign g[58545] = b[14] & g[25778];
assign g[42163] = a[14] & g[25779];
assign g[58546] = b[14] & g[25779];
assign g[42164] = a[14] & g[25780];
assign g[58547] = b[14] & g[25780];
assign g[42165] = a[14] & g[25781];
assign g[58548] = b[14] & g[25781];
assign g[42166] = a[14] & g[25782];
assign g[58549] = b[14] & g[25782];
assign g[42167] = a[14] & g[25783];
assign g[58550] = b[14] & g[25783];
assign g[42168] = a[14] & g[25784];
assign g[58551] = b[14] & g[25784];
assign g[42169] = a[14] & g[25785];
assign g[58552] = b[14] & g[25785];
assign g[42170] = a[14] & g[25786];
assign g[58553] = b[14] & g[25786];
assign g[42171] = a[14] & g[25787];
assign g[58554] = b[14] & g[25787];
assign g[42172] = a[14] & g[25788];
assign g[58555] = b[14] & g[25788];
assign g[42173] = a[14] & g[25789];
assign g[58556] = b[14] & g[25789];
assign g[42174] = a[14] & g[25790];
assign g[58557] = b[14] & g[25790];
assign g[42175] = a[14] & g[25791];
assign g[58558] = b[14] & g[25791];
assign g[42176] = a[14] & g[25792];
assign g[58559] = b[14] & g[25792];
assign g[42177] = a[14] & g[25793];
assign g[58560] = b[14] & g[25793];
assign g[42178] = a[14] & g[25794];
assign g[58561] = b[14] & g[25794];
assign g[42179] = a[14] & g[25795];
assign g[58562] = b[14] & g[25795];
assign g[42180] = a[14] & g[25796];
assign g[58563] = b[14] & g[25796];
assign g[42181] = a[14] & g[25797];
assign g[58564] = b[14] & g[25797];
assign g[42182] = a[14] & g[25798];
assign g[58565] = b[14] & g[25798];
assign g[42183] = a[14] & g[25799];
assign g[58566] = b[14] & g[25799];
assign g[42184] = a[14] & g[25800];
assign g[58567] = b[14] & g[25800];
assign g[42185] = a[14] & g[25801];
assign g[58568] = b[14] & g[25801];
assign g[42186] = a[14] & g[25802];
assign g[58569] = b[14] & g[25802];
assign g[42187] = a[14] & g[25803];
assign g[58570] = b[14] & g[25803];
assign g[42188] = a[14] & g[25804];
assign g[58571] = b[14] & g[25804];
assign g[42189] = a[14] & g[25805];
assign g[58572] = b[14] & g[25805];
assign g[42190] = a[14] & g[25806];
assign g[58573] = b[14] & g[25806];
assign g[42191] = a[14] & g[25807];
assign g[58574] = b[14] & g[25807];
assign g[42192] = a[14] & g[25808];
assign g[58575] = b[14] & g[25808];
assign g[42193] = a[14] & g[25809];
assign g[58576] = b[14] & g[25809];
assign g[42194] = a[14] & g[25810];
assign g[58577] = b[14] & g[25810];
assign g[42195] = a[14] & g[25811];
assign g[58578] = b[14] & g[25811];
assign g[42196] = a[14] & g[25812];
assign g[58579] = b[14] & g[25812];
assign g[42197] = a[14] & g[25813];
assign g[58580] = b[14] & g[25813];
assign g[42198] = a[14] & g[25814];
assign g[58581] = b[14] & g[25814];
assign g[42199] = a[14] & g[25815];
assign g[58582] = b[14] & g[25815];
assign g[42200] = a[14] & g[25816];
assign g[58583] = b[14] & g[25816];
assign g[42201] = a[14] & g[25817];
assign g[58584] = b[14] & g[25817];
assign g[42202] = a[14] & g[25818];
assign g[58585] = b[14] & g[25818];
assign g[42203] = a[14] & g[25819];
assign g[58586] = b[14] & g[25819];
assign g[42204] = a[14] & g[25820];
assign g[58587] = b[14] & g[25820];
assign g[42205] = a[14] & g[25821];
assign g[58588] = b[14] & g[25821];
assign g[42206] = a[14] & g[25822];
assign g[58589] = b[14] & g[25822];
assign g[42207] = a[14] & g[25823];
assign g[58590] = b[14] & g[25823];
assign g[42208] = a[14] & g[25824];
assign g[58591] = b[14] & g[25824];
assign g[42209] = a[14] & g[25825];
assign g[58592] = b[14] & g[25825];
assign g[42210] = a[14] & g[25826];
assign g[58593] = b[14] & g[25826];
assign g[42211] = a[14] & g[25827];
assign g[58594] = b[14] & g[25827];
assign g[42212] = a[14] & g[25828];
assign g[58595] = b[14] & g[25828];
assign g[42213] = a[14] & g[25829];
assign g[58596] = b[14] & g[25829];
assign g[42214] = a[14] & g[25830];
assign g[58597] = b[14] & g[25830];
assign g[42215] = a[14] & g[25831];
assign g[58598] = b[14] & g[25831];
assign g[42216] = a[14] & g[25832];
assign g[58599] = b[14] & g[25832];
assign g[42217] = a[14] & g[25833];
assign g[58600] = b[14] & g[25833];
assign g[42218] = a[14] & g[25834];
assign g[58601] = b[14] & g[25834];
assign g[42219] = a[14] & g[25835];
assign g[58602] = b[14] & g[25835];
assign g[42220] = a[14] & g[25836];
assign g[58603] = b[14] & g[25836];
assign g[42221] = a[14] & g[25837];
assign g[58604] = b[14] & g[25837];
assign g[42222] = a[14] & g[25838];
assign g[58605] = b[14] & g[25838];
assign g[42223] = a[14] & g[25839];
assign g[58606] = b[14] & g[25839];
assign g[42224] = a[14] & g[25840];
assign g[58607] = b[14] & g[25840];
assign g[42225] = a[14] & g[25841];
assign g[58608] = b[14] & g[25841];
assign g[42226] = a[14] & g[25842];
assign g[58609] = b[14] & g[25842];
assign g[42227] = a[14] & g[25843];
assign g[58610] = b[14] & g[25843];
assign g[42228] = a[14] & g[25844];
assign g[58611] = b[14] & g[25844];
assign g[42229] = a[14] & g[25845];
assign g[58612] = b[14] & g[25845];
assign g[42230] = a[14] & g[25846];
assign g[58613] = b[14] & g[25846];
assign g[42231] = a[14] & g[25847];
assign g[58614] = b[14] & g[25847];
assign g[42232] = a[14] & g[25848];
assign g[58615] = b[14] & g[25848];
assign g[42233] = a[14] & g[25849];
assign g[58616] = b[14] & g[25849];
assign g[42234] = a[14] & g[25850];
assign g[58617] = b[14] & g[25850];
assign g[42235] = a[14] & g[25851];
assign g[58618] = b[14] & g[25851];
assign g[42236] = a[14] & g[25852];
assign g[58619] = b[14] & g[25852];
assign g[42237] = a[14] & g[25853];
assign g[58620] = b[14] & g[25853];
assign g[42238] = a[14] & g[25854];
assign g[58621] = b[14] & g[25854];
assign g[42239] = a[14] & g[25855];
assign g[58622] = b[14] & g[25855];
assign g[42240] = a[14] & g[25856];
assign g[58623] = b[14] & g[25856];
assign g[42241] = a[14] & g[25857];
assign g[58624] = b[14] & g[25857];
assign g[42242] = a[14] & g[25858];
assign g[58625] = b[14] & g[25858];
assign g[42243] = a[14] & g[25859];
assign g[58626] = b[14] & g[25859];
assign g[42244] = a[14] & g[25860];
assign g[58627] = b[14] & g[25860];
assign g[42245] = a[14] & g[25861];
assign g[58628] = b[14] & g[25861];
assign g[42246] = a[14] & g[25862];
assign g[58629] = b[14] & g[25862];
assign g[42247] = a[14] & g[25863];
assign g[58630] = b[14] & g[25863];
assign g[42248] = a[14] & g[25864];
assign g[58631] = b[14] & g[25864];
assign g[42249] = a[14] & g[25865];
assign g[58632] = b[14] & g[25865];
assign g[42250] = a[14] & g[25866];
assign g[58633] = b[14] & g[25866];
assign g[42251] = a[14] & g[25867];
assign g[58634] = b[14] & g[25867];
assign g[42252] = a[14] & g[25868];
assign g[58635] = b[14] & g[25868];
assign g[42253] = a[14] & g[25869];
assign g[58636] = b[14] & g[25869];
assign g[42254] = a[14] & g[25870];
assign g[58637] = b[14] & g[25870];
assign g[42255] = a[14] & g[25871];
assign g[58638] = b[14] & g[25871];
assign g[42256] = a[14] & g[25872];
assign g[58639] = b[14] & g[25872];
assign g[42257] = a[14] & g[25873];
assign g[58640] = b[14] & g[25873];
assign g[42258] = a[14] & g[25874];
assign g[58641] = b[14] & g[25874];
assign g[42259] = a[14] & g[25875];
assign g[58642] = b[14] & g[25875];
assign g[42260] = a[14] & g[25876];
assign g[58643] = b[14] & g[25876];
assign g[42261] = a[14] & g[25877];
assign g[58644] = b[14] & g[25877];
assign g[42262] = a[14] & g[25878];
assign g[58645] = b[14] & g[25878];
assign g[42263] = a[14] & g[25879];
assign g[58646] = b[14] & g[25879];
assign g[42264] = a[14] & g[25880];
assign g[58647] = b[14] & g[25880];
assign g[42265] = a[14] & g[25881];
assign g[58648] = b[14] & g[25881];
assign g[42266] = a[14] & g[25882];
assign g[58649] = b[14] & g[25882];
assign g[42267] = a[14] & g[25883];
assign g[58650] = b[14] & g[25883];
assign g[42268] = a[14] & g[25884];
assign g[58651] = b[14] & g[25884];
assign g[42269] = a[14] & g[25885];
assign g[58652] = b[14] & g[25885];
assign g[42270] = a[14] & g[25886];
assign g[58653] = b[14] & g[25886];
assign g[42271] = a[14] & g[25887];
assign g[58654] = b[14] & g[25887];
assign g[42272] = a[14] & g[25888];
assign g[58655] = b[14] & g[25888];
assign g[42273] = a[14] & g[25889];
assign g[58656] = b[14] & g[25889];
assign g[42274] = a[14] & g[25890];
assign g[58657] = b[14] & g[25890];
assign g[42275] = a[14] & g[25891];
assign g[58658] = b[14] & g[25891];
assign g[42276] = a[14] & g[25892];
assign g[58659] = b[14] & g[25892];
assign g[42277] = a[14] & g[25893];
assign g[58660] = b[14] & g[25893];
assign g[42278] = a[14] & g[25894];
assign g[58661] = b[14] & g[25894];
assign g[42279] = a[14] & g[25895];
assign g[58662] = b[14] & g[25895];
assign g[42280] = a[14] & g[25896];
assign g[58663] = b[14] & g[25896];
assign g[42281] = a[14] & g[25897];
assign g[58664] = b[14] & g[25897];
assign g[42282] = a[14] & g[25898];
assign g[58665] = b[14] & g[25898];
assign g[42283] = a[14] & g[25899];
assign g[58666] = b[14] & g[25899];
assign g[42284] = a[14] & g[25900];
assign g[58667] = b[14] & g[25900];
assign g[42285] = a[14] & g[25901];
assign g[58668] = b[14] & g[25901];
assign g[42286] = a[14] & g[25902];
assign g[58669] = b[14] & g[25902];
assign g[42287] = a[14] & g[25903];
assign g[58670] = b[14] & g[25903];
assign g[42288] = a[14] & g[25904];
assign g[58671] = b[14] & g[25904];
assign g[42289] = a[14] & g[25905];
assign g[58672] = b[14] & g[25905];
assign g[42290] = a[14] & g[25906];
assign g[58673] = b[14] & g[25906];
assign g[42291] = a[14] & g[25907];
assign g[58674] = b[14] & g[25907];
assign g[42292] = a[14] & g[25908];
assign g[58675] = b[14] & g[25908];
assign g[42293] = a[14] & g[25909];
assign g[58676] = b[14] & g[25909];
assign g[42294] = a[14] & g[25910];
assign g[58677] = b[14] & g[25910];
assign g[42295] = a[14] & g[25911];
assign g[58678] = b[14] & g[25911];
assign g[42296] = a[14] & g[25912];
assign g[58679] = b[14] & g[25912];
assign g[42297] = a[14] & g[25913];
assign g[58680] = b[14] & g[25913];
assign g[42298] = a[14] & g[25914];
assign g[58681] = b[14] & g[25914];
assign g[42299] = a[14] & g[25915];
assign g[58682] = b[14] & g[25915];
assign g[42300] = a[14] & g[25916];
assign g[58683] = b[14] & g[25916];
assign g[42301] = a[14] & g[25917];
assign g[58684] = b[14] & g[25917];
assign g[42302] = a[14] & g[25918];
assign g[58685] = b[14] & g[25918];
assign g[42303] = a[14] & g[25919];
assign g[58686] = b[14] & g[25919];
assign g[42304] = a[14] & g[25920];
assign g[58687] = b[14] & g[25920];
assign g[42305] = a[14] & g[25921];
assign g[58688] = b[14] & g[25921];
assign g[42306] = a[14] & g[25922];
assign g[58689] = b[14] & g[25922];
assign g[42307] = a[14] & g[25923];
assign g[58690] = b[14] & g[25923];
assign g[42308] = a[14] & g[25924];
assign g[58691] = b[14] & g[25924];
assign g[42309] = a[14] & g[25925];
assign g[58692] = b[14] & g[25925];
assign g[42310] = a[14] & g[25926];
assign g[58693] = b[14] & g[25926];
assign g[42311] = a[14] & g[25927];
assign g[58694] = b[14] & g[25927];
assign g[42312] = a[14] & g[25928];
assign g[58695] = b[14] & g[25928];
assign g[42313] = a[14] & g[25929];
assign g[58696] = b[14] & g[25929];
assign g[42314] = a[14] & g[25930];
assign g[58697] = b[14] & g[25930];
assign g[42315] = a[14] & g[25931];
assign g[58698] = b[14] & g[25931];
assign g[42316] = a[14] & g[25932];
assign g[58699] = b[14] & g[25932];
assign g[42317] = a[14] & g[25933];
assign g[58700] = b[14] & g[25933];
assign g[42318] = a[14] & g[25934];
assign g[58701] = b[14] & g[25934];
assign g[42319] = a[14] & g[25935];
assign g[58702] = b[14] & g[25935];
assign g[42320] = a[14] & g[25936];
assign g[58703] = b[14] & g[25936];
assign g[42321] = a[14] & g[25937];
assign g[58704] = b[14] & g[25937];
assign g[42322] = a[14] & g[25938];
assign g[58705] = b[14] & g[25938];
assign g[42323] = a[14] & g[25939];
assign g[58706] = b[14] & g[25939];
assign g[42324] = a[14] & g[25940];
assign g[58707] = b[14] & g[25940];
assign g[42325] = a[14] & g[25941];
assign g[58708] = b[14] & g[25941];
assign g[42326] = a[14] & g[25942];
assign g[58709] = b[14] & g[25942];
assign g[42327] = a[14] & g[25943];
assign g[58710] = b[14] & g[25943];
assign g[42328] = a[14] & g[25944];
assign g[58711] = b[14] & g[25944];
assign g[42329] = a[14] & g[25945];
assign g[58712] = b[14] & g[25945];
assign g[42330] = a[14] & g[25946];
assign g[58713] = b[14] & g[25946];
assign g[42331] = a[14] & g[25947];
assign g[58714] = b[14] & g[25947];
assign g[42332] = a[14] & g[25948];
assign g[58715] = b[14] & g[25948];
assign g[42333] = a[14] & g[25949];
assign g[58716] = b[14] & g[25949];
assign g[42334] = a[14] & g[25950];
assign g[58717] = b[14] & g[25950];
assign g[42335] = a[14] & g[25951];
assign g[58718] = b[14] & g[25951];
assign g[42336] = a[14] & g[25952];
assign g[58719] = b[14] & g[25952];
assign g[42337] = a[14] & g[25953];
assign g[58720] = b[14] & g[25953];
assign g[42338] = a[14] & g[25954];
assign g[58721] = b[14] & g[25954];
assign g[42339] = a[14] & g[25955];
assign g[58722] = b[14] & g[25955];
assign g[42340] = a[14] & g[25956];
assign g[58723] = b[14] & g[25956];
assign g[42341] = a[14] & g[25957];
assign g[58724] = b[14] & g[25957];
assign g[42342] = a[14] & g[25958];
assign g[58725] = b[14] & g[25958];
assign g[42343] = a[14] & g[25959];
assign g[58726] = b[14] & g[25959];
assign g[42344] = a[14] & g[25960];
assign g[58727] = b[14] & g[25960];
assign g[42345] = a[14] & g[25961];
assign g[58728] = b[14] & g[25961];
assign g[42346] = a[14] & g[25962];
assign g[58729] = b[14] & g[25962];
assign g[42347] = a[14] & g[25963];
assign g[58730] = b[14] & g[25963];
assign g[42348] = a[14] & g[25964];
assign g[58731] = b[14] & g[25964];
assign g[42349] = a[14] & g[25965];
assign g[58732] = b[14] & g[25965];
assign g[42350] = a[14] & g[25966];
assign g[58733] = b[14] & g[25966];
assign g[42351] = a[14] & g[25967];
assign g[58734] = b[14] & g[25967];
assign g[42352] = a[14] & g[25968];
assign g[58735] = b[14] & g[25968];
assign g[42353] = a[14] & g[25969];
assign g[58736] = b[14] & g[25969];
assign g[42354] = a[14] & g[25970];
assign g[58737] = b[14] & g[25970];
assign g[42355] = a[14] & g[25971];
assign g[58738] = b[14] & g[25971];
assign g[42356] = a[14] & g[25972];
assign g[58739] = b[14] & g[25972];
assign g[42357] = a[14] & g[25973];
assign g[58740] = b[14] & g[25973];
assign g[42358] = a[14] & g[25974];
assign g[58741] = b[14] & g[25974];
assign g[42359] = a[14] & g[25975];
assign g[58742] = b[14] & g[25975];
assign g[42360] = a[14] & g[25976];
assign g[58743] = b[14] & g[25976];
assign g[42361] = a[14] & g[25977];
assign g[58744] = b[14] & g[25977];
assign g[42362] = a[14] & g[25978];
assign g[58745] = b[14] & g[25978];
assign g[42363] = a[14] & g[25979];
assign g[58746] = b[14] & g[25979];
assign g[42364] = a[14] & g[25980];
assign g[58747] = b[14] & g[25980];
assign g[42365] = a[14] & g[25981];
assign g[58748] = b[14] & g[25981];
assign g[42366] = a[14] & g[25982];
assign g[58749] = b[14] & g[25982];
assign g[42367] = a[14] & g[25983];
assign g[58750] = b[14] & g[25983];
assign g[42368] = a[14] & g[25984];
assign g[58751] = b[14] & g[25984];
assign g[42369] = a[14] & g[25985];
assign g[58752] = b[14] & g[25985];
assign g[42370] = a[14] & g[25986];
assign g[58753] = b[14] & g[25986];
assign g[42371] = a[14] & g[25987];
assign g[58754] = b[14] & g[25987];
assign g[42372] = a[14] & g[25988];
assign g[58755] = b[14] & g[25988];
assign g[42373] = a[14] & g[25989];
assign g[58756] = b[14] & g[25989];
assign g[42374] = a[14] & g[25990];
assign g[58757] = b[14] & g[25990];
assign g[42375] = a[14] & g[25991];
assign g[58758] = b[14] & g[25991];
assign g[42376] = a[14] & g[25992];
assign g[58759] = b[14] & g[25992];
assign g[42377] = a[14] & g[25993];
assign g[58760] = b[14] & g[25993];
assign g[42378] = a[14] & g[25994];
assign g[58761] = b[14] & g[25994];
assign g[42379] = a[14] & g[25995];
assign g[58762] = b[14] & g[25995];
assign g[42380] = a[14] & g[25996];
assign g[58763] = b[14] & g[25996];
assign g[42381] = a[14] & g[25997];
assign g[58764] = b[14] & g[25997];
assign g[42382] = a[14] & g[25998];
assign g[58765] = b[14] & g[25998];
assign g[42383] = a[14] & g[25999];
assign g[58766] = b[14] & g[25999];
assign g[42384] = a[14] & g[26000];
assign g[58767] = b[14] & g[26000];
assign g[42385] = a[14] & g[26001];
assign g[58768] = b[14] & g[26001];
assign g[42386] = a[14] & g[26002];
assign g[58769] = b[14] & g[26002];
assign g[42387] = a[14] & g[26003];
assign g[58770] = b[14] & g[26003];
assign g[42388] = a[14] & g[26004];
assign g[58771] = b[14] & g[26004];
assign g[42389] = a[14] & g[26005];
assign g[58772] = b[14] & g[26005];
assign g[42390] = a[14] & g[26006];
assign g[58773] = b[14] & g[26006];
assign g[42391] = a[14] & g[26007];
assign g[58774] = b[14] & g[26007];
assign g[42392] = a[14] & g[26008];
assign g[58775] = b[14] & g[26008];
assign g[42393] = a[14] & g[26009];
assign g[58776] = b[14] & g[26009];
assign g[42394] = a[14] & g[26010];
assign g[58777] = b[14] & g[26010];
assign g[42395] = a[14] & g[26011];
assign g[58778] = b[14] & g[26011];
assign g[42396] = a[14] & g[26012];
assign g[58779] = b[14] & g[26012];
assign g[42397] = a[14] & g[26013];
assign g[58780] = b[14] & g[26013];
assign g[42398] = a[14] & g[26014];
assign g[58781] = b[14] & g[26014];
assign g[42399] = a[14] & g[26015];
assign g[58782] = b[14] & g[26015];
assign g[42400] = a[14] & g[26016];
assign g[58783] = b[14] & g[26016];
assign g[42401] = a[14] & g[26017];
assign g[58784] = b[14] & g[26017];
assign g[42402] = a[14] & g[26018];
assign g[58785] = b[14] & g[26018];
assign g[42403] = a[14] & g[26019];
assign g[58786] = b[14] & g[26019];
assign g[42404] = a[14] & g[26020];
assign g[58787] = b[14] & g[26020];
assign g[42405] = a[14] & g[26021];
assign g[58788] = b[14] & g[26021];
assign g[42406] = a[14] & g[26022];
assign g[58789] = b[14] & g[26022];
assign g[42407] = a[14] & g[26023];
assign g[58790] = b[14] & g[26023];
assign g[42408] = a[14] & g[26024];
assign g[58791] = b[14] & g[26024];
assign g[42409] = a[14] & g[26025];
assign g[58792] = b[14] & g[26025];
assign g[42410] = a[14] & g[26026];
assign g[58793] = b[14] & g[26026];
assign g[42411] = a[14] & g[26027];
assign g[58794] = b[14] & g[26027];
assign g[42412] = a[14] & g[26028];
assign g[58795] = b[14] & g[26028];
assign g[42413] = a[14] & g[26029];
assign g[58796] = b[14] & g[26029];
assign g[42414] = a[14] & g[26030];
assign g[58797] = b[14] & g[26030];
assign g[42415] = a[14] & g[26031];
assign g[58798] = b[14] & g[26031];
assign g[42416] = a[14] & g[26032];
assign g[58799] = b[14] & g[26032];
assign g[42417] = a[14] & g[26033];
assign g[58800] = b[14] & g[26033];
assign g[42418] = a[14] & g[26034];
assign g[58801] = b[14] & g[26034];
assign g[42419] = a[14] & g[26035];
assign g[58802] = b[14] & g[26035];
assign g[42420] = a[14] & g[26036];
assign g[58803] = b[14] & g[26036];
assign g[42421] = a[14] & g[26037];
assign g[58804] = b[14] & g[26037];
assign g[42422] = a[14] & g[26038];
assign g[58805] = b[14] & g[26038];
assign g[42423] = a[14] & g[26039];
assign g[58806] = b[14] & g[26039];
assign g[42424] = a[14] & g[26040];
assign g[58807] = b[14] & g[26040];
assign g[42425] = a[14] & g[26041];
assign g[58808] = b[14] & g[26041];
assign g[42426] = a[14] & g[26042];
assign g[58809] = b[14] & g[26042];
assign g[42427] = a[14] & g[26043];
assign g[58810] = b[14] & g[26043];
assign g[42428] = a[14] & g[26044];
assign g[58811] = b[14] & g[26044];
assign g[42429] = a[14] & g[26045];
assign g[58812] = b[14] & g[26045];
assign g[42430] = a[14] & g[26046];
assign g[58813] = b[14] & g[26046];
assign g[42431] = a[14] & g[26047];
assign g[58814] = b[14] & g[26047];
assign g[42432] = a[14] & g[26048];
assign g[58815] = b[14] & g[26048];
assign g[42433] = a[14] & g[26049];
assign g[58816] = b[14] & g[26049];
assign g[42434] = a[14] & g[26050];
assign g[58817] = b[14] & g[26050];
assign g[42435] = a[14] & g[26051];
assign g[58818] = b[14] & g[26051];
assign g[42436] = a[14] & g[26052];
assign g[58819] = b[14] & g[26052];
assign g[42437] = a[14] & g[26053];
assign g[58820] = b[14] & g[26053];
assign g[42438] = a[14] & g[26054];
assign g[58821] = b[14] & g[26054];
assign g[42439] = a[14] & g[26055];
assign g[58822] = b[14] & g[26055];
assign g[42440] = a[14] & g[26056];
assign g[58823] = b[14] & g[26056];
assign g[42441] = a[14] & g[26057];
assign g[58824] = b[14] & g[26057];
assign g[42442] = a[14] & g[26058];
assign g[58825] = b[14] & g[26058];
assign g[42443] = a[14] & g[26059];
assign g[58826] = b[14] & g[26059];
assign g[42444] = a[14] & g[26060];
assign g[58827] = b[14] & g[26060];
assign g[42445] = a[14] & g[26061];
assign g[58828] = b[14] & g[26061];
assign g[42446] = a[14] & g[26062];
assign g[58829] = b[14] & g[26062];
assign g[42447] = a[14] & g[26063];
assign g[58830] = b[14] & g[26063];
assign g[42448] = a[14] & g[26064];
assign g[58831] = b[14] & g[26064];
assign g[42449] = a[14] & g[26065];
assign g[58832] = b[14] & g[26065];
assign g[42450] = a[14] & g[26066];
assign g[58833] = b[14] & g[26066];
assign g[42451] = a[14] & g[26067];
assign g[58834] = b[14] & g[26067];
assign g[42452] = a[14] & g[26068];
assign g[58835] = b[14] & g[26068];
assign g[42453] = a[14] & g[26069];
assign g[58836] = b[14] & g[26069];
assign g[42454] = a[14] & g[26070];
assign g[58837] = b[14] & g[26070];
assign g[42455] = a[14] & g[26071];
assign g[58838] = b[14] & g[26071];
assign g[42456] = a[14] & g[26072];
assign g[58839] = b[14] & g[26072];
assign g[42457] = a[14] & g[26073];
assign g[58840] = b[14] & g[26073];
assign g[42458] = a[14] & g[26074];
assign g[58841] = b[14] & g[26074];
assign g[42459] = a[14] & g[26075];
assign g[58842] = b[14] & g[26075];
assign g[42460] = a[14] & g[26076];
assign g[58843] = b[14] & g[26076];
assign g[42461] = a[14] & g[26077];
assign g[58844] = b[14] & g[26077];
assign g[42462] = a[14] & g[26078];
assign g[58845] = b[14] & g[26078];
assign g[42463] = a[14] & g[26079];
assign g[58846] = b[14] & g[26079];
assign g[42464] = a[14] & g[26080];
assign g[58847] = b[14] & g[26080];
assign g[42465] = a[14] & g[26081];
assign g[58848] = b[14] & g[26081];
assign g[42466] = a[14] & g[26082];
assign g[58849] = b[14] & g[26082];
assign g[42467] = a[14] & g[26083];
assign g[58850] = b[14] & g[26083];
assign g[42468] = a[14] & g[26084];
assign g[58851] = b[14] & g[26084];
assign g[42469] = a[14] & g[26085];
assign g[58852] = b[14] & g[26085];
assign g[42470] = a[14] & g[26086];
assign g[58853] = b[14] & g[26086];
assign g[42471] = a[14] & g[26087];
assign g[58854] = b[14] & g[26087];
assign g[42472] = a[14] & g[26088];
assign g[58855] = b[14] & g[26088];
assign g[42473] = a[14] & g[26089];
assign g[58856] = b[14] & g[26089];
assign g[42474] = a[14] & g[26090];
assign g[58857] = b[14] & g[26090];
assign g[42475] = a[14] & g[26091];
assign g[58858] = b[14] & g[26091];
assign g[42476] = a[14] & g[26092];
assign g[58859] = b[14] & g[26092];
assign g[42477] = a[14] & g[26093];
assign g[58860] = b[14] & g[26093];
assign g[42478] = a[14] & g[26094];
assign g[58861] = b[14] & g[26094];
assign g[42479] = a[14] & g[26095];
assign g[58862] = b[14] & g[26095];
assign g[42480] = a[14] & g[26096];
assign g[58863] = b[14] & g[26096];
assign g[42481] = a[14] & g[26097];
assign g[58864] = b[14] & g[26097];
assign g[42482] = a[14] & g[26098];
assign g[58865] = b[14] & g[26098];
assign g[42483] = a[14] & g[26099];
assign g[58866] = b[14] & g[26099];
assign g[42484] = a[14] & g[26100];
assign g[58867] = b[14] & g[26100];
assign g[42485] = a[14] & g[26101];
assign g[58868] = b[14] & g[26101];
assign g[42486] = a[14] & g[26102];
assign g[58869] = b[14] & g[26102];
assign g[42487] = a[14] & g[26103];
assign g[58870] = b[14] & g[26103];
assign g[42488] = a[14] & g[26104];
assign g[58871] = b[14] & g[26104];
assign g[42489] = a[14] & g[26105];
assign g[58872] = b[14] & g[26105];
assign g[42490] = a[14] & g[26106];
assign g[58873] = b[14] & g[26106];
assign g[42491] = a[14] & g[26107];
assign g[58874] = b[14] & g[26107];
assign g[42492] = a[14] & g[26108];
assign g[58875] = b[14] & g[26108];
assign g[42493] = a[14] & g[26109];
assign g[58876] = b[14] & g[26109];
assign g[42494] = a[14] & g[26110];
assign g[58877] = b[14] & g[26110];
assign g[42495] = a[14] & g[26111];
assign g[58878] = b[14] & g[26111];
assign g[42496] = a[14] & g[26112];
assign g[58879] = b[14] & g[26112];
assign g[42497] = a[14] & g[26113];
assign g[58880] = b[14] & g[26113];
assign g[42498] = a[14] & g[26114];
assign g[58881] = b[14] & g[26114];
assign g[42499] = a[14] & g[26115];
assign g[58882] = b[14] & g[26115];
assign g[42500] = a[14] & g[26116];
assign g[58883] = b[14] & g[26116];
assign g[42501] = a[14] & g[26117];
assign g[58884] = b[14] & g[26117];
assign g[42502] = a[14] & g[26118];
assign g[58885] = b[14] & g[26118];
assign g[42503] = a[14] & g[26119];
assign g[58886] = b[14] & g[26119];
assign g[42504] = a[14] & g[26120];
assign g[58887] = b[14] & g[26120];
assign g[42505] = a[14] & g[26121];
assign g[58888] = b[14] & g[26121];
assign g[42506] = a[14] & g[26122];
assign g[58889] = b[14] & g[26122];
assign g[42507] = a[14] & g[26123];
assign g[58890] = b[14] & g[26123];
assign g[42508] = a[14] & g[26124];
assign g[58891] = b[14] & g[26124];
assign g[42509] = a[14] & g[26125];
assign g[58892] = b[14] & g[26125];
assign g[42510] = a[14] & g[26126];
assign g[58893] = b[14] & g[26126];
assign g[42511] = a[14] & g[26127];
assign g[58894] = b[14] & g[26127];
assign g[42512] = a[14] & g[26128];
assign g[58895] = b[14] & g[26128];
assign g[42513] = a[14] & g[26129];
assign g[58896] = b[14] & g[26129];
assign g[42514] = a[14] & g[26130];
assign g[58897] = b[14] & g[26130];
assign g[42515] = a[14] & g[26131];
assign g[58898] = b[14] & g[26131];
assign g[42516] = a[14] & g[26132];
assign g[58899] = b[14] & g[26132];
assign g[42517] = a[14] & g[26133];
assign g[58900] = b[14] & g[26133];
assign g[42518] = a[14] & g[26134];
assign g[58901] = b[14] & g[26134];
assign g[42519] = a[14] & g[26135];
assign g[58902] = b[14] & g[26135];
assign g[42520] = a[14] & g[26136];
assign g[58903] = b[14] & g[26136];
assign g[42521] = a[14] & g[26137];
assign g[58904] = b[14] & g[26137];
assign g[42522] = a[14] & g[26138];
assign g[58905] = b[14] & g[26138];
assign g[42523] = a[14] & g[26139];
assign g[58906] = b[14] & g[26139];
assign g[42524] = a[14] & g[26140];
assign g[58907] = b[14] & g[26140];
assign g[42525] = a[14] & g[26141];
assign g[58908] = b[14] & g[26141];
assign g[42526] = a[14] & g[26142];
assign g[58909] = b[14] & g[26142];
assign g[42527] = a[14] & g[26143];
assign g[58910] = b[14] & g[26143];
assign g[42528] = a[14] & g[26144];
assign g[58911] = b[14] & g[26144];
assign g[42529] = a[14] & g[26145];
assign g[58912] = b[14] & g[26145];
assign g[42530] = a[14] & g[26146];
assign g[58913] = b[14] & g[26146];
assign g[42531] = a[14] & g[26147];
assign g[58914] = b[14] & g[26147];
assign g[42532] = a[14] & g[26148];
assign g[58915] = b[14] & g[26148];
assign g[42533] = a[14] & g[26149];
assign g[58916] = b[14] & g[26149];
assign g[42534] = a[14] & g[26150];
assign g[58917] = b[14] & g[26150];
assign g[42535] = a[14] & g[26151];
assign g[58918] = b[14] & g[26151];
assign g[42536] = a[14] & g[26152];
assign g[58919] = b[14] & g[26152];
assign g[42537] = a[14] & g[26153];
assign g[58920] = b[14] & g[26153];
assign g[42538] = a[14] & g[26154];
assign g[58921] = b[14] & g[26154];
assign g[42539] = a[14] & g[26155];
assign g[58922] = b[14] & g[26155];
assign g[42540] = a[14] & g[26156];
assign g[58923] = b[14] & g[26156];
assign g[42541] = a[14] & g[26157];
assign g[58924] = b[14] & g[26157];
assign g[42542] = a[14] & g[26158];
assign g[58925] = b[14] & g[26158];
assign g[42543] = a[14] & g[26159];
assign g[58926] = b[14] & g[26159];
assign g[42544] = a[14] & g[26160];
assign g[58927] = b[14] & g[26160];
assign g[42545] = a[14] & g[26161];
assign g[58928] = b[14] & g[26161];
assign g[42546] = a[14] & g[26162];
assign g[58929] = b[14] & g[26162];
assign g[42547] = a[14] & g[26163];
assign g[58930] = b[14] & g[26163];
assign g[42548] = a[14] & g[26164];
assign g[58931] = b[14] & g[26164];
assign g[42549] = a[14] & g[26165];
assign g[58932] = b[14] & g[26165];
assign g[42550] = a[14] & g[26166];
assign g[58933] = b[14] & g[26166];
assign g[42551] = a[14] & g[26167];
assign g[58934] = b[14] & g[26167];
assign g[42552] = a[14] & g[26168];
assign g[58935] = b[14] & g[26168];
assign g[42553] = a[14] & g[26169];
assign g[58936] = b[14] & g[26169];
assign g[42554] = a[14] & g[26170];
assign g[58937] = b[14] & g[26170];
assign g[42555] = a[14] & g[26171];
assign g[58938] = b[14] & g[26171];
assign g[42556] = a[14] & g[26172];
assign g[58939] = b[14] & g[26172];
assign g[42557] = a[14] & g[26173];
assign g[58940] = b[14] & g[26173];
assign g[42558] = a[14] & g[26174];
assign g[58941] = b[14] & g[26174];
assign g[42559] = a[14] & g[26175];
assign g[58942] = b[14] & g[26175];
assign g[42560] = a[14] & g[26176];
assign g[58943] = b[14] & g[26176];
assign g[42561] = a[14] & g[26177];
assign g[58944] = b[14] & g[26177];
assign g[42562] = a[14] & g[26178];
assign g[58945] = b[14] & g[26178];
assign g[42563] = a[14] & g[26179];
assign g[58946] = b[14] & g[26179];
assign g[42564] = a[14] & g[26180];
assign g[58947] = b[14] & g[26180];
assign g[42565] = a[14] & g[26181];
assign g[58948] = b[14] & g[26181];
assign g[42566] = a[14] & g[26182];
assign g[58949] = b[14] & g[26182];
assign g[42567] = a[14] & g[26183];
assign g[58950] = b[14] & g[26183];
assign g[42568] = a[14] & g[26184];
assign g[58951] = b[14] & g[26184];
assign g[42569] = a[14] & g[26185];
assign g[58952] = b[14] & g[26185];
assign g[42570] = a[14] & g[26186];
assign g[58953] = b[14] & g[26186];
assign g[42571] = a[14] & g[26187];
assign g[58954] = b[14] & g[26187];
assign g[42572] = a[14] & g[26188];
assign g[58955] = b[14] & g[26188];
assign g[42573] = a[14] & g[26189];
assign g[58956] = b[14] & g[26189];
assign g[42574] = a[14] & g[26190];
assign g[58957] = b[14] & g[26190];
assign g[42575] = a[14] & g[26191];
assign g[58958] = b[14] & g[26191];
assign g[42576] = a[14] & g[26192];
assign g[58959] = b[14] & g[26192];
assign g[42577] = a[14] & g[26193];
assign g[58960] = b[14] & g[26193];
assign g[42578] = a[14] & g[26194];
assign g[58961] = b[14] & g[26194];
assign g[42579] = a[14] & g[26195];
assign g[58962] = b[14] & g[26195];
assign g[42580] = a[14] & g[26196];
assign g[58963] = b[14] & g[26196];
assign g[42581] = a[14] & g[26197];
assign g[58964] = b[14] & g[26197];
assign g[42582] = a[14] & g[26198];
assign g[58965] = b[14] & g[26198];
assign g[42583] = a[14] & g[26199];
assign g[58966] = b[14] & g[26199];
assign g[42584] = a[14] & g[26200];
assign g[58967] = b[14] & g[26200];
assign g[42585] = a[14] & g[26201];
assign g[58968] = b[14] & g[26201];
assign g[42586] = a[14] & g[26202];
assign g[58969] = b[14] & g[26202];
assign g[42587] = a[14] & g[26203];
assign g[58970] = b[14] & g[26203];
assign g[42588] = a[14] & g[26204];
assign g[58971] = b[14] & g[26204];
assign g[42589] = a[14] & g[26205];
assign g[58972] = b[14] & g[26205];
assign g[42590] = a[14] & g[26206];
assign g[58973] = b[14] & g[26206];
assign g[42591] = a[14] & g[26207];
assign g[58974] = b[14] & g[26207];
assign g[42592] = a[14] & g[26208];
assign g[58975] = b[14] & g[26208];
assign g[42593] = a[14] & g[26209];
assign g[58976] = b[14] & g[26209];
assign g[42594] = a[14] & g[26210];
assign g[58977] = b[14] & g[26210];
assign g[42595] = a[14] & g[26211];
assign g[58978] = b[14] & g[26211];
assign g[42596] = a[14] & g[26212];
assign g[58979] = b[14] & g[26212];
assign g[42597] = a[14] & g[26213];
assign g[58980] = b[14] & g[26213];
assign g[42598] = a[14] & g[26214];
assign g[58981] = b[14] & g[26214];
assign g[42599] = a[14] & g[26215];
assign g[58982] = b[14] & g[26215];
assign g[42600] = a[14] & g[26216];
assign g[58983] = b[14] & g[26216];
assign g[42601] = a[14] & g[26217];
assign g[58984] = b[14] & g[26217];
assign g[42602] = a[14] & g[26218];
assign g[58985] = b[14] & g[26218];
assign g[42603] = a[14] & g[26219];
assign g[58986] = b[14] & g[26219];
assign g[42604] = a[14] & g[26220];
assign g[58987] = b[14] & g[26220];
assign g[42605] = a[14] & g[26221];
assign g[58988] = b[14] & g[26221];
assign g[42606] = a[14] & g[26222];
assign g[58989] = b[14] & g[26222];
assign g[42607] = a[14] & g[26223];
assign g[58990] = b[14] & g[26223];
assign g[42608] = a[14] & g[26224];
assign g[58991] = b[14] & g[26224];
assign g[42609] = a[14] & g[26225];
assign g[58992] = b[14] & g[26225];
assign g[42610] = a[14] & g[26226];
assign g[58993] = b[14] & g[26226];
assign g[42611] = a[14] & g[26227];
assign g[58994] = b[14] & g[26227];
assign g[42612] = a[14] & g[26228];
assign g[58995] = b[14] & g[26228];
assign g[42613] = a[14] & g[26229];
assign g[58996] = b[14] & g[26229];
assign g[42614] = a[14] & g[26230];
assign g[58997] = b[14] & g[26230];
assign g[42615] = a[14] & g[26231];
assign g[58998] = b[14] & g[26231];
assign g[42616] = a[14] & g[26232];
assign g[58999] = b[14] & g[26232];
assign g[42617] = a[14] & g[26233];
assign g[59000] = b[14] & g[26233];
assign g[42618] = a[14] & g[26234];
assign g[59001] = b[14] & g[26234];
assign g[42619] = a[14] & g[26235];
assign g[59002] = b[14] & g[26235];
assign g[42620] = a[14] & g[26236];
assign g[59003] = b[14] & g[26236];
assign g[42621] = a[14] & g[26237];
assign g[59004] = b[14] & g[26237];
assign g[42622] = a[14] & g[26238];
assign g[59005] = b[14] & g[26238];
assign g[42623] = a[14] & g[26239];
assign g[59006] = b[14] & g[26239];
assign g[42624] = a[14] & g[26240];
assign g[59007] = b[14] & g[26240];
assign g[42625] = a[14] & g[26241];
assign g[59008] = b[14] & g[26241];
assign g[42626] = a[14] & g[26242];
assign g[59009] = b[14] & g[26242];
assign g[42627] = a[14] & g[26243];
assign g[59010] = b[14] & g[26243];
assign g[42628] = a[14] & g[26244];
assign g[59011] = b[14] & g[26244];
assign g[42629] = a[14] & g[26245];
assign g[59012] = b[14] & g[26245];
assign g[42630] = a[14] & g[26246];
assign g[59013] = b[14] & g[26246];
assign g[42631] = a[14] & g[26247];
assign g[59014] = b[14] & g[26247];
assign g[42632] = a[14] & g[26248];
assign g[59015] = b[14] & g[26248];
assign g[42633] = a[14] & g[26249];
assign g[59016] = b[14] & g[26249];
assign g[42634] = a[14] & g[26250];
assign g[59017] = b[14] & g[26250];
assign g[42635] = a[14] & g[26251];
assign g[59018] = b[14] & g[26251];
assign g[42636] = a[14] & g[26252];
assign g[59019] = b[14] & g[26252];
assign g[42637] = a[14] & g[26253];
assign g[59020] = b[14] & g[26253];
assign g[42638] = a[14] & g[26254];
assign g[59021] = b[14] & g[26254];
assign g[42639] = a[14] & g[26255];
assign g[59022] = b[14] & g[26255];
assign g[42640] = a[14] & g[26256];
assign g[59023] = b[14] & g[26256];
assign g[42641] = a[14] & g[26257];
assign g[59024] = b[14] & g[26257];
assign g[42642] = a[14] & g[26258];
assign g[59025] = b[14] & g[26258];
assign g[42643] = a[14] & g[26259];
assign g[59026] = b[14] & g[26259];
assign g[42644] = a[14] & g[26260];
assign g[59027] = b[14] & g[26260];
assign g[42645] = a[14] & g[26261];
assign g[59028] = b[14] & g[26261];
assign g[42646] = a[14] & g[26262];
assign g[59029] = b[14] & g[26262];
assign g[42647] = a[14] & g[26263];
assign g[59030] = b[14] & g[26263];
assign g[42648] = a[14] & g[26264];
assign g[59031] = b[14] & g[26264];
assign g[42649] = a[14] & g[26265];
assign g[59032] = b[14] & g[26265];
assign g[42650] = a[14] & g[26266];
assign g[59033] = b[14] & g[26266];
assign g[42651] = a[14] & g[26267];
assign g[59034] = b[14] & g[26267];
assign g[42652] = a[14] & g[26268];
assign g[59035] = b[14] & g[26268];
assign g[42653] = a[14] & g[26269];
assign g[59036] = b[14] & g[26269];
assign g[42654] = a[14] & g[26270];
assign g[59037] = b[14] & g[26270];
assign g[42655] = a[14] & g[26271];
assign g[59038] = b[14] & g[26271];
assign g[42656] = a[14] & g[26272];
assign g[59039] = b[14] & g[26272];
assign g[42657] = a[14] & g[26273];
assign g[59040] = b[14] & g[26273];
assign g[42658] = a[14] & g[26274];
assign g[59041] = b[14] & g[26274];
assign g[42659] = a[14] & g[26275];
assign g[59042] = b[14] & g[26275];
assign g[42660] = a[14] & g[26276];
assign g[59043] = b[14] & g[26276];
assign g[42661] = a[14] & g[26277];
assign g[59044] = b[14] & g[26277];
assign g[42662] = a[14] & g[26278];
assign g[59045] = b[14] & g[26278];
assign g[42663] = a[14] & g[26279];
assign g[59046] = b[14] & g[26279];
assign g[42664] = a[14] & g[26280];
assign g[59047] = b[14] & g[26280];
assign g[42665] = a[14] & g[26281];
assign g[59048] = b[14] & g[26281];
assign g[42666] = a[14] & g[26282];
assign g[59049] = b[14] & g[26282];
assign g[42667] = a[14] & g[26283];
assign g[59050] = b[14] & g[26283];
assign g[42668] = a[14] & g[26284];
assign g[59051] = b[14] & g[26284];
assign g[42669] = a[14] & g[26285];
assign g[59052] = b[14] & g[26285];
assign g[42670] = a[14] & g[26286];
assign g[59053] = b[14] & g[26286];
assign g[42671] = a[14] & g[26287];
assign g[59054] = b[14] & g[26287];
assign g[42672] = a[14] & g[26288];
assign g[59055] = b[14] & g[26288];
assign g[42673] = a[14] & g[26289];
assign g[59056] = b[14] & g[26289];
assign g[42674] = a[14] & g[26290];
assign g[59057] = b[14] & g[26290];
assign g[42675] = a[14] & g[26291];
assign g[59058] = b[14] & g[26291];
assign g[42676] = a[14] & g[26292];
assign g[59059] = b[14] & g[26292];
assign g[42677] = a[14] & g[26293];
assign g[59060] = b[14] & g[26293];
assign g[42678] = a[14] & g[26294];
assign g[59061] = b[14] & g[26294];
assign g[42679] = a[14] & g[26295];
assign g[59062] = b[14] & g[26295];
assign g[42680] = a[14] & g[26296];
assign g[59063] = b[14] & g[26296];
assign g[42681] = a[14] & g[26297];
assign g[59064] = b[14] & g[26297];
assign g[42682] = a[14] & g[26298];
assign g[59065] = b[14] & g[26298];
assign g[42683] = a[14] & g[26299];
assign g[59066] = b[14] & g[26299];
assign g[42684] = a[14] & g[26300];
assign g[59067] = b[14] & g[26300];
assign g[42685] = a[14] & g[26301];
assign g[59068] = b[14] & g[26301];
assign g[42686] = a[14] & g[26302];
assign g[59069] = b[14] & g[26302];
assign g[42687] = a[14] & g[26303];
assign g[59070] = b[14] & g[26303];
assign g[42688] = a[14] & g[26304];
assign g[59071] = b[14] & g[26304];
assign g[42689] = a[14] & g[26305];
assign g[59072] = b[14] & g[26305];
assign g[42690] = a[14] & g[26306];
assign g[59073] = b[14] & g[26306];
assign g[42691] = a[14] & g[26307];
assign g[59074] = b[14] & g[26307];
assign g[42692] = a[14] & g[26308];
assign g[59075] = b[14] & g[26308];
assign g[42693] = a[14] & g[26309];
assign g[59076] = b[14] & g[26309];
assign g[42694] = a[14] & g[26310];
assign g[59077] = b[14] & g[26310];
assign g[42695] = a[14] & g[26311];
assign g[59078] = b[14] & g[26311];
assign g[42696] = a[14] & g[26312];
assign g[59079] = b[14] & g[26312];
assign g[42697] = a[14] & g[26313];
assign g[59080] = b[14] & g[26313];
assign g[42698] = a[14] & g[26314];
assign g[59081] = b[14] & g[26314];
assign g[42699] = a[14] & g[26315];
assign g[59082] = b[14] & g[26315];
assign g[42700] = a[14] & g[26316];
assign g[59083] = b[14] & g[26316];
assign g[42701] = a[14] & g[26317];
assign g[59084] = b[14] & g[26317];
assign g[42702] = a[14] & g[26318];
assign g[59085] = b[14] & g[26318];
assign g[42703] = a[14] & g[26319];
assign g[59086] = b[14] & g[26319];
assign g[42704] = a[14] & g[26320];
assign g[59087] = b[14] & g[26320];
assign g[42705] = a[14] & g[26321];
assign g[59088] = b[14] & g[26321];
assign g[42706] = a[14] & g[26322];
assign g[59089] = b[14] & g[26322];
assign g[42707] = a[14] & g[26323];
assign g[59090] = b[14] & g[26323];
assign g[42708] = a[14] & g[26324];
assign g[59091] = b[14] & g[26324];
assign g[42709] = a[14] & g[26325];
assign g[59092] = b[14] & g[26325];
assign g[42710] = a[14] & g[26326];
assign g[59093] = b[14] & g[26326];
assign g[42711] = a[14] & g[26327];
assign g[59094] = b[14] & g[26327];
assign g[42712] = a[14] & g[26328];
assign g[59095] = b[14] & g[26328];
assign g[42713] = a[14] & g[26329];
assign g[59096] = b[14] & g[26329];
assign g[42714] = a[14] & g[26330];
assign g[59097] = b[14] & g[26330];
assign g[42715] = a[14] & g[26331];
assign g[59098] = b[14] & g[26331];
assign g[42716] = a[14] & g[26332];
assign g[59099] = b[14] & g[26332];
assign g[42717] = a[14] & g[26333];
assign g[59100] = b[14] & g[26333];
assign g[42718] = a[14] & g[26334];
assign g[59101] = b[14] & g[26334];
assign g[42719] = a[14] & g[26335];
assign g[59102] = b[14] & g[26335];
assign g[42720] = a[14] & g[26336];
assign g[59103] = b[14] & g[26336];
assign g[42721] = a[14] & g[26337];
assign g[59104] = b[14] & g[26337];
assign g[42722] = a[14] & g[26338];
assign g[59105] = b[14] & g[26338];
assign g[42723] = a[14] & g[26339];
assign g[59106] = b[14] & g[26339];
assign g[42724] = a[14] & g[26340];
assign g[59107] = b[14] & g[26340];
assign g[42725] = a[14] & g[26341];
assign g[59108] = b[14] & g[26341];
assign g[42726] = a[14] & g[26342];
assign g[59109] = b[14] & g[26342];
assign g[42727] = a[14] & g[26343];
assign g[59110] = b[14] & g[26343];
assign g[42728] = a[14] & g[26344];
assign g[59111] = b[14] & g[26344];
assign g[42729] = a[14] & g[26345];
assign g[59112] = b[14] & g[26345];
assign g[42730] = a[14] & g[26346];
assign g[59113] = b[14] & g[26346];
assign g[42731] = a[14] & g[26347];
assign g[59114] = b[14] & g[26347];
assign g[42732] = a[14] & g[26348];
assign g[59115] = b[14] & g[26348];
assign g[42733] = a[14] & g[26349];
assign g[59116] = b[14] & g[26349];
assign g[42734] = a[14] & g[26350];
assign g[59117] = b[14] & g[26350];
assign g[42735] = a[14] & g[26351];
assign g[59118] = b[14] & g[26351];
assign g[42736] = a[14] & g[26352];
assign g[59119] = b[14] & g[26352];
assign g[42737] = a[14] & g[26353];
assign g[59120] = b[14] & g[26353];
assign g[42738] = a[14] & g[26354];
assign g[59121] = b[14] & g[26354];
assign g[42739] = a[14] & g[26355];
assign g[59122] = b[14] & g[26355];
assign g[42740] = a[14] & g[26356];
assign g[59123] = b[14] & g[26356];
assign g[42741] = a[14] & g[26357];
assign g[59124] = b[14] & g[26357];
assign g[42742] = a[14] & g[26358];
assign g[59125] = b[14] & g[26358];
assign g[42743] = a[14] & g[26359];
assign g[59126] = b[14] & g[26359];
assign g[42744] = a[14] & g[26360];
assign g[59127] = b[14] & g[26360];
assign g[42745] = a[14] & g[26361];
assign g[59128] = b[14] & g[26361];
assign g[42746] = a[14] & g[26362];
assign g[59129] = b[14] & g[26362];
assign g[42747] = a[14] & g[26363];
assign g[59130] = b[14] & g[26363];
assign g[42748] = a[14] & g[26364];
assign g[59131] = b[14] & g[26364];
assign g[42749] = a[14] & g[26365];
assign g[59132] = b[14] & g[26365];
assign g[42750] = a[14] & g[26366];
assign g[59133] = b[14] & g[26366];
assign g[42751] = a[14] & g[26367];
assign g[59134] = b[14] & g[26367];
assign g[42752] = a[14] & g[26368];
assign g[59135] = b[14] & g[26368];
assign g[42753] = a[14] & g[26369];
assign g[59136] = b[14] & g[26369];
assign g[42754] = a[14] & g[26370];
assign g[59137] = b[14] & g[26370];
assign g[42755] = a[14] & g[26371];
assign g[59138] = b[14] & g[26371];
assign g[42756] = a[14] & g[26372];
assign g[59139] = b[14] & g[26372];
assign g[42757] = a[14] & g[26373];
assign g[59140] = b[14] & g[26373];
assign g[42758] = a[14] & g[26374];
assign g[59141] = b[14] & g[26374];
assign g[42759] = a[14] & g[26375];
assign g[59142] = b[14] & g[26375];
assign g[42760] = a[14] & g[26376];
assign g[59143] = b[14] & g[26376];
assign g[42761] = a[14] & g[26377];
assign g[59144] = b[14] & g[26377];
assign g[42762] = a[14] & g[26378];
assign g[59145] = b[14] & g[26378];
assign g[42763] = a[14] & g[26379];
assign g[59146] = b[14] & g[26379];
assign g[42764] = a[14] & g[26380];
assign g[59147] = b[14] & g[26380];
assign g[42765] = a[14] & g[26381];
assign g[59148] = b[14] & g[26381];
assign g[42766] = a[14] & g[26382];
assign g[59149] = b[14] & g[26382];
assign g[42767] = a[14] & g[26383];
assign g[59150] = b[14] & g[26383];
assign g[42768] = a[14] & g[26384];
assign g[59151] = b[14] & g[26384];
assign g[42769] = a[14] & g[26385];
assign g[59152] = b[14] & g[26385];
assign g[42770] = a[14] & g[26386];
assign g[59153] = b[14] & g[26386];
assign g[42771] = a[14] & g[26387];
assign g[59154] = b[14] & g[26387];
assign g[42772] = a[14] & g[26388];
assign g[59155] = b[14] & g[26388];
assign g[42773] = a[14] & g[26389];
assign g[59156] = b[14] & g[26389];
assign g[42774] = a[14] & g[26390];
assign g[59157] = b[14] & g[26390];
assign g[42775] = a[14] & g[26391];
assign g[59158] = b[14] & g[26391];
assign g[42776] = a[14] & g[26392];
assign g[59159] = b[14] & g[26392];
assign g[42777] = a[14] & g[26393];
assign g[59160] = b[14] & g[26393];
assign g[42778] = a[14] & g[26394];
assign g[59161] = b[14] & g[26394];
assign g[42779] = a[14] & g[26395];
assign g[59162] = b[14] & g[26395];
assign g[42780] = a[14] & g[26396];
assign g[59163] = b[14] & g[26396];
assign g[42781] = a[14] & g[26397];
assign g[59164] = b[14] & g[26397];
assign g[42782] = a[14] & g[26398];
assign g[59165] = b[14] & g[26398];
assign g[42783] = a[14] & g[26399];
assign g[59166] = b[14] & g[26399];
assign g[42784] = a[14] & g[26400];
assign g[59167] = b[14] & g[26400];
assign g[42785] = a[14] & g[26401];
assign g[59168] = b[14] & g[26401];
assign g[42786] = a[14] & g[26402];
assign g[59169] = b[14] & g[26402];
assign g[42787] = a[14] & g[26403];
assign g[59170] = b[14] & g[26403];
assign g[42788] = a[14] & g[26404];
assign g[59171] = b[14] & g[26404];
assign g[42789] = a[14] & g[26405];
assign g[59172] = b[14] & g[26405];
assign g[42790] = a[14] & g[26406];
assign g[59173] = b[14] & g[26406];
assign g[42791] = a[14] & g[26407];
assign g[59174] = b[14] & g[26407];
assign g[42792] = a[14] & g[26408];
assign g[59175] = b[14] & g[26408];
assign g[42793] = a[14] & g[26409];
assign g[59176] = b[14] & g[26409];
assign g[42794] = a[14] & g[26410];
assign g[59177] = b[14] & g[26410];
assign g[42795] = a[14] & g[26411];
assign g[59178] = b[14] & g[26411];
assign g[42796] = a[14] & g[26412];
assign g[59179] = b[14] & g[26412];
assign g[42797] = a[14] & g[26413];
assign g[59180] = b[14] & g[26413];
assign g[42798] = a[14] & g[26414];
assign g[59181] = b[14] & g[26414];
assign g[42799] = a[14] & g[26415];
assign g[59182] = b[14] & g[26415];
assign g[42800] = a[14] & g[26416];
assign g[59183] = b[14] & g[26416];
assign g[42801] = a[14] & g[26417];
assign g[59184] = b[14] & g[26417];
assign g[42802] = a[14] & g[26418];
assign g[59185] = b[14] & g[26418];
assign g[42803] = a[14] & g[26419];
assign g[59186] = b[14] & g[26419];
assign g[42804] = a[14] & g[26420];
assign g[59187] = b[14] & g[26420];
assign g[42805] = a[14] & g[26421];
assign g[59188] = b[14] & g[26421];
assign g[42806] = a[14] & g[26422];
assign g[59189] = b[14] & g[26422];
assign g[42807] = a[14] & g[26423];
assign g[59190] = b[14] & g[26423];
assign g[42808] = a[14] & g[26424];
assign g[59191] = b[14] & g[26424];
assign g[42809] = a[14] & g[26425];
assign g[59192] = b[14] & g[26425];
assign g[42810] = a[14] & g[26426];
assign g[59193] = b[14] & g[26426];
assign g[42811] = a[14] & g[26427];
assign g[59194] = b[14] & g[26427];
assign g[42812] = a[14] & g[26428];
assign g[59195] = b[14] & g[26428];
assign g[42813] = a[14] & g[26429];
assign g[59196] = b[14] & g[26429];
assign g[42814] = a[14] & g[26430];
assign g[59197] = b[14] & g[26430];
assign g[42815] = a[14] & g[26431];
assign g[59198] = b[14] & g[26431];
assign g[42816] = a[14] & g[26432];
assign g[59199] = b[14] & g[26432];
assign g[42817] = a[14] & g[26433];
assign g[59200] = b[14] & g[26433];
assign g[42818] = a[14] & g[26434];
assign g[59201] = b[14] & g[26434];
assign g[42819] = a[14] & g[26435];
assign g[59202] = b[14] & g[26435];
assign g[42820] = a[14] & g[26436];
assign g[59203] = b[14] & g[26436];
assign g[42821] = a[14] & g[26437];
assign g[59204] = b[14] & g[26437];
assign g[42822] = a[14] & g[26438];
assign g[59205] = b[14] & g[26438];
assign g[42823] = a[14] & g[26439];
assign g[59206] = b[14] & g[26439];
assign g[42824] = a[14] & g[26440];
assign g[59207] = b[14] & g[26440];
assign g[42825] = a[14] & g[26441];
assign g[59208] = b[14] & g[26441];
assign g[42826] = a[14] & g[26442];
assign g[59209] = b[14] & g[26442];
assign g[42827] = a[14] & g[26443];
assign g[59210] = b[14] & g[26443];
assign g[42828] = a[14] & g[26444];
assign g[59211] = b[14] & g[26444];
assign g[42829] = a[14] & g[26445];
assign g[59212] = b[14] & g[26445];
assign g[42830] = a[14] & g[26446];
assign g[59213] = b[14] & g[26446];
assign g[42831] = a[14] & g[26447];
assign g[59214] = b[14] & g[26447];
assign g[42832] = a[14] & g[26448];
assign g[59215] = b[14] & g[26448];
assign g[42833] = a[14] & g[26449];
assign g[59216] = b[14] & g[26449];
assign g[42834] = a[14] & g[26450];
assign g[59217] = b[14] & g[26450];
assign g[42835] = a[14] & g[26451];
assign g[59218] = b[14] & g[26451];
assign g[42836] = a[14] & g[26452];
assign g[59219] = b[14] & g[26452];
assign g[42837] = a[14] & g[26453];
assign g[59220] = b[14] & g[26453];
assign g[42838] = a[14] & g[26454];
assign g[59221] = b[14] & g[26454];
assign g[42839] = a[14] & g[26455];
assign g[59222] = b[14] & g[26455];
assign g[42840] = a[14] & g[26456];
assign g[59223] = b[14] & g[26456];
assign g[42841] = a[14] & g[26457];
assign g[59224] = b[14] & g[26457];
assign g[42842] = a[14] & g[26458];
assign g[59225] = b[14] & g[26458];
assign g[42843] = a[14] & g[26459];
assign g[59226] = b[14] & g[26459];
assign g[42844] = a[14] & g[26460];
assign g[59227] = b[14] & g[26460];
assign g[42845] = a[14] & g[26461];
assign g[59228] = b[14] & g[26461];
assign g[42846] = a[14] & g[26462];
assign g[59229] = b[14] & g[26462];
assign g[42847] = a[14] & g[26463];
assign g[59230] = b[14] & g[26463];
assign g[42848] = a[14] & g[26464];
assign g[59231] = b[14] & g[26464];
assign g[42849] = a[14] & g[26465];
assign g[59232] = b[14] & g[26465];
assign g[42850] = a[14] & g[26466];
assign g[59233] = b[14] & g[26466];
assign g[42851] = a[14] & g[26467];
assign g[59234] = b[14] & g[26467];
assign g[42852] = a[14] & g[26468];
assign g[59235] = b[14] & g[26468];
assign g[42853] = a[14] & g[26469];
assign g[59236] = b[14] & g[26469];
assign g[42854] = a[14] & g[26470];
assign g[59237] = b[14] & g[26470];
assign g[42855] = a[14] & g[26471];
assign g[59238] = b[14] & g[26471];
assign g[42856] = a[14] & g[26472];
assign g[59239] = b[14] & g[26472];
assign g[42857] = a[14] & g[26473];
assign g[59240] = b[14] & g[26473];
assign g[42858] = a[14] & g[26474];
assign g[59241] = b[14] & g[26474];
assign g[42859] = a[14] & g[26475];
assign g[59242] = b[14] & g[26475];
assign g[42860] = a[14] & g[26476];
assign g[59243] = b[14] & g[26476];
assign g[42861] = a[14] & g[26477];
assign g[59244] = b[14] & g[26477];
assign g[42862] = a[14] & g[26478];
assign g[59245] = b[14] & g[26478];
assign g[42863] = a[14] & g[26479];
assign g[59246] = b[14] & g[26479];
assign g[42864] = a[14] & g[26480];
assign g[59247] = b[14] & g[26480];
assign g[42865] = a[14] & g[26481];
assign g[59248] = b[14] & g[26481];
assign g[42866] = a[14] & g[26482];
assign g[59249] = b[14] & g[26482];
assign g[42867] = a[14] & g[26483];
assign g[59250] = b[14] & g[26483];
assign g[42868] = a[14] & g[26484];
assign g[59251] = b[14] & g[26484];
assign g[42869] = a[14] & g[26485];
assign g[59252] = b[14] & g[26485];
assign g[42870] = a[14] & g[26486];
assign g[59253] = b[14] & g[26486];
assign g[42871] = a[14] & g[26487];
assign g[59254] = b[14] & g[26487];
assign g[42872] = a[14] & g[26488];
assign g[59255] = b[14] & g[26488];
assign g[42873] = a[14] & g[26489];
assign g[59256] = b[14] & g[26489];
assign g[42874] = a[14] & g[26490];
assign g[59257] = b[14] & g[26490];
assign g[42875] = a[14] & g[26491];
assign g[59258] = b[14] & g[26491];
assign g[42876] = a[14] & g[26492];
assign g[59259] = b[14] & g[26492];
assign g[42877] = a[14] & g[26493];
assign g[59260] = b[14] & g[26493];
assign g[42878] = a[14] & g[26494];
assign g[59261] = b[14] & g[26494];
assign g[42879] = a[14] & g[26495];
assign g[59262] = b[14] & g[26495];
assign g[42880] = a[14] & g[26496];
assign g[59263] = b[14] & g[26496];
assign g[42881] = a[14] & g[26497];
assign g[59264] = b[14] & g[26497];
assign g[42882] = a[14] & g[26498];
assign g[59265] = b[14] & g[26498];
assign g[42883] = a[14] & g[26499];
assign g[59266] = b[14] & g[26499];
assign g[42884] = a[14] & g[26500];
assign g[59267] = b[14] & g[26500];
assign g[42885] = a[14] & g[26501];
assign g[59268] = b[14] & g[26501];
assign g[42886] = a[14] & g[26502];
assign g[59269] = b[14] & g[26502];
assign g[42887] = a[14] & g[26503];
assign g[59270] = b[14] & g[26503];
assign g[42888] = a[14] & g[26504];
assign g[59271] = b[14] & g[26504];
assign g[42889] = a[14] & g[26505];
assign g[59272] = b[14] & g[26505];
assign g[42890] = a[14] & g[26506];
assign g[59273] = b[14] & g[26506];
assign g[42891] = a[14] & g[26507];
assign g[59274] = b[14] & g[26507];
assign g[42892] = a[14] & g[26508];
assign g[59275] = b[14] & g[26508];
assign g[42893] = a[14] & g[26509];
assign g[59276] = b[14] & g[26509];
assign g[42894] = a[14] & g[26510];
assign g[59277] = b[14] & g[26510];
assign g[42895] = a[14] & g[26511];
assign g[59278] = b[14] & g[26511];
assign g[42896] = a[14] & g[26512];
assign g[59279] = b[14] & g[26512];
assign g[42897] = a[14] & g[26513];
assign g[59280] = b[14] & g[26513];
assign g[42898] = a[14] & g[26514];
assign g[59281] = b[14] & g[26514];
assign g[42899] = a[14] & g[26515];
assign g[59282] = b[14] & g[26515];
assign g[42900] = a[14] & g[26516];
assign g[59283] = b[14] & g[26516];
assign g[42901] = a[14] & g[26517];
assign g[59284] = b[14] & g[26517];
assign g[42902] = a[14] & g[26518];
assign g[59285] = b[14] & g[26518];
assign g[42903] = a[14] & g[26519];
assign g[59286] = b[14] & g[26519];
assign g[42904] = a[14] & g[26520];
assign g[59287] = b[14] & g[26520];
assign g[42905] = a[14] & g[26521];
assign g[59288] = b[14] & g[26521];
assign g[42906] = a[14] & g[26522];
assign g[59289] = b[14] & g[26522];
assign g[42907] = a[14] & g[26523];
assign g[59290] = b[14] & g[26523];
assign g[42908] = a[14] & g[26524];
assign g[59291] = b[14] & g[26524];
assign g[42909] = a[14] & g[26525];
assign g[59292] = b[14] & g[26525];
assign g[42910] = a[14] & g[26526];
assign g[59293] = b[14] & g[26526];
assign g[42911] = a[14] & g[26527];
assign g[59294] = b[14] & g[26527];
assign g[42912] = a[14] & g[26528];
assign g[59295] = b[14] & g[26528];
assign g[42913] = a[14] & g[26529];
assign g[59296] = b[14] & g[26529];
assign g[42914] = a[14] & g[26530];
assign g[59297] = b[14] & g[26530];
assign g[42915] = a[14] & g[26531];
assign g[59298] = b[14] & g[26531];
assign g[42916] = a[14] & g[26532];
assign g[59299] = b[14] & g[26532];
assign g[42917] = a[14] & g[26533];
assign g[59300] = b[14] & g[26533];
assign g[42918] = a[14] & g[26534];
assign g[59301] = b[14] & g[26534];
assign g[42919] = a[14] & g[26535];
assign g[59302] = b[14] & g[26535];
assign g[42920] = a[14] & g[26536];
assign g[59303] = b[14] & g[26536];
assign g[42921] = a[14] & g[26537];
assign g[59304] = b[14] & g[26537];
assign g[42922] = a[14] & g[26538];
assign g[59305] = b[14] & g[26538];
assign g[42923] = a[14] & g[26539];
assign g[59306] = b[14] & g[26539];
assign g[42924] = a[14] & g[26540];
assign g[59307] = b[14] & g[26540];
assign g[42925] = a[14] & g[26541];
assign g[59308] = b[14] & g[26541];
assign g[42926] = a[14] & g[26542];
assign g[59309] = b[14] & g[26542];
assign g[42927] = a[14] & g[26543];
assign g[59310] = b[14] & g[26543];
assign g[42928] = a[14] & g[26544];
assign g[59311] = b[14] & g[26544];
assign g[42929] = a[14] & g[26545];
assign g[59312] = b[14] & g[26545];
assign g[42930] = a[14] & g[26546];
assign g[59313] = b[14] & g[26546];
assign g[42931] = a[14] & g[26547];
assign g[59314] = b[14] & g[26547];
assign g[42932] = a[14] & g[26548];
assign g[59315] = b[14] & g[26548];
assign g[42933] = a[14] & g[26549];
assign g[59316] = b[14] & g[26549];
assign g[42934] = a[14] & g[26550];
assign g[59317] = b[14] & g[26550];
assign g[42935] = a[14] & g[26551];
assign g[59318] = b[14] & g[26551];
assign g[42936] = a[14] & g[26552];
assign g[59319] = b[14] & g[26552];
assign g[42937] = a[14] & g[26553];
assign g[59320] = b[14] & g[26553];
assign g[42938] = a[14] & g[26554];
assign g[59321] = b[14] & g[26554];
assign g[42939] = a[14] & g[26555];
assign g[59322] = b[14] & g[26555];
assign g[42940] = a[14] & g[26556];
assign g[59323] = b[14] & g[26556];
assign g[42941] = a[14] & g[26557];
assign g[59324] = b[14] & g[26557];
assign g[42942] = a[14] & g[26558];
assign g[59325] = b[14] & g[26558];
assign g[42943] = a[14] & g[26559];
assign g[59326] = b[14] & g[26559];
assign g[42944] = a[14] & g[26560];
assign g[59327] = b[14] & g[26560];
assign g[42945] = a[14] & g[26561];
assign g[59328] = b[14] & g[26561];
assign g[42946] = a[14] & g[26562];
assign g[59329] = b[14] & g[26562];
assign g[42947] = a[14] & g[26563];
assign g[59330] = b[14] & g[26563];
assign g[42948] = a[14] & g[26564];
assign g[59331] = b[14] & g[26564];
assign g[42949] = a[14] & g[26565];
assign g[59332] = b[14] & g[26565];
assign g[42950] = a[14] & g[26566];
assign g[59333] = b[14] & g[26566];
assign g[42951] = a[14] & g[26567];
assign g[59334] = b[14] & g[26567];
assign g[42952] = a[14] & g[26568];
assign g[59335] = b[14] & g[26568];
assign g[42953] = a[14] & g[26569];
assign g[59336] = b[14] & g[26569];
assign g[42954] = a[14] & g[26570];
assign g[59337] = b[14] & g[26570];
assign g[42955] = a[14] & g[26571];
assign g[59338] = b[14] & g[26571];
assign g[42956] = a[14] & g[26572];
assign g[59339] = b[14] & g[26572];
assign g[42957] = a[14] & g[26573];
assign g[59340] = b[14] & g[26573];
assign g[42958] = a[14] & g[26574];
assign g[59341] = b[14] & g[26574];
assign g[42959] = a[14] & g[26575];
assign g[59342] = b[14] & g[26575];
assign g[42960] = a[14] & g[26576];
assign g[59343] = b[14] & g[26576];
assign g[42961] = a[14] & g[26577];
assign g[59344] = b[14] & g[26577];
assign g[42962] = a[14] & g[26578];
assign g[59345] = b[14] & g[26578];
assign g[42963] = a[14] & g[26579];
assign g[59346] = b[14] & g[26579];
assign g[42964] = a[14] & g[26580];
assign g[59347] = b[14] & g[26580];
assign g[42965] = a[14] & g[26581];
assign g[59348] = b[14] & g[26581];
assign g[42966] = a[14] & g[26582];
assign g[59349] = b[14] & g[26582];
assign g[42967] = a[14] & g[26583];
assign g[59350] = b[14] & g[26583];
assign g[42968] = a[14] & g[26584];
assign g[59351] = b[14] & g[26584];
assign g[42969] = a[14] & g[26585];
assign g[59352] = b[14] & g[26585];
assign g[42970] = a[14] & g[26586];
assign g[59353] = b[14] & g[26586];
assign g[42971] = a[14] & g[26587];
assign g[59354] = b[14] & g[26587];
assign g[42972] = a[14] & g[26588];
assign g[59355] = b[14] & g[26588];
assign g[42973] = a[14] & g[26589];
assign g[59356] = b[14] & g[26589];
assign g[42974] = a[14] & g[26590];
assign g[59357] = b[14] & g[26590];
assign g[42975] = a[14] & g[26591];
assign g[59358] = b[14] & g[26591];
assign g[42976] = a[14] & g[26592];
assign g[59359] = b[14] & g[26592];
assign g[42977] = a[14] & g[26593];
assign g[59360] = b[14] & g[26593];
assign g[42978] = a[14] & g[26594];
assign g[59361] = b[14] & g[26594];
assign g[42979] = a[14] & g[26595];
assign g[59362] = b[14] & g[26595];
assign g[42980] = a[14] & g[26596];
assign g[59363] = b[14] & g[26596];
assign g[42981] = a[14] & g[26597];
assign g[59364] = b[14] & g[26597];
assign g[42982] = a[14] & g[26598];
assign g[59365] = b[14] & g[26598];
assign g[42983] = a[14] & g[26599];
assign g[59366] = b[14] & g[26599];
assign g[42984] = a[14] & g[26600];
assign g[59367] = b[14] & g[26600];
assign g[42985] = a[14] & g[26601];
assign g[59368] = b[14] & g[26601];
assign g[42986] = a[14] & g[26602];
assign g[59369] = b[14] & g[26602];
assign g[42987] = a[14] & g[26603];
assign g[59370] = b[14] & g[26603];
assign g[42988] = a[14] & g[26604];
assign g[59371] = b[14] & g[26604];
assign g[42989] = a[14] & g[26605];
assign g[59372] = b[14] & g[26605];
assign g[42990] = a[14] & g[26606];
assign g[59373] = b[14] & g[26606];
assign g[42991] = a[14] & g[26607];
assign g[59374] = b[14] & g[26607];
assign g[42992] = a[14] & g[26608];
assign g[59375] = b[14] & g[26608];
assign g[42993] = a[14] & g[26609];
assign g[59376] = b[14] & g[26609];
assign g[42994] = a[14] & g[26610];
assign g[59377] = b[14] & g[26610];
assign g[42995] = a[14] & g[26611];
assign g[59378] = b[14] & g[26611];
assign g[42996] = a[14] & g[26612];
assign g[59379] = b[14] & g[26612];
assign g[42997] = a[14] & g[26613];
assign g[59380] = b[14] & g[26613];
assign g[42998] = a[14] & g[26614];
assign g[59381] = b[14] & g[26614];
assign g[42999] = a[14] & g[26615];
assign g[59382] = b[14] & g[26615];
assign g[43000] = a[14] & g[26616];
assign g[59383] = b[14] & g[26616];
assign g[43001] = a[14] & g[26617];
assign g[59384] = b[14] & g[26617];
assign g[43002] = a[14] & g[26618];
assign g[59385] = b[14] & g[26618];
assign g[43003] = a[14] & g[26619];
assign g[59386] = b[14] & g[26619];
assign g[43004] = a[14] & g[26620];
assign g[59387] = b[14] & g[26620];
assign g[43005] = a[14] & g[26621];
assign g[59388] = b[14] & g[26621];
assign g[43006] = a[14] & g[26622];
assign g[59389] = b[14] & g[26622];
assign g[43007] = a[14] & g[26623];
assign g[59390] = b[14] & g[26623];
assign g[43008] = a[14] & g[26624];
assign g[59391] = b[14] & g[26624];
assign g[43009] = a[14] & g[26625];
assign g[59392] = b[14] & g[26625];
assign g[43010] = a[14] & g[26626];
assign g[59393] = b[14] & g[26626];
assign g[43011] = a[14] & g[26627];
assign g[59394] = b[14] & g[26627];
assign g[43012] = a[14] & g[26628];
assign g[59395] = b[14] & g[26628];
assign g[43013] = a[14] & g[26629];
assign g[59396] = b[14] & g[26629];
assign g[43014] = a[14] & g[26630];
assign g[59397] = b[14] & g[26630];
assign g[43015] = a[14] & g[26631];
assign g[59398] = b[14] & g[26631];
assign g[43016] = a[14] & g[26632];
assign g[59399] = b[14] & g[26632];
assign g[43017] = a[14] & g[26633];
assign g[59400] = b[14] & g[26633];
assign g[43018] = a[14] & g[26634];
assign g[59401] = b[14] & g[26634];
assign g[43019] = a[14] & g[26635];
assign g[59402] = b[14] & g[26635];
assign g[43020] = a[14] & g[26636];
assign g[59403] = b[14] & g[26636];
assign g[43021] = a[14] & g[26637];
assign g[59404] = b[14] & g[26637];
assign g[43022] = a[14] & g[26638];
assign g[59405] = b[14] & g[26638];
assign g[43023] = a[14] & g[26639];
assign g[59406] = b[14] & g[26639];
assign g[43024] = a[14] & g[26640];
assign g[59407] = b[14] & g[26640];
assign g[43025] = a[14] & g[26641];
assign g[59408] = b[14] & g[26641];
assign g[43026] = a[14] & g[26642];
assign g[59409] = b[14] & g[26642];
assign g[43027] = a[14] & g[26643];
assign g[59410] = b[14] & g[26643];
assign g[43028] = a[14] & g[26644];
assign g[59411] = b[14] & g[26644];
assign g[43029] = a[14] & g[26645];
assign g[59412] = b[14] & g[26645];
assign g[43030] = a[14] & g[26646];
assign g[59413] = b[14] & g[26646];
assign g[43031] = a[14] & g[26647];
assign g[59414] = b[14] & g[26647];
assign g[43032] = a[14] & g[26648];
assign g[59415] = b[14] & g[26648];
assign g[43033] = a[14] & g[26649];
assign g[59416] = b[14] & g[26649];
assign g[43034] = a[14] & g[26650];
assign g[59417] = b[14] & g[26650];
assign g[43035] = a[14] & g[26651];
assign g[59418] = b[14] & g[26651];
assign g[43036] = a[14] & g[26652];
assign g[59419] = b[14] & g[26652];
assign g[43037] = a[14] & g[26653];
assign g[59420] = b[14] & g[26653];
assign g[43038] = a[14] & g[26654];
assign g[59421] = b[14] & g[26654];
assign g[43039] = a[14] & g[26655];
assign g[59422] = b[14] & g[26655];
assign g[43040] = a[14] & g[26656];
assign g[59423] = b[14] & g[26656];
assign g[43041] = a[14] & g[26657];
assign g[59424] = b[14] & g[26657];
assign g[43042] = a[14] & g[26658];
assign g[59425] = b[14] & g[26658];
assign g[43043] = a[14] & g[26659];
assign g[59426] = b[14] & g[26659];
assign g[43044] = a[14] & g[26660];
assign g[59427] = b[14] & g[26660];
assign g[43045] = a[14] & g[26661];
assign g[59428] = b[14] & g[26661];
assign g[43046] = a[14] & g[26662];
assign g[59429] = b[14] & g[26662];
assign g[43047] = a[14] & g[26663];
assign g[59430] = b[14] & g[26663];
assign g[43048] = a[14] & g[26664];
assign g[59431] = b[14] & g[26664];
assign g[43049] = a[14] & g[26665];
assign g[59432] = b[14] & g[26665];
assign g[43050] = a[14] & g[26666];
assign g[59433] = b[14] & g[26666];
assign g[43051] = a[14] & g[26667];
assign g[59434] = b[14] & g[26667];
assign g[43052] = a[14] & g[26668];
assign g[59435] = b[14] & g[26668];
assign g[43053] = a[14] & g[26669];
assign g[59436] = b[14] & g[26669];
assign g[43054] = a[14] & g[26670];
assign g[59437] = b[14] & g[26670];
assign g[43055] = a[14] & g[26671];
assign g[59438] = b[14] & g[26671];
assign g[43056] = a[14] & g[26672];
assign g[59439] = b[14] & g[26672];
assign g[43057] = a[14] & g[26673];
assign g[59440] = b[14] & g[26673];
assign g[43058] = a[14] & g[26674];
assign g[59441] = b[14] & g[26674];
assign g[43059] = a[14] & g[26675];
assign g[59442] = b[14] & g[26675];
assign g[43060] = a[14] & g[26676];
assign g[59443] = b[14] & g[26676];
assign g[43061] = a[14] & g[26677];
assign g[59444] = b[14] & g[26677];
assign g[43062] = a[14] & g[26678];
assign g[59445] = b[14] & g[26678];
assign g[43063] = a[14] & g[26679];
assign g[59446] = b[14] & g[26679];
assign g[43064] = a[14] & g[26680];
assign g[59447] = b[14] & g[26680];
assign g[43065] = a[14] & g[26681];
assign g[59448] = b[14] & g[26681];
assign g[43066] = a[14] & g[26682];
assign g[59449] = b[14] & g[26682];
assign g[43067] = a[14] & g[26683];
assign g[59450] = b[14] & g[26683];
assign g[43068] = a[14] & g[26684];
assign g[59451] = b[14] & g[26684];
assign g[43069] = a[14] & g[26685];
assign g[59452] = b[14] & g[26685];
assign g[43070] = a[14] & g[26686];
assign g[59453] = b[14] & g[26686];
assign g[43071] = a[14] & g[26687];
assign g[59454] = b[14] & g[26687];
assign g[43072] = a[14] & g[26688];
assign g[59455] = b[14] & g[26688];
assign g[43073] = a[14] & g[26689];
assign g[59456] = b[14] & g[26689];
assign g[43074] = a[14] & g[26690];
assign g[59457] = b[14] & g[26690];
assign g[43075] = a[14] & g[26691];
assign g[59458] = b[14] & g[26691];
assign g[43076] = a[14] & g[26692];
assign g[59459] = b[14] & g[26692];
assign g[43077] = a[14] & g[26693];
assign g[59460] = b[14] & g[26693];
assign g[43078] = a[14] & g[26694];
assign g[59461] = b[14] & g[26694];
assign g[43079] = a[14] & g[26695];
assign g[59462] = b[14] & g[26695];
assign g[43080] = a[14] & g[26696];
assign g[59463] = b[14] & g[26696];
assign g[43081] = a[14] & g[26697];
assign g[59464] = b[14] & g[26697];
assign g[43082] = a[14] & g[26698];
assign g[59465] = b[14] & g[26698];
assign g[43083] = a[14] & g[26699];
assign g[59466] = b[14] & g[26699];
assign g[43084] = a[14] & g[26700];
assign g[59467] = b[14] & g[26700];
assign g[43085] = a[14] & g[26701];
assign g[59468] = b[14] & g[26701];
assign g[43086] = a[14] & g[26702];
assign g[59469] = b[14] & g[26702];
assign g[43087] = a[14] & g[26703];
assign g[59470] = b[14] & g[26703];
assign g[43088] = a[14] & g[26704];
assign g[59471] = b[14] & g[26704];
assign g[43089] = a[14] & g[26705];
assign g[59472] = b[14] & g[26705];
assign g[43090] = a[14] & g[26706];
assign g[59473] = b[14] & g[26706];
assign g[43091] = a[14] & g[26707];
assign g[59474] = b[14] & g[26707];
assign g[43092] = a[14] & g[26708];
assign g[59475] = b[14] & g[26708];
assign g[43093] = a[14] & g[26709];
assign g[59476] = b[14] & g[26709];
assign g[43094] = a[14] & g[26710];
assign g[59477] = b[14] & g[26710];
assign g[43095] = a[14] & g[26711];
assign g[59478] = b[14] & g[26711];
assign g[43096] = a[14] & g[26712];
assign g[59479] = b[14] & g[26712];
assign g[43097] = a[14] & g[26713];
assign g[59480] = b[14] & g[26713];
assign g[43098] = a[14] & g[26714];
assign g[59481] = b[14] & g[26714];
assign g[43099] = a[14] & g[26715];
assign g[59482] = b[14] & g[26715];
assign g[43100] = a[14] & g[26716];
assign g[59483] = b[14] & g[26716];
assign g[43101] = a[14] & g[26717];
assign g[59484] = b[14] & g[26717];
assign g[43102] = a[14] & g[26718];
assign g[59485] = b[14] & g[26718];
assign g[43103] = a[14] & g[26719];
assign g[59486] = b[14] & g[26719];
assign g[43104] = a[14] & g[26720];
assign g[59487] = b[14] & g[26720];
assign g[43105] = a[14] & g[26721];
assign g[59488] = b[14] & g[26721];
assign g[43106] = a[14] & g[26722];
assign g[59489] = b[14] & g[26722];
assign g[43107] = a[14] & g[26723];
assign g[59490] = b[14] & g[26723];
assign g[43108] = a[14] & g[26724];
assign g[59491] = b[14] & g[26724];
assign g[43109] = a[14] & g[26725];
assign g[59492] = b[14] & g[26725];
assign g[43110] = a[14] & g[26726];
assign g[59493] = b[14] & g[26726];
assign g[43111] = a[14] & g[26727];
assign g[59494] = b[14] & g[26727];
assign g[43112] = a[14] & g[26728];
assign g[59495] = b[14] & g[26728];
assign g[43113] = a[14] & g[26729];
assign g[59496] = b[14] & g[26729];
assign g[43114] = a[14] & g[26730];
assign g[59497] = b[14] & g[26730];
assign g[43115] = a[14] & g[26731];
assign g[59498] = b[14] & g[26731];
assign g[43116] = a[14] & g[26732];
assign g[59499] = b[14] & g[26732];
assign g[43117] = a[14] & g[26733];
assign g[59500] = b[14] & g[26733];
assign g[43118] = a[14] & g[26734];
assign g[59501] = b[14] & g[26734];
assign g[43119] = a[14] & g[26735];
assign g[59502] = b[14] & g[26735];
assign g[43120] = a[14] & g[26736];
assign g[59503] = b[14] & g[26736];
assign g[43121] = a[14] & g[26737];
assign g[59504] = b[14] & g[26737];
assign g[43122] = a[14] & g[26738];
assign g[59505] = b[14] & g[26738];
assign g[43123] = a[14] & g[26739];
assign g[59506] = b[14] & g[26739];
assign g[43124] = a[14] & g[26740];
assign g[59507] = b[14] & g[26740];
assign g[43125] = a[14] & g[26741];
assign g[59508] = b[14] & g[26741];
assign g[43126] = a[14] & g[26742];
assign g[59509] = b[14] & g[26742];
assign g[43127] = a[14] & g[26743];
assign g[59510] = b[14] & g[26743];
assign g[43128] = a[14] & g[26744];
assign g[59511] = b[14] & g[26744];
assign g[43129] = a[14] & g[26745];
assign g[59512] = b[14] & g[26745];
assign g[43130] = a[14] & g[26746];
assign g[59513] = b[14] & g[26746];
assign g[43131] = a[14] & g[26747];
assign g[59514] = b[14] & g[26747];
assign g[43132] = a[14] & g[26748];
assign g[59515] = b[14] & g[26748];
assign g[43133] = a[14] & g[26749];
assign g[59516] = b[14] & g[26749];
assign g[43134] = a[14] & g[26750];
assign g[59517] = b[14] & g[26750];
assign g[43135] = a[14] & g[26751];
assign g[59518] = b[14] & g[26751];
assign g[43136] = a[14] & g[26752];
assign g[59519] = b[14] & g[26752];
assign g[43137] = a[14] & g[26753];
assign g[59520] = b[14] & g[26753];
assign g[43138] = a[14] & g[26754];
assign g[59521] = b[14] & g[26754];
assign g[43139] = a[14] & g[26755];
assign g[59522] = b[14] & g[26755];
assign g[43140] = a[14] & g[26756];
assign g[59523] = b[14] & g[26756];
assign g[43141] = a[14] & g[26757];
assign g[59524] = b[14] & g[26757];
assign g[43142] = a[14] & g[26758];
assign g[59525] = b[14] & g[26758];
assign g[43143] = a[14] & g[26759];
assign g[59526] = b[14] & g[26759];
assign g[43144] = a[14] & g[26760];
assign g[59527] = b[14] & g[26760];
assign g[43145] = a[14] & g[26761];
assign g[59528] = b[14] & g[26761];
assign g[43146] = a[14] & g[26762];
assign g[59529] = b[14] & g[26762];
assign g[43147] = a[14] & g[26763];
assign g[59530] = b[14] & g[26763];
assign g[43148] = a[14] & g[26764];
assign g[59531] = b[14] & g[26764];
assign g[43149] = a[14] & g[26765];
assign g[59532] = b[14] & g[26765];
assign g[43150] = a[14] & g[26766];
assign g[59533] = b[14] & g[26766];
assign g[43151] = a[14] & g[26767];
assign g[59534] = b[14] & g[26767];
assign g[43152] = a[14] & g[26768];
assign g[59535] = b[14] & g[26768];
assign g[43153] = a[14] & g[26769];
assign g[59536] = b[14] & g[26769];
assign g[43154] = a[14] & g[26770];
assign g[59537] = b[14] & g[26770];
assign g[43155] = a[14] & g[26771];
assign g[59538] = b[14] & g[26771];
assign g[43156] = a[14] & g[26772];
assign g[59539] = b[14] & g[26772];
assign g[43157] = a[14] & g[26773];
assign g[59540] = b[14] & g[26773];
assign g[43158] = a[14] & g[26774];
assign g[59541] = b[14] & g[26774];
assign g[43159] = a[14] & g[26775];
assign g[59542] = b[14] & g[26775];
assign g[43160] = a[14] & g[26776];
assign g[59543] = b[14] & g[26776];
assign g[43161] = a[14] & g[26777];
assign g[59544] = b[14] & g[26777];
assign g[43162] = a[14] & g[26778];
assign g[59545] = b[14] & g[26778];
assign g[43163] = a[14] & g[26779];
assign g[59546] = b[14] & g[26779];
assign g[43164] = a[14] & g[26780];
assign g[59547] = b[14] & g[26780];
assign g[43165] = a[14] & g[26781];
assign g[59548] = b[14] & g[26781];
assign g[43166] = a[14] & g[26782];
assign g[59549] = b[14] & g[26782];
assign g[43167] = a[14] & g[26783];
assign g[59550] = b[14] & g[26783];
assign g[43168] = a[14] & g[26784];
assign g[59551] = b[14] & g[26784];
assign g[43169] = a[14] & g[26785];
assign g[59552] = b[14] & g[26785];
assign g[43170] = a[14] & g[26786];
assign g[59553] = b[14] & g[26786];
assign g[43171] = a[14] & g[26787];
assign g[59554] = b[14] & g[26787];
assign g[43172] = a[14] & g[26788];
assign g[59555] = b[14] & g[26788];
assign g[43173] = a[14] & g[26789];
assign g[59556] = b[14] & g[26789];
assign g[43174] = a[14] & g[26790];
assign g[59557] = b[14] & g[26790];
assign g[43175] = a[14] & g[26791];
assign g[59558] = b[14] & g[26791];
assign g[43176] = a[14] & g[26792];
assign g[59559] = b[14] & g[26792];
assign g[43177] = a[14] & g[26793];
assign g[59560] = b[14] & g[26793];
assign g[43178] = a[14] & g[26794];
assign g[59561] = b[14] & g[26794];
assign g[43179] = a[14] & g[26795];
assign g[59562] = b[14] & g[26795];
assign g[43180] = a[14] & g[26796];
assign g[59563] = b[14] & g[26796];
assign g[43181] = a[14] & g[26797];
assign g[59564] = b[14] & g[26797];
assign g[43182] = a[14] & g[26798];
assign g[59565] = b[14] & g[26798];
assign g[43183] = a[14] & g[26799];
assign g[59566] = b[14] & g[26799];
assign g[43184] = a[14] & g[26800];
assign g[59567] = b[14] & g[26800];
assign g[43185] = a[14] & g[26801];
assign g[59568] = b[14] & g[26801];
assign g[43186] = a[14] & g[26802];
assign g[59569] = b[14] & g[26802];
assign g[43187] = a[14] & g[26803];
assign g[59570] = b[14] & g[26803];
assign g[43188] = a[14] & g[26804];
assign g[59571] = b[14] & g[26804];
assign g[43189] = a[14] & g[26805];
assign g[59572] = b[14] & g[26805];
assign g[43190] = a[14] & g[26806];
assign g[59573] = b[14] & g[26806];
assign g[43191] = a[14] & g[26807];
assign g[59574] = b[14] & g[26807];
assign g[43192] = a[14] & g[26808];
assign g[59575] = b[14] & g[26808];
assign g[43193] = a[14] & g[26809];
assign g[59576] = b[14] & g[26809];
assign g[43194] = a[14] & g[26810];
assign g[59577] = b[14] & g[26810];
assign g[43195] = a[14] & g[26811];
assign g[59578] = b[14] & g[26811];
assign g[43196] = a[14] & g[26812];
assign g[59579] = b[14] & g[26812];
assign g[43197] = a[14] & g[26813];
assign g[59580] = b[14] & g[26813];
assign g[43198] = a[14] & g[26814];
assign g[59581] = b[14] & g[26814];
assign g[43199] = a[14] & g[26815];
assign g[59582] = b[14] & g[26815];
assign g[43200] = a[14] & g[26816];
assign g[59583] = b[14] & g[26816];
assign g[43201] = a[14] & g[26817];
assign g[59584] = b[14] & g[26817];
assign g[43202] = a[14] & g[26818];
assign g[59585] = b[14] & g[26818];
assign g[43203] = a[14] & g[26819];
assign g[59586] = b[14] & g[26819];
assign g[43204] = a[14] & g[26820];
assign g[59587] = b[14] & g[26820];
assign g[43205] = a[14] & g[26821];
assign g[59588] = b[14] & g[26821];
assign g[43206] = a[14] & g[26822];
assign g[59589] = b[14] & g[26822];
assign g[43207] = a[14] & g[26823];
assign g[59590] = b[14] & g[26823];
assign g[43208] = a[14] & g[26824];
assign g[59591] = b[14] & g[26824];
assign g[43209] = a[14] & g[26825];
assign g[59592] = b[14] & g[26825];
assign g[43210] = a[14] & g[26826];
assign g[59593] = b[14] & g[26826];
assign g[43211] = a[14] & g[26827];
assign g[59594] = b[14] & g[26827];
assign g[43212] = a[14] & g[26828];
assign g[59595] = b[14] & g[26828];
assign g[43213] = a[14] & g[26829];
assign g[59596] = b[14] & g[26829];
assign g[43214] = a[14] & g[26830];
assign g[59597] = b[14] & g[26830];
assign g[43215] = a[14] & g[26831];
assign g[59598] = b[14] & g[26831];
assign g[43216] = a[14] & g[26832];
assign g[59599] = b[14] & g[26832];
assign g[43217] = a[14] & g[26833];
assign g[59600] = b[14] & g[26833];
assign g[43218] = a[14] & g[26834];
assign g[59601] = b[14] & g[26834];
assign g[43219] = a[14] & g[26835];
assign g[59602] = b[14] & g[26835];
assign g[43220] = a[14] & g[26836];
assign g[59603] = b[14] & g[26836];
assign g[43221] = a[14] & g[26837];
assign g[59604] = b[14] & g[26837];
assign g[43222] = a[14] & g[26838];
assign g[59605] = b[14] & g[26838];
assign g[43223] = a[14] & g[26839];
assign g[59606] = b[14] & g[26839];
assign g[43224] = a[14] & g[26840];
assign g[59607] = b[14] & g[26840];
assign g[43225] = a[14] & g[26841];
assign g[59608] = b[14] & g[26841];
assign g[43226] = a[14] & g[26842];
assign g[59609] = b[14] & g[26842];
assign g[43227] = a[14] & g[26843];
assign g[59610] = b[14] & g[26843];
assign g[43228] = a[14] & g[26844];
assign g[59611] = b[14] & g[26844];
assign g[43229] = a[14] & g[26845];
assign g[59612] = b[14] & g[26845];
assign g[43230] = a[14] & g[26846];
assign g[59613] = b[14] & g[26846];
assign g[43231] = a[14] & g[26847];
assign g[59614] = b[14] & g[26847];
assign g[43232] = a[14] & g[26848];
assign g[59615] = b[14] & g[26848];
assign g[43233] = a[14] & g[26849];
assign g[59616] = b[14] & g[26849];
assign g[43234] = a[14] & g[26850];
assign g[59617] = b[14] & g[26850];
assign g[43235] = a[14] & g[26851];
assign g[59618] = b[14] & g[26851];
assign g[43236] = a[14] & g[26852];
assign g[59619] = b[14] & g[26852];
assign g[43237] = a[14] & g[26853];
assign g[59620] = b[14] & g[26853];
assign g[43238] = a[14] & g[26854];
assign g[59621] = b[14] & g[26854];
assign g[43239] = a[14] & g[26855];
assign g[59622] = b[14] & g[26855];
assign g[43240] = a[14] & g[26856];
assign g[59623] = b[14] & g[26856];
assign g[43241] = a[14] & g[26857];
assign g[59624] = b[14] & g[26857];
assign g[43242] = a[14] & g[26858];
assign g[59625] = b[14] & g[26858];
assign g[43243] = a[14] & g[26859];
assign g[59626] = b[14] & g[26859];
assign g[43244] = a[14] & g[26860];
assign g[59627] = b[14] & g[26860];
assign g[43245] = a[14] & g[26861];
assign g[59628] = b[14] & g[26861];
assign g[43246] = a[14] & g[26862];
assign g[59629] = b[14] & g[26862];
assign g[43247] = a[14] & g[26863];
assign g[59630] = b[14] & g[26863];
assign g[43248] = a[14] & g[26864];
assign g[59631] = b[14] & g[26864];
assign g[43249] = a[14] & g[26865];
assign g[59632] = b[14] & g[26865];
assign g[43250] = a[14] & g[26866];
assign g[59633] = b[14] & g[26866];
assign g[43251] = a[14] & g[26867];
assign g[59634] = b[14] & g[26867];
assign g[43252] = a[14] & g[26868];
assign g[59635] = b[14] & g[26868];
assign g[43253] = a[14] & g[26869];
assign g[59636] = b[14] & g[26869];
assign g[43254] = a[14] & g[26870];
assign g[59637] = b[14] & g[26870];
assign g[43255] = a[14] & g[26871];
assign g[59638] = b[14] & g[26871];
assign g[43256] = a[14] & g[26872];
assign g[59639] = b[14] & g[26872];
assign g[43257] = a[14] & g[26873];
assign g[59640] = b[14] & g[26873];
assign g[43258] = a[14] & g[26874];
assign g[59641] = b[14] & g[26874];
assign g[43259] = a[14] & g[26875];
assign g[59642] = b[14] & g[26875];
assign g[43260] = a[14] & g[26876];
assign g[59643] = b[14] & g[26876];
assign g[43261] = a[14] & g[26877];
assign g[59644] = b[14] & g[26877];
assign g[43262] = a[14] & g[26878];
assign g[59645] = b[14] & g[26878];
assign g[43263] = a[14] & g[26879];
assign g[59646] = b[14] & g[26879];
assign g[43264] = a[14] & g[26880];
assign g[59647] = b[14] & g[26880];
assign g[43265] = a[14] & g[26881];
assign g[59648] = b[14] & g[26881];
assign g[43266] = a[14] & g[26882];
assign g[59649] = b[14] & g[26882];
assign g[43267] = a[14] & g[26883];
assign g[59650] = b[14] & g[26883];
assign g[43268] = a[14] & g[26884];
assign g[59651] = b[14] & g[26884];
assign g[43269] = a[14] & g[26885];
assign g[59652] = b[14] & g[26885];
assign g[43270] = a[14] & g[26886];
assign g[59653] = b[14] & g[26886];
assign g[43271] = a[14] & g[26887];
assign g[59654] = b[14] & g[26887];
assign g[43272] = a[14] & g[26888];
assign g[59655] = b[14] & g[26888];
assign g[43273] = a[14] & g[26889];
assign g[59656] = b[14] & g[26889];
assign g[43274] = a[14] & g[26890];
assign g[59657] = b[14] & g[26890];
assign g[43275] = a[14] & g[26891];
assign g[59658] = b[14] & g[26891];
assign g[43276] = a[14] & g[26892];
assign g[59659] = b[14] & g[26892];
assign g[43277] = a[14] & g[26893];
assign g[59660] = b[14] & g[26893];
assign g[43278] = a[14] & g[26894];
assign g[59661] = b[14] & g[26894];
assign g[43279] = a[14] & g[26895];
assign g[59662] = b[14] & g[26895];
assign g[43280] = a[14] & g[26896];
assign g[59663] = b[14] & g[26896];
assign g[43281] = a[14] & g[26897];
assign g[59664] = b[14] & g[26897];
assign g[43282] = a[14] & g[26898];
assign g[59665] = b[14] & g[26898];
assign g[43283] = a[14] & g[26899];
assign g[59666] = b[14] & g[26899];
assign g[43284] = a[14] & g[26900];
assign g[59667] = b[14] & g[26900];
assign g[43285] = a[14] & g[26901];
assign g[59668] = b[14] & g[26901];
assign g[43286] = a[14] & g[26902];
assign g[59669] = b[14] & g[26902];
assign g[43287] = a[14] & g[26903];
assign g[59670] = b[14] & g[26903];
assign g[43288] = a[14] & g[26904];
assign g[59671] = b[14] & g[26904];
assign g[43289] = a[14] & g[26905];
assign g[59672] = b[14] & g[26905];
assign g[43290] = a[14] & g[26906];
assign g[59673] = b[14] & g[26906];
assign g[43291] = a[14] & g[26907];
assign g[59674] = b[14] & g[26907];
assign g[43292] = a[14] & g[26908];
assign g[59675] = b[14] & g[26908];
assign g[43293] = a[14] & g[26909];
assign g[59676] = b[14] & g[26909];
assign g[43294] = a[14] & g[26910];
assign g[59677] = b[14] & g[26910];
assign g[43295] = a[14] & g[26911];
assign g[59678] = b[14] & g[26911];
assign g[43296] = a[14] & g[26912];
assign g[59679] = b[14] & g[26912];
assign g[43297] = a[14] & g[26913];
assign g[59680] = b[14] & g[26913];
assign g[43298] = a[14] & g[26914];
assign g[59681] = b[14] & g[26914];
assign g[43299] = a[14] & g[26915];
assign g[59682] = b[14] & g[26915];
assign g[43300] = a[14] & g[26916];
assign g[59683] = b[14] & g[26916];
assign g[43301] = a[14] & g[26917];
assign g[59684] = b[14] & g[26917];
assign g[43302] = a[14] & g[26918];
assign g[59685] = b[14] & g[26918];
assign g[43303] = a[14] & g[26919];
assign g[59686] = b[14] & g[26919];
assign g[43304] = a[14] & g[26920];
assign g[59687] = b[14] & g[26920];
assign g[43305] = a[14] & g[26921];
assign g[59688] = b[14] & g[26921];
assign g[43306] = a[14] & g[26922];
assign g[59689] = b[14] & g[26922];
assign g[43307] = a[14] & g[26923];
assign g[59690] = b[14] & g[26923];
assign g[43308] = a[14] & g[26924];
assign g[59691] = b[14] & g[26924];
assign g[43309] = a[14] & g[26925];
assign g[59692] = b[14] & g[26925];
assign g[43310] = a[14] & g[26926];
assign g[59693] = b[14] & g[26926];
assign g[43311] = a[14] & g[26927];
assign g[59694] = b[14] & g[26927];
assign g[43312] = a[14] & g[26928];
assign g[59695] = b[14] & g[26928];
assign g[43313] = a[14] & g[26929];
assign g[59696] = b[14] & g[26929];
assign g[43314] = a[14] & g[26930];
assign g[59697] = b[14] & g[26930];
assign g[43315] = a[14] & g[26931];
assign g[59698] = b[14] & g[26931];
assign g[43316] = a[14] & g[26932];
assign g[59699] = b[14] & g[26932];
assign g[43317] = a[14] & g[26933];
assign g[59700] = b[14] & g[26933];
assign g[43318] = a[14] & g[26934];
assign g[59701] = b[14] & g[26934];
assign g[43319] = a[14] & g[26935];
assign g[59702] = b[14] & g[26935];
assign g[43320] = a[14] & g[26936];
assign g[59703] = b[14] & g[26936];
assign g[43321] = a[14] & g[26937];
assign g[59704] = b[14] & g[26937];
assign g[43322] = a[14] & g[26938];
assign g[59705] = b[14] & g[26938];
assign g[43323] = a[14] & g[26939];
assign g[59706] = b[14] & g[26939];
assign g[43324] = a[14] & g[26940];
assign g[59707] = b[14] & g[26940];
assign g[43325] = a[14] & g[26941];
assign g[59708] = b[14] & g[26941];
assign g[43326] = a[14] & g[26942];
assign g[59709] = b[14] & g[26942];
assign g[43327] = a[14] & g[26943];
assign g[59710] = b[14] & g[26943];
assign g[43328] = a[14] & g[26944];
assign g[59711] = b[14] & g[26944];
assign g[43329] = a[14] & g[26945];
assign g[59712] = b[14] & g[26945];
assign g[43330] = a[14] & g[26946];
assign g[59713] = b[14] & g[26946];
assign g[43331] = a[14] & g[26947];
assign g[59714] = b[14] & g[26947];
assign g[43332] = a[14] & g[26948];
assign g[59715] = b[14] & g[26948];
assign g[43333] = a[14] & g[26949];
assign g[59716] = b[14] & g[26949];
assign g[43334] = a[14] & g[26950];
assign g[59717] = b[14] & g[26950];
assign g[43335] = a[14] & g[26951];
assign g[59718] = b[14] & g[26951];
assign g[43336] = a[14] & g[26952];
assign g[59719] = b[14] & g[26952];
assign g[43337] = a[14] & g[26953];
assign g[59720] = b[14] & g[26953];
assign g[43338] = a[14] & g[26954];
assign g[59721] = b[14] & g[26954];
assign g[43339] = a[14] & g[26955];
assign g[59722] = b[14] & g[26955];
assign g[43340] = a[14] & g[26956];
assign g[59723] = b[14] & g[26956];
assign g[43341] = a[14] & g[26957];
assign g[59724] = b[14] & g[26957];
assign g[43342] = a[14] & g[26958];
assign g[59725] = b[14] & g[26958];
assign g[43343] = a[14] & g[26959];
assign g[59726] = b[14] & g[26959];
assign g[43344] = a[14] & g[26960];
assign g[59727] = b[14] & g[26960];
assign g[43345] = a[14] & g[26961];
assign g[59728] = b[14] & g[26961];
assign g[43346] = a[14] & g[26962];
assign g[59729] = b[14] & g[26962];
assign g[43347] = a[14] & g[26963];
assign g[59730] = b[14] & g[26963];
assign g[43348] = a[14] & g[26964];
assign g[59731] = b[14] & g[26964];
assign g[43349] = a[14] & g[26965];
assign g[59732] = b[14] & g[26965];
assign g[43350] = a[14] & g[26966];
assign g[59733] = b[14] & g[26966];
assign g[43351] = a[14] & g[26967];
assign g[59734] = b[14] & g[26967];
assign g[43352] = a[14] & g[26968];
assign g[59735] = b[14] & g[26968];
assign g[43353] = a[14] & g[26969];
assign g[59736] = b[14] & g[26969];
assign g[43354] = a[14] & g[26970];
assign g[59737] = b[14] & g[26970];
assign g[43355] = a[14] & g[26971];
assign g[59738] = b[14] & g[26971];
assign g[43356] = a[14] & g[26972];
assign g[59739] = b[14] & g[26972];
assign g[43357] = a[14] & g[26973];
assign g[59740] = b[14] & g[26973];
assign g[43358] = a[14] & g[26974];
assign g[59741] = b[14] & g[26974];
assign g[43359] = a[14] & g[26975];
assign g[59742] = b[14] & g[26975];
assign g[43360] = a[14] & g[26976];
assign g[59743] = b[14] & g[26976];
assign g[43361] = a[14] & g[26977];
assign g[59744] = b[14] & g[26977];
assign g[43362] = a[14] & g[26978];
assign g[59745] = b[14] & g[26978];
assign g[43363] = a[14] & g[26979];
assign g[59746] = b[14] & g[26979];
assign g[43364] = a[14] & g[26980];
assign g[59747] = b[14] & g[26980];
assign g[43365] = a[14] & g[26981];
assign g[59748] = b[14] & g[26981];
assign g[43366] = a[14] & g[26982];
assign g[59749] = b[14] & g[26982];
assign g[43367] = a[14] & g[26983];
assign g[59750] = b[14] & g[26983];
assign g[43368] = a[14] & g[26984];
assign g[59751] = b[14] & g[26984];
assign g[43369] = a[14] & g[26985];
assign g[59752] = b[14] & g[26985];
assign g[43370] = a[14] & g[26986];
assign g[59753] = b[14] & g[26986];
assign g[43371] = a[14] & g[26987];
assign g[59754] = b[14] & g[26987];
assign g[43372] = a[14] & g[26988];
assign g[59755] = b[14] & g[26988];
assign g[43373] = a[14] & g[26989];
assign g[59756] = b[14] & g[26989];
assign g[43374] = a[14] & g[26990];
assign g[59757] = b[14] & g[26990];
assign g[43375] = a[14] & g[26991];
assign g[59758] = b[14] & g[26991];
assign g[43376] = a[14] & g[26992];
assign g[59759] = b[14] & g[26992];
assign g[43377] = a[14] & g[26993];
assign g[59760] = b[14] & g[26993];
assign g[43378] = a[14] & g[26994];
assign g[59761] = b[14] & g[26994];
assign g[43379] = a[14] & g[26995];
assign g[59762] = b[14] & g[26995];
assign g[43380] = a[14] & g[26996];
assign g[59763] = b[14] & g[26996];
assign g[43381] = a[14] & g[26997];
assign g[59764] = b[14] & g[26997];
assign g[43382] = a[14] & g[26998];
assign g[59765] = b[14] & g[26998];
assign g[43383] = a[14] & g[26999];
assign g[59766] = b[14] & g[26999];
assign g[43384] = a[14] & g[27000];
assign g[59767] = b[14] & g[27000];
assign g[43385] = a[14] & g[27001];
assign g[59768] = b[14] & g[27001];
assign g[43386] = a[14] & g[27002];
assign g[59769] = b[14] & g[27002];
assign g[43387] = a[14] & g[27003];
assign g[59770] = b[14] & g[27003];
assign g[43388] = a[14] & g[27004];
assign g[59771] = b[14] & g[27004];
assign g[43389] = a[14] & g[27005];
assign g[59772] = b[14] & g[27005];
assign g[43390] = a[14] & g[27006];
assign g[59773] = b[14] & g[27006];
assign g[43391] = a[14] & g[27007];
assign g[59774] = b[14] & g[27007];
assign g[43392] = a[14] & g[27008];
assign g[59775] = b[14] & g[27008];
assign g[43393] = a[14] & g[27009];
assign g[59776] = b[14] & g[27009];
assign g[43394] = a[14] & g[27010];
assign g[59777] = b[14] & g[27010];
assign g[43395] = a[14] & g[27011];
assign g[59778] = b[14] & g[27011];
assign g[43396] = a[14] & g[27012];
assign g[59779] = b[14] & g[27012];
assign g[43397] = a[14] & g[27013];
assign g[59780] = b[14] & g[27013];
assign g[43398] = a[14] & g[27014];
assign g[59781] = b[14] & g[27014];
assign g[43399] = a[14] & g[27015];
assign g[59782] = b[14] & g[27015];
assign g[43400] = a[14] & g[27016];
assign g[59783] = b[14] & g[27016];
assign g[43401] = a[14] & g[27017];
assign g[59784] = b[14] & g[27017];
assign g[43402] = a[14] & g[27018];
assign g[59785] = b[14] & g[27018];
assign g[43403] = a[14] & g[27019];
assign g[59786] = b[14] & g[27019];
assign g[43404] = a[14] & g[27020];
assign g[59787] = b[14] & g[27020];
assign g[43405] = a[14] & g[27021];
assign g[59788] = b[14] & g[27021];
assign g[43406] = a[14] & g[27022];
assign g[59789] = b[14] & g[27022];
assign g[43407] = a[14] & g[27023];
assign g[59790] = b[14] & g[27023];
assign g[43408] = a[14] & g[27024];
assign g[59791] = b[14] & g[27024];
assign g[43409] = a[14] & g[27025];
assign g[59792] = b[14] & g[27025];
assign g[43410] = a[14] & g[27026];
assign g[59793] = b[14] & g[27026];
assign g[43411] = a[14] & g[27027];
assign g[59794] = b[14] & g[27027];
assign g[43412] = a[14] & g[27028];
assign g[59795] = b[14] & g[27028];
assign g[43413] = a[14] & g[27029];
assign g[59796] = b[14] & g[27029];
assign g[43414] = a[14] & g[27030];
assign g[59797] = b[14] & g[27030];
assign g[43415] = a[14] & g[27031];
assign g[59798] = b[14] & g[27031];
assign g[43416] = a[14] & g[27032];
assign g[59799] = b[14] & g[27032];
assign g[43417] = a[14] & g[27033];
assign g[59800] = b[14] & g[27033];
assign g[43418] = a[14] & g[27034];
assign g[59801] = b[14] & g[27034];
assign g[43419] = a[14] & g[27035];
assign g[59802] = b[14] & g[27035];
assign g[43420] = a[14] & g[27036];
assign g[59803] = b[14] & g[27036];
assign g[43421] = a[14] & g[27037];
assign g[59804] = b[14] & g[27037];
assign g[43422] = a[14] & g[27038];
assign g[59805] = b[14] & g[27038];
assign g[43423] = a[14] & g[27039];
assign g[59806] = b[14] & g[27039];
assign g[43424] = a[14] & g[27040];
assign g[59807] = b[14] & g[27040];
assign g[43425] = a[14] & g[27041];
assign g[59808] = b[14] & g[27041];
assign g[43426] = a[14] & g[27042];
assign g[59809] = b[14] & g[27042];
assign g[43427] = a[14] & g[27043];
assign g[59810] = b[14] & g[27043];
assign g[43428] = a[14] & g[27044];
assign g[59811] = b[14] & g[27044];
assign g[43429] = a[14] & g[27045];
assign g[59812] = b[14] & g[27045];
assign g[43430] = a[14] & g[27046];
assign g[59813] = b[14] & g[27046];
assign g[43431] = a[14] & g[27047];
assign g[59814] = b[14] & g[27047];
assign g[43432] = a[14] & g[27048];
assign g[59815] = b[14] & g[27048];
assign g[43433] = a[14] & g[27049];
assign g[59816] = b[14] & g[27049];
assign g[43434] = a[14] & g[27050];
assign g[59817] = b[14] & g[27050];
assign g[43435] = a[14] & g[27051];
assign g[59818] = b[14] & g[27051];
assign g[43436] = a[14] & g[27052];
assign g[59819] = b[14] & g[27052];
assign g[43437] = a[14] & g[27053];
assign g[59820] = b[14] & g[27053];
assign g[43438] = a[14] & g[27054];
assign g[59821] = b[14] & g[27054];
assign g[43439] = a[14] & g[27055];
assign g[59822] = b[14] & g[27055];
assign g[43440] = a[14] & g[27056];
assign g[59823] = b[14] & g[27056];
assign g[43441] = a[14] & g[27057];
assign g[59824] = b[14] & g[27057];
assign g[43442] = a[14] & g[27058];
assign g[59825] = b[14] & g[27058];
assign g[43443] = a[14] & g[27059];
assign g[59826] = b[14] & g[27059];
assign g[43444] = a[14] & g[27060];
assign g[59827] = b[14] & g[27060];
assign g[43445] = a[14] & g[27061];
assign g[59828] = b[14] & g[27061];
assign g[43446] = a[14] & g[27062];
assign g[59829] = b[14] & g[27062];
assign g[43447] = a[14] & g[27063];
assign g[59830] = b[14] & g[27063];
assign g[43448] = a[14] & g[27064];
assign g[59831] = b[14] & g[27064];
assign g[43449] = a[14] & g[27065];
assign g[59832] = b[14] & g[27065];
assign g[43450] = a[14] & g[27066];
assign g[59833] = b[14] & g[27066];
assign g[43451] = a[14] & g[27067];
assign g[59834] = b[14] & g[27067];
assign g[43452] = a[14] & g[27068];
assign g[59835] = b[14] & g[27068];
assign g[43453] = a[14] & g[27069];
assign g[59836] = b[14] & g[27069];
assign g[43454] = a[14] & g[27070];
assign g[59837] = b[14] & g[27070];
assign g[43455] = a[14] & g[27071];
assign g[59838] = b[14] & g[27071];
assign g[43456] = a[14] & g[27072];
assign g[59839] = b[14] & g[27072];
assign g[43457] = a[14] & g[27073];
assign g[59840] = b[14] & g[27073];
assign g[43458] = a[14] & g[27074];
assign g[59841] = b[14] & g[27074];
assign g[43459] = a[14] & g[27075];
assign g[59842] = b[14] & g[27075];
assign g[43460] = a[14] & g[27076];
assign g[59843] = b[14] & g[27076];
assign g[43461] = a[14] & g[27077];
assign g[59844] = b[14] & g[27077];
assign g[43462] = a[14] & g[27078];
assign g[59845] = b[14] & g[27078];
assign g[43463] = a[14] & g[27079];
assign g[59846] = b[14] & g[27079];
assign g[43464] = a[14] & g[27080];
assign g[59847] = b[14] & g[27080];
assign g[43465] = a[14] & g[27081];
assign g[59848] = b[14] & g[27081];
assign g[43466] = a[14] & g[27082];
assign g[59849] = b[14] & g[27082];
assign g[43467] = a[14] & g[27083];
assign g[59850] = b[14] & g[27083];
assign g[43468] = a[14] & g[27084];
assign g[59851] = b[14] & g[27084];
assign g[43469] = a[14] & g[27085];
assign g[59852] = b[14] & g[27085];
assign g[43470] = a[14] & g[27086];
assign g[59853] = b[14] & g[27086];
assign g[43471] = a[14] & g[27087];
assign g[59854] = b[14] & g[27087];
assign g[43472] = a[14] & g[27088];
assign g[59855] = b[14] & g[27088];
assign g[43473] = a[14] & g[27089];
assign g[59856] = b[14] & g[27089];
assign g[43474] = a[14] & g[27090];
assign g[59857] = b[14] & g[27090];
assign g[43475] = a[14] & g[27091];
assign g[59858] = b[14] & g[27091];
assign g[43476] = a[14] & g[27092];
assign g[59859] = b[14] & g[27092];
assign g[43477] = a[14] & g[27093];
assign g[59860] = b[14] & g[27093];
assign g[43478] = a[14] & g[27094];
assign g[59861] = b[14] & g[27094];
assign g[43479] = a[14] & g[27095];
assign g[59862] = b[14] & g[27095];
assign g[43480] = a[14] & g[27096];
assign g[59863] = b[14] & g[27096];
assign g[43481] = a[14] & g[27097];
assign g[59864] = b[14] & g[27097];
assign g[43482] = a[14] & g[27098];
assign g[59865] = b[14] & g[27098];
assign g[43483] = a[14] & g[27099];
assign g[59866] = b[14] & g[27099];
assign g[43484] = a[14] & g[27100];
assign g[59867] = b[14] & g[27100];
assign g[43485] = a[14] & g[27101];
assign g[59868] = b[14] & g[27101];
assign g[43486] = a[14] & g[27102];
assign g[59869] = b[14] & g[27102];
assign g[43487] = a[14] & g[27103];
assign g[59870] = b[14] & g[27103];
assign g[43488] = a[14] & g[27104];
assign g[59871] = b[14] & g[27104];
assign g[43489] = a[14] & g[27105];
assign g[59872] = b[14] & g[27105];
assign g[43490] = a[14] & g[27106];
assign g[59873] = b[14] & g[27106];
assign g[43491] = a[14] & g[27107];
assign g[59874] = b[14] & g[27107];
assign g[43492] = a[14] & g[27108];
assign g[59875] = b[14] & g[27108];
assign g[43493] = a[14] & g[27109];
assign g[59876] = b[14] & g[27109];
assign g[43494] = a[14] & g[27110];
assign g[59877] = b[14] & g[27110];
assign g[43495] = a[14] & g[27111];
assign g[59878] = b[14] & g[27111];
assign g[43496] = a[14] & g[27112];
assign g[59879] = b[14] & g[27112];
assign g[43497] = a[14] & g[27113];
assign g[59880] = b[14] & g[27113];
assign g[43498] = a[14] & g[27114];
assign g[59881] = b[14] & g[27114];
assign g[43499] = a[14] & g[27115];
assign g[59882] = b[14] & g[27115];
assign g[43500] = a[14] & g[27116];
assign g[59883] = b[14] & g[27116];
assign g[43501] = a[14] & g[27117];
assign g[59884] = b[14] & g[27117];
assign g[43502] = a[14] & g[27118];
assign g[59885] = b[14] & g[27118];
assign g[43503] = a[14] & g[27119];
assign g[59886] = b[14] & g[27119];
assign g[43504] = a[14] & g[27120];
assign g[59887] = b[14] & g[27120];
assign g[43505] = a[14] & g[27121];
assign g[59888] = b[14] & g[27121];
assign g[43506] = a[14] & g[27122];
assign g[59889] = b[14] & g[27122];
assign g[43507] = a[14] & g[27123];
assign g[59890] = b[14] & g[27123];
assign g[43508] = a[14] & g[27124];
assign g[59891] = b[14] & g[27124];
assign g[43509] = a[14] & g[27125];
assign g[59892] = b[14] & g[27125];
assign g[43510] = a[14] & g[27126];
assign g[59893] = b[14] & g[27126];
assign g[43511] = a[14] & g[27127];
assign g[59894] = b[14] & g[27127];
assign g[43512] = a[14] & g[27128];
assign g[59895] = b[14] & g[27128];
assign g[43513] = a[14] & g[27129];
assign g[59896] = b[14] & g[27129];
assign g[43514] = a[14] & g[27130];
assign g[59897] = b[14] & g[27130];
assign g[43515] = a[14] & g[27131];
assign g[59898] = b[14] & g[27131];
assign g[43516] = a[14] & g[27132];
assign g[59899] = b[14] & g[27132];
assign g[43517] = a[14] & g[27133];
assign g[59900] = b[14] & g[27133];
assign g[43518] = a[14] & g[27134];
assign g[59901] = b[14] & g[27134];
assign g[43519] = a[14] & g[27135];
assign g[59902] = b[14] & g[27135];
assign g[43520] = a[14] & g[27136];
assign g[59903] = b[14] & g[27136];
assign g[43521] = a[14] & g[27137];
assign g[59904] = b[14] & g[27137];
assign g[43522] = a[14] & g[27138];
assign g[59905] = b[14] & g[27138];
assign g[43523] = a[14] & g[27139];
assign g[59906] = b[14] & g[27139];
assign g[43524] = a[14] & g[27140];
assign g[59907] = b[14] & g[27140];
assign g[43525] = a[14] & g[27141];
assign g[59908] = b[14] & g[27141];
assign g[43526] = a[14] & g[27142];
assign g[59909] = b[14] & g[27142];
assign g[43527] = a[14] & g[27143];
assign g[59910] = b[14] & g[27143];
assign g[43528] = a[14] & g[27144];
assign g[59911] = b[14] & g[27144];
assign g[43529] = a[14] & g[27145];
assign g[59912] = b[14] & g[27145];
assign g[43530] = a[14] & g[27146];
assign g[59913] = b[14] & g[27146];
assign g[43531] = a[14] & g[27147];
assign g[59914] = b[14] & g[27147];
assign g[43532] = a[14] & g[27148];
assign g[59915] = b[14] & g[27148];
assign g[43533] = a[14] & g[27149];
assign g[59916] = b[14] & g[27149];
assign g[43534] = a[14] & g[27150];
assign g[59917] = b[14] & g[27150];
assign g[43535] = a[14] & g[27151];
assign g[59918] = b[14] & g[27151];
assign g[43536] = a[14] & g[27152];
assign g[59919] = b[14] & g[27152];
assign g[43537] = a[14] & g[27153];
assign g[59920] = b[14] & g[27153];
assign g[43538] = a[14] & g[27154];
assign g[59921] = b[14] & g[27154];
assign g[43539] = a[14] & g[27155];
assign g[59922] = b[14] & g[27155];
assign g[43540] = a[14] & g[27156];
assign g[59923] = b[14] & g[27156];
assign g[43541] = a[14] & g[27157];
assign g[59924] = b[14] & g[27157];
assign g[43542] = a[14] & g[27158];
assign g[59925] = b[14] & g[27158];
assign g[43543] = a[14] & g[27159];
assign g[59926] = b[14] & g[27159];
assign g[43544] = a[14] & g[27160];
assign g[59927] = b[14] & g[27160];
assign g[43545] = a[14] & g[27161];
assign g[59928] = b[14] & g[27161];
assign g[43546] = a[14] & g[27162];
assign g[59929] = b[14] & g[27162];
assign g[43547] = a[14] & g[27163];
assign g[59930] = b[14] & g[27163];
assign g[43548] = a[14] & g[27164];
assign g[59931] = b[14] & g[27164];
assign g[43549] = a[14] & g[27165];
assign g[59932] = b[14] & g[27165];
assign g[43550] = a[14] & g[27166];
assign g[59933] = b[14] & g[27166];
assign g[43551] = a[14] & g[27167];
assign g[59934] = b[14] & g[27167];
assign g[43552] = a[14] & g[27168];
assign g[59935] = b[14] & g[27168];
assign g[43553] = a[14] & g[27169];
assign g[59936] = b[14] & g[27169];
assign g[43554] = a[14] & g[27170];
assign g[59937] = b[14] & g[27170];
assign g[43555] = a[14] & g[27171];
assign g[59938] = b[14] & g[27171];
assign g[43556] = a[14] & g[27172];
assign g[59939] = b[14] & g[27172];
assign g[43557] = a[14] & g[27173];
assign g[59940] = b[14] & g[27173];
assign g[43558] = a[14] & g[27174];
assign g[59941] = b[14] & g[27174];
assign g[43559] = a[14] & g[27175];
assign g[59942] = b[14] & g[27175];
assign g[43560] = a[14] & g[27176];
assign g[59943] = b[14] & g[27176];
assign g[43561] = a[14] & g[27177];
assign g[59944] = b[14] & g[27177];
assign g[43562] = a[14] & g[27178];
assign g[59945] = b[14] & g[27178];
assign g[43563] = a[14] & g[27179];
assign g[59946] = b[14] & g[27179];
assign g[43564] = a[14] & g[27180];
assign g[59947] = b[14] & g[27180];
assign g[43565] = a[14] & g[27181];
assign g[59948] = b[14] & g[27181];
assign g[43566] = a[14] & g[27182];
assign g[59949] = b[14] & g[27182];
assign g[43567] = a[14] & g[27183];
assign g[59950] = b[14] & g[27183];
assign g[43568] = a[14] & g[27184];
assign g[59951] = b[14] & g[27184];
assign g[43569] = a[14] & g[27185];
assign g[59952] = b[14] & g[27185];
assign g[43570] = a[14] & g[27186];
assign g[59953] = b[14] & g[27186];
assign g[43571] = a[14] & g[27187];
assign g[59954] = b[14] & g[27187];
assign g[43572] = a[14] & g[27188];
assign g[59955] = b[14] & g[27188];
assign g[43573] = a[14] & g[27189];
assign g[59956] = b[14] & g[27189];
assign g[43574] = a[14] & g[27190];
assign g[59957] = b[14] & g[27190];
assign g[43575] = a[14] & g[27191];
assign g[59958] = b[14] & g[27191];
assign g[43576] = a[14] & g[27192];
assign g[59959] = b[14] & g[27192];
assign g[43577] = a[14] & g[27193];
assign g[59960] = b[14] & g[27193];
assign g[43578] = a[14] & g[27194];
assign g[59961] = b[14] & g[27194];
assign g[43579] = a[14] & g[27195];
assign g[59962] = b[14] & g[27195];
assign g[43580] = a[14] & g[27196];
assign g[59963] = b[14] & g[27196];
assign g[43581] = a[14] & g[27197];
assign g[59964] = b[14] & g[27197];
assign g[43582] = a[14] & g[27198];
assign g[59965] = b[14] & g[27198];
assign g[43583] = a[14] & g[27199];
assign g[59966] = b[14] & g[27199];
assign g[43584] = a[14] & g[27200];
assign g[59967] = b[14] & g[27200];
assign g[43585] = a[14] & g[27201];
assign g[59968] = b[14] & g[27201];
assign g[43586] = a[14] & g[27202];
assign g[59969] = b[14] & g[27202];
assign g[43587] = a[14] & g[27203];
assign g[59970] = b[14] & g[27203];
assign g[43588] = a[14] & g[27204];
assign g[59971] = b[14] & g[27204];
assign g[43589] = a[14] & g[27205];
assign g[59972] = b[14] & g[27205];
assign g[43590] = a[14] & g[27206];
assign g[59973] = b[14] & g[27206];
assign g[43591] = a[14] & g[27207];
assign g[59974] = b[14] & g[27207];
assign g[43592] = a[14] & g[27208];
assign g[59975] = b[14] & g[27208];
assign g[43593] = a[14] & g[27209];
assign g[59976] = b[14] & g[27209];
assign g[43594] = a[14] & g[27210];
assign g[59977] = b[14] & g[27210];
assign g[43595] = a[14] & g[27211];
assign g[59978] = b[14] & g[27211];
assign g[43596] = a[14] & g[27212];
assign g[59979] = b[14] & g[27212];
assign g[43597] = a[14] & g[27213];
assign g[59980] = b[14] & g[27213];
assign g[43598] = a[14] & g[27214];
assign g[59981] = b[14] & g[27214];
assign g[43599] = a[14] & g[27215];
assign g[59982] = b[14] & g[27215];
assign g[43600] = a[14] & g[27216];
assign g[59983] = b[14] & g[27216];
assign g[43601] = a[14] & g[27217];
assign g[59984] = b[14] & g[27217];
assign g[43602] = a[14] & g[27218];
assign g[59985] = b[14] & g[27218];
assign g[43603] = a[14] & g[27219];
assign g[59986] = b[14] & g[27219];
assign g[43604] = a[14] & g[27220];
assign g[59987] = b[14] & g[27220];
assign g[43605] = a[14] & g[27221];
assign g[59988] = b[14] & g[27221];
assign g[43606] = a[14] & g[27222];
assign g[59989] = b[14] & g[27222];
assign g[43607] = a[14] & g[27223];
assign g[59990] = b[14] & g[27223];
assign g[43608] = a[14] & g[27224];
assign g[59991] = b[14] & g[27224];
assign g[43609] = a[14] & g[27225];
assign g[59992] = b[14] & g[27225];
assign g[43610] = a[14] & g[27226];
assign g[59993] = b[14] & g[27226];
assign g[43611] = a[14] & g[27227];
assign g[59994] = b[14] & g[27227];
assign g[43612] = a[14] & g[27228];
assign g[59995] = b[14] & g[27228];
assign g[43613] = a[14] & g[27229];
assign g[59996] = b[14] & g[27229];
assign g[43614] = a[14] & g[27230];
assign g[59997] = b[14] & g[27230];
assign g[43615] = a[14] & g[27231];
assign g[59998] = b[14] & g[27231];
assign g[43616] = a[14] & g[27232];
assign g[59999] = b[14] & g[27232];
assign g[43617] = a[14] & g[27233];
assign g[60000] = b[14] & g[27233];
assign g[43618] = a[14] & g[27234];
assign g[60001] = b[14] & g[27234];
assign g[43619] = a[14] & g[27235];
assign g[60002] = b[14] & g[27235];
assign g[43620] = a[14] & g[27236];
assign g[60003] = b[14] & g[27236];
assign g[43621] = a[14] & g[27237];
assign g[60004] = b[14] & g[27237];
assign g[43622] = a[14] & g[27238];
assign g[60005] = b[14] & g[27238];
assign g[43623] = a[14] & g[27239];
assign g[60006] = b[14] & g[27239];
assign g[43624] = a[14] & g[27240];
assign g[60007] = b[14] & g[27240];
assign g[43625] = a[14] & g[27241];
assign g[60008] = b[14] & g[27241];
assign g[43626] = a[14] & g[27242];
assign g[60009] = b[14] & g[27242];
assign g[43627] = a[14] & g[27243];
assign g[60010] = b[14] & g[27243];
assign g[43628] = a[14] & g[27244];
assign g[60011] = b[14] & g[27244];
assign g[43629] = a[14] & g[27245];
assign g[60012] = b[14] & g[27245];
assign g[43630] = a[14] & g[27246];
assign g[60013] = b[14] & g[27246];
assign g[43631] = a[14] & g[27247];
assign g[60014] = b[14] & g[27247];
assign g[43632] = a[14] & g[27248];
assign g[60015] = b[14] & g[27248];
assign g[43633] = a[14] & g[27249];
assign g[60016] = b[14] & g[27249];
assign g[43634] = a[14] & g[27250];
assign g[60017] = b[14] & g[27250];
assign g[43635] = a[14] & g[27251];
assign g[60018] = b[14] & g[27251];
assign g[43636] = a[14] & g[27252];
assign g[60019] = b[14] & g[27252];
assign g[43637] = a[14] & g[27253];
assign g[60020] = b[14] & g[27253];
assign g[43638] = a[14] & g[27254];
assign g[60021] = b[14] & g[27254];
assign g[43639] = a[14] & g[27255];
assign g[60022] = b[14] & g[27255];
assign g[43640] = a[14] & g[27256];
assign g[60023] = b[14] & g[27256];
assign g[43641] = a[14] & g[27257];
assign g[60024] = b[14] & g[27257];
assign g[43642] = a[14] & g[27258];
assign g[60025] = b[14] & g[27258];
assign g[43643] = a[14] & g[27259];
assign g[60026] = b[14] & g[27259];
assign g[43644] = a[14] & g[27260];
assign g[60027] = b[14] & g[27260];
assign g[43645] = a[14] & g[27261];
assign g[60028] = b[14] & g[27261];
assign g[43646] = a[14] & g[27262];
assign g[60029] = b[14] & g[27262];
assign g[43647] = a[14] & g[27263];
assign g[60030] = b[14] & g[27263];
assign g[43648] = a[14] & g[27264];
assign g[60031] = b[14] & g[27264];
assign g[43649] = a[14] & g[27265];
assign g[60032] = b[14] & g[27265];
assign g[43650] = a[14] & g[27266];
assign g[60033] = b[14] & g[27266];
assign g[43651] = a[14] & g[27267];
assign g[60034] = b[14] & g[27267];
assign g[43652] = a[14] & g[27268];
assign g[60035] = b[14] & g[27268];
assign g[43653] = a[14] & g[27269];
assign g[60036] = b[14] & g[27269];
assign g[43654] = a[14] & g[27270];
assign g[60037] = b[14] & g[27270];
assign g[43655] = a[14] & g[27271];
assign g[60038] = b[14] & g[27271];
assign g[43656] = a[14] & g[27272];
assign g[60039] = b[14] & g[27272];
assign g[43657] = a[14] & g[27273];
assign g[60040] = b[14] & g[27273];
assign g[43658] = a[14] & g[27274];
assign g[60041] = b[14] & g[27274];
assign g[43659] = a[14] & g[27275];
assign g[60042] = b[14] & g[27275];
assign g[43660] = a[14] & g[27276];
assign g[60043] = b[14] & g[27276];
assign g[43661] = a[14] & g[27277];
assign g[60044] = b[14] & g[27277];
assign g[43662] = a[14] & g[27278];
assign g[60045] = b[14] & g[27278];
assign g[43663] = a[14] & g[27279];
assign g[60046] = b[14] & g[27279];
assign g[43664] = a[14] & g[27280];
assign g[60047] = b[14] & g[27280];
assign g[43665] = a[14] & g[27281];
assign g[60048] = b[14] & g[27281];
assign g[43666] = a[14] & g[27282];
assign g[60049] = b[14] & g[27282];
assign g[43667] = a[14] & g[27283];
assign g[60050] = b[14] & g[27283];
assign g[43668] = a[14] & g[27284];
assign g[60051] = b[14] & g[27284];
assign g[43669] = a[14] & g[27285];
assign g[60052] = b[14] & g[27285];
assign g[43670] = a[14] & g[27286];
assign g[60053] = b[14] & g[27286];
assign g[43671] = a[14] & g[27287];
assign g[60054] = b[14] & g[27287];
assign g[43672] = a[14] & g[27288];
assign g[60055] = b[14] & g[27288];
assign g[43673] = a[14] & g[27289];
assign g[60056] = b[14] & g[27289];
assign g[43674] = a[14] & g[27290];
assign g[60057] = b[14] & g[27290];
assign g[43675] = a[14] & g[27291];
assign g[60058] = b[14] & g[27291];
assign g[43676] = a[14] & g[27292];
assign g[60059] = b[14] & g[27292];
assign g[43677] = a[14] & g[27293];
assign g[60060] = b[14] & g[27293];
assign g[43678] = a[14] & g[27294];
assign g[60061] = b[14] & g[27294];
assign g[43679] = a[14] & g[27295];
assign g[60062] = b[14] & g[27295];
assign g[43680] = a[14] & g[27296];
assign g[60063] = b[14] & g[27296];
assign g[43681] = a[14] & g[27297];
assign g[60064] = b[14] & g[27297];
assign g[43682] = a[14] & g[27298];
assign g[60065] = b[14] & g[27298];
assign g[43683] = a[14] & g[27299];
assign g[60066] = b[14] & g[27299];
assign g[43684] = a[14] & g[27300];
assign g[60067] = b[14] & g[27300];
assign g[43685] = a[14] & g[27301];
assign g[60068] = b[14] & g[27301];
assign g[43686] = a[14] & g[27302];
assign g[60069] = b[14] & g[27302];
assign g[43687] = a[14] & g[27303];
assign g[60070] = b[14] & g[27303];
assign g[43688] = a[14] & g[27304];
assign g[60071] = b[14] & g[27304];
assign g[43689] = a[14] & g[27305];
assign g[60072] = b[14] & g[27305];
assign g[43690] = a[14] & g[27306];
assign g[60073] = b[14] & g[27306];
assign g[43691] = a[14] & g[27307];
assign g[60074] = b[14] & g[27307];
assign g[43692] = a[14] & g[27308];
assign g[60075] = b[14] & g[27308];
assign g[43693] = a[14] & g[27309];
assign g[60076] = b[14] & g[27309];
assign g[43694] = a[14] & g[27310];
assign g[60077] = b[14] & g[27310];
assign g[43695] = a[14] & g[27311];
assign g[60078] = b[14] & g[27311];
assign g[43696] = a[14] & g[27312];
assign g[60079] = b[14] & g[27312];
assign g[43697] = a[14] & g[27313];
assign g[60080] = b[14] & g[27313];
assign g[43698] = a[14] & g[27314];
assign g[60081] = b[14] & g[27314];
assign g[43699] = a[14] & g[27315];
assign g[60082] = b[14] & g[27315];
assign g[43700] = a[14] & g[27316];
assign g[60083] = b[14] & g[27316];
assign g[43701] = a[14] & g[27317];
assign g[60084] = b[14] & g[27317];
assign g[43702] = a[14] & g[27318];
assign g[60085] = b[14] & g[27318];
assign g[43703] = a[14] & g[27319];
assign g[60086] = b[14] & g[27319];
assign g[43704] = a[14] & g[27320];
assign g[60087] = b[14] & g[27320];
assign g[43705] = a[14] & g[27321];
assign g[60088] = b[14] & g[27321];
assign g[43706] = a[14] & g[27322];
assign g[60089] = b[14] & g[27322];
assign g[43707] = a[14] & g[27323];
assign g[60090] = b[14] & g[27323];
assign g[43708] = a[14] & g[27324];
assign g[60091] = b[14] & g[27324];
assign g[43709] = a[14] & g[27325];
assign g[60092] = b[14] & g[27325];
assign g[43710] = a[14] & g[27326];
assign g[60093] = b[14] & g[27326];
assign g[43711] = a[14] & g[27327];
assign g[60094] = b[14] & g[27327];
assign g[43712] = a[14] & g[27328];
assign g[60095] = b[14] & g[27328];
assign g[43713] = a[14] & g[27329];
assign g[60096] = b[14] & g[27329];
assign g[43714] = a[14] & g[27330];
assign g[60097] = b[14] & g[27330];
assign g[43715] = a[14] & g[27331];
assign g[60098] = b[14] & g[27331];
assign g[43716] = a[14] & g[27332];
assign g[60099] = b[14] & g[27332];
assign g[43717] = a[14] & g[27333];
assign g[60100] = b[14] & g[27333];
assign g[43718] = a[14] & g[27334];
assign g[60101] = b[14] & g[27334];
assign g[43719] = a[14] & g[27335];
assign g[60102] = b[14] & g[27335];
assign g[43720] = a[14] & g[27336];
assign g[60103] = b[14] & g[27336];
assign g[43721] = a[14] & g[27337];
assign g[60104] = b[14] & g[27337];
assign g[43722] = a[14] & g[27338];
assign g[60105] = b[14] & g[27338];
assign g[43723] = a[14] & g[27339];
assign g[60106] = b[14] & g[27339];
assign g[43724] = a[14] & g[27340];
assign g[60107] = b[14] & g[27340];
assign g[43725] = a[14] & g[27341];
assign g[60108] = b[14] & g[27341];
assign g[43726] = a[14] & g[27342];
assign g[60109] = b[14] & g[27342];
assign g[43727] = a[14] & g[27343];
assign g[60110] = b[14] & g[27343];
assign g[43728] = a[14] & g[27344];
assign g[60111] = b[14] & g[27344];
assign g[43729] = a[14] & g[27345];
assign g[60112] = b[14] & g[27345];
assign g[43730] = a[14] & g[27346];
assign g[60113] = b[14] & g[27346];
assign g[43731] = a[14] & g[27347];
assign g[60114] = b[14] & g[27347];
assign g[43732] = a[14] & g[27348];
assign g[60115] = b[14] & g[27348];
assign g[43733] = a[14] & g[27349];
assign g[60116] = b[14] & g[27349];
assign g[43734] = a[14] & g[27350];
assign g[60117] = b[14] & g[27350];
assign g[43735] = a[14] & g[27351];
assign g[60118] = b[14] & g[27351];
assign g[43736] = a[14] & g[27352];
assign g[60119] = b[14] & g[27352];
assign g[43737] = a[14] & g[27353];
assign g[60120] = b[14] & g[27353];
assign g[43738] = a[14] & g[27354];
assign g[60121] = b[14] & g[27354];
assign g[43739] = a[14] & g[27355];
assign g[60122] = b[14] & g[27355];
assign g[43740] = a[14] & g[27356];
assign g[60123] = b[14] & g[27356];
assign g[43741] = a[14] & g[27357];
assign g[60124] = b[14] & g[27357];
assign g[43742] = a[14] & g[27358];
assign g[60125] = b[14] & g[27358];
assign g[43743] = a[14] & g[27359];
assign g[60126] = b[14] & g[27359];
assign g[43744] = a[14] & g[27360];
assign g[60127] = b[14] & g[27360];
assign g[43745] = a[14] & g[27361];
assign g[60128] = b[14] & g[27361];
assign g[43746] = a[14] & g[27362];
assign g[60129] = b[14] & g[27362];
assign g[43747] = a[14] & g[27363];
assign g[60130] = b[14] & g[27363];
assign g[43748] = a[14] & g[27364];
assign g[60131] = b[14] & g[27364];
assign g[43749] = a[14] & g[27365];
assign g[60132] = b[14] & g[27365];
assign g[43750] = a[14] & g[27366];
assign g[60133] = b[14] & g[27366];
assign g[43751] = a[14] & g[27367];
assign g[60134] = b[14] & g[27367];
assign g[43752] = a[14] & g[27368];
assign g[60135] = b[14] & g[27368];
assign g[43753] = a[14] & g[27369];
assign g[60136] = b[14] & g[27369];
assign g[43754] = a[14] & g[27370];
assign g[60137] = b[14] & g[27370];
assign g[43755] = a[14] & g[27371];
assign g[60138] = b[14] & g[27371];
assign g[43756] = a[14] & g[27372];
assign g[60139] = b[14] & g[27372];
assign g[43757] = a[14] & g[27373];
assign g[60140] = b[14] & g[27373];
assign g[43758] = a[14] & g[27374];
assign g[60141] = b[14] & g[27374];
assign g[43759] = a[14] & g[27375];
assign g[60142] = b[14] & g[27375];
assign g[43760] = a[14] & g[27376];
assign g[60143] = b[14] & g[27376];
assign g[43761] = a[14] & g[27377];
assign g[60144] = b[14] & g[27377];
assign g[43762] = a[14] & g[27378];
assign g[60145] = b[14] & g[27378];
assign g[43763] = a[14] & g[27379];
assign g[60146] = b[14] & g[27379];
assign g[43764] = a[14] & g[27380];
assign g[60147] = b[14] & g[27380];
assign g[43765] = a[14] & g[27381];
assign g[60148] = b[14] & g[27381];
assign g[43766] = a[14] & g[27382];
assign g[60149] = b[14] & g[27382];
assign g[43767] = a[14] & g[27383];
assign g[60150] = b[14] & g[27383];
assign g[43768] = a[14] & g[27384];
assign g[60151] = b[14] & g[27384];
assign g[43769] = a[14] & g[27385];
assign g[60152] = b[14] & g[27385];
assign g[43770] = a[14] & g[27386];
assign g[60153] = b[14] & g[27386];
assign g[43771] = a[14] & g[27387];
assign g[60154] = b[14] & g[27387];
assign g[43772] = a[14] & g[27388];
assign g[60155] = b[14] & g[27388];
assign g[43773] = a[14] & g[27389];
assign g[60156] = b[14] & g[27389];
assign g[43774] = a[14] & g[27390];
assign g[60157] = b[14] & g[27390];
assign g[43775] = a[14] & g[27391];
assign g[60158] = b[14] & g[27391];
assign g[43776] = a[14] & g[27392];
assign g[60159] = b[14] & g[27392];
assign g[43777] = a[14] & g[27393];
assign g[60160] = b[14] & g[27393];
assign g[43778] = a[14] & g[27394];
assign g[60161] = b[14] & g[27394];
assign g[43779] = a[14] & g[27395];
assign g[60162] = b[14] & g[27395];
assign g[43780] = a[14] & g[27396];
assign g[60163] = b[14] & g[27396];
assign g[43781] = a[14] & g[27397];
assign g[60164] = b[14] & g[27397];
assign g[43782] = a[14] & g[27398];
assign g[60165] = b[14] & g[27398];
assign g[43783] = a[14] & g[27399];
assign g[60166] = b[14] & g[27399];
assign g[43784] = a[14] & g[27400];
assign g[60167] = b[14] & g[27400];
assign g[43785] = a[14] & g[27401];
assign g[60168] = b[14] & g[27401];
assign g[43786] = a[14] & g[27402];
assign g[60169] = b[14] & g[27402];
assign g[43787] = a[14] & g[27403];
assign g[60170] = b[14] & g[27403];
assign g[43788] = a[14] & g[27404];
assign g[60171] = b[14] & g[27404];
assign g[43789] = a[14] & g[27405];
assign g[60172] = b[14] & g[27405];
assign g[43790] = a[14] & g[27406];
assign g[60173] = b[14] & g[27406];
assign g[43791] = a[14] & g[27407];
assign g[60174] = b[14] & g[27407];
assign g[43792] = a[14] & g[27408];
assign g[60175] = b[14] & g[27408];
assign g[43793] = a[14] & g[27409];
assign g[60176] = b[14] & g[27409];
assign g[43794] = a[14] & g[27410];
assign g[60177] = b[14] & g[27410];
assign g[43795] = a[14] & g[27411];
assign g[60178] = b[14] & g[27411];
assign g[43796] = a[14] & g[27412];
assign g[60179] = b[14] & g[27412];
assign g[43797] = a[14] & g[27413];
assign g[60180] = b[14] & g[27413];
assign g[43798] = a[14] & g[27414];
assign g[60181] = b[14] & g[27414];
assign g[43799] = a[14] & g[27415];
assign g[60182] = b[14] & g[27415];
assign g[43800] = a[14] & g[27416];
assign g[60183] = b[14] & g[27416];
assign g[43801] = a[14] & g[27417];
assign g[60184] = b[14] & g[27417];
assign g[43802] = a[14] & g[27418];
assign g[60185] = b[14] & g[27418];
assign g[43803] = a[14] & g[27419];
assign g[60186] = b[14] & g[27419];
assign g[43804] = a[14] & g[27420];
assign g[60187] = b[14] & g[27420];
assign g[43805] = a[14] & g[27421];
assign g[60188] = b[14] & g[27421];
assign g[43806] = a[14] & g[27422];
assign g[60189] = b[14] & g[27422];
assign g[43807] = a[14] & g[27423];
assign g[60190] = b[14] & g[27423];
assign g[43808] = a[14] & g[27424];
assign g[60191] = b[14] & g[27424];
assign g[43809] = a[14] & g[27425];
assign g[60192] = b[14] & g[27425];
assign g[43810] = a[14] & g[27426];
assign g[60193] = b[14] & g[27426];
assign g[43811] = a[14] & g[27427];
assign g[60194] = b[14] & g[27427];
assign g[43812] = a[14] & g[27428];
assign g[60195] = b[14] & g[27428];
assign g[43813] = a[14] & g[27429];
assign g[60196] = b[14] & g[27429];
assign g[43814] = a[14] & g[27430];
assign g[60197] = b[14] & g[27430];
assign g[43815] = a[14] & g[27431];
assign g[60198] = b[14] & g[27431];
assign g[43816] = a[14] & g[27432];
assign g[60199] = b[14] & g[27432];
assign g[43817] = a[14] & g[27433];
assign g[60200] = b[14] & g[27433];
assign g[43818] = a[14] & g[27434];
assign g[60201] = b[14] & g[27434];
assign g[43819] = a[14] & g[27435];
assign g[60202] = b[14] & g[27435];
assign g[43820] = a[14] & g[27436];
assign g[60203] = b[14] & g[27436];
assign g[43821] = a[14] & g[27437];
assign g[60204] = b[14] & g[27437];
assign g[43822] = a[14] & g[27438];
assign g[60205] = b[14] & g[27438];
assign g[43823] = a[14] & g[27439];
assign g[60206] = b[14] & g[27439];
assign g[43824] = a[14] & g[27440];
assign g[60207] = b[14] & g[27440];
assign g[43825] = a[14] & g[27441];
assign g[60208] = b[14] & g[27441];
assign g[43826] = a[14] & g[27442];
assign g[60209] = b[14] & g[27442];
assign g[43827] = a[14] & g[27443];
assign g[60210] = b[14] & g[27443];
assign g[43828] = a[14] & g[27444];
assign g[60211] = b[14] & g[27444];
assign g[43829] = a[14] & g[27445];
assign g[60212] = b[14] & g[27445];
assign g[43830] = a[14] & g[27446];
assign g[60213] = b[14] & g[27446];
assign g[43831] = a[14] & g[27447];
assign g[60214] = b[14] & g[27447];
assign g[43832] = a[14] & g[27448];
assign g[60215] = b[14] & g[27448];
assign g[43833] = a[14] & g[27449];
assign g[60216] = b[14] & g[27449];
assign g[43834] = a[14] & g[27450];
assign g[60217] = b[14] & g[27450];
assign g[43835] = a[14] & g[27451];
assign g[60218] = b[14] & g[27451];
assign g[43836] = a[14] & g[27452];
assign g[60219] = b[14] & g[27452];
assign g[43837] = a[14] & g[27453];
assign g[60220] = b[14] & g[27453];
assign g[43838] = a[14] & g[27454];
assign g[60221] = b[14] & g[27454];
assign g[43839] = a[14] & g[27455];
assign g[60222] = b[14] & g[27455];
assign g[43840] = a[14] & g[27456];
assign g[60223] = b[14] & g[27456];
assign g[43841] = a[14] & g[27457];
assign g[60224] = b[14] & g[27457];
assign g[43842] = a[14] & g[27458];
assign g[60225] = b[14] & g[27458];
assign g[43843] = a[14] & g[27459];
assign g[60226] = b[14] & g[27459];
assign g[43844] = a[14] & g[27460];
assign g[60227] = b[14] & g[27460];
assign g[43845] = a[14] & g[27461];
assign g[60228] = b[14] & g[27461];
assign g[43846] = a[14] & g[27462];
assign g[60229] = b[14] & g[27462];
assign g[43847] = a[14] & g[27463];
assign g[60230] = b[14] & g[27463];
assign g[43848] = a[14] & g[27464];
assign g[60231] = b[14] & g[27464];
assign g[43849] = a[14] & g[27465];
assign g[60232] = b[14] & g[27465];
assign g[43850] = a[14] & g[27466];
assign g[60233] = b[14] & g[27466];
assign g[43851] = a[14] & g[27467];
assign g[60234] = b[14] & g[27467];
assign g[43852] = a[14] & g[27468];
assign g[60235] = b[14] & g[27468];
assign g[43853] = a[14] & g[27469];
assign g[60236] = b[14] & g[27469];
assign g[43854] = a[14] & g[27470];
assign g[60237] = b[14] & g[27470];
assign g[43855] = a[14] & g[27471];
assign g[60238] = b[14] & g[27471];
assign g[43856] = a[14] & g[27472];
assign g[60239] = b[14] & g[27472];
assign g[43857] = a[14] & g[27473];
assign g[60240] = b[14] & g[27473];
assign g[43858] = a[14] & g[27474];
assign g[60241] = b[14] & g[27474];
assign g[43859] = a[14] & g[27475];
assign g[60242] = b[14] & g[27475];
assign g[43860] = a[14] & g[27476];
assign g[60243] = b[14] & g[27476];
assign g[43861] = a[14] & g[27477];
assign g[60244] = b[14] & g[27477];
assign g[43862] = a[14] & g[27478];
assign g[60245] = b[14] & g[27478];
assign g[43863] = a[14] & g[27479];
assign g[60246] = b[14] & g[27479];
assign g[43864] = a[14] & g[27480];
assign g[60247] = b[14] & g[27480];
assign g[43865] = a[14] & g[27481];
assign g[60248] = b[14] & g[27481];
assign g[43866] = a[14] & g[27482];
assign g[60249] = b[14] & g[27482];
assign g[43867] = a[14] & g[27483];
assign g[60250] = b[14] & g[27483];
assign g[43868] = a[14] & g[27484];
assign g[60251] = b[14] & g[27484];
assign g[43869] = a[14] & g[27485];
assign g[60252] = b[14] & g[27485];
assign g[43870] = a[14] & g[27486];
assign g[60253] = b[14] & g[27486];
assign g[43871] = a[14] & g[27487];
assign g[60254] = b[14] & g[27487];
assign g[43872] = a[14] & g[27488];
assign g[60255] = b[14] & g[27488];
assign g[43873] = a[14] & g[27489];
assign g[60256] = b[14] & g[27489];
assign g[43874] = a[14] & g[27490];
assign g[60257] = b[14] & g[27490];
assign g[43875] = a[14] & g[27491];
assign g[60258] = b[14] & g[27491];
assign g[43876] = a[14] & g[27492];
assign g[60259] = b[14] & g[27492];
assign g[43877] = a[14] & g[27493];
assign g[60260] = b[14] & g[27493];
assign g[43878] = a[14] & g[27494];
assign g[60261] = b[14] & g[27494];
assign g[43879] = a[14] & g[27495];
assign g[60262] = b[14] & g[27495];
assign g[43880] = a[14] & g[27496];
assign g[60263] = b[14] & g[27496];
assign g[43881] = a[14] & g[27497];
assign g[60264] = b[14] & g[27497];
assign g[43882] = a[14] & g[27498];
assign g[60265] = b[14] & g[27498];
assign g[43883] = a[14] & g[27499];
assign g[60266] = b[14] & g[27499];
assign g[43884] = a[14] & g[27500];
assign g[60267] = b[14] & g[27500];
assign g[43885] = a[14] & g[27501];
assign g[60268] = b[14] & g[27501];
assign g[43886] = a[14] & g[27502];
assign g[60269] = b[14] & g[27502];
assign g[43887] = a[14] & g[27503];
assign g[60270] = b[14] & g[27503];
assign g[43888] = a[14] & g[27504];
assign g[60271] = b[14] & g[27504];
assign g[43889] = a[14] & g[27505];
assign g[60272] = b[14] & g[27505];
assign g[43890] = a[14] & g[27506];
assign g[60273] = b[14] & g[27506];
assign g[43891] = a[14] & g[27507];
assign g[60274] = b[14] & g[27507];
assign g[43892] = a[14] & g[27508];
assign g[60275] = b[14] & g[27508];
assign g[43893] = a[14] & g[27509];
assign g[60276] = b[14] & g[27509];
assign g[43894] = a[14] & g[27510];
assign g[60277] = b[14] & g[27510];
assign g[43895] = a[14] & g[27511];
assign g[60278] = b[14] & g[27511];
assign g[43896] = a[14] & g[27512];
assign g[60279] = b[14] & g[27512];
assign g[43897] = a[14] & g[27513];
assign g[60280] = b[14] & g[27513];
assign g[43898] = a[14] & g[27514];
assign g[60281] = b[14] & g[27514];
assign g[43899] = a[14] & g[27515];
assign g[60282] = b[14] & g[27515];
assign g[43900] = a[14] & g[27516];
assign g[60283] = b[14] & g[27516];
assign g[43901] = a[14] & g[27517];
assign g[60284] = b[14] & g[27517];
assign g[43902] = a[14] & g[27518];
assign g[60285] = b[14] & g[27518];
assign g[43903] = a[14] & g[27519];
assign g[60286] = b[14] & g[27519];
assign g[43904] = a[14] & g[27520];
assign g[60287] = b[14] & g[27520];
assign g[43905] = a[14] & g[27521];
assign g[60288] = b[14] & g[27521];
assign g[43906] = a[14] & g[27522];
assign g[60289] = b[14] & g[27522];
assign g[43907] = a[14] & g[27523];
assign g[60290] = b[14] & g[27523];
assign g[43908] = a[14] & g[27524];
assign g[60291] = b[14] & g[27524];
assign g[43909] = a[14] & g[27525];
assign g[60292] = b[14] & g[27525];
assign g[43910] = a[14] & g[27526];
assign g[60293] = b[14] & g[27526];
assign g[43911] = a[14] & g[27527];
assign g[60294] = b[14] & g[27527];
assign g[43912] = a[14] & g[27528];
assign g[60295] = b[14] & g[27528];
assign g[43913] = a[14] & g[27529];
assign g[60296] = b[14] & g[27529];
assign g[43914] = a[14] & g[27530];
assign g[60297] = b[14] & g[27530];
assign g[43915] = a[14] & g[27531];
assign g[60298] = b[14] & g[27531];
assign g[43916] = a[14] & g[27532];
assign g[60299] = b[14] & g[27532];
assign g[43917] = a[14] & g[27533];
assign g[60300] = b[14] & g[27533];
assign g[43918] = a[14] & g[27534];
assign g[60301] = b[14] & g[27534];
assign g[43919] = a[14] & g[27535];
assign g[60302] = b[14] & g[27535];
assign g[43920] = a[14] & g[27536];
assign g[60303] = b[14] & g[27536];
assign g[43921] = a[14] & g[27537];
assign g[60304] = b[14] & g[27537];
assign g[43922] = a[14] & g[27538];
assign g[60305] = b[14] & g[27538];
assign g[43923] = a[14] & g[27539];
assign g[60306] = b[14] & g[27539];
assign g[43924] = a[14] & g[27540];
assign g[60307] = b[14] & g[27540];
assign g[43925] = a[14] & g[27541];
assign g[60308] = b[14] & g[27541];
assign g[43926] = a[14] & g[27542];
assign g[60309] = b[14] & g[27542];
assign g[43927] = a[14] & g[27543];
assign g[60310] = b[14] & g[27543];
assign g[43928] = a[14] & g[27544];
assign g[60311] = b[14] & g[27544];
assign g[43929] = a[14] & g[27545];
assign g[60312] = b[14] & g[27545];
assign g[43930] = a[14] & g[27546];
assign g[60313] = b[14] & g[27546];
assign g[43931] = a[14] & g[27547];
assign g[60314] = b[14] & g[27547];
assign g[43932] = a[14] & g[27548];
assign g[60315] = b[14] & g[27548];
assign g[43933] = a[14] & g[27549];
assign g[60316] = b[14] & g[27549];
assign g[43934] = a[14] & g[27550];
assign g[60317] = b[14] & g[27550];
assign g[43935] = a[14] & g[27551];
assign g[60318] = b[14] & g[27551];
assign g[43936] = a[14] & g[27552];
assign g[60319] = b[14] & g[27552];
assign g[43937] = a[14] & g[27553];
assign g[60320] = b[14] & g[27553];
assign g[43938] = a[14] & g[27554];
assign g[60321] = b[14] & g[27554];
assign g[43939] = a[14] & g[27555];
assign g[60322] = b[14] & g[27555];
assign g[43940] = a[14] & g[27556];
assign g[60323] = b[14] & g[27556];
assign g[43941] = a[14] & g[27557];
assign g[60324] = b[14] & g[27557];
assign g[43942] = a[14] & g[27558];
assign g[60325] = b[14] & g[27558];
assign g[43943] = a[14] & g[27559];
assign g[60326] = b[14] & g[27559];
assign g[43944] = a[14] & g[27560];
assign g[60327] = b[14] & g[27560];
assign g[43945] = a[14] & g[27561];
assign g[60328] = b[14] & g[27561];
assign g[43946] = a[14] & g[27562];
assign g[60329] = b[14] & g[27562];
assign g[43947] = a[14] & g[27563];
assign g[60330] = b[14] & g[27563];
assign g[43948] = a[14] & g[27564];
assign g[60331] = b[14] & g[27564];
assign g[43949] = a[14] & g[27565];
assign g[60332] = b[14] & g[27565];
assign g[43950] = a[14] & g[27566];
assign g[60333] = b[14] & g[27566];
assign g[43951] = a[14] & g[27567];
assign g[60334] = b[14] & g[27567];
assign g[43952] = a[14] & g[27568];
assign g[60335] = b[14] & g[27568];
assign g[43953] = a[14] & g[27569];
assign g[60336] = b[14] & g[27569];
assign g[43954] = a[14] & g[27570];
assign g[60337] = b[14] & g[27570];
assign g[43955] = a[14] & g[27571];
assign g[60338] = b[14] & g[27571];
assign g[43956] = a[14] & g[27572];
assign g[60339] = b[14] & g[27572];
assign g[43957] = a[14] & g[27573];
assign g[60340] = b[14] & g[27573];
assign g[43958] = a[14] & g[27574];
assign g[60341] = b[14] & g[27574];
assign g[43959] = a[14] & g[27575];
assign g[60342] = b[14] & g[27575];
assign g[43960] = a[14] & g[27576];
assign g[60343] = b[14] & g[27576];
assign g[43961] = a[14] & g[27577];
assign g[60344] = b[14] & g[27577];
assign g[43962] = a[14] & g[27578];
assign g[60345] = b[14] & g[27578];
assign g[43963] = a[14] & g[27579];
assign g[60346] = b[14] & g[27579];
assign g[43964] = a[14] & g[27580];
assign g[60347] = b[14] & g[27580];
assign g[43965] = a[14] & g[27581];
assign g[60348] = b[14] & g[27581];
assign g[43966] = a[14] & g[27582];
assign g[60349] = b[14] & g[27582];
assign g[43967] = a[14] & g[27583];
assign g[60350] = b[14] & g[27583];
assign g[43968] = a[14] & g[27584];
assign g[60351] = b[14] & g[27584];
assign g[43969] = a[14] & g[27585];
assign g[60352] = b[14] & g[27585];
assign g[43970] = a[14] & g[27586];
assign g[60353] = b[14] & g[27586];
assign g[43971] = a[14] & g[27587];
assign g[60354] = b[14] & g[27587];
assign g[43972] = a[14] & g[27588];
assign g[60355] = b[14] & g[27588];
assign g[43973] = a[14] & g[27589];
assign g[60356] = b[14] & g[27589];
assign g[43974] = a[14] & g[27590];
assign g[60357] = b[14] & g[27590];
assign g[43975] = a[14] & g[27591];
assign g[60358] = b[14] & g[27591];
assign g[43976] = a[14] & g[27592];
assign g[60359] = b[14] & g[27592];
assign g[43977] = a[14] & g[27593];
assign g[60360] = b[14] & g[27593];
assign g[43978] = a[14] & g[27594];
assign g[60361] = b[14] & g[27594];
assign g[43979] = a[14] & g[27595];
assign g[60362] = b[14] & g[27595];
assign g[43980] = a[14] & g[27596];
assign g[60363] = b[14] & g[27596];
assign g[43981] = a[14] & g[27597];
assign g[60364] = b[14] & g[27597];
assign g[43982] = a[14] & g[27598];
assign g[60365] = b[14] & g[27598];
assign g[43983] = a[14] & g[27599];
assign g[60366] = b[14] & g[27599];
assign g[43984] = a[14] & g[27600];
assign g[60367] = b[14] & g[27600];
assign g[43985] = a[14] & g[27601];
assign g[60368] = b[14] & g[27601];
assign g[43986] = a[14] & g[27602];
assign g[60369] = b[14] & g[27602];
assign g[43987] = a[14] & g[27603];
assign g[60370] = b[14] & g[27603];
assign g[43988] = a[14] & g[27604];
assign g[60371] = b[14] & g[27604];
assign g[43989] = a[14] & g[27605];
assign g[60372] = b[14] & g[27605];
assign g[43990] = a[14] & g[27606];
assign g[60373] = b[14] & g[27606];
assign g[43991] = a[14] & g[27607];
assign g[60374] = b[14] & g[27607];
assign g[43992] = a[14] & g[27608];
assign g[60375] = b[14] & g[27608];
assign g[43993] = a[14] & g[27609];
assign g[60376] = b[14] & g[27609];
assign g[43994] = a[14] & g[27610];
assign g[60377] = b[14] & g[27610];
assign g[43995] = a[14] & g[27611];
assign g[60378] = b[14] & g[27611];
assign g[43996] = a[14] & g[27612];
assign g[60379] = b[14] & g[27612];
assign g[43997] = a[14] & g[27613];
assign g[60380] = b[14] & g[27613];
assign g[43998] = a[14] & g[27614];
assign g[60381] = b[14] & g[27614];
assign g[43999] = a[14] & g[27615];
assign g[60382] = b[14] & g[27615];
assign g[44000] = a[14] & g[27616];
assign g[60383] = b[14] & g[27616];
assign g[44001] = a[14] & g[27617];
assign g[60384] = b[14] & g[27617];
assign g[44002] = a[14] & g[27618];
assign g[60385] = b[14] & g[27618];
assign g[44003] = a[14] & g[27619];
assign g[60386] = b[14] & g[27619];
assign g[44004] = a[14] & g[27620];
assign g[60387] = b[14] & g[27620];
assign g[44005] = a[14] & g[27621];
assign g[60388] = b[14] & g[27621];
assign g[44006] = a[14] & g[27622];
assign g[60389] = b[14] & g[27622];
assign g[44007] = a[14] & g[27623];
assign g[60390] = b[14] & g[27623];
assign g[44008] = a[14] & g[27624];
assign g[60391] = b[14] & g[27624];
assign g[44009] = a[14] & g[27625];
assign g[60392] = b[14] & g[27625];
assign g[44010] = a[14] & g[27626];
assign g[60393] = b[14] & g[27626];
assign g[44011] = a[14] & g[27627];
assign g[60394] = b[14] & g[27627];
assign g[44012] = a[14] & g[27628];
assign g[60395] = b[14] & g[27628];
assign g[44013] = a[14] & g[27629];
assign g[60396] = b[14] & g[27629];
assign g[44014] = a[14] & g[27630];
assign g[60397] = b[14] & g[27630];
assign g[44015] = a[14] & g[27631];
assign g[60398] = b[14] & g[27631];
assign g[44016] = a[14] & g[27632];
assign g[60399] = b[14] & g[27632];
assign g[44017] = a[14] & g[27633];
assign g[60400] = b[14] & g[27633];
assign g[44018] = a[14] & g[27634];
assign g[60401] = b[14] & g[27634];
assign g[44019] = a[14] & g[27635];
assign g[60402] = b[14] & g[27635];
assign g[44020] = a[14] & g[27636];
assign g[60403] = b[14] & g[27636];
assign g[44021] = a[14] & g[27637];
assign g[60404] = b[14] & g[27637];
assign g[44022] = a[14] & g[27638];
assign g[60405] = b[14] & g[27638];
assign g[44023] = a[14] & g[27639];
assign g[60406] = b[14] & g[27639];
assign g[44024] = a[14] & g[27640];
assign g[60407] = b[14] & g[27640];
assign g[44025] = a[14] & g[27641];
assign g[60408] = b[14] & g[27641];
assign g[44026] = a[14] & g[27642];
assign g[60409] = b[14] & g[27642];
assign g[44027] = a[14] & g[27643];
assign g[60410] = b[14] & g[27643];
assign g[44028] = a[14] & g[27644];
assign g[60411] = b[14] & g[27644];
assign g[44029] = a[14] & g[27645];
assign g[60412] = b[14] & g[27645];
assign g[44030] = a[14] & g[27646];
assign g[60413] = b[14] & g[27646];
assign g[44031] = a[14] & g[27647];
assign g[60414] = b[14] & g[27647];
assign g[44032] = a[14] & g[27648];
assign g[60415] = b[14] & g[27648];
assign g[44033] = a[14] & g[27649];
assign g[60416] = b[14] & g[27649];
assign g[44034] = a[14] & g[27650];
assign g[60417] = b[14] & g[27650];
assign g[44035] = a[14] & g[27651];
assign g[60418] = b[14] & g[27651];
assign g[44036] = a[14] & g[27652];
assign g[60419] = b[14] & g[27652];
assign g[44037] = a[14] & g[27653];
assign g[60420] = b[14] & g[27653];
assign g[44038] = a[14] & g[27654];
assign g[60421] = b[14] & g[27654];
assign g[44039] = a[14] & g[27655];
assign g[60422] = b[14] & g[27655];
assign g[44040] = a[14] & g[27656];
assign g[60423] = b[14] & g[27656];
assign g[44041] = a[14] & g[27657];
assign g[60424] = b[14] & g[27657];
assign g[44042] = a[14] & g[27658];
assign g[60425] = b[14] & g[27658];
assign g[44043] = a[14] & g[27659];
assign g[60426] = b[14] & g[27659];
assign g[44044] = a[14] & g[27660];
assign g[60427] = b[14] & g[27660];
assign g[44045] = a[14] & g[27661];
assign g[60428] = b[14] & g[27661];
assign g[44046] = a[14] & g[27662];
assign g[60429] = b[14] & g[27662];
assign g[44047] = a[14] & g[27663];
assign g[60430] = b[14] & g[27663];
assign g[44048] = a[14] & g[27664];
assign g[60431] = b[14] & g[27664];
assign g[44049] = a[14] & g[27665];
assign g[60432] = b[14] & g[27665];
assign g[44050] = a[14] & g[27666];
assign g[60433] = b[14] & g[27666];
assign g[44051] = a[14] & g[27667];
assign g[60434] = b[14] & g[27667];
assign g[44052] = a[14] & g[27668];
assign g[60435] = b[14] & g[27668];
assign g[44053] = a[14] & g[27669];
assign g[60436] = b[14] & g[27669];
assign g[44054] = a[14] & g[27670];
assign g[60437] = b[14] & g[27670];
assign g[44055] = a[14] & g[27671];
assign g[60438] = b[14] & g[27671];
assign g[44056] = a[14] & g[27672];
assign g[60439] = b[14] & g[27672];
assign g[44057] = a[14] & g[27673];
assign g[60440] = b[14] & g[27673];
assign g[44058] = a[14] & g[27674];
assign g[60441] = b[14] & g[27674];
assign g[44059] = a[14] & g[27675];
assign g[60442] = b[14] & g[27675];
assign g[44060] = a[14] & g[27676];
assign g[60443] = b[14] & g[27676];
assign g[44061] = a[14] & g[27677];
assign g[60444] = b[14] & g[27677];
assign g[44062] = a[14] & g[27678];
assign g[60445] = b[14] & g[27678];
assign g[44063] = a[14] & g[27679];
assign g[60446] = b[14] & g[27679];
assign g[44064] = a[14] & g[27680];
assign g[60447] = b[14] & g[27680];
assign g[44065] = a[14] & g[27681];
assign g[60448] = b[14] & g[27681];
assign g[44066] = a[14] & g[27682];
assign g[60449] = b[14] & g[27682];
assign g[44067] = a[14] & g[27683];
assign g[60450] = b[14] & g[27683];
assign g[44068] = a[14] & g[27684];
assign g[60451] = b[14] & g[27684];
assign g[44069] = a[14] & g[27685];
assign g[60452] = b[14] & g[27685];
assign g[44070] = a[14] & g[27686];
assign g[60453] = b[14] & g[27686];
assign g[44071] = a[14] & g[27687];
assign g[60454] = b[14] & g[27687];
assign g[44072] = a[14] & g[27688];
assign g[60455] = b[14] & g[27688];
assign g[44073] = a[14] & g[27689];
assign g[60456] = b[14] & g[27689];
assign g[44074] = a[14] & g[27690];
assign g[60457] = b[14] & g[27690];
assign g[44075] = a[14] & g[27691];
assign g[60458] = b[14] & g[27691];
assign g[44076] = a[14] & g[27692];
assign g[60459] = b[14] & g[27692];
assign g[44077] = a[14] & g[27693];
assign g[60460] = b[14] & g[27693];
assign g[44078] = a[14] & g[27694];
assign g[60461] = b[14] & g[27694];
assign g[44079] = a[14] & g[27695];
assign g[60462] = b[14] & g[27695];
assign g[44080] = a[14] & g[27696];
assign g[60463] = b[14] & g[27696];
assign g[44081] = a[14] & g[27697];
assign g[60464] = b[14] & g[27697];
assign g[44082] = a[14] & g[27698];
assign g[60465] = b[14] & g[27698];
assign g[44083] = a[14] & g[27699];
assign g[60466] = b[14] & g[27699];
assign g[44084] = a[14] & g[27700];
assign g[60467] = b[14] & g[27700];
assign g[44085] = a[14] & g[27701];
assign g[60468] = b[14] & g[27701];
assign g[44086] = a[14] & g[27702];
assign g[60469] = b[14] & g[27702];
assign g[44087] = a[14] & g[27703];
assign g[60470] = b[14] & g[27703];
assign g[44088] = a[14] & g[27704];
assign g[60471] = b[14] & g[27704];
assign g[44089] = a[14] & g[27705];
assign g[60472] = b[14] & g[27705];
assign g[44090] = a[14] & g[27706];
assign g[60473] = b[14] & g[27706];
assign g[44091] = a[14] & g[27707];
assign g[60474] = b[14] & g[27707];
assign g[44092] = a[14] & g[27708];
assign g[60475] = b[14] & g[27708];
assign g[44093] = a[14] & g[27709];
assign g[60476] = b[14] & g[27709];
assign g[44094] = a[14] & g[27710];
assign g[60477] = b[14] & g[27710];
assign g[44095] = a[14] & g[27711];
assign g[60478] = b[14] & g[27711];
assign g[44096] = a[14] & g[27712];
assign g[60479] = b[14] & g[27712];
assign g[44097] = a[14] & g[27713];
assign g[60480] = b[14] & g[27713];
assign g[44098] = a[14] & g[27714];
assign g[60481] = b[14] & g[27714];
assign g[44099] = a[14] & g[27715];
assign g[60482] = b[14] & g[27715];
assign g[44100] = a[14] & g[27716];
assign g[60483] = b[14] & g[27716];
assign g[44101] = a[14] & g[27717];
assign g[60484] = b[14] & g[27717];
assign g[44102] = a[14] & g[27718];
assign g[60485] = b[14] & g[27718];
assign g[44103] = a[14] & g[27719];
assign g[60486] = b[14] & g[27719];
assign g[44104] = a[14] & g[27720];
assign g[60487] = b[14] & g[27720];
assign g[44105] = a[14] & g[27721];
assign g[60488] = b[14] & g[27721];
assign g[44106] = a[14] & g[27722];
assign g[60489] = b[14] & g[27722];
assign g[44107] = a[14] & g[27723];
assign g[60490] = b[14] & g[27723];
assign g[44108] = a[14] & g[27724];
assign g[60491] = b[14] & g[27724];
assign g[44109] = a[14] & g[27725];
assign g[60492] = b[14] & g[27725];
assign g[44110] = a[14] & g[27726];
assign g[60493] = b[14] & g[27726];
assign g[44111] = a[14] & g[27727];
assign g[60494] = b[14] & g[27727];
assign g[44112] = a[14] & g[27728];
assign g[60495] = b[14] & g[27728];
assign g[44113] = a[14] & g[27729];
assign g[60496] = b[14] & g[27729];
assign g[44114] = a[14] & g[27730];
assign g[60497] = b[14] & g[27730];
assign g[44115] = a[14] & g[27731];
assign g[60498] = b[14] & g[27731];
assign g[44116] = a[14] & g[27732];
assign g[60499] = b[14] & g[27732];
assign g[44117] = a[14] & g[27733];
assign g[60500] = b[14] & g[27733];
assign g[44118] = a[14] & g[27734];
assign g[60501] = b[14] & g[27734];
assign g[44119] = a[14] & g[27735];
assign g[60502] = b[14] & g[27735];
assign g[44120] = a[14] & g[27736];
assign g[60503] = b[14] & g[27736];
assign g[44121] = a[14] & g[27737];
assign g[60504] = b[14] & g[27737];
assign g[44122] = a[14] & g[27738];
assign g[60505] = b[14] & g[27738];
assign g[44123] = a[14] & g[27739];
assign g[60506] = b[14] & g[27739];
assign g[44124] = a[14] & g[27740];
assign g[60507] = b[14] & g[27740];
assign g[44125] = a[14] & g[27741];
assign g[60508] = b[14] & g[27741];
assign g[44126] = a[14] & g[27742];
assign g[60509] = b[14] & g[27742];
assign g[44127] = a[14] & g[27743];
assign g[60510] = b[14] & g[27743];
assign g[44128] = a[14] & g[27744];
assign g[60511] = b[14] & g[27744];
assign g[44129] = a[14] & g[27745];
assign g[60512] = b[14] & g[27745];
assign g[44130] = a[14] & g[27746];
assign g[60513] = b[14] & g[27746];
assign g[44131] = a[14] & g[27747];
assign g[60514] = b[14] & g[27747];
assign g[44132] = a[14] & g[27748];
assign g[60515] = b[14] & g[27748];
assign g[44133] = a[14] & g[27749];
assign g[60516] = b[14] & g[27749];
assign g[44134] = a[14] & g[27750];
assign g[60517] = b[14] & g[27750];
assign g[44135] = a[14] & g[27751];
assign g[60518] = b[14] & g[27751];
assign g[44136] = a[14] & g[27752];
assign g[60519] = b[14] & g[27752];
assign g[44137] = a[14] & g[27753];
assign g[60520] = b[14] & g[27753];
assign g[44138] = a[14] & g[27754];
assign g[60521] = b[14] & g[27754];
assign g[44139] = a[14] & g[27755];
assign g[60522] = b[14] & g[27755];
assign g[44140] = a[14] & g[27756];
assign g[60523] = b[14] & g[27756];
assign g[44141] = a[14] & g[27757];
assign g[60524] = b[14] & g[27757];
assign g[44142] = a[14] & g[27758];
assign g[60525] = b[14] & g[27758];
assign g[44143] = a[14] & g[27759];
assign g[60526] = b[14] & g[27759];
assign g[44144] = a[14] & g[27760];
assign g[60527] = b[14] & g[27760];
assign g[44145] = a[14] & g[27761];
assign g[60528] = b[14] & g[27761];
assign g[44146] = a[14] & g[27762];
assign g[60529] = b[14] & g[27762];
assign g[44147] = a[14] & g[27763];
assign g[60530] = b[14] & g[27763];
assign g[44148] = a[14] & g[27764];
assign g[60531] = b[14] & g[27764];
assign g[44149] = a[14] & g[27765];
assign g[60532] = b[14] & g[27765];
assign g[44150] = a[14] & g[27766];
assign g[60533] = b[14] & g[27766];
assign g[44151] = a[14] & g[27767];
assign g[60534] = b[14] & g[27767];
assign g[44152] = a[14] & g[27768];
assign g[60535] = b[14] & g[27768];
assign g[44153] = a[14] & g[27769];
assign g[60536] = b[14] & g[27769];
assign g[44154] = a[14] & g[27770];
assign g[60537] = b[14] & g[27770];
assign g[44155] = a[14] & g[27771];
assign g[60538] = b[14] & g[27771];
assign g[44156] = a[14] & g[27772];
assign g[60539] = b[14] & g[27772];
assign g[44157] = a[14] & g[27773];
assign g[60540] = b[14] & g[27773];
assign g[44158] = a[14] & g[27774];
assign g[60541] = b[14] & g[27774];
assign g[44159] = a[14] & g[27775];
assign g[60542] = b[14] & g[27775];
assign g[44160] = a[14] & g[27776];
assign g[60543] = b[14] & g[27776];
assign g[44161] = a[14] & g[27777];
assign g[60544] = b[14] & g[27777];
assign g[44162] = a[14] & g[27778];
assign g[60545] = b[14] & g[27778];
assign g[44163] = a[14] & g[27779];
assign g[60546] = b[14] & g[27779];
assign g[44164] = a[14] & g[27780];
assign g[60547] = b[14] & g[27780];
assign g[44165] = a[14] & g[27781];
assign g[60548] = b[14] & g[27781];
assign g[44166] = a[14] & g[27782];
assign g[60549] = b[14] & g[27782];
assign g[44167] = a[14] & g[27783];
assign g[60550] = b[14] & g[27783];
assign g[44168] = a[14] & g[27784];
assign g[60551] = b[14] & g[27784];
assign g[44169] = a[14] & g[27785];
assign g[60552] = b[14] & g[27785];
assign g[44170] = a[14] & g[27786];
assign g[60553] = b[14] & g[27786];
assign g[44171] = a[14] & g[27787];
assign g[60554] = b[14] & g[27787];
assign g[44172] = a[14] & g[27788];
assign g[60555] = b[14] & g[27788];
assign g[44173] = a[14] & g[27789];
assign g[60556] = b[14] & g[27789];
assign g[44174] = a[14] & g[27790];
assign g[60557] = b[14] & g[27790];
assign g[44175] = a[14] & g[27791];
assign g[60558] = b[14] & g[27791];
assign g[44176] = a[14] & g[27792];
assign g[60559] = b[14] & g[27792];
assign g[44177] = a[14] & g[27793];
assign g[60560] = b[14] & g[27793];
assign g[44178] = a[14] & g[27794];
assign g[60561] = b[14] & g[27794];
assign g[44179] = a[14] & g[27795];
assign g[60562] = b[14] & g[27795];
assign g[44180] = a[14] & g[27796];
assign g[60563] = b[14] & g[27796];
assign g[44181] = a[14] & g[27797];
assign g[60564] = b[14] & g[27797];
assign g[44182] = a[14] & g[27798];
assign g[60565] = b[14] & g[27798];
assign g[44183] = a[14] & g[27799];
assign g[60566] = b[14] & g[27799];
assign g[44184] = a[14] & g[27800];
assign g[60567] = b[14] & g[27800];
assign g[44185] = a[14] & g[27801];
assign g[60568] = b[14] & g[27801];
assign g[44186] = a[14] & g[27802];
assign g[60569] = b[14] & g[27802];
assign g[44187] = a[14] & g[27803];
assign g[60570] = b[14] & g[27803];
assign g[44188] = a[14] & g[27804];
assign g[60571] = b[14] & g[27804];
assign g[44189] = a[14] & g[27805];
assign g[60572] = b[14] & g[27805];
assign g[44190] = a[14] & g[27806];
assign g[60573] = b[14] & g[27806];
assign g[44191] = a[14] & g[27807];
assign g[60574] = b[14] & g[27807];
assign g[44192] = a[14] & g[27808];
assign g[60575] = b[14] & g[27808];
assign g[44193] = a[14] & g[27809];
assign g[60576] = b[14] & g[27809];
assign g[44194] = a[14] & g[27810];
assign g[60577] = b[14] & g[27810];
assign g[44195] = a[14] & g[27811];
assign g[60578] = b[14] & g[27811];
assign g[44196] = a[14] & g[27812];
assign g[60579] = b[14] & g[27812];
assign g[44197] = a[14] & g[27813];
assign g[60580] = b[14] & g[27813];
assign g[44198] = a[14] & g[27814];
assign g[60581] = b[14] & g[27814];
assign g[44199] = a[14] & g[27815];
assign g[60582] = b[14] & g[27815];
assign g[44200] = a[14] & g[27816];
assign g[60583] = b[14] & g[27816];
assign g[44201] = a[14] & g[27817];
assign g[60584] = b[14] & g[27817];
assign g[44202] = a[14] & g[27818];
assign g[60585] = b[14] & g[27818];
assign g[44203] = a[14] & g[27819];
assign g[60586] = b[14] & g[27819];
assign g[44204] = a[14] & g[27820];
assign g[60587] = b[14] & g[27820];
assign g[44205] = a[14] & g[27821];
assign g[60588] = b[14] & g[27821];
assign g[44206] = a[14] & g[27822];
assign g[60589] = b[14] & g[27822];
assign g[44207] = a[14] & g[27823];
assign g[60590] = b[14] & g[27823];
assign g[44208] = a[14] & g[27824];
assign g[60591] = b[14] & g[27824];
assign g[44209] = a[14] & g[27825];
assign g[60592] = b[14] & g[27825];
assign g[44210] = a[14] & g[27826];
assign g[60593] = b[14] & g[27826];
assign g[44211] = a[14] & g[27827];
assign g[60594] = b[14] & g[27827];
assign g[44212] = a[14] & g[27828];
assign g[60595] = b[14] & g[27828];
assign g[44213] = a[14] & g[27829];
assign g[60596] = b[14] & g[27829];
assign g[44214] = a[14] & g[27830];
assign g[60597] = b[14] & g[27830];
assign g[44215] = a[14] & g[27831];
assign g[60598] = b[14] & g[27831];
assign g[44216] = a[14] & g[27832];
assign g[60599] = b[14] & g[27832];
assign g[44217] = a[14] & g[27833];
assign g[60600] = b[14] & g[27833];
assign g[44218] = a[14] & g[27834];
assign g[60601] = b[14] & g[27834];
assign g[44219] = a[14] & g[27835];
assign g[60602] = b[14] & g[27835];
assign g[44220] = a[14] & g[27836];
assign g[60603] = b[14] & g[27836];
assign g[44221] = a[14] & g[27837];
assign g[60604] = b[14] & g[27837];
assign g[44222] = a[14] & g[27838];
assign g[60605] = b[14] & g[27838];
assign g[44223] = a[14] & g[27839];
assign g[60606] = b[14] & g[27839];
assign g[44224] = a[14] & g[27840];
assign g[60607] = b[14] & g[27840];
assign g[44225] = a[14] & g[27841];
assign g[60608] = b[14] & g[27841];
assign g[44226] = a[14] & g[27842];
assign g[60609] = b[14] & g[27842];
assign g[44227] = a[14] & g[27843];
assign g[60610] = b[14] & g[27843];
assign g[44228] = a[14] & g[27844];
assign g[60611] = b[14] & g[27844];
assign g[44229] = a[14] & g[27845];
assign g[60612] = b[14] & g[27845];
assign g[44230] = a[14] & g[27846];
assign g[60613] = b[14] & g[27846];
assign g[44231] = a[14] & g[27847];
assign g[60614] = b[14] & g[27847];
assign g[44232] = a[14] & g[27848];
assign g[60615] = b[14] & g[27848];
assign g[44233] = a[14] & g[27849];
assign g[60616] = b[14] & g[27849];
assign g[44234] = a[14] & g[27850];
assign g[60617] = b[14] & g[27850];
assign g[44235] = a[14] & g[27851];
assign g[60618] = b[14] & g[27851];
assign g[44236] = a[14] & g[27852];
assign g[60619] = b[14] & g[27852];
assign g[44237] = a[14] & g[27853];
assign g[60620] = b[14] & g[27853];
assign g[44238] = a[14] & g[27854];
assign g[60621] = b[14] & g[27854];
assign g[44239] = a[14] & g[27855];
assign g[60622] = b[14] & g[27855];
assign g[44240] = a[14] & g[27856];
assign g[60623] = b[14] & g[27856];
assign g[44241] = a[14] & g[27857];
assign g[60624] = b[14] & g[27857];
assign g[44242] = a[14] & g[27858];
assign g[60625] = b[14] & g[27858];
assign g[44243] = a[14] & g[27859];
assign g[60626] = b[14] & g[27859];
assign g[44244] = a[14] & g[27860];
assign g[60627] = b[14] & g[27860];
assign g[44245] = a[14] & g[27861];
assign g[60628] = b[14] & g[27861];
assign g[44246] = a[14] & g[27862];
assign g[60629] = b[14] & g[27862];
assign g[44247] = a[14] & g[27863];
assign g[60630] = b[14] & g[27863];
assign g[44248] = a[14] & g[27864];
assign g[60631] = b[14] & g[27864];
assign g[44249] = a[14] & g[27865];
assign g[60632] = b[14] & g[27865];
assign g[44250] = a[14] & g[27866];
assign g[60633] = b[14] & g[27866];
assign g[44251] = a[14] & g[27867];
assign g[60634] = b[14] & g[27867];
assign g[44252] = a[14] & g[27868];
assign g[60635] = b[14] & g[27868];
assign g[44253] = a[14] & g[27869];
assign g[60636] = b[14] & g[27869];
assign g[44254] = a[14] & g[27870];
assign g[60637] = b[14] & g[27870];
assign g[44255] = a[14] & g[27871];
assign g[60638] = b[14] & g[27871];
assign g[44256] = a[14] & g[27872];
assign g[60639] = b[14] & g[27872];
assign g[44257] = a[14] & g[27873];
assign g[60640] = b[14] & g[27873];
assign g[44258] = a[14] & g[27874];
assign g[60641] = b[14] & g[27874];
assign g[44259] = a[14] & g[27875];
assign g[60642] = b[14] & g[27875];
assign g[44260] = a[14] & g[27876];
assign g[60643] = b[14] & g[27876];
assign g[44261] = a[14] & g[27877];
assign g[60644] = b[14] & g[27877];
assign g[44262] = a[14] & g[27878];
assign g[60645] = b[14] & g[27878];
assign g[44263] = a[14] & g[27879];
assign g[60646] = b[14] & g[27879];
assign g[44264] = a[14] & g[27880];
assign g[60647] = b[14] & g[27880];
assign g[44265] = a[14] & g[27881];
assign g[60648] = b[14] & g[27881];
assign g[44266] = a[14] & g[27882];
assign g[60649] = b[14] & g[27882];
assign g[44267] = a[14] & g[27883];
assign g[60650] = b[14] & g[27883];
assign g[44268] = a[14] & g[27884];
assign g[60651] = b[14] & g[27884];
assign g[44269] = a[14] & g[27885];
assign g[60652] = b[14] & g[27885];
assign g[44270] = a[14] & g[27886];
assign g[60653] = b[14] & g[27886];
assign g[44271] = a[14] & g[27887];
assign g[60654] = b[14] & g[27887];
assign g[44272] = a[14] & g[27888];
assign g[60655] = b[14] & g[27888];
assign g[44273] = a[14] & g[27889];
assign g[60656] = b[14] & g[27889];
assign g[44274] = a[14] & g[27890];
assign g[60657] = b[14] & g[27890];
assign g[44275] = a[14] & g[27891];
assign g[60658] = b[14] & g[27891];
assign g[44276] = a[14] & g[27892];
assign g[60659] = b[14] & g[27892];
assign g[44277] = a[14] & g[27893];
assign g[60660] = b[14] & g[27893];
assign g[44278] = a[14] & g[27894];
assign g[60661] = b[14] & g[27894];
assign g[44279] = a[14] & g[27895];
assign g[60662] = b[14] & g[27895];
assign g[44280] = a[14] & g[27896];
assign g[60663] = b[14] & g[27896];
assign g[44281] = a[14] & g[27897];
assign g[60664] = b[14] & g[27897];
assign g[44282] = a[14] & g[27898];
assign g[60665] = b[14] & g[27898];
assign g[44283] = a[14] & g[27899];
assign g[60666] = b[14] & g[27899];
assign g[44284] = a[14] & g[27900];
assign g[60667] = b[14] & g[27900];
assign g[44285] = a[14] & g[27901];
assign g[60668] = b[14] & g[27901];
assign g[44286] = a[14] & g[27902];
assign g[60669] = b[14] & g[27902];
assign g[44287] = a[14] & g[27903];
assign g[60670] = b[14] & g[27903];
assign g[44288] = a[14] & g[27904];
assign g[60671] = b[14] & g[27904];
assign g[44289] = a[14] & g[27905];
assign g[60672] = b[14] & g[27905];
assign g[44290] = a[14] & g[27906];
assign g[60673] = b[14] & g[27906];
assign g[44291] = a[14] & g[27907];
assign g[60674] = b[14] & g[27907];
assign g[44292] = a[14] & g[27908];
assign g[60675] = b[14] & g[27908];
assign g[44293] = a[14] & g[27909];
assign g[60676] = b[14] & g[27909];
assign g[44294] = a[14] & g[27910];
assign g[60677] = b[14] & g[27910];
assign g[44295] = a[14] & g[27911];
assign g[60678] = b[14] & g[27911];
assign g[44296] = a[14] & g[27912];
assign g[60679] = b[14] & g[27912];
assign g[44297] = a[14] & g[27913];
assign g[60680] = b[14] & g[27913];
assign g[44298] = a[14] & g[27914];
assign g[60681] = b[14] & g[27914];
assign g[44299] = a[14] & g[27915];
assign g[60682] = b[14] & g[27915];
assign g[44300] = a[14] & g[27916];
assign g[60683] = b[14] & g[27916];
assign g[44301] = a[14] & g[27917];
assign g[60684] = b[14] & g[27917];
assign g[44302] = a[14] & g[27918];
assign g[60685] = b[14] & g[27918];
assign g[44303] = a[14] & g[27919];
assign g[60686] = b[14] & g[27919];
assign g[44304] = a[14] & g[27920];
assign g[60687] = b[14] & g[27920];
assign g[44305] = a[14] & g[27921];
assign g[60688] = b[14] & g[27921];
assign g[44306] = a[14] & g[27922];
assign g[60689] = b[14] & g[27922];
assign g[44307] = a[14] & g[27923];
assign g[60690] = b[14] & g[27923];
assign g[44308] = a[14] & g[27924];
assign g[60691] = b[14] & g[27924];
assign g[44309] = a[14] & g[27925];
assign g[60692] = b[14] & g[27925];
assign g[44310] = a[14] & g[27926];
assign g[60693] = b[14] & g[27926];
assign g[44311] = a[14] & g[27927];
assign g[60694] = b[14] & g[27927];
assign g[44312] = a[14] & g[27928];
assign g[60695] = b[14] & g[27928];
assign g[44313] = a[14] & g[27929];
assign g[60696] = b[14] & g[27929];
assign g[44314] = a[14] & g[27930];
assign g[60697] = b[14] & g[27930];
assign g[44315] = a[14] & g[27931];
assign g[60698] = b[14] & g[27931];
assign g[44316] = a[14] & g[27932];
assign g[60699] = b[14] & g[27932];
assign g[44317] = a[14] & g[27933];
assign g[60700] = b[14] & g[27933];
assign g[44318] = a[14] & g[27934];
assign g[60701] = b[14] & g[27934];
assign g[44319] = a[14] & g[27935];
assign g[60702] = b[14] & g[27935];
assign g[44320] = a[14] & g[27936];
assign g[60703] = b[14] & g[27936];
assign g[44321] = a[14] & g[27937];
assign g[60704] = b[14] & g[27937];
assign g[44322] = a[14] & g[27938];
assign g[60705] = b[14] & g[27938];
assign g[44323] = a[14] & g[27939];
assign g[60706] = b[14] & g[27939];
assign g[44324] = a[14] & g[27940];
assign g[60707] = b[14] & g[27940];
assign g[44325] = a[14] & g[27941];
assign g[60708] = b[14] & g[27941];
assign g[44326] = a[14] & g[27942];
assign g[60709] = b[14] & g[27942];
assign g[44327] = a[14] & g[27943];
assign g[60710] = b[14] & g[27943];
assign g[44328] = a[14] & g[27944];
assign g[60711] = b[14] & g[27944];
assign g[44329] = a[14] & g[27945];
assign g[60712] = b[14] & g[27945];
assign g[44330] = a[14] & g[27946];
assign g[60713] = b[14] & g[27946];
assign g[44331] = a[14] & g[27947];
assign g[60714] = b[14] & g[27947];
assign g[44332] = a[14] & g[27948];
assign g[60715] = b[14] & g[27948];
assign g[44333] = a[14] & g[27949];
assign g[60716] = b[14] & g[27949];
assign g[44334] = a[14] & g[27950];
assign g[60717] = b[14] & g[27950];
assign g[44335] = a[14] & g[27951];
assign g[60718] = b[14] & g[27951];
assign g[44336] = a[14] & g[27952];
assign g[60719] = b[14] & g[27952];
assign g[44337] = a[14] & g[27953];
assign g[60720] = b[14] & g[27953];
assign g[44338] = a[14] & g[27954];
assign g[60721] = b[14] & g[27954];
assign g[44339] = a[14] & g[27955];
assign g[60722] = b[14] & g[27955];
assign g[44340] = a[14] & g[27956];
assign g[60723] = b[14] & g[27956];
assign g[44341] = a[14] & g[27957];
assign g[60724] = b[14] & g[27957];
assign g[44342] = a[14] & g[27958];
assign g[60725] = b[14] & g[27958];
assign g[44343] = a[14] & g[27959];
assign g[60726] = b[14] & g[27959];
assign g[44344] = a[14] & g[27960];
assign g[60727] = b[14] & g[27960];
assign g[44345] = a[14] & g[27961];
assign g[60728] = b[14] & g[27961];
assign g[44346] = a[14] & g[27962];
assign g[60729] = b[14] & g[27962];
assign g[44347] = a[14] & g[27963];
assign g[60730] = b[14] & g[27963];
assign g[44348] = a[14] & g[27964];
assign g[60731] = b[14] & g[27964];
assign g[44349] = a[14] & g[27965];
assign g[60732] = b[14] & g[27965];
assign g[44350] = a[14] & g[27966];
assign g[60733] = b[14] & g[27966];
assign g[44351] = a[14] & g[27967];
assign g[60734] = b[14] & g[27967];
assign g[44352] = a[14] & g[27968];
assign g[60735] = b[14] & g[27968];
assign g[44353] = a[14] & g[27969];
assign g[60736] = b[14] & g[27969];
assign g[44354] = a[14] & g[27970];
assign g[60737] = b[14] & g[27970];
assign g[44355] = a[14] & g[27971];
assign g[60738] = b[14] & g[27971];
assign g[44356] = a[14] & g[27972];
assign g[60739] = b[14] & g[27972];
assign g[44357] = a[14] & g[27973];
assign g[60740] = b[14] & g[27973];
assign g[44358] = a[14] & g[27974];
assign g[60741] = b[14] & g[27974];
assign g[44359] = a[14] & g[27975];
assign g[60742] = b[14] & g[27975];
assign g[44360] = a[14] & g[27976];
assign g[60743] = b[14] & g[27976];
assign g[44361] = a[14] & g[27977];
assign g[60744] = b[14] & g[27977];
assign g[44362] = a[14] & g[27978];
assign g[60745] = b[14] & g[27978];
assign g[44363] = a[14] & g[27979];
assign g[60746] = b[14] & g[27979];
assign g[44364] = a[14] & g[27980];
assign g[60747] = b[14] & g[27980];
assign g[44365] = a[14] & g[27981];
assign g[60748] = b[14] & g[27981];
assign g[44366] = a[14] & g[27982];
assign g[60749] = b[14] & g[27982];
assign g[44367] = a[14] & g[27983];
assign g[60750] = b[14] & g[27983];
assign g[44368] = a[14] & g[27984];
assign g[60751] = b[14] & g[27984];
assign g[44369] = a[14] & g[27985];
assign g[60752] = b[14] & g[27985];
assign g[44370] = a[14] & g[27986];
assign g[60753] = b[14] & g[27986];
assign g[44371] = a[14] & g[27987];
assign g[60754] = b[14] & g[27987];
assign g[44372] = a[14] & g[27988];
assign g[60755] = b[14] & g[27988];
assign g[44373] = a[14] & g[27989];
assign g[60756] = b[14] & g[27989];
assign g[44374] = a[14] & g[27990];
assign g[60757] = b[14] & g[27990];
assign g[44375] = a[14] & g[27991];
assign g[60758] = b[14] & g[27991];
assign g[44376] = a[14] & g[27992];
assign g[60759] = b[14] & g[27992];
assign g[44377] = a[14] & g[27993];
assign g[60760] = b[14] & g[27993];
assign g[44378] = a[14] & g[27994];
assign g[60761] = b[14] & g[27994];
assign g[44379] = a[14] & g[27995];
assign g[60762] = b[14] & g[27995];
assign g[44380] = a[14] & g[27996];
assign g[60763] = b[14] & g[27996];
assign g[44381] = a[14] & g[27997];
assign g[60764] = b[14] & g[27997];
assign g[44382] = a[14] & g[27998];
assign g[60765] = b[14] & g[27998];
assign g[44383] = a[14] & g[27999];
assign g[60766] = b[14] & g[27999];
assign g[44384] = a[14] & g[28000];
assign g[60767] = b[14] & g[28000];
assign g[44385] = a[14] & g[28001];
assign g[60768] = b[14] & g[28001];
assign g[44386] = a[14] & g[28002];
assign g[60769] = b[14] & g[28002];
assign g[44387] = a[14] & g[28003];
assign g[60770] = b[14] & g[28003];
assign g[44388] = a[14] & g[28004];
assign g[60771] = b[14] & g[28004];
assign g[44389] = a[14] & g[28005];
assign g[60772] = b[14] & g[28005];
assign g[44390] = a[14] & g[28006];
assign g[60773] = b[14] & g[28006];
assign g[44391] = a[14] & g[28007];
assign g[60774] = b[14] & g[28007];
assign g[44392] = a[14] & g[28008];
assign g[60775] = b[14] & g[28008];
assign g[44393] = a[14] & g[28009];
assign g[60776] = b[14] & g[28009];
assign g[44394] = a[14] & g[28010];
assign g[60777] = b[14] & g[28010];
assign g[44395] = a[14] & g[28011];
assign g[60778] = b[14] & g[28011];
assign g[44396] = a[14] & g[28012];
assign g[60779] = b[14] & g[28012];
assign g[44397] = a[14] & g[28013];
assign g[60780] = b[14] & g[28013];
assign g[44398] = a[14] & g[28014];
assign g[60781] = b[14] & g[28014];
assign g[44399] = a[14] & g[28015];
assign g[60782] = b[14] & g[28015];
assign g[44400] = a[14] & g[28016];
assign g[60783] = b[14] & g[28016];
assign g[44401] = a[14] & g[28017];
assign g[60784] = b[14] & g[28017];
assign g[44402] = a[14] & g[28018];
assign g[60785] = b[14] & g[28018];
assign g[44403] = a[14] & g[28019];
assign g[60786] = b[14] & g[28019];
assign g[44404] = a[14] & g[28020];
assign g[60787] = b[14] & g[28020];
assign g[44405] = a[14] & g[28021];
assign g[60788] = b[14] & g[28021];
assign g[44406] = a[14] & g[28022];
assign g[60789] = b[14] & g[28022];
assign g[44407] = a[14] & g[28023];
assign g[60790] = b[14] & g[28023];
assign g[44408] = a[14] & g[28024];
assign g[60791] = b[14] & g[28024];
assign g[44409] = a[14] & g[28025];
assign g[60792] = b[14] & g[28025];
assign g[44410] = a[14] & g[28026];
assign g[60793] = b[14] & g[28026];
assign g[44411] = a[14] & g[28027];
assign g[60794] = b[14] & g[28027];
assign g[44412] = a[14] & g[28028];
assign g[60795] = b[14] & g[28028];
assign g[44413] = a[14] & g[28029];
assign g[60796] = b[14] & g[28029];
assign g[44414] = a[14] & g[28030];
assign g[60797] = b[14] & g[28030];
assign g[44415] = a[14] & g[28031];
assign g[60798] = b[14] & g[28031];
assign g[44416] = a[14] & g[28032];
assign g[60799] = b[14] & g[28032];
assign g[44417] = a[14] & g[28033];
assign g[60800] = b[14] & g[28033];
assign g[44418] = a[14] & g[28034];
assign g[60801] = b[14] & g[28034];
assign g[44419] = a[14] & g[28035];
assign g[60802] = b[14] & g[28035];
assign g[44420] = a[14] & g[28036];
assign g[60803] = b[14] & g[28036];
assign g[44421] = a[14] & g[28037];
assign g[60804] = b[14] & g[28037];
assign g[44422] = a[14] & g[28038];
assign g[60805] = b[14] & g[28038];
assign g[44423] = a[14] & g[28039];
assign g[60806] = b[14] & g[28039];
assign g[44424] = a[14] & g[28040];
assign g[60807] = b[14] & g[28040];
assign g[44425] = a[14] & g[28041];
assign g[60808] = b[14] & g[28041];
assign g[44426] = a[14] & g[28042];
assign g[60809] = b[14] & g[28042];
assign g[44427] = a[14] & g[28043];
assign g[60810] = b[14] & g[28043];
assign g[44428] = a[14] & g[28044];
assign g[60811] = b[14] & g[28044];
assign g[44429] = a[14] & g[28045];
assign g[60812] = b[14] & g[28045];
assign g[44430] = a[14] & g[28046];
assign g[60813] = b[14] & g[28046];
assign g[44431] = a[14] & g[28047];
assign g[60814] = b[14] & g[28047];
assign g[44432] = a[14] & g[28048];
assign g[60815] = b[14] & g[28048];
assign g[44433] = a[14] & g[28049];
assign g[60816] = b[14] & g[28049];
assign g[44434] = a[14] & g[28050];
assign g[60817] = b[14] & g[28050];
assign g[44435] = a[14] & g[28051];
assign g[60818] = b[14] & g[28051];
assign g[44436] = a[14] & g[28052];
assign g[60819] = b[14] & g[28052];
assign g[44437] = a[14] & g[28053];
assign g[60820] = b[14] & g[28053];
assign g[44438] = a[14] & g[28054];
assign g[60821] = b[14] & g[28054];
assign g[44439] = a[14] & g[28055];
assign g[60822] = b[14] & g[28055];
assign g[44440] = a[14] & g[28056];
assign g[60823] = b[14] & g[28056];
assign g[44441] = a[14] & g[28057];
assign g[60824] = b[14] & g[28057];
assign g[44442] = a[14] & g[28058];
assign g[60825] = b[14] & g[28058];
assign g[44443] = a[14] & g[28059];
assign g[60826] = b[14] & g[28059];
assign g[44444] = a[14] & g[28060];
assign g[60827] = b[14] & g[28060];
assign g[44445] = a[14] & g[28061];
assign g[60828] = b[14] & g[28061];
assign g[44446] = a[14] & g[28062];
assign g[60829] = b[14] & g[28062];
assign g[44447] = a[14] & g[28063];
assign g[60830] = b[14] & g[28063];
assign g[44448] = a[14] & g[28064];
assign g[60831] = b[14] & g[28064];
assign g[44449] = a[14] & g[28065];
assign g[60832] = b[14] & g[28065];
assign g[44450] = a[14] & g[28066];
assign g[60833] = b[14] & g[28066];
assign g[44451] = a[14] & g[28067];
assign g[60834] = b[14] & g[28067];
assign g[44452] = a[14] & g[28068];
assign g[60835] = b[14] & g[28068];
assign g[44453] = a[14] & g[28069];
assign g[60836] = b[14] & g[28069];
assign g[44454] = a[14] & g[28070];
assign g[60837] = b[14] & g[28070];
assign g[44455] = a[14] & g[28071];
assign g[60838] = b[14] & g[28071];
assign g[44456] = a[14] & g[28072];
assign g[60839] = b[14] & g[28072];
assign g[44457] = a[14] & g[28073];
assign g[60840] = b[14] & g[28073];
assign g[44458] = a[14] & g[28074];
assign g[60841] = b[14] & g[28074];
assign g[44459] = a[14] & g[28075];
assign g[60842] = b[14] & g[28075];
assign g[44460] = a[14] & g[28076];
assign g[60843] = b[14] & g[28076];
assign g[44461] = a[14] & g[28077];
assign g[60844] = b[14] & g[28077];
assign g[44462] = a[14] & g[28078];
assign g[60845] = b[14] & g[28078];
assign g[44463] = a[14] & g[28079];
assign g[60846] = b[14] & g[28079];
assign g[44464] = a[14] & g[28080];
assign g[60847] = b[14] & g[28080];
assign g[44465] = a[14] & g[28081];
assign g[60848] = b[14] & g[28081];
assign g[44466] = a[14] & g[28082];
assign g[60849] = b[14] & g[28082];
assign g[44467] = a[14] & g[28083];
assign g[60850] = b[14] & g[28083];
assign g[44468] = a[14] & g[28084];
assign g[60851] = b[14] & g[28084];
assign g[44469] = a[14] & g[28085];
assign g[60852] = b[14] & g[28085];
assign g[44470] = a[14] & g[28086];
assign g[60853] = b[14] & g[28086];
assign g[44471] = a[14] & g[28087];
assign g[60854] = b[14] & g[28087];
assign g[44472] = a[14] & g[28088];
assign g[60855] = b[14] & g[28088];
assign g[44473] = a[14] & g[28089];
assign g[60856] = b[14] & g[28089];
assign g[44474] = a[14] & g[28090];
assign g[60857] = b[14] & g[28090];
assign g[44475] = a[14] & g[28091];
assign g[60858] = b[14] & g[28091];
assign g[44476] = a[14] & g[28092];
assign g[60859] = b[14] & g[28092];
assign g[44477] = a[14] & g[28093];
assign g[60860] = b[14] & g[28093];
assign g[44478] = a[14] & g[28094];
assign g[60861] = b[14] & g[28094];
assign g[44479] = a[14] & g[28095];
assign g[60862] = b[14] & g[28095];
assign g[44480] = a[14] & g[28096];
assign g[60863] = b[14] & g[28096];
assign g[44481] = a[14] & g[28097];
assign g[60864] = b[14] & g[28097];
assign g[44482] = a[14] & g[28098];
assign g[60865] = b[14] & g[28098];
assign g[44483] = a[14] & g[28099];
assign g[60866] = b[14] & g[28099];
assign g[44484] = a[14] & g[28100];
assign g[60867] = b[14] & g[28100];
assign g[44485] = a[14] & g[28101];
assign g[60868] = b[14] & g[28101];
assign g[44486] = a[14] & g[28102];
assign g[60869] = b[14] & g[28102];
assign g[44487] = a[14] & g[28103];
assign g[60870] = b[14] & g[28103];
assign g[44488] = a[14] & g[28104];
assign g[60871] = b[14] & g[28104];
assign g[44489] = a[14] & g[28105];
assign g[60872] = b[14] & g[28105];
assign g[44490] = a[14] & g[28106];
assign g[60873] = b[14] & g[28106];
assign g[44491] = a[14] & g[28107];
assign g[60874] = b[14] & g[28107];
assign g[44492] = a[14] & g[28108];
assign g[60875] = b[14] & g[28108];
assign g[44493] = a[14] & g[28109];
assign g[60876] = b[14] & g[28109];
assign g[44494] = a[14] & g[28110];
assign g[60877] = b[14] & g[28110];
assign g[44495] = a[14] & g[28111];
assign g[60878] = b[14] & g[28111];
assign g[44496] = a[14] & g[28112];
assign g[60879] = b[14] & g[28112];
assign g[44497] = a[14] & g[28113];
assign g[60880] = b[14] & g[28113];
assign g[44498] = a[14] & g[28114];
assign g[60881] = b[14] & g[28114];
assign g[44499] = a[14] & g[28115];
assign g[60882] = b[14] & g[28115];
assign g[44500] = a[14] & g[28116];
assign g[60883] = b[14] & g[28116];
assign g[44501] = a[14] & g[28117];
assign g[60884] = b[14] & g[28117];
assign g[44502] = a[14] & g[28118];
assign g[60885] = b[14] & g[28118];
assign g[44503] = a[14] & g[28119];
assign g[60886] = b[14] & g[28119];
assign g[44504] = a[14] & g[28120];
assign g[60887] = b[14] & g[28120];
assign g[44505] = a[14] & g[28121];
assign g[60888] = b[14] & g[28121];
assign g[44506] = a[14] & g[28122];
assign g[60889] = b[14] & g[28122];
assign g[44507] = a[14] & g[28123];
assign g[60890] = b[14] & g[28123];
assign g[44508] = a[14] & g[28124];
assign g[60891] = b[14] & g[28124];
assign g[44509] = a[14] & g[28125];
assign g[60892] = b[14] & g[28125];
assign g[44510] = a[14] & g[28126];
assign g[60893] = b[14] & g[28126];
assign g[44511] = a[14] & g[28127];
assign g[60894] = b[14] & g[28127];
assign g[44512] = a[14] & g[28128];
assign g[60895] = b[14] & g[28128];
assign g[44513] = a[14] & g[28129];
assign g[60896] = b[14] & g[28129];
assign g[44514] = a[14] & g[28130];
assign g[60897] = b[14] & g[28130];
assign g[44515] = a[14] & g[28131];
assign g[60898] = b[14] & g[28131];
assign g[44516] = a[14] & g[28132];
assign g[60899] = b[14] & g[28132];
assign g[44517] = a[14] & g[28133];
assign g[60900] = b[14] & g[28133];
assign g[44518] = a[14] & g[28134];
assign g[60901] = b[14] & g[28134];
assign g[44519] = a[14] & g[28135];
assign g[60902] = b[14] & g[28135];
assign g[44520] = a[14] & g[28136];
assign g[60903] = b[14] & g[28136];
assign g[44521] = a[14] & g[28137];
assign g[60904] = b[14] & g[28137];
assign g[44522] = a[14] & g[28138];
assign g[60905] = b[14] & g[28138];
assign g[44523] = a[14] & g[28139];
assign g[60906] = b[14] & g[28139];
assign g[44524] = a[14] & g[28140];
assign g[60907] = b[14] & g[28140];
assign g[44525] = a[14] & g[28141];
assign g[60908] = b[14] & g[28141];
assign g[44526] = a[14] & g[28142];
assign g[60909] = b[14] & g[28142];
assign g[44527] = a[14] & g[28143];
assign g[60910] = b[14] & g[28143];
assign g[44528] = a[14] & g[28144];
assign g[60911] = b[14] & g[28144];
assign g[44529] = a[14] & g[28145];
assign g[60912] = b[14] & g[28145];
assign g[44530] = a[14] & g[28146];
assign g[60913] = b[14] & g[28146];
assign g[44531] = a[14] & g[28147];
assign g[60914] = b[14] & g[28147];
assign g[44532] = a[14] & g[28148];
assign g[60915] = b[14] & g[28148];
assign g[44533] = a[14] & g[28149];
assign g[60916] = b[14] & g[28149];
assign g[44534] = a[14] & g[28150];
assign g[60917] = b[14] & g[28150];
assign g[44535] = a[14] & g[28151];
assign g[60918] = b[14] & g[28151];
assign g[44536] = a[14] & g[28152];
assign g[60919] = b[14] & g[28152];
assign g[44537] = a[14] & g[28153];
assign g[60920] = b[14] & g[28153];
assign g[44538] = a[14] & g[28154];
assign g[60921] = b[14] & g[28154];
assign g[44539] = a[14] & g[28155];
assign g[60922] = b[14] & g[28155];
assign g[44540] = a[14] & g[28156];
assign g[60923] = b[14] & g[28156];
assign g[44541] = a[14] & g[28157];
assign g[60924] = b[14] & g[28157];
assign g[44542] = a[14] & g[28158];
assign g[60925] = b[14] & g[28158];
assign g[44543] = a[14] & g[28159];
assign g[60926] = b[14] & g[28159];
assign g[44544] = a[14] & g[28160];
assign g[60927] = b[14] & g[28160];
assign g[44545] = a[14] & g[28161];
assign g[60928] = b[14] & g[28161];
assign g[44546] = a[14] & g[28162];
assign g[60929] = b[14] & g[28162];
assign g[44547] = a[14] & g[28163];
assign g[60930] = b[14] & g[28163];
assign g[44548] = a[14] & g[28164];
assign g[60931] = b[14] & g[28164];
assign g[44549] = a[14] & g[28165];
assign g[60932] = b[14] & g[28165];
assign g[44550] = a[14] & g[28166];
assign g[60933] = b[14] & g[28166];
assign g[44551] = a[14] & g[28167];
assign g[60934] = b[14] & g[28167];
assign g[44552] = a[14] & g[28168];
assign g[60935] = b[14] & g[28168];
assign g[44553] = a[14] & g[28169];
assign g[60936] = b[14] & g[28169];
assign g[44554] = a[14] & g[28170];
assign g[60937] = b[14] & g[28170];
assign g[44555] = a[14] & g[28171];
assign g[60938] = b[14] & g[28171];
assign g[44556] = a[14] & g[28172];
assign g[60939] = b[14] & g[28172];
assign g[44557] = a[14] & g[28173];
assign g[60940] = b[14] & g[28173];
assign g[44558] = a[14] & g[28174];
assign g[60941] = b[14] & g[28174];
assign g[44559] = a[14] & g[28175];
assign g[60942] = b[14] & g[28175];
assign g[44560] = a[14] & g[28176];
assign g[60943] = b[14] & g[28176];
assign g[44561] = a[14] & g[28177];
assign g[60944] = b[14] & g[28177];
assign g[44562] = a[14] & g[28178];
assign g[60945] = b[14] & g[28178];
assign g[44563] = a[14] & g[28179];
assign g[60946] = b[14] & g[28179];
assign g[44564] = a[14] & g[28180];
assign g[60947] = b[14] & g[28180];
assign g[44565] = a[14] & g[28181];
assign g[60948] = b[14] & g[28181];
assign g[44566] = a[14] & g[28182];
assign g[60949] = b[14] & g[28182];
assign g[44567] = a[14] & g[28183];
assign g[60950] = b[14] & g[28183];
assign g[44568] = a[14] & g[28184];
assign g[60951] = b[14] & g[28184];
assign g[44569] = a[14] & g[28185];
assign g[60952] = b[14] & g[28185];
assign g[44570] = a[14] & g[28186];
assign g[60953] = b[14] & g[28186];
assign g[44571] = a[14] & g[28187];
assign g[60954] = b[14] & g[28187];
assign g[44572] = a[14] & g[28188];
assign g[60955] = b[14] & g[28188];
assign g[44573] = a[14] & g[28189];
assign g[60956] = b[14] & g[28189];
assign g[44574] = a[14] & g[28190];
assign g[60957] = b[14] & g[28190];
assign g[44575] = a[14] & g[28191];
assign g[60958] = b[14] & g[28191];
assign g[44576] = a[14] & g[28192];
assign g[60959] = b[14] & g[28192];
assign g[44577] = a[14] & g[28193];
assign g[60960] = b[14] & g[28193];
assign g[44578] = a[14] & g[28194];
assign g[60961] = b[14] & g[28194];
assign g[44579] = a[14] & g[28195];
assign g[60962] = b[14] & g[28195];
assign g[44580] = a[14] & g[28196];
assign g[60963] = b[14] & g[28196];
assign g[44581] = a[14] & g[28197];
assign g[60964] = b[14] & g[28197];
assign g[44582] = a[14] & g[28198];
assign g[60965] = b[14] & g[28198];
assign g[44583] = a[14] & g[28199];
assign g[60966] = b[14] & g[28199];
assign g[44584] = a[14] & g[28200];
assign g[60967] = b[14] & g[28200];
assign g[44585] = a[14] & g[28201];
assign g[60968] = b[14] & g[28201];
assign g[44586] = a[14] & g[28202];
assign g[60969] = b[14] & g[28202];
assign g[44587] = a[14] & g[28203];
assign g[60970] = b[14] & g[28203];
assign g[44588] = a[14] & g[28204];
assign g[60971] = b[14] & g[28204];
assign g[44589] = a[14] & g[28205];
assign g[60972] = b[14] & g[28205];
assign g[44590] = a[14] & g[28206];
assign g[60973] = b[14] & g[28206];
assign g[44591] = a[14] & g[28207];
assign g[60974] = b[14] & g[28207];
assign g[44592] = a[14] & g[28208];
assign g[60975] = b[14] & g[28208];
assign g[44593] = a[14] & g[28209];
assign g[60976] = b[14] & g[28209];
assign g[44594] = a[14] & g[28210];
assign g[60977] = b[14] & g[28210];
assign g[44595] = a[14] & g[28211];
assign g[60978] = b[14] & g[28211];
assign g[44596] = a[14] & g[28212];
assign g[60979] = b[14] & g[28212];
assign g[44597] = a[14] & g[28213];
assign g[60980] = b[14] & g[28213];
assign g[44598] = a[14] & g[28214];
assign g[60981] = b[14] & g[28214];
assign g[44599] = a[14] & g[28215];
assign g[60982] = b[14] & g[28215];
assign g[44600] = a[14] & g[28216];
assign g[60983] = b[14] & g[28216];
assign g[44601] = a[14] & g[28217];
assign g[60984] = b[14] & g[28217];
assign g[44602] = a[14] & g[28218];
assign g[60985] = b[14] & g[28218];
assign g[44603] = a[14] & g[28219];
assign g[60986] = b[14] & g[28219];
assign g[44604] = a[14] & g[28220];
assign g[60987] = b[14] & g[28220];
assign g[44605] = a[14] & g[28221];
assign g[60988] = b[14] & g[28221];
assign g[44606] = a[14] & g[28222];
assign g[60989] = b[14] & g[28222];
assign g[44607] = a[14] & g[28223];
assign g[60990] = b[14] & g[28223];
assign g[44608] = a[14] & g[28224];
assign g[60991] = b[14] & g[28224];
assign g[44609] = a[14] & g[28225];
assign g[60992] = b[14] & g[28225];
assign g[44610] = a[14] & g[28226];
assign g[60993] = b[14] & g[28226];
assign g[44611] = a[14] & g[28227];
assign g[60994] = b[14] & g[28227];
assign g[44612] = a[14] & g[28228];
assign g[60995] = b[14] & g[28228];
assign g[44613] = a[14] & g[28229];
assign g[60996] = b[14] & g[28229];
assign g[44614] = a[14] & g[28230];
assign g[60997] = b[14] & g[28230];
assign g[44615] = a[14] & g[28231];
assign g[60998] = b[14] & g[28231];
assign g[44616] = a[14] & g[28232];
assign g[60999] = b[14] & g[28232];
assign g[44617] = a[14] & g[28233];
assign g[61000] = b[14] & g[28233];
assign g[44618] = a[14] & g[28234];
assign g[61001] = b[14] & g[28234];
assign g[44619] = a[14] & g[28235];
assign g[61002] = b[14] & g[28235];
assign g[44620] = a[14] & g[28236];
assign g[61003] = b[14] & g[28236];
assign g[44621] = a[14] & g[28237];
assign g[61004] = b[14] & g[28237];
assign g[44622] = a[14] & g[28238];
assign g[61005] = b[14] & g[28238];
assign g[44623] = a[14] & g[28239];
assign g[61006] = b[14] & g[28239];
assign g[44624] = a[14] & g[28240];
assign g[61007] = b[14] & g[28240];
assign g[44625] = a[14] & g[28241];
assign g[61008] = b[14] & g[28241];
assign g[44626] = a[14] & g[28242];
assign g[61009] = b[14] & g[28242];
assign g[44627] = a[14] & g[28243];
assign g[61010] = b[14] & g[28243];
assign g[44628] = a[14] & g[28244];
assign g[61011] = b[14] & g[28244];
assign g[44629] = a[14] & g[28245];
assign g[61012] = b[14] & g[28245];
assign g[44630] = a[14] & g[28246];
assign g[61013] = b[14] & g[28246];
assign g[44631] = a[14] & g[28247];
assign g[61014] = b[14] & g[28247];
assign g[44632] = a[14] & g[28248];
assign g[61015] = b[14] & g[28248];
assign g[44633] = a[14] & g[28249];
assign g[61016] = b[14] & g[28249];
assign g[44634] = a[14] & g[28250];
assign g[61017] = b[14] & g[28250];
assign g[44635] = a[14] & g[28251];
assign g[61018] = b[14] & g[28251];
assign g[44636] = a[14] & g[28252];
assign g[61019] = b[14] & g[28252];
assign g[44637] = a[14] & g[28253];
assign g[61020] = b[14] & g[28253];
assign g[44638] = a[14] & g[28254];
assign g[61021] = b[14] & g[28254];
assign g[44639] = a[14] & g[28255];
assign g[61022] = b[14] & g[28255];
assign g[44640] = a[14] & g[28256];
assign g[61023] = b[14] & g[28256];
assign g[44641] = a[14] & g[28257];
assign g[61024] = b[14] & g[28257];
assign g[44642] = a[14] & g[28258];
assign g[61025] = b[14] & g[28258];
assign g[44643] = a[14] & g[28259];
assign g[61026] = b[14] & g[28259];
assign g[44644] = a[14] & g[28260];
assign g[61027] = b[14] & g[28260];
assign g[44645] = a[14] & g[28261];
assign g[61028] = b[14] & g[28261];
assign g[44646] = a[14] & g[28262];
assign g[61029] = b[14] & g[28262];
assign g[44647] = a[14] & g[28263];
assign g[61030] = b[14] & g[28263];
assign g[44648] = a[14] & g[28264];
assign g[61031] = b[14] & g[28264];
assign g[44649] = a[14] & g[28265];
assign g[61032] = b[14] & g[28265];
assign g[44650] = a[14] & g[28266];
assign g[61033] = b[14] & g[28266];
assign g[44651] = a[14] & g[28267];
assign g[61034] = b[14] & g[28267];
assign g[44652] = a[14] & g[28268];
assign g[61035] = b[14] & g[28268];
assign g[44653] = a[14] & g[28269];
assign g[61036] = b[14] & g[28269];
assign g[44654] = a[14] & g[28270];
assign g[61037] = b[14] & g[28270];
assign g[44655] = a[14] & g[28271];
assign g[61038] = b[14] & g[28271];
assign g[44656] = a[14] & g[28272];
assign g[61039] = b[14] & g[28272];
assign g[44657] = a[14] & g[28273];
assign g[61040] = b[14] & g[28273];
assign g[44658] = a[14] & g[28274];
assign g[61041] = b[14] & g[28274];
assign g[44659] = a[14] & g[28275];
assign g[61042] = b[14] & g[28275];
assign g[44660] = a[14] & g[28276];
assign g[61043] = b[14] & g[28276];
assign g[44661] = a[14] & g[28277];
assign g[61044] = b[14] & g[28277];
assign g[44662] = a[14] & g[28278];
assign g[61045] = b[14] & g[28278];
assign g[44663] = a[14] & g[28279];
assign g[61046] = b[14] & g[28279];
assign g[44664] = a[14] & g[28280];
assign g[61047] = b[14] & g[28280];
assign g[44665] = a[14] & g[28281];
assign g[61048] = b[14] & g[28281];
assign g[44666] = a[14] & g[28282];
assign g[61049] = b[14] & g[28282];
assign g[44667] = a[14] & g[28283];
assign g[61050] = b[14] & g[28283];
assign g[44668] = a[14] & g[28284];
assign g[61051] = b[14] & g[28284];
assign g[44669] = a[14] & g[28285];
assign g[61052] = b[14] & g[28285];
assign g[44670] = a[14] & g[28286];
assign g[61053] = b[14] & g[28286];
assign g[44671] = a[14] & g[28287];
assign g[61054] = b[14] & g[28287];
assign g[44672] = a[14] & g[28288];
assign g[61055] = b[14] & g[28288];
assign g[44673] = a[14] & g[28289];
assign g[61056] = b[14] & g[28289];
assign g[44674] = a[14] & g[28290];
assign g[61057] = b[14] & g[28290];
assign g[44675] = a[14] & g[28291];
assign g[61058] = b[14] & g[28291];
assign g[44676] = a[14] & g[28292];
assign g[61059] = b[14] & g[28292];
assign g[44677] = a[14] & g[28293];
assign g[61060] = b[14] & g[28293];
assign g[44678] = a[14] & g[28294];
assign g[61061] = b[14] & g[28294];
assign g[44679] = a[14] & g[28295];
assign g[61062] = b[14] & g[28295];
assign g[44680] = a[14] & g[28296];
assign g[61063] = b[14] & g[28296];
assign g[44681] = a[14] & g[28297];
assign g[61064] = b[14] & g[28297];
assign g[44682] = a[14] & g[28298];
assign g[61065] = b[14] & g[28298];
assign g[44683] = a[14] & g[28299];
assign g[61066] = b[14] & g[28299];
assign g[44684] = a[14] & g[28300];
assign g[61067] = b[14] & g[28300];
assign g[44685] = a[14] & g[28301];
assign g[61068] = b[14] & g[28301];
assign g[44686] = a[14] & g[28302];
assign g[61069] = b[14] & g[28302];
assign g[44687] = a[14] & g[28303];
assign g[61070] = b[14] & g[28303];
assign g[44688] = a[14] & g[28304];
assign g[61071] = b[14] & g[28304];
assign g[44689] = a[14] & g[28305];
assign g[61072] = b[14] & g[28305];
assign g[44690] = a[14] & g[28306];
assign g[61073] = b[14] & g[28306];
assign g[44691] = a[14] & g[28307];
assign g[61074] = b[14] & g[28307];
assign g[44692] = a[14] & g[28308];
assign g[61075] = b[14] & g[28308];
assign g[44693] = a[14] & g[28309];
assign g[61076] = b[14] & g[28309];
assign g[44694] = a[14] & g[28310];
assign g[61077] = b[14] & g[28310];
assign g[44695] = a[14] & g[28311];
assign g[61078] = b[14] & g[28311];
assign g[44696] = a[14] & g[28312];
assign g[61079] = b[14] & g[28312];
assign g[44697] = a[14] & g[28313];
assign g[61080] = b[14] & g[28313];
assign g[44698] = a[14] & g[28314];
assign g[61081] = b[14] & g[28314];
assign g[44699] = a[14] & g[28315];
assign g[61082] = b[14] & g[28315];
assign g[44700] = a[14] & g[28316];
assign g[61083] = b[14] & g[28316];
assign g[44701] = a[14] & g[28317];
assign g[61084] = b[14] & g[28317];
assign g[44702] = a[14] & g[28318];
assign g[61085] = b[14] & g[28318];
assign g[44703] = a[14] & g[28319];
assign g[61086] = b[14] & g[28319];
assign g[44704] = a[14] & g[28320];
assign g[61087] = b[14] & g[28320];
assign g[44705] = a[14] & g[28321];
assign g[61088] = b[14] & g[28321];
assign g[44706] = a[14] & g[28322];
assign g[61089] = b[14] & g[28322];
assign g[44707] = a[14] & g[28323];
assign g[61090] = b[14] & g[28323];
assign g[44708] = a[14] & g[28324];
assign g[61091] = b[14] & g[28324];
assign g[44709] = a[14] & g[28325];
assign g[61092] = b[14] & g[28325];
assign g[44710] = a[14] & g[28326];
assign g[61093] = b[14] & g[28326];
assign g[44711] = a[14] & g[28327];
assign g[61094] = b[14] & g[28327];
assign g[44712] = a[14] & g[28328];
assign g[61095] = b[14] & g[28328];
assign g[44713] = a[14] & g[28329];
assign g[61096] = b[14] & g[28329];
assign g[44714] = a[14] & g[28330];
assign g[61097] = b[14] & g[28330];
assign g[44715] = a[14] & g[28331];
assign g[61098] = b[14] & g[28331];
assign g[44716] = a[14] & g[28332];
assign g[61099] = b[14] & g[28332];
assign g[44717] = a[14] & g[28333];
assign g[61100] = b[14] & g[28333];
assign g[44718] = a[14] & g[28334];
assign g[61101] = b[14] & g[28334];
assign g[44719] = a[14] & g[28335];
assign g[61102] = b[14] & g[28335];
assign g[44720] = a[14] & g[28336];
assign g[61103] = b[14] & g[28336];
assign g[44721] = a[14] & g[28337];
assign g[61104] = b[14] & g[28337];
assign g[44722] = a[14] & g[28338];
assign g[61105] = b[14] & g[28338];
assign g[44723] = a[14] & g[28339];
assign g[61106] = b[14] & g[28339];
assign g[44724] = a[14] & g[28340];
assign g[61107] = b[14] & g[28340];
assign g[44725] = a[14] & g[28341];
assign g[61108] = b[14] & g[28341];
assign g[44726] = a[14] & g[28342];
assign g[61109] = b[14] & g[28342];
assign g[44727] = a[14] & g[28343];
assign g[61110] = b[14] & g[28343];
assign g[44728] = a[14] & g[28344];
assign g[61111] = b[14] & g[28344];
assign g[44729] = a[14] & g[28345];
assign g[61112] = b[14] & g[28345];
assign g[44730] = a[14] & g[28346];
assign g[61113] = b[14] & g[28346];
assign g[44731] = a[14] & g[28347];
assign g[61114] = b[14] & g[28347];
assign g[44732] = a[14] & g[28348];
assign g[61115] = b[14] & g[28348];
assign g[44733] = a[14] & g[28349];
assign g[61116] = b[14] & g[28349];
assign g[44734] = a[14] & g[28350];
assign g[61117] = b[14] & g[28350];
assign g[44735] = a[14] & g[28351];
assign g[61118] = b[14] & g[28351];
assign g[44736] = a[14] & g[28352];
assign g[61119] = b[14] & g[28352];
assign g[44737] = a[14] & g[28353];
assign g[61120] = b[14] & g[28353];
assign g[44738] = a[14] & g[28354];
assign g[61121] = b[14] & g[28354];
assign g[44739] = a[14] & g[28355];
assign g[61122] = b[14] & g[28355];
assign g[44740] = a[14] & g[28356];
assign g[61123] = b[14] & g[28356];
assign g[44741] = a[14] & g[28357];
assign g[61124] = b[14] & g[28357];
assign g[44742] = a[14] & g[28358];
assign g[61125] = b[14] & g[28358];
assign g[44743] = a[14] & g[28359];
assign g[61126] = b[14] & g[28359];
assign g[44744] = a[14] & g[28360];
assign g[61127] = b[14] & g[28360];
assign g[44745] = a[14] & g[28361];
assign g[61128] = b[14] & g[28361];
assign g[44746] = a[14] & g[28362];
assign g[61129] = b[14] & g[28362];
assign g[44747] = a[14] & g[28363];
assign g[61130] = b[14] & g[28363];
assign g[44748] = a[14] & g[28364];
assign g[61131] = b[14] & g[28364];
assign g[44749] = a[14] & g[28365];
assign g[61132] = b[14] & g[28365];
assign g[44750] = a[14] & g[28366];
assign g[61133] = b[14] & g[28366];
assign g[44751] = a[14] & g[28367];
assign g[61134] = b[14] & g[28367];
assign g[44752] = a[14] & g[28368];
assign g[61135] = b[14] & g[28368];
assign g[44753] = a[14] & g[28369];
assign g[61136] = b[14] & g[28369];
assign g[44754] = a[14] & g[28370];
assign g[61137] = b[14] & g[28370];
assign g[44755] = a[14] & g[28371];
assign g[61138] = b[14] & g[28371];
assign g[44756] = a[14] & g[28372];
assign g[61139] = b[14] & g[28372];
assign g[44757] = a[14] & g[28373];
assign g[61140] = b[14] & g[28373];
assign g[44758] = a[14] & g[28374];
assign g[61141] = b[14] & g[28374];
assign g[44759] = a[14] & g[28375];
assign g[61142] = b[14] & g[28375];
assign g[44760] = a[14] & g[28376];
assign g[61143] = b[14] & g[28376];
assign g[44761] = a[14] & g[28377];
assign g[61144] = b[14] & g[28377];
assign g[44762] = a[14] & g[28378];
assign g[61145] = b[14] & g[28378];
assign g[44763] = a[14] & g[28379];
assign g[61146] = b[14] & g[28379];
assign g[44764] = a[14] & g[28380];
assign g[61147] = b[14] & g[28380];
assign g[44765] = a[14] & g[28381];
assign g[61148] = b[14] & g[28381];
assign g[44766] = a[14] & g[28382];
assign g[61149] = b[14] & g[28382];
assign g[44767] = a[14] & g[28383];
assign g[61150] = b[14] & g[28383];
assign g[44768] = a[14] & g[28384];
assign g[61151] = b[14] & g[28384];
assign g[44769] = a[14] & g[28385];
assign g[61152] = b[14] & g[28385];
assign g[44770] = a[14] & g[28386];
assign g[61153] = b[14] & g[28386];
assign g[44771] = a[14] & g[28387];
assign g[61154] = b[14] & g[28387];
assign g[44772] = a[14] & g[28388];
assign g[61155] = b[14] & g[28388];
assign g[44773] = a[14] & g[28389];
assign g[61156] = b[14] & g[28389];
assign g[44774] = a[14] & g[28390];
assign g[61157] = b[14] & g[28390];
assign g[44775] = a[14] & g[28391];
assign g[61158] = b[14] & g[28391];
assign g[44776] = a[14] & g[28392];
assign g[61159] = b[14] & g[28392];
assign g[44777] = a[14] & g[28393];
assign g[61160] = b[14] & g[28393];
assign g[44778] = a[14] & g[28394];
assign g[61161] = b[14] & g[28394];
assign g[44779] = a[14] & g[28395];
assign g[61162] = b[14] & g[28395];
assign g[44780] = a[14] & g[28396];
assign g[61163] = b[14] & g[28396];
assign g[44781] = a[14] & g[28397];
assign g[61164] = b[14] & g[28397];
assign g[44782] = a[14] & g[28398];
assign g[61165] = b[14] & g[28398];
assign g[44783] = a[14] & g[28399];
assign g[61166] = b[14] & g[28399];
assign g[44784] = a[14] & g[28400];
assign g[61167] = b[14] & g[28400];
assign g[44785] = a[14] & g[28401];
assign g[61168] = b[14] & g[28401];
assign g[44786] = a[14] & g[28402];
assign g[61169] = b[14] & g[28402];
assign g[44787] = a[14] & g[28403];
assign g[61170] = b[14] & g[28403];
assign g[44788] = a[14] & g[28404];
assign g[61171] = b[14] & g[28404];
assign g[44789] = a[14] & g[28405];
assign g[61172] = b[14] & g[28405];
assign g[44790] = a[14] & g[28406];
assign g[61173] = b[14] & g[28406];
assign g[44791] = a[14] & g[28407];
assign g[61174] = b[14] & g[28407];
assign g[44792] = a[14] & g[28408];
assign g[61175] = b[14] & g[28408];
assign g[44793] = a[14] & g[28409];
assign g[61176] = b[14] & g[28409];
assign g[44794] = a[14] & g[28410];
assign g[61177] = b[14] & g[28410];
assign g[44795] = a[14] & g[28411];
assign g[61178] = b[14] & g[28411];
assign g[44796] = a[14] & g[28412];
assign g[61179] = b[14] & g[28412];
assign g[44797] = a[14] & g[28413];
assign g[61180] = b[14] & g[28413];
assign g[44798] = a[14] & g[28414];
assign g[61181] = b[14] & g[28414];
assign g[44799] = a[14] & g[28415];
assign g[61182] = b[14] & g[28415];
assign g[44800] = a[14] & g[28416];
assign g[61183] = b[14] & g[28416];
assign g[44801] = a[14] & g[28417];
assign g[61184] = b[14] & g[28417];
assign g[44802] = a[14] & g[28418];
assign g[61185] = b[14] & g[28418];
assign g[44803] = a[14] & g[28419];
assign g[61186] = b[14] & g[28419];
assign g[44804] = a[14] & g[28420];
assign g[61187] = b[14] & g[28420];
assign g[44805] = a[14] & g[28421];
assign g[61188] = b[14] & g[28421];
assign g[44806] = a[14] & g[28422];
assign g[61189] = b[14] & g[28422];
assign g[44807] = a[14] & g[28423];
assign g[61190] = b[14] & g[28423];
assign g[44808] = a[14] & g[28424];
assign g[61191] = b[14] & g[28424];
assign g[44809] = a[14] & g[28425];
assign g[61192] = b[14] & g[28425];
assign g[44810] = a[14] & g[28426];
assign g[61193] = b[14] & g[28426];
assign g[44811] = a[14] & g[28427];
assign g[61194] = b[14] & g[28427];
assign g[44812] = a[14] & g[28428];
assign g[61195] = b[14] & g[28428];
assign g[44813] = a[14] & g[28429];
assign g[61196] = b[14] & g[28429];
assign g[44814] = a[14] & g[28430];
assign g[61197] = b[14] & g[28430];
assign g[44815] = a[14] & g[28431];
assign g[61198] = b[14] & g[28431];
assign g[44816] = a[14] & g[28432];
assign g[61199] = b[14] & g[28432];
assign g[44817] = a[14] & g[28433];
assign g[61200] = b[14] & g[28433];
assign g[44818] = a[14] & g[28434];
assign g[61201] = b[14] & g[28434];
assign g[44819] = a[14] & g[28435];
assign g[61202] = b[14] & g[28435];
assign g[44820] = a[14] & g[28436];
assign g[61203] = b[14] & g[28436];
assign g[44821] = a[14] & g[28437];
assign g[61204] = b[14] & g[28437];
assign g[44822] = a[14] & g[28438];
assign g[61205] = b[14] & g[28438];
assign g[44823] = a[14] & g[28439];
assign g[61206] = b[14] & g[28439];
assign g[44824] = a[14] & g[28440];
assign g[61207] = b[14] & g[28440];
assign g[44825] = a[14] & g[28441];
assign g[61208] = b[14] & g[28441];
assign g[44826] = a[14] & g[28442];
assign g[61209] = b[14] & g[28442];
assign g[44827] = a[14] & g[28443];
assign g[61210] = b[14] & g[28443];
assign g[44828] = a[14] & g[28444];
assign g[61211] = b[14] & g[28444];
assign g[44829] = a[14] & g[28445];
assign g[61212] = b[14] & g[28445];
assign g[44830] = a[14] & g[28446];
assign g[61213] = b[14] & g[28446];
assign g[44831] = a[14] & g[28447];
assign g[61214] = b[14] & g[28447];
assign g[44832] = a[14] & g[28448];
assign g[61215] = b[14] & g[28448];
assign g[44833] = a[14] & g[28449];
assign g[61216] = b[14] & g[28449];
assign g[44834] = a[14] & g[28450];
assign g[61217] = b[14] & g[28450];
assign g[44835] = a[14] & g[28451];
assign g[61218] = b[14] & g[28451];
assign g[44836] = a[14] & g[28452];
assign g[61219] = b[14] & g[28452];
assign g[44837] = a[14] & g[28453];
assign g[61220] = b[14] & g[28453];
assign g[44838] = a[14] & g[28454];
assign g[61221] = b[14] & g[28454];
assign g[44839] = a[14] & g[28455];
assign g[61222] = b[14] & g[28455];
assign g[44840] = a[14] & g[28456];
assign g[61223] = b[14] & g[28456];
assign g[44841] = a[14] & g[28457];
assign g[61224] = b[14] & g[28457];
assign g[44842] = a[14] & g[28458];
assign g[61225] = b[14] & g[28458];
assign g[44843] = a[14] & g[28459];
assign g[61226] = b[14] & g[28459];
assign g[44844] = a[14] & g[28460];
assign g[61227] = b[14] & g[28460];
assign g[44845] = a[14] & g[28461];
assign g[61228] = b[14] & g[28461];
assign g[44846] = a[14] & g[28462];
assign g[61229] = b[14] & g[28462];
assign g[44847] = a[14] & g[28463];
assign g[61230] = b[14] & g[28463];
assign g[44848] = a[14] & g[28464];
assign g[61231] = b[14] & g[28464];
assign g[44849] = a[14] & g[28465];
assign g[61232] = b[14] & g[28465];
assign g[44850] = a[14] & g[28466];
assign g[61233] = b[14] & g[28466];
assign g[44851] = a[14] & g[28467];
assign g[61234] = b[14] & g[28467];
assign g[44852] = a[14] & g[28468];
assign g[61235] = b[14] & g[28468];
assign g[44853] = a[14] & g[28469];
assign g[61236] = b[14] & g[28469];
assign g[44854] = a[14] & g[28470];
assign g[61237] = b[14] & g[28470];
assign g[44855] = a[14] & g[28471];
assign g[61238] = b[14] & g[28471];
assign g[44856] = a[14] & g[28472];
assign g[61239] = b[14] & g[28472];
assign g[44857] = a[14] & g[28473];
assign g[61240] = b[14] & g[28473];
assign g[44858] = a[14] & g[28474];
assign g[61241] = b[14] & g[28474];
assign g[44859] = a[14] & g[28475];
assign g[61242] = b[14] & g[28475];
assign g[44860] = a[14] & g[28476];
assign g[61243] = b[14] & g[28476];
assign g[44861] = a[14] & g[28477];
assign g[61244] = b[14] & g[28477];
assign g[44862] = a[14] & g[28478];
assign g[61245] = b[14] & g[28478];
assign g[44863] = a[14] & g[28479];
assign g[61246] = b[14] & g[28479];
assign g[44864] = a[14] & g[28480];
assign g[61247] = b[14] & g[28480];
assign g[44865] = a[14] & g[28481];
assign g[61248] = b[14] & g[28481];
assign g[44866] = a[14] & g[28482];
assign g[61249] = b[14] & g[28482];
assign g[44867] = a[14] & g[28483];
assign g[61250] = b[14] & g[28483];
assign g[44868] = a[14] & g[28484];
assign g[61251] = b[14] & g[28484];
assign g[44869] = a[14] & g[28485];
assign g[61252] = b[14] & g[28485];
assign g[44870] = a[14] & g[28486];
assign g[61253] = b[14] & g[28486];
assign g[44871] = a[14] & g[28487];
assign g[61254] = b[14] & g[28487];
assign g[44872] = a[14] & g[28488];
assign g[61255] = b[14] & g[28488];
assign g[44873] = a[14] & g[28489];
assign g[61256] = b[14] & g[28489];
assign g[44874] = a[14] & g[28490];
assign g[61257] = b[14] & g[28490];
assign g[44875] = a[14] & g[28491];
assign g[61258] = b[14] & g[28491];
assign g[44876] = a[14] & g[28492];
assign g[61259] = b[14] & g[28492];
assign g[44877] = a[14] & g[28493];
assign g[61260] = b[14] & g[28493];
assign g[44878] = a[14] & g[28494];
assign g[61261] = b[14] & g[28494];
assign g[44879] = a[14] & g[28495];
assign g[61262] = b[14] & g[28495];
assign g[44880] = a[14] & g[28496];
assign g[61263] = b[14] & g[28496];
assign g[44881] = a[14] & g[28497];
assign g[61264] = b[14] & g[28497];
assign g[44882] = a[14] & g[28498];
assign g[61265] = b[14] & g[28498];
assign g[44883] = a[14] & g[28499];
assign g[61266] = b[14] & g[28499];
assign g[44884] = a[14] & g[28500];
assign g[61267] = b[14] & g[28500];
assign g[44885] = a[14] & g[28501];
assign g[61268] = b[14] & g[28501];
assign g[44886] = a[14] & g[28502];
assign g[61269] = b[14] & g[28502];
assign g[44887] = a[14] & g[28503];
assign g[61270] = b[14] & g[28503];
assign g[44888] = a[14] & g[28504];
assign g[61271] = b[14] & g[28504];
assign g[44889] = a[14] & g[28505];
assign g[61272] = b[14] & g[28505];
assign g[44890] = a[14] & g[28506];
assign g[61273] = b[14] & g[28506];
assign g[44891] = a[14] & g[28507];
assign g[61274] = b[14] & g[28507];
assign g[44892] = a[14] & g[28508];
assign g[61275] = b[14] & g[28508];
assign g[44893] = a[14] & g[28509];
assign g[61276] = b[14] & g[28509];
assign g[44894] = a[14] & g[28510];
assign g[61277] = b[14] & g[28510];
assign g[44895] = a[14] & g[28511];
assign g[61278] = b[14] & g[28511];
assign g[44896] = a[14] & g[28512];
assign g[61279] = b[14] & g[28512];
assign g[44897] = a[14] & g[28513];
assign g[61280] = b[14] & g[28513];
assign g[44898] = a[14] & g[28514];
assign g[61281] = b[14] & g[28514];
assign g[44899] = a[14] & g[28515];
assign g[61282] = b[14] & g[28515];
assign g[44900] = a[14] & g[28516];
assign g[61283] = b[14] & g[28516];
assign g[44901] = a[14] & g[28517];
assign g[61284] = b[14] & g[28517];
assign g[44902] = a[14] & g[28518];
assign g[61285] = b[14] & g[28518];
assign g[44903] = a[14] & g[28519];
assign g[61286] = b[14] & g[28519];
assign g[44904] = a[14] & g[28520];
assign g[61287] = b[14] & g[28520];
assign g[44905] = a[14] & g[28521];
assign g[61288] = b[14] & g[28521];
assign g[44906] = a[14] & g[28522];
assign g[61289] = b[14] & g[28522];
assign g[44907] = a[14] & g[28523];
assign g[61290] = b[14] & g[28523];
assign g[44908] = a[14] & g[28524];
assign g[61291] = b[14] & g[28524];
assign g[44909] = a[14] & g[28525];
assign g[61292] = b[14] & g[28525];
assign g[44910] = a[14] & g[28526];
assign g[61293] = b[14] & g[28526];
assign g[44911] = a[14] & g[28527];
assign g[61294] = b[14] & g[28527];
assign g[44912] = a[14] & g[28528];
assign g[61295] = b[14] & g[28528];
assign g[44913] = a[14] & g[28529];
assign g[61296] = b[14] & g[28529];
assign g[44914] = a[14] & g[28530];
assign g[61297] = b[14] & g[28530];
assign g[44915] = a[14] & g[28531];
assign g[61298] = b[14] & g[28531];
assign g[44916] = a[14] & g[28532];
assign g[61299] = b[14] & g[28532];
assign g[44917] = a[14] & g[28533];
assign g[61300] = b[14] & g[28533];
assign g[44918] = a[14] & g[28534];
assign g[61301] = b[14] & g[28534];
assign g[44919] = a[14] & g[28535];
assign g[61302] = b[14] & g[28535];
assign g[44920] = a[14] & g[28536];
assign g[61303] = b[14] & g[28536];
assign g[44921] = a[14] & g[28537];
assign g[61304] = b[14] & g[28537];
assign g[44922] = a[14] & g[28538];
assign g[61305] = b[14] & g[28538];
assign g[44923] = a[14] & g[28539];
assign g[61306] = b[14] & g[28539];
assign g[44924] = a[14] & g[28540];
assign g[61307] = b[14] & g[28540];
assign g[44925] = a[14] & g[28541];
assign g[61308] = b[14] & g[28541];
assign g[44926] = a[14] & g[28542];
assign g[61309] = b[14] & g[28542];
assign g[44927] = a[14] & g[28543];
assign g[61310] = b[14] & g[28543];
assign g[44928] = a[14] & g[28544];
assign g[61311] = b[14] & g[28544];
assign g[44929] = a[14] & g[28545];
assign g[61312] = b[14] & g[28545];
assign g[44930] = a[14] & g[28546];
assign g[61313] = b[14] & g[28546];
assign g[44931] = a[14] & g[28547];
assign g[61314] = b[14] & g[28547];
assign g[44932] = a[14] & g[28548];
assign g[61315] = b[14] & g[28548];
assign g[44933] = a[14] & g[28549];
assign g[61316] = b[14] & g[28549];
assign g[44934] = a[14] & g[28550];
assign g[61317] = b[14] & g[28550];
assign g[44935] = a[14] & g[28551];
assign g[61318] = b[14] & g[28551];
assign g[44936] = a[14] & g[28552];
assign g[61319] = b[14] & g[28552];
assign g[44937] = a[14] & g[28553];
assign g[61320] = b[14] & g[28553];
assign g[44938] = a[14] & g[28554];
assign g[61321] = b[14] & g[28554];
assign g[44939] = a[14] & g[28555];
assign g[61322] = b[14] & g[28555];
assign g[44940] = a[14] & g[28556];
assign g[61323] = b[14] & g[28556];
assign g[44941] = a[14] & g[28557];
assign g[61324] = b[14] & g[28557];
assign g[44942] = a[14] & g[28558];
assign g[61325] = b[14] & g[28558];
assign g[44943] = a[14] & g[28559];
assign g[61326] = b[14] & g[28559];
assign g[44944] = a[14] & g[28560];
assign g[61327] = b[14] & g[28560];
assign g[44945] = a[14] & g[28561];
assign g[61328] = b[14] & g[28561];
assign g[44946] = a[14] & g[28562];
assign g[61329] = b[14] & g[28562];
assign g[44947] = a[14] & g[28563];
assign g[61330] = b[14] & g[28563];
assign g[44948] = a[14] & g[28564];
assign g[61331] = b[14] & g[28564];
assign g[44949] = a[14] & g[28565];
assign g[61332] = b[14] & g[28565];
assign g[44950] = a[14] & g[28566];
assign g[61333] = b[14] & g[28566];
assign g[44951] = a[14] & g[28567];
assign g[61334] = b[14] & g[28567];
assign g[44952] = a[14] & g[28568];
assign g[61335] = b[14] & g[28568];
assign g[44953] = a[14] & g[28569];
assign g[61336] = b[14] & g[28569];
assign g[44954] = a[14] & g[28570];
assign g[61337] = b[14] & g[28570];
assign g[44955] = a[14] & g[28571];
assign g[61338] = b[14] & g[28571];
assign g[44956] = a[14] & g[28572];
assign g[61339] = b[14] & g[28572];
assign g[44957] = a[14] & g[28573];
assign g[61340] = b[14] & g[28573];
assign g[44958] = a[14] & g[28574];
assign g[61341] = b[14] & g[28574];
assign g[44959] = a[14] & g[28575];
assign g[61342] = b[14] & g[28575];
assign g[44960] = a[14] & g[28576];
assign g[61343] = b[14] & g[28576];
assign g[44961] = a[14] & g[28577];
assign g[61344] = b[14] & g[28577];
assign g[44962] = a[14] & g[28578];
assign g[61345] = b[14] & g[28578];
assign g[44963] = a[14] & g[28579];
assign g[61346] = b[14] & g[28579];
assign g[44964] = a[14] & g[28580];
assign g[61347] = b[14] & g[28580];
assign g[44965] = a[14] & g[28581];
assign g[61348] = b[14] & g[28581];
assign g[44966] = a[14] & g[28582];
assign g[61349] = b[14] & g[28582];
assign g[44967] = a[14] & g[28583];
assign g[61350] = b[14] & g[28583];
assign g[44968] = a[14] & g[28584];
assign g[61351] = b[14] & g[28584];
assign g[44969] = a[14] & g[28585];
assign g[61352] = b[14] & g[28585];
assign g[44970] = a[14] & g[28586];
assign g[61353] = b[14] & g[28586];
assign g[44971] = a[14] & g[28587];
assign g[61354] = b[14] & g[28587];
assign g[44972] = a[14] & g[28588];
assign g[61355] = b[14] & g[28588];
assign g[44973] = a[14] & g[28589];
assign g[61356] = b[14] & g[28589];
assign g[44974] = a[14] & g[28590];
assign g[61357] = b[14] & g[28590];
assign g[44975] = a[14] & g[28591];
assign g[61358] = b[14] & g[28591];
assign g[44976] = a[14] & g[28592];
assign g[61359] = b[14] & g[28592];
assign g[44977] = a[14] & g[28593];
assign g[61360] = b[14] & g[28593];
assign g[44978] = a[14] & g[28594];
assign g[61361] = b[14] & g[28594];
assign g[44979] = a[14] & g[28595];
assign g[61362] = b[14] & g[28595];
assign g[44980] = a[14] & g[28596];
assign g[61363] = b[14] & g[28596];
assign g[44981] = a[14] & g[28597];
assign g[61364] = b[14] & g[28597];
assign g[44982] = a[14] & g[28598];
assign g[61365] = b[14] & g[28598];
assign g[44983] = a[14] & g[28599];
assign g[61366] = b[14] & g[28599];
assign g[44984] = a[14] & g[28600];
assign g[61367] = b[14] & g[28600];
assign g[44985] = a[14] & g[28601];
assign g[61368] = b[14] & g[28601];
assign g[44986] = a[14] & g[28602];
assign g[61369] = b[14] & g[28602];
assign g[44987] = a[14] & g[28603];
assign g[61370] = b[14] & g[28603];
assign g[44988] = a[14] & g[28604];
assign g[61371] = b[14] & g[28604];
assign g[44989] = a[14] & g[28605];
assign g[61372] = b[14] & g[28605];
assign g[44990] = a[14] & g[28606];
assign g[61373] = b[14] & g[28606];
assign g[44991] = a[14] & g[28607];
assign g[61374] = b[14] & g[28607];
assign g[44992] = a[14] & g[28608];
assign g[61375] = b[14] & g[28608];
assign g[44993] = a[14] & g[28609];
assign g[61376] = b[14] & g[28609];
assign g[44994] = a[14] & g[28610];
assign g[61377] = b[14] & g[28610];
assign g[44995] = a[14] & g[28611];
assign g[61378] = b[14] & g[28611];
assign g[44996] = a[14] & g[28612];
assign g[61379] = b[14] & g[28612];
assign g[44997] = a[14] & g[28613];
assign g[61380] = b[14] & g[28613];
assign g[44998] = a[14] & g[28614];
assign g[61381] = b[14] & g[28614];
assign g[44999] = a[14] & g[28615];
assign g[61382] = b[14] & g[28615];
assign g[45000] = a[14] & g[28616];
assign g[61383] = b[14] & g[28616];
assign g[45001] = a[14] & g[28617];
assign g[61384] = b[14] & g[28617];
assign g[45002] = a[14] & g[28618];
assign g[61385] = b[14] & g[28618];
assign g[45003] = a[14] & g[28619];
assign g[61386] = b[14] & g[28619];
assign g[45004] = a[14] & g[28620];
assign g[61387] = b[14] & g[28620];
assign g[45005] = a[14] & g[28621];
assign g[61388] = b[14] & g[28621];
assign g[45006] = a[14] & g[28622];
assign g[61389] = b[14] & g[28622];
assign g[45007] = a[14] & g[28623];
assign g[61390] = b[14] & g[28623];
assign g[45008] = a[14] & g[28624];
assign g[61391] = b[14] & g[28624];
assign g[45009] = a[14] & g[28625];
assign g[61392] = b[14] & g[28625];
assign g[45010] = a[14] & g[28626];
assign g[61393] = b[14] & g[28626];
assign g[45011] = a[14] & g[28627];
assign g[61394] = b[14] & g[28627];
assign g[45012] = a[14] & g[28628];
assign g[61395] = b[14] & g[28628];
assign g[45013] = a[14] & g[28629];
assign g[61396] = b[14] & g[28629];
assign g[45014] = a[14] & g[28630];
assign g[61397] = b[14] & g[28630];
assign g[45015] = a[14] & g[28631];
assign g[61398] = b[14] & g[28631];
assign g[45016] = a[14] & g[28632];
assign g[61399] = b[14] & g[28632];
assign g[45017] = a[14] & g[28633];
assign g[61400] = b[14] & g[28633];
assign g[45018] = a[14] & g[28634];
assign g[61401] = b[14] & g[28634];
assign g[45019] = a[14] & g[28635];
assign g[61402] = b[14] & g[28635];
assign g[45020] = a[14] & g[28636];
assign g[61403] = b[14] & g[28636];
assign g[45021] = a[14] & g[28637];
assign g[61404] = b[14] & g[28637];
assign g[45022] = a[14] & g[28638];
assign g[61405] = b[14] & g[28638];
assign g[45023] = a[14] & g[28639];
assign g[61406] = b[14] & g[28639];
assign g[45024] = a[14] & g[28640];
assign g[61407] = b[14] & g[28640];
assign g[45025] = a[14] & g[28641];
assign g[61408] = b[14] & g[28641];
assign g[45026] = a[14] & g[28642];
assign g[61409] = b[14] & g[28642];
assign g[45027] = a[14] & g[28643];
assign g[61410] = b[14] & g[28643];
assign g[45028] = a[14] & g[28644];
assign g[61411] = b[14] & g[28644];
assign g[45029] = a[14] & g[28645];
assign g[61412] = b[14] & g[28645];
assign g[45030] = a[14] & g[28646];
assign g[61413] = b[14] & g[28646];
assign g[45031] = a[14] & g[28647];
assign g[61414] = b[14] & g[28647];
assign g[45032] = a[14] & g[28648];
assign g[61415] = b[14] & g[28648];
assign g[45033] = a[14] & g[28649];
assign g[61416] = b[14] & g[28649];
assign g[45034] = a[14] & g[28650];
assign g[61417] = b[14] & g[28650];
assign g[45035] = a[14] & g[28651];
assign g[61418] = b[14] & g[28651];
assign g[45036] = a[14] & g[28652];
assign g[61419] = b[14] & g[28652];
assign g[45037] = a[14] & g[28653];
assign g[61420] = b[14] & g[28653];
assign g[45038] = a[14] & g[28654];
assign g[61421] = b[14] & g[28654];
assign g[45039] = a[14] & g[28655];
assign g[61422] = b[14] & g[28655];
assign g[45040] = a[14] & g[28656];
assign g[61423] = b[14] & g[28656];
assign g[45041] = a[14] & g[28657];
assign g[61424] = b[14] & g[28657];
assign g[45042] = a[14] & g[28658];
assign g[61425] = b[14] & g[28658];
assign g[45043] = a[14] & g[28659];
assign g[61426] = b[14] & g[28659];
assign g[45044] = a[14] & g[28660];
assign g[61427] = b[14] & g[28660];
assign g[45045] = a[14] & g[28661];
assign g[61428] = b[14] & g[28661];
assign g[45046] = a[14] & g[28662];
assign g[61429] = b[14] & g[28662];
assign g[45047] = a[14] & g[28663];
assign g[61430] = b[14] & g[28663];
assign g[45048] = a[14] & g[28664];
assign g[61431] = b[14] & g[28664];
assign g[45049] = a[14] & g[28665];
assign g[61432] = b[14] & g[28665];
assign g[45050] = a[14] & g[28666];
assign g[61433] = b[14] & g[28666];
assign g[45051] = a[14] & g[28667];
assign g[61434] = b[14] & g[28667];
assign g[45052] = a[14] & g[28668];
assign g[61435] = b[14] & g[28668];
assign g[45053] = a[14] & g[28669];
assign g[61436] = b[14] & g[28669];
assign g[45054] = a[14] & g[28670];
assign g[61437] = b[14] & g[28670];
assign g[45055] = a[14] & g[28671];
assign g[61438] = b[14] & g[28671];
assign g[45056] = a[14] & g[28672];
assign g[61439] = b[14] & g[28672];
assign g[45057] = a[14] & g[28673];
assign g[61440] = b[14] & g[28673];
assign g[45058] = a[14] & g[28674];
assign g[61441] = b[14] & g[28674];
assign g[45059] = a[14] & g[28675];
assign g[61442] = b[14] & g[28675];
assign g[45060] = a[14] & g[28676];
assign g[61443] = b[14] & g[28676];
assign g[45061] = a[14] & g[28677];
assign g[61444] = b[14] & g[28677];
assign g[45062] = a[14] & g[28678];
assign g[61445] = b[14] & g[28678];
assign g[45063] = a[14] & g[28679];
assign g[61446] = b[14] & g[28679];
assign g[45064] = a[14] & g[28680];
assign g[61447] = b[14] & g[28680];
assign g[45065] = a[14] & g[28681];
assign g[61448] = b[14] & g[28681];
assign g[45066] = a[14] & g[28682];
assign g[61449] = b[14] & g[28682];
assign g[45067] = a[14] & g[28683];
assign g[61450] = b[14] & g[28683];
assign g[45068] = a[14] & g[28684];
assign g[61451] = b[14] & g[28684];
assign g[45069] = a[14] & g[28685];
assign g[61452] = b[14] & g[28685];
assign g[45070] = a[14] & g[28686];
assign g[61453] = b[14] & g[28686];
assign g[45071] = a[14] & g[28687];
assign g[61454] = b[14] & g[28687];
assign g[45072] = a[14] & g[28688];
assign g[61455] = b[14] & g[28688];
assign g[45073] = a[14] & g[28689];
assign g[61456] = b[14] & g[28689];
assign g[45074] = a[14] & g[28690];
assign g[61457] = b[14] & g[28690];
assign g[45075] = a[14] & g[28691];
assign g[61458] = b[14] & g[28691];
assign g[45076] = a[14] & g[28692];
assign g[61459] = b[14] & g[28692];
assign g[45077] = a[14] & g[28693];
assign g[61460] = b[14] & g[28693];
assign g[45078] = a[14] & g[28694];
assign g[61461] = b[14] & g[28694];
assign g[45079] = a[14] & g[28695];
assign g[61462] = b[14] & g[28695];
assign g[45080] = a[14] & g[28696];
assign g[61463] = b[14] & g[28696];
assign g[45081] = a[14] & g[28697];
assign g[61464] = b[14] & g[28697];
assign g[45082] = a[14] & g[28698];
assign g[61465] = b[14] & g[28698];
assign g[45083] = a[14] & g[28699];
assign g[61466] = b[14] & g[28699];
assign g[45084] = a[14] & g[28700];
assign g[61467] = b[14] & g[28700];
assign g[45085] = a[14] & g[28701];
assign g[61468] = b[14] & g[28701];
assign g[45086] = a[14] & g[28702];
assign g[61469] = b[14] & g[28702];
assign g[45087] = a[14] & g[28703];
assign g[61470] = b[14] & g[28703];
assign g[45088] = a[14] & g[28704];
assign g[61471] = b[14] & g[28704];
assign g[45089] = a[14] & g[28705];
assign g[61472] = b[14] & g[28705];
assign g[45090] = a[14] & g[28706];
assign g[61473] = b[14] & g[28706];
assign g[45091] = a[14] & g[28707];
assign g[61474] = b[14] & g[28707];
assign g[45092] = a[14] & g[28708];
assign g[61475] = b[14] & g[28708];
assign g[45093] = a[14] & g[28709];
assign g[61476] = b[14] & g[28709];
assign g[45094] = a[14] & g[28710];
assign g[61477] = b[14] & g[28710];
assign g[45095] = a[14] & g[28711];
assign g[61478] = b[14] & g[28711];
assign g[45096] = a[14] & g[28712];
assign g[61479] = b[14] & g[28712];
assign g[45097] = a[14] & g[28713];
assign g[61480] = b[14] & g[28713];
assign g[45098] = a[14] & g[28714];
assign g[61481] = b[14] & g[28714];
assign g[45099] = a[14] & g[28715];
assign g[61482] = b[14] & g[28715];
assign g[45100] = a[14] & g[28716];
assign g[61483] = b[14] & g[28716];
assign g[45101] = a[14] & g[28717];
assign g[61484] = b[14] & g[28717];
assign g[45102] = a[14] & g[28718];
assign g[61485] = b[14] & g[28718];
assign g[45103] = a[14] & g[28719];
assign g[61486] = b[14] & g[28719];
assign g[45104] = a[14] & g[28720];
assign g[61487] = b[14] & g[28720];
assign g[45105] = a[14] & g[28721];
assign g[61488] = b[14] & g[28721];
assign g[45106] = a[14] & g[28722];
assign g[61489] = b[14] & g[28722];
assign g[45107] = a[14] & g[28723];
assign g[61490] = b[14] & g[28723];
assign g[45108] = a[14] & g[28724];
assign g[61491] = b[14] & g[28724];
assign g[45109] = a[14] & g[28725];
assign g[61492] = b[14] & g[28725];
assign g[45110] = a[14] & g[28726];
assign g[61493] = b[14] & g[28726];
assign g[45111] = a[14] & g[28727];
assign g[61494] = b[14] & g[28727];
assign g[45112] = a[14] & g[28728];
assign g[61495] = b[14] & g[28728];
assign g[45113] = a[14] & g[28729];
assign g[61496] = b[14] & g[28729];
assign g[45114] = a[14] & g[28730];
assign g[61497] = b[14] & g[28730];
assign g[45115] = a[14] & g[28731];
assign g[61498] = b[14] & g[28731];
assign g[45116] = a[14] & g[28732];
assign g[61499] = b[14] & g[28732];
assign g[45117] = a[14] & g[28733];
assign g[61500] = b[14] & g[28733];
assign g[45118] = a[14] & g[28734];
assign g[61501] = b[14] & g[28734];
assign g[45119] = a[14] & g[28735];
assign g[61502] = b[14] & g[28735];
assign g[45120] = a[14] & g[28736];
assign g[61503] = b[14] & g[28736];
assign g[45121] = a[14] & g[28737];
assign g[61504] = b[14] & g[28737];
assign g[45122] = a[14] & g[28738];
assign g[61505] = b[14] & g[28738];
assign g[45123] = a[14] & g[28739];
assign g[61506] = b[14] & g[28739];
assign g[45124] = a[14] & g[28740];
assign g[61507] = b[14] & g[28740];
assign g[45125] = a[14] & g[28741];
assign g[61508] = b[14] & g[28741];
assign g[45126] = a[14] & g[28742];
assign g[61509] = b[14] & g[28742];
assign g[45127] = a[14] & g[28743];
assign g[61510] = b[14] & g[28743];
assign g[45128] = a[14] & g[28744];
assign g[61511] = b[14] & g[28744];
assign g[45129] = a[14] & g[28745];
assign g[61512] = b[14] & g[28745];
assign g[45130] = a[14] & g[28746];
assign g[61513] = b[14] & g[28746];
assign g[45131] = a[14] & g[28747];
assign g[61514] = b[14] & g[28747];
assign g[45132] = a[14] & g[28748];
assign g[61515] = b[14] & g[28748];
assign g[45133] = a[14] & g[28749];
assign g[61516] = b[14] & g[28749];
assign g[45134] = a[14] & g[28750];
assign g[61517] = b[14] & g[28750];
assign g[45135] = a[14] & g[28751];
assign g[61518] = b[14] & g[28751];
assign g[45136] = a[14] & g[28752];
assign g[61519] = b[14] & g[28752];
assign g[45137] = a[14] & g[28753];
assign g[61520] = b[14] & g[28753];
assign g[45138] = a[14] & g[28754];
assign g[61521] = b[14] & g[28754];
assign g[45139] = a[14] & g[28755];
assign g[61522] = b[14] & g[28755];
assign g[45140] = a[14] & g[28756];
assign g[61523] = b[14] & g[28756];
assign g[45141] = a[14] & g[28757];
assign g[61524] = b[14] & g[28757];
assign g[45142] = a[14] & g[28758];
assign g[61525] = b[14] & g[28758];
assign g[45143] = a[14] & g[28759];
assign g[61526] = b[14] & g[28759];
assign g[45144] = a[14] & g[28760];
assign g[61527] = b[14] & g[28760];
assign g[45145] = a[14] & g[28761];
assign g[61528] = b[14] & g[28761];
assign g[45146] = a[14] & g[28762];
assign g[61529] = b[14] & g[28762];
assign g[45147] = a[14] & g[28763];
assign g[61530] = b[14] & g[28763];
assign g[45148] = a[14] & g[28764];
assign g[61531] = b[14] & g[28764];
assign g[45149] = a[14] & g[28765];
assign g[61532] = b[14] & g[28765];
assign g[45150] = a[14] & g[28766];
assign g[61533] = b[14] & g[28766];
assign g[45151] = a[14] & g[28767];
assign g[61534] = b[14] & g[28767];
assign g[45152] = a[14] & g[28768];
assign g[61535] = b[14] & g[28768];
assign g[45153] = a[14] & g[28769];
assign g[61536] = b[14] & g[28769];
assign g[45154] = a[14] & g[28770];
assign g[61537] = b[14] & g[28770];
assign g[45155] = a[14] & g[28771];
assign g[61538] = b[14] & g[28771];
assign g[45156] = a[14] & g[28772];
assign g[61539] = b[14] & g[28772];
assign g[45157] = a[14] & g[28773];
assign g[61540] = b[14] & g[28773];
assign g[45158] = a[14] & g[28774];
assign g[61541] = b[14] & g[28774];
assign g[45159] = a[14] & g[28775];
assign g[61542] = b[14] & g[28775];
assign g[45160] = a[14] & g[28776];
assign g[61543] = b[14] & g[28776];
assign g[45161] = a[14] & g[28777];
assign g[61544] = b[14] & g[28777];
assign g[45162] = a[14] & g[28778];
assign g[61545] = b[14] & g[28778];
assign g[45163] = a[14] & g[28779];
assign g[61546] = b[14] & g[28779];
assign g[45164] = a[14] & g[28780];
assign g[61547] = b[14] & g[28780];
assign g[45165] = a[14] & g[28781];
assign g[61548] = b[14] & g[28781];
assign g[45166] = a[14] & g[28782];
assign g[61549] = b[14] & g[28782];
assign g[45167] = a[14] & g[28783];
assign g[61550] = b[14] & g[28783];
assign g[45168] = a[14] & g[28784];
assign g[61551] = b[14] & g[28784];
assign g[45169] = a[14] & g[28785];
assign g[61552] = b[14] & g[28785];
assign g[45170] = a[14] & g[28786];
assign g[61553] = b[14] & g[28786];
assign g[45171] = a[14] & g[28787];
assign g[61554] = b[14] & g[28787];
assign g[45172] = a[14] & g[28788];
assign g[61555] = b[14] & g[28788];
assign g[45173] = a[14] & g[28789];
assign g[61556] = b[14] & g[28789];
assign g[45174] = a[14] & g[28790];
assign g[61557] = b[14] & g[28790];
assign g[45175] = a[14] & g[28791];
assign g[61558] = b[14] & g[28791];
assign g[45176] = a[14] & g[28792];
assign g[61559] = b[14] & g[28792];
assign g[45177] = a[14] & g[28793];
assign g[61560] = b[14] & g[28793];
assign g[45178] = a[14] & g[28794];
assign g[61561] = b[14] & g[28794];
assign g[45179] = a[14] & g[28795];
assign g[61562] = b[14] & g[28795];
assign g[45180] = a[14] & g[28796];
assign g[61563] = b[14] & g[28796];
assign g[45181] = a[14] & g[28797];
assign g[61564] = b[14] & g[28797];
assign g[45182] = a[14] & g[28798];
assign g[61565] = b[14] & g[28798];
assign g[45183] = a[14] & g[28799];
assign g[61566] = b[14] & g[28799];
assign g[45184] = a[14] & g[28800];
assign g[61567] = b[14] & g[28800];
assign g[45185] = a[14] & g[28801];
assign g[61568] = b[14] & g[28801];
assign g[45186] = a[14] & g[28802];
assign g[61569] = b[14] & g[28802];
assign g[45187] = a[14] & g[28803];
assign g[61570] = b[14] & g[28803];
assign g[45188] = a[14] & g[28804];
assign g[61571] = b[14] & g[28804];
assign g[45189] = a[14] & g[28805];
assign g[61572] = b[14] & g[28805];
assign g[45190] = a[14] & g[28806];
assign g[61573] = b[14] & g[28806];
assign g[45191] = a[14] & g[28807];
assign g[61574] = b[14] & g[28807];
assign g[45192] = a[14] & g[28808];
assign g[61575] = b[14] & g[28808];
assign g[45193] = a[14] & g[28809];
assign g[61576] = b[14] & g[28809];
assign g[45194] = a[14] & g[28810];
assign g[61577] = b[14] & g[28810];
assign g[45195] = a[14] & g[28811];
assign g[61578] = b[14] & g[28811];
assign g[45196] = a[14] & g[28812];
assign g[61579] = b[14] & g[28812];
assign g[45197] = a[14] & g[28813];
assign g[61580] = b[14] & g[28813];
assign g[45198] = a[14] & g[28814];
assign g[61581] = b[14] & g[28814];
assign g[45199] = a[14] & g[28815];
assign g[61582] = b[14] & g[28815];
assign g[45200] = a[14] & g[28816];
assign g[61583] = b[14] & g[28816];
assign g[45201] = a[14] & g[28817];
assign g[61584] = b[14] & g[28817];
assign g[45202] = a[14] & g[28818];
assign g[61585] = b[14] & g[28818];
assign g[45203] = a[14] & g[28819];
assign g[61586] = b[14] & g[28819];
assign g[45204] = a[14] & g[28820];
assign g[61587] = b[14] & g[28820];
assign g[45205] = a[14] & g[28821];
assign g[61588] = b[14] & g[28821];
assign g[45206] = a[14] & g[28822];
assign g[61589] = b[14] & g[28822];
assign g[45207] = a[14] & g[28823];
assign g[61590] = b[14] & g[28823];
assign g[45208] = a[14] & g[28824];
assign g[61591] = b[14] & g[28824];
assign g[45209] = a[14] & g[28825];
assign g[61592] = b[14] & g[28825];
assign g[45210] = a[14] & g[28826];
assign g[61593] = b[14] & g[28826];
assign g[45211] = a[14] & g[28827];
assign g[61594] = b[14] & g[28827];
assign g[45212] = a[14] & g[28828];
assign g[61595] = b[14] & g[28828];
assign g[45213] = a[14] & g[28829];
assign g[61596] = b[14] & g[28829];
assign g[45214] = a[14] & g[28830];
assign g[61597] = b[14] & g[28830];
assign g[45215] = a[14] & g[28831];
assign g[61598] = b[14] & g[28831];
assign g[45216] = a[14] & g[28832];
assign g[61599] = b[14] & g[28832];
assign g[45217] = a[14] & g[28833];
assign g[61600] = b[14] & g[28833];
assign g[45218] = a[14] & g[28834];
assign g[61601] = b[14] & g[28834];
assign g[45219] = a[14] & g[28835];
assign g[61602] = b[14] & g[28835];
assign g[45220] = a[14] & g[28836];
assign g[61603] = b[14] & g[28836];
assign g[45221] = a[14] & g[28837];
assign g[61604] = b[14] & g[28837];
assign g[45222] = a[14] & g[28838];
assign g[61605] = b[14] & g[28838];
assign g[45223] = a[14] & g[28839];
assign g[61606] = b[14] & g[28839];
assign g[45224] = a[14] & g[28840];
assign g[61607] = b[14] & g[28840];
assign g[45225] = a[14] & g[28841];
assign g[61608] = b[14] & g[28841];
assign g[45226] = a[14] & g[28842];
assign g[61609] = b[14] & g[28842];
assign g[45227] = a[14] & g[28843];
assign g[61610] = b[14] & g[28843];
assign g[45228] = a[14] & g[28844];
assign g[61611] = b[14] & g[28844];
assign g[45229] = a[14] & g[28845];
assign g[61612] = b[14] & g[28845];
assign g[45230] = a[14] & g[28846];
assign g[61613] = b[14] & g[28846];
assign g[45231] = a[14] & g[28847];
assign g[61614] = b[14] & g[28847];
assign g[45232] = a[14] & g[28848];
assign g[61615] = b[14] & g[28848];
assign g[45233] = a[14] & g[28849];
assign g[61616] = b[14] & g[28849];
assign g[45234] = a[14] & g[28850];
assign g[61617] = b[14] & g[28850];
assign g[45235] = a[14] & g[28851];
assign g[61618] = b[14] & g[28851];
assign g[45236] = a[14] & g[28852];
assign g[61619] = b[14] & g[28852];
assign g[45237] = a[14] & g[28853];
assign g[61620] = b[14] & g[28853];
assign g[45238] = a[14] & g[28854];
assign g[61621] = b[14] & g[28854];
assign g[45239] = a[14] & g[28855];
assign g[61622] = b[14] & g[28855];
assign g[45240] = a[14] & g[28856];
assign g[61623] = b[14] & g[28856];
assign g[45241] = a[14] & g[28857];
assign g[61624] = b[14] & g[28857];
assign g[45242] = a[14] & g[28858];
assign g[61625] = b[14] & g[28858];
assign g[45243] = a[14] & g[28859];
assign g[61626] = b[14] & g[28859];
assign g[45244] = a[14] & g[28860];
assign g[61627] = b[14] & g[28860];
assign g[45245] = a[14] & g[28861];
assign g[61628] = b[14] & g[28861];
assign g[45246] = a[14] & g[28862];
assign g[61629] = b[14] & g[28862];
assign g[45247] = a[14] & g[28863];
assign g[61630] = b[14] & g[28863];
assign g[45248] = a[14] & g[28864];
assign g[61631] = b[14] & g[28864];
assign g[45249] = a[14] & g[28865];
assign g[61632] = b[14] & g[28865];
assign g[45250] = a[14] & g[28866];
assign g[61633] = b[14] & g[28866];
assign g[45251] = a[14] & g[28867];
assign g[61634] = b[14] & g[28867];
assign g[45252] = a[14] & g[28868];
assign g[61635] = b[14] & g[28868];
assign g[45253] = a[14] & g[28869];
assign g[61636] = b[14] & g[28869];
assign g[45254] = a[14] & g[28870];
assign g[61637] = b[14] & g[28870];
assign g[45255] = a[14] & g[28871];
assign g[61638] = b[14] & g[28871];
assign g[45256] = a[14] & g[28872];
assign g[61639] = b[14] & g[28872];
assign g[45257] = a[14] & g[28873];
assign g[61640] = b[14] & g[28873];
assign g[45258] = a[14] & g[28874];
assign g[61641] = b[14] & g[28874];
assign g[45259] = a[14] & g[28875];
assign g[61642] = b[14] & g[28875];
assign g[45260] = a[14] & g[28876];
assign g[61643] = b[14] & g[28876];
assign g[45261] = a[14] & g[28877];
assign g[61644] = b[14] & g[28877];
assign g[45262] = a[14] & g[28878];
assign g[61645] = b[14] & g[28878];
assign g[45263] = a[14] & g[28879];
assign g[61646] = b[14] & g[28879];
assign g[45264] = a[14] & g[28880];
assign g[61647] = b[14] & g[28880];
assign g[45265] = a[14] & g[28881];
assign g[61648] = b[14] & g[28881];
assign g[45266] = a[14] & g[28882];
assign g[61649] = b[14] & g[28882];
assign g[45267] = a[14] & g[28883];
assign g[61650] = b[14] & g[28883];
assign g[45268] = a[14] & g[28884];
assign g[61651] = b[14] & g[28884];
assign g[45269] = a[14] & g[28885];
assign g[61652] = b[14] & g[28885];
assign g[45270] = a[14] & g[28886];
assign g[61653] = b[14] & g[28886];
assign g[45271] = a[14] & g[28887];
assign g[61654] = b[14] & g[28887];
assign g[45272] = a[14] & g[28888];
assign g[61655] = b[14] & g[28888];
assign g[45273] = a[14] & g[28889];
assign g[61656] = b[14] & g[28889];
assign g[45274] = a[14] & g[28890];
assign g[61657] = b[14] & g[28890];
assign g[45275] = a[14] & g[28891];
assign g[61658] = b[14] & g[28891];
assign g[45276] = a[14] & g[28892];
assign g[61659] = b[14] & g[28892];
assign g[45277] = a[14] & g[28893];
assign g[61660] = b[14] & g[28893];
assign g[45278] = a[14] & g[28894];
assign g[61661] = b[14] & g[28894];
assign g[45279] = a[14] & g[28895];
assign g[61662] = b[14] & g[28895];
assign g[45280] = a[14] & g[28896];
assign g[61663] = b[14] & g[28896];
assign g[45281] = a[14] & g[28897];
assign g[61664] = b[14] & g[28897];
assign g[45282] = a[14] & g[28898];
assign g[61665] = b[14] & g[28898];
assign g[45283] = a[14] & g[28899];
assign g[61666] = b[14] & g[28899];
assign g[45284] = a[14] & g[28900];
assign g[61667] = b[14] & g[28900];
assign g[45285] = a[14] & g[28901];
assign g[61668] = b[14] & g[28901];
assign g[45286] = a[14] & g[28902];
assign g[61669] = b[14] & g[28902];
assign g[45287] = a[14] & g[28903];
assign g[61670] = b[14] & g[28903];
assign g[45288] = a[14] & g[28904];
assign g[61671] = b[14] & g[28904];
assign g[45289] = a[14] & g[28905];
assign g[61672] = b[14] & g[28905];
assign g[45290] = a[14] & g[28906];
assign g[61673] = b[14] & g[28906];
assign g[45291] = a[14] & g[28907];
assign g[61674] = b[14] & g[28907];
assign g[45292] = a[14] & g[28908];
assign g[61675] = b[14] & g[28908];
assign g[45293] = a[14] & g[28909];
assign g[61676] = b[14] & g[28909];
assign g[45294] = a[14] & g[28910];
assign g[61677] = b[14] & g[28910];
assign g[45295] = a[14] & g[28911];
assign g[61678] = b[14] & g[28911];
assign g[45296] = a[14] & g[28912];
assign g[61679] = b[14] & g[28912];
assign g[45297] = a[14] & g[28913];
assign g[61680] = b[14] & g[28913];
assign g[45298] = a[14] & g[28914];
assign g[61681] = b[14] & g[28914];
assign g[45299] = a[14] & g[28915];
assign g[61682] = b[14] & g[28915];
assign g[45300] = a[14] & g[28916];
assign g[61683] = b[14] & g[28916];
assign g[45301] = a[14] & g[28917];
assign g[61684] = b[14] & g[28917];
assign g[45302] = a[14] & g[28918];
assign g[61685] = b[14] & g[28918];
assign g[45303] = a[14] & g[28919];
assign g[61686] = b[14] & g[28919];
assign g[45304] = a[14] & g[28920];
assign g[61687] = b[14] & g[28920];
assign g[45305] = a[14] & g[28921];
assign g[61688] = b[14] & g[28921];
assign g[45306] = a[14] & g[28922];
assign g[61689] = b[14] & g[28922];
assign g[45307] = a[14] & g[28923];
assign g[61690] = b[14] & g[28923];
assign g[45308] = a[14] & g[28924];
assign g[61691] = b[14] & g[28924];
assign g[45309] = a[14] & g[28925];
assign g[61692] = b[14] & g[28925];
assign g[45310] = a[14] & g[28926];
assign g[61693] = b[14] & g[28926];
assign g[45311] = a[14] & g[28927];
assign g[61694] = b[14] & g[28927];
assign g[45312] = a[14] & g[28928];
assign g[61695] = b[14] & g[28928];
assign g[45313] = a[14] & g[28929];
assign g[61696] = b[14] & g[28929];
assign g[45314] = a[14] & g[28930];
assign g[61697] = b[14] & g[28930];
assign g[45315] = a[14] & g[28931];
assign g[61698] = b[14] & g[28931];
assign g[45316] = a[14] & g[28932];
assign g[61699] = b[14] & g[28932];
assign g[45317] = a[14] & g[28933];
assign g[61700] = b[14] & g[28933];
assign g[45318] = a[14] & g[28934];
assign g[61701] = b[14] & g[28934];
assign g[45319] = a[14] & g[28935];
assign g[61702] = b[14] & g[28935];
assign g[45320] = a[14] & g[28936];
assign g[61703] = b[14] & g[28936];
assign g[45321] = a[14] & g[28937];
assign g[61704] = b[14] & g[28937];
assign g[45322] = a[14] & g[28938];
assign g[61705] = b[14] & g[28938];
assign g[45323] = a[14] & g[28939];
assign g[61706] = b[14] & g[28939];
assign g[45324] = a[14] & g[28940];
assign g[61707] = b[14] & g[28940];
assign g[45325] = a[14] & g[28941];
assign g[61708] = b[14] & g[28941];
assign g[45326] = a[14] & g[28942];
assign g[61709] = b[14] & g[28942];
assign g[45327] = a[14] & g[28943];
assign g[61710] = b[14] & g[28943];
assign g[45328] = a[14] & g[28944];
assign g[61711] = b[14] & g[28944];
assign g[45329] = a[14] & g[28945];
assign g[61712] = b[14] & g[28945];
assign g[45330] = a[14] & g[28946];
assign g[61713] = b[14] & g[28946];
assign g[45331] = a[14] & g[28947];
assign g[61714] = b[14] & g[28947];
assign g[45332] = a[14] & g[28948];
assign g[61715] = b[14] & g[28948];
assign g[45333] = a[14] & g[28949];
assign g[61716] = b[14] & g[28949];
assign g[45334] = a[14] & g[28950];
assign g[61717] = b[14] & g[28950];
assign g[45335] = a[14] & g[28951];
assign g[61718] = b[14] & g[28951];
assign g[45336] = a[14] & g[28952];
assign g[61719] = b[14] & g[28952];
assign g[45337] = a[14] & g[28953];
assign g[61720] = b[14] & g[28953];
assign g[45338] = a[14] & g[28954];
assign g[61721] = b[14] & g[28954];
assign g[45339] = a[14] & g[28955];
assign g[61722] = b[14] & g[28955];
assign g[45340] = a[14] & g[28956];
assign g[61723] = b[14] & g[28956];
assign g[45341] = a[14] & g[28957];
assign g[61724] = b[14] & g[28957];
assign g[45342] = a[14] & g[28958];
assign g[61725] = b[14] & g[28958];
assign g[45343] = a[14] & g[28959];
assign g[61726] = b[14] & g[28959];
assign g[45344] = a[14] & g[28960];
assign g[61727] = b[14] & g[28960];
assign g[45345] = a[14] & g[28961];
assign g[61728] = b[14] & g[28961];
assign g[45346] = a[14] & g[28962];
assign g[61729] = b[14] & g[28962];
assign g[45347] = a[14] & g[28963];
assign g[61730] = b[14] & g[28963];
assign g[45348] = a[14] & g[28964];
assign g[61731] = b[14] & g[28964];
assign g[45349] = a[14] & g[28965];
assign g[61732] = b[14] & g[28965];
assign g[45350] = a[14] & g[28966];
assign g[61733] = b[14] & g[28966];
assign g[45351] = a[14] & g[28967];
assign g[61734] = b[14] & g[28967];
assign g[45352] = a[14] & g[28968];
assign g[61735] = b[14] & g[28968];
assign g[45353] = a[14] & g[28969];
assign g[61736] = b[14] & g[28969];
assign g[45354] = a[14] & g[28970];
assign g[61737] = b[14] & g[28970];
assign g[45355] = a[14] & g[28971];
assign g[61738] = b[14] & g[28971];
assign g[45356] = a[14] & g[28972];
assign g[61739] = b[14] & g[28972];
assign g[45357] = a[14] & g[28973];
assign g[61740] = b[14] & g[28973];
assign g[45358] = a[14] & g[28974];
assign g[61741] = b[14] & g[28974];
assign g[45359] = a[14] & g[28975];
assign g[61742] = b[14] & g[28975];
assign g[45360] = a[14] & g[28976];
assign g[61743] = b[14] & g[28976];
assign g[45361] = a[14] & g[28977];
assign g[61744] = b[14] & g[28977];
assign g[45362] = a[14] & g[28978];
assign g[61745] = b[14] & g[28978];
assign g[45363] = a[14] & g[28979];
assign g[61746] = b[14] & g[28979];
assign g[45364] = a[14] & g[28980];
assign g[61747] = b[14] & g[28980];
assign g[45365] = a[14] & g[28981];
assign g[61748] = b[14] & g[28981];
assign g[45366] = a[14] & g[28982];
assign g[61749] = b[14] & g[28982];
assign g[45367] = a[14] & g[28983];
assign g[61750] = b[14] & g[28983];
assign g[45368] = a[14] & g[28984];
assign g[61751] = b[14] & g[28984];
assign g[45369] = a[14] & g[28985];
assign g[61752] = b[14] & g[28985];
assign g[45370] = a[14] & g[28986];
assign g[61753] = b[14] & g[28986];
assign g[45371] = a[14] & g[28987];
assign g[61754] = b[14] & g[28987];
assign g[45372] = a[14] & g[28988];
assign g[61755] = b[14] & g[28988];
assign g[45373] = a[14] & g[28989];
assign g[61756] = b[14] & g[28989];
assign g[45374] = a[14] & g[28990];
assign g[61757] = b[14] & g[28990];
assign g[45375] = a[14] & g[28991];
assign g[61758] = b[14] & g[28991];
assign g[45376] = a[14] & g[28992];
assign g[61759] = b[14] & g[28992];
assign g[45377] = a[14] & g[28993];
assign g[61760] = b[14] & g[28993];
assign g[45378] = a[14] & g[28994];
assign g[61761] = b[14] & g[28994];
assign g[45379] = a[14] & g[28995];
assign g[61762] = b[14] & g[28995];
assign g[45380] = a[14] & g[28996];
assign g[61763] = b[14] & g[28996];
assign g[45381] = a[14] & g[28997];
assign g[61764] = b[14] & g[28997];
assign g[45382] = a[14] & g[28998];
assign g[61765] = b[14] & g[28998];
assign g[45383] = a[14] & g[28999];
assign g[61766] = b[14] & g[28999];
assign g[45384] = a[14] & g[29000];
assign g[61767] = b[14] & g[29000];
assign g[45385] = a[14] & g[29001];
assign g[61768] = b[14] & g[29001];
assign g[45386] = a[14] & g[29002];
assign g[61769] = b[14] & g[29002];
assign g[45387] = a[14] & g[29003];
assign g[61770] = b[14] & g[29003];
assign g[45388] = a[14] & g[29004];
assign g[61771] = b[14] & g[29004];
assign g[45389] = a[14] & g[29005];
assign g[61772] = b[14] & g[29005];
assign g[45390] = a[14] & g[29006];
assign g[61773] = b[14] & g[29006];
assign g[45391] = a[14] & g[29007];
assign g[61774] = b[14] & g[29007];
assign g[45392] = a[14] & g[29008];
assign g[61775] = b[14] & g[29008];
assign g[45393] = a[14] & g[29009];
assign g[61776] = b[14] & g[29009];
assign g[45394] = a[14] & g[29010];
assign g[61777] = b[14] & g[29010];
assign g[45395] = a[14] & g[29011];
assign g[61778] = b[14] & g[29011];
assign g[45396] = a[14] & g[29012];
assign g[61779] = b[14] & g[29012];
assign g[45397] = a[14] & g[29013];
assign g[61780] = b[14] & g[29013];
assign g[45398] = a[14] & g[29014];
assign g[61781] = b[14] & g[29014];
assign g[45399] = a[14] & g[29015];
assign g[61782] = b[14] & g[29015];
assign g[45400] = a[14] & g[29016];
assign g[61783] = b[14] & g[29016];
assign g[45401] = a[14] & g[29017];
assign g[61784] = b[14] & g[29017];
assign g[45402] = a[14] & g[29018];
assign g[61785] = b[14] & g[29018];
assign g[45403] = a[14] & g[29019];
assign g[61786] = b[14] & g[29019];
assign g[45404] = a[14] & g[29020];
assign g[61787] = b[14] & g[29020];
assign g[45405] = a[14] & g[29021];
assign g[61788] = b[14] & g[29021];
assign g[45406] = a[14] & g[29022];
assign g[61789] = b[14] & g[29022];
assign g[45407] = a[14] & g[29023];
assign g[61790] = b[14] & g[29023];
assign g[45408] = a[14] & g[29024];
assign g[61791] = b[14] & g[29024];
assign g[45409] = a[14] & g[29025];
assign g[61792] = b[14] & g[29025];
assign g[45410] = a[14] & g[29026];
assign g[61793] = b[14] & g[29026];
assign g[45411] = a[14] & g[29027];
assign g[61794] = b[14] & g[29027];
assign g[45412] = a[14] & g[29028];
assign g[61795] = b[14] & g[29028];
assign g[45413] = a[14] & g[29029];
assign g[61796] = b[14] & g[29029];
assign g[45414] = a[14] & g[29030];
assign g[61797] = b[14] & g[29030];
assign g[45415] = a[14] & g[29031];
assign g[61798] = b[14] & g[29031];
assign g[45416] = a[14] & g[29032];
assign g[61799] = b[14] & g[29032];
assign g[45417] = a[14] & g[29033];
assign g[61800] = b[14] & g[29033];
assign g[45418] = a[14] & g[29034];
assign g[61801] = b[14] & g[29034];
assign g[45419] = a[14] & g[29035];
assign g[61802] = b[14] & g[29035];
assign g[45420] = a[14] & g[29036];
assign g[61803] = b[14] & g[29036];
assign g[45421] = a[14] & g[29037];
assign g[61804] = b[14] & g[29037];
assign g[45422] = a[14] & g[29038];
assign g[61805] = b[14] & g[29038];
assign g[45423] = a[14] & g[29039];
assign g[61806] = b[14] & g[29039];
assign g[45424] = a[14] & g[29040];
assign g[61807] = b[14] & g[29040];
assign g[45425] = a[14] & g[29041];
assign g[61808] = b[14] & g[29041];
assign g[45426] = a[14] & g[29042];
assign g[61809] = b[14] & g[29042];
assign g[45427] = a[14] & g[29043];
assign g[61810] = b[14] & g[29043];
assign g[45428] = a[14] & g[29044];
assign g[61811] = b[14] & g[29044];
assign g[45429] = a[14] & g[29045];
assign g[61812] = b[14] & g[29045];
assign g[45430] = a[14] & g[29046];
assign g[61813] = b[14] & g[29046];
assign g[45431] = a[14] & g[29047];
assign g[61814] = b[14] & g[29047];
assign g[45432] = a[14] & g[29048];
assign g[61815] = b[14] & g[29048];
assign g[45433] = a[14] & g[29049];
assign g[61816] = b[14] & g[29049];
assign g[45434] = a[14] & g[29050];
assign g[61817] = b[14] & g[29050];
assign g[45435] = a[14] & g[29051];
assign g[61818] = b[14] & g[29051];
assign g[45436] = a[14] & g[29052];
assign g[61819] = b[14] & g[29052];
assign g[45437] = a[14] & g[29053];
assign g[61820] = b[14] & g[29053];
assign g[45438] = a[14] & g[29054];
assign g[61821] = b[14] & g[29054];
assign g[45439] = a[14] & g[29055];
assign g[61822] = b[14] & g[29055];
assign g[45440] = a[14] & g[29056];
assign g[61823] = b[14] & g[29056];
assign g[45441] = a[14] & g[29057];
assign g[61824] = b[14] & g[29057];
assign g[45442] = a[14] & g[29058];
assign g[61825] = b[14] & g[29058];
assign g[45443] = a[14] & g[29059];
assign g[61826] = b[14] & g[29059];
assign g[45444] = a[14] & g[29060];
assign g[61827] = b[14] & g[29060];
assign g[45445] = a[14] & g[29061];
assign g[61828] = b[14] & g[29061];
assign g[45446] = a[14] & g[29062];
assign g[61829] = b[14] & g[29062];
assign g[45447] = a[14] & g[29063];
assign g[61830] = b[14] & g[29063];
assign g[45448] = a[14] & g[29064];
assign g[61831] = b[14] & g[29064];
assign g[45449] = a[14] & g[29065];
assign g[61832] = b[14] & g[29065];
assign g[45450] = a[14] & g[29066];
assign g[61833] = b[14] & g[29066];
assign g[45451] = a[14] & g[29067];
assign g[61834] = b[14] & g[29067];
assign g[45452] = a[14] & g[29068];
assign g[61835] = b[14] & g[29068];
assign g[45453] = a[14] & g[29069];
assign g[61836] = b[14] & g[29069];
assign g[45454] = a[14] & g[29070];
assign g[61837] = b[14] & g[29070];
assign g[45455] = a[14] & g[29071];
assign g[61838] = b[14] & g[29071];
assign g[45456] = a[14] & g[29072];
assign g[61839] = b[14] & g[29072];
assign g[45457] = a[14] & g[29073];
assign g[61840] = b[14] & g[29073];
assign g[45458] = a[14] & g[29074];
assign g[61841] = b[14] & g[29074];
assign g[45459] = a[14] & g[29075];
assign g[61842] = b[14] & g[29075];
assign g[45460] = a[14] & g[29076];
assign g[61843] = b[14] & g[29076];
assign g[45461] = a[14] & g[29077];
assign g[61844] = b[14] & g[29077];
assign g[45462] = a[14] & g[29078];
assign g[61845] = b[14] & g[29078];
assign g[45463] = a[14] & g[29079];
assign g[61846] = b[14] & g[29079];
assign g[45464] = a[14] & g[29080];
assign g[61847] = b[14] & g[29080];
assign g[45465] = a[14] & g[29081];
assign g[61848] = b[14] & g[29081];
assign g[45466] = a[14] & g[29082];
assign g[61849] = b[14] & g[29082];
assign g[45467] = a[14] & g[29083];
assign g[61850] = b[14] & g[29083];
assign g[45468] = a[14] & g[29084];
assign g[61851] = b[14] & g[29084];
assign g[45469] = a[14] & g[29085];
assign g[61852] = b[14] & g[29085];
assign g[45470] = a[14] & g[29086];
assign g[61853] = b[14] & g[29086];
assign g[45471] = a[14] & g[29087];
assign g[61854] = b[14] & g[29087];
assign g[45472] = a[14] & g[29088];
assign g[61855] = b[14] & g[29088];
assign g[45473] = a[14] & g[29089];
assign g[61856] = b[14] & g[29089];
assign g[45474] = a[14] & g[29090];
assign g[61857] = b[14] & g[29090];
assign g[45475] = a[14] & g[29091];
assign g[61858] = b[14] & g[29091];
assign g[45476] = a[14] & g[29092];
assign g[61859] = b[14] & g[29092];
assign g[45477] = a[14] & g[29093];
assign g[61860] = b[14] & g[29093];
assign g[45478] = a[14] & g[29094];
assign g[61861] = b[14] & g[29094];
assign g[45479] = a[14] & g[29095];
assign g[61862] = b[14] & g[29095];
assign g[45480] = a[14] & g[29096];
assign g[61863] = b[14] & g[29096];
assign g[45481] = a[14] & g[29097];
assign g[61864] = b[14] & g[29097];
assign g[45482] = a[14] & g[29098];
assign g[61865] = b[14] & g[29098];
assign g[45483] = a[14] & g[29099];
assign g[61866] = b[14] & g[29099];
assign g[45484] = a[14] & g[29100];
assign g[61867] = b[14] & g[29100];
assign g[45485] = a[14] & g[29101];
assign g[61868] = b[14] & g[29101];
assign g[45486] = a[14] & g[29102];
assign g[61869] = b[14] & g[29102];
assign g[45487] = a[14] & g[29103];
assign g[61870] = b[14] & g[29103];
assign g[45488] = a[14] & g[29104];
assign g[61871] = b[14] & g[29104];
assign g[45489] = a[14] & g[29105];
assign g[61872] = b[14] & g[29105];
assign g[45490] = a[14] & g[29106];
assign g[61873] = b[14] & g[29106];
assign g[45491] = a[14] & g[29107];
assign g[61874] = b[14] & g[29107];
assign g[45492] = a[14] & g[29108];
assign g[61875] = b[14] & g[29108];
assign g[45493] = a[14] & g[29109];
assign g[61876] = b[14] & g[29109];
assign g[45494] = a[14] & g[29110];
assign g[61877] = b[14] & g[29110];
assign g[45495] = a[14] & g[29111];
assign g[61878] = b[14] & g[29111];
assign g[45496] = a[14] & g[29112];
assign g[61879] = b[14] & g[29112];
assign g[45497] = a[14] & g[29113];
assign g[61880] = b[14] & g[29113];
assign g[45498] = a[14] & g[29114];
assign g[61881] = b[14] & g[29114];
assign g[45499] = a[14] & g[29115];
assign g[61882] = b[14] & g[29115];
assign g[45500] = a[14] & g[29116];
assign g[61883] = b[14] & g[29116];
assign g[45501] = a[14] & g[29117];
assign g[61884] = b[14] & g[29117];
assign g[45502] = a[14] & g[29118];
assign g[61885] = b[14] & g[29118];
assign g[45503] = a[14] & g[29119];
assign g[61886] = b[14] & g[29119];
assign g[45504] = a[14] & g[29120];
assign g[61887] = b[14] & g[29120];
assign g[45505] = a[14] & g[29121];
assign g[61888] = b[14] & g[29121];
assign g[45506] = a[14] & g[29122];
assign g[61889] = b[14] & g[29122];
assign g[45507] = a[14] & g[29123];
assign g[61890] = b[14] & g[29123];
assign g[45508] = a[14] & g[29124];
assign g[61891] = b[14] & g[29124];
assign g[45509] = a[14] & g[29125];
assign g[61892] = b[14] & g[29125];
assign g[45510] = a[14] & g[29126];
assign g[61893] = b[14] & g[29126];
assign g[45511] = a[14] & g[29127];
assign g[61894] = b[14] & g[29127];
assign g[45512] = a[14] & g[29128];
assign g[61895] = b[14] & g[29128];
assign g[45513] = a[14] & g[29129];
assign g[61896] = b[14] & g[29129];
assign g[45514] = a[14] & g[29130];
assign g[61897] = b[14] & g[29130];
assign g[45515] = a[14] & g[29131];
assign g[61898] = b[14] & g[29131];
assign g[45516] = a[14] & g[29132];
assign g[61899] = b[14] & g[29132];
assign g[45517] = a[14] & g[29133];
assign g[61900] = b[14] & g[29133];
assign g[45518] = a[14] & g[29134];
assign g[61901] = b[14] & g[29134];
assign g[45519] = a[14] & g[29135];
assign g[61902] = b[14] & g[29135];
assign g[45520] = a[14] & g[29136];
assign g[61903] = b[14] & g[29136];
assign g[45521] = a[14] & g[29137];
assign g[61904] = b[14] & g[29137];
assign g[45522] = a[14] & g[29138];
assign g[61905] = b[14] & g[29138];
assign g[45523] = a[14] & g[29139];
assign g[61906] = b[14] & g[29139];
assign g[45524] = a[14] & g[29140];
assign g[61907] = b[14] & g[29140];
assign g[45525] = a[14] & g[29141];
assign g[61908] = b[14] & g[29141];
assign g[45526] = a[14] & g[29142];
assign g[61909] = b[14] & g[29142];
assign g[45527] = a[14] & g[29143];
assign g[61910] = b[14] & g[29143];
assign g[45528] = a[14] & g[29144];
assign g[61911] = b[14] & g[29144];
assign g[45529] = a[14] & g[29145];
assign g[61912] = b[14] & g[29145];
assign g[45530] = a[14] & g[29146];
assign g[61913] = b[14] & g[29146];
assign g[45531] = a[14] & g[29147];
assign g[61914] = b[14] & g[29147];
assign g[45532] = a[14] & g[29148];
assign g[61915] = b[14] & g[29148];
assign g[45533] = a[14] & g[29149];
assign g[61916] = b[14] & g[29149];
assign g[45534] = a[14] & g[29150];
assign g[61917] = b[14] & g[29150];
assign g[45535] = a[14] & g[29151];
assign g[61918] = b[14] & g[29151];
assign g[45536] = a[14] & g[29152];
assign g[61919] = b[14] & g[29152];
assign g[45537] = a[14] & g[29153];
assign g[61920] = b[14] & g[29153];
assign g[45538] = a[14] & g[29154];
assign g[61921] = b[14] & g[29154];
assign g[45539] = a[14] & g[29155];
assign g[61922] = b[14] & g[29155];
assign g[45540] = a[14] & g[29156];
assign g[61923] = b[14] & g[29156];
assign g[45541] = a[14] & g[29157];
assign g[61924] = b[14] & g[29157];
assign g[45542] = a[14] & g[29158];
assign g[61925] = b[14] & g[29158];
assign g[45543] = a[14] & g[29159];
assign g[61926] = b[14] & g[29159];
assign g[45544] = a[14] & g[29160];
assign g[61927] = b[14] & g[29160];
assign g[45545] = a[14] & g[29161];
assign g[61928] = b[14] & g[29161];
assign g[45546] = a[14] & g[29162];
assign g[61929] = b[14] & g[29162];
assign g[45547] = a[14] & g[29163];
assign g[61930] = b[14] & g[29163];
assign g[45548] = a[14] & g[29164];
assign g[61931] = b[14] & g[29164];
assign g[45549] = a[14] & g[29165];
assign g[61932] = b[14] & g[29165];
assign g[45550] = a[14] & g[29166];
assign g[61933] = b[14] & g[29166];
assign g[45551] = a[14] & g[29167];
assign g[61934] = b[14] & g[29167];
assign g[45552] = a[14] & g[29168];
assign g[61935] = b[14] & g[29168];
assign g[45553] = a[14] & g[29169];
assign g[61936] = b[14] & g[29169];
assign g[45554] = a[14] & g[29170];
assign g[61937] = b[14] & g[29170];
assign g[45555] = a[14] & g[29171];
assign g[61938] = b[14] & g[29171];
assign g[45556] = a[14] & g[29172];
assign g[61939] = b[14] & g[29172];
assign g[45557] = a[14] & g[29173];
assign g[61940] = b[14] & g[29173];
assign g[45558] = a[14] & g[29174];
assign g[61941] = b[14] & g[29174];
assign g[45559] = a[14] & g[29175];
assign g[61942] = b[14] & g[29175];
assign g[45560] = a[14] & g[29176];
assign g[61943] = b[14] & g[29176];
assign g[45561] = a[14] & g[29177];
assign g[61944] = b[14] & g[29177];
assign g[45562] = a[14] & g[29178];
assign g[61945] = b[14] & g[29178];
assign g[45563] = a[14] & g[29179];
assign g[61946] = b[14] & g[29179];
assign g[45564] = a[14] & g[29180];
assign g[61947] = b[14] & g[29180];
assign g[45565] = a[14] & g[29181];
assign g[61948] = b[14] & g[29181];
assign g[45566] = a[14] & g[29182];
assign g[61949] = b[14] & g[29182];
assign g[45567] = a[14] & g[29183];
assign g[61950] = b[14] & g[29183];
assign g[45568] = a[14] & g[29184];
assign g[61951] = b[14] & g[29184];
assign g[45569] = a[14] & g[29185];
assign g[61952] = b[14] & g[29185];
assign g[45570] = a[14] & g[29186];
assign g[61953] = b[14] & g[29186];
assign g[45571] = a[14] & g[29187];
assign g[61954] = b[14] & g[29187];
assign g[45572] = a[14] & g[29188];
assign g[61955] = b[14] & g[29188];
assign g[45573] = a[14] & g[29189];
assign g[61956] = b[14] & g[29189];
assign g[45574] = a[14] & g[29190];
assign g[61957] = b[14] & g[29190];
assign g[45575] = a[14] & g[29191];
assign g[61958] = b[14] & g[29191];
assign g[45576] = a[14] & g[29192];
assign g[61959] = b[14] & g[29192];
assign g[45577] = a[14] & g[29193];
assign g[61960] = b[14] & g[29193];
assign g[45578] = a[14] & g[29194];
assign g[61961] = b[14] & g[29194];
assign g[45579] = a[14] & g[29195];
assign g[61962] = b[14] & g[29195];
assign g[45580] = a[14] & g[29196];
assign g[61963] = b[14] & g[29196];
assign g[45581] = a[14] & g[29197];
assign g[61964] = b[14] & g[29197];
assign g[45582] = a[14] & g[29198];
assign g[61965] = b[14] & g[29198];
assign g[45583] = a[14] & g[29199];
assign g[61966] = b[14] & g[29199];
assign g[45584] = a[14] & g[29200];
assign g[61967] = b[14] & g[29200];
assign g[45585] = a[14] & g[29201];
assign g[61968] = b[14] & g[29201];
assign g[45586] = a[14] & g[29202];
assign g[61969] = b[14] & g[29202];
assign g[45587] = a[14] & g[29203];
assign g[61970] = b[14] & g[29203];
assign g[45588] = a[14] & g[29204];
assign g[61971] = b[14] & g[29204];
assign g[45589] = a[14] & g[29205];
assign g[61972] = b[14] & g[29205];
assign g[45590] = a[14] & g[29206];
assign g[61973] = b[14] & g[29206];
assign g[45591] = a[14] & g[29207];
assign g[61974] = b[14] & g[29207];
assign g[45592] = a[14] & g[29208];
assign g[61975] = b[14] & g[29208];
assign g[45593] = a[14] & g[29209];
assign g[61976] = b[14] & g[29209];
assign g[45594] = a[14] & g[29210];
assign g[61977] = b[14] & g[29210];
assign g[45595] = a[14] & g[29211];
assign g[61978] = b[14] & g[29211];
assign g[45596] = a[14] & g[29212];
assign g[61979] = b[14] & g[29212];
assign g[45597] = a[14] & g[29213];
assign g[61980] = b[14] & g[29213];
assign g[45598] = a[14] & g[29214];
assign g[61981] = b[14] & g[29214];
assign g[45599] = a[14] & g[29215];
assign g[61982] = b[14] & g[29215];
assign g[45600] = a[14] & g[29216];
assign g[61983] = b[14] & g[29216];
assign g[45601] = a[14] & g[29217];
assign g[61984] = b[14] & g[29217];
assign g[45602] = a[14] & g[29218];
assign g[61985] = b[14] & g[29218];
assign g[45603] = a[14] & g[29219];
assign g[61986] = b[14] & g[29219];
assign g[45604] = a[14] & g[29220];
assign g[61987] = b[14] & g[29220];
assign g[45605] = a[14] & g[29221];
assign g[61988] = b[14] & g[29221];
assign g[45606] = a[14] & g[29222];
assign g[61989] = b[14] & g[29222];
assign g[45607] = a[14] & g[29223];
assign g[61990] = b[14] & g[29223];
assign g[45608] = a[14] & g[29224];
assign g[61991] = b[14] & g[29224];
assign g[45609] = a[14] & g[29225];
assign g[61992] = b[14] & g[29225];
assign g[45610] = a[14] & g[29226];
assign g[61993] = b[14] & g[29226];
assign g[45611] = a[14] & g[29227];
assign g[61994] = b[14] & g[29227];
assign g[45612] = a[14] & g[29228];
assign g[61995] = b[14] & g[29228];
assign g[45613] = a[14] & g[29229];
assign g[61996] = b[14] & g[29229];
assign g[45614] = a[14] & g[29230];
assign g[61997] = b[14] & g[29230];
assign g[45615] = a[14] & g[29231];
assign g[61998] = b[14] & g[29231];
assign g[45616] = a[14] & g[29232];
assign g[61999] = b[14] & g[29232];
assign g[45617] = a[14] & g[29233];
assign g[62000] = b[14] & g[29233];
assign g[45618] = a[14] & g[29234];
assign g[62001] = b[14] & g[29234];
assign g[45619] = a[14] & g[29235];
assign g[62002] = b[14] & g[29235];
assign g[45620] = a[14] & g[29236];
assign g[62003] = b[14] & g[29236];
assign g[45621] = a[14] & g[29237];
assign g[62004] = b[14] & g[29237];
assign g[45622] = a[14] & g[29238];
assign g[62005] = b[14] & g[29238];
assign g[45623] = a[14] & g[29239];
assign g[62006] = b[14] & g[29239];
assign g[45624] = a[14] & g[29240];
assign g[62007] = b[14] & g[29240];
assign g[45625] = a[14] & g[29241];
assign g[62008] = b[14] & g[29241];
assign g[45626] = a[14] & g[29242];
assign g[62009] = b[14] & g[29242];
assign g[45627] = a[14] & g[29243];
assign g[62010] = b[14] & g[29243];
assign g[45628] = a[14] & g[29244];
assign g[62011] = b[14] & g[29244];
assign g[45629] = a[14] & g[29245];
assign g[62012] = b[14] & g[29245];
assign g[45630] = a[14] & g[29246];
assign g[62013] = b[14] & g[29246];
assign g[45631] = a[14] & g[29247];
assign g[62014] = b[14] & g[29247];
assign g[45632] = a[14] & g[29248];
assign g[62015] = b[14] & g[29248];
assign g[45633] = a[14] & g[29249];
assign g[62016] = b[14] & g[29249];
assign g[45634] = a[14] & g[29250];
assign g[62017] = b[14] & g[29250];
assign g[45635] = a[14] & g[29251];
assign g[62018] = b[14] & g[29251];
assign g[45636] = a[14] & g[29252];
assign g[62019] = b[14] & g[29252];
assign g[45637] = a[14] & g[29253];
assign g[62020] = b[14] & g[29253];
assign g[45638] = a[14] & g[29254];
assign g[62021] = b[14] & g[29254];
assign g[45639] = a[14] & g[29255];
assign g[62022] = b[14] & g[29255];
assign g[45640] = a[14] & g[29256];
assign g[62023] = b[14] & g[29256];
assign g[45641] = a[14] & g[29257];
assign g[62024] = b[14] & g[29257];
assign g[45642] = a[14] & g[29258];
assign g[62025] = b[14] & g[29258];
assign g[45643] = a[14] & g[29259];
assign g[62026] = b[14] & g[29259];
assign g[45644] = a[14] & g[29260];
assign g[62027] = b[14] & g[29260];
assign g[45645] = a[14] & g[29261];
assign g[62028] = b[14] & g[29261];
assign g[45646] = a[14] & g[29262];
assign g[62029] = b[14] & g[29262];
assign g[45647] = a[14] & g[29263];
assign g[62030] = b[14] & g[29263];
assign g[45648] = a[14] & g[29264];
assign g[62031] = b[14] & g[29264];
assign g[45649] = a[14] & g[29265];
assign g[62032] = b[14] & g[29265];
assign g[45650] = a[14] & g[29266];
assign g[62033] = b[14] & g[29266];
assign g[45651] = a[14] & g[29267];
assign g[62034] = b[14] & g[29267];
assign g[45652] = a[14] & g[29268];
assign g[62035] = b[14] & g[29268];
assign g[45653] = a[14] & g[29269];
assign g[62036] = b[14] & g[29269];
assign g[45654] = a[14] & g[29270];
assign g[62037] = b[14] & g[29270];
assign g[45655] = a[14] & g[29271];
assign g[62038] = b[14] & g[29271];
assign g[45656] = a[14] & g[29272];
assign g[62039] = b[14] & g[29272];
assign g[45657] = a[14] & g[29273];
assign g[62040] = b[14] & g[29273];
assign g[45658] = a[14] & g[29274];
assign g[62041] = b[14] & g[29274];
assign g[45659] = a[14] & g[29275];
assign g[62042] = b[14] & g[29275];
assign g[45660] = a[14] & g[29276];
assign g[62043] = b[14] & g[29276];
assign g[45661] = a[14] & g[29277];
assign g[62044] = b[14] & g[29277];
assign g[45662] = a[14] & g[29278];
assign g[62045] = b[14] & g[29278];
assign g[45663] = a[14] & g[29279];
assign g[62046] = b[14] & g[29279];
assign g[45664] = a[14] & g[29280];
assign g[62047] = b[14] & g[29280];
assign g[45665] = a[14] & g[29281];
assign g[62048] = b[14] & g[29281];
assign g[45666] = a[14] & g[29282];
assign g[62049] = b[14] & g[29282];
assign g[45667] = a[14] & g[29283];
assign g[62050] = b[14] & g[29283];
assign g[45668] = a[14] & g[29284];
assign g[62051] = b[14] & g[29284];
assign g[45669] = a[14] & g[29285];
assign g[62052] = b[14] & g[29285];
assign g[45670] = a[14] & g[29286];
assign g[62053] = b[14] & g[29286];
assign g[45671] = a[14] & g[29287];
assign g[62054] = b[14] & g[29287];
assign g[45672] = a[14] & g[29288];
assign g[62055] = b[14] & g[29288];
assign g[45673] = a[14] & g[29289];
assign g[62056] = b[14] & g[29289];
assign g[45674] = a[14] & g[29290];
assign g[62057] = b[14] & g[29290];
assign g[45675] = a[14] & g[29291];
assign g[62058] = b[14] & g[29291];
assign g[45676] = a[14] & g[29292];
assign g[62059] = b[14] & g[29292];
assign g[45677] = a[14] & g[29293];
assign g[62060] = b[14] & g[29293];
assign g[45678] = a[14] & g[29294];
assign g[62061] = b[14] & g[29294];
assign g[45679] = a[14] & g[29295];
assign g[62062] = b[14] & g[29295];
assign g[45680] = a[14] & g[29296];
assign g[62063] = b[14] & g[29296];
assign g[45681] = a[14] & g[29297];
assign g[62064] = b[14] & g[29297];
assign g[45682] = a[14] & g[29298];
assign g[62065] = b[14] & g[29298];
assign g[45683] = a[14] & g[29299];
assign g[62066] = b[14] & g[29299];
assign g[45684] = a[14] & g[29300];
assign g[62067] = b[14] & g[29300];
assign g[45685] = a[14] & g[29301];
assign g[62068] = b[14] & g[29301];
assign g[45686] = a[14] & g[29302];
assign g[62069] = b[14] & g[29302];
assign g[45687] = a[14] & g[29303];
assign g[62070] = b[14] & g[29303];
assign g[45688] = a[14] & g[29304];
assign g[62071] = b[14] & g[29304];
assign g[45689] = a[14] & g[29305];
assign g[62072] = b[14] & g[29305];
assign g[45690] = a[14] & g[29306];
assign g[62073] = b[14] & g[29306];
assign g[45691] = a[14] & g[29307];
assign g[62074] = b[14] & g[29307];
assign g[45692] = a[14] & g[29308];
assign g[62075] = b[14] & g[29308];
assign g[45693] = a[14] & g[29309];
assign g[62076] = b[14] & g[29309];
assign g[45694] = a[14] & g[29310];
assign g[62077] = b[14] & g[29310];
assign g[45695] = a[14] & g[29311];
assign g[62078] = b[14] & g[29311];
assign g[45696] = a[14] & g[29312];
assign g[62079] = b[14] & g[29312];
assign g[45697] = a[14] & g[29313];
assign g[62080] = b[14] & g[29313];
assign g[45698] = a[14] & g[29314];
assign g[62081] = b[14] & g[29314];
assign g[45699] = a[14] & g[29315];
assign g[62082] = b[14] & g[29315];
assign g[45700] = a[14] & g[29316];
assign g[62083] = b[14] & g[29316];
assign g[45701] = a[14] & g[29317];
assign g[62084] = b[14] & g[29317];
assign g[45702] = a[14] & g[29318];
assign g[62085] = b[14] & g[29318];
assign g[45703] = a[14] & g[29319];
assign g[62086] = b[14] & g[29319];
assign g[45704] = a[14] & g[29320];
assign g[62087] = b[14] & g[29320];
assign g[45705] = a[14] & g[29321];
assign g[62088] = b[14] & g[29321];
assign g[45706] = a[14] & g[29322];
assign g[62089] = b[14] & g[29322];
assign g[45707] = a[14] & g[29323];
assign g[62090] = b[14] & g[29323];
assign g[45708] = a[14] & g[29324];
assign g[62091] = b[14] & g[29324];
assign g[45709] = a[14] & g[29325];
assign g[62092] = b[14] & g[29325];
assign g[45710] = a[14] & g[29326];
assign g[62093] = b[14] & g[29326];
assign g[45711] = a[14] & g[29327];
assign g[62094] = b[14] & g[29327];
assign g[45712] = a[14] & g[29328];
assign g[62095] = b[14] & g[29328];
assign g[45713] = a[14] & g[29329];
assign g[62096] = b[14] & g[29329];
assign g[45714] = a[14] & g[29330];
assign g[62097] = b[14] & g[29330];
assign g[45715] = a[14] & g[29331];
assign g[62098] = b[14] & g[29331];
assign g[45716] = a[14] & g[29332];
assign g[62099] = b[14] & g[29332];
assign g[45717] = a[14] & g[29333];
assign g[62100] = b[14] & g[29333];
assign g[45718] = a[14] & g[29334];
assign g[62101] = b[14] & g[29334];
assign g[45719] = a[14] & g[29335];
assign g[62102] = b[14] & g[29335];
assign g[45720] = a[14] & g[29336];
assign g[62103] = b[14] & g[29336];
assign g[45721] = a[14] & g[29337];
assign g[62104] = b[14] & g[29337];
assign g[45722] = a[14] & g[29338];
assign g[62105] = b[14] & g[29338];
assign g[45723] = a[14] & g[29339];
assign g[62106] = b[14] & g[29339];
assign g[45724] = a[14] & g[29340];
assign g[62107] = b[14] & g[29340];
assign g[45725] = a[14] & g[29341];
assign g[62108] = b[14] & g[29341];
assign g[45726] = a[14] & g[29342];
assign g[62109] = b[14] & g[29342];
assign g[45727] = a[14] & g[29343];
assign g[62110] = b[14] & g[29343];
assign g[45728] = a[14] & g[29344];
assign g[62111] = b[14] & g[29344];
assign g[45729] = a[14] & g[29345];
assign g[62112] = b[14] & g[29345];
assign g[45730] = a[14] & g[29346];
assign g[62113] = b[14] & g[29346];
assign g[45731] = a[14] & g[29347];
assign g[62114] = b[14] & g[29347];
assign g[45732] = a[14] & g[29348];
assign g[62115] = b[14] & g[29348];
assign g[45733] = a[14] & g[29349];
assign g[62116] = b[14] & g[29349];
assign g[45734] = a[14] & g[29350];
assign g[62117] = b[14] & g[29350];
assign g[45735] = a[14] & g[29351];
assign g[62118] = b[14] & g[29351];
assign g[45736] = a[14] & g[29352];
assign g[62119] = b[14] & g[29352];
assign g[45737] = a[14] & g[29353];
assign g[62120] = b[14] & g[29353];
assign g[45738] = a[14] & g[29354];
assign g[62121] = b[14] & g[29354];
assign g[45739] = a[14] & g[29355];
assign g[62122] = b[14] & g[29355];
assign g[45740] = a[14] & g[29356];
assign g[62123] = b[14] & g[29356];
assign g[45741] = a[14] & g[29357];
assign g[62124] = b[14] & g[29357];
assign g[45742] = a[14] & g[29358];
assign g[62125] = b[14] & g[29358];
assign g[45743] = a[14] & g[29359];
assign g[62126] = b[14] & g[29359];
assign g[45744] = a[14] & g[29360];
assign g[62127] = b[14] & g[29360];
assign g[45745] = a[14] & g[29361];
assign g[62128] = b[14] & g[29361];
assign g[45746] = a[14] & g[29362];
assign g[62129] = b[14] & g[29362];
assign g[45747] = a[14] & g[29363];
assign g[62130] = b[14] & g[29363];
assign g[45748] = a[14] & g[29364];
assign g[62131] = b[14] & g[29364];
assign g[45749] = a[14] & g[29365];
assign g[62132] = b[14] & g[29365];
assign g[45750] = a[14] & g[29366];
assign g[62133] = b[14] & g[29366];
assign g[45751] = a[14] & g[29367];
assign g[62134] = b[14] & g[29367];
assign g[45752] = a[14] & g[29368];
assign g[62135] = b[14] & g[29368];
assign g[45753] = a[14] & g[29369];
assign g[62136] = b[14] & g[29369];
assign g[45754] = a[14] & g[29370];
assign g[62137] = b[14] & g[29370];
assign g[45755] = a[14] & g[29371];
assign g[62138] = b[14] & g[29371];
assign g[45756] = a[14] & g[29372];
assign g[62139] = b[14] & g[29372];
assign g[45757] = a[14] & g[29373];
assign g[62140] = b[14] & g[29373];
assign g[45758] = a[14] & g[29374];
assign g[62141] = b[14] & g[29374];
assign g[45759] = a[14] & g[29375];
assign g[62142] = b[14] & g[29375];
assign g[45760] = a[14] & g[29376];
assign g[62143] = b[14] & g[29376];
assign g[45761] = a[14] & g[29377];
assign g[62144] = b[14] & g[29377];
assign g[45762] = a[14] & g[29378];
assign g[62145] = b[14] & g[29378];
assign g[45763] = a[14] & g[29379];
assign g[62146] = b[14] & g[29379];
assign g[45764] = a[14] & g[29380];
assign g[62147] = b[14] & g[29380];
assign g[45765] = a[14] & g[29381];
assign g[62148] = b[14] & g[29381];
assign g[45766] = a[14] & g[29382];
assign g[62149] = b[14] & g[29382];
assign g[45767] = a[14] & g[29383];
assign g[62150] = b[14] & g[29383];
assign g[45768] = a[14] & g[29384];
assign g[62151] = b[14] & g[29384];
assign g[45769] = a[14] & g[29385];
assign g[62152] = b[14] & g[29385];
assign g[45770] = a[14] & g[29386];
assign g[62153] = b[14] & g[29386];
assign g[45771] = a[14] & g[29387];
assign g[62154] = b[14] & g[29387];
assign g[45772] = a[14] & g[29388];
assign g[62155] = b[14] & g[29388];
assign g[45773] = a[14] & g[29389];
assign g[62156] = b[14] & g[29389];
assign g[45774] = a[14] & g[29390];
assign g[62157] = b[14] & g[29390];
assign g[45775] = a[14] & g[29391];
assign g[62158] = b[14] & g[29391];
assign g[45776] = a[14] & g[29392];
assign g[62159] = b[14] & g[29392];
assign g[45777] = a[14] & g[29393];
assign g[62160] = b[14] & g[29393];
assign g[45778] = a[14] & g[29394];
assign g[62161] = b[14] & g[29394];
assign g[45779] = a[14] & g[29395];
assign g[62162] = b[14] & g[29395];
assign g[45780] = a[14] & g[29396];
assign g[62163] = b[14] & g[29396];
assign g[45781] = a[14] & g[29397];
assign g[62164] = b[14] & g[29397];
assign g[45782] = a[14] & g[29398];
assign g[62165] = b[14] & g[29398];
assign g[45783] = a[14] & g[29399];
assign g[62166] = b[14] & g[29399];
assign g[45784] = a[14] & g[29400];
assign g[62167] = b[14] & g[29400];
assign g[45785] = a[14] & g[29401];
assign g[62168] = b[14] & g[29401];
assign g[45786] = a[14] & g[29402];
assign g[62169] = b[14] & g[29402];
assign g[45787] = a[14] & g[29403];
assign g[62170] = b[14] & g[29403];
assign g[45788] = a[14] & g[29404];
assign g[62171] = b[14] & g[29404];
assign g[45789] = a[14] & g[29405];
assign g[62172] = b[14] & g[29405];
assign g[45790] = a[14] & g[29406];
assign g[62173] = b[14] & g[29406];
assign g[45791] = a[14] & g[29407];
assign g[62174] = b[14] & g[29407];
assign g[45792] = a[14] & g[29408];
assign g[62175] = b[14] & g[29408];
assign g[45793] = a[14] & g[29409];
assign g[62176] = b[14] & g[29409];
assign g[45794] = a[14] & g[29410];
assign g[62177] = b[14] & g[29410];
assign g[45795] = a[14] & g[29411];
assign g[62178] = b[14] & g[29411];
assign g[45796] = a[14] & g[29412];
assign g[62179] = b[14] & g[29412];
assign g[45797] = a[14] & g[29413];
assign g[62180] = b[14] & g[29413];
assign g[45798] = a[14] & g[29414];
assign g[62181] = b[14] & g[29414];
assign g[45799] = a[14] & g[29415];
assign g[62182] = b[14] & g[29415];
assign g[45800] = a[14] & g[29416];
assign g[62183] = b[14] & g[29416];
assign g[45801] = a[14] & g[29417];
assign g[62184] = b[14] & g[29417];
assign g[45802] = a[14] & g[29418];
assign g[62185] = b[14] & g[29418];
assign g[45803] = a[14] & g[29419];
assign g[62186] = b[14] & g[29419];
assign g[45804] = a[14] & g[29420];
assign g[62187] = b[14] & g[29420];
assign g[45805] = a[14] & g[29421];
assign g[62188] = b[14] & g[29421];
assign g[45806] = a[14] & g[29422];
assign g[62189] = b[14] & g[29422];
assign g[45807] = a[14] & g[29423];
assign g[62190] = b[14] & g[29423];
assign g[45808] = a[14] & g[29424];
assign g[62191] = b[14] & g[29424];
assign g[45809] = a[14] & g[29425];
assign g[62192] = b[14] & g[29425];
assign g[45810] = a[14] & g[29426];
assign g[62193] = b[14] & g[29426];
assign g[45811] = a[14] & g[29427];
assign g[62194] = b[14] & g[29427];
assign g[45812] = a[14] & g[29428];
assign g[62195] = b[14] & g[29428];
assign g[45813] = a[14] & g[29429];
assign g[62196] = b[14] & g[29429];
assign g[45814] = a[14] & g[29430];
assign g[62197] = b[14] & g[29430];
assign g[45815] = a[14] & g[29431];
assign g[62198] = b[14] & g[29431];
assign g[45816] = a[14] & g[29432];
assign g[62199] = b[14] & g[29432];
assign g[45817] = a[14] & g[29433];
assign g[62200] = b[14] & g[29433];
assign g[45818] = a[14] & g[29434];
assign g[62201] = b[14] & g[29434];
assign g[45819] = a[14] & g[29435];
assign g[62202] = b[14] & g[29435];
assign g[45820] = a[14] & g[29436];
assign g[62203] = b[14] & g[29436];
assign g[45821] = a[14] & g[29437];
assign g[62204] = b[14] & g[29437];
assign g[45822] = a[14] & g[29438];
assign g[62205] = b[14] & g[29438];
assign g[45823] = a[14] & g[29439];
assign g[62206] = b[14] & g[29439];
assign g[45824] = a[14] & g[29440];
assign g[62207] = b[14] & g[29440];
assign g[45825] = a[14] & g[29441];
assign g[62208] = b[14] & g[29441];
assign g[45826] = a[14] & g[29442];
assign g[62209] = b[14] & g[29442];
assign g[45827] = a[14] & g[29443];
assign g[62210] = b[14] & g[29443];
assign g[45828] = a[14] & g[29444];
assign g[62211] = b[14] & g[29444];
assign g[45829] = a[14] & g[29445];
assign g[62212] = b[14] & g[29445];
assign g[45830] = a[14] & g[29446];
assign g[62213] = b[14] & g[29446];
assign g[45831] = a[14] & g[29447];
assign g[62214] = b[14] & g[29447];
assign g[45832] = a[14] & g[29448];
assign g[62215] = b[14] & g[29448];
assign g[45833] = a[14] & g[29449];
assign g[62216] = b[14] & g[29449];
assign g[45834] = a[14] & g[29450];
assign g[62217] = b[14] & g[29450];
assign g[45835] = a[14] & g[29451];
assign g[62218] = b[14] & g[29451];
assign g[45836] = a[14] & g[29452];
assign g[62219] = b[14] & g[29452];
assign g[45837] = a[14] & g[29453];
assign g[62220] = b[14] & g[29453];
assign g[45838] = a[14] & g[29454];
assign g[62221] = b[14] & g[29454];
assign g[45839] = a[14] & g[29455];
assign g[62222] = b[14] & g[29455];
assign g[45840] = a[14] & g[29456];
assign g[62223] = b[14] & g[29456];
assign g[45841] = a[14] & g[29457];
assign g[62224] = b[14] & g[29457];
assign g[45842] = a[14] & g[29458];
assign g[62225] = b[14] & g[29458];
assign g[45843] = a[14] & g[29459];
assign g[62226] = b[14] & g[29459];
assign g[45844] = a[14] & g[29460];
assign g[62227] = b[14] & g[29460];
assign g[45845] = a[14] & g[29461];
assign g[62228] = b[14] & g[29461];
assign g[45846] = a[14] & g[29462];
assign g[62229] = b[14] & g[29462];
assign g[45847] = a[14] & g[29463];
assign g[62230] = b[14] & g[29463];
assign g[45848] = a[14] & g[29464];
assign g[62231] = b[14] & g[29464];
assign g[45849] = a[14] & g[29465];
assign g[62232] = b[14] & g[29465];
assign g[45850] = a[14] & g[29466];
assign g[62233] = b[14] & g[29466];
assign g[45851] = a[14] & g[29467];
assign g[62234] = b[14] & g[29467];
assign g[45852] = a[14] & g[29468];
assign g[62235] = b[14] & g[29468];
assign g[45853] = a[14] & g[29469];
assign g[62236] = b[14] & g[29469];
assign g[45854] = a[14] & g[29470];
assign g[62237] = b[14] & g[29470];
assign g[45855] = a[14] & g[29471];
assign g[62238] = b[14] & g[29471];
assign g[45856] = a[14] & g[29472];
assign g[62239] = b[14] & g[29472];
assign g[45857] = a[14] & g[29473];
assign g[62240] = b[14] & g[29473];
assign g[45858] = a[14] & g[29474];
assign g[62241] = b[14] & g[29474];
assign g[45859] = a[14] & g[29475];
assign g[62242] = b[14] & g[29475];
assign g[45860] = a[14] & g[29476];
assign g[62243] = b[14] & g[29476];
assign g[45861] = a[14] & g[29477];
assign g[62244] = b[14] & g[29477];
assign g[45862] = a[14] & g[29478];
assign g[62245] = b[14] & g[29478];
assign g[45863] = a[14] & g[29479];
assign g[62246] = b[14] & g[29479];
assign g[45864] = a[14] & g[29480];
assign g[62247] = b[14] & g[29480];
assign g[45865] = a[14] & g[29481];
assign g[62248] = b[14] & g[29481];
assign g[45866] = a[14] & g[29482];
assign g[62249] = b[14] & g[29482];
assign g[45867] = a[14] & g[29483];
assign g[62250] = b[14] & g[29483];
assign g[45868] = a[14] & g[29484];
assign g[62251] = b[14] & g[29484];
assign g[45869] = a[14] & g[29485];
assign g[62252] = b[14] & g[29485];
assign g[45870] = a[14] & g[29486];
assign g[62253] = b[14] & g[29486];
assign g[45871] = a[14] & g[29487];
assign g[62254] = b[14] & g[29487];
assign g[45872] = a[14] & g[29488];
assign g[62255] = b[14] & g[29488];
assign g[45873] = a[14] & g[29489];
assign g[62256] = b[14] & g[29489];
assign g[45874] = a[14] & g[29490];
assign g[62257] = b[14] & g[29490];
assign g[45875] = a[14] & g[29491];
assign g[62258] = b[14] & g[29491];
assign g[45876] = a[14] & g[29492];
assign g[62259] = b[14] & g[29492];
assign g[45877] = a[14] & g[29493];
assign g[62260] = b[14] & g[29493];
assign g[45878] = a[14] & g[29494];
assign g[62261] = b[14] & g[29494];
assign g[45879] = a[14] & g[29495];
assign g[62262] = b[14] & g[29495];
assign g[45880] = a[14] & g[29496];
assign g[62263] = b[14] & g[29496];
assign g[45881] = a[14] & g[29497];
assign g[62264] = b[14] & g[29497];
assign g[45882] = a[14] & g[29498];
assign g[62265] = b[14] & g[29498];
assign g[45883] = a[14] & g[29499];
assign g[62266] = b[14] & g[29499];
assign g[45884] = a[14] & g[29500];
assign g[62267] = b[14] & g[29500];
assign g[45885] = a[14] & g[29501];
assign g[62268] = b[14] & g[29501];
assign g[45886] = a[14] & g[29502];
assign g[62269] = b[14] & g[29502];
assign g[45887] = a[14] & g[29503];
assign g[62270] = b[14] & g[29503];
assign g[45888] = a[14] & g[29504];
assign g[62271] = b[14] & g[29504];
assign g[45889] = a[14] & g[29505];
assign g[62272] = b[14] & g[29505];
assign g[45890] = a[14] & g[29506];
assign g[62273] = b[14] & g[29506];
assign g[45891] = a[14] & g[29507];
assign g[62274] = b[14] & g[29507];
assign g[45892] = a[14] & g[29508];
assign g[62275] = b[14] & g[29508];
assign g[45893] = a[14] & g[29509];
assign g[62276] = b[14] & g[29509];
assign g[45894] = a[14] & g[29510];
assign g[62277] = b[14] & g[29510];
assign g[45895] = a[14] & g[29511];
assign g[62278] = b[14] & g[29511];
assign g[45896] = a[14] & g[29512];
assign g[62279] = b[14] & g[29512];
assign g[45897] = a[14] & g[29513];
assign g[62280] = b[14] & g[29513];
assign g[45898] = a[14] & g[29514];
assign g[62281] = b[14] & g[29514];
assign g[45899] = a[14] & g[29515];
assign g[62282] = b[14] & g[29515];
assign g[45900] = a[14] & g[29516];
assign g[62283] = b[14] & g[29516];
assign g[45901] = a[14] & g[29517];
assign g[62284] = b[14] & g[29517];
assign g[45902] = a[14] & g[29518];
assign g[62285] = b[14] & g[29518];
assign g[45903] = a[14] & g[29519];
assign g[62286] = b[14] & g[29519];
assign g[45904] = a[14] & g[29520];
assign g[62287] = b[14] & g[29520];
assign g[45905] = a[14] & g[29521];
assign g[62288] = b[14] & g[29521];
assign g[45906] = a[14] & g[29522];
assign g[62289] = b[14] & g[29522];
assign g[45907] = a[14] & g[29523];
assign g[62290] = b[14] & g[29523];
assign g[45908] = a[14] & g[29524];
assign g[62291] = b[14] & g[29524];
assign g[45909] = a[14] & g[29525];
assign g[62292] = b[14] & g[29525];
assign g[45910] = a[14] & g[29526];
assign g[62293] = b[14] & g[29526];
assign g[45911] = a[14] & g[29527];
assign g[62294] = b[14] & g[29527];
assign g[45912] = a[14] & g[29528];
assign g[62295] = b[14] & g[29528];
assign g[45913] = a[14] & g[29529];
assign g[62296] = b[14] & g[29529];
assign g[45914] = a[14] & g[29530];
assign g[62297] = b[14] & g[29530];
assign g[45915] = a[14] & g[29531];
assign g[62298] = b[14] & g[29531];
assign g[45916] = a[14] & g[29532];
assign g[62299] = b[14] & g[29532];
assign g[45917] = a[14] & g[29533];
assign g[62300] = b[14] & g[29533];
assign g[45918] = a[14] & g[29534];
assign g[62301] = b[14] & g[29534];
assign g[45919] = a[14] & g[29535];
assign g[62302] = b[14] & g[29535];
assign g[45920] = a[14] & g[29536];
assign g[62303] = b[14] & g[29536];
assign g[45921] = a[14] & g[29537];
assign g[62304] = b[14] & g[29537];
assign g[45922] = a[14] & g[29538];
assign g[62305] = b[14] & g[29538];
assign g[45923] = a[14] & g[29539];
assign g[62306] = b[14] & g[29539];
assign g[45924] = a[14] & g[29540];
assign g[62307] = b[14] & g[29540];
assign g[45925] = a[14] & g[29541];
assign g[62308] = b[14] & g[29541];
assign g[45926] = a[14] & g[29542];
assign g[62309] = b[14] & g[29542];
assign g[45927] = a[14] & g[29543];
assign g[62310] = b[14] & g[29543];
assign g[45928] = a[14] & g[29544];
assign g[62311] = b[14] & g[29544];
assign g[45929] = a[14] & g[29545];
assign g[62312] = b[14] & g[29545];
assign g[45930] = a[14] & g[29546];
assign g[62313] = b[14] & g[29546];
assign g[45931] = a[14] & g[29547];
assign g[62314] = b[14] & g[29547];
assign g[45932] = a[14] & g[29548];
assign g[62315] = b[14] & g[29548];
assign g[45933] = a[14] & g[29549];
assign g[62316] = b[14] & g[29549];
assign g[45934] = a[14] & g[29550];
assign g[62317] = b[14] & g[29550];
assign g[45935] = a[14] & g[29551];
assign g[62318] = b[14] & g[29551];
assign g[45936] = a[14] & g[29552];
assign g[62319] = b[14] & g[29552];
assign g[45937] = a[14] & g[29553];
assign g[62320] = b[14] & g[29553];
assign g[45938] = a[14] & g[29554];
assign g[62321] = b[14] & g[29554];
assign g[45939] = a[14] & g[29555];
assign g[62322] = b[14] & g[29555];
assign g[45940] = a[14] & g[29556];
assign g[62323] = b[14] & g[29556];
assign g[45941] = a[14] & g[29557];
assign g[62324] = b[14] & g[29557];
assign g[45942] = a[14] & g[29558];
assign g[62325] = b[14] & g[29558];
assign g[45943] = a[14] & g[29559];
assign g[62326] = b[14] & g[29559];
assign g[45944] = a[14] & g[29560];
assign g[62327] = b[14] & g[29560];
assign g[45945] = a[14] & g[29561];
assign g[62328] = b[14] & g[29561];
assign g[45946] = a[14] & g[29562];
assign g[62329] = b[14] & g[29562];
assign g[45947] = a[14] & g[29563];
assign g[62330] = b[14] & g[29563];
assign g[45948] = a[14] & g[29564];
assign g[62331] = b[14] & g[29564];
assign g[45949] = a[14] & g[29565];
assign g[62332] = b[14] & g[29565];
assign g[45950] = a[14] & g[29566];
assign g[62333] = b[14] & g[29566];
assign g[45951] = a[14] & g[29567];
assign g[62334] = b[14] & g[29567];
assign g[45952] = a[14] & g[29568];
assign g[62335] = b[14] & g[29568];
assign g[45953] = a[14] & g[29569];
assign g[62336] = b[14] & g[29569];
assign g[45954] = a[14] & g[29570];
assign g[62337] = b[14] & g[29570];
assign g[45955] = a[14] & g[29571];
assign g[62338] = b[14] & g[29571];
assign g[45956] = a[14] & g[29572];
assign g[62339] = b[14] & g[29572];
assign g[45957] = a[14] & g[29573];
assign g[62340] = b[14] & g[29573];
assign g[45958] = a[14] & g[29574];
assign g[62341] = b[14] & g[29574];
assign g[45959] = a[14] & g[29575];
assign g[62342] = b[14] & g[29575];
assign g[45960] = a[14] & g[29576];
assign g[62343] = b[14] & g[29576];
assign g[45961] = a[14] & g[29577];
assign g[62344] = b[14] & g[29577];
assign g[45962] = a[14] & g[29578];
assign g[62345] = b[14] & g[29578];
assign g[45963] = a[14] & g[29579];
assign g[62346] = b[14] & g[29579];
assign g[45964] = a[14] & g[29580];
assign g[62347] = b[14] & g[29580];
assign g[45965] = a[14] & g[29581];
assign g[62348] = b[14] & g[29581];
assign g[45966] = a[14] & g[29582];
assign g[62349] = b[14] & g[29582];
assign g[45967] = a[14] & g[29583];
assign g[62350] = b[14] & g[29583];
assign g[45968] = a[14] & g[29584];
assign g[62351] = b[14] & g[29584];
assign g[45969] = a[14] & g[29585];
assign g[62352] = b[14] & g[29585];
assign g[45970] = a[14] & g[29586];
assign g[62353] = b[14] & g[29586];
assign g[45971] = a[14] & g[29587];
assign g[62354] = b[14] & g[29587];
assign g[45972] = a[14] & g[29588];
assign g[62355] = b[14] & g[29588];
assign g[45973] = a[14] & g[29589];
assign g[62356] = b[14] & g[29589];
assign g[45974] = a[14] & g[29590];
assign g[62357] = b[14] & g[29590];
assign g[45975] = a[14] & g[29591];
assign g[62358] = b[14] & g[29591];
assign g[45976] = a[14] & g[29592];
assign g[62359] = b[14] & g[29592];
assign g[45977] = a[14] & g[29593];
assign g[62360] = b[14] & g[29593];
assign g[45978] = a[14] & g[29594];
assign g[62361] = b[14] & g[29594];
assign g[45979] = a[14] & g[29595];
assign g[62362] = b[14] & g[29595];
assign g[45980] = a[14] & g[29596];
assign g[62363] = b[14] & g[29596];
assign g[45981] = a[14] & g[29597];
assign g[62364] = b[14] & g[29597];
assign g[45982] = a[14] & g[29598];
assign g[62365] = b[14] & g[29598];
assign g[45983] = a[14] & g[29599];
assign g[62366] = b[14] & g[29599];
assign g[45984] = a[14] & g[29600];
assign g[62367] = b[14] & g[29600];
assign g[45985] = a[14] & g[29601];
assign g[62368] = b[14] & g[29601];
assign g[45986] = a[14] & g[29602];
assign g[62369] = b[14] & g[29602];
assign g[45987] = a[14] & g[29603];
assign g[62370] = b[14] & g[29603];
assign g[45988] = a[14] & g[29604];
assign g[62371] = b[14] & g[29604];
assign g[45989] = a[14] & g[29605];
assign g[62372] = b[14] & g[29605];
assign g[45990] = a[14] & g[29606];
assign g[62373] = b[14] & g[29606];
assign g[45991] = a[14] & g[29607];
assign g[62374] = b[14] & g[29607];
assign g[45992] = a[14] & g[29608];
assign g[62375] = b[14] & g[29608];
assign g[45993] = a[14] & g[29609];
assign g[62376] = b[14] & g[29609];
assign g[45994] = a[14] & g[29610];
assign g[62377] = b[14] & g[29610];
assign g[45995] = a[14] & g[29611];
assign g[62378] = b[14] & g[29611];
assign g[45996] = a[14] & g[29612];
assign g[62379] = b[14] & g[29612];
assign g[45997] = a[14] & g[29613];
assign g[62380] = b[14] & g[29613];
assign g[45998] = a[14] & g[29614];
assign g[62381] = b[14] & g[29614];
assign g[45999] = a[14] & g[29615];
assign g[62382] = b[14] & g[29615];
assign g[46000] = a[14] & g[29616];
assign g[62383] = b[14] & g[29616];
assign g[46001] = a[14] & g[29617];
assign g[62384] = b[14] & g[29617];
assign g[46002] = a[14] & g[29618];
assign g[62385] = b[14] & g[29618];
assign g[46003] = a[14] & g[29619];
assign g[62386] = b[14] & g[29619];
assign g[46004] = a[14] & g[29620];
assign g[62387] = b[14] & g[29620];
assign g[46005] = a[14] & g[29621];
assign g[62388] = b[14] & g[29621];
assign g[46006] = a[14] & g[29622];
assign g[62389] = b[14] & g[29622];
assign g[46007] = a[14] & g[29623];
assign g[62390] = b[14] & g[29623];
assign g[46008] = a[14] & g[29624];
assign g[62391] = b[14] & g[29624];
assign g[46009] = a[14] & g[29625];
assign g[62392] = b[14] & g[29625];
assign g[46010] = a[14] & g[29626];
assign g[62393] = b[14] & g[29626];
assign g[46011] = a[14] & g[29627];
assign g[62394] = b[14] & g[29627];
assign g[46012] = a[14] & g[29628];
assign g[62395] = b[14] & g[29628];
assign g[46013] = a[14] & g[29629];
assign g[62396] = b[14] & g[29629];
assign g[46014] = a[14] & g[29630];
assign g[62397] = b[14] & g[29630];
assign g[46015] = a[14] & g[29631];
assign g[62398] = b[14] & g[29631];
assign g[46016] = a[14] & g[29632];
assign g[62399] = b[14] & g[29632];
assign g[46017] = a[14] & g[29633];
assign g[62400] = b[14] & g[29633];
assign g[46018] = a[14] & g[29634];
assign g[62401] = b[14] & g[29634];
assign g[46019] = a[14] & g[29635];
assign g[62402] = b[14] & g[29635];
assign g[46020] = a[14] & g[29636];
assign g[62403] = b[14] & g[29636];
assign g[46021] = a[14] & g[29637];
assign g[62404] = b[14] & g[29637];
assign g[46022] = a[14] & g[29638];
assign g[62405] = b[14] & g[29638];
assign g[46023] = a[14] & g[29639];
assign g[62406] = b[14] & g[29639];
assign g[46024] = a[14] & g[29640];
assign g[62407] = b[14] & g[29640];
assign g[46025] = a[14] & g[29641];
assign g[62408] = b[14] & g[29641];
assign g[46026] = a[14] & g[29642];
assign g[62409] = b[14] & g[29642];
assign g[46027] = a[14] & g[29643];
assign g[62410] = b[14] & g[29643];
assign g[46028] = a[14] & g[29644];
assign g[62411] = b[14] & g[29644];
assign g[46029] = a[14] & g[29645];
assign g[62412] = b[14] & g[29645];
assign g[46030] = a[14] & g[29646];
assign g[62413] = b[14] & g[29646];
assign g[46031] = a[14] & g[29647];
assign g[62414] = b[14] & g[29647];
assign g[46032] = a[14] & g[29648];
assign g[62415] = b[14] & g[29648];
assign g[46033] = a[14] & g[29649];
assign g[62416] = b[14] & g[29649];
assign g[46034] = a[14] & g[29650];
assign g[62417] = b[14] & g[29650];
assign g[46035] = a[14] & g[29651];
assign g[62418] = b[14] & g[29651];
assign g[46036] = a[14] & g[29652];
assign g[62419] = b[14] & g[29652];
assign g[46037] = a[14] & g[29653];
assign g[62420] = b[14] & g[29653];
assign g[46038] = a[14] & g[29654];
assign g[62421] = b[14] & g[29654];
assign g[46039] = a[14] & g[29655];
assign g[62422] = b[14] & g[29655];
assign g[46040] = a[14] & g[29656];
assign g[62423] = b[14] & g[29656];
assign g[46041] = a[14] & g[29657];
assign g[62424] = b[14] & g[29657];
assign g[46042] = a[14] & g[29658];
assign g[62425] = b[14] & g[29658];
assign g[46043] = a[14] & g[29659];
assign g[62426] = b[14] & g[29659];
assign g[46044] = a[14] & g[29660];
assign g[62427] = b[14] & g[29660];
assign g[46045] = a[14] & g[29661];
assign g[62428] = b[14] & g[29661];
assign g[46046] = a[14] & g[29662];
assign g[62429] = b[14] & g[29662];
assign g[46047] = a[14] & g[29663];
assign g[62430] = b[14] & g[29663];
assign g[46048] = a[14] & g[29664];
assign g[62431] = b[14] & g[29664];
assign g[46049] = a[14] & g[29665];
assign g[62432] = b[14] & g[29665];
assign g[46050] = a[14] & g[29666];
assign g[62433] = b[14] & g[29666];
assign g[46051] = a[14] & g[29667];
assign g[62434] = b[14] & g[29667];
assign g[46052] = a[14] & g[29668];
assign g[62435] = b[14] & g[29668];
assign g[46053] = a[14] & g[29669];
assign g[62436] = b[14] & g[29669];
assign g[46054] = a[14] & g[29670];
assign g[62437] = b[14] & g[29670];
assign g[46055] = a[14] & g[29671];
assign g[62438] = b[14] & g[29671];
assign g[46056] = a[14] & g[29672];
assign g[62439] = b[14] & g[29672];
assign g[46057] = a[14] & g[29673];
assign g[62440] = b[14] & g[29673];
assign g[46058] = a[14] & g[29674];
assign g[62441] = b[14] & g[29674];
assign g[46059] = a[14] & g[29675];
assign g[62442] = b[14] & g[29675];
assign g[46060] = a[14] & g[29676];
assign g[62443] = b[14] & g[29676];
assign g[46061] = a[14] & g[29677];
assign g[62444] = b[14] & g[29677];
assign g[46062] = a[14] & g[29678];
assign g[62445] = b[14] & g[29678];
assign g[46063] = a[14] & g[29679];
assign g[62446] = b[14] & g[29679];
assign g[46064] = a[14] & g[29680];
assign g[62447] = b[14] & g[29680];
assign g[46065] = a[14] & g[29681];
assign g[62448] = b[14] & g[29681];
assign g[46066] = a[14] & g[29682];
assign g[62449] = b[14] & g[29682];
assign g[46067] = a[14] & g[29683];
assign g[62450] = b[14] & g[29683];
assign g[46068] = a[14] & g[29684];
assign g[62451] = b[14] & g[29684];
assign g[46069] = a[14] & g[29685];
assign g[62452] = b[14] & g[29685];
assign g[46070] = a[14] & g[29686];
assign g[62453] = b[14] & g[29686];
assign g[46071] = a[14] & g[29687];
assign g[62454] = b[14] & g[29687];
assign g[46072] = a[14] & g[29688];
assign g[62455] = b[14] & g[29688];
assign g[46073] = a[14] & g[29689];
assign g[62456] = b[14] & g[29689];
assign g[46074] = a[14] & g[29690];
assign g[62457] = b[14] & g[29690];
assign g[46075] = a[14] & g[29691];
assign g[62458] = b[14] & g[29691];
assign g[46076] = a[14] & g[29692];
assign g[62459] = b[14] & g[29692];
assign g[46077] = a[14] & g[29693];
assign g[62460] = b[14] & g[29693];
assign g[46078] = a[14] & g[29694];
assign g[62461] = b[14] & g[29694];
assign g[46079] = a[14] & g[29695];
assign g[62462] = b[14] & g[29695];
assign g[46080] = a[14] & g[29696];
assign g[62463] = b[14] & g[29696];
assign g[46081] = a[14] & g[29697];
assign g[62464] = b[14] & g[29697];
assign g[46082] = a[14] & g[29698];
assign g[62465] = b[14] & g[29698];
assign g[46083] = a[14] & g[29699];
assign g[62466] = b[14] & g[29699];
assign g[46084] = a[14] & g[29700];
assign g[62467] = b[14] & g[29700];
assign g[46085] = a[14] & g[29701];
assign g[62468] = b[14] & g[29701];
assign g[46086] = a[14] & g[29702];
assign g[62469] = b[14] & g[29702];
assign g[46087] = a[14] & g[29703];
assign g[62470] = b[14] & g[29703];
assign g[46088] = a[14] & g[29704];
assign g[62471] = b[14] & g[29704];
assign g[46089] = a[14] & g[29705];
assign g[62472] = b[14] & g[29705];
assign g[46090] = a[14] & g[29706];
assign g[62473] = b[14] & g[29706];
assign g[46091] = a[14] & g[29707];
assign g[62474] = b[14] & g[29707];
assign g[46092] = a[14] & g[29708];
assign g[62475] = b[14] & g[29708];
assign g[46093] = a[14] & g[29709];
assign g[62476] = b[14] & g[29709];
assign g[46094] = a[14] & g[29710];
assign g[62477] = b[14] & g[29710];
assign g[46095] = a[14] & g[29711];
assign g[62478] = b[14] & g[29711];
assign g[46096] = a[14] & g[29712];
assign g[62479] = b[14] & g[29712];
assign g[46097] = a[14] & g[29713];
assign g[62480] = b[14] & g[29713];
assign g[46098] = a[14] & g[29714];
assign g[62481] = b[14] & g[29714];
assign g[46099] = a[14] & g[29715];
assign g[62482] = b[14] & g[29715];
assign g[46100] = a[14] & g[29716];
assign g[62483] = b[14] & g[29716];
assign g[46101] = a[14] & g[29717];
assign g[62484] = b[14] & g[29717];
assign g[46102] = a[14] & g[29718];
assign g[62485] = b[14] & g[29718];
assign g[46103] = a[14] & g[29719];
assign g[62486] = b[14] & g[29719];
assign g[46104] = a[14] & g[29720];
assign g[62487] = b[14] & g[29720];
assign g[46105] = a[14] & g[29721];
assign g[62488] = b[14] & g[29721];
assign g[46106] = a[14] & g[29722];
assign g[62489] = b[14] & g[29722];
assign g[46107] = a[14] & g[29723];
assign g[62490] = b[14] & g[29723];
assign g[46108] = a[14] & g[29724];
assign g[62491] = b[14] & g[29724];
assign g[46109] = a[14] & g[29725];
assign g[62492] = b[14] & g[29725];
assign g[46110] = a[14] & g[29726];
assign g[62493] = b[14] & g[29726];
assign g[46111] = a[14] & g[29727];
assign g[62494] = b[14] & g[29727];
assign g[46112] = a[14] & g[29728];
assign g[62495] = b[14] & g[29728];
assign g[46113] = a[14] & g[29729];
assign g[62496] = b[14] & g[29729];
assign g[46114] = a[14] & g[29730];
assign g[62497] = b[14] & g[29730];
assign g[46115] = a[14] & g[29731];
assign g[62498] = b[14] & g[29731];
assign g[46116] = a[14] & g[29732];
assign g[62499] = b[14] & g[29732];
assign g[46117] = a[14] & g[29733];
assign g[62500] = b[14] & g[29733];
assign g[46118] = a[14] & g[29734];
assign g[62501] = b[14] & g[29734];
assign g[46119] = a[14] & g[29735];
assign g[62502] = b[14] & g[29735];
assign g[46120] = a[14] & g[29736];
assign g[62503] = b[14] & g[29736];
assign g[46121] = a[14] & g[29737];
assign g[62504] = b[14] & g[29737];
assign g[46122] = a[14] & g[29738];
assign g[62505] = b[14] & g[29738];
assign g[46123] = a[14] & g[29739];
assign g[62506] = b[14] & g[29739];
assign g[46124] = a[14] & g[29740];
assign g[62507] = b[14] & g[29740];
assign g[46125] = a[14] & g[29741];
assign g[62508] = b[14] & g[29741];
assign g[46126] = a[14] & g[29742];
assign g[62509] = b[14] & g[29742];
assign g[46127] = a[14] & g[29743];
assign g[62510] = b[14] & g[29743];
assign g[46128] = a[14] & g[29744];
assign g[62511] = b[14] & g[29744];
assign g[46129] = a[14] & g[29745];
assign g[62512] = b[14] & g[29745];
assign g[46130] = a[14] & g[29746];
assign g[62513] = b[14] & g[29746];
assign g[46131] = a[14] & g[29747];
assign g[62514] = b[14] & g[29747];
assign g[46132] = a[14] & g[29748];
assign g[62515] = b[14] & g[29748];
assign g[46133] = a[14] & g[29749];
assign g[62516] = b[14] & g[29749];
assign g[46134] = a[14] & g[29750];
assign g[62517] = b[14] & g[29750];
assign g[46135] = a[14] & g[29751];
assign g[62518] = b[14] & g[29751];
assign g[46136] = a[14] & g[29752];
assign g[62519] = b[14] & g[29752];
assign g[46137] = a[14] & g[29753];
assign g[62520] = b[14] & g[29753];
assign g[46138] = a[14] & g[29754];
assign g[62521] = b[14] & g[29754];
assign g[46139] = a[14] & g[29755];
assign g[62522] = b[14] & g[29755];
assign g[46140] = a[14] & g[29756];
assign g[62523] = b[14] & g[29756];
assign g[46141] = a[14] & g[29757];
assign g[62524] = b[14] & g[29757];
assign g[46142] = a[14] & g[29758];
assign g[62525] = b[14] & g[29758];
assign g[46143] = a[14] & g[29759];
assign g[62526] = b[14] & g[29759];
assign g[46144] = a[14] & g[29760];
assign g[62527] = b[14] & g[29760];
assign g[46145] = a[14] & g[29761];
assign g[62528] = b[14] & g[29761];
assign g[46146] = a[14] & g[29762];
assign g[62529] = b[14] & g[29762];
assign g[46147] = a[14] & g[29763];
assign g[62530] = b[14] & g[29763];
assign g[46148] = a[14] & g[29764];
assign g[62531] = b[14] & g[29764];
assign g[46149] = a[14] & g[29765];
assign g[62532] = b[14] & g[29765];
assign g[46150] = a[14] & g[29766];
assign g[62533] = b[14] & g[29766];
assign g[46151] = a[14] & g[29767];
assign g[62534] = b[14] & g[29767];
assign g[46152] = a[14] & g[29768];
assign g[62535] = b[14] & g[29768];
assign g[46153] = a[14] & g[29769];
assign g[62536] = b[14] & g[29769];
assign g[46154] = a[14] & g[29770];
assign g[62537] = b[14] & g[29770];
assign g[46155] = a[14] & g[29771];
assign g[62538] = b[14] & g[29771];
assign g[46156] = a[14] & g[29772];
assign g[62539] = b[14] & g[29772];
assign g[46157] = a[14] & g[29773];
assign g[62540] = b[14] & g[29773];
assign g[46158] = a[14] & g[29774];
assign g[62541] = b[14] & g[29774];
assign g[46159] = a[14] & g[29775];
assign g[62542] = b[14] & g[29775];
assign g[46160] = a[14] & g[29776];
assign g[62543] = b[14] & g[29776];
assign g[46161] = a[14] & g[29777];
assign g[62544] = b[14] & g[29777];
assign g[46162] = a[14] & g[29778];
assign g[62545] = b[14] & g[29778];
assign g[46163] = a[14] & g[29779];
assign g[62546] = b[14] & g[29779];
assign g[46164] = a[14] & g[29780];
assign g[62547] = b[14] & g[29780];
assign g[46165] = a[14] & g[29781];
assign g[62548] = b[14] & g[29781];
assign g[46166] = a[14] & g[29782];
assign g[62549] = b[14] & g[29782];
assign g[46167] = a[14] & g[29783];
assign g[62550] = b[14] & g[29783];
assign g[46168] = a[14] & g[29784];
assign g[62551] = b[14] & g[29784];
assign g[46169] = a[14] & g[29785];
assign g[62552] = b[14] & g[29785];
assign g[46170] = a[14] & g[29786];
assign g[62553] = b[14] & g[29786];
assign g[46171] = a[14] & g[29787];
assign g[62554] = b[14] & g[29787];
assign g[46172] = a[14] & g[29788];
assign g[62555] = b[14] & g[29788];
assign g[46173] = a[14] & g[29789];
assign g[62556] = b[14] & g[29789];
assign g[46174] = a[14] & g[29790];
assign g[62557] = b[14] & g[29790];
assign g[46175] = a[14] & g[29791];
assign g[62558] = b[14] & g[29791];
assign g[46176] = a[14] & g[29792];
assign g[62559] = b[14] & g[29792];
assign g[46177] = a[14] & g[29793];
assign g[62560] = b[14] & g[29793];
assign g[46178] = a[14] & g[29794];
assign g[62561] = b[14] & g[29794];
assign g[46179] = a[14] & g[29795];
assign g[62562] = b[14] & g[29795];
assign g[46180] = a[14] & g[29796];
assign g[62563] = b[14] & g[29796];
assign g[46181] = a[14] & g[29797];
assign g[62564] = b[14] & g[29797];
assign g[46182] = a[14] & g[29798];
assign g[62565] = b[14] & g[29798];
assign g[46183] = a[14] & g[29799];
assign g[62566] = b[14] & g[29799];
assign g[46184] = a[14] & g[29800];
assign g[62567] = b[14] & g[29800];
assign g[46185] = a[14] & g[29801];
assign g[62568] = b[14] & g[29801];
assign g[46186] = a[14] & g[29802];
assign g[62569] = b[14] & g[29802];
assign g[46187] = a[14] & g[29803];
assign g[62570] = b[14] & g[29803];
assign g[46188] = a[14] & g[29804];
assign g[62571] = b[14] & g[29804];
assign g[46189] = a[14] & g[29805];
assign g[62572] = b[14] & g[29805];
assign g[46190] = a[14] & g[29806];
assign g[62573] = b[14] & g[29806];
assign g[46191] = a[14] & g[29807];
assign g[62574] = b[14] & g[29807];
assign g[46192] = a[14] & g[29808];
assign g[62575] = b[14] & g[29808];
assign g[46193] = a[14] & g[29809];
assign g[62576] = b[14] & g[29809];
assign g[46194] = a[14] & g[29810];
assign g[62577] = b[14] & g[29810];
assign g[46195] = a[14] & g[29811];
assign g[62578] = b[14] & g[29811];
assign g[46196] = a[14] & g[29812];
assign g[62579] = b[14] & g[29812];
assign g[46197] = a[14] & g[29813];
assign g[62580] = b[14] & g[29813];
assign g[46198] = a[14] & g[29814];
assign g[62581] = b[14] & g[29814];
assign g[46199] = a[14] & g[29815];
assign g[62582] = b[14] & g[29815];
assign g[46200] = a[14] & g[29816];
assign g[62583] = b[14] & g[29816];
assign g[46201] = a[14] & g[29817];
assign g[62584] = b[14] & g[29817];
assign g[46202] = a[14] & g[29818];
assign g[62585] = b[14] & g[29818];
assign g[46203] = a[14] & g[29819];
assign g[62586] = b[14] & g[29819];
assign g[46204] = a[14] & g[29820];
assign g[62587] = b[14] & g[29820];
assign g[46205] = a[14] & g[29821];
assign g[62588] = b[14] & g[29821];
assign g[46206] = a[14] & g[29822];
assign g[62589] = b[14] & g[29822];
assign g[46207] = a[14] & g[29823];
assign g[62590] = b[14] & g[29823];
assign g[46208] = a[14] & g[29824];
assign g[62591] = b[14] & g[29824];
assign g[46209] = a[14] & g[29825];
assign g[62592] = b[14] & g[29825];
assign g[46210] = a[14] & g[29826];
assign g[62593] = b[14] & g[29826];
assign g[46211] = a[14] & g[29827];
assign g[62594] = b[14] & g[29827];
assign g[46212] = a[14] & g[29828];
assign g[62595] = b[14] & g[29828];
assign g[46213] = a[14] & g[29829];
assign g[62596] = b[14] & g[29829];
assign g[46214] = a[14] & g[29830];
assign g[62597] = b[14] & g[29830];
assign g[46215] = a[14] & g[29831];
assign g[62598] = b[14] & g[29831];
assign g[46216] = a[14] & g[29832];
assign g[62599] = b[14] & g[29832];
assign g[46217] = a[14] & g[29833];
assign g[62600] = b[14] & g[29833];
assign g[46218] = a[14] & g[29834];
assign g[62601] = b[14] & g[29834];
assign g[46219] = a[14] & g[29835];
assign g[62602] = b[14] & g[29835];
assign g[46220] = a[14] & g[29836];
assign g[62603] = b[14] & g[29836];
assign g[46221] = a[14] & g[29837];
assign g[62604] = b[14] & g[29837];
assign g[46222] = a[14] & g[29838];
assign g[62605] = b[14] & g[29838];
assign g[46223] = a[14] & g[29839];
assign g[62606] = b[14] & g[29839];
assign g[46224] = a[14] & g[29840];
assign g[62607] = b[14] & g[29840];
assign g[46225] = a[14] & g[29841];
assign g[62608] = b[14] & g[29841];
assign g[46226] = a[14] & g[29842];
assign g[62609] = b[14] & g[29842];
assign g[46227] = a[14] & g[29843];
assign g[62610] = b[14] & g[29843];
assign g[46228] = a[14] & g[29844];
assign g[62611] = b[14] & g[29844];
assign g[46229] = a[14] & g[29845];
assign g[62612] = b[14] & g[29845];
assign g[46230] = a[14] & g[29846];
assign g[62613] = b[14] & g[29846];
assign g[46231] = a[14] & g[29847];
assign g[62614] = b[14] & g[29847];
assign g[46232] = a[14] & g[29848];
assign g[62615] = b[14] & g[29848];
assign g[46233] = a[14] & g[29849];
assign g[62616] = b[14] & g[29849];
assign g[46234] = a[14] & g[29850];
assign g[62617] = b[14] & g[29850];
assign g[46235] = a[14] & g[29851];
assign g[62618] = b[14] & g[29851];
assign g[46236] = a[14] & g[29852];
assign g[62619] = b[14] & g[29852];
assign g[46237] = a[14] & g[29853];
assign g[62620] = b[14] & g[29853];
assign g[46238] = a[14] & g[29854];
assign g[62621] = b[14] & g[29854];
assign g[46239] = a[14] & g[29855];
assign g[62622] = b[14] & g[29855];
assign g[46240] = a[14] & g[29856];
assign g[62623] = b[14] & g[29856];
assign g[46241] = a[14] & g[29857];
assign g[62624] = b[14] & g[29857];
assign g[46242] = a[14] & g[29858];
assign g[62625] = b[14] & g[29858];
assign g[46243] = a[14] & g[29859];
assign g[62626] = b[14] & g[29859];
assign g[46244] = a[14] & g[29860];
assign g[62627] = b[14] & g[29860];
assign g[46245] = a[14] & g[29861];
assign g[62628] = b[14] & g[29861];
assign g[46246] = a[14] & g[29862];
assign g[62629] = b[14] & g[29862];
assign g[46247] = a[14] & g[29863];
assign g[62630] = b[14] & g[29863];
assign g[46248] = a[14] & g[29864];
assign g[62631] = b[14] & g[29864];
assign g[46249] = a[14] & g[29865];
assign g[62632] = b[14] & g[29865];
assign g[46250] = a[14] & g[29866];
assign g[62633] = b[14] & g[29866];
assign g[46251] = a[14] & g[29867];
assign g[62634] = b[14] & g[29867];
assign g[46252] = a[14] & g[29868];
assign g[62635] = b[14] & g[29868];
assign g[46253] = a[14] & g[29869];
assign g[62636] = b[14] & g[29869];
assign g[46254] = a[14] & g[29870];
assign g[62637] = b[14] & g[29870];
assign g[46255] = a[14] & g[29871];
assign g[62638] = b[14] & g[29871];
assign g[46256] = a[14] & g[29872];
assign g[62639] = b[14] & g[29872];
assign g[46257] = a[14] & g[29873];
assign g[62640] = b[14] & g[29873];
assign g[46258] = a[14] & g[29874];
assign g[62641] = b[14] & g[29874];
assign g[46259] = a[14] & g[29875];
assign g[62642] = b[14] & g[29875];
assign g[46260] = a[14] & g[29876];
assign g[62643] = b[14] & g[29876];
assign g[46261] = a[14] & g[29877];
assign g[62644] = b[14] & g[29877];
assign g[46262] = a[14] & g[29878];
assign g[62645] = b[14] & g[29878];
assign g[46263] = a[14] & g[29879];
assign g[62646] = b[14] & g[29879];
assign g[46264] = a[14] & g[29880];
assign g[62647] = b[14] & g[29880];
assign g[46265] = a[14] & g[29881];
assign g[62648] = b[14] & g[29881];
assign g[46266] = a[14] & g[29882];
assign g[62649] = b[14] & g[29882];
assign g[46267] = a[14] & g[29883];
assign g[62650] = b[14] & g[29883];
assign g[46268] = a[14] & g[29884];
assign g[62651] = b[14] & g[29884];
assign g[46269] = a[14] & g[29885];
assign g[62652] = b[14] & g[29885];
assign g[46270] = a[14] & g[29886];
assign g[62653] = b[14] & g[29886];
assign g[46271] = a[14] & g[29887];
assign g[62654] = b[14] & g[29887];
assign g[46272] = a[14] & g[29888];
assign g[62655] = b[14] & g[29888];
assign g[46273] = a[14] & g[29889];
assign g[62656] = b[14] & g[29889];
assign g[46274] = a[14] & g[29890];
assign g[62657] = b[14] & g[29890];
assign g[46275] = a[14] & g[29891];
assign g[62658] = b[14] & g[29891];
assign g[46276] = a[14] & g[29892];
assign g[62659] = b[14] & g[29892];
assign g[46277] = a[14] & g[29893];
assign g[62660] = b[14] & g[29893];
assign g[46278] = a[14] & g[29894];
assign g[62661] = b[14] & g[29894];
assign g[46279] = a[14] & g[29895];
assign g[62662] = b[14] & g[29895];
assign g[46280] = a[14] & g[29896];
assign g[62663] = b[14] & g[29896];
assign g[46281] = a[14] & g[29897];
assign g[62664] = b[14] & g[29897];
assign g[46282] = a[14] & g[29898];
assign g[62665] = b[14] & g[29898];
assign g[46283] = a[14] & g[29899];
assign g[62666] = b[14] & g[29899];
assign g[46284] = a[14] & g[29900];
assign g[62667] = b[14] & g[29900];
assign g[46285] = a[14] & g[29901];
assign g[62668] = b[14] & g[29901];
assign g[46286] = a[14] & g[29902];
assign g[62669] = b[14] & g[29902];
assign g[46287] = a[14] & g[29903];
assign g[62670] = b[14] & g[29903];
assign g[46288] = a[14] & g[29904];
assign g[62671] = b[14] & g[29904];
assign g[46289] = a[14] & g[29905];
assign g[62672] = b[14] & g[29905];
assign g[46290] = a[14] & g[29906];
assign g[62673] = b[14] & g[29906];
assign g[46291] = a[14] & g[29907];
assign g[62674] = b[14] & g[29907];
assign g[46292] = a[14] & g[29908];
assign g[62675] = b[14] & g[29908];
assign g[46293] = a[14] & g[29909];
assign g[62676] = b[14] & g[29909];
assign g[46294] = a[14] & g[29910];
assign g[62677] = b[14] & g[29910];
assign g[46295] = a[14] & g[29911];
assign g[62678] = b[14] & g[29911];
assign g[46296] = a[14] & g[29912];
assign g[62679] = b[14] & g[29912];
assign g[46297] = a[14] & g[29913];
assign g[62680] = b[14] & g[29913];
assign g[46298] = a[14] & g[29914];
assign g[62681] = b[14] & g[29914];
assign g[46299] = a[14] & g[29915];
assign g[62682] = b[14] & g[29915];
assign g[46300] = a[14] & g[29916];
assign g[62683] = b[14] & g[29916];
assign g[46301] = a[14] & g[29917];
assign g[62684] = b[14] & g[29917];
assign g[46302] = a[14] & g[29918];
assign g[62685] = b[14] & g[29918];
assign g[46303] = a[14] & g[29919];
assign g[62686] = b[14] & g[29919];
assign g[46304] = a[14] & g[29920];
assign g[62687] = b[14] & g[29920];
assign g[46305] = a[14] & g[29921];
assign g[62688] = b[14] & g[29921];
assign g[46306] = a[14] & g[29922];
assign g[62689] = b[14] & g[29922];
assign g[46307] = a[14] & g[29923];
assign g[62690] = b[14] & g[29923];
assign g[46308] = a[14] & g[29924];
assign g[62691] = b[14] & g[29924];
assign g[46309] = a[14] & g[29925];
assign g[62692] = b[14] & g[29925];
assign g[46310] = a[14] & g[29926];
assign g[62693] = b[14] & g[29926];
assign g[46311] = a[14] & g[29927];
assign g[62694] = b[14] & g[29927];
assign g[46312] = a[14] & g[29928];
assign g[62695] = b[14] & g[29928];
assign g[46313] = a[14] & g[29929];
assign g[62696] = b[14] & g[29929];
assign g[46314] = a[14] & g[29930];
assign g[62697] = b[14] & g[29930];
assign g[46315] = a[14] & g[29931];
assign g[62698] = b[14] & g[29931];
assign g[46316] = a[14] & g[29932];
assign g[62699] = b[14] & g[29932];
assign g[46317] = a[14] & g[29933];
assign g[62700] = b[14] & g[29933];
assign g[46318] = a[14] & g[29934];
assign g[62701] = b[14] & g[29934];
assign g[46319] = a[14] & g[29935];
assign g[62702] = b[14] & g[29935];
assign g[46320] = a[14] & g[29936];
assign g[62703] = b[14] & g[29936];
assign g[46321] = a[14] & g[29937];
assign g[62704] = b[14] & g[29937];
assign g[46322] = a[14] & g[29938];
assign g[62705] = b[14] & g[29938];
assign g[46323] = a[14] & g[29939];
assign g[62706] = b[14] & g[29939];
assign g[46324] = a[14] & g[29940];
assign g[62707] = b[14] & g[29940];
assign g[46325] = a[14] & g[29941];
assign g[62708] = b[14] & g[29941];
assign g[46326] = a[14] & g[29942];
assign g[62709] = b[14] & g[29942];
assign g[46327] = a[14] & g[29943];
assign g[62710] = b[14] & g[29943];
assign g[46328] = a[14] & g[29944];
assign g[62711] = b[14] & g[29944];
assign g[46329] = a[14] & g[29945];
assign g[62712] = b[14] & g[29945];
assign g[46330] = a[14] & g[29946];
assign g[62713] = b[14] & g[29946];
assign g[46331] = a[14] & g[29947];
assign g[62714] = b[14] & g[29947];
assign g[46332] = a[14] & g[29948];
assign g[62715] = b[14] & g[29948];
assign g[46333] = a[14] & g[29949];
assign g[62716] = b[14] & g[29949];
assign g[46334] = a[14] & g[29950];
assign g[62717] = b[14] & g[29950];
assign g[46335] = a[14] & g[29951];
assign g[62718] = b[14] & g[29951];
assign g[46336] = a[14] & g[29952];
assign g[62719] = b[14] & g[29952];
assign g[46337] = a[14] & g[29953];
assign g[62720] = b[14] & g[29953];
assign g[46338] = a[14] & g[29954];
assign g[62721] = b[14] & g[29954];
assign g[46339] = a[14] & g[29955];
assign g[62722] = b[14] & g[29955];
assign g[46340] = a[14] & g[29956];
assign g[62723] = b[14] & g[29956];
assign g[46341] = a[14] & g[29957];
assign g[62724] = b[14] & g[29957];
assign g[46342] = a[14] & g[29958];
assign g[62725] = b[14] & g[29958];
assign g[46343] = a[14] & g[29959];
assign g[62726] = b[14] & g[29959];
assign g[46344] = a[14] & g[29960];
assign g[62727] = b[14] & g[29960];
assign g[46345] = a[14] & g[29961];
assign g[62728] = b[14] & g[29961];
assign g[46346] = a[14] & g[29962];
assign g[62729] = b[14] & g[29962];
assign g[46347] = a[14] & g[29963];
assign g[62730] = b[14] & g[29963];
assign g[46348] = a[14] & g[29964];
assign g[62731] = b[14] & g[29964];
assign g[46349] = a[14] & g[29965];
assign g[62732] = b[14] & g[29965];
assign g[46350] = a[14] & g[29966];
assign g[62733] = b[14] & g[29966];
assign g[46351] = a[14] & g[29967];
assign g[62734] = b[14] & g[29967];
assign g[46352] = a[14] & g[29968];
assign g[62735] = b[14] & g[29968];
assign g[46353] = a[14] & g[29969];
assign g[62736] = b[14] & g[29969];
assign g[46354] = a[14] & g[29970];
assign g[62737] = b[14] & g[29970];
assign g[46355] = a[14] & g[29971];
assign g[62738] = b[14] & g[29971];
assign g[46356] = a[14] & g[29972];
assign g[62739] = b[14] & g[29972];
assign g[46357] = a[14] & g[29973];
assign g[62740] = b[14] & g[29973];
assign g[46358] = a[14] & g[29974];
assign g[62741] = b[14] & g[29974];
assign g[46359] = a[14] & g[29975];
assign g[62742] = b[14] & g[29975];
assign g[46360] = a[14] & g[29976];
assign g[62743] = b[14] & g[29976];
assign g[46361] = a[14] & g[29977];
assign g[62744] = b[14] & g[29977];
assign g[46362] = a[14] & g[29978];
assign g[62745] = b[14] & g[29978];
assign g[46363] = a[14] & g[29979];
assign g[62746] = b[14] & g[29979];
assign g[46364] = a[14] & g[29980];
assign g[62747] = b[14] & g[29980];
assign g[46365] = a[14] & g[29981];
assign g[62748] = b[14] & g[29981];
assign g[46366] = a[14] & g[29982];
assign g[62749] = b[14] & g[29982];
assign g[46367] = a[14] & g[29983];
assign g[62750] = b[14] & g[29983];
assign g[46368] = a[14] & g[29984];
assign g[62751] = b[14] & g[29984];
assign g[46369] = a[14] & g[29985];
assign g[62752] = b[14] & g[29985];
assign g[46370] = a[14] & g[29986];
assign g[62753] = b[14] & g[29986];
assign g[46371] = a[14] & g[29987];
assign g[62754] = b[14] & g[29987];
assign g[46372] = a[14] & g[29988];
assign g[62755] = b[14] & g[29988];
assign g[46373] = a[14] & g[29989];
assign g[62756] = b[14] & g[29989];
assign g[46374] = a[14] & g[29990];
assign g[62757] = b[14] & g[29990];
assign g[46375] = a[14] & g[29991];
assign g[62758] = b[14] & g[29991];
assign g[46376] = a[14] & g[29992];
assign g[62759] = b[14] & g[29992];
assign g[46377] = a[14] & g[29993];
assign g[62760] = b[14] & g[29993];
assign g[46378] = a[14] & g[29994];
assign g[62761] = b[14] & g[29994];
assign g[46379] = a[14] & g[29995];
assign g[62762] = b[14] & g[29995];
assign g[46380] = a[14] & g[29996];
assign g[62763] = b[14] & g[29996];
assign g[46381] = a[14] & g[29997];
assign g[62764] = b[14] & g[29997];
assign g[46382] = a[14] & g[29998];
assign g[62765] = b[14] & g[29998];
assign g[46383] = a[14] & g[29999];
assign g[62766] = b[14] & g[29999];
assign g[46384] = a[14] & g[30000];
assign g[62767] = b[14] & g[30000];
assign g[46385] = a[14] & g[30001];
assign g[62768] = b[14] & g[30001];
assign g[46386] = a[14] & g[30002];
assign g[62769] = b[14] & g[30002];
assign g[46387] = a[14] & g[30003];
assign g[62770] = b[14] & g[30003];
assign g[46388] = a[14] & g[30004];
assign g[62771] = b[14] & g[30004];
assign g[46389] = a[14] & g[30005];
assign g[62772] = b[14] & g[30005];
assign g[46390] = a[14] & g[30006];
assign g[62773] = b[14] & g[30006];
assign g[46391] = a[14] & g[30007];
assign g[62774] = b[14] & g[30007];
assign g[46392] = a[14] & g[30008];
assign g[62775] = b[14] & g[30008];
assign g[46393] = a[14] & g[30009];
assign g[62776] = b[14] & g[30009];
assign g[46394] = a[14] & g[30010];
assign g[62777] = b[14] & g[30010];
assign g[46395] = a[14] & g[30011];
assign g[62778] = b[14] & g[30011];
assign g[46396] = a[14] & g[30012];
assign g[62779] = b[14] & g[30012];
assign g[46397] = a[14] & g[30013];
assign g[62780] = b[14] & g[30013];
assign g[46398] = a[14] & g[30014];
assign g[62781] = b[14] & g[30014];
assign g[46399] = a[14] & g[30015];
assign g[62782] = b[14] & g[30015];
assign g[46400] = a[14] & g[30016];
assign g[62783] = b[14] & g[30016];
assign g[46401] = a[14] & g[30017];
assign g[62784] = b[14] & g[30017];
assign g[46402] = a[14] & g[30018];
assign g[62785] = b[14] & g[30018];
assign g[46403] = a[14] & g[30019];
assign g[62786] = b[14] & g[30019];
assign g[46404] = a[14] & g[30020];
assign g[62787] = b[14] & g[30020];
assign g[46405] = a[14] & g[30021];
assign g[62788] = b[14] & g[30021];
assign g[46406] = a[14] & g[30022];
assign g[62789] = b[14] & g[30022];
assign g[46407] = a[14] & g[30023];
assign g[62790] = b[14] & g[30023];
assign g[46408] = a[14] & g[30024];
assign g[62791] = b[14] & g[30024];
assign g[46409] = a[14] & g[30025];
assign g[62792] = b[14] & g[30025];
assign g[46410] = a[14] & g[30026];
assign g[62793] = b[14] & g[30026];
assign g[46411] = a[14] & g[30027];
assign g[62794] = b[14] & g[30027];
assign g[46412] = a[14] & g[30028];
assign g[62795] = b[14] & g[30028];
assign g[46413] = a[14] & g[30029];
assign g[62796] = b[14] & g[30029];
assign g[46414] = a[14] & g[30030];
assign g[62797] = b[14] & g[30030];
assign g[46415] = a[14] & g[30031];
assign g[62798] = b[14] & g[30031];
assign g[46416] = a[14] & g[30032];
assign g[62799] = b[14] & g[30032];
assign g[46417] = a[14] & g[30033];
assign g[62800] = b[14] & g[30033];
assign g[46418] = a[14] & g[30034];
assign g[62801] = b[14] & g[30034];
assign g[46419] = a[14] & g[30035];
assign g[62802] = b[14] & g[30035];
assign g[46420] = a[14] & g[30036];
assign g[62803] = b[14] & g[30036];
assign g[46421] = a[14] & g[30037];
assign g[62804] = b[14] & g[30037];
assign g[46422] = a[14] & g[30038];
assign g[62805] = b[14] & g[30038];
assign g[46423] = a[14] & g[30039];
assign g[62806] = b[14] & g[30039];
assign g[46424] = a[14] & g[30040];
assign g[62807] = b[14] & g[30040];
assign g[46425] = a[14] & g[30041];
assign g[62808] = b[14] & g[30041];
assign g[46426] = a[14] & g[30042];
assign g[62809] = b[14] & g[30042];
assign g[46427] = a[14] & g[30043];
assign g[62810] = b[14] & g[30043];
assign g[46428] = a[14] & g[30044];
assign g[62811] = b[14] & g[30044];
assign g[46429] = a[14] & g[30045];
assign g[62812] = b[14] & g[30045];
assign g[46430] = a[14] & g[30046];
assign g[62813] = b[14] & g[30046];
assign g[46431] = a[14] & g[30047];
assign g[62814] = b[14] & g[30047];
assign g[46432] = a[14] & g[30048];
assign g[62815] = b[14] & g[30048];
assign g[46433] = a[14] & g[30049];
assign g[62816] = b[14] & g[30049];
assign g[46434] = a[14] & g[30050];
assign g[62817] = b[14] & g[30050];
assign g[46435] = a[14] & g[30051];
assign g[62818] = b[14] & g[30051];
assign g[46436] = a[14] & g[30052];
assign g[62819] = b[14] & g[30052];
assign g[46437] = a[14] & g[30053];
assign g[62820] = b[14] & g[30053];
assign g[46438] = a[14] & g[30054];
assign g[62821] = b[14] & g[30054];
assign g[46439] = a[14] & g[30055];
assign g[62822] = b[14] & g[30055];
assign g[46440] = a[14] & g[30056];
assign g[62823] = b[14] & g[30056];
assign g[46441] = a[14] & g[30057];
assign g[62824] = b[14] & g[30057];
assign g[46442] = a[14] & g[30058];
assign g[62825] = b[14] & g[30058];
assign g[46443] = a[14] & g[30059];
assign g[62826] = b[14] & g[30059];
assign g[46444] = a[14] & g[30060];
assign g[62827] = b[14] & g[30060];
assign g[46445] = a[14] & g[30061];
assign g[62828] = b[14] & g[30061];
assign g[46446] = a[14] & g[30062];
assign g[62829] = b[14] & g[30062];
assign g[46447] = a[14] & g[30063];
assign g[62830] = b[14] & g[30063];
assign g[46448] = a[14] & g[30064];
assign g[62831] = b[14] & g[30064];
assign g[46449] = a[14] & g[30065];
assign g[62832] = b[14] & g[30065];
assign g[46450] = a[14] & g[30066];
assign g[62833] = b[14] & g[30066];
assign g[46451] = a[14] & g[30067];
assign g[62834] = b[14] & g[30067];
assign g[46452] = a[14] & g[30068];
assign g[62835] = b[14] & g[30068];
assign g[46453] = a[14] & g[30069];
assign g[62836] = b[14] & g[30069];
assign g[46454] = a[14] & g[30070];
assign g[62837] = b[14] & g[30070];
assign g[46455] = a[14] & g[30071];
assign g[62838] = b[14] & g[30071];
assign g[46456] = a[14] & g[30072];
assign g[62839] = b[14] & g[30072];
assign g[46457] = a[14] & g[30073];
assign g[62840] = b[14] & g[30073];
assign g[46458] = a[14] & g[30074];
assign g[62841] = b[14] & g[30074];
assign g[46459] = a[14] & g[30075];
assign g[62842] = b[14] & g[30075];
assign g[46460] = a[14] & g[30076];
assign g[62843] = b[14] & g[30076];
assign g[46461] = a[14] & g[30077];
assign g[62844] = b[14] & g[30077];
assign g[46462] = a[14] & g[30078];
assign g[62845] = b[14] & g[30078];
assign g[46463] = a[14] & g[30079];
assign g[62846] = b[14] & g[30079];
assign g[46464] = a[14] & g[30080];
assign g[62847] = b[14] & g[30080];
assign g[46465] = a[14] & g[30081];
assign g[62848] = b[14] & g[30081];
assign g[46466] = a[14] & g[30082];
assign g[62849] = b[14] & g[30082];
assign g[46467] = a[14] & g[30083];
assign g[62850] = b[14] & g[30083];
assign g[46468] = a[14] & g[30084];
assign g[62851] = b[14] & g[30084];
assign g[46469] = a[14] & g[30085];
assign g[62852] = b[14] & g[30085];
assign g[46470] = a[14] & g[30086];
assign g[62853] = b[14] & g[30086];
assign g[46471] = a[14] & g[30087];
assign g[62854] = b[14] & g[30087];
assign g[46472] = a[14] & g[30088];
assign g[62855] = b[14] & g[30088];
assign g[46473] = a[14] & g[30089];
assign g[62856] = b[14] & g[30089];
assign g[46474] = a[14] & g[30090];
assign g[62857] = b[14] & g[30090];
assign g[46475] = a[14] & g[30091];
assign g[62858] = b[14] & g[30091];
assign g[46476] = a[14] & g[30092];
assign g[62859] = b[14] & g[30092];
assign g[46477] = a[14] & g[30093];
assign g[62860] = b[14] & g[30093];
assign g[46478] = a[14] & g[30094];
assign g[62861] = b[14] & g[30094];
assign g[46479] = a[14] & g[30095];
assign g[62862] = b[14] & g[30095];
assign g[46480] = a[14] & g[30096];
assign g[62863] = b[14] & g[30096];
assign g[46481] = a[14] & g[30097];
assign g[62864] = b[14] & g[30097];
assign g[46482] = a[14] & g[30098];
assign g[62865] = b[14] & g[30098];
assign g[46483] = a[14] & g[30099];
assign g[62866] = b[14] & g[30099];
assign g[46484] = a[14] & g[30100];
assign g[62867] = b[14] & g[30100];
assign g[46485] = a[14] & g[30101];
assign g[62868] = b[14] & g[30101];
assign g[46486] = a[14] & g[30102];
assign g[62869] = b[14] & g[30102];
assign g[46487] = a[14] & g[30103];
assign g[62870] = b[14] & g[30103];
assign g[46488] = a[14] & g[30104];
assign g[62871] = b[14] & g[30104];
assign g[46489] = a[14] & g[30105];
assign g[62872] = b[14] & g[30105];
assign g[46490] = a[14] & g[30106];
assign g[62873] = b[14] & g[30106];
assign g[46491] = a[14] & g[30107];
assign g[62874] = b[14] & g[30107];
assign g[46492] = a[14] & g[30108];
assign g[62875] = b[14] & g[30108];
assign g[46493] = a[14] & g[30109];
assign g[62876] = b[14] & g[30109];
assign g[46494] = a[14] & g[30110];
assign g[62877] = b[14] & g[30110];
assign g[46495] = a[14] & g[30111];
assign g[62878] = b[14] & g[30111];
assign g[46496] = a[14] & g[30112];
assign g[62879] = b[14] & g[30112];
assign g[46497] = a[14] & g[30113];
assign g[62880] = b[14] & g[30113];
assign g[46498] = a[14] & g[30114];
assign g[62881] = b[14] & g[30114];
assign g[46499] = a[14] & g[30115];
assign g[62882] = b[14] & g[30115];
assign g[46500] = a[14] & g[30116];
assign g[62883] = b[14] & g[30116];
assign g[46501] = a[14] & g[30117];
assign g[62884] = b[14] & g[30117];
assign g[46502] = a[14] & g[30118];
assign g[62885] = b[14] & g[30118];
assign g[46503] = a[14] & g[30119];
assign g[62886] = b[14] & g[30119];
assign g[46504] = a[14] & g[30120];
assign g[62887] = b[14] & g[30120];
assign g[46505] = a[14] & g[30121];
assign g[62888] = b[14] & g[30121];
assign g[46506] = a[14] & g[30122];
assign g[62889] = b[14] & g[30122];
assign g[46507] = a[14] & g[30123];
assign g[62890] = b[14] & g[30123];
assign g[46508] = a[14] & g[30124];
assign g[62891] = b[14] & g[30124];
assign g[46509] = a[14] & g[30125];
assign g[62892] = b[14] & g[30125];
assign g[46510] = a[14] & g[30126];
assign g[62893] = b[14] & g[30126];
assign g[46511] = a[14] & g[30127];
assign g[62894] = b[14] & g[30127];
assign g[46512] = a[14] & g[30128];
assign g[62895] = b[14] & g[30128];
assign g[46513] = a[14] & g[30129];
assign g[62896] = b[14] & g[30129];
assign g[46514] = a[14] & g[30130];
assign g[62897] = b[14] & g[30130];
assign g[46515] = a[14] & g[30131];
assign g[62898] = b[14] & g[30131];
assign g[46516] = a[14] & g[30132];
assign g[62899] = b[14] & g[30132];
assign g[46517] = a[14] & g[30133];
assign g[62900] = b[14] & g[30133];
assign g[46518] = a[14] & g[30134];
assign g[62901] = b[14] & g[30134];
assign g[46519] = a[14] & g[30135];
assign g[62902] = b[14] & g[30135];
assign g[46520] = a[14] & g[30136];
assign g[62903] = b[14] & g[30136];
assign g[46521] = a[14] & g[30137];
assign g[62904] = b[14] & g[30137];
assign g[46522] = a[14] & g[30138];
assign g[62905] = b[14] & g[30138];
assign g[46523] = a[14] & g[30139];
assign g[62906] = b[14] & g[30139];
assign g[46524] = a[14] & g[30140];
assign g[62907] = b[14] & g[30140];
assign g[46525] = a[14] & g[30141];
assign g[62908] = b[14] & g[30141];
assign g[46526] = a[14] & g[30142];
assign g[62909] = b[14] & g[30142];
assign g[46527] = a[14] & g[30143];
assign g[62910] = b[14] & g[30143];
assign g[46528] = a[14] & g[30144];
assign g[62911] = b[14] & g[30144];
assign g[46529] = a[14] & g[30145];
assign g[62912] = b[14] & g[30145];
assign g[46530] = a[14] & g[30146];
assign g[62913] = b[14] & g[30146];
assign g[46531] = a[14] & g[30147];
assign g[62914] = b[14] & g[30147];
assign g[46532] = a[14] & g[30148];
assign g[62915] = b[14] & g[30148];
assign g[46533] = a[14] & g[30149];
assign g[62916] = b[14] & g[30149];
assign g[46534] = a[14] & g[30150];
assign g[62917] = b[14] & g[30150];
assign g[46535] = a[14] & g[30151];
assign g[62918] = b[14] & g[30151];
assign g[46536] = a[14] & g[30152];
assign g[62919] = b[14] & g[30152];
assign g[46537] = a[14] & g[30153];
assign g[62920] = b[14] & g[30153];
assign g[46538] = a[14] & g[30154];
assign g[62921] = b[14] & g[30154];
assign g[46539] = a[14] & g[30155];
assign g[62922] = b[14] & g[30155];
assign g[46540] = a[14] & g[30156];
assign g[62923] = b[14] & g[30156];
assign g[46541] = a[14] & g[30157];
assign g[62924] = b[14] & g[30157];
assign g[46542] = a[14] & g[30158];
assign g[62925] = b[14] & g[30158];
assign g[46543] = a[14] & g[30159];
assign g[62926] = b[14] & g[30159];
assign g[46544] = a[14] & g[30160];
assign g[62927] = b[14] & g[30160];
assign g[46545] = a[14] & g[30161];
assign g[62928] = b[14] & g[30161];
assign g[46546] = a[14] & g[30162];
assign g[62929] = b[14] & g[30162];
assign g[46547] = a[14] & g[30163];
assign g[62930] = b[14] & g[30163];
assign g[46548] = a[14] & g[30164];
assign g[62931] = b[14] & g[30164];
assign g[46549] = a[14] & g[30165];
assign g[62932] = b[14] & g[30165];
assign g[46550] = a[14] & g[30166];
assign g[62933] = b[14] & g[30166];
assign g[46551] = a[14] & g[30167];
assign g[62934] = b[14] & g[30167];
assign g[46552] = a[14] & g[30168];
assign g[62935] = b[14] & g[30168];
assign g[46553] = a[14] & g[30169];
assign g[62936] = b[14] & g[30169];
assign g[46554] = a[14] & g[30170];
assign g[62937] = b[14] & g[30170];
assign g[46555] = a[14] & g[30171];
assign g[62938] = b[14] & g[30171];
assign g[46556] = a[14] & g[30172];
assign g[62939] = b[14] & g[30172];
assign g[46557] = a[14] & g[30173];
assign g[62940] = b[14] & g[30173];
assign g[46558] = a[14] & g[30174];
assign g[62941] = b[14] & g[30174];
assign g[46559] = a[14] & g[30175];
assign g[62942] = b[14] & g[30175];
assign g[46560] = a[14] & g[30176];
assign g[62943] = b[14] & g[30176];
assign g[46561] = a[14] & g[30177];
assign g[62944] = b[14] & g[30177];
assign g[46562] = a[14] & g[30178];
assign g[62945] = b[14] & g[30178];
assign g[46563] = a[14] & g[30179];
assign g[62946] = b[14] & g[30179];
assign g[46564] = a[14] & g[30180];
assign g[62947] = b[14] & g[30180];
assign g[46565] = a[14] & g[30181];
assign g[62948] = b[14] & g[30181];
assign g[46566] = a[14] & g[30182];
assign g[62949] = b[14] & g[30182];
assign g[46567] = a[14] & g[30183];
assign g[62950] = b[14] & g[30183];
assign g[46568] = a[14] & g[30184];
assign g[62951] = b[14] & g[30184];
assign g[46569] = a[14] & g[30185];
assign g[62952] = b[14] & g[30185];
assign g[46570] = a[14] & g[30186];
assign g[62953] = b[14] & g[30186];
assign g[46571] = a[14] & g[30187];
assign g[62954] = b[14] & g[30187];
assign g[46572] = a[14] & g[30188];
assign g[62955] = b[14] & g[30188];
assign g[46573] = a[14] & g[30189];
assign g[62956] = b[14] & g[30189];
assign g[46574] = a[14] & g[30190];
assign g[62957] = b[14] & g[30190];
assign g[46575] = a[14] & g[30191];
assign g[62958] = b[14] & g[30191];
assign g[46576] = a[14] & g[30192];
assign g[62959] = b[14] & g[30192];
assign g[46577] = a[14] & g[30193];
assign g[62960] = b[14] & g[30193];
assign g[46578] = a[14] & g[30194];
assign g[62961] = b[14] & g[30194];
assign g[46579] = a[14] & g[30195];
assign g[62962] = b[14] & g[30195];
assign g[46580] = a[14] & g[30196];
assign g[62963] = b[14] & g[30196];
assign g[46581] = a[14] & g[30197];
assign g[62964] = b[14] & g[30197];
assign g[46582] = a[14] & g[30198];
assign g[62965] = b[14] & g[30198];
assign g[46583] = a[14] & g[30199];
assign g[62966] = b[14] & g[30199];
assign g[46584] = a[14] & g[30200];
assign g[62967] = b[14] & g[30200];
assign g[46585] = a[14] & g[30201];
assign g[62968] = b[14] & g[30201];
assign g[46586] = a[14] & g[30202];
assign g[62969] = b[14] & g[30202];
assign g[46587] = a[14] & g[30203];
assign g[62970] = b[14] & g[30203];
assign g[46588] = a[14] & g[30204];
assign g[62971] = b[14] & g[30204];
assign g[46589] = a[14] & g[30205];
assign g[62972] = b[14] & g[30205];
assign g[46590] = a[14] & g[30206];
assign g[62973] = b[14] & g[30206];
assign g[46591] = a[14] & g[30207];
assign g[62974] = b[14] & g[30207];
assign g[46592] = a[14] & g[30208];
assign g[62975] = b[14] & g[30208];
assign g[46593] = a[14] & g[30209];
assign g[62976] = b[14] & g[30209];
assign g[46594] = a[14] & g[30210];
assign g[62977] = b[14] & g[30210];
assign g[46595] = a[14] & g[30211];
assign g[62978] = b[14] & g[30211];
assign g[46596] = a[14] & g[30212];
assign g[62979] = b[14] & g[30212];
assign g[46597] = a[14] & g[30213];
assign g[62980] = b[14] & g[30213];
assign g[46598] = a[14] & g[30214];
assign g[62981] = b[14] & g[30214];
assign g[46599] = a[14] & g[30215];
assign g[62982] = b[14] & g[30215];
assign g[46600] = a[14] & g[30216];
assign g[62983] = b[14] & g[30216];
assign g[46601] = a[14] & g[30217];
assign g[62984] = b[14] & g[30217];
assign g[46602] = a[14] & g[30218];
assign g[62985] = b[14] & g[30218];
assign g[46603] = a[14] & g[30219];
assign g[62986] = b[14] & g[30219];
assign g[46604] = a[14] & g[30220];
assign g[62987] = b[14] & g[30220];
assign g[46605] = a[14] & g[30221];
assign g[62988] = b[14] & g[30221];
assign g[46606] = a[14] & g[30222];
assign g[62989] = b[14] & g[30222];
assign g[46607] = a[14] & g[30223];
assign g[62990] = b[14] & g[30223];
assign g[46608] = a[14] & g[30224];
assign g[62991] = b[14] & g[30224];
assign g[46609] = a[14] & g[30225];
assign g[62992] = b[14] & g[30225];
assign g[46610] = a[14] & g[30226];
assign g[62993] = b[14] & g[30226];
assign g[46611] = a[14] & g[30227];
assign g[62994] = b[14] & g[30227];
assign g[46612] = a[14] & g[30228];
assign g[62995] = b[14] & g[30228];
assign g[46613] = a[14] & g[30229];
assign g[62996] = b[14] & g[30229];
assign g[46614] = a[14] & g[30230];
assign g[62997] = b[14] & g[30230];
assign g[46615] = a[14] & g[30231];
assign g[62998] = b[14] & g[30231];
assign g[46616] = a[14] & g[30232];
assign g[62999] = b[14] & g[30232];
assign g[46617] = a[14] & g[30233];
assign g[63000] = b[14] & g[30233];
assign g[46618] = a[14] & g[30234];
assign g[63001] = b[14] & g[30234];
assign g[46619] = a[14] & g[30235];
assign g[63002] = b[14] & g[30235];
assign g[46620] = a[14] & g[30236];
assign g[63003] = b[14] & g[30236];
assign g[46621] = a[14] & g[30237];
assign g[63004] = b[14] & g[30237];
assign g[46622] = a[14] & g[30238];
assign g[63005] = b[14] & g[30238];
assign g[46623] = a[14] & g[30239];
assign g[63006] = b[14] & g[30239];
assign g[46624] = a[14] & g[30240];
assign g[63007] = b[14] & g[30240];
assign g[46625] = a[14] & g[30241];
assign g[63008] = b[14] & g[30241];
assign g[46626] = a[14] & g[30242];
assign g[63009] = b[14] & g[30242];
assign g[46627] = a[14] & g[30243];
assign g[63010] = b[14] & g[30243];
assign g[46628] = a[14] & g[30244];
assign g[63011] = b[14] & g[30244];
assign g[46629] = a[14] & g[30245];
assign g[63012] = b[14] & g[30245];
assign g[46630] = a[14] & g[30246];
assign g[63013] = b[14] & g[30246];
assign g[46631] = a[14] & g[30247];
assign g[63014] = b[14] & g[30247];
assign g[46632] = a[14] & g[30248];
assign g[63015] = b[14] & g[30248];
assign g[46633] = a[14] & g[30249];
assign g[63016] = b[14] & g[30249];
assign g[46634] = a[14] & g[30250];
assign g[63017] = b[14] & g[30250];
assign g[46635] = a[14] & g[30251];
assign g[63018] = b[14] & g[30251];
assign g[46636] = a[14] & g[30252];
assign g[63019] = b[14] & g[30252];
assign g[46637] = a[14] & g[30253];
assign g[63020] = b[14] & g[30253];
assign g[46638] = a[14] & g[30254];
assign g[63021] = b[14] & g[30254];
assign g[46639] = a[14] & g[30255];
assign g[63022] = b[14] & g[30255];
assign g[46640] = a[14] & g[30256];
assign g[63023] = b[14] & g[30256];
assign g[46641] = a[14] & g[30257];
assign g[63024] = b[14] & g[30257];
assign g[46642] = a[14] & g[30258];
assign g[63025] = b[14] & g[30258];
assign g[46643] = a[14] & g[30259];
assign g[63026] = b[14] & g[30259];
assign g[46644] = a[14] & g[30260];
assign g[63027] = b[14] & g[30260];
assign g[46645] = a[14] & g[30261];
assign g[63028] = b[14] & g[30261];
assign g[46646] = a[14] & g[30262];
assign g[63029] = b[14] & g[30262];
assign g[46647] = a[14] & g[30263];
assign g[63030] = b[14] & g[30263];
assign g[46648] = a[14] & g[30264];
assign g[63031] = b[14] & g[30264];
assign g[46649] = a[14] & g[30265];
assign g[63032] = b[14] & g[30265];
assign g[46650] = a[14] & g[30266];
assign g[63033] = b[14] & g[30266];
assign g[46651] = a[14] & g[30267];
assign g[63034] = b[14] & g[30267];
assign g[46652] = a[14] & g[30268];
assign g[63035] = b[14] & g[30268];
assign g[46653] = a[14] & g[30269];
assign g[63036] = b[14] & g[30269];
assign g[46654] = a[14] & g[30270];
assign g[63037] = b[14] & g[30270];
assign g[46655] = a[14] & g[30271];
assign g[63038] = b[14] & g[30271];
assign g[46656] = a[14] & g[30272];
assign g[63039] = b[14] & g[30272];
assign g[46657] = a[14] & g[30273];
assign g[63040] = b[14] & g[30273];
assign g[46658] = a[14] & g[30274];
assign g[63041] = b[14] & g[30274];
assign g[46659] = a[14] & g[30275];
assign g[63042] = b[14] & g[30275];
assign g[46660] = a[14] & g[30276];
assign g[63043] = b[14] & g[30276];
assign g[46661] = a[14] & g[30277];
assign g[63044] = b[14] & g[30277];
assign g[46662] = a[14] & g[30278];
assign g[63045] = b[14] & g[30278];
assign g[46663] = a[14] & g[30279];
assign g[63046] = b[14] & g[30279];
assign g[46664] = a[14] & g[30280];
assign g[63047] = b[14] & g[30280];
assign g[46665] = a[14] & g[30281];
assign g[63048] = b[14] & g[30281];
assign g[46666] = a[14] & g[30282];
assign g[63049] = b[14] & g[30282];
assign g[46667] = a[14] & g[30283];
assign g[63050] = b[14] & g[30283];
assign g[46668] = a[14] & g[30284];
assign g[63051] = b[14] & g[30284];
assign g[46669] = a[14] & g[30285];
assign g[63052] = b[14] & g[30285];
assign g[46670] = a[14] & g[30286];
assign g[63053] = b[14] & g[30286];
assign g[46671] = a[14] & g[30287];
assign g[63054] = b[14] & g[30287];
assign g[46672] = a[14] & g[30288];
assign g[63055] = b[14] & g[30288];
assign g[46673] = a[14] & g[30289];
assign g[63056] = b[14] & g[30289];
assign g[46674] = a[14] & g[30290];
assign g[63057] = b[14] & g[30290];
assign g[46675] = a[14] & g[30291];
assign g[63058] = b[14] & g[30291];
assign g[46676] = a[14] & g[30292];
assign g[63059] = b[14] & g[30292];
assign g[46677] = a[14] & g[30293];
assign g[63060] = b[14] & g[30293];
assign g[46678] = a[14] & g[30294];
assign g[63061] = b[14] & g[30294];
assign g[46679] = a[14] & g[30295];
assign g[63062] = b[14] & g[30295];
assign g[46680] = a[14] & g[30296];
assign g[63063] = b[14] & g[30296];
assign g[46681] = a[14] & g[30297];
assign g[63064] = b[14] & g[30297];
assign g[46682] = a[14] & g[30298];
assign g[63065] = b[14] & g[30298];
assign g[46683] = a[14] & g[30299];
assign g[63066] = b[14] & g[30299];
assign g[46684] = a[14] & g[30300];
assign g[63067] = b[14] & g[30300];
assign g[46685] = a[14] & g[30301];
assign g[63068] = b[14] & g[30301];
assign g[46686] = a[14] & g[30302];
assign g[63069] = b[14] & g[30302];
assign g[46687] = a[14] & g[30303];
assign g[63070] = b[14] & g[30303];
assign g[46688] = a[14] & g[30304];
assign g[63071] = b[14] & g[30304];
assign g[46689] = a[14] & g[30305];
assign g[63072] = b[14] & g[30305];
assign g[46690] = a[14] & g[30306];
assign g[63073] = b[14] & g[30306];
assign g[46691] = a[14] & g[30307];
assign g[63074] = b[14] & g[30307];
assign g[46692] = a[14] & g[30308];
assign g[63075] = b[14] & g[30308];
assign g[46693] = a[14] & g[30309];
assign g[63076] = b[14] & g[30309];
assign g[46694] = a[14] & g[30310];
assign g[63077] = b[14] & g[30310];
assign g[46695] = a[14] & g[30311];
assign g[63078] = b[14] & g[30311];
assign g[46696] = a[14] & g[30312];
assign g[63079] = b[14] & g[30312];
assign g[46697] = a[14] & g[30313];
assign g[63080] = b[14] & g[30313];
assign g[46698] = a[14] & g[30314];
assign g[63081] = b[14] & g[30314];
assign g[46699] = a[14] & g[30315];
assign g[63082] = b[14] & g[30315];
assign g[46700] = a[14] & g[30316];
assign g[63083] = b[14] & g[30316];
assign g[46701] = a[14] & g[30317];
assign g[63084] = b[14] & g[30317];
assign g[46702] = a[14] & g[30318];
assign g[63085] = b[14] & g[30318];
assign g[46703] = a[14] & g[30319];
assign g[63086] = b[14] & g[30319];
assign g[46704] = a[14] & g[30320];
assign g[63087] = b[14] & g[30320];
assign g[46705] = a[14] & g[30321];
assign g[63088] = b[14] & g[30321];
assign g[46706] = a[14] & g[30322];
assign g[63089] = b[14] & g[30322];
assign g[46707] = a[14] & g[30323];
assign g[63090] = b[14] & g[30323];
assign g[46708] = a[14] & g[30324];
assign g[63091] = b[14] & g[30324];
assign g[46709] = a[14] & g[30325];
assign g[63092] = b[14] & g[30325];
assign g[46710] = a[14] & g[30326];
assign g[63093] = b[14] & g[30326];
assign g[46711] = a[14] & g[30327];
assign g[63094] = b[14] & g[30327];
assign g[46712] = a[14] & g[30328];
assign g[63095] = b[14] & g[30328];
assign g[46713] = a[14] & g[30329];
assign g[63096] = b[14] & g[30329];
assign g[46714] = a[14] & g[30330];
assign g[63097] = b[14] & g[30330];
assign g[46715] = a[14] & g[30331];
assign g[63098] = b[14] & g[30331];
assign g[46716] = a[14] & g[30332];
assign g[63099] = b[14] & g[30332];
assign g[46717] = a[14] & g[30333];
assign g[63100] = b[14] & g[30333];
assign g[46718] = a[14] & g[30334];
assign g[63101] = b[14] & g[30334];
assign g[46719] = a[14] & g[30335];
assign g[63102] = b[14] & g[30335];
assign g[46720] = a[14] & g[30336];
assign g[63103] = b[14] & g[30336];
assign g[46721] = a[14] & g[30337];
assign g[63104] = b[14] & g[30337];
assign g[46722] = a[14] & g[30338];
assign g[63105] = b[14] & g[30338];
assign g[46723] = a[14] & g[30339];
assign g[63106] = b[14] & g[30339];
assign g[46724] = a[14] & g[30340];
assign g[63107] = b[14] & g[30340];
assign g[46725] = a[14] & g[30341];
assign g[63108] = b[14] & g[30341];
assign g[46726] = a[14] & g[30342];
assign g[63109] = b[14] & g[30342];
assign g[46727] = a[14] & g[30343];
assign g[63110] = b[14] & g[30343];
assign g[46728] = a[14] & g[30344];
assign g[63111] = b[14] & g[30344];
assign g[46729] = a[14] & g[30345];
assign g[63112] = b[14] & g[30345];
assign g[46730] = a[14] & g[30346];
assign g[63113] = b[14] & g[30346];
assign g[46731] = a[14] & g[30347];
assign g[63114] = b[14] & g[30347];
assign g[46732] = a[14] & g[30348];
assign g[63115] = b[14] & g[30348];
assign g[46733] = a[14] & g[30349];
assign g[63116] = b[14] & g[30349];
assign g[46734] = a[14] & g[30350];
assign g[63117] = b[14] & g[30350];
assign g[46735] = a[14] & g[30351];
assign g[63118] = b[14] & g[30351];
assign g[46736] = a[14] & g[30352];
assign g[63119] = b[14] & g[30352];
assign g[46737] = a[14] & g[30353];
assign g[63120] = b[14] & g[30353];
assign g[46738] = a[14] & g[30354];
assign g[63121] = b[14] & g[30354];
assign g[46739] = a[14] & g[30355];
assign g[63122] = b[14] & g[30355];
assign g[46740] = a[14] & g[30356];
assign g[63123] = b[14] & g[30356];
assign g[46741] = a[14] & g[30357];
assign g[63124] = b[14] & g[30357];
assign g[46742] = a[14] & g[30358];
assign g[63125] = b[14] & g[30358];
assign g[46743] = a[14] & g[30359];
assign g[63126] = b[14] & g[30359];
assign g[46744] = a[14] & g[30360];
assign g[63127] = b[14] & g[30360];
assign g[46745] = a[14] & g[30361];
assign g[63128] = b[14] & g[30361];
assign g[46746] = a[14] & g[30362];
assign g[63129] = b[14] & g[30362];
assign g[46747] = a[14] & g[30363];
assign g[63130] = b[14] & g[30363];
assign g[46748] = a[14] & g[30364];
assign g[63131] = b[14] & g[30364];
assign g[46749] = a[14] & g[30365];
assign g[63132] = b[14] & g[30365];
assign g[46750] = a[14] & g[30366];
assign g[63133] = b[14] & g[30366];
assign g[46751] = a[14] & g[30367];
assign g[63134] = b[14] & g[30367];
assign g[46752] = a[14] & g[30368];
assign g[63135] = b[14] & g[30368];
assign g[46753] = a[14] & g[30369];
assign g[63136] = b[14] & g[30369];
assign g[46754] = a[14] & g[30370];
assign g[63137] = b[14] & g[30370];
assign g[46755] = a[14] & g[30371];
assign g[63138] = b[14] & g[30371];
assign g[46756] = a[14] & g[30372];
assign g[63139] = b[14] & g[30372];
assign g[46757] = a[14] & g[30373];
assign g[63140] = b[14] & g[30373];
assign g[46758] = a[14] & g[30374];
assign g[63141] = b[14] & g[30374];
assign g[46759] = a[14] & g[30375];
assign g[63142] = b[14] & g[30375];
assign g[46760] = a[14] & g[30376];
assign g[63143] = b[14] & g[30376];
assign g[46761] = a[14] & g[30377];
assign g[63144] = b[14] & g[30377];
assign g[46762] = a[14] & g[30378];
assign g[63145] = b[14] & g[30378];
assign g[46763] = a[14] & g[30379];
assign g[63146] = b[14] & g[30379];
assign g[46764] = a[14] & g[30380];
assign g[63147] = b[14] & g[30380];
assign g[46765] = a[14] & g[30381];
assign g[63148] = b[14] & g[30381];
assign g[46766] = a[14] & g[30382];
assign g[63149] = b[14] & g[30382];
assign g[46767] = a[14] & g[30383];
assign g[63150] = b[14] & g[30383];
assign g[46768] = a[14] & g[30384];
assign g[63151] = b[14] & g[30384];
assign g[46769] = a[14] & g[30385];
assign g[63152] = b[14] & g[30385];
assign g[46770] = a[14] & g[30386];
assign g[63153] = b[14] & g[30386];
assign g[46771] = a[14] & g[30387];
assign g[63154] = b[14] & g[30387];
assign g[46772] = a[14] & g[30388];
assign g[63155] = b[14] & g[30388];
assign g[46773] = a[14] & g[30389];
assign g[63156] = b[14] & g[30389];
assign g[46774] = a[14] & g[30390];
assign g[63157] = b[14] & g[30390];
assign g[46775] = a[14] & g[30391];
assign g[63158] = b[14] & g[30391];
assign g[46776] = a[14] & g[30392];
assign g[63159] = b[14] & g[30392];
assign g[46777] = a[14] & g[30393];
assign g[63160] = b[14] & g[30393];
assign g[46778] = a[14] & g[30394];
assign g[63161] = b[14] & g[30394];
assign g[46779] = a[14] & g[30395];
assign g[63162] = b[14] & g[30395];
assign g[46780] = a[14] & g[30396];
assign g[63163] = b[14] & g[30396];
assign g[46781] = a[14] & g[30397];
assign g[63164] = b[14] & g[30397];
assign g[46782] = a[14] & g[30398];
assign g[63165] = b[14] & g[30398];
assign g[46783] = a[14] & g[30399];
assign g[63166] = b[14] & g[30399];
assign g[46784] = a[14] & g[30400];
assign g[63167] = b[14] & g[30400];
assign g[46785] = a[14] & g[30401];
assign g[63168] = b[14] & g[30401];
assign g[46786] = a[14] & g[30402];
assign g[63169] = b[14] & g[30402];
assign g[46787] = a[14] & g[30403];
assign g[63170] = b[14] & g[30403];
assign g[46788] = a[14] & g[30404];
assign g[63171] = b[14] & g[30404];
assign g[46789] = a[14] & g[30405];
assign g[63172] = b[14] & g[30405];
assign g[46790] = a[14] & g[30406];
assign g[63173] = b[14] & g[30406];
assign g[46791] = a[14] & g[30407];
assign g[63174] = b[14] & g[30407];
assign g[46792] = a[14] & g[30408];
assign g[63175] = b[14] & g[30408];
assign g[46793] = a[14] & g[30409];
assign g[63176] = b[14] & g[30409];
assign g[46794] = a[14] & g[30410];
assign g[63177] = b[14] & g[30410];
assign g[46795] = a[14] & g[30411];
assign g[63178] = b[14] & g[30411];
assign g[46796] = a[14] & g[30412];
assign g[63179] = b[14] & g[30412];
assign g[46797] = a[14] & g[30413];
assign g[63180] = b[14] & g[30413];
assign g[46798] = a[14] & g[30414];
assign g[63181] = b[14] & g[30414];
assign g[46799] = a[14] & g[30415];
assign g[63182] = b[14] & g[30415];
assign g[46800] = a[14] & g[30416];
assign g[63183] = b[14] & g[30416];
assign g[46801] = a[14] & g[30417];
assign g[63184] = b[14] & g[30417];
assign g[46802] = a[14] & g[30418];
assign g[63185] = b[14] & g[30418];
assign g[46803] = a[14] & g[30419];
assign g[63186] = b[14] & g[30419];
assign g[46804] = a[14] & g[30420];
assign g[63187] = b[14] & g[30420];
assign g[46805] = a[14] & g[30421];
assign g[63188] = b[14] & g[30421];
assign g[46806] = a[14] & g[30422];
assign g[63189] = b[14] & g[30422];
assign g[46807] = a[14] & g[30423];
assign g[63190] = b[14] & g[30423];
assign g[46808] = a[14] & g[30424];
assign g[63191] = b[14] & g[30424];
assign g[46809] = a[14] & g[30425];
assign g[63192] = b[14] & g[30425];
assign g[46810] = a[14] & g[30426];
assign g[63193] = b[14] & g[30426];
assign g[46811] = a[14] & g[30427];
assign g[63194] = b[14] & g[30427];
assign g[46812] = a[14] & g[30428];
assign g[63195] = b[14] & g[30428];
assign g[46813] = a[14] & g[30429];
assign g[63196] = b[14] & g[30429];
assign g[46814] = a[14] & g[30430];
assign g[63197] = b[14] & g[30430];
assign g[46815] = a[14] & g[30431];
assign g[63198] = b[14] & g[30431];
assign g[46816] = a[14] & g[30432];
assign g[63199] = b[14] & g[30432];
assign g[46817] = a[14] & g[30433];
assign g[63200] = b[14] & g[30433];
assign g[46818] = a[14] & g[30434];
assign g[63201] = b[14] & g[30434];
assign g[46819] = a[14] & g[30435];
assign g[63202] = b[14] & g[30435];
assign g[46820] = a[14] & g[30436];
assign g[63203] = b[14] & g[30436];
assign g[46821] = a[14] & g[30437];
assign g[63204] = b[14] & g[30437];
assign g[46822] = a[14] & g[30438];
assign g[63205] = b[14] & g[30438];
assign g[46823] = a[14] & g[30439];
assign g[63206] = b[14] & g[30439];
assign g[46824] = a[14] & g[30440];
assign g[63207] = b[14] & g[30440];
assign g[46825] = a[14] & g[30441];
assign g[63208] = b[14] & g[30441];
assign g[46826] = a[14] & g[30442];
assign g[63209] = b[14] & g[30442];
assign g[46827] = a[14] & g[30443];
assign g[63210] = b[14] & g[30443];
assign g[46828] = a[14] & g[30444];
assign g[63211] = b[14] & g[30444];
assign g[46829] = a[14] & g[30445];
assign g[63212] = b[14] & g[30445];
assign g[46830] = a[14] & g[30446];
assign g[63213] = b[14] & g[30446];
assign g[46831] = a[14] & g[30447];
assign g[63214] = b[14] & g[30447];
assign g[46832] = a[14] & g[30448];
assign g[63215] = b[14] & g[30448];
assign g[46833] = a[14] & g[30449];
assign g[63216] = b[14] & g[30449];
assign g[46834] = a[14] & g[30450];
assign g[63217] = b[14] & g[30450];
assign g[46835] = a[14] & g[30451];
assign g[63218] = b[14] & g[30451];
assign g[46836] = a[14] & g[30452];
assign g[63219] = b[14] & g[30452];
assign g[46837] = a[14] & g[30453];
assign g[63220] = b[14] & g[30453];
assign g[46838] = a[14] & g[30454];
assign g[63221] = b[14] & g[30454];
assign g[46839] = a[14] & g[30455];
assign g[63222] = b[14] & g[30455];
assign g[46840] = a[14] & g[30456];
assign g[63223] = b[14] & g[30456];
assign g[46841] = a[14] & g[30457];
assign g[63224] = b[14] & g[30457];
assign g[46842] = a[14] & g[30458];
assign g[63225] = b[14] & g[30458];
assign g[46843] = a[14] & g[30459];
assign g[63226] = b[14] & g[30459];
assign g[46844] = a[14] & g[30460];
assign g[63227] = b[14] & g[30460];
assign g[46845] = a[14] & g[30461];
assign g[63228] = b[14] & g[30461];
assign g[46846] = a[14] & g[30462];
assign g[63229] = b[14] & g[30462];
assign g[46847] = a[14] & g[30463];
assign g[63230] = b[14] & g[30463];
assign g[46848] = a[14] & g[30464];
assign g[63231] = b[14] & g[30464];
assign g[46849] = a[14] & g[30465];
assign g[63232] = b[14] & g[30465];
assign g[46850] = a[14] & g[30466];
assign g[63233] = b[14] & g[30466];
assign g[46851] = a[14] & g[30467];
assign g[63234] = b[14] & g[30467];
assign g[46852] = a[14] & g[30468];
assign g[63235] = b[14] & g[30468];
assign g[46853] = a[14] & g[30469];
assign g[63236] = b[14] & g[30469];
assign g[46854] = a[14] & g[30470];
assign g[63237] = b[14] & g[30470];
assign g[46855] = a[14] & g[30471];
assign g[63238] = b[14] & g[30471];
assign g[46856] = a[14] & g[30472];
assign g[63239] = b[14] & g[30472];
assign g[46857] = a[14] & g[30473];
assign g[63240] = b[14] & g[30473];
assign g[46858] = a[14] & g[30474];
assign g[63241] = b[14] & g[30474];
assign g[46859] = a[14] & g[30475];
assign g[63242] = b[14] & g[30475];
assign g[46860] = a[14] & g[30476];
assign g[63243] = b[14] & g[30476];
assign g[46861] = a[14] & g[30477];
assign g[63244] = b[14] & g[30477];
assign g[46862] = a[14] & g[30478];
assign g[63245] = b[14] & g[30478];
assign g[46863] = a[14] & g[30479];
assign g[63246] = b[14] & g[30479];
assign g[46864] = a[14] & g[30480];
assign g[63247] = b[14] & g[30480];
assign g[46865] = a[14] & g[30481];
assign g[63248] = b[14] & g[30481];
assign g[46866] = a[14] & g[30482];
assign g[63249] = b[14] & g[30482];
assign g[46867] = a[14] & g[30483];
assign g[63250] = b[14] & g[30483];
assign g[46868] = a[14] & g[30484];
assign g[63251] = b[14] & g[30484];
assign g[46869] = a[14] & g[30485];
assign g[63252] = b[14] & g[30485];
assign g[46870] = a[14] & g[30486];
assign g[63253] = b[14] & g[30486];
assign g[46871] = a[14] & g[30487];
assign g[63254] = b[14] & g[30487];
assign g[46872] = a[14] & g[30488];
assign g[63255] = b[14] & g[30488];
assign g[46873] = a[14] & g[30489];
assign g[63256] = b[14] & g[30489];
assign g[46874] = a[14] & g[30490];
assign g[63257] = b[14] & g[30490];
assign g[46875] = a[14] & g[30491];
assign g[63258] = b[14] & g[30491];
assign g[46876] = a[14] & g[30492];
assign g[63259] = b[14] & g[30492];
assign g[46877] = a[14] & g[30493];
assign g[63260] = b[14] & g[30493];
assign g[46878] = a[14] & g[30494];
assign g[63261] = b[14] & g[30494];
assign g[46879] = a[14] & g[30495];
assign g[63262] = b[14] & g[30495];
assign g[46880] = a[14] & g[30496];
assign g[63263] = b[14] & g[30496];
assign g[46881] = a[14] & g[30497];
assign g[63264] = b[14] & g[30497];
assign g[46882] = a[14] & g[30498];
assign g[63265] = b[14] & g[30498];
assign g[46883] = a[14] & g[30499];
assign g[63266] = b[14] & g[30499];
assign g[46884] = a[14] & g[30500];
assign g[63267] = b[14] & g[30500];
assign g[46885] = a[14] & g[30501];
assign g[63268] = b[14] & g[30501];
assign g[46886] = a[14] & g[30502];
assign g[63269] = b[14] & g[30502];
assign g[46887] = a[14] & g[30503];
assign g[63270] = b[14] & g[30503];
assign g[46888] = a[14] & g[30504];
assign g[63271] = b[14] & g[30504];
assign g[46889] = a[14] & g[30505];
assign g[63272] = b[14] & g[30505];
assign g[46890] = a[14] & g[30506];
assign g[63273] = b[14] & g[30506];
assign g[46891] = a[14] & g[30507];
assign g[63274] = b[14] & g[30507];
assign g[46892] = a[14] & g[30508];
assign g[63275] = b[14] & g[30508];
assign g[46893] = a[14] & g[30509];
assign g[63276] = b[14] & g[30509];
assign g[46894] = a[14] & g[30510];
assign g[63277] = b[14] & g[30510];
assign g[46895] = a[14] & g[30511];
assign g[63278] = b[14] & g[30511];
assign g[46896] = a[14] & g[30512];
assign g[63279] = b[14] & g[30512];
assign g[46897] = a[14] & g[30513];
assign g[63280] = b[14] & g[30513];
assign g[46898] = a[14] & g[30514];
assign g[63281] = b[14] & g[30514];
assign g[46899] = a[14] & g[30515];
assign g[63282] = b[14] & g[30515];
assign g[46900] = a[14] & g[30516];
assign g[63283] = b[14] & g[30516];
assign g[46901] = a[14] & g[30517];
assign g[63284] = b[14] & g[30517];
assign g[46902] = a[14] & g[30518];
assign g[63285] = b[14] & g[30518];
assign g[46903] = a[14] & g[30519];
assign g[63286] = b[14] & g[30519];
assign g[46904] = a[14] & g[30520];
assign g[63287] = b[14] & g[30520];
assign g[46905] = a[14] & g[30521];
assign g[63288] = b[14] & g[30521];
assign g[46906] = a[14] & g[30522];
assign g[63289] = b[14] & g[30522];
assign g[46907] = a[14] & g[30523];
assign g[63290] = b[14] & g[30523];
assign g[46908] = a[14] & g[30524];
assign g[63291] = b[14] & g[30524];
assign g[46909] = a[14] & g[30525];
assign g[63292] = b[14] & g[30525];
assign g[46910] = a[14] & g[30526];
assign g[63293] = b[14] & g[30526];
assign g[46911] = a[14] & g[30527];
assign g[63294] = b[14] & g[30527];
assign g[46912] = a[14] & g[30528];
assign g[63295] = b[14] & g[30528];
assign g[46913] = a[14] & g[30529];
assign g[63296] = b[14] & g[30529];
assign g[46914] = a[14] & g[30530];
assign g[63297] = b[14] & g[30530];
assign g[46915] = a[14] & g[30531];
assign g[63298] = b[14] & g[30531];
assign g[46916] = a[14] & g[30532];
assign g[63299] = b[14] & g[30532];
assign g[46917] = a[14] & g[30533];
assign g[63300] = b[14] & g[30533];
assign g[46918] = a[14] & g[30534];
assign g[63301] = b[14] & g[30534];
assign g[46919] = a[14] & g[30535];
assign g[63302] = b[14] & g[30535];
assign g[46920] = a[14] & g[30536];
assign g[63303] = b[14] & g[30536];
assign g[46921] = a[14] & g[30537];
assign g[63304] = b[14] & g[30537];
assign g[46922] = a[14] & g[30538];
assign g[63305] = b[14] & g[30538];
assign g[46923] = a[14] & g[30539];
assign g[63306] = b[14] & g[30539];
assign g[46924] = a[14] & g[30540];
assign g[63307] = b[14] & g[30540];
assign g[46925] = a[14] & g[30541];
assign g[63308] = b[14] & g[30541];
assign g[46926] = a[14] & g[30542];
assign g[63309] = b[14] & g[30542];
assign g[46927] = a[14] & g[30543];
assign g[63310] = b[14] & g[30543];
assign g[46928] = a[14] & g[30544];
assign g[63311] = b[14] & g[30544];
assign g[46929] = a[14] & g[30545];
assign g[63312] = b[14] & g[30545];
assign g[46930] = a[14] & g[30546];
assign g[63313] = b[14] & g[30546];
assign g[46931] = a[14] & g[30547];
assign g[63314] = b[14] & g[30547];
assign g[46932] = a[14] & g[30548];
assign g[63315] = b[14] & g[30548];
assign g[46933] = a[14] & g[30549];
assign g[63316] = b[14] & g[30549];
assign g[46934] = a[14] & g[30550];
assign g[63317] = b[14] & g[30550];
assign g[46935] = a[14] & g[30551];
assign g[63318] = b[14] & g[30551];
assign g[46936] = a[14] & g[30552];
assign g[63319] = b[14] & g[30552];
assign g[46937] = a[14] & g[30553];
assign g[63320] = b[14] & g[30553];
assign g[46938] = a[14] & g[30554];
assign g[63321] = b[14] & g[30554];
assign g[46939] = a[14] & g[30555];
assign g[63322] = b[14] & g[30555];
assign g[46940] = a[14] & g[30556];
assign g[63323] = b[14] & g[30556];
assign g[46941] = a[14] & g[30557];
assign g[63324] = b[14] & g[30557];
assign g[46942] = a[14] & g[30558];
assign g[63325] = b[14] & g[30558];
assign g[46943] = a[14] & g[30559];
assign g[63326] = b[14] & g[30559];
assign g[46944] = a[14] & g[30560];
assign g[63327] = b[14] & g[30560];
assign g[46945] = a[14] & g[30561];
assign g[63328] = b[14] & g[30561];
assign g[46946] = a[14] & g[30562];
assign g[63329] = b[14] & g[30562];
assign g[46947] = a[14] & g[30563];
assign g[63330] = b[14] & g[30563];
assign g[46948] = a[14] & g[30564];
assign g[63331] = b[14] & g[30564];
assign g[46949] = a[14] & g[30565];
assign g[63332] = b[14] & g[30565];
assign g[46950] = a[14] & g[30566];
assign g[63333] = b[14] & g[30566];
assign g[46951] = a[14] & g[30567];
assign g[63334] = b[14] & g[30567];
assign g[46952] = a[14] & g[30568];
assign g[63335] = b[14] & g[30568];
assign g[46953] = a[14] & g[30569];
assign g[63336] = b[14] & g[30569];
assign g[46954] = a[14] & g[30570];
assign g[63337] = b[14] & g[30570];
assign g[46955] = a[14] & g[30571];
assign g[63338] = b[14] & g[30571];
assign g[46956] = a[14] & g[30572];
assign g[63339] = b[14] & g[30572];
assign g[46957] = a[14] & g[30573];
assign g[63340] = b[14] & g[30573];
assign g[46958] = a[14] & g[30574];
assign g[63341] = b[14] & g[30574];
assign g[46959] = a[14] & g[30575];
assign g[63342] = b[14] & g[30575];
assign g[46960] = a[14] & g[30576];
assign g[63343] = b[14] & g[30576];
assign g[46961] = a[14] & g[30577];
assign g[63344] = b[14] & g[30577];
assign g[46962] = a[14] & g[30578];
assign g[63345] = b[14] & g[30578];
assign g[46963] = a[14] & g[30579];
assign g[63346] = b[14] & g[30579];
assign g[46964] = a[14] & g[30580];
assign g[63347] = b[14] & g[30580];
assign g[46965] = a[14] & g[30581];
assign g[63348] = b[14] & g[30581];
assign g[46966] = a[14] & g[30582];
assign g[63349] = b[14] & g[30582];
assign g[46967] = a[14] & g[30583];
assign g[63350] = b[14] & g[30583];
assign g[46968] = a[14] & g[30584];
assign g[63351] = b[14] & g[30584];
assign g[46969] = a[14] & g[30585];
assign g[63352] = b[14] & g[30585];
assign g[46970] = a[14] & g[30586];
assign g[63353] = b[14] & g[30586];
assign g[46971] = a[14] & g[30587];
assign g[63354] = b[14] & g[30587];
assign g[46972] = a[14] & g[30588];
assign g[63355] = b[14] & g[30588];
assign g[46973] = a[14] & g[30589];
assign g[63356] = b[14] & g[30589];
assign g[46974] = a[14] & g[30590];
assign g[63357] = b[14] & g[30590];
assign g[46975] = a[14] & g[30591];
assign g[63358] = b[14] & g[30591];
assign g[46976] = a[14] & g[30592];
assign g[63359] = b[14] & g[30592];
assign g[46977] = a[14] & g[30593];
assign g[63360] = b[14] & g[30593];
assign g[46978] = a[14] & g[30594];
assign g[63361] = b[14] & g[30594];
assign g[46979] = a[14] & g[30595];
assign g[63362] = b[14] & g[30595];
assign g[46980] = a[14] & g[30596];
assign g[63363] = b[14] & g[30596];
assign g[46981] = a[14] & g[30597];
assign g[63364] = b[14] & g[30597];
assign g[46982] = a[14] & g[30598];
assign g[63365] = b[14] & g[30598];
assign g[46983] = a[14] & g[30599];
assign g[63366] = b[14] & g[30599];
assign g[46984] = a[14] & g[30600];
assign g[63367] = b[14] & g[30600];
assign g[46985] = a[14] & g[30601];
assign g[63368] = b[14] & g[30601];
assign g[46986] = a[14] & g[30602];
assign g[63369] = b[14] & g[30602];
assign g[46987] = a[14] & g[30603];
assign g[63370] = b[14] & g[30603];
assign g[46988] = a[14] & g[30604];
assign g[63371] = b[14] & g[30604];
assign g[46989] = a[14] & g[30605];
assign g[63372] = b[14] & g[30605];
assign g[46990] = a[14] & g[30606];
assign g[63373] = b[14] & g[30606];
assign g[46991] = a[14] & g[30607];
assign g[63374] = b[14] & g[30607];
assign g[46992] = a[14] & g[30608];
assign g[63375] = b[14] & g[30608];
assign g[46993] = a[14] & g[30609];
assign g[63376] = b[14] & g[30609];
assign g[46994] = a[14] & g[30610];
assign g[63377] = b[14] & g[30610];
assign g[46995] = a[14] & g[30611];
assign g[63378] = b[14] & g[30611];
assign g[46996] = a[14] & g[30612];
assign g[63379] = b[14] & g[30612];
assign g[46997] = a[14] & g[30613];
assign g[63380] = b[14] & g[30613];
assign g[46998] = a[14] & g[30614];
assign g[63381] = b[14] & g[30614];
assign g[46999] = a[14] & g[30615];
assign g[63382] = b[14] & g[30615];
assign g[47000] = a[14] & g[30616];
assign g[63383] = b[14] & g[30616];
assign g[47001] = a[14] & g[30617];
assign g[63384] = b[14] & g[30617];
assign g[47002] = a[14] & g[30618];
assign g[63385] = b[14] & g[30618];
assign g[47003] = a[14] & g[30619];
assign g[63386] = b[14] & g[30619];
assign g[47004] = a[14] & g[30620];
assign g[63387] = b[14] & g[30620];
assign g[47005] = a[14] & g[30621];
assign g[63388] = b[14] & g[30621];
assign g[47006] = a[14] & g[30622];
assign g[63389] = b[14] & g[30622];
assign g[47007] = a[14] & g[30623];
assign g[63390] = b[14] & g[30623];
assign g[47008] = a[14] & g[30624];
assign g[63391] = b[14] & g[30624];
assign g[47009] = a[14] & g[30625];
assign g[63392] = b[14] & g[30625];
assign g[47010] = a[14] & g[30626];
assign g[63393] = b[14] & g[30626];
assign g[47011] = a[14] & g[30627];
assign g[63394] = b[14] & g[30627];
assign g[47012] = a[14] & g[30628];
assign g[63395] = b[14] & g[30628];
assign g[47013] = a[14] & g[30629];
assign g[63396] = b[14] & g[30629];
assign g[47014] = a[14] & g[30630];
assign g[63397] = b[14] & g[30630];
assign g[47015] = a[14] & g[30631];
assign g[63398] = b[14] & g[30631];
assign g[47016] = a[14] & g[30632];
assign g[63399] = b[14] & g[30632];
assign g[47017] = a[14] & g[30633];
assign g[63400] = b[14] & g[30633];
assign g[47018] = a[14] & g[30634];
assign g[63401] = b[14] & g[30634];
assign g[47019] = a[14] & g[30635];
assign g[63402] = b[14] & g[30635];
assign g[47020] = a[14] & g[30636];
assign g[63403] = b[14] & g[30636];
assign g[47021] = a[14] & g[30637];
assign g[63404] = b[14] & g[30637];
assign g[47022] = a[14] & g[30638];
assign g[63405] = b[14] & g[30638];
assign g[47023] = a[14] & g[30639];
assign g[63406] = b[14] & g[30639];
assign g[47024] = a[14] & g[30640];
assign g[63407] = b[14] & g[30640];
assign g[47025] = a[14] & g[30641];
assign g[63408] = b[14] & g[30641];
assign g[47026] = a[14] & g[30642];
assign g[63409] = b[14] & g[30642];
assign g[47027] = a[14] & g[30643];
assign g[63410] = b[14] & g[30643];
assign g[47028] = a[14] & g[30644];
assign g[63411] = b[14] & g[30644];
assign g[47029] = a[14] & g[30645];
assign g[63412] = b[14] & g[30645];
assign g[47030] = a[14] & g[30646];
assign g[63413] = b[14] & g[30646];
assign g[47031] = a[14] & g[30647];
assign g[63414] = b[14] & g[30647];
assign g[47032] = a[14] & g[30648];
assign g[63415] = b[14] & g[30648];
assign g[47033] = a[14] & g[30649];
assign g[63416] = b[14] & g[30649];
assign g[47034] = a[14] & g[30650];
assign g[63417] = b[14] & g[30650];
assign g[47035] = a[14] & g[30651];
assign g[63418] = b[14] & g[30651];
assign g[47036] = a[14] & g[30652];
assign g[63419] = b[14] & g[30652];
assign g[47037] = a[14] & g[30653];
assign g[63420] = b[14] & g[30653];
assign g[47038] = a[14] & g[30654];
assign g[63421] = b[14] & g[30654];
assign g[47039] = a[14] & g[30655];
assign g[63422] = b[14] & g[30655];
assign g[47040] = a[14] & g[30656];
assign g[63423] = b[14] & g[30656];
assign g[47041] = a[14] & g[30657];
assign g[63424] = b[14] & g[30657];
assign g[47042] = a[14] & g[30658];
assign g[63425] = b[14] & g[30658];
assign g[47043] = a[14] & g[30659];
assign g[63426] = b[14] & g[30659];
assign g[47044] = a[14] & g[30660];
assign g[63427] = b[14] & g[30660];
assign g[47045] = a[14] & g[30661];
assign g[63428] = b[14] & g[30661];
assign g[47046] = a[14] & g[30662];
assign g[63429] = b[14] & g[30662];
assign g[47047] = a[14] & g[30663];
assign g[63430] = b[14] & g[30663];
assign g[47048] = a[14] & g[30664];
assign g[63431] = b[14] & g[30664];
assign g[47049] = a[14] & g[30665];
assign g[63432] = b[14] & g[30665];
assign g[47050] = a[14] & g[30666];
assign g[63433] = b[14] & g[30666];
assign g[47051] = a[14] & g[30667];
assign g[63434] = b[14] & g[30667];
assign g[47052] = a[14] & g[30668];
assign g[63435] = b[14] & g[30668];
assign g[47053] = a[14] & g[30669];
assign g[63436] = b[14] & g[30669];
assign g[47054] = a[14] & g[30670];
assign g[63437] = b[14] & g[30670];
assign g[47055] = a[14] & g[30671];
assign g[63438] = b[14] & g[30671];
assign g[47056] = a[14] & g[30672];
assign g[63439] = b[14] & g[30672];
assign g[47057] = a[14] & g[30673];
assign g[63440] = b[14] & g[30673];
assign g[47058] = a[14] & g[30674];
assign g[63441] = b[14] & g[30674];
assign g[47059] = a[14] & g[30675];
assign g[63442] = b[14] & g[30675];
assign g[47060] = a[14] & g[30676];
assign g[63443] = b[14] & g[30676];
assign g[47061] = a[14] & g[30677];
assign g[63444] = b[14] & g[30677];
assign g[47062] = a[14] & g[30678];
assign g[63445] = b[14] & g[30678];
assign g[47063] = a[14] & g[30679];
assign g[63446] = b[14] & g[30679];
assign g[47064] = a[14] & g[30680];
assign g[63447] = b[14] & g[30680];
assign g[47065] = a[14] & g[30681];
assign g[63448] = b[14] & g[30681];
assign g[47066] = a[14] & g[30682];
assign g[63449] = b[14] & g[30682];
assign g[47067] = a[14] & g[30683];
assign g[63450] = b[14] & g[30683];
assign g[47068] = a[14] & g[30684];
assign g[63451] = b[14] & g[30684];
assign g[47069] = a[14] & g[30685];
assign g[63452] = b[14] & g[30685];
assign g[47070] = a[14] & g[30686];
assign g[63453] = b[14] & g[30686];
assign g[47071] = a[14] & g[30687];
assign g[63454] = b[14] & g[30687];
assign g[47072] = a[14] & g[30688];
assign g[63455] = b[14] & g[30688];
assign g[47073] = a[14] & g[30689];
assign g[63456] = b[14] & g[30689];
assign g[47074] = a[14] & g[30690];
assign g[63457] = b[14] & g[30690];
assign g[47075] = a[14] & g[30691];
assign g[63458] = b[14] & g[30691];
assign g[47076] = a[14] & g[30692];
assign g[63459] = b[14] & g[30692];
assign g[47077] = a[14] & g[30693];
assign g[63460] = b[14] & g[30693];
assign g[47078] = a[14] & g[30694];
assign g[63461] = b[14] & g[30694];
assign g[47079] = a[14] & g[30695];
assign g[63462] = b[14] & g[30695];
assign g[47080] = a[14] & g[30696];
assign g[63463] = b[14] & g[30696];
assign g[47081] = a[14] & g[30697];
assign g[63464] = b[14] & g[30697];
assign g[47082] = a[14] & g[30698];
assign g[63465] = b[14] & g[30698];
assign g[47083] = a[14] & g[30699];
assign g[63466] = b[14] & g[30699];
assign g[47084] = a[14] & g[30700];
assign g[63467] = b[14] & g[30700];
assign g[47085] = a[14] & g[30701];
assign g[63468] = b[14] & g[30701];
assign g[47086] = a[14] & g[30702];
assign g[63469] = b[14] & g[30702];
assign g[47087] = a[14] & g[30703];
assign g[63470] = b[14] & g[30703];
assign g[47088] = a[14] & g[30704];
assign g[63471] = b[14] & g[30704];
assign g[47089] = a[14] & g[30705];
assign g[63472] = b[14] & g[30705];
assign g[47090] = a[14] & g[30706];
assign g[63473] = b[14] & g[30706];
assign g[47091] = a[14] & g[30707];
assign g[63474] = b[14] & g[30707];
assign g[47092] = a[14] & g[30708];
assign g[63475] = b[14] & g[30708];
assign g[47093] = a[14] & g[30709];
assign g[63476] = b[14] & g[30709];
assign g[47094] = a[14] & g[30710];
assign g[63477] = b[14] & g[30710];
assign g[47095] = a[14] & g[30711];
assign g[63478] = b[14] & g[30711];
assign g[47096] = a[14] & g[30712];
assign g[63479] = b[14] & g[30712];
assign g[47097] = a[14] & g[30713];
assign g[63480] = b[14] & g[30713];
assign g[47098] = a[14] & g[30714];
assign g[63481] = b[14] & g[30714];
assign g[47099] = a[14] & g[30715];
assign g[63482] = b[14] & g[30715];
assign g[47100] = a[14] & g[30716];
assign g[63483] = b[14] & g[30716];
assign g[47101] = a[14] & g[30717];
assign g[63484] = b[14] & g[30717];
assign g[47102] = a[14] & g[30718];
assign g[63485] = b[14] & g[30718];
assign g[47103] = a[14] & g[30719];
assign g[63486] = b[14] & g[30719];
assign g[47104] = a[14] & g[30720];
assign g[63487] = b[14] & g[30720];
assign g[47105] = a[14] & g[30721];
assign g[63488] = b[14] & g[30721];
assign g[47106] = a[14] & g[30722];
assign g[63489] = b[14] & g[30722];
assign g[47107] = a[14] & g[30723];
assign g[63490] = b[14] & g[30723];
assign g[47108] = a[14] & g[30724];
assign g[63491] = b[14] & g[30724];
assign g[47109] = a[14] & g[30725];
assign g[63492] = b[14] & g[30725];
assign g[47110] = a[14] & g[30726];
assign g[63493] = b[14] & g[30726];
assign g[47111] = a[14] & g[30727];
assign g[63494] = b[14] & g[30727];
assign g[47112] = a[14] & g[30728];
assign g[63495] = b[14] & g[30728];
assign g[47113] = a[14] & g[30729];
assign g[63496] = b[14] & g[30729];
assign g[47114] = a[14] & g[30730];
assign g[63497] = b[14] & g[30730];
assign g[47115] = a[14] & g[30731];
assign g[63498] = b[14] & g[30731];
assign g[47116] = a[14] & g[30732];
assign g[63499] = b[14] & g[30732];
assign g[47117] = a[14] & g[30733];
assign g[63500] = b[14] & g[30733];
assign g[47118] = a[14] & g[30734];
assign g[63501] = b[14] & g[30734];
assign g[47119] = a[14] & g[30735];
assign g[63502] = b[14] & g[30735];
assign g[47120] = a[14] & g[30736];
assign g[63503] = b[14] & g[30736];
assign g[47121] = a[14] & g[30737];
assign g[63504] = b[14] & g[30737];
assign g[47122] = a[14] & g[30738];
assign g[63505] = b[14] & g[30738];
assign g[47123] = a[14] & g[30739];
assign g[63506] = b[14] & g[30739];
assign g[47124] = a[14] & g[30740];
assign g[63507] = b[14] & g[30740];
assign g[47125] = a[14] & g[30741];
assign g[63508] = b[14] & g[30741];
assign g[47126] = a[14] & g[30742];
assign g[63509] = b[14] & g[30742];
assign g[47127] = a[14] & g[30743];
assign g[63510] = b[14] & g[30743];
assign g[47128] = a[14] & g[30744];
assign g[63511] = b[14] & g[30744];
assign g[47129] = a[14] & g[30745];
assign g[63512] = b[14] & g[30745];
assign g[47130] = a[14] & g[30746];
assign g[63513] = b[14] & g[30746];
assign g[47131] = a[14] & g[30747];
assign g[63514] = b[14] & g[30747];
assign g[47132] = a[14] & g[30748];
assign g[63515] = b[14] & g[30748];
assign g[47133] = a[14] & g[30749];
assign g[63516] = b[14] & g[30749];
assign g[47134] = a[14] & g[30750];
assign g[63517] = b[14] & g[30750];
assign g[47135] = a[14] & g[30751];
assign g[63518] = b[14] & g[30751];
assign g[47136] = a[14] & g[30752];
assign g[63519] = b[14] & g[30752];
assign g[47137] = a[14] & g[30753];
assign g[63520] = b[14] & g[30753];
assign g[47138] = a[14] & g[30754];
assign g[63521] = b[14] & g[30754];
assign g[47139] = a[14] & g[30755];
assign g[63522] = b[14] & g[30755];
assign g[47140] = a[14] & g[30756];
assign g[63523] = b[14] & g[30756];
assign g[47141] = a[14] & g[30757];
assign g[63524] = b[14] & g[30757];
assign g[47142] = a[14] & g[30758];
assign g[63525] = b[14] & g[30758];
assign g[47143] = a[14] & g[30759];
assign g[63526] = b[14] & g[30759];
assign g[47144] = a[14] & g[30760];
assign g[63527] = b[14] & g[30760];
assign g[47145] = a[14] & g[30761];
assign g[63528] = b[14] & g[30761];
assign g[47146] = a[14] & g[30762];
assign g[63529] = b[14] & g[30762];
assign g[47147] = a[14] & g[30763];
assign g[63530] = b[14] & g[30763];
assign g[47148] = a[14] & g[30764];
assign g[63531] = b[14] & g[30764];
assign g[47149] = a[14] & g[30765];
assign g[63532] = b[14] & g[30765];
assign g[47150] = a[14] & g[30766];
assign g[63533] = b[14] & g[30766];
assign g[47151] = a[14] & g[30767];
assign g[63534] = b[14] & g[30767];
assign g[47152] = a[14] & g[30768];
assign g[63535] = b[14] & g[30768];
assign g[47153] = a[14] & g[30769];
assign g[63536] = b[14] & g[30769];
assign g[47154] = a[14] & g[30770];
assign g[63537] = b[14] & g[30770];
assign g[47155] = a[14] & g[30771];
assign g[63538] = b[14] & g[30771];
assign g[47156] = a[14] & g[30772];
assign g[63539] = b[14] & g[30772];
assign g[47157] = a[14] & g[30773];
assign g[63540] = b[14] & g[30773];
assign g[47158] = a[14] & g[30774];
assign g[63541] = b[14] & g[30774];
assign g[47159] = a[14] & g[30775];
assign g[63542] = b[14] & g[30775];
assign g[47160] = a[14] & g[30776];
assign g[63543] = b[14] & g[30776];
assign g[47161] = a[14] & g[30777];
assign g[63544] = b[14] & g[30777];
assign g[47162] = a[14] & g[30778];
assign g[63545] = b[14] & g[30778];
assign g[47163] = a[14] & g[30779];
assign g[63546] = b[14] & g[30779];
assign g[47164] = a[14] & g[30780];
assign g[63547] = b[14] & g[30780];
assign g[47165] = a[14] & g[30781];
assign g[63548] = b[14] & g[30781];
assign g[47166] = a[14] & g[30782];
assign g[63549] = b[14] & g[30782];
assign g[47167] = a[14] & g[30783];
assign g[63550] = b[14] & g[30783];
assign g[47168] = a[14] & g[30784];
assign g[63551] = b[14] & g[30784];
assign g[47169] = a[14] & g[30785];
assign g[63552] = b[14] & g[30785];
assign g[47170] = a[14] & g[30786];
assign g[63553] = b[14] & g[30786];
assign g[47171] = a[14] & g[30787];
assign g[63554] = b[14] & g[30787];
assign g[47172] = a[14] & g[30788];
assign g[63555] = b[14] & g[30788];
assign g[47173] = a[14] & g[30789];
assign g[63556] = b[14] & g[30789];
assign g[47174] = a[14] & g[30790];
assign g[63557] = b[14] & g[30790];
assign g[47175] = a[14] & g[30791];
assign g[63558] = b[14] & g[30791];
assign g[47176] = a[14] & g[30792];
assign g[63559] = b[14] & g[30792];
assign g[47177] = a[14] & g[30793];
assign g[63560] = b[14] & g[30793];
assign g[47178] = a[14] & g[30794];
assign g[63561] = b[14] & g[30794];
assign g[47179] = a[14] & g[30795];
assign g[63562] = b[14] & g[30795];
assign g[47180] = a[14] & g[30796];
assign g[63563] = b[14] & g[30796];
assign g[47181] = a[14] & g[30797];
assign g[63564] = b[14] & g[30797];
assign g[47182] = a[14] & g[30798];
assign g[63565] = b[14] & g[30798];
assign g[47183] = a[14] & g[30799];
assign g[63566] = b[14] & g[30799];
assign g[47184] = a[14] & g[30800];
assign g[63567] = b[14] & g[30800];
assign g[47185] = a[14] & g[30801];
assign g[63568] = b[14] & g[30801];
assign g[47186] = a[14] & g[30802];
assign g[63569] = b[14] & g[30802];
assign g[47187] = a[14] & g[30803];
assign g[63570] = b[14] & g[30803];
assign g[47188] = a[14] & g[30804];
assign g[63571] = b[14] & g[30804];
assign g[47189] = a[14] & g[30805];
assign g[63572] = b[14] & g[30805];
assign g[47190] = a[14] & g[30806];
assign g[63573] = b[14] & g[30806];
assign g[47191] = a[14] & g[30807];
assign g[63574] = b[14] & g[30807];
assign g[47192] = a[14] & g[30808];
assign g[63575] = b[14] & g[30808];
assign g[47193] = a[14] & g[30809];
assign g[63576] = b[14] & g[30809];
assign g[47194] = a[14] & g[30810];
assign g[63577] = b[14] & g[30810];
assign g[47195] = a[14] & g[30811];
assign g[63578] = b[14] & g[30811];
assign g[47196] = a[14] & g[30812];
assign g[63579] = b[14] & g[30812];
assign g[47197] = a[14] & g[30813];
assign g[63580] = b[14] & g[30813];
assign g[47198] = a[14] & g[30814];
assign g[63581] = b[14] & g[30814];
assign g[47199] = a[14] & g[30815];
assign g[63582] = b[14] & g[30815];
assign g[47200] = a[14] & g[30816];
assign g[63583] = b[14] & g[30816];
assign g[47201] = a[14] & g[30817];
assign g[63584] = b[14] & g[30817];
assign g[47202] = a[14] & g[30818];
assign g[63585] = b[14] & g[30818];
assign g[47203] = a[14] & g[30819];
assign g[63586] = b[14] & g[30819];
assign g[47204] = a[14] & g[30820];
assign g[63587] = b[14] & g[30820];
assign g[47205] = a[14] & g[30821];
assign g[63588] = b[14] & g[30821];
assign g[47206] = a[14] & g[30822];
assign g[63589] = b[14] & g[30822];
assign g[47207] = a[14] & g[30823];
assign g[63590] = b[14] & g[30823];
assign g[47208] = a[14] & g[30824];
assign g[63591] = b[14] & g[30824];
assign g[47209] = a[14] & g[30825];
assign g[63592] = b[14] & g[30825];
assign g[47210] = a[14] & g[30826];
assign g[63593] = b[14] & g[30826];
assign g[47211] = a[14] & g[30827];
assign g[63594] = b[14] & g[30827];
assign g[47212] = a[14] & g[30828];
assign g[63595] = b[14] & g[30828];
assign g[47213] = a[14] & g[30829];
assign g[63596] = b[14] & g[30829];
assign g[47214] = a[14] & g[30830];
assign g[63597] = b[14] & g[30830];
assign g[47215] = a[14] & g[30831];
assign g[63598] = b[14] & g[30831];
assign g[47216] = a[14] & g[30832];
assign g[63599] = b[14] & g[30832];
assign g[47217] = a[14] & g[30833];
assign g[63600] = b[14] & g[30833];
assign g[47218] = a[14] & g[30834];
assign g[63601] = b[14] & g[30834];
assign g[47219] = a[14] & g[30835];
assign g[63602] = b[14] & g[30835];
assign g[47220] = a[14] & g[30836];
assign g[63603] = b[14] & g[30836];
assign g[47221] = a[14] & g[30837];
assign g[63604] = b[14] & g[30837];
assign g[47222] = a[14] & g[30838];
assign g[63605] = b[14] & g[30838];
assign g[47223] = a[14] & g[30839];
assign g[63606] = b[14] & g[30839];
assign g[47224] = a[14] & g[30840];
assign g[63607] = b[14] & g[30840];
assign g[47225] = a[14] & g[30841];
assign g[63608] = b[14] & g[30841];
assign g[47226] = a[14] & g[30842];
assign g[63609] = b[14] & g[30842];
assign g[47227] = a[14] & g[30843];
assign g[63610] = b[14] & g[30843];
assign g[47228] = a[14] & g[30844];
assign g[63611] = b[14] & g[30844];
assign g[47229] = a[14] & g[30845];
assign g[63612] = b[14] & g[30845];
assign g[47230] = a[14] & g[30846];
assign g[63613] = b[14] & g[30846];
assign g[47231] = a[14] & g[30847];
assign g[63614] = b[14] & g[30847];
assign g[47232] = a[14] & g[30848];
assign g[63615] = b[14] & g[30848];
assign g[47233] = a[14] & g[30849];
assign g[63616] = b[14] & g[30849];
assign g[47234] = a[14] & g[30850];
assign g[63617] = b[14] & g[30850];
assign g[47235] = a[14] & g[30851];
assign g[63618] = b[14] & g[30851];
assign g[47236] = a[14] & g[30852];
assign g[63619] = b[14] & g[30852];
assign g[47237] = a[14] & g[30853];
assign g[63620] = b[14] & g[30853];
assign g[47238] = a[14] & g[30854];
assign g[63621] = b[14] & g[30854];
assign g[47239] = a[14] & g[30855];
assign g[63622] = b[14] & g[30855];
assign g[47240] = a[14] & g[30856];
assign g[63623] = b[14] & g[30856];
assign g[47241] = a[14] & g[30857];
assign g[63624] = b[14] & g[30857];
assign g[47242] = a[14] & g[30858];
assign g[63625] = b[14] & g[30858];
assign g[47243] = a[14] & g[30859];
assign g[63626] = b[14] & g[30859];
assign g[47244] = a[14] & g[30860];
assign g[63627] = b[14] & g[30860];
assign g[47245] = a[14] & g[30861];
assign g[63628] = b[14] & g[30861];
assign g[47246] = a[14] & g[30862];
assign g[63629] = b[14] & g[30862];
assign g[47247] = a[14] & g[30863];
assign g[63630] = b[14] & g[30863];
assign g[47248] = a[14] & g[30864];
assign g[63631] = b[14] & g[30864];
assign g[47249] = a[14] & g[30865];
assign g[63632] = b[14] & g[30865];
assign g[47250] = a[14] & g[30866];
assign g[63633] = b[14] & g[30866];
assign g[47251] = a[14] & g[30867];
assign g[63634] = b[14] & g[30867];
assign g[47252] = a[14] & g[30868];
assign g[63635] = b[14] & g[30868];
assign g[47253] = a[14] & g[30869];
assign g[63636] = b[14] & g[30869];
assign g[47254] = a[14] & g[30870];
assign g[63637] = b[14] & g[30870];
assign g[47255] = a[14] & g[30871];
assign g[63638] = b[14] & g[30871];
assign g[47256] = a[14] & g[30872];
assign g[63639] = b[14] & g[30872];
assign g[47257] = a[14] & g[30873];
assign g[63640] = b[14] & g[30873];
assign g[47258] = a[14] & g[30874];
assign g[63641] = b[14] & g[30874];
assign g[47259] = a[14] & g[30875];
assign g[63642] = b[14] & g[30875];
assign g[47260] = a[14] & g[30876];
assign g[63643] = b[14] & g[30876];
assign g[47261] = a[14] & g[30877];
assign g[63644] = b[14] & g[30877];
assign g[47262] = a[14] & g[30878];
assign g[63645] = b[14] & g[30878];
assign g[47263] = a[14] & g[30879];
assign g[63646] = b[14] & g[30879];
assign g[47264] = a[14] & g[30880];
assign g[63647] = b[14] & g[30880];
assign g[47265] = a[14] & g[30881];
assign g[63648] = b[14] & g[30881];
assign g[47266] = a[14] & g[30882];
assign g[63649] = b[14] & g[30882];
assign g[47267] = a[14] & g[30883];
assign g[63650] = b[14] & g[30883];
assign g[47268] = a[14] & g[30884];
assign g[63651] = b[14] & g[30884];
assign g[47269] = a[14] & g[30885];
assign g[63652] = b[14] & g[30885];
assign g[47270] = a[14] & g[30886];
assign g[63653] = b[14] & g[30886];
assign g[47271] = a[14] & g[30887];
assign g[63654] = b[14] & g[30887];
assign g[47272] = a[14] & g[30888];
assign g[63655] = b[14] & g[30888];
assign g[47273] = a[14] & g[30889];
assign g[63656] = b[14] & g[30889];
assign g[47274] = a[14] & g[30890];
assign g[63657] = b[14] & g[30890];
assign g[47275] = a[14] & g[30891];
assign g[63658] = b[14] & g[30891];
assign g[47276] = a[14] & g[30892];
assign g[63659] = b[14] & g[30892];
assign g[47277] = a[14] & g[30893];
assign g[63660] = b[14] & g[30893];
assign g[47278] = a[14] & g[30894];
assign g[63661] = b[14] & g[30894];
assign g[47279] = a[14] & g[30895];
assign g[63662] = b[14] & g[30895];
assign g[47280] = a[14] & g[30896];
assign g[63663] = b[14] & g[30896];
assign g[47281] = a[14] & g[30897];
assign g[63664] = b[14] & g[30897];
assign g[47282] = a[14] & g[30898];
assign g[63665] = b[14] & g[30898];
assign g[47283] = a[14] & g[30899];
assign g[63666] = b[14] & g[30899];
assign g[47284] = a[14] & g[30900];
assign g[63667] = b[14] & g[30900];
assign g[47285] = a[14] & g[30901];
assign g[63668] = b[14] & g[30901];
assign g[47286] = a[14] & g[30902];
assign g[63669] = b[14] & g[30902];
assign g[47287] = a[14] & g[30903];
assign g[63670] = b[14] & g[30903];
assign g[47288] = a[14] & g[30904];
assign g[63671] = b[14] & g[30904];
assign g[47289] = a[14] & g[30905];
assign g[63672] = b[14] & g[30905];
assign g[47290] = a[14] & g[30906];
assign g[63673] = b[14] & g[30906];
assign g[47291] = a[14] & g[30907];
assign g[63674] = b[14] & g[30907];
assign g[47292] = a[14] & g[30908];
assign g[63675] = b[14] & g[30908];
assign g[47293] = a[14] & g[30909];
assign g[63676] = b[14] & g[30909];
assign g[47294] = a[14] & g[30910];
assign g[63677] = b[14] & g[30910];
assign g[47295] = a[14] & g[30911];
assign g[63678] = b[14] & g[30911];
assign g[47296] = a[14] & g[30912];
assign g[63679] = b[14] & g[30912];
assign g[47297] = a[14] & g[30913];
assign g[63680] = b[14] & g[30913];
assign g[47298] = a[14] & g[30914];
assign g[63681] = b[14] & g[30914];
assign g[47299] = a[14] & g[30915];
assign g[63682] = b[14] & g[30915];
assign g[47300] = a[14] & g[30916];
assign g[63683] = b[14] & g[30916];
assign g[47301] = a[14] & g[30917];
assign g[63684] = b[14] & g[30917];
assign g[47302] = a[14] & g[30918];
assign g[63685] = b[14] & g[30918];
assign g[47303] = a[14] & g[30919];
assign g[63686] = b[14] & g[30919];
assign g[47304] = a[14] & g[30920];
assign g[63687] = b[14] & g[30920];
assign g[47305] = a[14] & g[30921];
assign g[63688] = b[14] & g[30921];
assign g[47306] = a[14] & g[30922];
assign g[63689] = b[14] & g[30922];
assign g[47307] = a[14] & g[30923];
assign g[63690] = b[14] & g[30923];
assign g[47308] = a[14] & g[30924];
assign g[63691] = b[14] & g[30924];
assign g[47309] = a[14] & g[30925];
assign g[63692] = b[14] & g[30925];
assign g[47310] = a[14] & g[30926];
assign g[63693] = b[14] & g[30926];
assign g[47311] = a[14] & g[30927];
assign g[63694] = b[14] & g[30927];
assign g[47312] = a[14] & g[30928];
assign g[63695] = b[14] & g[30928];
assign g[47313] = a[14] & g[30929];
assign g[63696] = b[14] & g[30929];
assign g[47314] = a[14] & g[30930];
assign g[63697] = b[14] & g[30930];
assign g[47315] = a[14] & g[30931];
assign g[63698] = b[14] & g[30931];
assign g[47316] = a[14] & g[30932];
assign g[63699] = b[14] & g[30932];
assign g[47317] = a[14] & g[30933];
assign g[63700] = b[14] & g[30933];
assign g[47318] = a[14] & g[30934];
assign g[63701] = b[14] & g[30934];
assign g[47319] = a[14] & g[30935];
assign g[63702] = b[14] & g[30935];
assign g[47320] = a[14] & g[30936];
assign g[63703] = b[14] & g[30936];
assign g[47321] = a[14] & g[30937];
assign g[63704] = b[14] & g[30937];
assign g[47322] = a[14] & g[30938];
assign g[63705] = b[14] & g[30938];
assign g[47323] = a[14] & g[30939];
assign g[63706] = b[14] & g[30939];
assign g[47324] = a[14] & g[30940];
assign g[63707] = b[14] & g[30940];
assign g[47325] = a[14] & g[30941];
assign g[63708] = b[14] & g[30941];
assign g[47326] = a[14] & g[30942];
assign g[63709] = b[14] & g[30942];
assign g[47327] = a[14] & g[30943];
assign g[63710] = b[14] & g[30943];
assign g[47328] = a[14] & g[30944];
assign g[63711] = b[14] & g[30944];
assign g[47329] = a[14] & g[30945];
assign g[63712] = b[14] & g[30945];
assign g[47330] = a[14] & g[30946];
assign g[63713] = b[14] & g[30946];
assign g[47331] = a[14] & g[30947];
assign g[63714] = b[14] & g[30947];
assign g[47332] = a[14] & g[30948];
assign g[63715] = b[14] & g[30948];
assign g[47333] = a[14] & g[30949];
assign g[63716] = b[14] & g[30949];
assign g[47334] = a[14] & g[30950];
assign g[63717] = b[14] & g[30950];
assign g[47335] = a[14] & g[30951];
assign g[63718] = b[14] & g[30951];
assign g[47336] = a[14] & g[30952];
assign g[63719] = b[14] & g[30952];
assign g[47337] = a[14] & g[30953];
assign g[63720] = b[14] & g[30953];
assign g[47338] = a[14] & g[30954];
assign g[63721] = b[14] & g[30954];
assign g[47339] = a[14] & g[30955];
assign g[63722] = b[14] & g[30955];
assign g[47340] = a[14] & g[30956];
assign g[63723] = b[14] & g[30956];
assign g[47341] = a[14] & g[30957];
assign g[63724] = b[14] & g[30957];
assign g[47342] = a[14] & g[30958];
assign g[63725] = b[14] & g[30958];
assign g[47343] = a[14] & g[30959];
assign g[63726] = b[14] & g[30959];
assign g[47344] = a[14] & g[30960];
assign g[63727] = b[14] & g[30960];
assign g[47345] = a[14] & g[30961];
assign g[63728] = b[14] & g[30961];
assign g[47346] = a[14] & g[30962];
assign g[63729] = b[14] & g[30962];
assign g[47347] = a[14] & g[30963];
assign g[63730] = b[14] & g[30963];
assign g[47348] = a[14] & g[30964];
assign g[63731] = b[14] & g[30964];
assign g[47349] = a[14] & g[30965];
assign g[63732] = b[14] & g[30965];
assign g[47350] = a[14] & g[30966];
assign g[63733] = b[14] & g[30966];
assign g[47351] = a[14] & g[30967];
assign g[63734] = b[14] & g[30967];
assign g[47352] = a[14] & g[30968];
assign g[63735] = b[14] & g[30968];
assign g[47353] = a[14] & g[30969];
assign g[63736] = b[14] & g[30969];
assign g[47354] = a[14] & g[30970];
assign g[63737] = b[14] & g[30970];
assign g[47355] = a[14] & g[30971];
assign g[63738] = b[14] & g[30971];
assign g[47356] = a[14] & g[30972];
assign g[63739] = b[14] & g[30972];
assign g[47357] = a[14] & g[30973];
assign g[63740] = b[14] & g[30973];
assign g[47358] = a[14] & g[30974];
assign g[63741] = b[14] & g[30974];
assign g[47359] = a[14] & g[30975];
assign g[63742] = b[14] & g[30975];
assign g[47360] = a[14] & g[30976];
assign g[63743] = b[14] & g[30976];
assign g[47361] = a[14] & g[30977];
assign g[63744] = b[14] & g[30977];
assign g[47362] = a[14] & g[30978];
assign g[63745] = b[14] & g[30978];
assign g[47363] = a[14] & g[30979];
assign g[63746] = b[14] & g[30979];
assign g[47364] = a[14] & g[30980];
assign g[63747] = b[14] & g[30980];
assign g[47365] = a[14] & g[30981];
assign g[63748] = b[14] & g[30981];
assign g[47366] = a[14] & g[30982];
assign g[63749] = b[14] & g[30982];
assign g[47367] = a[14] & g[30983];
assign g[63750] = b[14] & g[30983];
assign g[47368] = a[14] & g[30984];
assign g[63751] = b[14] & g[30984];
assign g[47369] = a[14] & g[30985];
assign g[63752] = b[14] & g[30985];
assign g[47370] = a[14] & g[30986];
assign g[63753] = b[14] & g[30986];
assign g[47371] = a[14] & g[30987];
assign g[63754] = b[14] & g[30987];
assign g[47372] = a[14] & g[30988];
assign g[63755] = b[14] & g[30988];
assign g[47373] = a[14] & g[30989];
assign g[63756] = b[14] & g[30989];
assign g[47374] = a[14] & g[30990];
assign g[63757] = b[14] & g[30990];
assign g[47375] = a[14] & g[30991];
assign g[63758] = b[14] & g[30991];
assign g[47376] = a[14] & g[30992];
assign g[63759] = b[14] & g[30992];
assign g[47377] = a[14] & g[30993];
assign g[63760] = b[14] & g[30993];
assign g[47378] = a[14] & g[30994];
assign g[63761] = b[14] & g[30994];
assign g[47379] = a[14] & g[30995];
assign g[63762] = b[14] & g[30995];
assign g[47380] = a[14] & g[30996];
assign g[63763] = b[14] & g[30996];
assign g[47381] = a[14] & g[30997];
assign g[63764] = b[14] & g[30997];
assign g[47382] = a[14] & g[30998];
assign g[63765] = b[14] & g[30998];
assign g[47383] = a[14] & g[30999];
assign g[63766] = b[14] & g[30999];
assign g[47384] = a[14] & g[31000];
assign g[63767] = b[14] & g[31000];
assign g[47385] = a[14] & g[31001];
assign g[63768] = b[14] & g[31001];
assign g[47386] = a[14] & g[31002];
assign g[63769] = b[14] & g[31002];
assign g[47387] = a[14] & g[31003];
assign g[63770] = b[14] & g[31003];
assign g[47388] = a[14] & g[31004];
assign g[63771] = b[14] & g[31004];
assign g[47389] = a[14] & g[31005];
assign g[63772] = b[14] & g[31005];
assign g[47390] = a[14] & g[31006];
assign g[63773] = b[14] & g[31006];
assign g[47391] = a[14] & g[31007];
assign g[63774] = b[14] & g[31007];
assign g[47392] = a[14] & g[31008];
assign g[63775] = b[14] & g[31008];
assign g[47393] = a[14] & g[31009];
assign g[63776] = b[14] & g[31009];
assign g[47394] = a[14] & g[31010];
assign g[63777] = b[14] & g[31010];
assign g[47395] = a[14] & g[31011];
assign g[63778] = b[14] & g[31011];
assign g[47396] = a[14] & g[31012];
assign g[63779] = b[14] & g[31012];
assign g[47397] = a[14] & g[31013];
assign g[63780] = b[14] & g[31013];
assign g[47398] = a[14] & g[31014];
assign g[63781] = b[14] & g[31014];
assign g[47399] = a[14] & g[31015];
assign g[63782] = b[14] & g[31015];
assign g[47400] = a[14] & g[31016];
assign g[63783] = b[14] & g[31016];
assign g[47401] = a[14] & g[31017];
assign g[63784] = b[14] & g[31017];
assign g[47402] = a[14] & g[31018];
assign g[63785] = b[14] & g[31018];
assign g[47403] = a[14] & g[31019];
assign g[63786] = b[14] & g[31019];
assign g[47404] = a[14] & g[31020];
assign g[63787] = b[14] & g[31020];
assign g[47405] = a[14] & g[31021];
assign g[63788] = b[14] & g[31021];
assign g[47406] = a[14] & g[31022];
assign g[63789] = b[14] & g[31022];
assign g[47407] = a[14] & g[31023];
assign g[63790] = b[14] & g[31023];
assign g[47408] = a[14] & g[31024];
assign g[63791] = b[14] & g[31024];
assign g[47409] = a[14] & g[31025];
assign g[63792] = b[14] & g[31025];
assign g[47410] = a[14] & g[31026];
assign g[63793] = b[14] & g[31026];
assign g[47411] = a[14] & g[31027];
assign g[63794] = b[14] & g[31027];
assign g[47412] = a[14] & g[31028];
assign g[63795] = b[14] & g[31028];
assign g[47413] = a[14] & g[31029];
assign g[63796] = b[14] & g[31029];
assign g[47414] = a[14] & g[31030];
assign g[63797] = b[14] & g[31030];
assign g[47415] = a[14] & g[31031];
assign g[63798] = b[14] & g[31031];
assign g[47416] = a[14] & g[31032];
assign g[63799] = b[14] & g[31032];
assign g[47417] = a[14] & g[31033];
assign g[63800] = b[14] & g[31033];
assign g[47418] = a[14] & g[31034];
assign g[63801] = b[14] & g[31034];
assign g[47419] = a[14] & g[31035];
assign g[63802] = b[14] & g[31035];
assign g[47420] = a[14] & g[31036];
assign g[63803] = b[14] & g[31036];
assign g[47421] = a[14] & g[31037];
assign g[63804] = b[14] & g[31037];
assign g[47422] = a[14] & g[31038];
assign g[63805] = b[14] & g[31038];
assign g[47423] = a[14] & g[31039];
assign g[63806] = b[14] & g[31039];
assign g[47424] = a[14] & g[31040];
assign g[63807] = b[14] & g[31040];
assign g[47425] = a[14] & g[31041];
assign g[63808] = b[14] & g[31041];
assign g[47426] = a[14] & g[31042];
assign g[63809] = b[14] & g[31042];
assign g[47427] = a[14] & g[31043];
assign g[63810] = b[14] & g[31043];
assign g[47428] = a[14] & g[31044];
assign g[63811] = b[14] & g[31044];
assign g[47429] = a[14] & g[31045];
assign g[63812] = b[14] & g[31045];
assign g[47430] = a[14] & g[31046];
assign g[63813] = b[14] & g[31046];
assign g[47431] = a[14] & g[31047];
assign g[63814] = b[14] & g[31047];
assign g[47432] = a[14] & g[31048];
assign g[63815] = b[14] & g[31048];
assign g[47433] = a[14] & g[31049];
assign g[63816] = b[14] & g[31049];
assign g[47434] = a[14] & g[31050];
assign g[63817] = b[14] & g[31050];
assign g[47435] = a[14] & g[31051];
assign g[63818] = b[14] & g[31051];
assign g[47436] = a[14] & g[31052];
assign g[63819] = b[14] & g[31052];
assign g[47437] = a[14] & g[31053];
assign g[63820] = b[14] & g[31053];
assign g[47438] = a[14] & g[31054];
assign g[63821] = b[14] & g[31054];
assign g[47439] = a[14] & g[31055];
assign g[63822] = b[14] & g[31055];
assign g[47440] = a[14] & g[31056];
assign g[63823] = b[14] & g[31056];
assign g[47441] = a[14] & g[31057];
assign g[63824] = b[14] & g[31057];
assign g[47442] = a[14] & g[31058];
assign g[63825] = b[14] & g[31058];
assign g[47443] = a[14] & g[31059];
assign g[63826] = b[14] & g[31059];
assign g[47444] = a[14] & g[31060];
assign g[63827] = b[14] & g[31060];
assign g[47445] = a[14] & g[31061];
assign g[63828] = b[14] & g[31061];
assign g[47446] = a[14] & g[31062];
assign g[63829] = b[14] & g[31062];
assign g[47447] = a[14] & g[31063];
assign g[63830] = b[14] & g[31063];
assign g[47448] = a[14] & g[31064];
assign g[63831] = b[14] & g[31064];
assign g[47449] = a[14] & g[31065];
assign g[63832] = b[14] & g[31065];
assign g[47450] = a[14] & g[31066];
assign g[63833] = b[14] & g[31066];
assign g[47451] = a[14] & g[31067];
assign g[63834] = b[14] & g[31067];
assign g[47452] = a[14] & g[31068];
assign g[63835] = b[14] & g[31068];
assign g[47453] = a[14] & g[31069];
assign g[63836] = b[14] & g[31069];
assign g[47454] = a[14] & g[31070];
assign g[63837] = b[14] & g[31070];
assign g[47455] = a[14] & g[31071];
assign g[63838] = b[14] & g[31071];
assign g[47456] = a[14] & g[31072];
assign g[63839] = b[14] & g[31072];
assign g[47457] = a[14] & g[31073];
assign g[63840] = b[14] & g[31073];
assign g[47458] = a[14] & g[31074];
assign g[63841] = b[14] & g[31074];
assign g[47459] = a[14] & g[31075];
assign g[63842] = b[14] & g[31075];
assign g[47460] = a[14] & g[31076];
assign g[63843] = b[14] & g[31076];
assign g[47461] = a[14] & g[31077];
assign g[63844] = b[14] & g[31077];
assign g[47462] = a[14] & g[31078];
assign g[63845] = b[14] & g[31078];
assign g[47463] = a[14] & g[31079];
assign g[63846] = b[14] & g[31079];
assign g[47464] = a[14] & g[31080];
assign g[63847] = b[14] & g[31080];
assign g[47465] = a[14] & g[31081];
assign g[63848] = b[14] & g[31081];
assign g[47466] = a[14] & g[31082];
assign g[63849] = b[14] & g[31082];
assign g[47467] = a[14] & g[31083];
assign g[63850] = b[14] & g[31083];
assign g[47468] = a[14] & g[31084];
assign g[63851] = b[14] & g[31084];
assign g[47469] = a[14] & g[31085];
assign g[63852] = b[14] & g[31085];
assign g[47470] = a[14] & g[31086];
assign g[63853] = b[14] & g[31086];
assign g[47471] = a[14] & g[31087];
assign g[63854] = b[14] & g[31087];
assign g[47472] = a[14] & g[31088];
assign g[63855] = b[14] & g[31088];
assign g[47473] = a[14] & g[31089];
assign g[63856] = b[14] & g[31089];
assign g[47474] = a[14] & g[31090];
assign g[63857] = b[14] & g[31090];
assign g[47475] = a[14] & g[31091];
assign g[63858] = b[14] & g[31091];
assign g[47476] = a[14] & g[31092];
assign g[63859] = b[14] & g[31092];
assign g[47477] = a[14] & g[31093];
assign g[63860] = b[14] & g[31093];
assign g[47478] = a[14] & g[31094];
assign g[63861] = b[14] & g[31094];
assign g[47479] = a[14] & g[31095];
assign g[63862] = b[14] & g[31095];
assign g[47480] = a[14] & g[31096];
assign g[63863] = b[14] & g[31096];
assign g[47481] = a[14] & g[31097];
assign g[63864] = b[14] & g[31097];
assign g[47482] = a[14] & g[31098];
assign g[63865] = b[14] & g[31098];
assign g[47483] = a[14] & g[31099];
assign g[63866] = b[14] & g[31099];
assign g[47484] = a[14] & g[31100];
assign g[63867] = b[14] & g[31100];
assign g[47485] = a[14] & g[31101];
assign g[63868] = b[14] & g[31101];
assign g[47486] = a[14] & g[31102];
assign g[63869] = b[14] & g[31102];
assign g[47487] = a[14] & g[31103];
assign g[63870] = b[14] & g[31103];
assign g[47488] = a[14] & g[31104];
assign g[63871] = b[14] & g[31104];
assign g[47489] = a[14] & g[31105];
assign g[63872] = b[14] & g[31105];
assign g[47490] = a[14] & g[31106];
assign g[63873] = b[14] & g[31106];
assign g[47491] = a[14] & g[31107];
assign g[63874] = b[14] & g[31107];
assign g[47492] = a[14] & g[31108];
assign g[63875] = b[14] & g[31108];
assign g[47493] = a[14] & g[31109];
assign g[63876] = b[14] & g[31109];
assign g[47494] = a[14] & g[31110];
assign g[63877] = b[14] & g[31110];
assign g[47495] = a[14] & g[31111];
assign g[63878] = b[14] & g[31111];
assign g[47496] = a[14] & g[31112];
assign g[63879] = b[14] & g[31112];
assign g[47497] = a[14] & g[31113];
assign g[63880] = b[14] & g[31113];
assign g[47498] = a[14] & g[31114];
assign g[63881] = b[14] & g[31114];
assign g[47499] = a[14] & g[31115];
assign g[63882] = b[14] & g[31115];
assign g[47500] = a[14] & g[31116];
assign g[63883] = b[14] & g[31116];
assign g[47501] = a[14] & g[31117];
assign g[63884] = b[14] & g[31117];
assign g[47502] = a[14] & g[31118];
assign g[63885] = b[14] & g[31118];
assign g[47503] = a[14] & g[31119];
assign g[63886] = b[14] & g[31119];
assign g[47504] = a[14] & g[31120];
assign g[63887] = b[14] & g[31120];
assign g[47505] = a[14] & g[31121];
assign g[63888] = b[14] & g[31121];
assign g[47506] = a[14] & g[31122];
assign g[63889] = b[14] & g[31122];
assign g[47507] = a[14] & g[31123];
assign g[63890] = b[14] & g[31123];
assign g[47508] = a[14] & g[31124];
assign g[63891] = b[14] & g[31124];
assign g[47509] = a[14] & g[31125];
assign g[63892] = b[14] & g[31125];
assign g[47510] = a[14] & g[31126];
assign g[63893] = b[14] & g[31126];
assign g[47511] = a[14] & g[31127];
assign g[63894] = b[14] & g[31127];
assign g[47512] = a[14] & g[31128];
assign g[63895] = b[14] & g[31128];
assign g[47513] = a[14] & g[31129];
assign g[63896] = b[14] & g[31129];
assign g[47514] = a[14] & g[31130];
assign g[63897] = b[14] & g[31130];
assign g[47515] = a[14] & g[31131];
assign g[63898] = b[14] & g[31131];
assign g[47516] = a[14] & g[31132];
assign g[63899] = b[14] & g[31132];
assign g[47517] = a[14] & g[31133];
assign g[63900] = b[14] & g[31133];
assign g[47518] = a[14] & g[31134];
assign g[63901] = b[14] & g[31134];
assign g[47519] = a[14] & g[31135];
assign g[63902] = b[14] & g[31135];
assign g[47520] = a[14] & g[31136];
assign g[63903] = b[14] & g[31136];
assign g[47521] = a[14] & g[31137];
assign g[63904] = b[14] & g[31137];
assign g[47522] = a[14] & g[31138];
assign g[63905] = b[14] & g[31138];
assign g[47523] = a[14] & g[31139];
assign g[63906] = b[14] & g[31139];
assign g[47524] = a[14] & g[31140];
assign g[63907] = b[14] & g[31140];
assign g[47525] = a[14] & g[31141];
assign g[63908] = b[14] & g[31141];
assign g[47526] = a[14] & g[31142];
assign g[63909] = b[14] & g[31142];
assign g[47527] = a[14] & g[31143];
assign g[63910] = b[14] & g[31143];
assign g[47528] = a[14] & g[31144];
assign g[63911] = b[14] & g[31144];
assign g[47529] = a[14] & g[31145];
assign g[63912] = b[14] & g[31145];
assign g[47530] = a[14] & g[31146];
assign g[63913] = b[14] & g[31146];
assign g[47531] = a[14] & g[31147];
assign g[63914] = b[14] & g[31147];
assign g[47532] = a[14] & g[31148];
assign g[63915] = b[14] & g[31148];
assign g[47533] = a[14] & g[31149];
assign g[63916] = b[14] & g[31149];
assign g[47534] = a[14] & g[31150];
assign g[63917] = b[14] & g[31150];
assign g[47535] = a[14] & g[31151];
assign g[63918] = b[14] & g[31151];
assign g[47536] = a[14] & g[31152];
assign g[63919] = b[14] & g[31152];
assign g[47537] = a[14] & g[31153];
assign g[63920] = b[14] & g[31153];
assign g[47538] = a[14] & g[31154];
assign g[63921] = b[14] & g[31154];
assign g[47539] = a[14] & g[31155];
assign g[63922] = b[14] & g[31155];
assign g[47540] = a[14] & g[31156];
assign g[63923] = b[14] & g[31156];
assign g[47541] = a[14] & g[31157];
assign g[63924] = b[14] & g[31157];
assign g[47542] = a[14] & g[31158];
assign g[63925] = b[14] & g[31158];
assign g[47543] = a[14] & g[31159];
assign g[63926] = b[14] & g[31159];
assign g[47544] = a[14] & g[31160];
assign g[63927] = b[14] & g[31160];
assign g[47545] = a[14] & g[31161];
assign g[63928] = b[14] & g[31161];
assign g[47546] = a[14] & g[31162];
assign g[63929] = b[14] & g[31162];
assign g[47547] = a[14] & g[31163];
assign g[63930] = b[14] & g[31163];
assign g[47548] = a[14] & g[31164];
assign g[63931] = b[14] & g[31164];
assign g[47549] = a[14] & g[31165];
assign g[63932] = b[14] & g[31165];
assign g[47550] = a[14] & g[31166];
assign g[63933] = b[14] & g[31166];
assign g[47551] = a[14] & g[31167];
assign g[63934] = b[14] & g[31167];
assign g[47552] = a[14] & g[31168];
assign g[63935] = b[14] & g[31168];
assign g[47553] = a[14] & g[31169];
assign g[63936] = b[14] & g[31169];
assign g[47554] = a[14] & g[31170];
assign g[63937] = b[14] & g[31170];
assign g[47555] = a[14] & g[31171];
assign g[63938] = b[14] & g[31171];
assign g[47556] = a[14] & g[31172];
assign g[63939] = b[14] & g[31172];
assign g[47557] = a[14] & g[31173];
assign g[63940] = b[14] & g[31173];
assign g[47558] = a[14] & g[31174];
assign g[63941] = b[14] & g[31174];
assign g[47559] = a[14] & g[31175];
assign g[63942] = b[14] & g[31175];
assign g[47560] = a[14] & g[31176];
assign g[63943] = b[14] & g[31176];
assign g[47561] = a[14] & g[31177];
assign g[63944] = b[14] & g[31177];
assign g[47562] = a[14] & g[31178];
assign g[63945] = b[14] & g[31178];
assign g[47563] = a[14] & g[31179];
assign g[63946] = b[14] & g[31179];
assign g[47564] = a[14] & g[31180];
assign g[63947] = b[14] & g[31180];
assign g[47565] = a[14] & g[31181];
assign g[63948] = b[14] & g[31181];
assign g[47566] = a[14] & g[31182];
assign g[63949] = b[14] & g[31182];
assign g[47567] = a[14] & g[31183];
assign g[63950] = b[14] & g[31183];
assign g[47568] = a[14] & g[31184];
assign g[63951] = b[14] & g[31184];
assign g[47569] = a[14] & g[31185];
assign g[63952] = b[14] & g[31185];
assign g[47570] = a[14] & g[31186];
assign g[63953] = b[14] & g[31186];
assign g[47571] = a[14] & g[31187];
assign g[63954] = b[14] & g[31187];
assign g[47572] = a[14] & g[31188];
assign g[63955] = b[14] & g[31188];
assign g[47573] = a[14] & g[31189];
assign g[63956] = b[14] & g[31189];
assign g[47574] = a[14] & g[31190];
assign g[63957] = b[14] & g[31190];
assign g[47575] = a[14] & g[31191];
assign g[63958] = b[14] & g[31191];
assign g[47576] = a[14] & g[31192];
assign g[63959] = b[14] & g[31192];
assign g[47577] = a[14] & g[31193];
assign g[63960] = b[14] & g[31193];
assign g[47578] = a[14] & g[31194];
assign g[63961] = b[14] & g[31194];
assign g[47579] = a[14] & g[31195];
assign g[63962] = b[14] & g[31195];
assign g[47580] = a[14] & g[31196];
assign g[63963] = b[14] & g[31196];
assign g[47581] = a[14] & g[31197];
assign g[63964] = b[14] & g[31197];
assign g[47582] = a[14] & g[31198];
assign g[63965] = b[14] & g[31198];
assign g[47583] = a[14] & g[31199];
assign g[63966] = b[14] & g[31199];
assign g[47584] = a[14] & g[31200];
assign g[63967] = b[14] & g[31200];
assign g[47585] = a[14] & g[31201];
assign g[63968] = b[14] & g[31201];
assign g[47586] = a[14] & g[31202];
assign g[63969] = b[14] & g[31202];
assign g[47587] = a[14] & g[31203];
assign g[63970] = b[14] & g[31203];
assign g[47588] = a[14] & g[31204];
assign g[63971] = b[14] & g[31204];
assign g[47589] = a[14] & g[31205];
assign g[63972] = b[14] & g[31205];
assign g[47590] = a[14] & g[31206];
assign g[63973] = b[14] & g[31206];
assign g[47591] = a[14] & g[31207];
assign g[63974] = b[14] & g[31207];
assign g[47592] = a[14] & g[31208];
assign g[63975] = b[14] & g[31208];
assign g[47593] = a[14] & g[31209];
assign g[63976] = b[14] & g[31209];
assign g[47594] = a[14] & g[31210];
assign g[63977] = b[14] & g[31210];
assign g[47595] = a[14] & g[31211];
assign g[63978] = b[14] & g[31211];
assign g[47596] = a[14] & g[31212];
assign g[63979] = b[14] & g[31212];
assign g[47597] = a[14] & g[31213];
assign g[63980] = b[14] & g[31213];
assign g[47598] = a[14] & g[31214];
assign g[63981] = b[14] & g[31214];
assign g[47599] = a[14] & g[31215];
assign g[63982] = b[14] & g[31215];
assign g[47600] = a[14] & g[31216];
assign g[63983] = b[14] & g[31216];
assign g[47601] = a[14] & g[31217];
assign g[63984] = b[14] & g[31217];
assign g[47602] = a[14] & g[31218];
assign g[63985] = b[14] & g[31218];
assign g[47603] = a[14] & g[31219];
assign g[63986] = b[14] & g[31219];
assign g[47604] = a[14] & g[31220];
assign g[63987] = b[14] & g[31220];
assign g[47605] = a[14] & g[31221];
assign g[63988] = b[14] & g[31221];
assign g[47606] = a[14] & g[31222];
assign g[63989] = b[14] & g[31222];
assign g[47607] = a[14] & g[31223];
assign g[63990] = b[14] & g[31223];
assign g[47608] = a[14] & g[31224];
assign g[63991] = b[14] & g[31224];
assign g[47609] = a[14] & g[31225];
assign g[63992] = b[14] & g[31225];
assign g[47610] = a[14] & g[31226];
assign g[63993] = b[14] & g[31226];
assign g[47611] = a[14] & g[31227];
assign g[63994] = b[14] & g[31227];
assign g[47612] = a[14] & g[31228];
assign g[63995] = b[14] & g[31228];
assign g[47613] = a[14] & g[31229];
assign g[63996] = b[14] & g[31229];
assign g[47614] = a[14] & g[31230];
assign g[63997] = b[14] & g[31230];
assign g[47615] = a[14] & g[31231];
assign g[63998] = b[14] & g[31231];
assign g[47616] = a[14] & g[31232];
assign g[63999] = b[14] & g[31232];
assign g[47617] = a[14] & g[31233];
assign g[64000] = b[14] & g[31233];
assign g[47618] = a[14] & g[31234];
assign g[64001] = b[14] & g[31234];
assign g[47619] = a[14] & g[31235];
assign g[64002] = b[14] & g[31235];
assign g[47620] = a[14] & g[31236];
assign g[64003] = b[14] & g[31236];
assign g[47621] = a[14] & g[31237];
assign g[64004] = b[14] & g[31237];
assign g[47622] = a[14] & g[31238];
assign g[64005] = b[14] & g[31238];
assign g[47623] = a[14] & g[31239];
assign g[64006] = b[14] & g[31239];
assign g[47624] = a[14] & g[31240];
assign g[64007] = b[14] & g[31240];
assign g[47625] = a[14] & g[31241];
assign g[64008] = b[14] & g[31241];
assign g[47626] = a[14] & g[31242];
assign g[64009] = b[14] & g[31242];
assign g[47627] = a[14] & g[31243];
assign g[64010] = b[14] & g[31243];
assign g[47628] = a[14] & g[31244];
assign g[64011] = b[14] & g[31244];
assign g[47629] = a[14] & g[31245];
assign g[64012] = b[14] & g[31245];
assign g[47630] = a[14] & g[31246];
assign g[64013] = b[14] & g[31246];
assign g[47631] = a[14] & g[31247];
assign g[64014] = b[14] & g[31247];
assign g[47632] = a[14] & g[31248];
assign g[64015] = b[14] & g[31248];
assign g[47633] = a[14] & g[31249];
assign g[64016] = b[14] & g[31249];
assign g[47634] = a[14] & g[31250];
assign g[64017] = b[14] & g[31250];
assign g[47635] = a[14] & g[31251];
assign g[64018] = b[14] & g[31251];
assign g[47636] = a[14] & g[31252];
assign g[64019] = b[14] & g[31252];
assign g[47637] = a[14] & g[31253];
assign g[64020] = b[14] & g[31253];
assign g[47638] = a[14] & g[31254];
assign g[64021] = b[14] & g[31254];
assign g[47639] = a[14] & g[31255];
assign g[64022] = b[14] & g[31255];
assign g[47640] = a[14] & g[31256];
assign g[64023] = b[14] & g[31256];
assign g[47641] = a[14] & g[31257];
assign g[64024] = b[14] & g[31257];
assign g[47642] = a[14] & g[31258];
assign g[64025] = b[14] & g[31258];
assign g[47643] = a[14] & g[31259];
assign g[64026] = b[14] & g[31259];
assign g[47644] = a[14] & g[31260];
assign g[64027] = b[14] & g[31260];
assign g[47645] = a[14] & g[31261];
assign g[64028] = b[14] & g[31261];
assign g[47646] = a[14] & g[31262];
assign g[64029] = b[14] & g[31262];
assign g[47647] = a[14] & g[31263];
assign g[64030] = b[14] & g[31263];
assign g[47648] = a[14] & g[31264];
assign g[64031] = b[14] & g[31264];
assign g[47649] = a[14] & g[31265];
assign g[64032] = b[14] & g[31265];
assign g[47650] = a[14] & g[31266];
assign g[64033] = b[14] & g[31266];
assign g[47651] = a[14] & g[31267];
assign g[64034] = b[14] & g[31267];
assign g[47652] = a[14] & g[31268];
assign g[64035] = b[14] & g[31268];
assign g[47653] = a[14] & g[31269];
assign g[64036] = b[14] & g[31269];
assign g[47654] = a[14] & g[31270];
assign g[64037] = b[14] & g[31270];
assign g[47655] = a[14] & g[31271];
assign g[64038] = b[14] & g[31271];
assign g[47656] = a[14] & g[31272];
assign g[64039] = b[14] & g[31272];
assign g[47657] = a[14] & g[31273];
assign g[64040] = b[14] & g[31273];
assign g[47658] = a[14] & g[31274];
assign g[64041] = b[14] & g[31274];
assign g[47659] = a[14] & g[31275];
assign g[64042] = b[14] & g[31275];
assign g[47660] = a[14] & g[31276];
assign g[64043] = b[14] & g[31276];
assign g[47661] = a[14] & g[31277];
assign g[64044] = b[14] & g[31277];
assign g[47662] = a[14] & g[31278];
assign g[64045] = b[14] & g[31278];
assign g[47663] = a[14] & g[31279];
assign g[64046] = b[14] & g[31279];
assign g[47664] = a[14] & g[31280];
assign g[64047] = b[14] & g[31280];
assign g[47665] = a[14] & g[31281];
assign g[64048] = b[14] & g[31281];
assign g[47666] = a[14] & g[31282];
assign g[64049] = b[14] & g[31282];
assign g[47667] = a[14] & g[31283];
assign g[64050] = b[14] & g[31283];
assign g[47668] = a[14] & g[31284];
assign g[64051] = b[14] & g[31284];
assign g[47669] = a[14] & g[31285];
assign g[64052] = b[14] & g[31285];
assign g[47670] = a[14] & g[31286];
assign g[64053] = b[14] & g[31286];
assign g[47671] = a[14] & g[31287];
assign g[64054] = b[14] & g[31287];
assign g[47672] = a[14] & g[31288];
assign g[64055] = b[14] & g[31288];
assign g[47673] = a[14] & g[31289];
assign g[64056] = b[14] & g[31289];
assign g[47674] = a[14] & g[31290];
assign g[64057] = b[14] & g[31290];
assign g[47675] = a[14] & g[31291];
assign g[64058] = b[14] & g[31291];
assign g[47676] = a[14] & g[31292];
assign g[64059] = b[14] & g[31292];
assign g[47677] = a[14] & g[31293];
assign g[64060] = b[14] & g[31293];
assign g[47678] = a[14] & g[31294];
assign g[64061] = b[14] & g[31294];
assign g[47679] = a[14] & g[31295];
assign g[64062] = b[14] & g[31295];
assign g[47680] = a[14] & g[31296];
assign g[64063] = b[14] & g[31296];
assign g[47681] = a[14] & g[31297];
assign g[64064] = b[14] & g[31297];
assign g[47682] = a[14] & g[31298];
assign g[64065] = b[14] & g[31298];
assign g[47683] = a[14] & g[31299];
assign g[64066] = b[14] & g[31299];
assign g[47684] = a[14] & g[31300];
assign g[64067] = b[14] & g[31300];
assign g[47685] = a[14] & g[31301];
assign g[64068] = b[14] & g[31301];
assign g[47686] = a[14] & g[31302];
assign g[64069] = b[14] & g[31302];
assign g[47687] = a[14] & g[31303];
assign g[64070] = b[14] & g[31303];
assign g[47688] = a[14] & g[31304];
assign g[64071] = b[14] & g[31304];
assign g[47689] = a[14] & g[31305];
assign g[64072] = b[14] & g[31305];
assign g[47690] = a[14] & g[31306];
assign g[64073] = b[14] & g[31306];
assign g[47691] = a[14] & g[31307];
assign g[64074] = b[14] & g[31307];
assign g[47692] = a[14] & g[31308];
assign g[64075] = b[14] & g[31308];
assign g[47693] = a[14] & g[31309];
assign g[64076] = b[14] & g[31309];
assign g[47694] = a[14] & g[31310];
assign g[64077] = b[14] & g[31310];
assign g[47695] = a[14] & g[31311];
assign g[64078] = b[14] & g[31311];
assign g[47696] = a[14] & g[31312];
assign g[64079] = b[14] & g[31312];
assign g[47697] = a[14] & g[31313];
assign g[64080] = b[14] & g[31313];
assign g[47698] = a[14] & g[31314];
assign g[64081] = b[14] & g[31314];
assign g[47699] = a[14] & g[31315];
assign g[64082] = b[14] & g[31315];
assign g[47700] = a[14] & g[31316];
assign g[64083] = b[14] & g[31316];
assign g[47701] = a[14] & g[31317];
assign g[64084] = b[14] & g[31317];
assign g[47702] = a[14] & g[31318];
assign g[64085] = b[14] & g[31318];
assign g[47703] = a[14] & g[31319];
assign g[64086] = b[14] & g[31319];
assign g[47704] = a[14] & g[31320];
assign g[64087] = b[14] & g[31320];
assign g[47705] = a[14] & g[31321];
assign g[64088] = b[14] & g[31321];
assign g[47706] = a[14] & g[31322];
assign g[64089] = b[14] & g[31322];
assign g[47707] = a[14] & g[31323];
assign g[64090] = b[14] & g[31323];
assign g[47708] = a[14] & g[31324];
assign g[64091] = b[14] & g[31324];
assign g[47709] = a[14] & g[31325];
assign g[64092] = b[14] & g[31325];
assign g[47710] = a[14] & g[31326];
assign g[64093] = b[14] & g[31326];
assign g[47711] = a[14] & g[31327];
assign g[64094] = b[14] & g[31327];
assign g[47712] = a[14] & g[31328];
assign g[64095] = b[14] & g[31328];
assign g[47713] = a[14] & g[31329];
assign g[64096] = b[14] & g[31329];
assign g[47714] = a[14] & g[31330];
assign g[64097] = b[14] & g[31330];
assign g[47715] = a[14] & g[31331];
assign g[64098] = b[14] & g[31331];
assign g[47716] = a[14] & g[31332];
assign g[64099] = b[14] & g[31332];
assign g[47717] = a[14] & g[31333];
assign g[64100] = b[14] & g[31333];
assign g[47718] = a[14] & g[31334];
assign g[64101] = b[14] & g[31334];
assign g[47719] = a[14] & g[31335];
assign g[64102] = b[14] & g[31335];
assign g[47720] = a[14] & g[31336];
assign g[64103] = b[14] & g[31336];
assign g[47721] = a[14] & g[31337];
assign g[64104] = b[14] & g[31337];
assign g[47722] = a[14] & g[31338];
assign g[64105] = b[14] & g[31338];
assign g[47723] = a[14] & g[31339];
assign g[64106] = b[14] & g[31339];
assign g[47724] = a[14] & g[31340];
assign g[64107] = b[14] & g[31340];
assign g[47725] = a[14] & g[31341];
assign g[64108] = b[14] & g[31341];
assign g[47726] = a[14] & g[31342];
assign g[64109] = b[14] & g[31342];
assign g[47727] = a[14] & g[31343];
assign g[64110] = b[14] & g[31343];
assign g[47728] = a[14] & g[31344];
assign g[64111] = b[14] & g[31344];
assign g[47729] = a[14] & g[31345];
assign g[64112] = b[14] & g[31345];
assign g[47730] = a[14] & g[31346];
assign g[64113] = b[14] & g[31346];
assign g[47731] = a[14] & g[31347];
assign g[64114] = b[14] & g[31347];
assign g[47732] = a[14] & g[31348];
assign g[64115] = b[14] & g[31348];
assign g[47733] = a[14] & g[31349];
assign g[64116] = b[14] & g[31349];
assign g[47734] = a[14] & g[31350];
assign g[64117] = b[14] & g[31350];
assign g[47735] = a[14] & g[31351];
assign g[64118] = b[14] & g[31351];
assign g[47736] = a[14] & g[31352];
assign g[64119] = b[14] & g[31352];
assign g[47737] = a[14] & g[31353];
assign g[64120] = b[14] & g[31353];
assign g[47738] = a[14] & g[31354];
assign g[64121] = b[14] & g[31354];
assign g[47739] = a[14] & g[31355];
assign g[64122] = b[14] & g[31355];
assign g[47740] = a[14] & g[31356];
assign g[64123] = b[14] & g[31356];
assign g[47741] = a[14] & g[31357];
assign g[64124] = b[14] & g[31357];
assign g[47742] = a[14] & g[31358];
assign g[64125] = b[14] & g[31358];
assign g[47743] = a[14] & g[31359];
assign g[64126] = b[14] & g[31359];
assign g[47744] = a[14] & g[31360];
assign g[64127] = b[14] & g[31360];
assign g[47745] = a[14] & g[31361];
assign g[64128] = b[14] & g[31361];
assign g[47746] = a[14] & g[31362];
assign g[64129] = b[14] & g[31362];
assign g[47747] = a[14] & g[31363];
assign g[64130] = b[14] & g[31363];
assign g[47748] = a[14] & g[31364];
assign g[64131] = b[14] & g[31364];
assign g[47749] = a[14] & g[31365];
assign g[64132] = b[14] & g[31365];
assign g[47750] = a[14] & g[31366];
assign g[64133] = b[14] & g[31366];
assign g[47751] = a[14] & g[31367];
assign g[64134] = b[14] & g[31367];
assign g[47752] = a[14] & g[31368];
assign g[64135] = b[14] & g[31368];
assign g[47753] = a[14] & g[31369];
assign g[64136] = b[14] & g[31369];
assign g[47754] = a[14] & g[31370];
assign g[64137] = b[14] & g[31370];
assign g[47755] = a[14] & g[31371];
assign g[64138] = b[14] & g[31371];
assign g[47756] = a[14] & g[31372];
assign g[64139] = b[14] & g[31372];
assign g[47757] = a[14] & g[31373];
assign g[64140] = b[14] & g[31373];
assign g[47758] = a[14] & g[31374];
assign g[64141] = b[14] & g[31374];
assign g[47759] = a[14] & g[31375];
assign g[64142] = b[14] & g[31375];
assign g[47760] = a[14] & g[31376];
assign g[64143] = b[14] & g[31376];
assign g[47761] = a[14] & g[31377];
assign g[64144] = b[14] & g[31377];
assign g[47762] = a[14] & g[31378];
assign g[64145] = b[14] & g[31378];
assign g[47763] = a[14] & g[31379];
assign g[64146] = b[14] & g[31379];
assign g[47764] = a[14] & g[31380];
assign g[64147] = b[14] & g[31380];
assign g[47765] = a[14] & g[31381];
assign g[64148] = b[14] & g[31381];
assign g[47766] = a[14] & g[31382];
assign g[64149] = b[14] & g[31382];
assign g[47767] = a[14] & g[31383];
assign g[64150] = b[14] & g[31383];
assign g[47768] = a[14] & g[31384];
assign g[64151] = b[14] & g[31384];
assign g[47769] = a[14] & g[31385];
assign g[64152] = b[14] & g[31385];
assign g[47770] = a[14] & g[31386];
assign g[64153] = b[14] & g[31386];
assign g[47771] = a[14] & g[31387];
assign g[64154] = b[14] & g[31387];
assign g[47772] = a[14] & g[31388];
assign g[64155] = b[14] & g[31388];
assign g[47773] = a[14] & g[31389];
assign g[64156] = b[14] & g[31389];
assign g[47774] = a[14] & g[31390];
assign g[64157] = b[14] & g[31390];
assign g[47775] = a[14] & g[31391];
assign g[64158] = b[14] & g[31391];
assign g[47776] = a[14] & g[31392];
assign g[64159] = b[14] & g[31392];
assign g[47777] = a[14] & g[31393];
assign g[64160] = b[14] & g[31393];
assign g[47778] = a[14] & g[31394];
assign g[64161] = b[14] & g[31394];
assign g[47779] = a[14] & g[31395];
assign g[64162] = b[14] & g[31395];
assign g[47780] = a[14] & g[31396];
assign g[64163] = b[14] & g[31396];
assign g[47781] = a[14] & g[31397];
assign g[64164] = b[14] & g[31397];
assign g[47782] = a[14] & g[31398];
assign g[64165] = b[14] & g[31398];
assign g[47783] = a[14] & g[31399];
assign g[64166] = b[14] & g[31399];
assign g[47784] = a[14] & g[31400];
assign g[64167] = b[14] & g[31400];
assign g[47785] = a[14] & g[31401];
assign g[64168] = b[14] & g[31401];
assign g[47786] = a[14] & g[31402];
assign g[64169] = b[14] & g[31402];
assign g[47787] = a[14] & g[31403];
assign g[64170] = b[14] & g[31403];
assign g[47788] = a[14] & g[31404];
assign g[64171] = b[14] & g[31404];
assign g[47789] = a[14] & g[31405];
assign g[64172] = b[14] & g[31405];
assign g[47790] = a[14] & g[31406];
assign g[64173] = b[14] & g[31406];
assign g[47791] = a[14] & g[31407];
assign g[64174] = b[14] & g[31407];
assign g[47792] = a[14] & g[31408];
assign g[64175] = b[14] & g[31408];
assign g[47793] = a[14] & g[31409];
assign g[64176] = b[14] & g[31409];
assign g[47794] = a[14] & g[31410];
assign g[64177] = b[14] & g[31410];
assign g[47795] = a[14] & g[31411];
assign g[64178] = b[14] & g[31411];
assign g[47796] = a[14] & g[31412];
assign g[64179] = b[14] & g[31412];
assign g[47797] = a[14] & g[31413];
assign g[64180] = b[14] & g[31413];
assign g[47798] = a[14] & g[31414];
assign g[64181] = b[14] & g[31414];
assign g[47799] = a[14] & g[31415];
assign g[64182] = b[14] & g[31415];
assign g[47800] = a[14] & g[31416];
assign g[64183] = b[14] & g[31416];
assign g[47801] = a[14] & g[31417];
assign g[64184] = b[14] & g[31417];
assign g[47802] = a[14] & g[31418];
assign g[64185] = b[14] & g[31418];
assign g[47803] = a[14] & g[31419];
assign g[64186] = b[14] & g[31419];
assign g[47804] = a[14] & g[31420];
assign g[64187] = b[14] & g[31420];
assign g[47805] = a[14] & g[31421];
assign g[64188] = b[14] & g[31421];
assign g[47806] = a[14] & g[31422];
assign g[64189] = b[14] & g[31422];
assign g[47807] = a[14] & g[31423];
assign g[64190] = b[14] & g[31423];
assign g[47808] = a[14] & g[31424];
assign g[64191] = b[14] & g[31424];
assign g[47809] = a[14] & g[31425];
assign g[64192] = b[14] & g[31425];
assign g[47810] = a[14] & g[31426];
assign g[64193] = b[14] & g[31426];
assign g[47811] = a[14] & g[31427];
assign g[64194] = b[14] & g[31427];
assign g[47812] = a[14] & g[31428];
assign g[64195] = b[14] & g[31428];
assign g[47813] = a[14] & g[31429];
assign g[64196] = b[14] & g[31429];
assign g[47814] = a[14] & g[31430];
assign g[64197] = b[14] & g[31430];
assign g[47815] = a[14] & g[31431];
assign g[64198] = b[14] & g[31431];
assign g[47816] = a[14] & g[31432];
assign g[64199] = b[14] & g[31432];
assign g[47817] = a[14] & g[31433];
assign g[64200] = b[14] & g[31433];
assign g[47818] = a[14] & g[31434];
assign g[64201] = b[14] & g[31434];
assign g[47819] = a[14] & g[31435];
assign g[64202] = b[14] & g[31435];
assign g[47820] = a[14] & g[31436];
assign g[64203] = b[14] & g[31436];
assign g[47821] = a[14] & g[31437];
assign g[64204] = b[14] & g[31437];
assign g[47822] = a[14] & g[31438];
assign g[64205] = b[14] & g[31438];
assign g[47823] = a[14] & g[31439];
assign g[64206] = b[14] & g[31439];
assign g[47824] = a[14] & g[31440];
assign g[64207] = b[14] & g[31440];
assign g[47825] = a[14] & g[31441];
assign g[64208] = b[14] & g[31441];
assign g[47826] = a[14] & g[31442];
assign g[64209] = b[14] & g[31442];
assign g[47827] = a[14] & g[31443];
assign g[64210] = b[14] & g[31443];
assign g[47828] = a[14] & g[31444];
assign g[64211] = b[14] & g[31444];
assign g[47829] = a[14] & g[31445];
assign g[64212] = b[14] & g[31445];
assign g[47830] = a[14] & g[31446];
assign g[64213] = b[14] & g[31446];
assign g[47831] = a[14] & g[31447];
assign g[64214] = b[14] & g[31447];
assign g[47832] = a[14] & g[31448];
assign g[64215] = b[14] & g[31448];
assign g[47833] = a[14] & g[31449];
assign g[64216] = b[14] & g[31449];
assign g[47834] = a[14] & g[31450];
assign g[64217] = b[14] & g[31450];
assign g[47835] = a[14] & g[31451];
assign g[64218] = b[14] & g[31451];
assign g[47836] = a[14] & g[31452];
assign g[64219] = b[14] & g[31452];
assign g[47837] = a[14] & g[31453];
assign g[64220] = b[14] & g[31453];
assign g[47838] = a[14] & g[31454];
assign g[64221] = b[14] & g[31454];
assign g[47839] = a[14] & g[31455];
assign g[64222] = b[14] & g[31455];
assign g[47840] = a[14] & g[31456];
assign g[64223] = b[14] & g[31456];
assign g[47841] = a[14] & g[31457];
assign g[64224] = b[14] & g[31457];
assign g[47842] = a[14] & g[31458];
assign g[64225] = b[14] & g[31458];
assign g[47843] = a[14] & g[31459];
assign g[64226] = b[14] & g[31459];
assign g[47844] = a[14] & g[31460];
assign g[64227] = b[14] & g[31460];
assign g[47845] = a[14] & g[31461];
assign g[64228] = b[14] & g[31461];
assign g[47846] = a[14] & g[31462];
assign g[64229] = b[14] & g[31462];
assign g[47847] = a[14] & g[31463];
assign g[64230] = b[14] & g[31463];
assign g[47848] = a[14] & g[31464];
assign g[64231] = b[14] & g[31464];
assign g[47849] = a[14] & g[31465];
assign g[64232] = b[14] & g[31465];
assign g[47850] = a[14] & g[31466];
assign g[64233] = b[14] & g[31466];
assign g[47851] = a[14] & g[31467];
assign g[64234] = b[14] & g[31467];
assign g[47852] = a[14] & g[31468];
assign g[64235] = b[14] & g[31468];
assign g[47853] = a[14] & g[31469];
assign g[64236] = b[14] & g[31469];
assign g[47854] = a[14] & g[31470];
assign g[64237] = b[14] & g[31470];
assign g[47855] = a[14] & g[31471];
assign g[64238] = b[14] & g[31471];
assign g[47856] = a[14] & g[31472];
assign g[64239] = b[14] & g[31472];
assign g[47857] = a[14] & g[31473];
assign g[64240] = b[14] & g[31473];
assign g[47858] = a[14] & g[31474];
assign g[64241] = b[14] & g[31474];
assign g[47859] = a[14] & g[31475];
assign g[64242] = b[14] & g[31475];
assign g[47860] = a[14] & g[31476];
assign g[64243] = b[14] & g[31476];
assign g[47861] = a[14] & g[31477];
assign g[64244] = b[14] & g[31477];
assign g[47862] = a[14] & g[31478];
assign g[64245] = b[14] & g[31478];
assign g[47863] = a[14] & g[31479];
assign g[64246] = b[14] & g[31479];
assign g[47864] = a[14] & g[31480];
assign g[64247] = b[14] & g[31480];
assign g[47865] = a[14] & g[31481];
assign g[64248] = b[14] & g[31481];
assign g[47866] = a[14] & g[31482];
assign g[64249] = b[14] & g[31482];
assign g[47867] = a[14] & g[31483];
assign g[64250] = b[14] & g[31483];
assign g[47868] = a[14] & g[31484];
assign g[64251] = b[14] & g[31484];
assign g[47869] = a[14] & g[31485];
assign g[64252] = b[14] & g[31485];
assign g[47870] = a[14] & g[31486];
assign g[64253] = b[14] & g[31486];
assign g[47871] = a[14] & g[31487];
assign g[64254] = b[14] & g[31487];
assign g[47872] = a[14] & g[31488];
assign g[64255] = b[14] & g[31488];
assign g[47873] = a[14] & g[31489];
assign g[64256] = b[14] & g[31489];
assign g[47874] = a[14] & g[31490];
assign g[64257] = b[14] & g[31490];
assign g[47875] = a[14] & g[31491];
assign g[64258] = b[14] & g[31491];
assign g[47876] = a[14] & g[31492];
assign g[64259] = b[14] & g[31492];
assign g[47877] = a[14] & g[31493];
assign g[64260] = b[14] & g[31493];
assign g[47878] = a[14] & g[31494];
assign g[64261] = b[14] & g[31494];
assign g[47879] = a[14] & g[31495];
assign g[64262] = b[14] & g[31495];
assign g[47880] = a[14] & g[31496];
assign g[64263] = b[14] & g[31496];
assign g[47881] = a[14] & g[31497];
assign g[64264] = b[14] & g[31497];
assign g[47882] = a[14] & g[31498];
assign g[64265] = b[14] & g[31498];
assign g[47883] = a[14] & g[31499];
assign g[64266] = b[14] & g[31499];
assign g[47884] = a[14] & g[31500];
assign g[64267] = b[14] & g[31500];
assign g[47885] = a[14] & g[31501];
assign g[64268] = b[14] & g[31501];
assign g[47886] = a[14] & g[31502];
assign g[64269] = b[14] & g[31502];
assign g[47887] = a[14] & g[31503];
assign g[64270] = b[14] & g[31503];
assign g[47888] = a[14] & g[31504];
assign g[64271] = b[14] & g[31504];
assign g[47889] = a[14] & g[31505];
assign g[64272] = b[14] & g[31505];
assign g[47890] = a[14] & g[31506];
assign g[64273] = b[14] & g[31506];
assign g[47891] = a[14] & g[31507];
assign g[64274] = b[14] & g[31507];
assign g[47892] = a[14] & g[31508];
assign g[64275] = b[14] & g[31508];
assign g[47893] = a[14] & g[31509];
assign g[64276] = b[14] & g[31509];
assign g[47894] = a[14] & g[31510];
assign g[64277] = b[14] & g[31510];
assign g[47895] = a[14] & g[31511];
assign g[64278] = b[14] & g[31511];
assign g[47896] = a[14] & g[31512];
assign g[64279] = b[14] & g[31512];
assign g[47897] = a[14] & g[31513];
assign g[64280] = b[14] & g[31513];
assign g[47898] = a[14] & g[31514];
assign g[64281] = b[14] & g[31514];
assign g[47899] = a[14] & g[31515];
assign g[64282] = b[14] & g[31515];
assign g[47900] = a[14] & g[31516];
assign g[64283] = b[14] & g[31516];
assign g[47901] = a[14] & g[31517];
assign g[64284] = b[14] & g[31517];
assign g[47902] = a[14] & g[31518];
assign g[64285] = b[14] & g[31518];
assign g[47903] = a[14] & g[31519];
assign g[64286] = b[14] & g[31519];
assign g[47904] = a[14] & g[31520];
assign g[64287] = b[14] & g[31520];
assign g[47905] = a[14] & g[31521];
assign g[64288] = b[14] & g[31521];
assign g[47906] = a[14] & g[31522];
assign g[64289] = b[14] & g[31522];
assign g[47907] = a[14] & g[31523];
assign g[64290] = b[14] & g[31523];
assign g[47908] = a[14] & g[31524];
assign g[64291] = b[14] & g[31524];
assign g[47909] = a[14] & g[31525];
assign g[64292] = b[14] & g[31525];
assign g[47910] = a[14] & g[31526];
assign g[64293] = b[14] & g[31526];
assign g[47911] = a[14] & g[31527];
assign g[64294] = b[14] & g[31527];
assign g[47912] = a[14] & g[31528];
assign g[64295] = b[14] & g[31528];
assign g[47913] = a[14] & g[31529];
assign g[64296] = b[14] & g[31529];
assign g[47914] = a[14] & g[31530];
assign g[64297] = b[14] & g[31530];
assign g[47915] = a[14] & g[31531];
assign g[64298] = b[14] & g[31531];
assign g[47916] = a[14] & g[31532];
assign g[64299] = b[14] & g[31532];
assign g[47917] = a[14] & g[31533];
assign g[64300] = b[14] & g[31533];
assign g[47918] = a[14] & g[31534];
assign g[64301] = b[14] & g[31534];
assign g[47919] = a[14] & g[31535];
assign g[64302] = b[14] & g[31535];
assign g[47920] = a[14] & g[31536];
assign g[64303] = b[14] & g[31536];
assign g[47921] = a[14] & g[31537];
assign g[64304] = b[14] & g[31537];
assign g[47922] = a[14] & g[31538];
assign g[64305] = b[14] & g[31538];
assign g[47923] = a[14] & g[31539];
assign g[64306] = b[14] & g[31539];
assign g[47924] = a[14] & g[31540];
assign g[64307] = b[14] & g[31540];
assign g[47925] = a[14] & g[31541];
assign g[64308] = b[14] & g[31541];
assign g[47926] = a[14] & g[31542];
assign g[64309] = b[14] & g[31542];
assign g[47927] = a[14] & g[31543];
assign g[64310] = b[14] & g[31543];
assign g[47928] = a[14] & g[31544];
assign g[64311] = b[14] & g[31544];
assign g[47929] = a[14] & g[31545];
assign g[64312] = b[14] & g[31545];
assign g[47930] = a[14] & g[31546];
assign g[64313] = b[14] & g[31546];
assign g[47931] = a[14] & g[31547];
assign g[64314] = b[14] & g[31547];
assign g[47932] = a[14] & g[31548];
assign g[64315] = b[14] & g[31548];
assign g[47933] = a[14] & g[31549];
assign g[64316] = b[14] & g[31549];
assign g[47934] = a[14] & g[31550];
assign g[64317] = b[14] & g[31550];
assign g[47935] = a[14] & g[31551];
assign g[64318] = b[14] & g[31551];
assign g[47936] = a[14] & g[31552];
assign g[64319] = b[14] & g[31552];
assign g[47937] = a[14] & g[31553];
assign g[64320] = b[14] & g[31553];
assign g[47938] = a[14] & g[31554];
assign g[64321] = b[14] & g[31554];
assign g[47939] = a[14] & g[31555];
assign g[64322] = b[14] & g[31555];
assign g[47940] = a[14] & g[31556];
assign g[64323] = b[14] & g[31556];
assign g[47941] = a[14] & g[31557];
assign g[64324] = b[14] & g[31557];
assign g[47942] = a[14] & g[31558];
assign g[64325] = b[14] & g[31558];
assign g[47943] = a[14] & g[31559];
assign g[64326] = b[14] & g[31559];
assign g[47944] = a[14] & g[31560];
assign g[64327] = b[14] & g[31560];
assign g[47945] = a[14] & g[31561];
assign g[64328] = b[14] & g[31561];
assign g[47946] = a[14] & g[31562];
assign g[64329] = b[14] & g[31562];
assign g[47947] = a[14] & g[31563];
assign g[64330] = b[14] & g[31563];
assign g[47948] = a[14] & g[31564];
assign g[64331] = b[14] & g[31564];
assign g[47949] = a[14] & g[31565];
assign g[64332] = b[14] & g[31565];
assign g[47950] = a[14] & g[31566];
assign g[64333] = b[14] & g[31566];
assign g[47951] = a[14] & g[31567];
assign g[64334] = b[14] & g[31567];
assign g[47952] = a[14] & g[31568];
assign g[64335] = b[14] & g[31568];
assign g[47953] = a[14] & g[31569];
assign g[64336] = b[14] & g[31569];
assign g[47954] = a[14] & g[31570];
assign g[64337] = b[14] & g[31570];
assign g[47955] = a[14] & g[31571];
assign g[64338] = b[14] & g[31571];
assign g[47956] = a[14] & g[31572];
assign g[64339] = b[14] & g[31572];
assign g[47957] = a[14] & g[31573];
assign g[64340] = b[14] & g[31573];
assign g[47958] = a[14] & g[31574];
assign g[64341] = b[14] & g[31574];
assign g[47959] = a[14] & g[31575];
assign g[64342] = b[14] & g[31575];
assign g[47960] = a[14] & g[31576];
assign g[64343] = b[14] & g[31576];
assign g[47961] = a[14] & g[31577];
assign g[64344] = b[14] & g[31577];
assign g[47962] = a[14] & g[31578];
assign g[64345] = b[14] & g[31578];
assign g[47963] = a[14] & g[31579];
assign g[64346] = b[14] & g[31579];
assign g[47964] = a[14] & g[31580];
assign g[64347] = b[14] & g[31580];
assign g[47965] = a[14] & g[31581];
assign g[64348] = b[14] & g[31581];
assign g[47966] = a[14] & g[31582];
assign g[64349] = b[14] & g[31582];
assign g[47967] = a[14] & g[31583];
assign g[64350] = b[14] & g[31583];
assign g[47968] = a[14] & g[31584];
assign g[64351] = b[14] & g[31584];
assign g[47969] = a[14] & g[31585];
assign g[64352] = b[14] & g[31585];
assign g[47970] = a[14] & g[31586];
assign g[64353] = b[14] & g[31586];
assign g[47971] = a[14] & g[31587];
assign g[64354] = b[14] & g[31587];
assign g[47972] = a[14] & g[31588];
assign g[64355] = b[14] & g[31588];
assign g[47973] = a[14] & g[31589];
assign g[64356] = b[14] & g[31589];
assign g[47974] = a[14] & g[31590];
assign g[64357] = b[14] & g[31590];
assign g[47975] = a[14] & g[31591];
assign g[64358] = b[14] & g[31591];
assign g[47976] = a[14] & g[31592];
assign g[64359] = b[14] & g[31592];
assign g[47977] = a[14] & g[31593];
assign g[64360] = b[14] & g[31593];
assign g[47978] = a[14] & g[31594];
assign g[64361] = b[14] & g[31594];
assign g[47979] = a[14] & g[31595];
assign g[64362] = b[14] & g[31595];
assign g[47980] = a[14] & g[31596];
assign g[64363] = b[14] & g[31596];
assign g[47981] = a[14] & g[31597];
assign g[64364] = b[14] & g[31597];
assign g[47982] = a[14] & g[31598];
assign g[64365] = b[14] & g[31598];
assign g[47983] = a[14] & g[31599];
assign g[64366] = b[14] & g[31599];
assign g[47984] = a[14] & g[31600];
assign g[64367] = b[14] & g[31600];
assign g[47985] = a[14] & g[31601];
assign g[64368] = b[14] & g[31601];
assign g[47986] = a[14] & g[31602];
assign g[64369] = b[14] & g[31602];
assign g[47987] = a[14] & g[31603];
assign g[64370] = b[14] & g[31603];
assign g[47988] = a[14] & g[31604];
assign g[64371] = b[14] & g[31604];
assign g[47989] = a[14] & g[31605];
assign g[64372] = b[14] & g[31605];
assign g[47990] = a[14] & g[31606];
assign g[64373] = b[14] & g[31606];
assign g[47991] = a[14] & g[31607];
assign g[64374] = b[14] & g[31607];
assign g[47992] = a[14] & g[31608];
assign g[64375] = b[14] & g[31608];
assign g[47993] = a[14] & g[31609];
assign g[64376] = b[14] & g[31609];
assign g[47994] = a[14] & g[31610];
assign g[64377] = b[14] & g[31610];
assign g[47995] = a[14] & g[31611];
assign g[64378] = b[14] & g[31611];
assign g[47996] = a[14] & g[31612];
assign g[64379] = b[14] & g[31612];
assign g[47997] = a[14] & g[31613];
assign g[64380] = b[14] & g[31613];
assign g[47998] = a[14] & g[31614];
assign g[64381] = b[14] & g[31614];
assign g[47999] = a[14] & g[31615];
assign g[64382] = b[14] & g[31615];
assign g[48000] = a[14] & g[31616];
assign g[64383] = b[14] & g[31616];
assign g[48001] = a[14] & g[31617];
assign g[64384] = b[14] & g[31617];
assign g[48002] = a[14] & g[31618];
assign g[64385] = b[14] & g[31618];
assign g[48003] = a[14] & g[31619];
assign g[64386] = b[14] & g[31619];
assign g[48004] = a[14] & g[31620];
assign g[64387] = b[14] & g[31620];
assign g[48005] = a[14] & g[31621];
assign g[64388] = b[14] & g[31621];
assign g[48006] = a[14] & g[31622];
assign g[64389] = b[14] & g[31622];
assign g[48007] = a[14] & g[31623];
assign g[64390] = b[14] & g[31623];
assign g[48008] = a[14] & g[31624];
assign g[64391] = b[14] & g[31624];
assign g[48009] = a[14] & g[31625];
assign g[64392] = b[14] & g[31625];
assign g[48010] = a[14] & g[31626];
assign g[64393] = b[14] & g[31626];
assign g[48011] = a[14] & g[31627];
assign g[64394] = b[14] & g[31627];
assign g[48012] = a[14] & g[31628];
assign g[64395] = b[14] & g[31628];
assign g[48013] = a[14] & g[31629];
assign g[64396] = b[14] & g[31629];
assign g[48014] = a[14] & g[31630];
assign g[64397] = b[14] & g[31630];
assign g[48015] = a[14] & g[31631];
assign g[64398] = b[14] & g[31631];
assign g[48016] = a[14] & g[31632];
assign g[64399] = b[14] & g[31632];
assign g[48017] = a[14] & g[31633];
assign g[64400] = b[14] & g[31633];
assign g[48018] = a[14] & g[31634];
assign g[64401] = b[14] & g[31634];
assign g[48019] = a[14] & g[31635];
assign g[64402] = b[14] & g[31635];
assign g[48020] = a[14] & g[31636];
assign g[64403] = b[14] & g[31636];
assign g[48021] = a[14] & g[31637];
assign g[64404] = b[14] & g[31637];
assign g[48022] = a[14] & g[31638];
assign g[64405] = b[14] & g[31638];
assign g[48023] = a[14] & g[31639];
assign g[64406] = b[14] & g[31639];
assign g[48024] = a[14] & g[31640];
assign g[64407] = b[14] & g[31640];
assign g[48025] = a[14] & g[31641];
assign g[64408] = b[14] & g[31641];
assign g[48026] = a[14] & g[31642];
assign g[64409] = b[14] & g[31642];
assign g[48027] = a[14] & g[31643];
assign g[64410] = b[14] & g[31643];
assign g[48028] = a[14] & g[31644];
assign g[64411] = b[14] & g[31644];
assign g[48029] = a[14] & g[31645];
assign g[64412] = b[14] & g[31645];
assign g[48030] = a[14] & g[31646];
assign g[64413] = b[14] & g[31646];
assign g[48031] = a[14] & g[31647];
assign g[64414] = b[14] & g[31647];
assign g[48032] = a[14] & g[31648];
assign g[64415] = b[14] & g[31648];
assign g[48033] = a[14] & g[31649];
assign g[64416] = b[14] & g[31649];
assign g[48034] = a[14] & g[31650];
assign g[64417] = b[14] & g[31650];
assign g[48035] = a[14] & g[31651];
assign g[64418] = b[14] & g[31651];
assign g[48036] = a[14] & g[31652];
assign g[64419] = b[14] & g[31652];
assign g[48037] = a[14] & g[31653];
assign g[64420] = b[14] & g[31653];
assign g[48038] = a[14] & g[31654];
assign g[64421] = b[14] & g[31654];
assign g[48039] = a[14] & g[31655];
assign g[64422] = b[14] & g[31655];
assign g[48040] = a[14] & g[31656];
assign g[64423] = b[14] & g[31656];
assign g[48041] = a[14] & g[31657];
assign g[64424] = b[14] & g[31657];
assign g[48042] = a[14] & g[31658];
assign g[64425] = b[14] & g[31658];
assign g[48043] = a[14] & g[31659];
assign g[64426] = b[14] & g[31659];
assign g[48044] = a[14] & g[31660];
assign g[64427] = b[14] & g[31660];
assign g[48045] = a[14] & g[31661];
assign g[64428] = b[14] & g[31661];
assign g[48046] = a[14] & g[31662];
assign g[64429] = b[14] & g[31662];
assign g[48047] = a[14] & g[31663];
assign g[64430] = b[14] & g[31663];
assign g[48048] = a[14] & g[31664];
assign g[64431] = b[14] & g[31664];
assign g[48049] = a[14] & g[31665];
assign g[64432] = b[14] & g[31665];
assign g[48050] = a[14] & g[31666];
assign g[64433] = b[14] & g[31666];
assign g[48051] = a[14] & g[31667];
assign g[64434] = b[14] & g[31667];
assign g[48052] = a[14] & g[31668];
assign g[64435] = b[14] & g[31668];
assign g[48053] = a[14] & g[31669];
assign g[64436] = b[14] & g[31669];
assign g[48054] = a[14] & g[31670];
assign g[64437] = b[14] & g[31670];
assign g[48055] = a[14] & g[31671];
assign g[64438] = b[14] & g[31671];
assign g[48056] = a[14] & g[31672];
assign g[64439] = b[14] & g[31672];
assign g[48057] = a[14] & g[31673];
assign g[64440] = b[14] & g[31673];
assign g[48058] = a[14] & g[31674];
assign g[64441] = b[14] & g[31674];
assign g[48059] = a[14] & g[31675];
assign g[64442] = b[14] & g[31675];
assign g[48060] = a[14] & g[31676];
assign g[64443] = b[14] & g[31676];
assign g[48061] = a[14] & g[31677];
assign g[64444] = b[14] & g[31677];
assign g[48062] = a[14] & g[31678];
assign g[64445] = b[14] & g[31678];
assign g[48063] = a[14] & g[31679];
assign g[64446] = b[14] & g[31679];
assign g[48064] = a[14] & g[31680];
assign g[64447] = b[14] & g[31680];
assign g[48065] = a[14] & g[31681];
assign g[64448] = b[14] & g[31681];
assign g[48066] = a[14] & g[31682];
assign g[64449] = b[14] & g[31682];
assign g[48067] = a[14] & g[31683];
assign g[64450] = b[14] & g[31683];
assign g[48068] = a[14] & g[31684];
assign g[64451] = b[14] & g[31684];
assign g[48069] = a[14] & g[31685];
assign g[64452] = b[14] & g[31685];
assign g[48070] = a[14] & g[31686];
assign g[64453] = b[14] & g[31686];
assign g[48071] = a[14] & g[31687];
assign g[64454] = b[14] & g[31687];
assign g[48072] = a[14] & g[31688];
assign g[64455] = b[14] & g[31688];
assign g[48073] = a[14] & g[31689];
assign g[64456] = b[14] & g[31689];
assign g[48074] = a[14] & g[31690];
assign g[64457] = b[14] & g[31690];
assign g[48075] = a[14] & g[31691];
assign g[64458] = b[14] & g[31691];
assign g[48076] = a[14] & g[31692];
assign g[64459] = b[14] & g[31692];
assign g[48077] = a[14] & g[31693];
assign g[64460] = b[14] & g[31693];
assign g[48078] = a[14] & g[31694];
assign g[64461] = b[14] & g[31694];
assign g[48079] = a[14] & g[31695];
assign g[64462] = b[14] & g[31695];
assign g[48080] = a[14] & g[31696];
assign g[64463] = b[14] & g[31696];
assign g[48081] = a[14] & g[31697];
assign g[64464] = b[14] & g[31697];
assign g[48082] = a[14] & g[31698];
assign g[64465] = b[14] & g[31698];
assign g[48083] = a[14] & g[31699];
assign g[64466] = b[14] & g[31699];
assign g[48084] = a[14] & g[31700];
assign g[64467] = b[14] & g[31700];
assign g[48085] = a[14] & g[31701];
assign g[64468] = b[14] & g[31701];
assign g[48086] = a[14] & g[31702];
assign g[64469] = b[14] & g[31702];
assign g[48087] = a[14] & g[31703];
assign g[64470] = b[14] & g[31703];
assign g[48088] = a[14] & g[31704];
assign g[64471] = b[14] & g[31704];
assign g[48089] = a[14] & g[31705];
assign g[64472] = b[14] & g[31705];
assign g[48090] = a[14] & g[31706];
assign g[64473] = b[14] & g[31706];
assign g[48091] = a[14] & g[31707];
assign g[64474] = b[14] & g[31707];
assign g[48092] = a[14] & g[31708];
assign g[64475] = b[14] & g[31708];
assign g[48093] = a[14] & g[31709];
assign g[64476] = b[14] & g[31709];
assign g[48094] = a[14] & g[31710];
assign g[64477] = b[14] & g[31710];
assign g[48095] = a[14] & g[31711];
assign g[64478] = b[14] & g[31711];
assign g[48096] = a[14] & g[31712];
assign g[64479] = b[14] & g[31712];
assign g[48097] = a[14] & g[31713];
assign g[64480] = b[14] & g[31713];
assign g[48098] = a[14] & g[31714];
assign g[64481] = b[14] & g[31714];
assign g[48099] = a[14] & g[31715];
assign g[64482] = b[14] & g[31715];
assign g[48100] = a[14] & g[31716];
assign g[64483] = b[14] & g[31716];
assign g[48101] = a[14] & g[31717];
assign g[64484] = b[14] & g[31717];
assign g[48102] = a[14] & g[31718];
assign g[64485] = b[14] & g[31718];
assign g[48103] = a[14] & g[31719];
assign g[64486] = b[14] & g[31719];
assign g[48104] = a[14] & g[31720];
assign g[64487] = b[14] & g[31720];
assign g[48105] = a[14] & g[31721];
assign g[64488] = b[14] & g[31721];
assign g[48106] = a[14] & g[31722];
assign g[64489] = b[14] & g[31722];
assign g[48107] = a[14] & g[31723];
assign g[64490] = b[14] & g[31723];
assign g[48108] = a[14] & g[31724];
assign g[64491] = b[14] & g[31724];
assign g[48109] = a[14] & g[31725];
assign g[64492] = b[14] & g[31725];
assign g[48110] = a[14] & g[31726];
assign g[64493] = b[14] & g[31726];
assign g[48111] = a[14] & g[31727];
assign g[64494] = b[14] & g[31727];
assign g[48112] = a[14] & g[31728];
assign g[64495] = b[14] & g[31728];
assign g[48113] = a[14] & g[31729];
assign g[64496] = b[14] & g[31729];
assign g[48114] = a[14] & g[31730];
assign g[64497] = b[14] & g[31730];
assign g[48115] = a[14] & g[31731];
assign g[64498] = b[14] & g[31731];
assign g[48116] = a[14] & g[31732];
assign g[64499] = b[14] & g[31732];
assign g[48117] = a[14] & g[31733];
assign g[64500] = b[14] & g[31733];
assign g[48118] = a[14] & g[31734];
assign g[64501] = b[14] & g[31734];
assign g[48119] = a[14] & g[31735];
assign g[64502] = b[14] & g[31735];
assign g[48120] = a[14] & g[31736];
assign g[64503] = b[14] & g[31736];
assign g[48121] = a[14] & g[31737];
assign g[64504] = b[14] & g[31737];
assign g[48122] = a[14] & g[31738];
assign g[64505] = b[14] & g[31738];
assign g[48123] = a[14] & g[31739];
assign g[64506] = b[14] & g[31739];
assign g[48124] = a[14] & g[31740];
assign g[64507] = b[14] & g[31740];
assign g[48125] = a[14] & g[31741];
assign g[64508] = b[14] & g[31741];
assign g[48126] = a[14] & g[31742];
assign g[64509] = b[14] & g[31742];
assign g[48127] = a[14] & g[31743];
assign g[64510] = b[14] & g[31743];
assign g[48128] = a[14] & g[31744];
assign g[64511] = b[14] & g[31744];
assign g[48129] = a[14] & g[31745];
assign g[64512] = b[14] & g[31745];
assign g[48130] = a[14] & g[31746];
assign g[64513] = b[14] & g[31746];
assign g[48131] = a[14] & g[31747];
assign g[64514] = b[14] & g[31747];
assign g[48132] = a[14] & g[31748];
assign g[64515] = b[14] & g[31748];
assign g[48133] = a[14] & g[31749];
assign g[64516] = b[14] & g[31749];
assign g[48134] = a[14] & g[31750];
assign g[64517] = b[14] & g[31750];
assign g[48135] = a[14] & g[31751];
assign g[64518] = b[14] & g[31751];
assign g[48136] = a[14] & g[31752];
assign g[64519] = b[14] & g[31752];
assign g[48137] = a[14] & g[31753];
assign g[64520] = b[14] & g[31753];
assign g[48138] = a[14] & g[31754];
assign g[64521] = b[14] & g[31754];
assign g[48139] = a[14] & g[31755];
assign g[64522] = b[14] & g[31755];
assign g[48140] = a[14] & g[31756];
assign g[64523] = b[14] & g[31756];
assign g[48141] = a[14] & g[31757];
assign g[64524] = b[14] & g[31757];
assign g[48142] = a[14] & g[31758];
assign g[64525] = b[14] & g[31758];
assign g[48143] = a[14] & g[31759];
assign g[64526] = b[14] & g[31759];
assign g[48144] = a[14] & g[31760];
assign g[64527] = b[14] & g[31760];
assign g[48145] = a[14] & g[31761];
assign g[64528] = b[14] & g[31761];
assign g[48146] = a[14] & g[31762];
assign g[64529] = b[14] & g[31762];
assign g[48147] = a[14] & g[31763];
assign g[64530] = b[14] & g[31763];
assign g[48148] = a[14] & g[31764];
assign g[64531] = b[14] & g[31764];
assign g[48149] = a[14] & g[31765];
assign g[64532] = b[14] & g[31765];
assign g[48150] = a[14] & g[31766];
assign g[64533] = b[14] & g[31766];
assign g[48151] = a[14] & g[31767];
assign g[64534] = b[14] & g[31767];
assign g[48152] = a[14] & g[31768];
assign g[64535] = b[14] & g[31768];
assign g[48153] = a[14] & g[31769];
assign g[64536] = b[14] & g[31769];
assign g[48154] = a[14] & g[31770];
assign g[64537] = b[14] & g[31770];
assign g[48155] = a[14] & g[31771];
assign g[64538] = b[14] & g[31771];
assign g[48156] = a[14] & g[31772];
assign g[64539] = b[14] & g[31772];
assign g[48157] = a[14] & g[31773];
assign g[64540] = b[14] & g[31773];
assign g[48158] = a[14] & g[31774];
assign g[64541] = b[14] & g[31774];
assign g[48159] = a[14] & g[31775];
assign g[64542] = b[14] & g[31775];
assign g[48160] = a[14] & g[31776];
assign g[64543] = b[14] & g[31776];
assign g[48161] = a[14] & g[31777];
assign g[64544] = b[14] & g[31777];
assign g[48162] = a[14] & g[31778];
assign g[64545] = b[14] & g[31778];
assign g[48163] = a[14] & g[31779];
assign g[64546] = b[14] & g[31779];
assign g[48164] = a[14] & g[31780];
assign g[64547] = b[14] & g[31780];
assign g[48165] = a[14] & g[31781];
assign g[64548] = b[14] & g[31781];
assign g[48166] = a[14] & g[31782];
assign g[64549] = b[14] & g[31782];
assign g[48167] = a[14] & g[31783];
assign g[64550] = b[14] & g[31783];
assign g[48168] = a[14] & g[31784];
assign g[64551] = b[14] & g[31784];
assign g[48169] = a[14] & g[31785];
assign g[64552] = b[14] & g[31785];
assign g[48170] = a[14] & g[31786];
assign g[64553] = b[14] & g[31786];
assign g[48171] = a[14] & g[31787];
assign g[64554] = b[14] & g[31787];
assign g[48172] = a[14] & g[31788];
assign g[64555] = b[14] & g[31788];
assign g[48173] = a[14] & g[31789];
assign g[64556] = b[14] & g[31789];
assign g[48174] = a[14] & g[31790];
assign g[64557] = b[14] & g[31790];
assign g[48175] = a[14] & g[31791];
assign g[64558] = b[14] & g[31791];
assign g[48176] = a[14] & g[31792];
assign g[64559] = b[14] & g[31792];
assign g[48177] = a[14] & g[31793];
assign g[64560] = b[14] & g[31793];
assign g[48178] = a[14] & g[31794];
assign g[64561] = b[14] & g[31794];
assign g[48179] = a[14] & g[31795];
assign g[64562] = b[14] & g[31795];
assign g[48180] = a[14] & g[31796];
assign g[64563] = b[14] & g[31796];
assign g[48181] = a[14] & g[31797];
assign g[64564] = b[14] & g[31797];
assign g[48182] = a[14] & g[31798];
assign g[64565] = b[14] & g[31798];
assign g[48183] = a[14] & g[31799];
assign g[64566] = b[14] & g[31799];
assign g[48184] = a[14] & g[31800];
assign g[64567] = b[14] & g[31800];
assign g[48185] = a[14] & g[31801];
assign g[64568] = b[14] & g[31801];
assign g[48186] = a[14] & g[31802];
assign g[64569] = b[14] & g[31802];
assign g[48187] = a[14] & g[31803];
assign g[64570] = b[14] & g[31803];
assign g[48188] = a[14] & g[31804];
assign g[64571] = b[14] & g[31804];
assign g[48189] = a[14] & g[31805];
assign g[64572] = b[14] & g[31805];
assign g[48190] = a[14] & g[31806];
assign g[64573] = b[14] & g[31806];
assign g[48191] = a[14] & g[31807];
assign g[64574] = b[14] & g[31807];
assign g[48192] = a[14] & g[31808];
assign g[64575] = b[14] & g[31808];
assign g[48193] = a[14] & g[31809];
assign g[64576] = b[14] & g[31809];
assign g[48194] = a[14] & g[31810];
assign g[64577] = b[14] & g[31810];
assign g[48195] = a[14] & g[31811];
assign g[64578] = b[14] & g[31811];
assign g[48196] = a[14] & g[31812];
assign g[64579] = b[14] & g[31812];
assign g[48197] = a[14] & g[31813];
assign g[64580] = b[14] & g[31813];
assign g[48198] = a[14] & g[31814];
assign g[64581] = b[14] & g[31814];
assign g[48199] = a[14] & g[31815];
assign g[64582] = b[14] & g[31815];
assign g[48200] = a[14] & g[31816];
assign g[64583] = b[14] & g[31816];
assign g[48201] = a[14] & g[31817];
assign g[64584] = b[14] & g[31817];
assign g[48202] = a[14] & g[31818];
assign g[64585] = b[14] & g[31818];
assign g[48203] = a[14] & g[31819];
assign g[64586] = b[14] & g[31819];
assign g[48204] = a[14] & g[31820];
assign g[64587] = b[14] & g[31820];
assign g[48205] = a[14] & g[31821];
assign g[64588] = b[14] & g[31821];
assign g[48206] = a[14] & g[31822];
assign g[64589] = b[14] & g[31822];
assign g[48207] = a[14] & g[31823];
assign g[64590] = b[14] & g[31823];
assign g[48208] = a[14] & g[31824];
assign g[64591] = b[14] & g[31824];
assign g[48209] = a[14] & g[31825];
assign g[64592] = b[14] & g[31825];
assign g[48210] = a[14] & g[31826];
assign g[64593] = b[14] & g[31826];
assign g[48211] = a[14] & g[31827];
assign g[64594] = b[14] & g[31827];
assign g[48212] = a[14] & g[31828];
assign g[64595] = b[14] & g[31828];
assign g[48213] = a[14] & g[31829];
assign g[64596] = b[14] & g[31829];
assign g[48214] = a[14] & g[31830];
assign g[64597] = b[14] & g[31830];
assign g[48215] = a[14] & g[31831];
assign g[64598] = b[14] & g[31831];
assign g[48216] = a[14] & g[31832];
assign g[64599] = b[14] & g[31832];
assign g[48217] = a[14] & g[31833];
assign g[64600] = b[14] & g[31833];
assign g[48218] = a[14] & g[31834];
assign g[64601] = b[14] & g[31834];
assign g[48219] = a[14] & g[31835];
assign g[64602] = b[14] & g[31835];
assign g[48220] = a[14] & g[31836];
assign g[64603] = b[14] & g[31836];
assign g[48221] = a[14] & g[31837];
assign g[64604] = b[14] & g[31837];
assign g[48222] = a[14] & g[31838];
assign g[64605] = b[14] & g[31838];
assign g[48223] = a[14] & g[31839];
assign g[64606] = b[14] & g[31839];
assign g[48224] = a[14] & g[31840];
assign g[64607] = b[14] & g[31840];
assign g[48225] = a[14] & g[31841];
assign g[64608] = b[14] & g[31841];
assign g[48226] = a[14] & g[31842];
assign g[64609] = b[14] & g[31842];
assign g[48227] = a[14] & g[31843];
assign g[64610] = b[14] & g[31843];
assign g[48228] = a[14] & g[31844];
assign g[64611] = b[14] & g[31844];
assign g[48229] = a[14] & g[31845];
assign g[64612] = b[14] & g[31845];
assign g[48230] = a[14] & g[31846];
assign g[64613] = b[14] & g[31846];
assign g[48231] = a[14] & g[31847];
assign g[64614] = b[14] & g[31847];
assign g[48232] = a[14] & g[31848];
assign g[64615] = b[14] & g[31848];
assign g[48233] = a[14] & g[31849];
assign g[64616] = b[14] & g[31849];
assign g[48234] = a[14] & g[31850];
assign g[64617] = b[14] & g[31850];
assign g[48235] = a[14] & g[31851];
assign g[64618] = b[14] & g[31851];
assign g[48236] = a[14] & g[31852];
assign g[64619] = b[14] & g[31852];
assign g[48237] = a[14] & g[31853];
assign g[64620] = b[14] & g[31853];
assign g[48238] = a[14] & g[31854];
assign g[64621] = b[14] & g[31854];
assign g[48239] = a[14] & g[31855];
assign g[64622] = b[14] & g[31855];
assign g[48240] = a[14] & g[31856];
assign g[64623] = b[14] & g[31856];
assign g[48241] = a[14] & g[31857];
assign g[64624] = b[14] & g[31857];
assign g[48242] = a[14] & g[31858];
assign g[64625] = b[14] & g[31858];
assign g[48243] = a[14] & g[31859];
assign g[64626] = b[14] & g[31859];
assign g[48244] = a[14] & g[31860];
assign g[64627] = b[14] & g[31860];
assign g[48245] = a[14] & g[31861];
assign g[64628] = b[14] & g[31861];
assign g[48246] = a[14] & g[31862];
assign g[64629] = b[14] & g[31862];
assign g[48247] = a[14] & g[31863];
assign g[64630] = b[14] & g[31863];
assign g[48248] = a[14] & g[31864];
assign g[64631] = b[14] & g[31864];
assign g[48249] = a[14] & g[31865];
assign g[64632] = b[14] & g[31865];
assign g[48250] = a[14] & g[31866];
assign g[64633] = b[14] & g[31866];
assign g[48251] = a[14] & g[31867];
assign g[64634] = b[14] & g[31867];
assign g[48252] = a[14] & g[31868];
assign g[64635] = b[14] & g[31868];
assign g[48253] = a[14] & g[31869];
assign g[64636] = b[14] & g[31869];
assign g[48254] = a[14] & g[31870];
assign g[64637] = b[14] & g[31870];
assign g[48255] = a[14] & g[31871];
assign g[64638] = b[14] & g[31871];
assign g[48256] = a[14] & g[31872];
assign g[64639] = b[14] & g[31872];
assign g[48257] = a[14] & g[31873];
assign g[64640] = b[14] & g[31873];
assign g[48258] = a[14] & g[31874];
assign g[64641] = b[14] & g[31874];
assign g[48259] = a[14] & g[31875];
assign g[64642] = b[14] & g[31875];
assign g[48260] = a[14] & g[31876];
assign g[64643] = b[14] & g[31876];
assign g[48261] = a[14] & g[31877];
assign g[64644] = b[14] & g[31877];
assign g[48262] = a[14] & g[31878];
assign g[64645] = b[14] & g[31878];
assign g[48263] = a[14] & g[31879];
assign g[64646] = b[14] & g[31879];
assign g[48264] = a[14] & g[31880];
assign g[64647] = b[14] & g[31880];
assign g[48265] = a[14] & g[31881];
assign g[64648] = b[14] & g[31881];
assign g[48266] = a[14] & g[31882];
assign g[64649] = b[14] & g[31882];
assign g[48267] = a[14] & g[31883];
assign g[64650] = b[14] & g[31883];
assign g[48268] = a[14] & g[31884];
assign g[64651] = b[14] & g[31884];
assign g[48269] = a[14] & g[31885];
assign g[64652] = b[14] & g[31885];
assign g[48270] = a[14] & g[31886];
assign g[64653] = b[14] & g[31886];
assign g[48271] = a[14] & g[31887];
assign g[64654] = b[14] & g[31887];
assign g[48272] = a[14] & g[31888];
assign g[64655] = b[14] & g[31888];
assign g[48273] = a[14] & g[31889];
assign g[64656] = b[14] & g[31889];
assign g[48274] = a[14] & g[31890];
assign g[64657] = b[14] & g[31890];
assign g[48275] = a[14] & g[31891];
assign g[64658] = b[14] & g[31891];
assign g[48276] = a[14] & g[31892];
assign g[64659] = b[14] & g[31892];
assign g[48277] = a[14] & g[31893];
assign g[64660] = b[14] & g[31893];
assign g[48278] = a[14] & g[31894];
assign g[64661] = b[14] & g[31894];
assign g[48279] = a[14] & g[31895];
assign g[64662] = b[14] & g[31895];
assign g[48280] = a[14] & g[31896];
assign g[64663] = b[14] & g[31896];
assign g[48281] = a[14] & g[31897];
assign g[64664] = b[14] & g[31897];
assign g[48282] = a[14] & g[31898];
assign g[64665] = b[14] & g[31898];
assign g[48283] = a[14] & g[31899];
assign g[64666] = b[14] & g[31899];
assign g[48284] = a[14] & g[31900];
assign g[64667] = b[14] & g[31900];
assign g[48285] = a[14] & g[31901];
assign g[64668] = b[14] & g[31901];
assign g[48286] = a[14] & g[31902];
assign g[64669] = b[14] & g[31902];
assign g[48287] = a[14] & g[31903];
assign g[64670] = b[14] & g[31903];
assign g[48288] = a[14] & g[31904];
assign g[64671] = b[14] & g[31904];
assign g[48289] = a[14] & g[31905];
assign g[64672] = b[14] & g[31905];
assign g[48290] = a[14] & g[31906];
assign g[64673] = b[14] & g[31906];
assign g[48291] = a[14] & g[31907];
assign g[64674] = b[14] & g[31907];
assign g[48292] = a[14] & g[31908];
assign g[64675] = b[14] & g[31908];
assign g[48293] = a[14] & g[31909];
assign g[64676] = b[14] & g[31909];
assign g[48294] = a[14] & g[31910];
assign g[64677] = b[14] & g[31910];
assign g[48295] = a[14] & g[31911];
assign g[64678] = b[14] & g[31911];
assign g[48296] = a[14] & g[31912];
assign g[64679] = b[14] & g[31912];
assign g[48297] = a[14] & g[31913];
assign g[64680] = b[14] & g[31913];
assign g[48298] = a[14] & g[31914];
assign g[64681] = b[14] & g[31914];
assign g[48299] = a[14] & g[31915];
assign g[64682] = b[14] & g[31915];
assign g[48300] = a[14] & g[31916];
assign g[64683] = b[14] & g[31916];
assign g[48301] = a[14] & g[31917];
assign g[64684] = b[14] & g[31917];
assign g[48302] = a[14] & g[31918];
assign g[64685] = b[14] & g[31918];
assign g[48303] = a[14] & g[31919];
assign g[64686] = b[14] & g[31919];
assign g[48304] = a[14] & g[31920];
assign g[64687] = b[14] & g[31920];
assign g[48305] = a[14] & g[31921];
assign g[64688] = b[14] & g[31921];
assign g[48306] = a[14] & g[31922];
assign g[64689] = b[14] & g[31922];
assign g[48307] = a[14] & g[31923];
assign g[64690] = b[14] & g[31923];
assign g[48308] = a[14] & g[31924];
assign g[64691] = b[14] & g[31924];
assign g[48309] = a[14] & g[31925];
assign g[64692] = b[14] & g[31925];
assign g[48310] = a[14] & g[31926];
assign g[64693] = b[14] & g[31926];
assign g[48311] = a[14] & g[31927];
assign g[64694] = b[14] & g[31927];
assign g[48312] = a[14] & g[31928];
assign g[64695] = b[14] & g[31928];
assign g[48313] = a[14] & g[31929];
assign g[64696] = b[14] & g[31929];
assign g[48314] = a[14] & g[31930];
assign g[64697] = b[14] & g[31930];
assign g[48315] = a[14] & g[31931];
assign g[64698] = b[14] & g[31931];
assign g[48316] = a[14] & g[31932];
assign g[64699] = b[14] & g[31932];
assign g[48317] = a[14] & g[31933];
assign g[64700] = b[14] & g[31933];
assign g[48318] = a[14] & g[31934];
assign g[64701] = b[14] & g[31934];
assign g[48319] = a[14] & g[31935];
assign g[64702] = b[14] & g[31935];
assign g[48320] = a[14] & g[31936];
assign g[64703] = b[14] & g[31936];
assign g[48321] = a[14] & g[31937];
assign g[64704] = b[14] & g[31937];
assign g[48322] = a[14] & g[31938];
assign g[64705] = b[14] & g[31938];
assign g[48323] = a[14] & g[31939];
assign g[64706] = b[14] & g[31939];
assign g[48324] = a[14] & g[31940];
assign g[64707] = b[14] & g[31940];
assign g[48325] = a[14] & g[31941];
assign g[64708] = b[14] & g[31941];
assign g[48326] = a[14] & g[31942];
assign g[64709] = b[14] & g[31942];
assign g[48327] = a[14] & g[31943];
assign g[64710] = b[14] & g[31943];
assign g[48328] = a[14] & g[31944];
assign g[64711] = b[14] & g[31944];
assign g[48329] = a[14] & g[31945];
assign g[64712] = b[14] & g[31945];
assign g[48330] = a[14] & g[31946];
assign g[64713] = b[14] & g[31946];
assign g[48331] = a[14] & g[31947];
assign g[64714] = b[14] & g[31947];
assign g[48332] = a[14] & g[31948];
assign g[64715] = b[14] & g[31948];
assign g[48333] = a[14] & g[31949];
assign g[64716] = b[14] & g[31949];
assign g[48334] = a[14] & g[31950];
assign g[64717] = b[14] & g[31950];
assign g[48335] = a[14] & g[31951];
assign g[64718] = b[14] & g[31951];
assign g[48336] = a[14] & g[31952];
assign g[64719] = b[14] & g[31952];
assign g[48337] = a[14] & g[31953];
assign g[64720] = b[14] & g[31953];
assign g[48338] = a[14] & g[31954];
assign g[64721] = b[14] & g[31954];
assign g[48339] = a[14] & g[31955];
assign g[64722] = b[14] & g[31955];
assign g[48340] = a[14] & g[31956];
assign g[64723] = b[14] & g[31956];
assign g[48341] = a[14] & g[31957];
assign g[64724] = b[14] & g[31957];
assign g[48342] = a[14] & g[31958];
assign g[64725] = b[14] & g[31958];
assign g[48343] = a[14] & g[31959];
assign g[64726] = b[14] & g[31959];
assign g[48344] = a[14] & g[31960];
assign g[64727] = b[14] & g[31960];
assign g[48345] = a[14] & g[31961];
assign g[64728] = b[14] & g[31961];
assign g[48346] = a[14] & g[31962];
assign g[64729] = b[14] & g[31962];
assign g[48347] = a[14] & g[31963];
assign g[64730] = b[14] & g[31963];
assign g[48348] = a[14] & g[31964];
assign g[64731] = b[14] & g[31964];
assign g[48349] = a[14] & g[31965];
assign g[64732] = b[14] & g[31965];
assign g[48350] = a[14] & g[31966];
assign g[64733] = b[14] & g[31966];
assign g[48351] = a[14] & g[31967];
assign g[64734] = b[14] & g[31967];
assign g[48352] = a[14] & g[31968];
assign g[64735] = b[14] & g[31968];
assign g[48353] = a[14] & g[31969];
assign g[64736] = b[14] & g[31969];
assign g[48354] = a[14] & g[31970];
assign g[64737] = b[14] & g[31970];
assign g[48355] = a[14] & g[31971];
assign g[64738] = b[14] & g[31971];
assign g[48356] = a[14] & g[31972];
assign g[64739] = b[14] & g[31972];
assign g[48357] = a[14] & g[31973];
assign g[64740] = b[14] & g[31973];
assign g[48358] = a[14] & g[31974];
assign g[64741] = b[14] & g[31974];
assign g[48359] = a[14] & g[31975];
assign g[64742] = b[14] & g[31975];
assign g[48360] = a[14] & g[31976];
assign g[64743] = b[14] & g[31976];
assign g[48361] = a[14] & g[31977];
assign g[64744] = b[14] & g[31977];
assign g[48362] = a[14] & g[31978];
assign g[64745] = b[14] & g[31978];
assign g[48363] = a[14] & g[31979];
assign g[64746] = b[14] & g[31979];
assign g[48364] = a[14] & g[31980];
assign g[64747] = b[14] & g[31980];
assign g[48365] = a[14] & g[31981];
assign g[64748] = b[14] & g[31981];
assign g[48366] = a[14] & g[31982];
assign g[64749] = b[14] & g[31982];
assign g[48367] = a[14] & g[31983];
assign g[64750] = b[14] & g[31983];
assign g[48368] = a[14] & g[31984];
assign g[64751] = b[14] & g[31984];
assign g[48369] = a[14] & g[31985];
assign g[64752] = b[14] & g[31985];
assign g[48370] = a[14] & g[31986];
assign g[64753] = b[14] & g[31986];
assign g[48371] = a[14] & g[31987];
assign g[64754] = b[14] & g[31987];
assign g[48372] = a[14] & g[31988];
assign g[64755] = b[14] & g[31988];
assign g[48373] = a[14] & g[31989];
assign g[64756] = b[14] & g[31989];
assign g[48374] = a[14] & g[31990];
assign g[64757] = b[14] & g[31990];
assign g[48375] = a[14] & g[31991];
assign g[64758] = b[14] & g[31991];
assign g[48376] = a[14] & g[31992];
assign g[64759] = b[14] & g[31992];
assign g[48377] = a[14] & g[31993];
assign g[64760] = b[14] & g[31993];
assign g[48378] = a[14] & g[31994];
assign g[64761] = b[14] & g[31994];
assign g[48379] = a[14] & g[31995];
assign g[64762] = b[14] & g[31995];
assign g[48380] = a[14] & g[31996];
assign g[64763] = b[14] & g[31996];
assign g[48381] = a[14] & g[31997];
assign g[64764] = b[14] & g[31997];
assign g[48382] = a[14] & g[31998];
assign g[64765] = b[14] & g[31998];
assign g[48383] = a[14] & g[31999];
assign g[64766] = b[14] & g[31999];
assign g[48384] = a[14] & g[32000];
assign g[64767] = b[14] & g[32000];
assign g[48385] = a[14] & g[32001];
assign g[64768] = b[14] & g[32001];
assign g[48386] = a[14] & g[32002];
assign g[64769] = b[14] & g[32002];
assign g[48387] = a[14] & g[32003];
assign g[64770] = b[14] & g[32003];
assign g[48388] = a[14] & g[32004];
assign g[64771] = b[14] & g[32004];
assign g[48389] = a[14] & g[32005];
assign g[64772] = b[14] & g[32005];
assign g[48390] = a[14] & g[32006];
assign g[64773] = b[14] & g[32006];
assign g[48391] = a[14] & g[32007];
assign g[64774] = b[14] & g[32007];
assign g[48392] = a[14] & g[32008];
assign g[64775] = b[14] & g[32008];
assign g[48393] = a[14] & g[32009];
assign g[64776] = b[14] & g[32009];
assign g[48394] = a[14] & g[32010];
assign g[64777] = b[14] & g[32010];
assign g[48395] = a[14] & g[32011];
assign g[64778] = b[14] & g[32011];
assign g[48396] = a[14] & g[32012];
assign g[64779] = b[14] & g[32012];
assign g[48397] = a[14] & g[32013];
assign g[64780] = b[14] & g[32013];
assign g[48398] = a[14] & g[32014];
assign g[64781] = b[14] & g[32014];
assign g[48399] = a[14] & g[32015];
assign g[64782] = b[14] & g[32015];
assign g[48400] = a[14] & g[32016];
assign g[64783] = b[14] & g[32016];
assign g[48401] = a[14] & g[32017];
assign g[64784] = b[14] & g[32017];
assign g[48402] = a[14] & g[32018];
assign g[64785] = b[14] & g[32018];
assign g[48403] = a[14] & g[32019];
assign g[64786] = b[14] & g[32019];
assign g[48404] = a[14] & g[32020];
assign g[64787] = b[14] & g[32020];
assign g[48405] = a[14] & g[32021];
assign g[64788] = b[14] & g[32021];
assign g[48406] = a[14] & g[32022];
assign g[64789] = b[14] & g[32022];
assign g[48407] = a[14] & g[32023];
assign g[64790] = b[14] & g[32023];
assign g[48408] = a[14] & g[32024];
assign g[64791] = b[14] & g[32024];
assign g[48409] = a[14] & g[32025];
assign g[64792] = b[14] & g[32025];
assign g[48410] = a[14] & g[32026];
assign g[64793] = b[14] & g[32026];
assign g[48411] = a[14] & g[32027];
assign g[64794] = b[14] & g[32027];
assign g[48412] = a[14] & g[32028];
assign g[64795] = b[14] & g[32028];
assign g[48413] = a[14] & g[32029];
assign g[64796] = b[14] & g[32029];
assign g[48414] = a[14] & g[32030];
assign g[64797] = b[14] & g[32030];
assign g[48415] = a[14] & g[32031];
assign g[64798] = b[14] & g[32031];
assign g[48416] = a[14] & g[32032];
assign g[64799] = b[14] & g[32032];
assign g[48417] = a[14] & g[32033];
assign g[64800] = b[14] & g[32033];
assign g[48418] = a[14] & g[32034];
assign g[64801] = b[14] & g[32034];
assign g[48419] = a[14] & g[32035];
assign g[64802] = b[14] & g[32035];
assign g[48420] = a[14] & g[32036];
assign g[64803] = b[14] & g[32036];
assign g[48421] = a[14] & g[32037];
assign g[64804] = b[14] & g[32037];
assign g[48422] = a[14] & g[32038];
assign g[64805] = b[14] & g[32038];
assign g[48423] = a[14] & g[32039];
assign g[64806] = b[14] & g[32039];
assign g[48424] = a[14] & g[32040];
assign g[64807] = b[14] & g[32040];
assign g[48425] = a[14] & g[32041];
assign g[64808] = b[14] & g[32041];
assign g[48426] = a[14] & g[32042];
assign g[64809] = b[14] & g[32042];
assign g[48427] = a[14] & g[32043];
assign g[64810] = b[14] & g[32043];
assign g[48428] = a[14] & g[32044];
assign g[64811] = b[14] & g[32044];
assign g[48429] = a[14] & g[32045];
assign g[64812] = b[14] & g[32045];
assign g[48430] = a[14] & g[32046];
assign g[64813] = b[14] & g[32046];
assign g[48431] = a[14] & g[32047];
assign g[64814] = b[14] & g[32047];
assign g[48432] = a[14] & g[32048];
assign g[64815] = b[14] & g[32048];
assign g[48433] = a[14] & g[32049];
assign g[64816] = b[14] & g[32049];
assign g[48434] = a[14] & g[32050];
assign g[64817] = b[14] & g[32050];
assign g[48435] = a[14] & g[32051];
assign g[64818] = b[14] & g[32051];
assign g[48436] = a[14] & g[32052];
assign g[64819] = b[14] & g[32052];
assign g[48437] = a[14] & g[32053];
assign g[64820] = b[14] & g[32053];
assign g[48438] = a[14] & g[32054];
assign g[64821] = b[14] & g[32054];
assign g[48439] = a[14] & g[32055];
assign g[64822] = b[14] & g[32055];
assign g[48440] = a[14] & g[32056];
assign g[64823] = b[14] & g[32056];
assign g[48441] = a[14] & g[32057];
assign g[64824] = b[14] & g[32057];
assign g[48442] = a[14] & g[32058];
assign g[64825] = b[14] & g[32058];
assign g[48443] = a[14] & g[32059];
assign g[64826] = b[14] & g[32059];
assign g[48444] = a[14] & g[32060];
assign g[64827] = b[14] & g[32060];
assign g[48445] = a[14] & g[32061];
assign g[64828] = b[14] & g[32061];
assign g[48446] = a[14] & g[32062];
assign g[64829] = b[14] & g[32062];
assign g[48447] = a[14] & g[32063];
assign g[64830] = b[14] & g[32063];
assign g[48448] = a[14] & g[32064];
assign g[64831] = b[14] & g[32064];
assign g[48449] = a[14] & g[32065];
assign g[64832] = b[14] & g[32065];
assign g[48450] = a[14] & g[32066];
assign g[64833] = b[14] & g[32066];
assign g[48451] = a[14] & g[32067];
assign g[64834] = b[14] & g[32067];
assign g[48452] = a[14] & g[32068];
assign g[64835] = b[14] & g[32068];
assign g[48453] = a[14] & g[32069];
assign g[64836] = b[14] & g[32069];
assign g[48454] = a[14] & g[32070];
assign g[64837] = b[14] & g[32070];
assign g[48455] = a[14] & g[32071];
assign g[64838] = b[14] & g[32071];
assign g[48456] = a[14] & g[32072];
assign g[64839] = b[14] & g[32072];
assign g[48457] = a[14] & g[32073];
assign g[64840] = b[14] & g[32073];
assign g[48458] = a[14] & g[32074];
assign g[64841] = b[14] & g[32074];
assign g[48459] = a[14] & g[32075];
assign g[64842] = b[14] & g[32075];
assign g[48460] = a[14] & g[32076];
assign g[64843] = b[14] & g[32076];
assign g[48461] = a[14] & g[32077];
assign g[64844] = b[14] & g[32077];
assign g[48462] = a[14] & g[32078];
assign g[64845] = b[14] & g[32078];
assign g[48463] = a[14] & g[32079];
assign g[64846] = b[14] & g[32079];
assign g[48464] = a[14] & g[32080];
assign g[64847] = b[14] & g[32080];
assign g[48465] = a[14] & g[32081];
assign g[64848] = b[14] & g[32081];
assign g[48466] = a[14] & g[32082];
assign g[64849] = b[14] & g[32082];
assign g[48467] = a[14] & g[32083];
assign g[64850] = b[14] & g[32083];
assign g[48468] = a[14] & g[32084];
assign g[64851] = b[14] & g[32084];
assign g[48469] = a[14] & g[32085];
assign g[64852] = b[14] & g[32085];
assign g[48470] = a[14] & g[32086];
assign g[64853] = b[14] & g[32086];
assign g[48471] = a[14] & g[32087];
assign g[64854] = b[14] & g[32087];
assign g[48472] = a[14] & g[32088];
assign g[64855] = b[14] & g[32088];
assign g[48473] = a[14] & g[32089];
assign g[64856] = b[14] & g[32089];
assign g[48474] = a[14] & g[32090];
assign g[64857] = b[14] & g[32090];
assign g[48475] = a[14] & g[32091];
assign g[64858] = b[14] & g[32091];
assign g[48476] = a[14] & g[32092];
assign g[64859] = b[14] & g[32092];
assign g[48477] = a[14] & g[32093];
assign g[64860] = b[14] & g[32093];
assign g[48478] = a[14] & g[32094];
assign g[64861] = b[14] & g[32094];
assign g[48479] = a[14] & g[32095];
assign g[64862] = b[14] & g[32095];
assign g[48480] = a[14] & g[32096];
assign g[64863] = b[14] & g[32096];
assign g[48481] = a[14] & g[32097];
assign g[64864] = b[14] & g[32097];
assign g[48482] = a[14] & g[32098];
assign g[64865] = b[14] & g[32098];
assign g[48483] = a[14] & g[32099];
assign g[64866] = b[14] & g[32099];
assign g[48484] = a[14] & g[32100];
assign g[64867] = b[14] & g[32100];
assign g[48485] = a[14] & g[32101];
assign g[64868] = b[14] & g[32101];
assign g[48486] = a[14] & g[32102];
assign g[64869] = b[14] & g[32102];
assign g[48487] = a[14] & g[32103];
assign g[64870] = b[14] & g[32103];
assign g[48488] = a[14] & g[32104];
assign g[64871] = b[14] & g[32104];
assign g[48489] = a[14] & g[32105];
assign g[64872] = b[14] & g[32105];
assign g[48490] = a[14] & g[32106];
assign g[64873] = b[14] & g[32106];
assign g[48491] = a[14] & g[32107];
assign g[64874] = b[14] & g[32107];
assign g[48492] = a[14] & g[32108];
assign g[64875] = b[14] & g[32108];
assign g[48493] = a[14] & g[32109];
assign g[64876] = b[14] & g[32109];
assign g[48494] = a[14] & g[32110];
assign g[64877] = b[14] & g[32110];
assign g[48495] = a[14] & g[32111];
assign g[64878] = b[14] & g[32111];
assign g[48496] = a[14] & g[32112];
assign g[64879] = b[14] & g[32112];
assign g[48497] = a[14] & g[32113];
assign g[64880] = b[14] & g[32113];
assign g[48498] = a[14] & g[32114];
assign g[64881] = b[14] & g[32114];
assign g[48499] = a[14] & g[32115];
assign g[64882] = b[14] & g[32115];
assign g[48500] = a[14] & g[32116];
assign g[64883] = b[14] & g[32116];
assign g[48501] = a[14] & g[32117];
assign g[64884] = b[14] & g[32117];
assign g[48502] = a[14] & g[32118];
assign g[64885] = b[14] & g[32118];
assign g[48503] = a[14] & g[32119];
assign g[64886] = b[14] & g[32119];
assign g[48504] = a[14] & g[32120];
assign g[64887] = b[14] & g[32120];
assign g[48505] = a[14] & g[32121];
assign g[64888] = b[14] & g[32121];
assign g[48506] = a[14] & g[32122];
assign g[64889] = b[14] & g[32122];
assign g[48507] = a[14] & g[32123];
assign g[64890] = b[14] & g[32123];
assign g[48508] = a[14] & g[32124];
assign g[64891] = b[14] & g[32124];
assign g[48509] = a[14] & g[32125];
assign g[64892] = b[14] & g[32125];
assign g[48510] = a[14] & g[32126];
assign g[64893] = b[14] & g[32126];
assign g[48511] = a[14] & g[32127];
assign g[64894] = b[14] & g[32127];
assign g[48512] = a[14] & g[32128];
assign g[64895] = b[14] & g[32128];
assign g[48513] = a[14] & g[32129];
assign g[64896] = b[14] & g[32129];
assign g[48514] = a[14] & g[32130];
assign g[64897] = b[14] & g[32130];
assign g[48515] = a[14] & g[32131];
assign g[64898] = b[14] & g[32131];
assign g[48516] = a[14] & g[32132];
assign g[64899] = b[14] & g[32132];
assign g[48517] = a[14] & g[32133];
assign g[64900] = b[14] & g[32133];
assign g[48518] = a[14] & g[32134];
assign g[64901] = b[14] & g[32134];
assign g[48519] = a[14] & g[32135];
assign g[64902] = b[14] & g[32135];
assign g[48520] = a[14] & g[32136];
assign g[64903] = b[14] & g[32136];
assign g[48521] = a[14] & g[32137];
assign g[64904] = b[14] & g[32137];
assign g[48522] = a[14] & g[32138];
assign g[64905] = b[14] & g[32138];
assign g[48523] = a[14] & g[32139];
assign g[64906] = b[14] & g[32139];
assign g[48524] = a[14] & g[32140];
assign g[64907] = b[14] & g[32140];
assign g[48525] = a[14] & g[32141];
assign g[64908] = b[14] & g[32141];
assign g[48526] = a[14] & g[32142];
assign g[64909] = b[14] & g[32142];
assign g[48527] = a[14] & g[32143];
assign g[64910] = b[14] & g[32143];
assign g[48528] = a[14] & g[32144];
assign g[64911] = b[14] & g[32144];
assign g[48529] = a[14] & g[32145];
assign g[64912] = b[14] & g[32145];
assign g[48530] = a[14] & g[32146];
assign g[64913] = b[14] & g[32146];
assign g[48531] = a[14] & g[32147];
assign g[64914] = b[14] & g[32147];
assign g[48532] = a[14] & g[32148];
assign g[64915] = b[14] & g[32148];
assign g[48533] = a[14] & g[32149];
assign g[64916] = b[14] & g[32149];
assign g[48534] = a[14] & g[32150];
assign g[64917] = b[14] & g[32150];
assign g[48535] = a[14] & g[32151];
assign g[64918] = b[14] & g[32151];
assign g[48536] = a[14] & g[32152];
assign g[64919] = b[14] & g[32152];
assign g[48537] = a[14] & g[32153];
assign g[64920] = b[14] & g[32153];
assign g[48538] = a[14] & g[32154];
assign g[64921] = b[14] & g[32154];
assign g[48539] = a[14] & g[32155];
assign g[64922] = b[14] & g[32155];
assign g[48540] = a[14] & g[32156];
assign g[64923] = b[14] & g[32156];
assign g[48541] = a[14] & g[32157];
assign g[64924] = b[14] & g[32157];
assign g[48542] = a[14] & g[32158];
assign g[64925] = b[14] & g[32158];
assign g[48543] = a[14] & g[32159];
assign g[64926] = b[14] & g[32159];
assign g[48544] = a[14] & g[32160];
assign g[64927] = b[14] & g[32160];
assign g[48545] = a[14] & g[32161];
assign g[64928] = b[14] & g[32161];
assign g[48546] = a[14] & g[32162];
assign g[64929] = b[14] & g[32162];
assign g[48547] = a[14] & g[32163];
assign g[64930] = b[14] & g[32163];
assign g[48548] = a[14] & g[32164];
assign g[64931] = b[14] & g[32164];
assign g[48549] = a[14] & g[32165];
assign g[64932] = b[14] & g[32165];
assign g[48550] = a[14] & g[32166];
assign g[64933] = b[14] & g[32166];
assign g[48551] = a[14] & g[32167];
assign g[64934] = b[14] & g[32167];
assign g[48552] = a[14] & g[32168];
assign g[64935] = b[14] & g[32168];
assign g[48553] = a[14] & g[32169];
assign g[64936] = b[14] & g[32169];
assign g[48554] = a[14] & g[32170];
assign g[64937] = b[14] & g[32170];
assign g[48555] = a[14] & g[32171];
assign g[64938] = b[14] & g[32171];
assign g[48556] = a[14] & g[32172];
assign g[64939] = b[14] & g[32172];
assign g[48557] = a[14] & g[32173];
assign g[64940] = b[14] & g[32173];
assign g[48558] = a[14] & g[32174];
assign g[64941] = b[14] & g[32174];
assign g[48559] = a[14] & g[32175];
assign g[64942] = b[14] & g[32175];
assign g[48560] = a[14] & g[32176];
assign g[64943] = b[14] & g[32176];
assign g[48561] = a[14] & g[32177];
assign g[64944] = b[14] & g[32177];
assign g[48562] = a[14] & g[32178];
assign g[64945] = b[14] & g[32178];
assign g[48563] = a[14] & g[32179];
assign g[64946] = b[14] & g[32179];
assign g[48564] = a[14] & g[32180];
assign g[64947] = b[14] & g[32180];
assign g[48565] = a[14] & g[32181];
assign g[64948] = b[14] & g[32181];
assign g[48566] = a[14] & g[32182];
assign g[64949] = b[14] & g[32182];
assign g[48567] = a[14] & g[32183];
assign g[64950] = b[14] & g[32183];
assign g[48568] = a[14] & g[32184];
assign g[64951] = b[14] & g[32184];
assign g[48569] = a[14] & g[32185];
assign g[64952] = b[14] & g[32185];
assign g[48570] = a[14] & g[32186];
assign g[64953] = b[14] & g[32186];
assign g[48571] = a[14] & g[32187];
assign g[64954] = b[14] & g[32187];
assign g[48572] = a[14] & g[32188];
assign g[64955] = b[14] & g[32188];
assign g[48573] = a[14] & g[32189];
assign g[64956] = b[14] & g[32189];
assign g[48574] = a[14] & g[32190];
assign g[64957] = b[14] & g[32190];
assign g[48575] = a[14] & g[32191];
assign g[64958] = b[14] & g[32191];
assign g[48576] = a[14] & g[32192];
assign g[64959] = b[14] & g[32192];
assign g[48577] = a[14] & g[32193];
assign g[64960] = b[14] & g[32193];
assign g[48578] = a[14] & g[32194];
assign g[64961] = b[14] & g[32194];
assign g[48579] = a[14] & g[32195];
assign g[64962] = b[14] & g[32195];
assign g[48580] = a[14] & g[32196];
assign g[64963] = b[14] & g[32196];
assign g[48581] = a[14] & g[32197];
assign g[64964] = b[14] & g[32197];
assign g[48582] = a[14] & g[32198];
assign g[64965] = b[14] & g[32198];
assign g[48583] = a[14] & g[32199];
assign g[64966] = b[14] & g[32199];
assign g[48584] = a[14] & g[32200];
assign g[64967] = b[14] & g[32200];
assign g[48585] = a[14] & g[32201];
assign g[64968] = b[14] & g[32201];
assign g[48586] = a[14] & g[32202];
assign g[64969] = b[14] & g[32202];
assign g[48587] = a[14] & g[32203];
assign g[64970] = b[14] & g[32203];
assign g[48588] = a[14] & g[32204];
assign g[64971] = b[14] & g[32204];
assign g[48589] = a[14] & g[32205];
assign g[64972] = b[14] & g[32205];
assign g[48590] = a[14] & g[32206];
assign g[64973] = b[14] & g[32206];
assign g[48591] = a[14] & g[32207];
assign g[64974] = b[14] & g[32207];
assign g[48592] = a[14] & g[32208];
assign g[64975] = b[14] & g[32208];
assign g[48593] = a[14] & g[32209];
assign g[64976] = b[14] & g[32209];
assign g[48594] = a[14] & g[32210];
assign g[64977] = b[14] & g[32210];
assign g[48595] = a[14] & g[32211];
assign g[64978] = b[14] & g[32211];
assign g[48596] = a[14] & g[32212];
assign g[64979] = b[14] & g[32212];
assign g[48597] = a[14] & g[32213];
assign g[64980] = b[14] & g[32213];
assign g[48598] = a[14] & g[32214];
assign g[64981] = b[14] & g[32214];
assign g[48599] = a[14] & g[32215];
assign g[64982] = b[14] & g[32215];
assign g[48600] = a[14] & g[32216];
assign g[64983] = b[14] & g[32216];
assign g[48601] = a[14] & g[32217];
assign g[64984] = b[14] & g[32217];
assign g[48602] = a[14] & g[32218];
assign g[64985] = b[14] & g[32218];
assign g[48603] = a[14] & g[32219];
assign g[64986] = b[14] & g[32219];
assign g[48604] = a[14] & g[32220];
assign g[64987] = b[14] & g[32220];
assign g[48605] = a[14] & g[32221];
assign g[64988] = b[14] & g[32221];
assign g[48606] = a[14] & g[32222];
assign g[64989] = b[14] & g[32222];
assign g[48607] = a[14] & g[32223];
assign g[64990] = b[14] & g[32223];
assign g[48608] = a[14] & g[32224];
assign g[64991] = b[14] & g[32224];
assign g[48609] = a[14] & g[32225];
assign g[64992] = b[14] & g[32225];
assign g[48610] = a[14] & g[32226];
assign g[64993] = b[14] & g[32226];
assign g[48611] = a[14] & g[32227];
assign g[64994] = b[14] & g[32227];
assign g[48612] = a[14] & g[32228];
assign g[64995] = b[14] & g[32228];
assign g[48613] = a[14] & g[32229];
assign g[64996] = b[14] & g[32229];
assign g[48614] = a[14] & g[32230];
assign g[64997] = b[14] & g[32230];
assign g[48615] = a[14] & g[32231];
assign g[64998] = b[14] & g[32231];
assign g[48616] = a[14] & g[32232];
assign g[64999] = b[14] & g[32232];
assign g[48617] = a[14] & g[32233];
assign g[65000] = b[14] & g[32233];
assign g[48618] = a[14] & g[32234];
assign g[65001] = b[14] & g[32234];
assign g[48619] = a[14] & g[32235];
assign g[65002] = b[14] & g[32235];
assign g[48620] = a[14] & g[32236];
assign g[65003] = b[14] & g[32236];
assign g[48621] = a[14] & g[32237];
assign g[65004] = b[14] & g[32237];
assign g[48622] = a[14] & g[32238];
assign g[65005] = b[14] & g[32238];
assign g[48623] = a[14] & g[32239];
assign g[65006] = b[14] & g[32239];
assign g[48624] = a[14] & g[32240];
assign g[65007] = b[14] & g[32240];
assign g[48625] = a[14] & g[32241];
assign g[65008] = b[14] & g[32241];
assign g[48626] = a[14] & g[32242];
assign g[65009] = b[14] & g[32242];
assign g[48627] = a[14] & g[32243];
assign g[65010] = b[14] & g[32243];
assign g[48628] = a[14] & g[32244];
assign g[65011] = b[14] & g[32244];
assign g[48629] = a[14] & g[32245];
assign g[65012] = b[14] & g[32245];
assign g[48630] = a[14] & g[32246];
assign g[65013] = b[14] & g[32246];
assign g[48631] = a[14] & g[32247];
assign g[65014] = b[14] & g[32247];
assign g[48632] = a[14] & g[32248];
assign g[65015] = b[14] & g[32248];
assign g[48633] = a[14] & g[32249];
assign g[65016] = b[14] & g[32249];
assign g[48634] = a[14] & g[32250];
assign g[65017] = b[14] & g[32250];
assign g[48635] = a[14] & g[32251];
assign g[65018] = b[14] & g[32251];
assign g[48636] = a[14] & g[32252];
assign g[65019] = b[14] & g[32252];
assign g[48637] = a[14] & g[32253];
assign g[65020] = b[14] & g[32253];
assign g[48638] = a[14] & g[32254];
assign g[65021] = b[14] & g[32254];
assign g[48639] = a[14] & g[32255];
assign g[65022] = b[14] & g[32255];
assign g[48640] = a[14] & g[32256];
assign g[65023] = b[14] & g[32256];
assign g[48641] = a[14] & g[32257];
assign g[65024] = b[14] & g[32257];
assign g[48642] = a[14] & g[32258];
assign g[65025] = b[14] & g[32258];
assign g[48643] = a[14] & g[32259];
assign g[65026] = b[14] & g[32259];
assign g[48644] = a[14] & g[32260];
assign g[65027] = b[14] & g[32260];
assign g[48645] = a[14] & g[32261];
assign g[65028] = b[14] & g[32261];
assign g[48646] = a[14] & g[32262];
assign g[65029] = b[14] & g[32262];
assign g[48647] = a[14] & g[32263];
assign g[65030] = b[14] & g[32263];
assign g[48648] = a[14] & g[32264];
assign g[65031] = b[14] & g[32264];
assign g[48649] = a[14] & g[32265];
assign g[65032] = b[14] & g[32265];
assign g[48650] = a[14] & g[32266];
assign g[65033] = b[14] & g[32266];
assign g[48651] = a[14] & g[32267];
assign g[65034] = b[14] & g[32267];
assign g[48652] = a[14] & g[32268];
assign g[65035] = b[14] & g[32268];
assign g[48653] = a[14] & g[32269];
assign g[65036] = b[14] & g[32269];
assign g[48654] = a[14] & g[32270];
assign g[65037] = b[14] & g[32270];
assign g[48655] = a[14] & g[32271];
assign g[65038] = b[14] & g[32271];
assign g[48656] = a[14] & g[32272];
assign g[65039] = b[14] & g[32272];
assign g[48657] = a[14] & g[32273];
assign g[65040] = b[14] & g[32273];
assign g[48658] = a[14] & g[32274];
assign g[65041] = b[14] & g[32274];
assign g[48659] = a[14] & g[32275];
assign g[65042] = b[14] & g[32275];
assign g[48660] = a[14] & g[32276];
assign g[65043] = b[14] & g[32276];
assign g[48661] = a[14] & g[32277];
assign g[65044] = b[14] & g[32277];
assign g[48662] = a[14] & g[32278];
assign g[65045] = b[14] & g[32278];
assign g[48663] = a[14] & g[32279];
assign g[65046] = b[14] & g[32279];
assign g[48664] = a[14] & g[32280];
assign g[65047] = b[14] & g[32280];
assign g[48665] = a[14] & g[32281];
assign g[65048] = b[14] & g[32281];
assign g[48666] = a[14] & g[32282];
assign g[65049] = b[14] & g[32282];
assign g[48667] = a[14] & g[32283];
assign g[65050] = b[14] & g[32283];
assign g[48668] = a[14] & g[32284];
assign g[65051] = b[14] & g[32284];
assign g[48669] = a[14] & g[32285];
assign g[65052] = b[14] & g[32285];
assign g[48670] = a[14] & g[32286];
assign g[65053] = b[14] & g[32286];
assign g[48671] = a[14] & g[32287];
assign g[65054] = b[14] & g[32287];
assign g[48672] = a[14] & g[32288];
assign g[65055] = b[14] & g[32288];
assign g[48673] = a[14] & g[32289];
assign g[65056] = b[14] & g[32289];
assign g[48674] = a[14] & g[32290];
assign g[65057] = b[14] & g[32290];
assign g[48675] = a[14] & g[32291];
assign g[65058] = b[14] & g[32291];
assign g[48676] = a[14] & g[32292];
assign g[65059] = b[14] & g[32292];
assign g[48677] = a[14] & g[32293];
assign g[65060] = b[14] & g[32293];
assign g[48678] = a[14] & g[32294];
assign g[65061] = b[14] & g[32294];
assign g[48679] = a[14] & g[32295];
assign g[65062] = b[14] & g[32295];
assign g[48680] = a[14] & g[32296];
assign g[65063] = b[14] & g[32296];
assign g[48681] = a[14] & g[32297];
assign g[65064] = b[14] & g[32297];
assign g[48682] = a[14] & g[32298];
assign g[65065] = b[14] & g[32298];
assign g[48683] = a[14] & g[32299];
assign g[65066] = b[14] & g[32299];
assign g[48684] = a[14] & g[32300];
assign g[65067] = b[14] & g[32300];
assign g[48685] = a[14] & g[32301];
assign g[65068] = b[14] & g[32301];
assign g[48686] = a[14] & g[32302];
assign g[65069] = b[14] & g[32302];
assign g[48687] = a[14] & g[32303];
assign g[65070] = b[14] & g[32303];
assign g[48688] = a[14] & g[32304];
assign g[65071] = b[14] & g[32304];
assign g[48689] = a[14] & g[32305];
assign g[65072] = b[14] & g[32305];
assign g[48690] = a[14] & g[32306];
assign g[65073] = b[14] & g[32306];
assign g[48691] = a[14] & g[32307];
assign g[65074] = b[14] & g[32307];
assign g[48692] = a[14] & g[32308];
assign g[65075] = b[14] & g[32308];
assign g[48693] = a[14] & g[32309];
assign g[65076] = b[14] & g[32309];
assign g[48694] = a[14] & g[32310];
assign g[65077] = b[14] & g[32310];
assign g[48695] = a[14] & g[32311];
assign g[65078] = b[14] & g[32311];
assign g[48696] = a[14] & g[32312];
assign g[65079] = b[14] & g[32312];
assign g[48697] = a[14] & g[32313];
assign g[65080] = b[14] & g[32313];
assign g[48698] = a[14] & g[32314];
assign g[65081] = b[14] & g[32314];
assign g[48699] = a[14] & g[32315];
assign g[65082] = b[14] & g[32315];
assign g[48700] = a[14] & g[32316];
assign g[65083] = b[14] & g[32316];
assign g[48701] = a[14] & g[32317];
assign g[65084] = b[14] & g[32317];
assign g[48702] = a[14] & g[32318];
assign g[65085] = b[14] & g[32318];
assign g[48703] = a[14] & g[32319];
assign g[65086] = b[14] & g[32319];
assign g[48704] = a[14] & g[32320];
assign g[65087] = b[14] & g[32320];
assign g[48705] = a[14] & g[32321];
assign g[65088] = b[14] & g[32321];
assign g[48706] = a[14] & g[32322];
assign g[65089] = b[14] & g[32322];
assign g[48707] = a[14] & g[32323];
assign g[65090] = b[14] & g[32323];
assign g[48708] = a[14] & g[32324];
assign g[65091] = b[14] & g[32324];
assign g[48709] = a[14] & g[32325];
assign g[65092] = b[14] & g[32325];
assign g[48710] = a[14] & g[32326];
assign g[65093] = b[14] & g[32326];
assign g[48711] = a[14] & g[32327];
assign g[65094] = b[14] & g[32327];
assign g[48712] = a[14] & g[32328];
assign g[65095] = b[14] & g[32328];
assign g[48713] = a[14] & g[32329];
assign g[65096] = b[14] & g[32329];
assign g[48714] = a[14] & g[32330];
assign g[65097] = b[14] & g[32330];
assign g[48715] = a[14] & g[32331];
assign g[65098] = b[14] & g[32331];
assign g[48716] = a[14] & g[32332];
assign g[65099] = b[14] & g[32332];
assign g[48717] = a[14] & g[32333];
assign g[65100] = b[14] & g[32333];
assign g[48718] = a[14] & g[32334];
assign g[65101] = b[14] & g[32334];
assign g[48719] = a[14] & g[32335];
assign g[65102] = b[14] & g[32335];
assign g[48720] = a[14] & g[32336];
assign g[65103] = b[14] & g[32336];
assign g[48721] = a[14] & g[32337];
assign g[65104] = b[14] & g[32337];
assign g[48722] = a[14] & g[32338];
assign g[65105] = b[14] & g[32338];
assign g[48723] = a[14] & g[32339];
assign g[65106] = b[14] & g[32339];
assign g[48724] = a[14] & g[32340];
assign g[65107] = b[14] & g[32340];
assign g[48725] = a[14] & g[32341];
assign g[65108] = b[14] & g[32341];
assign g[48726] = a[14] & g[32342];
assign g[65109] = b[14] & g[32342];
assign g[48727] = a[14] & g[32343];
assign g[65110] = b[14] & g[32343];
assign g[48728] = a[14] & g[32344];
assign g[65111] = b[14] & g[32344];
assign g[48729] = a[14] & g[32345];
assign g[65112] = b[14] & g[32345];
assign g[48730] = a[14] & g[32346];
assign g[65113] = b[14] & g[32346];
assign g[48731] = a[14] & g[32347];
assign g[65114] = b[14] & g[32347];
assign g[48732] = a[14] & g[32348];
assign g[65115] = b[14] & g[32348];
assign g[48733] = a[14] & g[32349];
assign g[65116] = b[14] & g[32349];
assign g[48734] = a[14] & g[32350];
assign g[65117] = b[14] & g[32350];
assign g[48735] = a[14] & g[32351];
assign g[65118] = b[14] & g[32351];
assign g[48736] = a[14] & g[32352];
assign g[65119] = b[14] & g[32352];
assign g[48737] = a[14] & g[32353];
assign g[65120] = b[14] & g[32353];
assign g[48738] = a[14] & g[32354];
assign g[65121] = b[14] & g[32354];
assign g[48739] = a[14] & g[32355];
assign g[65122] = b[14] & g[32355];
assign g[48740] = a[14] & g[32356];
assign g[65123] = b[14] & g[32356];
assign g[48741] = a[14] & g[32357];
assign g[65124] = b[14] & g[32357];
assign g[48742] = a[14] & g[32358];
assign g[65125] = b[14] & g[32358];
assign g[48743] = a[14] & g[32359];
assign g[65126] = b[14] & g[32359];
assign g[48744] = a[14] & g[32360];
assign g[65127] = b[14] & g[32360];
assign g[48745] = a[14] & g[32361];
assign g[65128] = b[14] & g[32361];
assign g[48746] = a[14] & g[32362];
assign g[65129] = b[14] & g[32362];
assign g[48747] = a[14] & g[32363];
assign g[65130] = b[14] & g[32363];
assign g[48748] = a[14] & g[32364];
assign g[65131] = b[14] & g[32364];
assign g[48749] = a[14] & g[32365];
assign g[65132] = b[14] & g[32365];
assign g[48750] = a[14] & g[32366];
assign g[65133] = b[14] & g[32366];
assign g[48751] = a[14] & g[32367];
assign g[65134] = b[14] & g[32367];
assign g[48752] = a[14] & g[32368];
assign g[65135] = b[14] & g[32368];
assign g[48753] = a[14] & g[32369];
assign g[65136] = b[14] & g[32369];
assign g[48754] = a[14] & g[32370];
assign g[65137] = b[14] & g[32370];
assign g[48755] = a[14] & g[32371];
assign g[65138] = b[14] & g[32371];
assign g[48756] = a[14] & g[32372];
assign g[65139] = b[14] & g[32372];
assign g[48757] = a[14] & g[32373];
assign g[65140] = b[14] & g[32373];
assign g[48758] = a[14] & g[32374];
assign g[65141] = b[14] & g[32374];
assign g[48759] = a[14] & g[32375];
assign g[65142] = b[14] & g[32375];
assign g[48760] = a[14] & g[32376];
assign g[65143] = b[14] & g[32376];
assign g[48761] = a[14] & g[32377];
assign g[65144] = b[14] & g[32377];
assign g[48762] = a[14] & g[32378];
assign g[65145] = b[14] & g[32378];
assign g[48763] = a[14] & g[32379];
assign g[65146] = b[14] & g[32379];
assign g[48764] = a[14] & g[32380];
assign g[65147] = b[14] & g[32380];
assign g[48765] = a[14] & g[32381];
assign g[65148] = b[14] & g[32381];
assign g[48766] = a[14] & g[32382];
assign g[65149] = b[14] & g[32382];
assign g[48767] = a[14] & g[32383];
assign g[65150] = b[14] & g[32383];
assign g[48768] = a[14] & g[32384];
assign g[65151] = b[14] & g[32384];
assign g[48769] = a[14] & g[32385];
assign g[65152] = b[14] & g[32385];
assign g[48770] = a[14] & g[32386];
assign g[65153] = b[14] & g[32386];
assign g[48771] = a[14] & g[32387];
assign g[65154] = b[14] & g[32387];
assign g[48772] = a[14] & g[32388];
assign g[65155] = b[14] & g[32388];
assign g[48773] = a[14] & g[32389];
assign g[65156] = b[14] & g[32389];
assign g[48774] = a[14] & g[32390];
assign g[65157] = b[14] & g[32390];
assign g[48775] = a[14] & g[32391];
assign g[65158] = b[14] & g[32391];
assign g[48776] = a[14] & g[32392];
assign g[65159] = b[14] & g[32392];
assign g[48777] = a[14] & g[32393];
assign g[65160] = b[14] & g[32393];
assign g[48778] = a[14] & g[32394];
assign g[65161] = b[14] & g[32394];
assign g[48779] = a[14] & g[32395];
assign g[65162] = b[14] & g[32395];
assign g[48780] = a[14] & g[32396];
assign g[65163] = b[14] & g[32396];
assign g[48781] = a[14] & g[32397];
assign g[65164] = b[14] & g[32397];
assign g[48782] = a[14] & g[32398];
assign g[65165] = b[14] & g[32398];
assign g[48783] = a[14] & g[32399];
assign g[65166] = b[14] & g[32399];
assign g[48784] = a[14] & g[32400];
assign g[65167] = b[14] & g[32400];
assign g[48785] = a[14] & g[32401];
assign g[65168] = b[14] & g[32401];
assign g[48786] = a[14] & g[32402];
assign g[65169] = b[14] & g[32402];
assign g[48787] = a[14] & g[32403];
assign g[65170] = b[14] & g[32403];
assign g[48788] = a[14] & g[32404];
assign g[65171] = b[14] & g[32404];
assign g[48789] = a[14] & g[32405];
assign g[65172] = b[14] & g[32405];
assign g[48790] = a[14] & g[32406];
assign g[65173] = b[14] & g[32406];
assign g[48791] = a[14] & g[32407];
assign g[65174] = b[14] & g[32407];
assign g[48792] = a[14] & g[32408];
assign g[65175] = b[14] & g[32408];
assign g[48793] = a[14] & g[32409];
assign g[65176] = b[14] & g[32409];
assign g[48794] = a[14] & g[32410];
assign g[65177] = b[14] & g[32410];
assign g[48795] = a[14] & g[32411];
assign g[65178] = b[14] & g[32411];
assign g[48796] = a[14] & g[32412];
assign g[65179] = b[14] & g[32412];
assign g[48797] = a[14] & g[32413];
assign g[65180] = b[14] & g[32413];
assign g[48798] = a[14] & g[32414];
assign g[65181] = b[14] & g[32414];
assign g[48799] = a[14] & g[32415];
assign g[65182] = b[14] & g[32415];
assign g[48800] = a[14] & g[32416];
assign g[65183] = b[14] & g[32416];
assign g[48801] = a[14] & g[32417];
assign g[65184] = b[14] & g[32417];
assign g[48802] = a[14] & g[32418];
assign g[65185] = b[14] & g[32418];
assign g[48803] = a[14] & g[32419];
assign g[65186] = b[14] & g[32419];
assign g[48804] = a[14] & g[32420];
assign g[65187] = b[14] & g[32420];
assign g[48805] = a[14] & g[32421];
assign g[65188] = b[14] & g[32421];
assign g[48806] = a[14] & g[32422];
assign g[65189] = b[14] & g[32422];
assign g[48807] = a[14] & g[32423];
assign g[65190] = b[14] & g[32423];
assign g[48808] = a[14] & g[32424];
assign g[65191] = b[14] & g[32424];
assign g[48809] = a[14] & g[32425];
assign g[65192] = b[14] & g[32425];
assign g[48810] = a[14] & g[32426];
assign g[65193] = b[14] & g[32426];
assign g[48811] = a[14] & g[32427];
assign g[65194] = b[14] & g[32427];
assign g[48812] = a[14] & g[32428];
assign g[65195] = b[14] & g[32428];
assign g[48813] = a[14] & g[32429];
assign g[65196] = b[14] & g[32429];
assign g[48814] = a[14] & g[32430];
assign g[65197] = b[14] & g[32430];
assign g[48815] = a[14] & g[32431];
assign g[65198] = b[14] & g[32431];
assign g[48816] = a[14] & g[32432];
assign g[65199] = b[14] & g[32432];
assign g[48817] = a[14] & g[32433];
assign g[65200] = b[14] & g[32433];
assign g[48818] = a[14] & g[32434];
assign g[65201] = b[14] & g[32434];
assign g[48819] = a[14] & g[32435];
assign g[65202] = b[14] & g[32435];
assign g[48820] = a[14] & g[32436];
assign g[65203] = b[14] & g[32436];
assign g[48821] = a[14] & g[32437];
assign g[65204] = b[14] & g[32437];
assign g[48822] = a[14] & g[32438];
assign g[65205] = b[14] & g[32438];
assign g[48823] = a[14] & g[32439];
assign g[65206] = b[14] & g[32439];
assign g[48824] = a[14] & g[32440];
assign g[65207] = b[14] & g[32440];
assign g[48825] = a[14] & g[32441];
assign g[65208] = b[14] & g[32441];
assign g[48826] = a[14] & g[32442];
assign g[65209] = b[14] & g[32442];
assign g[48827] = a[14] & g[32443];
assign g[65210] = b[14] & g[32443];
assign g[48828] = a[14] & g[32444];
assign g[65211] = b[14] & g[32444];
assign g[48829] = a[14] & g[32445];
assign g[65212] = b[14] & g[32445];
assign g[48830] = a[14] & g[32446];
assign g[65213] = b[14] & g[32446];
assign g[48831] = a[14] & g[32447];
assign g[65214] = b[14] & g[32447];
assign g[48832] = a[14] & g[32448];
assign g[65215] = b[14] & g[32448];
assign g[48833] = a[14] & g[32449];
assign g[65216] = b[14] & g[32449];
assign g[48834] = a[14] & g[32450];
assign g[65217] = b[14] & g[32450];
assign g[48835] = a[14] & g[32451];
assign g[65218] = b[14] & g[32451];
assign g[48836] = a[14] & g[32452];
assign g[65219] = b[14] & g[32452];
assign g[48837] = a[14] & g[32453];
assign g[65220] = b[14] & g[32453];
assign g[48838] = a[14] & g[32454];
assign g[65221] = b[14] & g[32454];
assign g[48839] = a[14] & g[32455];
assign g[65222] = b[14] & g[32455];
assign g[48840] = a[14] & g[32456];
assign g[65223] = b[14] & g[32456];
assign g[48841] = a[14] & g[32457];
assign g[65224] = b[14] & g[32457];
assign g[48842] = a[14] & g[32458];
assign g[65225] = b[14] & g[32458];
assign g[48843] = a[14] & g[32459];
assign g[65226] = b[14] & g[32459];
assign g[48844] = a[14] & g[32460];
assign g[65227] = b[14] & g[32460];
assign g[48845] = a[14] & g[32461];
assign g[65228] = b[14] & g[32461];
assign g[48846] = a[14] & g[32462];
assign g[65229] = b[14] & g[32462];
assign g[48847] = a[14] & g[32463];
assign g[65230] = b[14] & g[32463];
assign g[48848] = a[14] & g[32464];
assign g[65231] = b[14] & g[32464];
assign g[48849] = a[14] & g[32465];
assign g[65232] = b[14] & g[32465];
assign g[48850] = a[14] & g[32466];
assign g[65233] = b[14] & g[32466];
assign g[48851] = a[14] & g[32467];
assign g[65234] = b[14] & g[32467];
assign g[48852] = a[14] & g[32468];
assign g[65235] = b[14] & g[32468];
assign g[48853] = a[14] & g[32469];
assign g[65236] = b[14] & g[32469];
assign g[48854] = a[14] & g[32470];
assign g[65237] = b[14] & g[32470];
assign g[48855] = a[14] & g[32471];
assign g[65238] = b[14] & g[32471];
assign g[48856] = a[14] & g[32472];
assign g[65239] = b[14] & g[32472];
assign g[48857] = a[14] & g[32473];
assign g[65240] = b[14] & g[32473];
assign g[48858] = a[14] & g[32474];
assign g[65241] = b[14] & g[32474];
assign g[48859] = a[14] & g[32475];
assign g[65242] = b[14] & g[32475];
assign g[48860] = a[14] & g[32476];
assign g[65243] = b[14] & g[32476];
assign g[48861] = a[14] & g[32477];
assign g[65244] = b[14] & g[32477];
assign g[48862] = a[14] & g[32478];
assign g[65245] = b[14] & g[32478];
assign g[48863] = a[14] & g[32479];
assign g[65246] = b[14] & g[32479];
assign g[48864] = a[14] & g[32480];
assign g[65247] = b[14] & g[32480];
assign g[48865] = a[14] & g[32481];
assign g[65248] = b[14] & g[32481];
assign g[48866] = a[14] & g[32482];
assign g[65249] = b[14] & g[32482];
assign g[48867] = a[14] & g[32483];
assign g[65250] = b[14] & g[32483];
assign g[48868] = a[14] & g[32484];
assign g[65251] = b[14] & g[32484];
assign g[48869] = a[14] & g[32485];
assign g[65252] = b[14] & g[32485];
assign g[48870] = a[14] & g[32486];
assign g[65253] = b[14] & g[32486];
assign g[48871] = a[14] & g[32487];
assign g[65254] = b[14] & g[32487];
assign g[48872] = a[14] & g[32488];
assign g[65255] = b[14] & g[32488];
assign g[48873] = a[14] & g[32489];
assign g[65256] = b[14] & g[32489];
assign g[48874] = a[14] & g[32490];
assign g[65257] = b[14] & g[32490];
assign g[48875] = a[14] & g[32491];
assign g[65258] = b[14] & g[32491];
assign g[48876] = a[14] & g[32492];
assign g[65259] = b[14] & g[32492];
assign g[48877] = a[14] & g[32493];
assign g[65260] = b[14] & g[32493];
assign g[48878] = a[14] & g[32494];
assign g[65261] = b[14] & g[32494];
assign g[48879] = a[14] & g[32495];
assign g[65262] = b[14] & g[32495];
assign g[48880] = a[14] & g[32496];
assign g[65263] = b[14] & g[32496];
assign g[48881] = a[14] & g[32497];
assign g[65264] = b[14] & g[32497];
assign g[48882] = a[14] & g[32498];
assign g[65265] = b[14] & g[32498];
assign g[48883] = a[14] & g[32499];
assign g[65266] = b[14] & g[32499];
assign g[48884] = a[14] & g[32500];
assign g[65267] = b[14] & g[32500];
assign g[48885] = a[14] & g[32501];
assign g[65268] = b[14] & g[32501];
assign g[48886] = a[14] & g[32502];
assign g[65269] = b[14] & g[32502];
assign g[48887] = a[14] & g[32503];
assign g[65270] = b[14] & g[32503];
assign g[48888] = a[14] & g[32504];
assign g[65271] = b[14] & g[32504];
assign g[48889] = a[14] & g[32505];
assign g[65272] = b[14] & g[32505];
assign g[48890] = a[14] & g[32506];
assign g[65273] = b[14] & g[32506];
assign g[48891] = a[14] & g[32507];
assign g[65274] = b[14] & g[32507];
assign g[48892] = a[14] & g[32508];
assign g[65275] = b[14] & g[32508];
assign g[48893] = a[14] & g[32509];
assign g[65276] = b[14] & g[32509];
assign g[48894] = a[14] & g[32510];
assign g[65277] = b[14] & g[32510];
assign g[48895] = a[14] & g[32511];
assign g[65278] = b[14] & g[32511];
assign g[48896] = a[14] & g[32512];
assign g[65279] = b[14] & g[32512];
assign g[48897] = a[14] & g[32513];
assign g[65280] = b[14] & g[32513];
assign g[48898] = a[14] & g[32514];
assign g[65281] = b[14] & g[32514];
assign g[48899] = a[14] & g[32515];
assign g[65282] = b[14] & g[32515];
assign g[48900] = a[14] & g[32516];
assign g[65283] = b[14] & g[32516];
assign g[48901] = a[14] & g[32517];
assign g[65284] = b[14] & g[32517];
assign g[48902] = a[14] & g[32518];
assign g[65285] = b[14] & g[32518];
assign g[48903] = a[14] & g[32519];
assign g[65286] = b[14] & g[32519];
assign g[48904] = a[14] & g[32520];
assign g[65287] = b[14] & g[32520];
assign g[48905] = a[14] & g[32521];
assign g[65288] = b[14] & g[32521];
assign g[48906] = a[14] & g[32522];
assign g[65289] = b[14] & g[32522];
assign g[48907] = a[14] & g[32523];
assign g[65290] = b[14] & g[32523];
assign g[48908] = a[14] & g[32524];
assign g[65291] = b[14] & g[32524];
assign g[48909] = a[14] & g[32525];
assign g[65292] = b[14] & g[32525];
assign g[48910] = a[14] & g[32526];
assign g[65293] = b[14] & g[32526];
assign g[48911] = a[14] & g[32527];
assign g[65294] = b[14] & g[32527];
assign g[48912] = a[14] & g[32528];
assign g[65295] = b[14] & g[32528];
assign g[48913] = a[14] & g[32529];
assign g[65296] = b[14] & g[32529];
assign g[48914] = a[14] & g[32530];
assign g[65297] = b[14] & g[32530];
assign g[48915] = a[14] & g[32531];
assign g[65298] = b[14] & g[32531];
assign g[48916] = a[14] & g[32532];
assign g[65299] = b[14] & g[32532];
assign g[48917] = a[14] & g[32533];
assign g[65300] = b[14] & g[32533];
assign g[48918] = a[14] & g[32534];
assign g[65301] = b[14] & g[32534];
assign g[48919] = a[14] & g[32535];
assign g[65302] = b[14] & g[32535];
assign g[48920] = a[14] & g[32536];
assign g[65303] = b[14] & g[32536];
assign g[48921] = a[14] & g[32537];
assign g[65304] = b[14] & g[32537];
assign g[48922] = a[14] & g[32538];
assign g[65305] = b[14] & g[32538];
assign g[48923] = a[14] & g[32539];
assign g[65306] = b[14] & g[32539];
assign g[48924] = a[14] & g[32540];
assign g[65307] = b[14] & g[32540];
assign g[48925] = a[14] & g[32541];
assign g[65308] = b[14] & g[32541];
assign g[48926] = a[14] & g[32542];
assign g[65309] = b[14] & g[32542];
assign g[48927] = a[14] & g[32543];
assign g[65310] = b[14] & g[32543];
assign g[48928] = a[14] & g[32544];
assign g[65311] = b[14] & g[32544];
assign g[48929] = a[14] & g[32545];
assign g[65312] = b[14] & g[32545];
assign g[48930] = a[14] & g[32546];
assign g[65313] = b[14] & g[32546];
assign g[48931] = a[14] & g[32547];
assign g[65314] = b[14] & g[32547];
assign g[48932] = a[14] & g[32548];
assign g[65315] = b[14] & g[32548];
assign g[48933] = a[14] & g[32549];
assign g[65316] = b[14] & g[32549];
assign g[48934] = a[14] & g[32550];
assign g[65317] = b[14] & g[32550];
assign g[48935] = a[14] & g[32551];
assign g[65318] = b[14] & g[32551];
assign g[48936] = a[14] & g[32552];
assign g[65319] = b[14] & g[32552];
assign g[48937] = a[14] & g[32553];
assign g[65320] = b[14] & g[32553];
assign g[48938] = a[14] & g[32554];
assign g[65321] = b[14] & g[32554];
assign g[48939] = a[14] & g[32555];
assign g[65322] = b[14] & g[32555];
assign g[48940] = a[14] & g[32556];
assign g[65323] = b[14] & g[32556];
assign g[48941] = a[14] & g[32557];
assign g[65324] = b[14] & g[32557];
assign g[48942] = a[14] & g[32558];
assign g[65325] = b[14] & g[32558];
assign g[48943] = a[14] & g[32559];
assign g[65326] = b[14] & g[32559];
assign g[48944] = a[14] & g[32560];
assign g[65327] = b[14] & g[32560];
assign g[48945] = a[14] & g[32561];
assign g[65328] = b[14] & g[32561];
assign g[48946] = a[14] & g[32562];
assign g[65329] = b[14] & g[32562];
assign g[48947] = a[14] & g[32563];
assign g[65330] = b[14] & g[32563];
assign g[48948] = a[14] & g[32564];
assign g[65331] = b[14] & g[32564];
assign g[48949] = a[14] & g[32565];
assign g[65332] = b[14] & g[32565];
assign g[48950] = a[14] & g[32566];
assign g[65333] = b[14] & g[32566];
assign g[48951] = a[14] & g[32567];
assign g[65334] = b[14] & g[32567];
assign g[48952] = a[14] & g[32568];
assign g[65335] = b[14] & g[32568];
assign g[48953] = a[14] & g[32569];
assign g[65336] = b[14] & g[32569];
assign g[48954] = a[14] & g[32570];
assign g[65337] = b[14] & g[32570];
assign g[48955] = a[14] & g[32571];
assign g[65338] = b[14] & g[32571];
assign g[48956] = a[14] & g[32572];
assign g[65339] = b[14] & g[32572];
assign g[48957] = a[14] & g[32573];
assign g[65340] = b[14] & g[32573];
assign g[48958] = a[14] & g[32574];
assign g[65341] = b[14] & g[32574];
assign g[48959] = a[14] & g[32575];
assign g[65342] = b[14] & g[32575];
assign g[48960] = a[14] & g[32576];
assign g[65343] = b[14] & g[32576];
assign g[48961] = a[14] & g[32577];
assign g[65344] = b[14] & g[32577];
assign g[48962] = a[14] & g[32578];
assign g[65345] = b[14] & g[32578];
assign g[48963] = a[14] & g[32579];
assign g[65346] = b[14] & g[32579];
assign g[48964] = a[14] & g[32580];
assign g[65347] = b[14] & g[32580];
assign g[48965] = a[14] & g[32581];
assign g[65348] = b[14] & g[32581];
assign g[48966] = a[14] & g[32582];
assign g[65349] = b[14] & g[32582];
assign g[48967] = a[14] & g[32583];
assign g[65350] = b[14] & g[32583];
assign g[48968] = a[14] & g[32584];
assign g[65351] = b[14] & g[32584];
assign g[48969] = a[14] & g[32585];
assign g[65352] = b[14] & g[32585];
assign g[48970] = a[14] & g[32586];
assign g[65353] = b[14] & g[32586];
assign g[48971] = a[14] & g[32587];
assign g[65354] = b[14] & g[32587];
assign g[48972] = a[14] & g[32588];
assign g[65355] = b[14] & g[32588];
assign g[48973] = a[14] & g[32589];
assign g[65356] = b[14] & g[32589];
assign g[48974] = a[14] & g[32590];
assign g[65357] = b[14] & g[32590];
assign g[48975] = a[14] & g[32591];
assign g[65358] = b[14] & g[32591];
assign g[48976] = a[14] & g[32592];
assign g[65359] = b[14] & g[32592];
assign g[48977] = a[14] & g[32593];
assign g[65360] = b[14] & g[32593];
assign g[48978] = a[14] & g[32594];
assign g[65361] = b[14] & g[32594];
assign g[48979] = a[14] & g[32595];
assign g[65362] = b[14] & g[32595];
assign g[48980] = a[14] & g[32596];
assign g[65363] = b[14] & g[32596];
assign g[48981] = a[14] & g[32597];
assign g[65364] = b[14] & g[32597];
assign g[48982] = a[14] & g[32598];
assign g[65365] = b[14] & g[32598];
assign g[48983] = a[14] & g[32599];
assign g[65366] = b[14] & g[32599];
assign g[48984] = a[14] & g[32600];
assign g[65367] = b[14] & g[32600];
assign g[48985] = a[14] & g[32601];
assign g[65368] = b[14] & g[32601];
assign g[48986] = a[14] & g[32602];
assign g[65369] = b[14] & g[32602];
assign g[48987] = a[14] & g[32603];
assign g[65370] = b[14] & g[32603];
assign g[48988] = a[14] & g[32604];
assign g[65371] = b[14] & g[32604];
assign g[48989] = a[14] & g[32605];
assign g[65372] = b[14] & g[32605];
assign g[48990] = a[14] & g[32606];
assign g[65373] = b[14] & g[32606];
assign g[48991] = a[14] & g[32607];
assign g[65374] = b[14] & g[32607];
assign g[48992] = a[14] & g[32608];
assign g[65375] = b[14] & g[32608];
assign g[48993] = a[14] & g[32609];
assign g[65376] = b[14] & g[32609];
assign g[48994] = a[14] & g[32610];
assign g[65377] = b[14] & g[32610];
assign g[48995] = a[14] & g[32611];
assign g[65378] = b[14] & g[32611];
assign g[48996] = a[14] & g[32612];
assign g[65379] = b[14] & g[32612];
assign g[48997] = a[14] & g[32613];
assign g[65380] = b[14] & g[32613];
assign g[48998] = a[14] & g[32614];
assign g[65381] = b[14] & g[32614];
assign g[48999] = a[14] & g[32615];
assign g[65382] = b[14] & g[32615];
assign g[49000] = a[14] & g[32616];
assign g[65383] = b[14] & g[32616];
assign g[49001] = a[14] & g[32617];
assign g[65384] = b[14] & g[32617];
assign g[49002] = a[14] & g[32618];
assign g[65385] = b[14] & g[32618];
assign g[49003] = a[14] & g[32619];
assign g[65386] = b[14] & g[32619];
assign g[49004] = a[14] & g[32620];
assign g[65387] = b[14] & g[32620];
assign g[49005] = a[14] & g[32621];
assign g[65388] = b[14] & g[32621];
assign g[49006] = a[14] & g[32622];
assign g[65389] = b[14] & g[32622];
assign g[49007] = a[14] & g[32623];
assign g[65390] = b[14] & g[32623];
assign g[49008] = a[14] & g[32624];
assign g[65391] = b[14] & g[32624];
assign g[49009] = a[14] & g[32625];
assign g[65392] = b[14] & g[32625];
assign g[49010] = a[14] & g[32626];
assign g[65393] = b[14] & g[32626];
assign g[49011] = a[14] & g[32627];
assign g[65394] = b[14] & g[32627];
assign g[49012] = a[14] & g[32628];
assign g[65395] = b[14] & g[32628];
assign g[49013] = a[14] & g[32629];
assign g[65396] = b[14] & g[32629];
assign g[49014] = a[14] & g[32630];
assign g[65397] = b[14] & g[32630];
assign g[49015] = a[14] & g[32631];
assign g[65398] = b[14] & g[32631];
assign g[49016] = a[14] & g[32632];
assign g[65399] = b[14] & g[32632];
assign g[49017] = a[14] & g[32633];
assign g[65400] = b[14] & g[32633];
assign g[49018] = a[14] & g[32634];
assign g[65401] = b[14] & g[32634];
assign g[49019] = a[14] & g[32635];
assign g[65402] = b[14] & g[32635];
assign g[49020] = a[14] & g[32636];
assign g[65403] = b[14] & g[32636];
assign g[49021] = a[14] & g[32637];
assign g[65404] = b[14] & g[32637];
assign g[49022] = a[14] & g[32638];
assign g[65405] = b[14] & g[32638];
assign g[49023] = a[14] & g[32639];
assign g[65406] = b[14] & g[32639];
assign g[49024] = a[14] & g[32640];
assign g[65407] = b[14] & g[32640];
assign g[49025] = a[14] & g[32641];
assign g[65408] = b[14] & g[32641];
assign g[49026] = a[14] & g[32642];
assign g[65409] = b[14] & g[32642];
assign g[49027] = a[14] & g[32643];
assign g[65410] = b[14] & g[32643];
assign g[49028] = a[14] & g[32644];
assign g[65411] = b[14] & g[32644];
assign g[49029] = a[14] & g[32645];
assign g[65412] = b[14] & g[32645];
assign g[49030] = a[14] & g[32646];
assign g[65413] = b[14] & g[32646];
assign g[49031] = a[14] & g[32647];
assign g[65414] = b[14] & g[32647];
assign g[49032] = a[14] & g[32648];
assign g[65415] = b[14] & g[32648];
assign g[49033] = a[14] & g[32649];
assign g[65416] = b[14] & g[32649];
assign g[49034] = a[14] & g[32650];
assign g[65417] = b[14] & g[32650];
assign g[49035] = a[14] & g[32651];
assign g[65418] = b[14] & g[32651];
assign g[49036] = a[14] & g[32652];
assign g[65419] = b[14] & g[32652];
assign g[49037] = a[14] & g[32653];
assign g[65420] = b[14] & g[32653];
assign g[49038] = a[14] & g[32654];
assign g[65421] = b[14] & g[32654];
assign g[49039] = a[14] & g[32655];
assign g[65422] = b[14] & g[32655];
assign g[49040] = a[14] & g[32656];
assign g[65423] = b[14] & g[32656];
assign g[49041] = a[14] & g[32657];
assign g[65424] = b[14] & g[32657];
assign g[49042] = a[14] & g[32658];
assign g[65425] = b[14] & g[32658];
assign g[49043] = a[14] & g[32659];
assign g[65426] = b[14] & g[32659];
assign g[49044] = a[14] & g[32660];
assign g[65427] = b[14] & g[32660];
assign g[49045] = a[14] & g[32661];
assign g[65428] = b[14] & g[32661];
assign g[49046] = a[14] & g[32662];
assign g[65429] = b[14] & g[32662];
assign g[49047] = a[14] & g[32663];
assign g[65430] = b[14] & g[32663];
assign g[49048] = a[14] & g[32664];
assign g[65431] = b[14] & g[32664];
assign g[49049] = a[14] & g[32665];
assign g[65432] = b[14] & g[32665];
assign g[49050] = a[14] & g[32666];
assign g[65433] = b[14] & g[32666];
assign g[49051] = a[14] & g[32667];
assign g[65434] = b[14] & g[32667];
assign g[49052] = a[14] & g[32668];
assign g[65435] = b[14] & g[32668];
assign g[49053] = a[14] & g[32669];
assign g[65436] = b[14] & g[32669];
assign g[49054] = a[14] & g[32670];
assign g[65437] = b[14] & g[32670];
assign g[49055] = a[14] & g[32671];
assign g[65438] = b[14] & g[32671];
assign g[49056] = a[14] & g[32672];
assign g[65439] = b[14] & g[32672];
assign g[49057] = a[14] & g[32673];
assign g[65440] = b[14] & g[32673];
assign g[49058] = a[14] & g[32674];
assign g[65441] = b[14] & g[32674];
assign g[49059] = a[14] & g[32675];
assign g[65442] = b[14] & g[32675];
assign g[49060] = a[14] & g[32676];
assign g[65443] = b[14] & g[32676];
assign g[49061] = a[14] & g[32677];
assign g[65444] = b[14] & g[32677];
assign g[49062] = a[14] & g[32678];
assign g[65445] = b[14] & g[32678];
assign g[49063] = a[14] & g[32679];
assign g[65446] = b[14] & g[32679];
assign g[49064] = a[14] & g[32680];
assign g[65447] = b[14] & g[32680];
assign g[49065] = a[14] & g[32681];
assign g[65448] = b[14] & g[32681];
assign g[49066] = a[14] & g[32682];
assign g[65449] = b[14] & g[32682];
assign g[49067] = a[14] & g[32683];
assign g[65450] = b[14] & g[32683];
assign g[49068] = a[14] & g[32684];
assign g[65451] = b[14] & g[32684];
assign g[49069] = a[14] & g[32685];
assign g[65452] = b[14] & g[32685];
assign g[49070] = a[14] & g[32686];
assign g[65453] = b[14] & g[32686];
assign g[49071] = a[14] & g[32687];
assign g[65454] = b[14] & g[32687];
assign g[49072] = a[14] & g[32688];
assign g[65455] = b[14] & g[32688];
assign g[49073] = a[14] & g[32689];
assign g[65456] = b[14] & g[32689];
assign g[49074] = a[14] & g[32690];
assign g[65457] = b[14] & g[32690];
assign g[49075] = a[14] & g[32691];
assign g[65458] = b[14] & g[32691];
assign g[49076] = a[14] & g[32692];
assign g[65459] = b[14] & g[32692];
assign g[49077] = a[14] & g[32693];
assign g[65460] = b[14] & g[32693];
assign g[49078] = a[14] & g[32694];
assign g[65461] = b[14] & g[32694];
assign g[49079] = a[14] & g[32695];
assign g[65462] = b[14] & g[32695];
assign g[49080] = a[14] & g[32696];
assign g[65463] = b[14] & g[32696];
assign g[49081] = a[14] & g[32697];
assign g[65464] = b[14] & g[32697];
assign g[49082] = a[14] & g[32698];
assign g[65465] = b[14] & g[32698];
assign g[49083] = a[14] & g[32699];
assign g[65466] = b[14] & g[32699];
assign g[49084] = a[14] & g[32700];
assign g[65467] = b[14] & g[32700];
assign g[49085] = a[14] & g[32701];
assign g[65468] = b[14] & g[32701];
assign g[49086] = a[14] & g[32702];
assign g[65469] = b[14] & g[32702];
assign g[49087] = a[14] & g[32703];
assign g[65470] = b[14] & g[32703];
assign g[49088] = a[14] & g[32704];
assign g[65471] = b[14] & g[32704];
assign g[49089] = a[14] & g[32705];
assign g[65472] = b[14] & g[32705];
assign g[49090] = a[14] & g[32706];
assign g[65473] = b[14] & g[32706];
assign g[49091] = a[14] & g[32707];
assign g[65474] = b[14] & g[32707];
assign g[49092] = a[14] & g[32708];
assign g[65475] = b[14] & g[32708];
assign g[49093] = a[14] & g[32709];
assign g[65476] = b[14] & g[32709];
assign g[49094] = a[14] & g[32710];
assign g[65477] = b[14] & g[32710];
assign g[49095] = a[14] & g[32711];
assign g[65478] = b[14] & g[32711];
assign g[49096] = a[14] & g[32712];
assign g[65479] = b[14] & g[32712];
assign g[49097] = a[14] & g[32713];
assign g[65480] = b[14] & g[32713];
assign g[49098] = a[14] & g[32714];
assign g[65481] = b[14] & g[32714];
assign g[49099] = a[14] & g[32715];
assign g[65482] = b[14] & g[32715];
assign g[49100] = a[14] & g[32716];
assign g[65483] = b[14] & g[32716];
assign g[49101] = a[14] & g[32717];
assign g[65484] = b[14] & g[32717];
assign g[49102] = a[14] & g[32718];
assign g[65485] = b[14] & g[32718];
assign g[49103] = a[14] & g[32719];
assign g[65486] = b[14] & g[32719];
assign g[49104] = a[14] & g[32720];
assign g[65487] = b[14] & g[32720];
assign g[49105] = a[14] & g[32721];
assign g[65488] = b[14] & g[32721];
assign g[49106] = a[14] & g[32722];
assign g[65489] = b[14] & g[32722];
assign g[49107] = a[14] & g[32723];
assign g[65490] = b[14] & g[32723];
assign g[49108] = a[14] & g[32724];
assign g[65491] = b[14] & g[32724];
assign g[49109] = a[14] & g[32725];
assign g[65492] = b[14] & g[32725];
assign g[49110] = a[14] & g[32726];
assign g[65493] = b[14] & g[32726];
assign g[49111] = a[14] & g[32727];
assign g[65494] = b[14] & g[32727];
assign g[49112] = a[14] & g[32728];
assign g[65495] = b[14] & g[32728];
assign g[49113] = a[14] & g[32729];
assign g[65496] = b[14] & g[32729];
assign g[49114] = a[14] & g[32730];
assign g[65497] = b[14] & g[32730];
assign g[49115] = a[14] & g[32731];
assign g[65498] = b[14] & g[32731];
assign g[49116] = a[14] & g[32732];
assign g[65499] = b[14] & g[32732];
assign g[49117] = a[14] & g[32733];
assign g[65500] = b[14] & g[32733];
assign g[49118] = a[14] & g[32734];
assign g[65501] = b[14] & g[32734];
assign g[49119] = a[14] & g[32735];
assign g[65502] = b[14] & g[32735];
assign g[49120] = a[14] & g[32736];
assign g[65503] = b[14] & g[32736];
assign g[49121] = a[14] & g[32737];
assign g[65504] = b[14] & g[32737];
assign g[49122] = a[14] & g[32738];
assign g[65505] = b[14] & g[32738];
assign g[49123] = a[14] & g[32739];
assign g[65506] = b[14] & g[32739];
assign g[49124] = a[14] & g[32740];
assign g[65507] = b[14] & g[32740];
assign g[49125] = a[14] & g[32741];
assign g[65508] = b[14] & g[32741];
assign g[49126] = a[14] & g[32742];
assign g[65509] = b[14] & g[32742];
assign g[49127] = a[14] & g[32743];
assign g[65510] = b[14] & g[32743];
assign g[49128] = a[14] & g[32744];
assign g[65511] = b[14] & g[32744];
assign g[49129] = a[14] & g[32745];
assign g[65512] = b[14] & g[32745];
assign g[49130] = a[14] & g[32746];
assign g[65513] = b[14] & g[32746];
assign g[49131] = a[14] & g[32747];
assign g[65514] = b[14] & g[32747];
assign g[49132] = a[14] & g[32748];
assign g[65515] = b[14] & g[32748];
assign g[49133] = a[14] & g[32749];
assign g[65516] = b[14] & g[32749];
assign g[49134] = a[14] & g[32750];
assign g[65517] = b[14] & g[32750];
assign g[49135] = a[14] & g[32751];
assign g[65518] = b[14] & g[32751];
endmodule