
module gen_linear_part ( a, b, n, s );
  input [5:0] a;
  input [5:0] b;
  input [118:0] n;
  output [5:0] s;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41;

  XOR3D0 U1 ( .A1(n1), .A2(n2), .A3(n[118]), .Z(s[5]) );
  XOR4D0 U2 ( .A1(a[5]), .A2(n3), .A3(n[113]), .A4(b[5]), .Z(n2) );
  XOR4D0 U3 ( .A1(n[108]), .A2(n[107]), .A3(n4), .A4(n5), .Z(n3) );
  XOR3D0 U4 ( .A1(n6), .A2(n7), .A3(n[106]), .Z(n5) );
  XOR4D0 U5 ( .A1(n[100]), .A2(n8), .A3(n[102]), .A4(n[101]), .Z(n7) );
  XOR4D0 U6 ( .A1(n[94]), .A2(n[93]), .A3(n9), .A4(n10), .Z(n8) );
  XOR3D0 U7 ( .A1(n11), .A2(n12), .A3(n[92]), .Z(n10) );
  XOR4D0 U8 ( .A1(n[85]), .A2(n13), .A3(n[87]), .A4(n[86]), .Z(n12) );
  XOR4D0 U9 ( .A1(n[80]), .A2(n[79]), .A3(n14), .A4(n15), .Z(n13) );
  XOR3D0 U10 ( .A1(n16), .A2(n17), .A3(n[78]), .Z(n15) );
  XOR4D0 U11 ( .A1(n[71]), .A2(n18), .A3(n[73]), .A4(n[72]), .Z(n17) );
  XOR4D0 U12 ( .A1(n[66]), .A2(n[65]), .A3(n19), .A4(n20), .Z(n18) );
  XOR3D0 U13 ( .A1(n21), .A2(n22), .A3(n[64]), .Z(n20) );
  XOR4D0 U14 ( .A1(n[57]), .A2(n[56]), .A3(n[59]), .A4(n[58]), .Z(n22) );
  XOR4D0 U15 ( .A1(n[61]), .A2(n[60]), .A3(n[63]), .A4(n[62]), .Z(n21) );
  XOR4D0 U16 ( .A1(n[68]), .A2(n[67]), .A3(n[70]), .A4(n[69]), .Z(n19) );
  XOR4D0 U17 ( .A1(n[75]), .A2(n[74]), .A3(n[77]), .A4(n[76]), .Z(n16) );
  XOR4D0 U18 ( .A1(n[82]), .A2(n[81]), .A3(n[84]), .A4(n[83]), .Z(n14) );
  XOR4D0 U19 ( .A1(n[89]), .A2(n[88]), .A3(n[91]), .A4(n[90]), .Z(n11) );
  XOR4D0 U20 ( .A1(n[96]), .A2(n[95]), .A3(n[98]), .A4(n[97]), .Z(n9) );
  XOR4D0 U21 ( .A1(n[104]), .A2(n[103]), .A3(n[99]), .A4(n[105]), .Z(n6) );
  XOR4D0 U22 ( .A1(n[110]), .A2(n[109]), .A3(n[112]), .A4(n[111]), .Z(n4) );
  XOR4D0 U23 ( .A1(n[115]), .A2(n[114]), .A3(n[117]), .A4(n[116]), .Z(n1) );
  XOR4D0 U24 ( .A1(n23), .A2(n24), .A3(n25), .A4(n[50]), .Z(s[4]) );
  XOR3D0 U25 ( .A1(n[53]), .A2(n[52]), .A3(n[51]), .Z(n25) );
  XOR4D0 U26 ( .A1(a[4]), .A2(n26), .A3(n[47]), .A4(b[4]), .Z(n24) );
  XOR4D0 U27 ( .A1(n[42]), .A2(n[41]), .A3(n27), .A4(n28), .Z(n26) );
  XOR3D0 U28 ( .A1(n29), .A2(n30), .A3(n[40]), .Z(n28) );
  XOR3D0 U29 ( .A1(n[35]), .A2(n[34]), .A3(n31), .Z(n30) );
  XOR3D0 U30 ( .A1(n32), .A2(n33), .A3(n[33]), .Z(n31) );
  XOR4D0 U31 ( .A1(n[26]), .A2(n[25]), .A3(n[28]), .A4(n[27]), .Z(n33) );
  XOR4D0 U32 ( .A1(n[30]), .A2(n[29]), .A3(n[32]), .A4(n[31]), .Z(n32) );
  XOR4D0 U33 ( .A1(n[37]), .A2(n[36]), .A3(n[39]), .A4(n[38]), .Z(n29) );
  XOR4D0 U34 ( .A1(n[44]), .A2(n[43]), .A3(n[46]), .A4(n[45]), .Z(n27) );
  XOR4D0 U35 ( .A1(n[49]), .A2(n[48]), .A3(n[55]), .A4(n[54]), .Z(n23) );
  XOR4D0 U36 ( .A1(b[3]), .A2(a[3]), .A3(n34), .A4(n35), .Z(s[3]) );
  XOR3D0 U37 ( .A1(n[20]), .A2(n[19]), .A3(n36), .Z(n35) );
  XOR3D0 U38 ( .A1(n37), .A2(n38), .A3(n[18]), .Z(n36) );
  XOR4D0 U39 ( .A1(n[11]), .A2(n[10]), .A3(n[13]), .A4(n[12]), .Z(n38) );
  XOR4D0 U40 ( .A1(n[15]), .A2(n[14]), .A3(n[17]), .A4(n[16]), .Z(n37) );
  XOR4D0 U41 ( .A1(n[22]), .A2(n[21]), .A3(n[24]), .A4(n[23]), .Z(n34) );
  XOR3D0 U42 ( .A1(n39), .A2(n40), .A3(n[9]), .Z(s[2]) );
  XOR4D0 U43 ( .A1(b[2]), .A2(a[2]), .A3(n[4]), .A4(n[3]), .Z(n40) );
  XOR4D0 U44 ( .A1(n[6]), .A2(n[5]), .A3(n[8]), .A4(n[7]), .Z(n39) );
  XOR3D0 U45 ( .A1(b[1]), .A2(a[1]), .A3(n41), .Z(s[1]) );
  XOR3D0 U46 ( .A1(n[2]), .A2(n[1]), .A3(n[0]), .Z(n41) );
  XOR2D0 U47 ( .A1(b[0]), .A2(a[0]), .Z(s[0]) );
endmodule


module gen_nonlinear_part ( a, b, n );
  input [5:0] a;
  input [5:0] b;
  output [118:0] n;


  INVD0 U2 ( .I(1'b1), .ZN(n[1]) );
  INVD0 U4 ( .I(1'b1), .ZN(n[2]) );
  INVD0 U6 ( .I(1'b1), .ZN(n[5]) );
  INVD0 U8 ( .I(1'b1), .ZN(n[6]) );
  INVD0 U10 ( .I(1'b1), .ZN(n[8]) );
  INVD0 U12 ( .I(1'b1), .ZN(n[9]) );
  INVD0 U14 ( .I(1'b1), .ZN(n[13]) );
  INVD0 U16 ( .I(1'b1), .ZN(n[14]) );
  INVD0 U18 ( .I(1'b1), .ZN(n[16]) );
  INVD0 U20 ( .I(1'b1), .ZN(n[17]) );
  INVD0 U22 ( .I(1'b1), .ZN(n[20]) );
  INVD0 U24 ( .I(1'b1), .ZN(n[21]) );
  INVD0 U26 ( .I(1'b1), .ZN(n[23]) );
  INVD0 U28 ( .I(1'b1), .ZN(n[24]) );
  INVD0 U30 ( .I(1'b1), .ZN(n[29]) );
  INVD0 U32 ( .I(1'b1), .ZN(n[30]) );
  INVD0 U34 ( .I(1'b1), .ZN(n[32]) );
  INVD0 U36 ( .I(1'b1), .ZN(n[33]) );
  INVD0 U38 ( .I(1'b1), .ZN(n[36]) );
  INVD0 U40 ( .I(1'b1), .ZN(n[37]) );
  INVD0 U42 ( .I(1'b1), .ZN(n[39]) );
  INVD0 U44 ( .I(1'b1), .ZN(n[40]) );
  INVD0 U46 ( .I(1'b1), .ZN(n[44]) );
  INVD0 U48 ( .I(1'b1), .ZN(n[45]) );
  INVD0 U50 ( .I(1'b1), .ZN(n[47]) );
  INVD0 U52 ( .I(1'b1), .ZN(n[48]) );
  INVD0 U54 ( .I(1'b1), .ZN(n[51]) );
  INVD0 U56 ( .I(1'b1), .ZN(n[52]) );
  INVD0 U58 ( .I(1'b1), .ZN(n[54]) );
  INVD0 U61 ( .I(1'b1), .ZN(n[55]) );
  INVD0 U63 ( .I(1'b1), .ZN(n[61]) );
  INVD0 U65 ( .I(1'b1), .ZN(n[62]) );
  INVD0 U67 ( .I(1'b1), .ZN(n[64]) );
  INVD0 U69 ( .I(1'b1), .ZN(n[65]) );
  INVD0 U71 ( .I(1'b1), .ZN(n[68]) );
  INVD0 U73 ( .I(1'b1), .ZN(n[69]) );
  INVD0 U75 ( .I(1'b1), .ZN(n[71]) );
  INVD0 U77 ( .I(1'b1), .ZN(n[72]) );
  INVD0 U79 ( .I(1'b1), .ZN(n[76]) );
  INVD0 U81 ( .I(1'b1), .ZN(n[77]) );
  INVD0 U83 ( .I(1'b1), .ZN(n[79]) );
  INVD0 U85 ( .I(1'b1), .ZN(n[80]) );
  INVD0 U87 ( .I(1'b1), .ZN(n[83]) );
  INVD0 U89 ( .I(1'b1), .ZN(n[84]) );
  INVD0 U91 ( .I(1'b1), .ZN(n[86]) );
  INVD0 U93 ( .I(1'b1), .ZN(n[87]) );
  INVD0 U95 ( .I(1'b1), .ZN(n[92]) );
  INVD0 U97 ( .I(1'b1), .ZN(n[93]) );
  INVD0 U99 ( .I(1'b1), .ZN(n[95]) );
  INVD0 U101 ( .I(1'b1), .ZN(n[96]) );
  INVD0 U103 ( .I(1'b1), .ZN(n[99]) );
  INVD0 U105 ( .I(1'b1), .ZN(n[100]) );
  INVD0 U107 ( .I(1'b1), .ZN(n[102]) );
  INVD0 U109 ( .I(1'b1), .ZN(n[103]) );
  INVD0 U111 ( .I(1'b1), .ZN(n[107]) );
  INVD0 U113 ( .I(1'b1), .ZN(n[108]) );
  INVD0 U115 ( .I(1'b1), .ZN(n[110]) );
  INVD0 U117 ( .I(1'b1), .ZN(n[111]) );
  INVD0 U119 ( .I(1'b1), .ZN(n[114]) );
  INVD0 U121 ( .I(1'b1), .ZN(n[115]) );
  INVD0 U123 ( .I(1'b1), .ZN(n[117]) );
  INVD0 U125 ( .I(1'b1), .ZN(n[118]) );
  AN2D0 U127 ( .A1(b[4]), .A2(n[35]), .Z(n[98]) );
  AN2D0 U128 ( .A1(n[34]), .A2(b[4]), .Z(n[97]) );
  AN2D0 U129 ( .A1(n[31]), .A2(b[4]), .Z(n[94]) );
  AN2D0 U130 ( .A1(n[28]), .A2(b[4]), .Z(n[91]) );
  AN2D0 U131 ( .A1(n[27]), .A2(b[4]), .Z(n[90]) );
  AN2D0 U132 ( .A1(n[26]), .A2(b[4]), .Z(n[89]) );
  AN2D0 U133 ( .A1(n[25]), .A2(b[4]), .Z(n[88]) );
  AN2D0 U134 ( .A1(a[4]), .A2(n[53]), .Z(n[85]) );
  AN2D0 U135 ( .A1(n[50]), .A2(a[4]), .Z(n[82]) );
  AN2D0 U136 ( .A1(n[49]), .A2(a[4]), .Z(n[81]) );
  AN2D0 U137 ( .A1(n[46]), .A2(a[4]), .Z(n[78]) );
  AN2D0 U138 ( .A1(n[43]), .A2(a[4]), .Z(n[75]) );
  AN2D0 U139 ( .A1(n[42]), .A2(a[4]), .Z(n[74]) );
  AN2D0 U140 ( .A1(n[41]), .A2(a[4]), .Z(n[73]) );
  AN2D0 U141 ( .A1(n[38]), .A2(a[4]), .Z(n[70]) );
  AN2D0 U142 ( .A1(a[4]), .A2(n[35]), .Z(n[67]) );
  AN2D0 U143 ( .A1(a[4]), .A2(n[34]), .Z(n[66]) );
  AN2D0 U144 ( .A1(a[4]), .A2(n[31]), .Z(n[63]) );
  AN2D0 U145 ( .A1(a[4]), .A2(n[28]), .Z(n[60]) );
  AN2D0 U146 ( .A1(a[4]), .A2(n[27]), .Z(n[59]) );
  AN2D0 U147 ( .A1(a[4]), .A2(n[26]), .Z(n[58]) );
  AN2D0 U148 ( .A1(a[4]), .A2(n[25]), .Z(n[57]) );
  AN2D0 U149 ( .A1(a[4]), .A2(b[4]), .Z(n[56]) );
  AN2D0 U150 ( .A1(n[19]), .A2(a[3]), .Z(n[35]) );
  AN2D0 U151 ( .A1(a[3]), .A2(n[18]), .Z(n[34]) );
  AN2D0 U152 ( .A1(a[3]), .A2(n[15]), .Z(n[31]) );
  AN2D0 U153 ( .A1(a[3]), .A2(n[12]), .Z(n[28]) );
  AN2D0 U154 ( .A1(a[3]), .A2(n[11]), .Z(n[27]) );
  AN2D0 U155 ( .A1(a[3]), .A2(n[10]), .Z(n[26]) );
  AN2D0 U156 ( .A1(a[3]), .A2(b[3]), .Z(n[25]) );
  AN2D0 U157 ( .A1(n[53]), .A2(b[4]), .Z(n[116]) );
  AN2D0 U158 ( .A1(b[3]), .A2(n[22]), .Z(n[53]) );
  AN2D0 U159 ( .A1(n[50]), .A2(b[4]), .Z(n[113]) );
  AN2D0 U160 ( .A1(n[19]), .A2(b[3]), .Z(n[50]) );
  AN2D0 U161 ( .A1(n[4]), .A2(b[2]), .Z(n[19]) );
  AN2D0 U162 ( .A1(n[49]), .A2(b[4]), .Z(n[112]) );
  AN2D0 U163 ( .A1(n[18]), .A2(b[3]), .Z(n[49]) );
  AN2D0 U164 ( .A1(b[2]), .A2(n[3]), .Z(n[18]) );
  AN2D0 U165 ( .A1(n[46]), .A2(b[4]), .Z(n[109]) );
  AN2D0 U166 ( .A1(n[15]), .A2(b[3]), .Z(n[46]) );
  AN2D0 U167 ( .A1(n[7]), .A2(a[2]), .Z(n[15]) );
  AN2D0 U168 ( .A1(n[43]), .A2(b[4]), .Z(n[106]) );
  AN2D0 U169 ( .A1(n[12]), .A2(b[3]), .Z(n[43]) );
  AN2D0 U170 ( .A1(n[4]), .A2(a[2]), .Z(n[12]) );
  AN2D0 U171 ( .A1(n[0]), .A2(a[1]), .Z(n[4]) );
  AN2D0 U172 ( .A1(n[42]), .A2(b[4]), .Z(n[105]) );
  AN2D0 U173 ( .A1(n[11]), .A2(b[3]), .Z(n[42]) );
  AN2D0 U174 ( .A1(n[3]), .A2(a[2]), .Z(n[11]) );
  AN2D0 U175 ( .A1(a[1]), .A2(b[1]), .Z(n[3]) );
  AN2D0 U176 ( .A1(n[41]), .A2(b[4]), .Z(n[104]) );
  AN2D0 U177 ( .A1(n[10]), .A2(b[3]), .Z(n[41]) );
  AN2D0 U178 ( .A1(b[2]), .A2(a[2]), .Z(n[10]) );
  AN2D0 U179 ( .A1(n[38]), .A2(b[4]), .Z(n[101]) );
  AN2D0 U180 ( .A1(a[3]), .A2(n[22]), .Z(n[38]) );
  AN2D0 U181 ( .A1(b[2]), .A2(n[7]), .Z(n[22]) );
  AN2D0 U182 ( .A1(n[0]), .A2(b[1]), .Z(n[7]) );
  AN2D0 U183 ( .A1(b[0]), .A2(a[0]), .Z(n[0]) );
endmodule


module gen_cla_decomposed ( a, b, s );
  input [5:0] a;
  input [5:0] b;
  output [5:0] s;

  wire   [118:0] n;

  gen_nonlinear_part NLIN ( .a(a), .b(b), .n(n) );
  gen_linear_part LIN ( .a(a), .b(b), .n({1'b0, 1'b0, n[116], 1'b0, 1'b0, 
        n[113:112], 1'b0, 1'b0, n[109], 1'b0, 1'b0, n[106:104], 1'b0, 1'b0, 
        n[101], 1'b0, 1'b0, n[98:97], 1'b0, 1'b0, n[94], 1'b0, 1'b0, n[91:88], 
        1'b0, 1'b0, n[85], 1'b0, 1'b0, n[82:81], 1'b0, 1'b0, n[78], 1'b0, 1'b0, 
        n[75:73], 1'b0, 1'b0, n[70], 1'b0, 1'b0, n[67:66], 1'b0, 1'b0, n[63], 
        1'b0, 1'b0, n[60:56], 1'b0, 1'b0, n[53], 1'b0, 1'b0, n[50:49], 1'b0, 
        1'b0, n[46], 1'b0, 1'b0, n[43:41], 1'b0, 1'b0, n[38], 1'b0, 1'b0, 
        n[35:34], 1'b0, 1'b0, n[31], 1'b0, 1'b0, n[28:25], 1'b0, 1'b0, n[22], 
        1'b0, 1'b0, n[19:18], 1'b0, 1'b0, n[15], 1'b0, 1'b0, n[12:10], 1'b0, 
        1'b0, n[7], 1'b0, 1'b0, n[4:3], 1'b0, 1'b0, n[0]}), .s(s) );
endmodule

