module nonlin_mapped(n__0, n__1, n__2, n__3, n__4, n__5, n__6, n__7, n__8, n__9, n__10, n__11, n__12, n__13, n__14, n__15, n__16, n__17, n__18, n__19, n__20, n__21, n__22, n__23, n__24, n__25, n__26, n__27, n__28, n__29, n__30, n__31, n__32, n__33, n__34, n__35, n__36, n__37, n__38, n__39, n__40, n__41, n__42, n__43, n__44, n__45, n__46, n__47, n__48, n__49, n__50, n__51, n__52, n__53, n__54, n__55, n__56, n__57, n__58, n__59, n__60, n__61, n__62, n__63, n__64, n__65, n__66, n__67, n__68, n__69, n__70, n__71, n__72, n__73, n__74, n__75, n__76, n__77, n__78, n__79, n__80, n__81, n__82, n__83, n__84, n__85, n__86, n__87, n__88, n__89, n__90, n__91, n__92, n__93, n__94, n__95, n__96, n__97, n__98, n__99, n__100, n__101, n__102, n__103, n__104, n__105, n__106, n__107, n__108, n__109, n__110, n__111, n__112, n__113, n__114, n__115, n__116, n__117, n__118, n__119, n__120, n__121, n__122, n__123, n__124, n__125, n__126, n__127, n__128, n__129, n__130, n__131, n__132, n__133, n__134, n__135, n__136, n__137, n__138, n__139, n__140, n__141, n__142, n__143, n__144, n__145, n__146, n__147, n__148, n__149, n__150, n__151, n__152, n__153, n__154, n__155, n__156, n__157, n__158, n__159, n__160, n__161, n__162, n__163, n__164, n__165, n__166, n__167, n__168, n__169, n__170, n__171, n__172, n__173, n__174, n__175, n__176, n__177, n__178, n__179, n__180, n__181, n__182, n__183, n__184, n__185, n__186, n__187, n__188, n__189, n__190, n__191, n__192, n__193, n__194, n__195, n__196, n__197, n__198, n__199, n__200, n__201, n__202, n__203, n__204, n__205, n__206, n__207, n__208, n__209, n__210, n__211, n__212, n__213, n__214, n__215, n__216, n__217, n__218, n__219, n__220, n__221, n__222, n__223, n__224, n__225, n__226, n__227, n__228, n__229, n__230, n__231, n__232, n__233, n__234, n__235, n__236, n__237, n__238, n__239, n__240, n__241, n__242, n__243, n__244, n__245, n__246, n__247, n__248, n__249, n__250, n__251, n__252, n__253, n__254, n__255, n__256, n__257, n__258, n__259, n__260, n__261, n__262, n__263, n__264, n__265, n__266, n__267, n__268, n__269, n__270, n__271, n__272, n__273, n__274, n__275, n__276, n__277, n__278, n__279, n__280, n__281, n__282, n__283, n__284, n__285, n__286, n__287, n__288, n__289, n__290, n__291, n__292, n__293, n__294, n__295, n__296, n__297, n__298, n__299, n__300, n__301, n__302, n__303, n__304, n__305, n__306, n__307, n__308, n__309, n__310, n__311, n__312, n__313, n__314, n__315, n__316, n__317, n__318, n__319, n__320, n__321, n__322, n__323, n__324, n__325, n__326, n__327, n__328, n__329, n__330, n__331, n__332, n__333, n__334, n__335, n__336, n__337, n__338, n__339, n__340, n__341, n__342, n__343, n__344, n__345, n__346, n__347, n__348, n__349, n__350, n__351, n__352, n__353, n__354, n__355, n__356, n__357, n__358, n__359, n__360, n__361, n__362, n__363, n__364, n__365, n__366, n__367, n__368, n__369, n__370, n__371, n__372, n__373, n__374, n__375, n__376, n__377, n__378, n__379, n__380, n__381, n__382, n__383, n__384, n__385, n__386, n__387, n__388, n__389, n__390, n__391, n__392, n__393, n__394, n__395, n__396, n__397, n__398, n__399, n__400, n__401, n__402, n__403, n__404, n__405, n__406, n__407, n__408, n__409, n__410, n__411, n__412, n__413, n__414, n__415, n__416, n__417, n__418, n__419, n__420, n__421, n__422, n__423, n__424, n__425, n__426, n__427, n__428, n__429, n__430, n__431, n__432, n__433, n__434, n__435, n__436, n__437, n__438, n__439, n__440, n__441, n__442, n__443, n__444, n__445, n__446, n__447, n__448, n__449, n__450, n__451, n__452, n__453, n__454, n__455, n__456, n__457, n__458, n__459, n__460, n__461, n__462, n__463, n__464, n__465, n__466, n__467, n__468, n__469, n__470, n__471, n__472, n__473, n__474, n__475, n__476, n__477, n__478, n__479, n__480, n__481, n__482, n__483, n__484, n__485, n__486, n__487, n__488, n__489, n__490, n__491, n__492, n__493, n__494, n__495, n__496, n__497, n__498, n__499, n__500, a__0, a__1, a__2, a__3, a__4, a__5, a__6, b__0, b__1, b__2, b__3, b__4, b__5, b__6, c);
  input a__0, a__1, a__2, a__3, a__4, a__5, a__6, b__0, b__1, b__2, b__3, b__4, b__5, b__6, c;
  output n__0, n__1, n__2, n__3, n__4, n__5, n__6, n__7, n__8, n__9, n__10, n__11, n__12, n__13, n__14, n__15, n__16, n__17, n__18, n__19, n__20, n__21, n__22, n__23, n__24, n__25, n__26, n__27, n__28, n__29, n__30, n__31, n__32, n__33, n__34, n__35, n__36, n__37, n__38, n__39, n__40, n__41, n__42, n__43, n__44, n__45, n__46, n__47, n__48, n__49, n__50, n__51, n__52, n__53, n__54, n__55, n__56, n__57, n__58, n__59, n__60, n__61, n__62, n__63, n__64, n__65, n__66, n__67, n__68, n__69, n__70, n__71, n__72, n__73, n__74, n__75, n__76, n__77, n__78, n__79, n__80, n__81, n__82, n__83, n__84, n__85, n__86, n__87, n__88, n__89, n__90, n__91, n__92, n__93, n__94, n__95, n__96, n__97, n__98, n__99, n__100, n__101, n__102, n__103, n__104, n__105, n__106, n__107, n__108, n__109, n__110, n__111, n__112, n__113, n__114, n__115, n__116, n__117, n__118, n__119, n__120, n__121, n__122, n__123, n__124, n__125, n__126, n__127, n__128, n__129, n__130, n__131, n__132, n__133, n__134, n__135, n__136, n__137, n__138, n__139, n__140, n__141, n__142, n__143, n__144, n__145, n__146, n__147, n__148, n__149, n__150, n__151, n__152, n__153, n__154, n__155, n__156, n__157, n__158, n__159, n__160, n__161, n__162, n__163, n__164, n__165, n__166, n__167, n__168, n__169, n__170, n__171, n__172, n__173, n__174, n__175, n__176, n__177, n__178, n__179, n__180, n__181, n__182, n__183, n__184, n__185, n__186, n__187, n__188, n__189, n__190, n__191, n__192, n__193, n__194, n__195, n__196, n__197, n__198, n__199, n__200, n__201, n__202, n__203, n__204, n__205, n__206, n__207, n__208, n__209, n__210, n__211, n__212, n__213, n__214, n__215, n__216, n__217, n__218, n__219, n__220, n__221, n__222, n__223, n__224, n__225, n__226, n__227, n__228, n__229, n__230, n__231, n__232, n__233, n__234, n__235, n__236, n__237, n__238, n__239, n__240, n__241, n__242, n__243, n__244, n__245, n__246, n__247, n__248, n__249, n__250, n__251, n__252, n__253, n__254, n__255, n__256, n__257, n__258, n__259, n__260, n__261, n__262, n__263, n__264, n__265, n__266, n__267, n__268, n__269, n__270, n__271, n__272, n__273, n__274, n__275, n__276, n__277, n__278, n__279, n__280, n__281, n__282, n__283, n__284, n__285, n__286, n__287, n__288, n__289, n__290, n__291, n__292, n__293, n__294, n__295, n__296, n__297, n__298, n__299, n__300, n__301, n__302, n__303, n__304, n__305, n__306, n__307, n__308, n__309, n__310, n__311, n__312, n__313, n__314, n__315, n__316, n__317, n__318, n__319, n__320, n__321, n__322, n__323, n__324, n__325, n__326, n__327, n__328, n__329, n__330, n__331, n__332, n__333, n__334, n__335, n__336, n__337, n__338, n__339, n__340, n__341, n__342, n__343, n__344, n__345, n__346, n__347, n__348, n__349, n__350, n__351, n__352, n__353, n__354, n__355, n__356, n__357, n__358, n__359, n__360, n__361, n__362, n__363, n__364, n__365, n__366, n__367, n__368, n__369, n__370, n__371, n__372, n__373, n__374, n__375, n__376, n__377, n__378, n__379, n__380, n__381, n__382, n__383, n__384, n__385, n__386, n__387, n__388, n__389, n__390, n__391, n__392, n__393, n__394, n__395, n__396, n__397, n__398, n__399, n__400, n__401, n__402, n__403, n__404, n__405, n__406, n__407, n__408, n__409, n__410, n__411, n__412, n__413, n__414, n__415, n__416, n__417, n__418, n__419, n__420, n__421, n__422, n__423, n__424, n__425, n__426, n__427, n__428, n__429, n__430, n__431, n__432, n__433, n__434, n__435, n__436, n__437, n__438, n__439, n__440, n__441, n__442, n__443, n__444, n__445, n__446, n__447, n__448, n__449, n__450, n__451, n__452, n__453, n__454, n__455, n__456, n__457, n__458, n__459, n__460, n__461, n__462, n__463, n__464, n__465, n__466, n__467, n__468, n__469, n__470, n__471, n__472, n__473, n__474, n__475, n__476, n__477, n__478, n__479, n__480, n__481, n__482, n__483, n__484, n__485, n__486, n__487, n__488, n__489, n__490, n__491, n__492, n__493, n__494, n__495, n__496, n__497, n__498, n__499, n__500;

  wire   n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,         n654;
  assign n423 = ~b__6;
  assign n424 = ~b__6;
  assign n425 = ~b__6;
  assign n426 = ~b__6;
  assign n427 = ~b__6;
  assign n428 = ~b__6;
  assign n429 = ~b__6;
  assign n430 = ~b__6;
  assign n431 = ~b__6;
  assign n432 = ~b__6;
  assign n433 = ~a__6;
  assign n434 = ~a__6;
  assign n435 = ~a__6;
  assign n436 = ~a__6;
  assign n437 = ~a__6;
  assign n438 = ~a__6;
  assign n439 = ~a__6;
  assign n440 = ~a__6;
  assign n441 = ~a__6;
  assign n442 = ~a__6;
  assign n__500 = ~(n443 | n432);
  assign n__499 = ~(n432 | n444);
  assign n__498 = ~(n432 | n445);
  assign n__497 = ~(n432 | n446);
  assign n__496 = ~(n432 | n447);
  assign n__495 = ~(n432 | n448);
  assign n__494 = ~(n432 | n449);
  assign n__493 = ~(n432 | n450);
  assign n__492 = ~(n432 | n451);
  assign n__491 = ~(n432 | n452);
  assign n__490 = ~(n432 | n453);
  assign n__489 = ~(n431 | n454);
  assign n__488 = ~(n431 | n455);
  assign n__487 = ~(n431 | n456);
  assign n__486 = ~(n431 | n457);
  assign n__485 = ~(n431 | n458);
  assign n__484 = ~(n431 | n459);
  assign n__483 = ~(n431 | n460);
  assign n__482 = ~(n431 | n461);
  assign n__481 = ~(n431 | n462);
  assign n__480 = ~(n431 | n463);
  assign n__479 = ~(n431 | n464);
  assign n__478 = ~(n431 | n465);
  assign n__477 = ~(n431 | n466);
  assign n__476 = ~(n430 | n467);
  assign n__475 = ~(n430 | n468);
  assign n__474 = ~(n430 | n469);
  assign n__473 = ~(n430 | n470);
  assign n__472 = ~(n430 | n471);
  assign n__471 = ~(n430 | n472);
  assign n__470 = ~(n430 | n473);
  assign n__469 = ~(n430 | n474);
  assign n__468 = ~(n430 | n475);
  assign n__467 = ~(n430 | n476);
  assign n__466 = ~(n430 | n477);
  assign n__465 = ~(n430 | n478);
  assign n__464 = ~(n430 | n479);
  assign n__463 = ~(n429 | n480);
  assign n__462 = ~(n429 | n481);
  assign n__461 = ~(n429 | n482);
  assign n__460 = ~(n429 | n483);
  assign n__459 = ~(n429 | n484);
  assign n__458 = ~(n429 | n485);
  assign n__457 = ~(n429 | n486);
  assign n__456 = ~(n429 | n487);
  assign n__455 = ~(n429 | n488);
  assign n__454 = ~(n429 | n489);
  assign n__453 = ~(n429 | n490);
  assign n__452 = ~(n429 | n491);
  assign n__451 = ~(n429 | n492);
  assign n__450 = ~(n428 | n493);
  assign n__449 = ~(n428 | n494);
  assign n__448 = ~(n428 | n495);
  assign n__447 = ~(n428 | n496);
  assign n__446 = ~(n428 | n497);
  assign n__445 = ~(n428 | n498);
  assign n__444 = ~(n428 | n499);
  assign n__443 = ~(n428 | n500);
  assign n__442 = ~(n428 | n501);
  assign n__441 = ~(n428 | n502);
  assign n__440 = ~(n428 | n503);
  assign n__439 = ~(n428 | n504);
  assign n__438 = ~(n428 | n505);
  assign n__437 = ~(n427 | n506);
  assign n__436 = ~(n427 | n507);
  assign n__435 = ~(n427 | n508);
  assign n__434 = ~(n427 | n509);
  assign n__433 = ~(n427 | n510);
  assign n__432 = ~(n427 | n511);
  assign n__431 = ~(n427 | n512);
  assign n__430 = ~(n427 | n513);
  assign n__429 = ~(n427 | n514);
  assign n__428 = ~(n427 | n515);
  assign n__427 = ~(n427 | n516);
  assign n__426 = ~(n427 | n517);
  assign n__425 = ~(n427 | n518);
  assign n__424 = ~(n426 | n519);
  assign n__423 = ~(n426 | n520);
  assign n__422 = ~(n426 | n521);
  assign n__421 = ~(n426 | n522);
  assign n__420 = ~(n426 | n523);
  assign n__419 = ~(n426 | n524);
  assign n__418 = ~(n426 | n525);
  assign n__417 = ~(n426 | n526);
  assign n__416 = ~(n426 | n527);
  assign n__415 = ~(n426 | n528);
  assign n__414 = ~(n426 | n529);
  assign n__413 = ~(n426 | n530);
  assign n__412 = ~(n426 | n531);
  assign n__411 = ~(n425 | n532);
  assign n__410 = ~(n425 | n533);
  assign n__409 = ~(n425 | n534);
  assign n__408 = ~(n425 | n535);
  assign n__407 = ~(n425 | n536);
  assign n__406 = ~(n425 | n537);
  assign n__405 = ~(n425 | n538);
  assign n__404 = ~(n425 | n539);
  assign n__403 = ~(n425 | n540);
  assign n__402 = ~(n425 | n541);
  assign n__401 = ~(n425 | n542);
  assign n__400 = ~(n425 | n543);
  assign n__399 = ~(n425 | n544);
  assign n__398 = ~(n424 | n545);
  assign n__397 = ~(n424 | n546);
  assign n__396 = ~(n424 | n547);
  assign n__395 = ~(n424 | n548);
  assign n__394 = ~(n424 | n549);
  assign n__393 = ~(n424 | n550);
  assign n__392 = ~(n424 | n551);
  assign n__391 = ~(n424 | n552);
  assign n__390 = ~(n424 | n553);
  assign n__389 = ~(n424 | n554);
  assign n__388 = ~(n424 | n555);
  assign n__387 = ~(n424 | n556);
  assign n__386 = ~(n424 | n557);
  assign n__385 = ~(n423 | n558);
  assign n__384 = ~(n423 | n559);
  assign n__383 = ~(n423 | n560);
  assign n__382 = ~(n423 | n561);
  assign n__381 = ~(n423 | n562);
  assign n__380 = ~(n423 | n563);
  assign n__379 = ~(n423 | n564);
  assign n__378 = ~(n423 | n565);
  assign n__377 = ~(n423 | n566);
  assign n__376 = ~(n423 | n567);
  assign n__375 = ~(n423 | n568);
  assign n__374 = ~(n423 | n569);
  assign n__373 = ~(n443 | n442);
  assign n__372 = ~(n444 | n442);
  assign n__371 = ~(n445 | n442);
  assign n__370 = ~(n446 | n442);
  assign n__369 = ~(n447 | n442);
  assign n__368 = ~(n448 | n442);
  assign n__367 = ~(n449 | n442);
  assign n__366 = ~(n450 | n442);
  assign n__365 = ~(n451 | n442);
  assign n__364 = ~(n452 | n442);
  assign n__363 = ~(n453 | n442);
  assign n__362 = ~(n454 | n441);
  assign n__361 = ~(n455 | n441);
  assign n__360 = ~(n456 | n441);
  assign n__359 = ~(n457 | n441);
  assign n__358 = ~(n458 | n441);
  assign n__357 = ~(n459 | n441);
  assign n__356 = ~(n460 | n441);
  assign n__355 = ~(n461 | n441);
  assign n__354 = ~(n462 | n441);
  assign n__353 = ~(n463 | n441);
  assign n__352 = ~(n464 | n441);
  assign n__351 = ~(n465 | n441);
  assign n__350 = ~(n466 | n441);
  assign n__349 = ~(n467 | n440);
  assign n__348 = ~(n468 | n440);
  assign n__347 = ~(n469 | n440);
  assign n__346 = ~(n470 | n440);
  assign n__345 = ~(n471 | n440);
  assign n__344 = ~(n472 | n440);
  assign n__343 = ~(n473 | n440);
  assign n__342 = ~(n474 | n440);
  assign n__341 = ~(n475 | n440);
  assign n__340 = ~(n476 | n440);
  assign n__339 = ~(n477 | n440);
  assign n__338 = ~(n478 | n440);
  assign n__337 = ~(n479 | n440);
  assign n__336 = ~(n480 | n439);
  assign n__335 = ~(n481 | n439);
  assign n__334 = ~(n482 | n439);
  assign n__333 = ~(n483 | n439);
  assign n__332 = ~(n484 | n439);
  assign n__331 = ~(n485 | n439);
  assign n__330 = ~(n486 | n439);
  assign n__329 = ~(n487 | n439);
  assign n__328 = ~(n488 | n439);
  assign n__327 = ~(n489 | n439);
  assign n__326 = ~(n490 | n439);
  assign n__325 = ~(n491 | n439);
  assign n__324 = ~(n492 | n439);
  assign n__323 = ~(n493 | n438);
  assign n__322 = ~(n494 | n438);
  assign n__321 = ~(n495 | n438);
  assign n__320 = ~(n496 | n438);
  assign n__319 = ~(n497 | n438);
  assign n__318 = ~(n498 | n438);
  assign n__317 = ~(n499 | n438);
  assign n__316 = ~(n500 | n438);
  assign n__315 = ~(n501 | n438);
  assign n__314 = ~(n502 | n438);
  assign n__313 = ~(n503 | n438);
  assign n__312 = ~(n504 | n438);
  assign n__311 = ~(n505 | n438);
  assign n__310 = ~(n506 | n437);
  assign n__309 = ~(n507 | n437);
  assign n__308 = ~(n508 | n437);
  assign n__307 = ~(n509 | n437);
  assign n__306 = ~(n510 | n437);
  assign n__305 = ~(n511 | n437);
  assign n__304 = ~(n512 | n437);
  assign n__303 = ~(n513 | n437);
  assign n__302 = ~(n514 | n437);
  assign n__301 = ~(n515 | n437);
  assign n__300 = ~(n516 | n437);
  assign n__2 = ~n570;
  assign n__299 = ~(n517 | n437);
  assign n__298 = ~(n518 | n437);
  assign n__297 = ~(n519 | n436);
  assign n__296 = ~(n520 | n436);
  assign n__295 = ~(n521 | n436);
  assign n__294 = ~(n522 | n436);
  assign n__293 = ~(n523 | n436);
  assign n__292 = ~(n524 | n436);
  assign n__291 = ~(n525 | n436);
  assign n__290 = ~(n526 | n436);
  assign n__289 = ~(n527 | n436);
  assign n__288 = ~(n528 | n436);
  assign n__287 = ~(n529 | n436);
  assign n__286 = ~(n530 | n436);
  assign n__285 = ~(n531 | n436);
  assign n__284 = ~(n532 | n435);
  assign n__283 = ~(n533 | n435);
  assign n__282 = ~(n534 | n435);
  assign n__281 = ~(n535 | n435);
  assign n__280 = ~(n536 | n435);
  assign n__279 = ~(n537 | n435);
  assign n__278 = ~(n538 | n435);
  assign n__277 = ~(n539 | n435);
  assign n__276 = ~(n540 | n435);
  assign n__275 = ~(n541 | n435);
  assign n__274 = ~(n542 | n435);
  assign n__273 = ~(n543 | n435);
  assign n__272 = ~(n544 | n435);
  assign n__271 = ~(n545 | n434);
  assign n__270 = ~(n546 | n434);
  assign n__269 = ~(n547 | n434);
  assign n__268 = ~(n548 | n434);
  assign n__267 = ~(n549 | n434);
  assign n__266 = ~(n550 | n434);
  assign n__265 = ~(n551 | n434);
  assign n__264 = ~(n552 | n434);
  assign n__263 = ~(n553 | n434);
  assign n__262 = ~(n554 | n434);
  assign n__261 = ~(n555 | n434);
  assign n__260 = ~(n556 | n434);
  assign n__259 = ~(n557 | n434);
  assign n__258 = ~(n558 | n433);
  assign n__257 = ~(n559 | n433);
  assign n__256 = ~(n560 | n433);
  assign n__255 = ~(n561 | n433);
  assign n__254 = ~(n562 | n433);
  assign n__253 = ~(n563 | n433);
  assign n__252 = ~(n564 | n433);
  assign n__251 = ~(n565 | n433);
  assign n__250 = ~(n566 | n433);
  assign n__24 = ~n571;
  assign n__249 = ~(n567 | n433);
  assign n__248 = ~(n568 | n433);
  assign n__247 = ~(n569 | n433);
  assign n__246 = ~(n423 | n433);
  assign n__245 = ~n443;
  assign n443 = ~(b__5 & n__118);
  assign n__244 = ~n444;
  assign n444 = ~(n__117 & b__5);
  assign n__243 = ~n445;
  assign n445 = ~(n__116 & b__5);
  assign n__242 = ~n446;
  assign n446 = ~(n__115 & b__5);
  assign n__241 = ~n447;
  assign n447 = ~(n__114 & b__5);
  assign n__240 = ~n448;
  assign n448 = ~(n__113 & b__5);
  assign n__23 = ~n572;
  assign n__239 = ~n449;
  assign n449 = ~(n__112 & b__5);
  assign n__238 = ~n450;
  assign n450 = ~(n__111 & b__5);
  assign n__237 = ~n451;
  assign n451 = ~(n__110 & b__5);
  assign n__236 = ~n452;
  assign n452 = ~(n__109 & b__5);
  assign n__235 = ~n453;
  assign n453 = ~(n__108 & b__5);
  assign n__234 = ~n454;
  assign n454 = ~(n__107 & b__5);
  assign n__233 = ~n455;
  assign n455 = ~(n__106 & b__5);
  assign n__232 = ~n456;
  assign n456 = ~(n__105 & b__5);
  assign n__231 = ~n457;
  assign n457 = ~(n__104 & b__5);
  assign n__230 = ~n458;
  assign n458 = ~(n__103 & b__5);
  assign n__22 = ~n573;
  assign n__229 = ~n459;
  assign n459 = ~(n__102 & b__5);
  assign n__228 = ~n460;
  assign n460 = ~(n__101 & b__5);
  assign n__227 = ~n461;
  assign n461 = ~(n__100 & b__5);
  assign n__226 = ~n462;
  assign n462 = ~(n__99 & b__5);
  assign n__225 = ~n463;
  assign n463 = ~(n__98 & b__5);
  assign n__224 = ~n464;
  assign n464 = ~(n__97 & b__5);
  assign n__223 = ~n465;
  assign n465 = ~(n__96 & b__5);
  assign n__222 = ~n466;
  assign n466 = ~(n__95 & b__5);
  assign n__221 = ~n467;
  assign n467 = ~(n__94 & b__5);
  assign n__220 = ~n468;
  assign n468 = ~(n__93 & b__5);
  assign n__21 = ~n574;
  assign n__219 = ~n469;
  assign n469 = ~(n__92 & b__5);
  assign n__218 = ~n470;
  assign n470 = ~(n__91 & b__5);
  assign n__217 = ~n471;
  assign n471 = ~(n__90 & b__5);
  assign n__216 = ~n472;
  assign n472 = ~(n__89 & b__5);
  assign n__215 = ~n473;
  assign n473 = ~(n__88 & b__5);
  assign n__214 = ~n474;
  assign n474 = ~(n__87 & b__5);
  assign n__213 = ~n475;
  assign n475 = ~(n__86 & b__5);
  assign n__212 = ~n476;
  assign n476 = ~(n__85 & b__5);
  assign n__211 = ~n477;
  assign n477 = ~(n__84 & b__5);
  assign n__210 = ~n478;
  assign n478 = ~(n__83 & b__5);
  assign n__20 = ~n575;
  assign n__209 = ~n479;
  assign n479 = ~(n__82 & b__5);
  assign n__208 = ~n480;
  assign n480 = ~(n__81 & b__5);
  assign n__207 = ~n481;
  assign n481 = ~(n__80 & b__5);
  assign n__206 = ~n482;
  assign n482 = ~(n__79 & b__5);
  assign n__205 = ~n483;
  assign n483 = ~(n__78 & b__5);
  assign n__204 = ~n484;
  assign n484 = ~(n__77 & b__5);
  assign n__203 = ~n485;
  assign n485 = ~(n__76 & b__5);
  assign n__202 = ~n486;
  assign n486 = ~(n__75 & b__5);
  assign n__201 = ~n487;
  assign n487 = ~(n__74 & b__5);
  assign n__200 = ~n488;
  assign n488 = ~(n__73 & b__5);
  assign n__1 = ~n576;
  assign n__19 = ~n577;
  assign n__199 = ~n489;
  assign n489 = ~(n__72 & b__5);
  assign n__198 = ~n490;
  assign n490 = ~(n__71 & b__5);
  assign n__197 = ~n491;
  assign n491 = ~(n__70 & b__5);
  assign n__196 = ~n492;
  assign n492 = ~(n__69 & b__5);
  assign n__195 = ~n493;
  assign n493 = ~(n__68 & b__5);
  assign n__194 = ~n494;
  assign n494 = ~(n__67 & b__5);
  assign n__193 = ~n495;
  assign n495 = ~(n__66 & b__5);
  assign n__192 = ~n496;
  assign n496 = ~(n__65 & b__5);
  assign n__191 = ~n497;
  assign n497 = ~(n__64 & b__5);
  assign n__190 = ~n498;
  assign n498 = ~(n__63 & b__5);
  assign n__18 = ~n578;
  assign n__189 = ~n499;
  assign n499 = ~(n__62 & b__5);
  assign n__188 = ~n500;
  assign n500 = ~(n__61 & b__5);
  assign n__187 = ~n501;
  assign n501 = ~(n__60 & b__5);
  assign n__186 = ~n502;
  assign n502 = ~(n__59 & b__5);
  assign n__185 = ~n503;
  assign n503 = ~(n__58 & b__5);
  assign n__184 = ~n504;
  assign n504 = ~(n__57 & b__5);
  assign n__183 = ~n505;
  assign n505 = ~(n__56 & b__5);
  assign n__182 = ~n506;
  assign n506 = ~(a__5 & n__118);
  assign n__181 = ~n507;
  assign n507 = ~(a__5 & n__117);
  assign n__180 = ~n508;
  assign n508 = ~(a__5 & n__116);
  assign n__17 = ~n579;
  assign n__179 = ~n509;
  assign n509 = ~(a__5 & n__115);
  assign n__178 = ~n510;
  assign n510 = ~(a__5 & n__114);
  assign n__177 = ~n511;
  assign n511 = ~(a__5 & n__113);
  assign n__176 = ~n512;
  assign n512 = ~(a__5 & n__112);
  assign n__175 = ~n513;
  assign n513 = ~(a__5 & n__111);
  assign n__174 = ~n514;
  assign n514 = ~(a__5 & n__110);
  assign n__173 = ~n515;
  assign n515 = ~(a__5 & n__109);
  assign n__172 = ~n516;
  assign n516 = ~(a__5 & n__108);
  assign n__171 = ~n517;
  assign n517 = ~(a__5 & n__107);
  assign n__170 = ~n518;
  assign n518 = ~(a__5 & n__106);
  assign n__16 = ~n580;
  assign n__169 = ~n519;
  assign n519 = ~(a__5 & n__105);
  assign n__168 = ~n520;
  assign n520 = ~(a__5 & n__104);
  assign n__167 = ~n521;
  assign n521 = ~(a__5 & n__103);
  assign n__166 = ~n522;
  assign n522 = ~(a__5 & n__102);
  assign n__165 = ~n523;
  assign n523 = ~(a__5 & n__101);
  assign n__164 = ~n524;
  assign n524 = ~(a__5 & n__100);
  assign n__163 = ~n525;
  assign n525 = ~(a__5 & n__99);
  assign n__99 = ~n581;
  assign n581 = ~(b__4 & n__36);
  assign n__162 = ~n526;
  assign n526 = ~(a__5 & n__98);
  assign n__98 = ~n582;
  assign n582 = ~(n__35 & b__4);
  assign n__161 = ~n527;
  assign n527 = ~(a__5 & n__97);
  assign n__97 = ~n583;
  assign n583 = ~(n__34 & b__4);
  assign n__160 = ~n528;
  assign n528 = ~(a__5 & n__96);
  assign n__96 = ~n584;
  assign n584 = ~(n__33 & b__4);
  assign n__15 = ~n585;
  assign n__159 = ~n529;
  assign n529 = ~(a__5 & n__95);
  assign n__95 = ~n586;
  assign n586 = ~(n__32 & b__4);
  assign n__158 = ~n530;
  assign n530 = ~(a__5 & n__94);
  assign n__94 = ~n587;
  assign n587 = ~(n__31 & b__4);
  assign n__157 = ~n531;
  assign n531 = ~(a__5 & n__93);
  assign n__93 = ~n588;
  assign n588 = ~(n__30 & b__4);
  assign n__156 = ~n532;
  assign n532 = ~(a__5 & n__92);
  assign n__92 = ~n589;
  assign n589 = ~(n__29 & b__4);
  assign n__155 = ~n533;
  assign n533 = ~(a__5 & n__91);
  assign n__91 = ~n590;
  assign n590 = ~(n__28 & b__4);
  assign n__154 = ~n534;
  assign n534 = ~(a__5 & n__90);
  assign n__90 = ~n591;
  assign n591 = ~(n__27 & b__4);
  assign n__153 = ~n535;
  assign n535 = ~(a__5 & n__89);
  assign n__89 = ~n592;
  assign n592 = ~(n__26 & b__4);
  assign n__152 = ~n536;
  assign n536 = ~(a__5 & n__88);
  assign n__88 = ~n593;
  assign n593 = ~(n__25 & b__4);
  assign n__151 = ~n537;
  assign n537 = ~(a__5 & n__87);
  assign n__87 = ~n594;
  assign n594 = ~(a__4 & n__55);
  assign n__150 = ~n538;
  assign n538 = ~(a__5 & n__86);
  assign n__86 = ~n595;
  assign n595 = ~(n__54 & a__4);
  assign n__14 = ~n596;
  assign n__149 = ~n539;
  assign n539 = ~(a__5 & n__85);
  assign n__85 = ~n597;
  assign n597 = ~(n__53 & a__4);
  assign n__148 = ~n540;
  assign n540 = ~(a__5 & n__84);
  assign n__84 = ~n598;
  assign n598 = ~(n__52 & a__4);
  assign n__147 = ~n541;
  assign n541 = ~(a__5 & n__83);
  assign n__83 = ~n599;
  assign n599 = ~(n__51 & a__4);
  assign n__146 = ~n542;
  assign n542 = ~(a__5 & n__82);
  assign n__82 = ~n600;
  assign n600 = ~(n__50 & a__4);
  assign n__145 = ~n543;
  assign n543 = ~(a__5 & n__81);
  assign n__81 = ~n601;
  assign n601 = ~(n__49 & a__4);
  assign n__144 = ~n544;
  assign n544 = ~(a__5 & n__80);
  assign n__80 = ~n602;
  assign n602 = ~(n__48 & a__4);
  assign n__143 = ~n545;
  assign n545 = ~(a__5 & n__79);
  assign n__79 = ~n603;
  assign n603 = ~(n__47 & a__4);
  assign n__142 = ~n546;
  assign n546 = ~(a__5 & n__78);
  assign n__78 = ~n604;
  assign n604 = ~(n__46 & a__4);
  assign n__141 = ~n547;
  assign n547 = ~(a__5 & n__77);
  assign n__77 = ~n605;
  assign n605 = ~(n__45 & a__4);
  assign n__140 = ~n548;
  assign n548 = ~(a__5 & n__76);
  assign n__76 = ~n606;
  assign n606 = ~(n__44 & a__4);
  assign n__13 = ~n607;
  assign n__139 = ~n549;
  assign n549 = ~(a__5 & n__75);
  assign n__75 = ~n608;
  assign n608 = ~(n__43 & a__4);
  assign n__138 = ~n550;
  assign n550 = ~(a__5 & n__74);
  assign n__74 = ~n609;
  assign n609 = ~(n__42 & a__4);
  assign n__137 = ~n551;
  assign n551 = ~(a__5 & n__73);
  assign n__73 = ~n610;
  assign n610 = ~(n__41 & a__4);
  assign n__136 = ~n552;
  assign n552 = ~(a__5 & n__72);
  assign n__72 = ~n611;
  assign n611 = ~(n__40 & a__4);
  assign n__135 = ~n553;
  assign n553 = ~(a__5 & n__71);
  assign n__71 = ~n612;
  assign n612 = ~(n__39 & a__4);
  assign n__134 = ~n554;
  assign n554 = ~(a__5 & n__70);
  assign n__70 = ~n613;
  assign n613 = ~(n__38 & a__4);
  assign n__133 = ~n555;
  assign n555 = ~(a__5 & n__69);
  assign n__69 = ~n614;
  assign n614 = ~(n__37 & a__4);
  assign n__132 = ~n556;
  assign n556 = ~(a__5 & n__68);
  assign n__68 = ~n615;
  assign n615 = ~(a__4 & n__36);
  assign n__36 = ~(n616 | n575);
  assign n__131 = ~n557;
  assign n557 = ~(a__5 & n__67);
  assign n__67 = ~n617;
  assign n617 = ~(a__4 & n__35);
  assign n__35 = ~(n577 | n616);
  assign n__130 = ~n558;
  assign n558 = ~(a__5 & n__66);
  assign n__66 = ~n618;
  assign n618 = ~(a__4 & n__34);
  assign n__34 = ~(n578 | n616);
  assign n__12 = ~n619;
  assign n__129 = ~n559;
  assign n559 = ~(a__5 & n__65);
  assign n__65 = ~n620;
  assign n620 = ~(a__4 & n__33);
  assign n__33 = ~(n579 | n616);
  assign n__128 = ~n560;
  assign n560 = ~(a__5 & n__64);
  assign n__64 = ~n621;
  assign n621 = ~(a__4 & n__32);
  assign n__32 = ~(n580 | n616);
  assign n__127 = ~n561;
  assign n561 = ~(a__5 & n__63);
  assign n__63 = ~n622;
  assign n622 = ~(a__4 & n__31);
  assign n__31 = ~(n585 | n616);
  assign n__126 = ~n562;
  assign n562 = ~(a__5 & n__62);
  assign n__62 = ~n623;
  assign n623 = ~(a__4 & n__30);
  assign n__30 = ~(n596 | n616);
  assign n__125 = ~n563;
  assign n563 = ~(a__5 & n__61);
  assign n__61 = ~n624;
  assign n624 = ~(a__4 & n__29);
  assign n__29 = ~(n607 | n616);
  assign n__124 = ~n564;
  assign n564 = ~(a__5 & n__60);
  assign n__60 = ~n625;
  assign n625 = ~(a__4 & n__28);
  assign n__28 = ~(n619 | n616);
  assign n__123 = ~n565;
  assign n565 = ~(a__5 & n__59);
  assign n__59 = ~n626;
  assign n626 = ~(a__4 & n__27);
  assign n__27 = ~(n627 | n616);
  assign n__122 = ~n566;
  assign n566 = ~(a__5 & n__58);
  assign n__58 = ~n628;
  assign n628 = ~(a__4 & n__26);
  assign n__26 = ~(n629 | n616);
  assign n__121 = ~n567;
  assign n567 = ~(a__5 & n__57);
  assign n__57 = ~n630;
  assign n630 = ~(a__4 & n__25);
  assign n__25 = ~(n631 | n616);
  assign n__120 = ~n568;
  assign n568 = ~(a__5 & n__56);
  assign n__56 = ~n632;
  assign n632 = ~(a__4 & b__4);
  assign n__11 = ~n627;
  assign n__119 = ~n569;
  assign n569 = ~(a__5 & b__5);
  assign n__118 = ~n633;
  assign n633 = ~(n__55 & b__4);
  assign n__55 = ~(n571 | n631);
  assign n__117 = ~n634;
  assign n634 = ~(n__54 & b__4);
  assign n__54 = ~(n572 | n631);
  assign n__116 = ~n635;
  assign n635 = ~(n__53 & b__4);
  assign n__53 = ~(n573 | n631);
  assign n__115 = ~n636;
  assign n636 = ~(n__52 & b__4);
  assign n__52 = ~(n574 | n631);
  assign n__114 = ~n637;
  assign n637 = ~(n__51 & b__4);
  assign n__51 = ~(n631 | n575);
  assign n575 = ~(b__2 & n__5);
  assign n__113 = ~n638;
  assign n638 = ~(n__50 & b__4);
  assign n__50 = ~(n631 | n577);
  assign n577 = ~(n__4 & b__2);
  assign n__112 = ~n639;
  assign n639 = ~(n__49 & b__4);
  assign n__49 = ~(n631 | n578);
  assign n578 = ~(n__3 & b__2);
  assign n__111 = ~n640;
  assign n640 = ~(n__48 & b__4);
  assign n__48 = ~(n631 | n579);
  assign n579 = ~(a__2 & n__9);
  assign n__110 = ~n641;
  assign n641 = ~(n__47 & b__4);
  assign n__47 = ~(n631 | n580);
  assign n580 = ~(n__8 & a__2);
  assign n__10 = ~n629;
  assign n__109 = ~n642;
  assign n642 = ~(n__46 & b__4);
  assign n__46 = ~(n631 | n585);
  assign n585 = ~(n__7 & a__2);
  assign n__108 = ~n643;
  assign n643 = ~(n__45 & b__4);
  assign n__45 = ~(n631 | n596);
  assign n596 = ~(n__6 & a__2);
  assign n__107 = ~n644;
  assign n644 = ~(n__44 & b__4);
  assign n__44 = ~(n631 | n607);
  assign n607 = ~(a__2 & n__5);
  assign n__5 = ~(n645 | n576);
  assign n__106 = ~n646;
  assign n646 = ~(n__43 & b__4);
  assign n__43 = ~(n631 | n619);
  assign n619 = ~(a__2 & n__4);
  assign n__4 = ~(n647 | n645);
  assign n__105 = ~n648;
  assign n648 = ~(n__42 & b__4);
  assign n__42 = ~(n631 | n627);
  assign n627 = ~(a__2 & n__3);
  assign n__3 = ~(n645 | n649);
  assign n__104 = ~n650;
  assign n650 = ~(n__41 & b__4);
  assign n__41 = ~(n631 | n629);
  assign n629 = ~(a__2 & b__2);
  assign n631 = ~b__3;
  assign n__103 = ~n651;
  assign n651 = ~(n__40 & b__4);
  assign n__40 = ~(n571 | n616);
  assign n571 = ~(n__9 & b__2);
  assign n__9 = ~(n649 | n570);
  assign n__102 = ~n652;
  assign n652 = ~(n__39 & b__4);
  assign n__39 = ~(n572 | n616);
  assign n572 = ~(n__8 & b__2);
  assign n__8 = ~(n576 | n649);
  assign n576 = ~(a__0 & c);
  assign n__101 = ~n653;
  assign n653 = ~(n__38 & b__4);
  assign n__38 = ~(n573 | n616);
  assign n573 = ~(n__7 & b__2);
  assign n__7 = ~(n647 | n649);
  assign n649 = ~b__1;
  assign n__100 = ~n654;
  assign n654 = ~(n__37 & b__4);
  assign n__37 = ~(n574 | n616);
  assign n616 = ~a__3;
  assign n574 = ~(n__6 & b__2);
  assign n__6 = ~(n645 | n570);
  assign n570 = ~(c & b__0);
  assign n645 = ~a__1;
  assign n__0 = ~n647;
  assign n647 = ~(a__0 & b__0);
endmodule