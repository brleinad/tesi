
module generator ( i, c );
  input [6:0] i;
  output [14:0] c;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13;
  assign c[6] = i[6];
  assign c[5] = i[5];
  assign c[4] = i[4];
  assign c[3] = i[3];
  assign c[2] = i[2];
  assign c[1] = i[1];
  assign c[0] = i[0];

  GTECH_XOR2 __tmp100_1 ( .A(c[0]), .B(c[1]), .Z(N0) );
  GTECH_XOR2 __tmp100_2 ( .A(N0), .B(c[3]), .Z(c[7]) );
  GTECH_XOR2 __tmp101_1 ( .A(c[1]), .B(c[2]), .Z(N1) );
  GTECH_XOR2 __tmp101_2 ( .A(N1), .B(c[4]), .Z(c[8]) );
  GTECH_XOR2 __tmp102_1 ( .A(c[2]), .B(c[3]), .Z(N2) );
  GTECH_XOR2 __tmp102_2 ( .A(N2), .B(c[5]), .Z(c[9]) );
  GTECH_XOR2 __tmp103_1 ( .A(c[3]), .B(c[4]), .Z(N3) );
  GTECH_XOR2 __tmp103_2 ( .A(N3), .B(c[6]), .Z(c[10]) );
  GTECH_XOR2 __tmp104_1 ( .A(c[0]), .B(c[1]), .Z(N4) );
  GTECH_XOR2 __tmp104_2 ( .A(N4), .B(c[3]), .Z(N5) );
  GTECH_XOR2 __tmp104_3 ( .A(N5), .B(c[4]), .Z(N6) );
  GTECH_XOR2 __tmp104_4 ( .A(N6), .B(c[5]), .Z(c[11]) );
  GTECH_XOR2 __tmp105_1 ( .A(c[1]), .B(c[2]), .Z(N7) );
  GTECH_XOR2 __tmp105_2 ( .A(N7), .B(c[4]), .Z(N8) );
  GTECH_XOR2 __tmp105_3 ( .A(N8), .B(c[5]), .Z(N9) );
  GTECH_XOR2 __tmp105_4 ( .A(N9), .B(c[6]), .Z(c[12]) );
  GTECH_XOR2 __tmp106_1 ( .A(c[0]), .B(c[1]), .Z(N10) );
  GTECH_XOR2 __tmp106_2 ( .A(N10), .B(c[2]), .Z(N11) );
  GTECH_XOR2 __tmp106_3 ( .A(N11), .B(c[5]), .Z(N12) );
  GTECH_XOR2 __tmp106_4 ( .A(N12), .B(c[6]), .Z(c[13]) );
  GTECH_XOR2 __tmp107_1 ( .A(c[0]), .B(c[2]), .Z(N13) );
  GTECH_XOR2 __tmp107_2 ( .A(N13), .B(c[6]), .Z(c[14]) );
endmodule


module gen_linear_part ( a, b, c_in, n, s );
  input [6:0] a;
  input [6:0] b;
  input [500:0] n;
  output [7:0] s;
  input c_in;
  wire   t_245, t_244, t_243, t_242, t_241, t_240, t_239, t_238, t_237, t_236,
         t_235, t_234, t_233, t_232, t_231, t_230, t_229, t_228, t_227, t_226,
         t_225, t_224, t_223, t_222, t_221, t_220, t_219, t_218, t_217, t_216,
         t_215, t_214, t_213, t_212, t_211, t_210, t_209, t_208, t_207, t_206,
         t_205, t_204, t_203, t_202, t_201, t_200, t_199, t_198, t_197, t_196,
         t_195, t_194, t_193, t_192, t_191, t_190, t_189, t_188, t_187, t_186,
         t_185, t_184, t_183, t_182, t_181, t_180, t_179, t_178, t_177, t_176,
         t_175, t_174, t_173, t_172, t_171, t_170, t_169, t_168, t_167, t_166,
         t_165, t_164, t_163, t_162, t_161, t_160, t_159, t_158, t_157, t_156,
         t_155, t_154, t_153, t_152, t_151, t_150, t_149, t_148, t_147, t_146,
         t_145, t_144, t_143, t_142, t_141, t_140, t_139, t_138, t_137, t_136,
         t_135, t_134, t_133, t_132, t_131, t_130, t_129, t_128, t_127, t_126,
         t_125, t_124, t_123, t_122, t_121, t_120, t_118, t_117, t_116, t_115,
         t_114, t_113, t_112, t_111, t_110, t_109, t_108, t_107, t_106, t_105,
         t_104, t_103, t_102, t_101, t_100, t_99, t_98, t_97, t_96, t_95, t_94,
         t_93, t_92, t_91, t_90, t_89, t_88, t_87, t_86, t_85, t_84, t_83,
         t_82, t_81, t_80, t_79, t_78, t_77, t_76, t_75, t_74, t_73, t_72,
         t_71, t_70, t_69, t_68, t_67, t_66, t_65, t_64, t_63, t_62, t_61,
         t_60, t_59, t_58, t_57, t_55, t_54, t_53, t_52, t_51, t_50, t_49,
         t_48, t_47, t_46, t_45, t_44, t_43, t_42, t_41, t_40, t_39, t_38,
         t_37, t_36, t_35, t_34, t_33, t_32, t_31, t_30, t_29, t_28, t_27,
         t_26, t_24, t_23, t_22, t_21, t_20, t_19, t_18, t_17, t_16, t_15,
         t_14, t_13, t_12, t_11, t_9, t_8, t_7, t_6, t_5, t_4, t_2, t_1, N0,
         N1, N2, N3, N4, N5, N6;
  wire   [499:247] t;

  GTECH_XOR2 C507 ( .A(N0), .B(c_in), .Z(s[0]) );
  GTECH_XOR2 C508 ( .A(a[0]), .B(b[0]), .Z(N0) );
  GTECH_XOR2 C509 ( .A(n[0]), .B(n[1]), .Z(t_1) );
  GTECH_XOR2 C510 ( .A(t_1), .B(n[2]), .Z(t_2) );
  GTECH_XOR2 C511 ( .A(N1), .B(t_2), .Z(s[1]) );
  GTECH_XOR2 C512 ( .A(a[1]), .B(b[1]), .Z(N1) );
  GTECH_XOR2 C513 ( .A(n[3]), .B(n[4]), .Z(t_4) );
  GTECH_XOR2 C514 ( .A(t_4), .B(n[5]), .Z(t_5) );
  GTECH_XOR2 C515 ( .A(t_5), .B(n[6]), .Z(t_6) );
  GTECH_XOR2 C516 ( .A(t_6), .B(n[7]), .Z(t_7) );
  GTECH_XOR2 C517 ( .A(t_7), .B(n[8]), .Z(t_8) );
  GTECH_XOR2 C518 ( .A(t_8), .B(n[9]), .Z(t_9) );
  GTECH_XOR2 C519 ( .A(N2), .B(t_9), .Z(s[2]) );
  GTECH_XOR2 C520 ( .A(a[2]), .B(b[2]), .Z(N2) );
  GTECH_XOR2 C521 ( .A(n[10]), .B(n[11]), .Z(t_11) );
  GTECH_XOR2 C522 ( .A(t_11), .B(n[12]), .Z(t_12) );
  GTECH_XOR2 C523 ( .A(t_12), .B(n[13]), .Z(t_13) );
  GTECH_XOR2 C524 ( .A(t_13), .B(n[14]), .Z(t_14) );
  GTECH_XOR2 C525 ( .A(t_14), .B(n[15]), .Z(t_15) );
  GTECH_XOR2 C526 ( .A(t_15), .B(n[16]), .Z(t_16) );
  GTECH_XOR2 C527 ( .A(t_16), .B(n[17]), .Z(t_17) );
  GTECH_XOR2 C528 ( .A(t_17), .B(n[18]), .Z(t_18) );
  GTECH_XOR2 C529 ( .A(t_18), .B(n[19]), .Z(t_19) );
  GTECH_XOR2 C530 ( .A(t_19), .B(n[20]), .Z(t_20) );
  GTECH_XOR2 C531 ( .A(t_20), .B(n[21]), .Z(t_21) );
  GTECH_XOR2 C532 ( .A(t_21), .B(n[22]), .Z(t_22) );
  GTECH_XOR2 C533 ( .A(t_22), .B(n[23]), .Z(t_23) );
  GTECH_XOR2 C534 ( .A(t_23), .B(n[24]), .Z(t_24) );
  GTECH_XOR2 C535 ( .A(N3), .B(t_24), .Z(s[3]) );
  GTECH_XOR2 C536 ( .A(a[3]), .B(b[3]), .Z(N3) );
  GTECH_XOR2 C537 ( .A(n[25]), .B(n[26]), .Z(t_26) );
  GTECH_XOR2 C538 ( .A(t_26), .B(n[27]), .Z(t_27) );
  GTECH_XOR2 C539 ( .A(t_27), .B(n[28]), .Z(t_28) );
  GTECH_XOR2 C540 ( .A(t_28), .B(n[29]), .Z(t_29) );
  GTECH_XOR2 C541 ( .A(t_29), .B(n[30]), .Z(t_30) );
  GTECH_XOR2 C542 ( .A(t_30), .B(n[31]), .Z(t_31) );
  GTECH_XOR2 C543 ( .A(t_31), .B(n[32]), .Z(t_32) );
  GTECH_XOR2 C544 ( .A(t_32), .B(n[33]), .Z(t_33) );
  GTECH_XOR2 C545 ( .A(t_33), .B(n[34]), .Z(t_34) );
  GTECH_XOR2 C546 ( .A(t_34), .B(n[35]), .Z(t_35) );
  GTECH_XOR2 C547 ( .A(t_35), .B(n[36]), .Z(t_36) );
  GTECH_XOR2 C548 ( .A(t_36), .B(n[37]), .Z(t_37) );
  GTECH_XOR2 C549 ( .A(t_37), .B(n[38]), .Z(t_38) );
  GTECH_XOR2 C550 ( .A(t_38), .B(n[39]), .Z(t_39) );
  GTECH_XOR2 C551 ( .A(t_39), .B(n[40]), .Z(t_40) );
  GTECH_XOR2 C552 ( .A(t_40), .B(n[41]), .Z(t_41) );
  GTECH_XOR2 C553 ( .A(t_41), .B(n[42]), .Z(t_42) );
  GTECH_XOR2 C554 ( .A(t_42), .B(n[43]), .Z(t_43) );
  GTECH_XOR2 C555 ( .A(t_43), .B(n[44]), .Z(t_44) );
  GTECH_XOR2 C556 ( .A(t_44), .B(n[45]), .Z(t_45) );
  GTECH_XOR2 C557 ( .A(t_45), .B(n[46]), .Z(t_46) );
  GTECH_XOR2 C558 ( .A(t_46), .B(n[47]), .Z(t_47) );
  GTECH_XOR2 C559 ( .A(t_47), .B(n[48]), .Z(t_48) );
  GTECH_XOR2 C560 ( .A(t_48), .B(n[49]), .Z(t_49) );
  GTECH_XOR2 C561 ( .A(t_49), .B(n[50]), .Z(t_50) );
  GTECH_XOR2 C562 ( .A(t_50), .B(n[51]), .Z(t_51) );
  GTECH_XOR2 C563 ( .A(t_51), .B(n[52]), .Z(t_52) );
  GTECH_XOR2 C564 ( .A(t_52), .B(n[53]), .Z(t_53) );
  GTECH_XOR2 C565 ( .A(t_53), .B(n[54]), .Z(t_54) );
  GTECH_XOR2 C566 ( .A(t_54), .B(n[55]), .Z(t_55) );
  GTECH_XOR2 C567 ( .A(N4), .B(t_55), .Z(s[4]) );
  GTECH_XOR2 C568 ( .A(a[4]), .B(b[4]), .Z(N4) );
  GTECH_XOR2 C569 ( .A(n[56]), .B(n[57]), .Z(t_57) );
  GTECH_XOR2 C570 ( .A(t_57), .B(n[58]), .Z(t_58) );
  GTECH_XOR2 C571 ( .A(t_58), .B(n[59]), .Z(t_59) );
  GTECH_XOR2 C572 ( .A(t_59), .B(n[60]), .Z(t_60) );
  GTECH_XOR2 C573 ( .A(t_60), .B(n[61]), .Z(t_61) );
  GTECH_XOR2 C574 ( .A(t_61), .B(n[62]), .Z(t_62) );
  GTECH_XOR2 C575 ( .A(t_62), .B(n[63]), .Z(t_63) );
  GTECH_XOR2 C576 ( .A(t_63), .B(n[64]), .Z(t_64) );
  GTECH_XOR2 C577 ( .A(t_64), .B(n[65]), .Z(t_65) );
  GTECH_XOR2 C578 ( .A(t_65), .B(n[66]), .Z(t_66) );
  GTECH_XOR2 C579 ( .A(t_66), .B(n[67]), .Z(t_67) );
  GTECH_XOR2 C580 ( .A(t_67), .B(n[68]), .Z(t_68) );
  GTECH_XOR2 C581 ( .A(t_68), .B(n[69]), .Z(t_69) );
  GTECH_XOR2 C582 ( .A(t_69), .B(n[70]), .Z(t_70) );
  GTECH_XOR2 C583 ( .A(t_70), .B(n[71]), .Z(t_71) );
  GTECH_XOR2 C584 ( .A(t_71), .B(n[72]), .Z(t_72) );
  GTECH_XOR2 C585 ( .A(t_72), .B(n[73]), .Z(t_73) );
  GTECH_XOR2 C586 ( .A(t_73), .B(n[74]), .Z(t_74) );
  GTECH_XOR2 C587 ( .A(t_74), .B(n[75]), .Z(t_75) );
  GTECH_XOR2 C588 ( .A(t_75), .B(n[76]), .Z(t_76) );
  GTECH_XOR2 C589 ( .A(t_76), .B(n[77]), .Z(t_77) );
  GTECH_XOR2 C590 ( .A(t_77), .B(n[78]), .Z(t_78) );
  GTECH_XOR2 C591 ( .A(t_78), .B(n[79]), .Z(t_79) );
  GTECH_XOR2 C592 ( .A(t_79), .B(n[80]), .Z(t_80) );
  GTECH_XOR2 C593 ( .A(t_80), .B(n[81]), .Z(t_81) );
  GTECH_XOR2 C594 ( .A(t_81), .B(n[82]), .Z(t_82) );
  GTECH_XOR2 C595 ( .A(t_82), .B(n[83]), .Z(t_83) );
  GTECH_XOR2 C596 ( .A(t_83), .B(n[84]), .Z(t_84) );
  GTECH_XOR2 C597 ( .A(t_84), .B(n[85]), .Z(t_85) );
  GTECH_XOR2 C598 ( .A(t_85), .B(n[86]), .Z(t_86) );
  GTECH_XOR2 C599 ( .A(t_86), .B(n[87]), .Z(t_87) );
  GTECH_XOR2 C600 ( .A(t_87), .B(n[88]), .Z(t_88) );
  GTECH_XOR2 C601 ( .A(t_88), .B(n[89]), .Z(t_89) );
  GTECH_XOR2 C602 ( .A(t_89), .B(n[90]), .Z(t_90) );
  GTECH_XOR2 C603 ( .A(t_90), .B(n[91]), .Z(t_91) );
  GTECH_XOR2 C604 ( .A(t_91), .B(n[92]), .Z(t_92) );
  GTECH_XOR2 C605 ( .A(t_92), .B(n[93]), .Z(t_93) );
  GTECH_XOR2 C606 ( .A(t_93), .B(n[94]), .Z(t_94) );
  GTECH_XOR2 C607 ( .A(t_94), .B(n[95]), .Z(t_95) );
  GTECH_XOR2 C608 ( .A(t_95), .B(n[96]), .Z(t_96) );
  GTECH_XOR2 C609 ( .A(t_96), .B(n[97]), .Z(t_97) );
  GTECH_XOR2 C610 ( .A(t_97), .B(n[98]), .Z(t_98) );
  GTECH_XOR2 C611 ( .A(t_98), .B(n[99]), .Z(t_99) );
  GTECH_XOR2 C612 ( .A(t_99), .B(n[100]), .Z(t_100) );
  GTECH_XOR2 C613 ( .A(t_100), .B(n[101]), .Z(t_101) );
  GTECH_XOR2 C614 ( .A(t_101), .B(n[102]), .Z(t_102) );
  GTECH_XOR2 C615 ( .A(t_102), .B(n[103]), .Z(t_103) );
  GTECH_XOR2 C616 ( .A(t_103), .B(n[104]), .Z(t_104) );
  GTECH_XOR2 C617 ( .A(t_104), .B(n[105]), .Z(t_105) );
  GTECH_XOR2 C618 ( .A(t_105), .B(n[106]), .Z(t_106) );
  GTECH_XOR2 C619 ( .A(t_106), .B(n[107]), .Z(t_107) );
  GTECH_XOR2 C620 ( .A(t_107), .B(n[108]), .Z(t_108) );
  GTECH_XOR2 C621 ( .A(t_108), .B(n[109]), .Z(t_109) );
  GTECH_XOR2 C622 ( .A(t_109), .B(n[110]), .Z(t_110) );
  GTECH_XOR2 C623 ( .A(t_110), .B(n[111]), .Z(t_111) );
  GTECH_XOR2 C624 ( .A(t_111), .B(n[112]), .Z(t_112) );
  GTECH_XOR2 C625 ( .A(t_112), .B(n[113]), .Z(t_113) );
  GTECH_XOR2 C626 ( .A(t_113), .B(n[114]), .Z(t_114) );
  GTECH_XOR2 C627 ( .A(t_114), .B(n[115]), .Z(t_115) );
  GTECH_XOR2 C628 ( .A(t_115), .B(n[116]), .Z(t_116) );
  GTECH_XOR2 C629 ( .A(t_116), .B(n[117]), .Z(t_117) );
  GTECH_XOR2 C630 ( .A(t_117), .B(n[118]), .Z(t_118) );
  GTECH_XOR2 C631 ( .A(N5), .B(t_118), .Z(s[5]) );
  GTECH_XOR2 C632 ( .A(a[5]), .B(b[5]), .Z(N5) );
  GTECH_XOR2 C633 ( .A(n[119]), .B(n[120]), .Z(t_120) );
  GTECH_XOR2 C634 ( .A(t_120), .B(n[121]), .Z(t_121) );
  GTECH_XOR2 C635 ( .A(t_121), .B(n[122]), .Z(t_122) );
  GTECH_XOR2 C636 ( .A(t_122), .B(n[123]), .Z(t_123) );
  GTECH_XOR2 C637 ( .A(t_123), .B(n[124]), .Z(t_124) );
  GTECH_XOR2 C638 ( .A(t_124), .B(n[125]), .Z(t_125) );
  GTECH_XOR2 C639 ( .A(t_125), .B(n[126]), .Z(t_126) );
  GTECH_XOR2 C640 ( .A(t_126), .B(n[127]), .Z(t_127) );
  GTECH_XOR2 C641 ( .A(t_127), .B(n[128]), .Z(t_128) );
  GTECH_XOR2 C642 ( .A(t_128), .B(n[129]), .Z(t_129) );
  GTECH_XOR2 C643 ( .A(t_129), .B(n[130]), .Z(t_130) );
  GTECH_XOR2 C644 ( .A(t_130), .B(n[131]), .Z(t_131) );
  GTECH_XOR2 C645 ( .A(t_131), .B(n[132]), .Z(t_132) );
  GTECH_XOR2 C646 ( .A(t_132), .B(n[133]), .Z(t_133) );
  GTECH_XOR2 C647 ( .A(t_133), .B(n[134]), .Z(t_134) );
  GTECH_XOR2 C648 ( .A(t_134), .B(n[135]), .Z(t_135) );
  GTECH_XOR2 C649 ( .A(t_135), .B(n[136]), .Z(t_136) );
  GTECH_XOR2 C650 ( .A(t_136), .B(n[137]), .Z(t_137) );
  GTECH_XOR2 C651 ( .A(t_137), .B(n[138]), .Z(t_138) );
  GTECH_XOR2 C652 ( .A(t_138), .B(n[139]), .Z(t_139) );
  GTECH_XOR2 C653 ( .A(t_139), .B(n[140]), .Z(t_140) );
  GTECH_XOR2 C654 ( .A(t_140), .B(n[141]), .Z(t_141) );
  GTECH_XOR2 C655 ( .A(t_141), .B(n[142]), .Z(t_142) );
  GTECH_XOR2 C656 ( .A(t_142), .B(n[143]), .Z(t_143) );
  GTECH_XOR2 C657 ( .A(t_143), .B(n[144]), .Z(t_144) );
  GTECH_XOR2 C658 ( .A(t_144), .B(n[145]), .Z(t_145) );
  GTECH_XOR2 C659 ( .A(t_145), .B(n[146]), .Z(t_146) );
  GTECH_XOR2 C660 ( .A(t_146), .B(n[147]), .Z(t_147) );
  GTECH_XOR2 C661 ( .A(t_147), .B(n[148]), .Z(t_148) );
  GTECH_XOR2 C662 ( .A(t_148), .B(n[149]), .Z(t_149) );
  GTECH_XOR2 C663 ( .A(t_149), .B(n[150]), .Z(t_150) );
  GTECH_XOR2 C664 ( .A(t_150), .B(n[151]), .Z(t_151) );
  GTECH_XOR2 C665 ( .A(t_151), .B(n[152]), .Z(t_152) );
  GTECH_XOR2 C666 ( .A(t_152), .B(n[153]), .Z(t_153) );
  GTECH_XOR2 C667 ( .A(t_153), .B(n[154]), .Z(t_154) );
  GTECH_XOR2 C668 ( .A(t_154), .B(n[155]), .Z(t_155) );
  GTECH_XOR2 C669 ( .A(t_155), .B(n[156]), .Z(t_156) );
  GTECH_XOR2 C670 ( .A(t_156), .B(n[157]), .Z(t_157) );
  GTECH_XOR2 C671 ( .A(t_157), .B(n[158]), .Z(t_158) );
  GTECH_XOR2 C672 ( .A(t_158), .B(n[159]), .Z(t_159) );
  GTECH_XOR2 C673 ( .A(t_159), .B(n[160]), .Z(t_160) );
  GTECH_XOR2 C674 ( .A(t_160), .B(n[161]), .Z(t_161) );
  GTECH_XOR2 C675 ( .A(t_161), .B(n[162]), .Z(t_162) );
  GTECH_XOR2 C676 ( .A(t_162), .B(n[163]), .Z(t_163) );
  GTECH_XOR2 C677 ( .A(t_163), .B(n[164]), .Z(t_164) );
  GTECH_XOR2 C678 ( .A(t_164), .B(n[165]), .Z(t_165) );
  GTECH_XOR2 C679 ( .A(t_165), .B(n[166]), .Z(t_166) );
  GTECH_XOR2 C680 ( .A(t_166), .B(n[167]), .Z(t_167) );
  GTECH_XOR2 C681 ( .A(t_167), .B(n[168]), .Z(t_168) );
  GTECH_XOR2 C682 ( .A(t_168), .B(n[169]), .Z(t_169) );
  GTECH_XOR2 C683 ( .A(t_169), .B(n[170]), .Z(t_170) );
  GTECH_XOR2 C684 ( .A(t_170), .B(n[171]), .Z(t_171) );
  GTECH_XOR2 C685 ( .A(t_171), .B(n[172]), .Z(t_172) );
  GTECH_XOR2 C686 ( .A(t_172), .B(n[173]), .Z(t_173) );
  GTECH_XOR2 C687 ( .A(t_173), .B(n[174]), .Z(t_174) );
  GTECH_XOR2 C688 ( .A(t_174), .B(n[175]), .Z(t_175) );
  GTECH_XOR2 C689 ( .A(t_175), .B(n[176]), .Z(t_176) );
  GTECH_XOR2 C690 ( .A(t_176), .B(n[177]), .Z(t_177) );
  GTECH_XOR2 C691 ( .A(t_177), .B(n[178]), .Z(t_178) );
  GTECH_XOR2 C692 ( .A(t_178), .B(n[179]), .Z(t_179) );
  GTECH_XOR2 C693 ( .A(t_179), .B(n[180]), .Z(t_180) );
  GTECH_XOR2 C694 ( .A(t_180), .B(n[181]), .Z(t_181) );
  GTECH_XOR2 C695 ( .A(t_181), .B(n[182]), .Z(t_182) );
  GTECH_XOR2 C696 ( .A(t_182), .B(n[183]), .Z(t_183) );
  GTECH_XOR2 C697 ( .A(t_183), .B(n[184]), .Z(t_184) );
  GTECH_XOR2 C698 ( .A(t_184), .B(n[185]), .Z(t_185) );
  GTECH_XOR2 C699 ( .A(t_185), .B(n[186]), .Z(t_186) );
  GTECH_XOR2 C700 ( .A(t_186), .B(n[187]), .Z(t_187) );
  GTECH_XOR2 C701 ( .A(t_187), .B(n[188]), .Z(t_188) );
  GTECH_XOR2 C702 ( .A(t_188), .B(n[189]), .Z(t_189) );
  GTECH_XOR2 C703 ( .A(t_189), .B(n[190]), .Z(t_190) );
  GTECH_XOR2 C704 ( .A(t_190), .B(n[191]), .Z(t_191) );
  GTECH_XOR2 C705 ( .A(t_191), .B(n[192]), .Z(t_192) );
  GTECH_XOR2 C706 ( .A(t_192), .B(n[193]), .Z(t_193) );
  GTECH_XOR2 C707 ( .A(t_193), .B(n[194]), .Z(t_194) );
  GTECH_XOR2 C708 ( .A(t_194), .B(n[195]), .Z(t_195) );
  GTECH_XOR2 C709 ( .A(t_195), .B(n[196]), .Z(t_196) );
  GTECH_XOR2 C710 ( .A(t_196), .B(n[197]), .Z(t_197) );
  GTECH_XOR2 C711 ( .A(t_197), .B(n[198]), .Z(t_198) );
  GTECH_XOR2 C712 ( .A(t_198), .B(n[199]), .Z(t_199) );
  GTECH_XOR2 C713 ( .A(t_199), .B(n[200]), .Z(t_200) );
  GTECH_XOR2 C714 ( .A(t_200), .B(n[201]), .Z(t_201) );
  GTECH_XOR2 C715 ( .A(t_201), .B(n[202]), .Z(t_202) );
  GTECH_XOR2 C716 ( .A(t_202), .B(n[203]), .Z(t_203) );
  GTECH_XOR2 C717 ( .A(t_203), .B(n[204]), .Z(t_204) );
  GTECH_XOR2 C718 ( .A(t_204), .B(n[205]), .Z(t_205) );
  GTECH_XOR2 C719 ( .A(t_205), .B(n[206]), .Z(t_206) );
  GTECH_XOR2 C720 ( .A(t_206), .B(n[207]), .Z(t_207) );
  GTECH_XOR2 C721 ( .A(t_207), .B(n[208]), .Z(t_208) );
  GTECH_XOR2 C722 ( .A(t_208), .B(n[209]), .Z(t_209) );
  GTECH_XOR2 C723 ( .A(t_209), .B(n[210]), .Z(t_210) );
  GTECH_XOR2 C724 ( .A(t_210), .B(n[211]), .Z(t_211) );
  GTECH_XOR2 C725 ( .A(t_211), .B(n[212]), .Z(t_212) );
  GTECH_XOR2 C726 ( .A(t_212), .B(n[213]), .Z(t_213) );
  GTECH_XOR2 C727 ( .A(t_213), .B(n[214]), .Z(t_214) );
  GTECH_XOR2 C728 ( .A(t_214), .B(n[215]), .Z(t_215) );
  GTECH_XOR2 C729 ( .A(t_215), .B(n[216]), .Z(t_216) );
  GTECH_XOR2 C730 ( .A(t_216), .B(n[217]), .Z(t_217) );
  GTECH_XOR2 C731 ( .A(t_217), .B(n[218]), .Z(t_218) );
  GTECH_XOR2 C732 ( .A(t_218), .B(n[219]), .Z(t_219) );
  GTECH_XOR2 C733 ( .A(t_219), .B(n[220]), .Z(t_220) );
  GTECH_XOR2 C734 ( .A(t_220), .B(n[221]), .Z(t_221) );
  GTECH_XOR2 C735 ( .A(t_221), .B(n[222]), .Z(t_222) );
  GTECH_XOR2 C736 ( .A(t_222), .B(n[223]), .Z(t_223) );
  GTECH_XOR2 C737 ( .A(t_223), .B(n[224]), .Z(t_224) );
  GTECH_XOR2 C738 ( .A(t_224), .B(n[225]), .Z(t_225) );
  GTECH_XOR2 C739 ( .A(t_225), .B(n[226]), .Z(t_226) );
  GTECH_XOR2 C740 ( .A(t_226), .B(n[227]), .Z(t_227) );
  GTECH_XOR2 C741 ( .A(t_227), .B(n[228]), .Z(t_228) );
  GTECH_XOR2 C742 ( .A(t_228), .B(n[229]), .Z(t_229) );
  GTECH_XOR2 C743 ( .A(t_229), .B(n[230]), .Z(t_230) );
  GTECH_XOR2 C744 ( .A(t_230), .B(n[231]), .Z(t_231) );
  GTECH_XOR2 C745 ( .A(t_231), .B(n[232]), .Z(t_232) );
  GTECH_XOR2 C746 ( .A(t_232), .B(n[233]), .Z(t_233) );
  GTECH_XOR2 C747 ( .A(t_233), .B(n[234]), .Z(t_234) );
  GTECH_XOR2 C748 ( .A(t_234), .B(n[235]), .Z(t_235) );
  GTECH_XOR2 C749 ( .A(t_235), .B(n[236]), .Z(t_236) );
  GTECH_XOR2 C750 ( .A(t_236), .B(n[237]), .Z(t_237) );
  GTECH_XOR2 C751 ( .A(t_237), .B(n[238]), .Z(t_238) );
  GTECH_XOR2 C752 ( .A(t_238), .B(n[239]), .Z(t_239) );
  GTECH_XOR2 C753 ( .A(t_239), .B(n[240]), .Z(t_240) );
  GTECH_XOR2 C754 ( .A(t_240), .B(n[241]), .Z(t_241) );
  GTECH_XOR2 C755 ( .A(t_241), .B(n[242]), .Z(t_242) );
  GTECH_XOR2 C756 ( .A(t_242), .B(n[243]), .Z(t_243) );
  GTECH_XOR2 C757 ( .A(t_243), .B(n[244]), .Z(t_244) );
  GTECH_XOR2 C758 ( .A(t_244), .B(n[245]), .Z(t_245) );
  GTECH_XOR2 C759 ( .A(N6), .B(t_245), .Z(s[6]) );
  GTECH_XOR2 C760 ( .A(a[6]), .B(b[6]), .Z(N6) );
  GTECH_XOR2 C761 ( .A(n[246]), .B(n[247]), .Z(t[247]) );
  GTECH_XOR2 C762 ( .A(t[247]), .B(n[248]), .Z(t[248]) );
  GTECH_XOR2 C763 ( .A(t[248]), .B(n[249]), .Z(t[249]) );
  GTECH_XOR2 C764 ( .A(t[249]), .B(n[250]), .Z(t[250]) );
  GTECH_XOR2 C765 ( .A(t[250]), .B(n[251]), .Z(t[251]) );
  GTECH_XOR2 C766 ( .A(t[251]), .B(n[252]), .Z(t[252]) );
  GTECH_XOR2 C767 ( .A(t[252]), .B(n[253]), .Z(t[253]) );
  GTECH_XOR2 C768 ( .A(t[253]), .B(n[254]), .Z(t[254]) );
  GTECH_XOR2 C769 ( .A(t[254]), .B(n[255]), .Z(t[255]) );
  GTECH_XOR2 C770 ( .A(t[255]), .B(n[256]), .Z(t[256]) );
  GTECH_XOR2 C771 ( .A(t[256]), .B(n[257]), .Z(t[257]) );
  GTECH_XOR2 C772 ( .A(t[257]), .B(n[258]), .Z(t[258]) );
  GTECH_XOR2 C773 ( .A(t[258]), .B(n[259]), .Z(t[259]) );
  GTECH_XOR2 C774 ( .A(t[259]), .B(n[260]), .Z(t[260]) );
  GTECH_XOR2 C775 ( .A(t[260]), .B(n[261]), .Z(t[261]) );
  GTECH_XOR2 C776 ( .A(t[261]), .B(n[262]), .Z(t[262]) );
  GTECH_XOR2 C777 ( .A(t[262]), .B(n[263]), .Z(t[263]) );
  GTECH_XOR2 C778 ( .A(t[263]), .B(n[264]), .Z(t[264]) );
  GTECH_XOR2 C779 ( .A(t[264]), .B(n[265]), .Z(t[265]) );
  GTECH_XOR2 C780 ( .A(t[265]), .B(n[266]), .Z(t[266]) );
  GTECH_XOR2 C781 ( .A(t[266]), .B(n[267]), .Z(t[267]) );
  GTECH_XOR2 C782 ( .A(t[267]), .B(n[268]), .Z(t[268]) );
  GTECH_XOR2 C783 ( .A(t[268]), .B(n[269]), .Z(t[269]) );
  GTECH_XOR2 C784 ( .A(t[269]), .B(n[270]), .Z(t[270]) );
  GTECH_XOR2 C785 ( .A(t[270]), .B(n[271]), .Z(t[271]) );
  GTECH_XOR2 C786 ( .A(t[271]), .B(n[272]), .Z(t[272]) );
  GTECH_XOR2 C787 ( .A(t[272]), .B(n[273]), .Z(t[273]) );
  GTECH_XOR2 C788 ( .A(t[273]), .B(n[274]), .Z(t[274]) );
  GTECH_XOR2 C789 ( .A(t[274]), .B(n[275]), .Z(t[275]) );
  GTECH_XOR2 C790 ( .A(t[275]), .B(n[276]), .Z(t[276]) );
  GTECH_XOR2 C791 ( .A(t[276]), .B(n[277]), .Z(t[277]) );
  GTECH_XOR2 C792 ( .A(t[277]), .B(n[278]), .Z(t[278]) );
  GTECH_XOR2 C793 ( .A(t[278]), .B(n[279]), .Z(t[279]) );
  GTECH_XOR2 C794 ( .A(t[279]), .B(n[280]), .Z(t[280]) );
  GTECH_XOR2 C795 ( .A(t[280]), .B(n[281]), .Z(t[281]) );
  GTECH_XOR2 C796 ( .A(t[281]), .B(n[282]), .Z(t[282]) );
  GTECH_XOR2 C797 ( .A(t[282]), .B(n[283]), .Z(t[283]) );
  GTECH_XOR2 C798 ( .A(t[283]), .B(n[284]), .Z(t[284]) );
  GTECH_XOR2 C799 ( .A(t[284]), .B(n[285]), .Z(t[285]) );
  GTECH_XOR2 C800 ( .A(t[285]), .B(n[286]), .Z(t[286]) );
  GTECH_XOR2 C801 ( .A(t[286]), .B(n[287]), .Z(t[287]) );
  GTECH_XOR2 C802 ( .A(t[287]), .B(n[288]), .Z(t[288]) );
  GTECH_XOR2 C803 ( .A(t[288]), .B(n[289]), .Z(t[289]) );
  GTECH_XOR2 C804 ( .A(t[289]), .B(n[290]), .Z(t[290]) );
  GTECH_XOR2 C805 ( .A(t[290]), .B(n[291]), .Z(t[291]) );
  GTECH_XOR2 C806 ( .A(t[291]), .B(n[292]), .Z(t[292]) );
  GTECH_XOR2 C807 ( .A(t[292]), .B(n[293]), .Z(t[293]) );
  GTECH_XOR2 C808 ( .A(t[293]), .B(n[294]), .Z(t[294]) );
  GTECH_XOR2 C809 ( .A(t[294]), .B(n[295]), .Z(t[295]) );
  GTECH_XOR2 C810 ( .A(t[295]), .B(n[296]), .Z(t[296]) );
  GTECH_XOR2 C811 ( .A(t[296]), .B(n[297]), .Z(t[297]) );
  GTECH_XOR2 C812 ( .A(t[297]), .B(n[298]), .Z(t[298]) );
  GTECH_XOR2 C813 ( .A(t[298]), .B(n[299]), .Z(t[299]) );
  GTECH_XOR2 C814 ( .A(t[299]), .B(n[300]), .Z(t[300]) );
  GTECH_XOR2 C815 ( .A(t[300]), .B(n[301]), .Z(t[301]) );
  GTECH_XOR2 C816 ( .A(t[301]), .B(n[302]), .Z(t[302]) );
  GTECH_XOR2 C817 ( .A(t[302]), .B(n[303]), .Z(t[303]) );
  GTECH_XOR2 C818 ( .A(t[303]), .B(n[304]), .Z(t[304]) );
  GTECH_XOR2 C819 ( .A(t[304]), .B(n[305]), .Z(t[305]) );
  GTECH_XOR2 C820 ( .A(t[305]), .B(n[306]), .Z(t[306]) );
  GTECH_XOR2 C821 ( .A(t[306]), .B(n[307]), .Z(t[307]) );
  GTECH_XOR2 C822 ( .A(t[307]), .B(n[308]), .Z(t[308]) );
  GTECH_XOR2 C823 ( .A(t[308]), .B(n[309]), .Z(t[309]) );
  GTECH_XOR2 C824 ( .A(t[309]), .B(n[310]), .Z(t[310]) );
  GTECH_XOR2 C825 ( .A(t[310]), .B(n[311]), .Z(t[311]) );
  GTECH_XOR2 C826 ( .A(t[311]), .B(n[312]), .Z(t[312]) );
  GTECH_XOR2 C827 ( .A(t[312]), .B(n[313]), .Z(t[313]) );
  GTECH_XOR2 C828 ( .A(t[313]), .B(n[314]), .Z(t[314]) );
  GTECH_XOR2 C829 ( .A(t[314]), .B(n[315]), .Z(t[315]) );
  GTECH_XOR2 C830 ( .A(t[315]), .B(n[316]), .Z(t[316]) );
  GTECH_XOR2 C831 ( .A(t[316]), .B(n[317]), .Z(t[317]) );
  GTECH_XOR2 C832 ( .A(t[317]), .B(n[318]), .Z(t[318]) );
  GTECH_XOR2 C833 ( .A(t[318]), .B(n[319]), .Z(t[319]) );
  GTECH_XOR2 C834 ( .A(t[319]), .B(n[320]), .Z(t[320]) );
  GTECH_XOR2 C835 ( .A(t[320]), .B(n[321]), .Z(t[321]) );
  GTECH_XOR2 C836 ( .A(t[321]), .B(n[322]), .Z(t[322]) );
  GTECH_XOR2 C837 ( .A(t[322]), .B(n[323]), .Z(t[323]) );
  GTECH_XOR2 C838 ( .A(t[323]), .B(n[324]), .Z(t[324]) );
  GTECH_XOR2 C839 ( .A(t[324]), .B(n[325]), .Z(t[325]) );
  GTECH_XOR2 C840 ( .A(t[325]), .B(n[326]), .Z(t[326]) );
  GTECH_XOR2 C841 ( .A(t[326]), .B(n[327]), .Z(t[327]) );
  GTECH_XOR2 C842 ( .A(t[327]), .B(n[328]), .Z(t[328]) );
  GTECH_XOR2 C843 ( .A(t[328]), .B(n[329]), .Z(t[329]) );
  GTECH_XOR2 C844 ( .A(t[329]), .B(n[330]), .Z(t[330]) );
  GTECH_XOR2 C845 ( .A(t[330]), .B(n[331]), .Z(t[331]) );
  GTECH_XOR2 C846 ( .A(t[331]), .B(n[332]), .Z(t[332]) );
  GTECH_XOR2 C847 ( .A(t[332]), .B(n[333]), .Z(t[333]) );
  GTECH_XOR2 C848 ( .A(t[333]), .B(n[334]), .Z(t[334]) );
  GTECH_XOR2 C849 ( .A(t[334]), .B(n[335]), .Z(t[335]) );
  GTECH_XOR2 C850 ( .A(t[335]), .B(n[336]), .Z(t[336]) );
  GTECH_XOR2 C851 ( .A(t[336]), .B(n[337]), .Z(t[337]) );
  GTECH_XOR2 C852 ( .A(t[337]), .B(n[338]), .Z(t[338]) );
  GTECH_XOR2 C853 ( .A(t[338]), .B(n[339]), .Z(t[339]) );
  GTECH_XOR2 C854 ( .A(t[339]), .B(n[340]), .Z(t[340]) );
  GTECH_XOR2 C855 ( .A(t[340]), .B(n[341]), .Z(t[341]) );
  GTECH_XOR2 C856 ( .A(t[341]), .B(n[342]), .Z(t[342]) );
  GTECH_XOR2 C857 ( .A(t[342]), .B(n[343]), .Z(t[343]) );
  GTECH_XOR2 C858 ( .A(t[343]), .B(n[344]), .Z(t[344]) );
  GTECH_XOR2 C859 ( .A(t[344]), .B(n[345]), .Z(t[345]) );
  GTECH_XOR2 C860 ( .A(t[345]), .B(n[346]), .Z(t[346]) );
  GTECH_XOR2 C861 ( .A(t[346]), .B(n[347]), .Z(t[347]) );
  GTECH_XOR2 C862 ( .A(t[347]), .B(n[348]), .Z(t[348]) );
  GTECH_XOR2 C863 ( .A(t[348]), .B(n[349]), .Z(t[349]) );
  GTECH_XOR2 C864 ( .A(t[349]), .B(n[350]), .Z(t[350]) );
  GTECH_XOR2 C865 ( .A(t[350]), .B(n[351]), .Z(t[351]) );
  GTECH_XOR2 C866 ( .A(t[351]), .B(n[352]), .Z(t[352]) );
  GTECH_XOR2 C867 ( .A(t[352]), .B(n[353]), .Z(t[353]) );
  GTECH_XOR2 C868 ( .A(t[353]), .B(n[354]), .Z(t[354]) );
  GTECH_XOR2 C869 ( .A(t[354]), .B(n[355]), .Z(t[355]) );
  GTECH_XOR2 C870 ( .A(t[355]), .B(n[356]), .Z(t[356]) );
  GTECH_XOR2 C871 ( .A(t[356]), .B(n[357]), .Z(t[357]) );
  GTECH_XOR2 C872 ( .A(t[357]), .B(n[358]), .Z(t[358]) );
  GTECH_XOR2 C873 ( .A(t[358]), .B(n[359]), .Z(t[359]) );
  GTECH_XOR2 C874 ( .A(t[359]), .B(n[360]), .Z(t[360]) );
  GTECH_XOR2 C875 ( .A(t[360]), .B(n[361]), .Z(t[361]) );
  GTECH_XOR2 C876 ( .A(t[361]), .B(n[362]), .Z(t[362]) );
  GTECH_XOR2 C877 ( .A(t[362]), .B(n[363]), .Z(t[363]) );
  GTECH_XOR2 C878 ( .A(t[363]), .B(n[364]), .Z(t[364]) );
  GTECH_XOR2 C879 ( .A(t[364]), .B(n[365]), .Z(t[365]) );
  GTECH_XOR2 C880 ( .A(t[365]), .B(n[366]), .Z(t[366]) );
  GTECH_XOR2 C881 ( .A(t[366]), .B(n[367]), .Z(t[367]) );
  GTECH_XOR2 C882 ( .A(t[367]), .B(n[368]), .Z(t[368]) );
  GTECH_XOR2 C883 ( .A(t[368]), .B(n[369]), .Z(t[369]) );
  GTECH_XOR2 C884 ( .A(t[369]), .B(n[370]), .Z(t[370]) );
  GTECH_XOR2 C885 ( .A(t[370]), .B(n[371]), .Z(t[371]) );
  GTECH_XOR2 C886 ( .A(t[371]), .B(n[372]), .Z(t[372]) );
  GTECH_XOR2 C887 ( .A(t[372]), .B(n[373]), .Z(t[373]) );
  GTECH_XOR2 C888 ( .A(t[373]), .B(n[374]), .Z(t[374]) );
  GTECH_XOR2 C889 ( .A(t[374]), .B(n[375]), .Z(t[375]) );
  GTECH_XOR2 C890 ( .A(t[375]), .B(n[376]), .Z(t[376]) );
  GTECH_XOR2 C891 ( .A(t[376]), .B(n[377]), .Z(t[377]) );
  GTECH_XOR2 C892 ( .A(t[377]), .B(n[378]), .Z(t[378]) );
  GTECH_XOR2 C893 ( .A(t[378]), .B(n[379]), .Z(t[379]) );
  GTECH_XOR2 C894 ( .A(t[379]), .B(n[380]), .Z(t[380]) );
  GTECH_XOR2 C895 ( .A(t[380]), .B(n[381]), .Z(t[381]) );
  GTECH_XOR2 C896 ( .A(t[381]), .B(n[382]), .Z(t[382]) );
  GTECH_XOR2 C897 ( .A(t[382]), .B(n[383]), .Z(t[383]) );
  GTECH_XOR2 C898 ( .A(t[383]), .B(n[384]), .Z(t[384]) );
  GTECH_XOR2 C899 ( .A(t[384]), .B(n[385]), .Z(t[385]) );
  GTECH_XOR2 C900 ( .A(t[385]), .B(n[386]), .Z(t[386]) );
  GTECH_XOR2 C901 ( .A(t[386]), .B(n[387]), .Z(t[387]) );
  GTECH_XOR2 C902 ( .A(t[387]), .B(n[388]), .Z(t[388]) );
  GTECH_XOR2 C903 ( .A(t[388]), .B(n[389]), .Z(t[389]) );
  GTECH_XOR2 C904 ( .A(t[389]), .B(n[390]), .Z(t[390]) );
  GTECH_XOR2 C905 ( .A(t[390]), .B(n[391]), .Z(t[391]) );
  GTECH_XOR2 C906 ( .A(t[391]), .B(n[392]), .Z(t[392]) );
  GTECH_XOR2 C907 ( .A(t[392]), .B(n[393]), .Z(t[393]) );
  GTECH_XOR2 C908 ( .A(t[393]), .B(n[394]), .Z(t[394]) );
  GTECH_XOR2 C909 ( .A(t[394]), .B(n[395]), .Z(t[395]) );
  GTECH_XOR2 C910 ( .A(t[395]), .B(n[396]), .Z(t[396]) );
  GTECH_XOR2 C911 ( .A(t[396]), .B(n[397]), .Z(t[397]) );
  GTECH_XOR2 C912 ( .A(t[397]), .B(n[398]), .Z(t[398]) );
  GTECH_XOR2 C913 ( .A(t[398]), .B(n[399]), .Z(t[399]) );
  GTECH_XOR2 C914 ( .A(t[399]), .B(n[400]), .Z(t[400]) );
  GTECH_XOR2 C915 ( .A(t[400]), .B(n[401]), .Z(t[401]) );
  GTECH_XOR2 C916 ( .A(t[401]), .B(n[402]), .Z(t[402]) );
  GTECH_XOR2 C917 ( .A(t[402]), .B(n[403]), .Z(t[403]) );
  GTECH_XOR2 C918 ( .A(t[403]), .B(n[404]), .Z(t[404]) );
  GTECH_XOR2 C919 ( .A(t[404]), .B(n[405]), .Z(t[405]) );
  GTECH_XOR2 C920 ( .A(t[405]), .B(n[406]), .Z(t[406]) );
  GTECH_XOR2 C921 ( .A(t[406]), .B(n[407]), .Z(t[407]) );
  GTECH_XOR2 C922 ( .A(t[407]), .B(n[408]), .Z(t[408]) );
  GTECH_XOR2 C923 ( .A(t[408]), .B(n[409]), .Z(t[409]) );
  GTECH_XOR2 C924 ( .A(t[409]), .B(n[410]), .Z(t[410]) );
  GTECH_XOR2 C925 ( .A(t[410]), .B(n[411]), .Z(t[411]) );
  GTECH_XOR2 C926 ( .A(t[411]), .B(n[412]), .Z(t[412]) );
  GTECH_XOR2 C927 ( .A(t[412]), .B(n[413]), .Z(t[413]) );
  GTECH_XOR2 C928 ( .A(t[413]), .B(n[414]), .Z(t[414]) );
  GTECH_XOR2 C929 ( .A(t[414]), .B(n[415]), .Z(t[415]) );
  GTECH_XOR2 C930 ( .A(t[415]), .B(n[416]), .Z(t[416]) );
  GTECH_XOR2 C931 ( .A(t[416]), .B(n[417]), .Z(t[417]) );
  GTECH_XOR2 C932 ( .A(t[417]), .B(n[418]), .Z(t[418]) );
  GTECH_XOR2 C933 ( .A(t[418]), .B(n[419]), .Z(t[419]) );
  GTECH_XOR2 C934 ( .A(t[419]), .B(n[420]), .Z(t[420]) );
  GTECH_XOR2 C935 ( .A(t[420]), .B(n[421]), .Z(t[421]) );
  GTECH_XOR2 C936 ( .A(t[421]), .B(n[422]), .Z(t[422]) );
  GTECH_XOR2 C937 ( .A(t[422]), .B(n[423]), .Z(t[423]) );
  GTECH_XOR2 C938 ( .A(t[423]), .B(n[424]), .Z(t[424]) );
  GTECH_XOR2 C939 ( .A(t[424]), .B(n[425]), .Z(t[425]) );
  GTECH_XOR2 C940 ( .A(t[425]), .B(n[426]), .Z(t[426]) );
  GTECH_XOR2 C941 ( .A(t[426]), .B(n[427]), .Z(t[427]) );
  GTECH_XOR2 C942 ( .A(t[427]), .B(n[428]), .Z(t[428]) );
  GTECH_XOR2 C943 ( .A(t[428]), .B(n[429]), .Z(t[429]) );
  GTECH_XOR2 C944 ( .A(t[429]), .B(n[430]), .Z(t[430]) );
  GTECH_XOR2 C945 ( .A(t[430]), .B(n[431]), .Z(t[431]) );
  GTECH_XOR2 C946 ( .A(t[431]), .B(n[432]), .Z(t[432]) );
  GTECH_XOR2 C947 ( .A(t[432]), .B(n[433]), .Z(t[433]) );
  GTECH_XOR2 C948 ( .A(t[433]), .B(n[434]), .Z(t[434]) );
  GTECH_XOR2 C949 ( .A(t[434]), .B(n[435]), .Z(t[435]) );
  GTECH_XOR2 C950 ( .A(t[435]), .B(n[436]), .Z(t[436]) );
  GTECH_XOR2 C951 ( .A(t[436]), .B(n[437]), .Z(t[437]) );
  GTECH_XOR2 C952 ( .A(t[437]), .B(n[438]), .Z(t[438]) );
  GTECH_XOR2 C953 ( .A(t[438]), .B(n[439]), .Z(t[439]) );
  GTECH_XOR2 C954 ( .A(t[439]), .B(n[440]), .Z(t[440]) );
  GTECH_XOR2 C955 ( .A(t[440]), .B(n[441]), .Z(t[441]) );
  GTECH_XOR2 C956 ( .A(t[441]), .B(n[442]), .Z(t[442]) );
  GTECH_XOR2 C957 ( .A(t[442]), .B(n[443]), .Z(t[443]) );
  GTECH_XOR2 C958 ( .A(t[443]), .B(n[444]), .Z(t[444]) );
  GTECH_XOR2 C959 ( .A(t[444]), .B(n[445]), .Z(t[445]) );
  GTECH_XOR2 C960 ( .A(t[445]), .B(n[446]), .Z(t[446]) );
  GTECH_XOR2 C961 ( .A(t[446]), .B(n[447]), .Z(t[447]) );
  GTECH_XOR2 C962 ( .A(t[447]), .B(n[448]), .Z(t[448]) );
  GTECH_XOR2 C963 ( .A(t[448]), .B(n[449]), .Z(t[449]) );
  GTECH_XOR2 C964 ( .A(t[449]), .B(n[450]), .Z(t[450]) );
  GTECH_XOR2 C965 ( .A(t[450]), .B(n[451]), .Z(t[451]) );
  GTECH_XOR2 C966 ( .A(t[451]), .B(n[452]), .Z(t[452]) );
  GTECH_XOR2 C967 ( .A(t[452]), .B(n[453]), .Z(t[453]) );
  GTECH_XOR2 C968 ( .A(t[453]), .B(n[454]), .Z(t[454]) );
  GTECH_XOR2 C969 ( .A(t[454]), .B(n[455]), .Z(t[455]) );
  GTECH_XOR2 C970 ( .A(t[455]), .B(n[456]), .Z(t[456]) );
  GTECH_XOR2 C971 ( .A(t[456]), .B(n[457]), .Z(t[457]) );
  GTECH_XOR2 C972 ( .A(t[457]), .B(n[458]), .Z(t[458]) );
  GTECH_XOR2 C973 ( .A(t[458]), .B(n[459]), .Z(t[459]) );
  GTECH_XOR2 C974 ( .A(t[459]), .B(n[460]), .Z(t[460]) );
  GTECH_XOR2 C975 ( .A(t[460]), .B(n[461]), .Z(t[461]) );
  GTECH_XOR2 C976 ( .A(t[461]), .B(n[462]), .Z(t[462]) );
  GTECH_XOR2 C977 ( .A(t[462]), .B(n[463]), .Z(t[463]) );
  GTECH_XOR2 C978 ( .A(t[463]), .B(n[464]), .Z(t[464]) );
  GTECH_XOR2 C979 ( .A(t[464]), .B(n[465]), .Z(t[465]) );
  GTECH_XOR2 C980 ( .A(t[465]), .B(n[466]), .Z(t[466]) );
  GTECH_XOR2 C981 ( .A(t[466]), .B(n[467]), .Z(t[467]) );
  GTECH_XOR2 C982 ( .A(t[467]), .B(n[468]), .Z(t[468]) );
  GTECH_XOR2 C983 ( .A(t[468]), .B(n[469]), .Z(t[469]) );
  GTECH_XOR2 C984 ( .A(t[469]), .B(n[470]), .Z(t[470]) );
  GTECH_XOR2 C985 ( .A(t[470]), .B(n[471]), .Z(t[471]) );
  GTECH_XOR2 C986 ( .A(t[471]), .B(n[472]), .Z(t[472]) );
  GTECH_XOR2 C987 ( .A(t[472]), .B(n[473]), .Z(t[473]) );
  GTECH_XOR2 C988 ( .A(t[473]), .B(n[474]), .Z(t[474]) );
  GTECH_XOR2 C989 ( .A(t[474]), .B(n[475]), .Z(t[475]) );
  GTECH_XOR2 C990 ( .A(t[475]), .B(n[476]), .Z(t[476]) );
  GTECH_XOR2 C991 ( .A(t[476]), .B(n[477]), .Z(t[477]) );
  GTECH_XOR2 C992 ( .A(t[477]), .B(n[478]), .Z(t[478]) );
  GTECH_XOR2 C993 ( .A(t[478]), .B(n[479]), .Z(t[479]) );
  GTECH_XOR2 C994 ( .A(t[479]), .B(n[480]), .Z(t[480]) );
  GTECH_XOR2 C995 ( .A(t[480]), .B(n[481]), .Z(t[481]) );
  GTECH_XOR2 C996 ( .A(t[481]), .B(n[482]), .Z(t[482]) );
  GTECH_XOR2 C997 ( .A(t[482]), .B(n[483]), .Z(t[483]) );
  GTECH_XOR2 C998 ( .A(t[483]), .B(n[484]), .Z(t[484]) );
  GTECH_XOR2 C999 ( .A(t[484]), .B(n[485]), .Z(t[485]) );
  GTECH_XOR2 C1000 ( .A(t[485]), .B(n[486]), .Z(t[486]) );
  GTECH_XOR2 C1001 ( .A(t[486]), .B(n[487]), .Z(t[487]) );
  GTECH_XOR2 C1002 ( .A(t[487]), .B(n[488]), .Z(t[488]) );
  GTECH_XOR2 C1003 ( .A(t[488]), .B(n[489]), .Z(t[489]) );
  GTECH_XOR2 C1004 ( .A(t[489]), .B(n[490]), .Z(t[490]) );
  GTECH_XOR2 C1005 ( .A(t[490]), .B(n[491]), .Z(t[491]) );
  GTECH_XOR2 C1006 ( .A(t[491]), .B(n[492]), .Z(t[492]) );
  GTECH_XOR2 C1007 ( .A(t[492]), .B(n[493]), .Z(t[493]) );
  GTECH_XOR2 C1008 ( .A(t[493]), .B(n[494]), .Z(t[494]) );
  GTECH_XOR2 C1009 ( .A(t[494]), .B(n[495]), .Z(t[495]) );
  GTECH_XOR2 C1010 ( .A(t[495]), .B(n[496]), .Z(t[496]) );
  GTECH_XOR2 C1011 ( .A(t[496]), .B(n[497]), .Z(t[497]) );
  GTECH_XOR2 C1012 ( .A(t[497]), .B(n[498]), .Z(t[498]) );
  GTECH_XOR2 C1013 ( .A(t[498]), .B(n[499]), .Z(t[499]) );
  GTECH_XOR2 C1014 ( .A(t[499]), .B(n[500]), .Z(s[7]) );
endmodule


module gen_nonlinear_part ( a, b, c, n );
  input [6:0] a;
  input [6:0] b;
  output [500:0] n;
  input c;


  GTECH_AND2 C507 ( .A(a[0]), .B(b[0]), .Z(n[0]) );
  GTECH_AND2 C508 ( .A(a[0]), .B(c), .Z(n[1]) );
  GTECH_AND2 C509 ( .A(b[0]), .B(c), .Z(n[2]) );
  GTECH_AND2 C510 ( .A(a[1]), .B(b[1]), .Z(n[3]) );
  GTECH_AND2 C511 ( .A(a[1]), .B(n[0]), .Z(n[4]) );
  GTECH_AND2 C512 ( .A(b[1]), .B(n[0]), .Z(n[7]) );
  GTECH_AND2 C513 ( .A(a[1]), .B(n[1]), .Z(n[5]) );
  GTECH_AND2 C514 ( .A(b[1]), .B(n[1]), .Z(n[8]) );
  GTECH_AND2 C515 ( .A(a[1]), .B(n[2]), .Z(n[6]) );
  GTECH_AND2 C516 ( .A(b[1]), .B(n[2]), .Z(n[9]) );
  GTECH_AND2 C517 ( .A(a[2]), .B(b[2]), .Z(n[10]) );
  GTECH_AND2 C518 ( .A(a[2]), .B(n[3]), .Z(n[11]) );
  GTECH_AND2 C519 ( .A(b[2]), .B(n[3]), .Z(n[18]) );
  GTECH_AND2 C520 ( .A(a[2]), .B(n[4]), .Z(n[12]) );
  GTECH_AND2 C521 ( .A(b[2]), .B(n[4]), .Z(n[19]) );
  GTECH_AND2 C522 ( .A(a[2]), .B(n[5]), .Z(n[13]) );
  GTECH_AND2 C523 ( .A(b[2]), .B(n[5]), .Z(n[20]) );
  GTECH_AND2 C524 ( .A(a[2]), .B(n[6]), .Z(n[14]) );
  GTECH_AND2 C525 ( .A(b[2]), .B(n[6]), .Z(n[21]) );
  GTECH_AND2 C526 ( .A(a[2]), .B(n[7]), .Z(n[15]) );
  GTECH_AND2 C527 ( .A(b[2]), .B(n[7]), .Z(n[22]) );
  GTECH_AND2 C528 ( .A(a[2]), .B(n[8]), .Z(n[16]) );
  GTECH_AND2 C529 ( .A(b[2]), .B(n[8]), .Z(n[23]) );
  GTECH_AND2 C530 ( .A(a[2]), .B(n[9]), .Z(n[17]) );
  GTECH_AND2 C531 ( .A(b[2]), .B(n[9]), .Z(n[24]) );
  GTECH_AND2 C532 ( .A(a[3]), .B(b[3]), .Z(n[25]) );
  GTECH_AND2 C533 ( .A(a[3]), .B(n[10]), .Z(n[26]) );
  GTECH_AND2 C534 ( .A(b[3]), .B(n[10]), .Z(n[41]) );
  GTECH_AND2 C535 ( .A(a[3]), .B(n[11]), .Z(n[27]) );
  GTECH_AND2 C536 ( .A(b[3]), .B(n[11]), .Z(n[42]) );
  GTECH_AND2 C537 ( .A(a[3]), .B(n[12]), .Z(n[28]) );
  GTECH_AND2 C538 ( .A(b[3]), .B(n[12]), .Z(n[43]) );
  GTECH_AND2 C539 ( .A(a[3]), .B(n[13]), .Z(n[29]) );
  GTECH_AND2 C540 ( .A(b[3]), .B(n[13]), .Z(n[44]) );
  GTECH_AND2 C541 ( .A(a[3]), .B(n[14]), .Z(n[30]) );
  GTECH_AND2 C542 ( .A(b[3]), .B(n[14]), .Z(n[45]) );
  GTECH_AND2 C543 ( .A(a[3]), .B(n[15]), .Z(n[31]) );
  GTECH_AND2 C544 ( .A(b[3]), .B(n[15]), .Z(n[46]) );
  GTECH_AND2 C545 ( .A(a[3]), .B(n[16]), .Z(n[32]) );
  GTECH_AND2 C546 ( .A(b[3]), .B(n[16]), .Z(n[47]) );
  GTECH_AND2 C547 ( .A(a[3]), .B(n[17]), .Z(n[33]) );
  GTECH_AND2 C548 ( .A(b[3]), .B(n[17]), .Z(n[48]) );
  GTECH_AND2 C549 ( .A(a[3]), .B(n[18]), .Z(n[34]) );
  GTECH_AND2 C550 ( .A(b[3]), .B(n[18]), .Z(n[49]) );
  GTECH_AND2 C551 ( .A(a[3]), .B(n[19]), .Z(n[35]) );
  GTECH_AND2 C552 ( .A(b[3]), .B(n[19]), .Z(n[50]) );
  GTECH_AND2 C553 ( .A(a[3]), .B(n[20]), .Z(n[36]) );
  GTECH_AND2 C554 ( .A(b[3]), .B(n[20]), .Z(n[51]) );
  GTECH_AND2 C555 ( .A(a[3]), .B(n[21]), .Z(n[37]) );
  GTECH_AND2 C556 ( .A(b[3]), .B(n[21]), .Z(n[52]) );
  GTECH_AND2 C557 ( .A(a[3]), .B(n[22]), .Z(n[38]) );
  GTECH_AND2 C558 ( .A(b[3]), .B(n[22]), .Z(n[53]) );
  GTECH_AND2 C559 ( .A(a[3]), .B(n[23]), .Z(n[39]) );
  GTECH_AND2 C560 ( .A(b[3]), .B(n[23]), .Z(n[54]) );
  GTECH_AND2 C561 ( .A(a[3]), .B(n[24]), .Z(n[40]) );
  GTECH_AND2 C562 ( .A(b[3]), .B(n[24]), .Z(n[55]) );
  GTECH_AND2 C563 ( .A(a[4]), .B(b[4]), .Z(n[56]) );
  GTECH_AND2 C564 ( .A(a[4]), .B(n[25]), .Z(n[57]) );
  GTECH_AND2 C565 ( .A(b[4]), .B(n[25]), .Z(n[88]) );
  GTECH_AND2 C566 ( .A(a[4]), .B(n[26]), .Z(n[58]) );
  GTECH_AND2 C567 ( .A(b[4]), .B(n[26]), .Z(n[89]) );
  GTECH_AND2 C568 ( .A(a[4]), .B(n[27]), .Z(n[59]) );
  GTECH_AND2 C569 ( .A(b[4]), .B(n[27]), .Z(n[90]) );
  GTECH_AND2 C570 ( .A(a[4]), .B(n[28]), .Z(n[60]) );
  GTECH_AND2 C571 ( .A(b[4]), .B(n[28]), .Z(n[91]) );
  GTECH_AND2 C572 ( .A(a[4]), .B(n[29]), .Z(n[61]) );
  GTECH_AND2 C573 ( .A(b[4]), .B(n[29]), .Z(n[92]) );
  GTECH_AND2 C574 ( .A(a[4]), .B(n[30]), .Z(n[62]) );
  GTECH_AND2 C575 ( .A(b[4]), .B(n[30]), .Z(n[93]) );
  GTECH_AND2 C576 ( .A(a[4]), .B(n[31]), .Z(n[63]) );
  GTECH_AND2 C577 ( .A(b[4]), .B(n[31]), .Z(n[94]) );
  GTECH_AND2 C578 ( .A(a[4]), .B(n[32]), .Z(n[64]) );
  GTECH_AND2 C579 ( .A(b[4]), .B(n[32]), .Z(n[95]) );
  GTECH_AND2 C580 ( .A(a[4]), .B(n[33]), .Z(n[65]) );
  GTECH_AND2 C581 ( .A(b[4]), .B(n[33]), .Z(n[96]) );
  GTECH_AND2 C582 ( .A(a[4]), .B(n[34]), .Z(n[66]) );
  GTECH_AND2 C583 ( .A(b[4]), .B(n[34]), .Z(n[97]) );
  GTECH_AND2 C584 ( .A(a[4]), .B(n[35]), .Z(n[67]) );
  GTECH_AND2 C585 ( .A(b[4]), .B(n[35]), .Z(n[98]) );
  GTECH_AND2 C586 ( .A(a[4]), .B(n[36]), .Z(n[68]) );
  GTECH_AND2 C587 ( .A(b[4]), .B(n[36]), .Z(n[99]) );
  GTECH_AND2 C588 ( .A(a[4]), .B(n[37]), .Z(n[69]) );
  GTECH_AND2 C589 ( .A(b[4]), .B(n[37]), .Z(n[100]) );
  GTECH_AND2 C590 ( .A(a[4]), .B(n[38]), .Z(n[70]) );
  GTECH_AND2 C591 ( .A(b[4]), .B(n[38]), .Z(n[101]) );
  GTECH_AND2 C592 ( .A(a[4]), .B(n[39]), .Z(n[71]) );
  GTECH_AND2 C593 ( .A(b[4]), .B(n[39]), .Z(n[102]) );
  GTECH_AND2 C594 ( .A(a[4]), .B(n[40]), .Z(n[72]) );
  GTECH_AND2 C595 ( .A(b[4]), .B(n[40]), .Z(n[103]) );
  GTECH_AND2 C596 ( .A(a[4]), .B(n[41]), .Z(n[73]) );
  GTECH_AND2 C597 ( .A(b[4]), .B(n[41]), .Z(n[104]) );
  GTECH_AND2 C598 ( .A(a[4]), .B(n[42]), .Z(n[74]) );
  GTECH_AND2 C599 ( .A(b[4]), .B(n[42]), .Z(n[105]) );
  GTECH_AND2 C600 ( .A(a[4]), .B(n[43]), .Z(n[75]) );
  GTECH_AND2 C601 ( .A(b[4]), .B(n[43]), .Z(n[106]) );
  GTECH_AND2 C602 ( .A(a[4]), .B(n[44]), .Z(n[76]) );
  GTECH_AND2 C603 ( .A(b[4]), .B(n[44]), .Z(n[107]) );
  GTECH_AND2 C604 ( .A(a[4]), .B(n[45]), .Z(n[77]) );
  GTECH_AND2 C605 ( .A(b[4]), .B(n[45]), .Z(n[108]) );
  GTECH_AND2 C606 ( .A(a[4]), .B(n[46]), .Z(n[78]) );
  GTECH_AND2 C607 ( .A(b[4]), .B(n[46]), .Z(n[109]) );
  GTECH_AND2 C608 ( .A(a[4]), .B(n[47]), .Z(n[79]) );
  GTECH_AND2 C609 ( .A(b[4]), .B(n[47]), .Z(n[110]) );
  GTECH_AND2 C610 ( .A(a[4]), .B(n[48]), .Z(n[80]) );
  GTECH_AND2 C611 ( .A(b[4]), .B(n[48]), .Z(n[111]) );
  GTECH_AND2 C612 ( .A(a[4]), .B(n[49]), .Z(n[81]) );
  GTECH_AND2 C613 ( .A(b[4]), .B(n[49]), .Z(n[112]) );
  GTECH_AND2 C614 ( .A(a[4]), .B(n[50]), .Z(n[82]) );
  GTECH_AND2 C615 ( .A(b[4]), .B(n[50]), .Z(n[113]) );
  GTECH_AND2 C616 ( .A(a[4]), .B(n[51]), .Z(n[83]) );
  GTECH_AND2 C617 ( .A(b[4]), .B(n[51]), .Z(n[114]) );
  GTECH_AND2 C618 ( .A(a[4]), .B(n[52]), .Z(n[84]) );
  GTECH_AND2 C619 ( .A(b[4]), .B(n[52]), .Z(n[115]) );
  GTECH_AND2 C620 ( .A(a[4]), .B(n[53]), .Z(n[85]) );
  GTECH_AND2 C621 ( .A(b[4]), .B(n[53]), .Z(n[116]) );
  GTECH_AND2 C622 ( .A(a[4]), .B(n[54]), .Z(n[86]) );
  GTECH_AND2 C623 ( .A(b[4]), .B(n[54]), .Z(n[117]) );
  GTECH_AND2 C624 ( .A(a[4]), .B(n[55]), .Z(n[87]) );
  GTECH_AND2 C625 ( .A(b[4]), .B(n[55]), .Z(n[118]) );
  GTECH_AND2 C626 ( .A(a[5]), .B(b[5]), .Z(n[119]) );
  GTECH_AND2 C627 ( .A(a[5]), .B(n[56]), .Z(n[120]) );
  GTECH_AND2 C628 ( .A(b[5]), .B(n[56]), .Z(n[183]) );
  GTECH_AND2 C629 ( .A(a[5]), .B(n[57]), .Z(n[121]) );
  GTECH_AND2 C630 ( .A(b[5]), .B(n[57]), .Z(n[184]) );
  GTECH_AND2 C631 ( .A(a[5]), .B(n[58]), .Z(n[122]) );
  GTECH_AND2 C632 ( .A(b[5]), .B(n[58]), .Z(n[185]) );
  GTECH_AND2 C633 ( .A(a[5]), .B(n[59]), .Z(n[123]) );
  GTECH_AND2 C634 ( .A(b[5]), .B(n[59]), .Z(n[186]) );
  GTECH_AND2 C635 ( .A(a[5]), .B(n[60]), .Z(n[124]) );
  GTECH_AND2 C636 ( .A(b[5]), .B(n[60]), .Z(n[187]) );
  GTECH_AND2 C637 ( .A(a[5]), .B(n[61]), .Z(n[125]) );
  GTECH_AND2 C638 ( .A(b[5]), .B(n[61]), .Z(n[188]) );
  GTECH_AND2 C639 ( .A(a[5]), .B(n[62]), .Z(n[126]) );
  GTECH_AND2 C640 ( .A(b[5]), .B(n[62]), .Z(n[189]) );
  GTECH_AND2 C641 ( .A(a[5]), .B(n[63]), .Z(n[127]) );
  GTECH_AND2 C642 ( .A(b[5]), .B(n[63]), .Z(n[190]) );
  GTECH_AND2 C643 ( .A(a[5]), .B(n[64]), .Z(n[128]) );
  GTECH_AND2 C644 ( .A(b[5]), .B(n[64]), .Z(n[191]) );
  GTECH_AND2 C645 ( .A(a[5]), .B(n[65]), .Z(n[129]) );
  GTECH_AND2 C646 ( .A(b[5]), .B(n[65]), .Z(n[192]) );
  GTECH_AND2 C647 ( .A(a[5]), .B(n[66]), .Z(n[130]) );
  GTECH_AND2 C648 ( .A(b[5]), .B(n[66]), .Z(n[193]) );
  GTECH_AND2 C649 ( .A(a[5]), .B(n[67]), .Z(n[131]) );
  GTECH_AND2 C650 ( .A(b[5]), .B(n[67]), .Z(n[194]) );
  GTECH_AND2 C651 ( .A(a[5]), .B(n[68]), .Z(n[132]) );
  GTECH_AND2 C652 ( .A(b[5]), .B(n[68]), .Z(n[195]) );
  GTECH_AND2 C653 ( .A(a[5]), .B(n[69]), .Z(n[133]) );
  GTECH_AND2 C654 ( .A(b[5]), .B(n[69]), .Z(n[196]) );
  GTECH_AND2 C655 ( .A(a[5]), .B(n[70]), .Z(n[134]) );
  GTECH_AND2 C656 ( .A(b[5]), .B(n[70]), .Z(n[197]) );
  GTECH_AND2 C657 ( .A(a[5]), .B(n[71]), .Z(n[135]) );
  GTECH_AND2 C658 ( .A(b[5]), .B(n[71]), .Z(n[198]) );
  GTECH_AND2 C659 ( .A(a[5]), .B(n[72]), .Z(n[136]) );
  GTECH_AND2 C660 ( .A(b[5]), .B(n[72]), .Z(n[199]) );
  GTECH_AND2 C661 ( .A(a[5]), .B(n[73]), .Z(n[137]) );
  GTECH_AND2 C662 ( .A(b[5]), .B(n[73]), .Z(n[200]) );
  GTECH_AND2 C663 ( .A(a[5]), .B(n[74]), .Z(n[138]) );
  GTECH_AND2 C664 ( .A(b[5]), .B(n[74]), .Z(n[201]) );
  GTECH_AND2 C665 ( .A(a[5]), .B(n[75]), .Z(n[139]) );
  GTECH_AND2 C666 ( .A(b[5]), .B(n[75]), .Z(n[202]) );
  GTECH_AND2 C667 ( .A(a[5]), .B(n[76]), .Z(n[140]) );
  GTECH_AND2 C668 ( .A(b[5]), .B(n[76]), .Z(n[203]) );
  GTECH_AND2 C669 ( .A(a[5]), .B(n[77]), .Z(n[141]) );
  GTECH_AND2 C670 ( .A(b[5]), .B(n[77]), .Z(n[204]) );
  GTECH_AND2 C671 ( .A(a[5]), .B(n[78]), .Z(n[142]) );
  GTECH_AND2 C672 ( .A(b[5]), .B(n[78]), .Z(n[205]) );
  GTECH_AND2 C673 ( .A(a[5]), .B(n[79]), .Z(n[143]) );
  GTECH_AND2 C674 ( .A(b[5]), .B(n[79]), .Z(n[206]) );
  GTECH_AND2 C675 ( .A(a[5]), .B(n[80]), .Z(n[144]) );
  GTECH_AND2 C676 ( .A(b[5]), .B(n[80]), .Z(n[207]) );
  GTECH_AND2 C677 ( .A(a[5]), .B(n[81]), .Z(n[145]) );
  GTECH_AND2 C678 ( .A(b[5]), .B(n[81]), .Z(n[208]) );
  GTECH_AND2 C679 ( .A(a[5]), .B(n[82]), .Z(n[146]) );
  GTECH_AND2 C680 ( .A(b[5]), .B(n[82]), .Z(n[209]) );
  GTECH_AND2 C681 ( .A(a[5]), .B(n[83]), .Z(n[147]) );
  GTECH_AND2 C682 ( .A(b[5]), .B(n[83]), .Z(n[210]) );
  GTECH_AND2 C683 ( .A(a[5]), .B(n[84]), .Z(n[148]) );
  GTECH_AND2 C684 ( .A(b[5]), .B(n[84]), .Z(n[211]) );
  GTECH_AND2 C685 ( .A(a[5]), .B(n[85]), .Z(n[149]) );
  GTECH_AND2 C686 ( .A(b[5]), .B(n[85]), .Z(n[212]) );
  GTECH_AND2 C687 ( .A(a[5]), .B(n[86]), .Z(n[150]) );
  GTECH_AND2 C688 ( .A(b[5]), .B(n[86]), .Z(n[213]) );
  GTECH_AND2 C689 ( .A(a[5]), .B(n[87]), .Z(n[151]) );
  GTECH_AND2 C690 ( .A(b[5]), .B(n[87]), .Z(n[214]) );
  GTECH_AND2 C691 ( .A(a[5]), .B(n[88]), .Z(n[152]) );
  GTECH_AND2 C692 ( .A(b[5]), .B(n[88]), .Z(n[215]) );
  GTECH_AND2 C693 ( .A(a[5]), .B(n[89]), .Z(n[153]) );
  GTECH_AND2 C694 ( .A(b[5]), .B(n[89]), .Z(n[216]) );
  GTECH_AND2 C695 ( .A(a[5]), .B(n[90]), .Z(n[154]) );
  GTECH_AND2 C696 ( .A(b[5]), .B(n[90]), .Z(n[217]) );
  GTECH_AND2 C697 ( .A(a[5]), .B(n[91]), .Z(n[155]) );
  GTECH_AND2 C698 ( .A(b[5]), .B(n[91]), .Z(n[218]) );
  GTECH_AND2 C699 ( .A(a[5]), .B(n[92]), .Z(n[156]) );
  GTECH_AND2 C700 ( .A(b[5]), .B(n[92]), .Z(n[219]) );
  GTECH_AND2 C701 ( .A(a[5]), .B(n[93]), .Z(n[157]) );
  GTECH_AND2 C702 ( .A(b[5]), .B(n[93]), .Z(n[220]) );
  GTECH_AND2 C703 ( .A(a[5]), .B(n[94]), .Z(n[158]) );
  GTECH_AND2 C704 ( .A(b[5]), .B(n[94]), .Z(n[221]) );
  GTECH_AND2 C705 ( .A(a[5]), .B(n[95]), .Z(n[159]) );
  GTECH_AND2 C706 ( .A(b[5]), .B(n[95]), .Z(n[222]) );
  GTECH_AND2 C707 ( .A(a[5]), .B(n[96]), .Z(n[160]) );
  GTECH_AND2 C708 ( .A(b[5]), .B(n[96]), .Z(n[223]) );
  GTECH_AND2 C709 ( .A(a[5]), .B(n[97]), .Z(n[161]) );
  GTECH_AND2 C710 ( .A(b[5]), .B(n[97]), .Z(n[224]) );
  GTECH_AND2 C711 ( .A(a[5]), .B(n[98]), .Z(n[162]) );
  GTECH_AND2 C712 ( .A(b[5]), .B(n[98]), .Z(n[225]) );
  GTECH_AND2 C713 ( .A(a[5]), .B(n[99]), .Z(n[163]) );
  GTECH_AND2 C714 ( .A(b[5]), .B(n[99]), .Z(n[226]) );
  GTECH_AND2 C715 ( .A(a[5]), .B(n[100]), .Z(n[164]) );
  GTECH_AND2 C716 ( .A(b[5]), .B(n[100]), .Z(n[227]) );
  GTECH_AND2 C717 ( .A(a[5]), .B(n[101]), .Z(n[165]) );
  GTECH_AND2 C718 ( .A(b[5]), .B(n[101]), .Z(n[228]) );
  GTECH_AND2 C719 ( .A(a[5]), .B(n[102]), .Z(n[166]) );
  GTECH_AND2 C720 ( .A(b[5]), .B(n[102]), .Z(n[229]) );
  GTECH_AND2 C721 ( .A(a[5]), .B(n[103]), .Z(n[167]) );
  GTECH_AND2 C722 ( .A(b[5]), .B(n[103]), .Z(n[230]) );
  GTECH_AND2 C723 ( .A(a[5]), .B(n[104]), .Z(n[168]) );
  GTECH_AND2 C724 ( .A(b[5]), .B(n[104]), .Z(n[231]) );
  GTECH_AND2 C725 ( .A(a[5]), .B(n[105]), .Z(n[169]) );
  GTECH_AND2 C726 ( .A(b[5]), .B(n[105]), .Z(n[232]) );
  GTECH_AND2 C727 ( .A(a[5]), .B(n[106]), .Z(n[170]) );
  GTECH_AND2 C728 ( .A(b[5]), .B(n[106]), .Z(n[233]) );
  GTECH_AND2 C729 ( .A(a[5]), .B(n[107]), .Z(n[171]) );
  GTECH_AND2 C730 ( .A(b[5]), .B(n[107]), .Z(n[234]) );
  GTECH_AND2 C731 ( .A(a[5]), .B(n[108]), .Z(n[172]) );
  GTECH_AND2 C732 ( .A(b[5]), .B(n[108]), .Z(n[235]) );
  GTECH_AND2 C733 ( .A(a[5]), .B(n[109]), .Z(n[173]) );
  GTECH_AND2 C734 ( .A(b[5]), .B(n[109]), .Z(n[236]) );
  GTECH_AND2 C735 ( .A(a[5]), .B(n[110]), .Z(n[174]) );
  GTECH_AND2 C736 ( .A(b[5]), .B(n[110]), .Z(n[237]) );
  GTECH_AND2 C737 ( .A(a[5]), .B(n[111]), .Z(n[175]) );
  GTECH_AND2 C738 ( .A(b[5]), .B(n[111]), .Z(n[238]) );
  GTECH_AND2 C739 ( .A(a[5]), .B(n[112]), .Z(n[176]) );
  GTECH_AND2 C740 ( .A(b[5]), .B(n[112]), .Z(n[239]) );
  GTECH_AND2 C741 ( .A(a[5]), .B(n[113]), .Z(n[177]) );
  GTECH_AND2 C742 ( .A(b[5]), .B(n[113]), .Z(n[240]) );
  GTECH_AND2 C743 ( .A(a[5]), .B(n[114]), .Z(n[178]) );
  GTECH_AND2 C744 ( .A(b[5]), .B(n[114]), .Z(n[241]) );
  GTECH_AND2 C745 ( .A(a[5]), .B(n[115]), .Z(n[179]) );
  GTECH_AND2 C746 ( .A(b[5]), .B(n[115]), .Z(n[242]) );
  GTECH_AND2 C747 ( .A(a[5]), .B(n[116]), .Z(n[180]) );
  GTECH_AND2 C748 ( .A(b[5]), .B(n[116]), .Z(n[243]) );
  GTECH_AND2 C749 ( .A(a[5]), .B(n[117]), .Z(n[181]) );
  GTECH_AND2 C750 ( .A(b[5]), .B(n[117]), .Z(n[244]) );
  GTECH_AND2 C751 ( .A(a[5]), .B(n[118]), .Z(n[182]) );
  GTECH_AND2 C752 ( .A(b[5]), .B(n[118]), .Z(n[245]) );
  GTECH_AND2 C753 ( .A(a[6]), .B(b[6]), .Z(n[246]) );
  GTECH_AND2 C754 ( .A(a[6]), .B(n[119]), .Z(n[247]) );
  GTECH_AND2 C755 ( .A(b[6]), .B(n[119]), .Z(n[374]) );
  GTECH_AND2 C756 ( .A(a[6]), .B(n[120]), .Z(n[248]) );
  GTECH_AND2 C757 ( .A(b[6]), .B(n[120]), .Z(n[375]) );
  GTECH_AND2 C758 ( .A(a[6]), .B(n[121]), .Z(n[249]) );
  GTECH_AND2 C759 ( .A(b[6]), .B(n[121]), .Z(n[376]) );
  GTECH_AND2 C760 ( .A(a[6]), .B(n[122]), .Z(n[250]) );
  GTECH_AND2 C761 ( .A(b[6]), .B(n[122]), .Z(n[377]) );
  GTECH_AND2 C762 ( .A(a[6]), .B(n[123]), .Z(n[251]) );
  GTECH_AND2 C763 ( .A(b[6]), .B(n[123]), .Z(n[378]) );
  GTECH_AND2 C764 ( .A(a[6]), .B(n[124]), .Z(n[252]) );
  GTECH_AND2 C765 ( .A(b[6]), .B(n[124]), .Z(n[379]) );
  GTECH_AND2 C766 ( .A(a[6]), .B(n[125]), .Z(n[253]) );
  GTECH_AND2 C767 ( .A(b[6]), .B(n[125]), .Z(n[380]) );
  GTECH_AND2 C768 ( .A(a[6]), .B(n[126]), .Z(n[254]) );
  GTECH_AND2 C769 ( .A(b[6]), .B(n[126]), .Z(n[381]) );
  GTECH_AND2 C770 ( .A(a[6]), .B(n[127]), .Z(n[255]) );
  GTECH_AND2 C771 ( .A(b[6]), .B(n[127]), .Z(n[382]) );
  GTECH_AND2 C772 ( .A(a[6]), .B(n[128]), .Z(n[256]) );
  GTECH_AND2 C773 ( .A(b[6]), .B(n[128]), .Z(n[383]) );
  GTECH_AND2 C774 ( .A(a[6]), .B(n[129]), .Z(n[257]) );
  GTECH_AND2 C775 ( .A(b[6]), .B(n[129]), .Z(n[384]) );
  GTECH_AND2 C776 ( .A(a[6]), .B(n[130]), .Z(n[258]) );
  GTECH_AND2 C777 ( .A(b[6]), .B(n[130]), .Z(n[385]) );
  GTECH_AND2 C778 ( .A(a[6]), .B(n[131]), .Z(n[259]) );
  GTECH_AND2 C779 ( .A(b[6]), .B(n[131]), .Z(n[386]) );
  GTECH_AND2 C780 ( .A(a[6]), .B(n[132]), .Z(n[260]) );
  GTECH_AND2 C781 ( .A(b[6]), .B(n[132]), .Z(n[387]) );
  GTECH_AND2 C782 ( .A(a[6]), .B(n[133]), .Z(n[261]) );
  GTECH_AND2 C783 ( .A(b[6]), .B(n[133]), .Z(n[388]) );
  GTECH_AND2 C784 ( .A(a[6]), .B(n[134]), .Z(n[262]) );
  GTECH_AND2 C785 ( .A(b[6]), .B(n[134]), .Z(n[389]) );
  GTECH_AND2 C786 ( .A(a[6]), .B(n[135]), .Z(n[263]) );
  GTECH_AND2 C787 ( .A(b[6]), .B(n[135]), .Z(n[390]) );
  GTECH_AND2 C788 ( .A(a[6]), .B(n[136]), .Z(n[264]) );
  GTECH_AND2 C789 ( .A(b[6]), .B(n[136]), .Z(n[391]) );
  GTECH_AND2 C790 ( .A(a[6]), .B(n[137]), .Z(n[265]) );
  GTECH_AND2 C791 ( .A(b[6]), .B(n[137]), .Z(n[392]) );
  GTECH_AND2 C792 ( .A(a[6]), .B(n[138]), .Z(n[266]) );
  GTECH_AND2 C793 ( .A(b[6]), .B(n[138]), .Z(n[393]) );
  GTECH_AND2 C794 ( .A(a[6]), .B(n[139]), .Z(n[267]) );
  GTECH_AND2 C795 ( .A(b[6]), .B(n[139]), .Z(n[394]) );
  GTECH_AND2 C796 ( .A(a[6]), .B(n[140]), .Z(n[268]) );
  GTECH_AND2 C797 ( .A(b[6]), .B(n[140]), .Z(n[395]) );
  GTECH_AND2 C798 ( .A(a[6]), .B(n[141]), .Z(n[269]) );
  GTECH_AND2 C799 ( .A(b[6]), .B(n[141]), .Z(n[396]) );
  GTECH_AND2 C800 ( .A(a[6]), .B(n[142]), .Z(n[270]) );
  GTECH_AND2 C801 ( .A(b[6]), .B(n[142]), .Z(n[397]) );
  GTECH_AND2 C802 ( .A(a[6]), .B(n[143]), .Z(n[271]) );
  GTECH_AND2 C803 ( .A(b[6]), .B(n[143]), .Z(n[398]) );
  GTECH_AND2 C804 ( .A(a[6]), .B(n[144]), .Z(n[272]) );
  GTECH_AND2 C805 ( .A(b[6]), .B(n[144]), .Z(n[399]) );
  GTECH_AND2 C806 ( .A(a[6]), .B(n[145]), .Z(n[273]) );
  GTECH_AND2 C807 ( .A(b[6]), .B(n[145]), .Z(n[400]) );
  GTECH_AND2 C808 ( .A(a[6]), .B(n[146]), .Z(n[274]) );
  GTECH_AND2 C809 ( .A(b[6]), .B(n[146]), .Z(n[401]) );
  GTECH_AND2 C810 ( .A(a[6]), .B(n[147]), .Z(n[275]) );
  GTECH_AND2 C811 ( .A(b[6]), .B(n[147]), .Z(n[402]) );
  GTECH_AND2 C812 ( .A(a[6]), .B(n[148]), .Z(n[276]) );
  GTECH_AND2 C813 ( .A(b[6]), .B(n[148]), .Z(n[403]) );
  GTECH_AND2 C814 ( .A(a[6]), .B(n[149]), .Z(n[277]) );
  GTECH_AND2 C815 ( .A(b[6]), .B(n[149]), .Z(n[404]) );
  GTECH_AND2 C816 ( .A(a[6]), .B(n[150]), .Z(n[278]) );
  GTECH_AND2 C817 ( .A(b[6]), .B(n[150]), .Z(n[405]) );
  GTECH_AND2 C818 ( .A(a[6]), .B(n[151]), .Z(n[279]) );
  GTECH_AND2 C819 ( .A(b[6]), .B(n[151]), .Z(n[406]) );
  GTECH_AND2 C820 ( .A(a[6]), .B(n[152]), .Z(n[280]) );
  GTECH_AND2 C821 ( .A(b[6]), .B(n[152]), .Z(n[407]) );
  GTECH_AND2 C822 ( .A(a[6]), .B(n[153]), .Z(n[281]) );
  GTECH_AND2 C823 ( .A(b[6]), .B(n[153]), .Z(n[408]) );
  GTECH_AND2 C824 ( .A(a[6]), .B(n[154]), .Z(n[282]) );
  GTECH_AND2 C825 ( .A(b[6]), .B(n[154]), .Z(n[409]) );
  GTECH_AND2 C826 ( .A(a[6]), .B(n[155]), .Z(n[283]) );
  GTECH_AND2 C827 ( .A(b[6]), .B(n[155]), .Z(n[410]) );
  GTECH_AND2 C828 ( .A(a[6]), .B(n[156]), .Z(n[284]) );
  GTECH_AND2 C829 ( .A(b[6]), .B(n[156]), .Z(n[411]) );
  GTECH_AND2 C830 ( .A(a[6]), .B(n[157]), .Z(n[285]) );
  GTECH_AND2 C831 ( .A(b[6]), .B(n[157]), .Z(n[412]) );
  GTECH_AND2 C832 ( .A(a[6]), .B(n[158]), .Z(n[286]) );
  GTECH_AND2 C833 ( .A(b[6]), .B(n[158]), .Z(n[413]) );
  GTECH_AND2 C834 ( .A(a[6]), .B(n[159]), .Z(n[287]) );
  GTECH_AND2 C835 ( .A(b[6]), .B(n[159]), .Z(n[414]) );
  GTECH_AND2 C836 ( .A(a[6]), .B(n[160]), .Z(n[288]) );
  GTECH_AND2 C837 ( .A(b[6]), .B(n[160]), .Z(n[415]) );
  GTECH_AND2 C838 ( .A(a[6]), .B(n[161]), .Z(n[289]) );
  GTECH_AND2 C839 ( .A(b[6]), .B(n[161]), .Z(n[416]) );
  GTECH_AND2 C840 ( .A(a[6]), .B(n[162]), .Z(n[290]) );
  GTECH_AND2 C841 ( .A(b[6]), .B(n[162]), .Z(n[417]) );
  GTECH_AND2 C842 ( .A(a[6]), .B(n[163]), .Z(n[291]) );
  GTECH_AND2 C843 ( .A(b[6]), .B(n[163]), .Z(n[418]) );
  GTECH_AND2 C844 ( .A(a[6]), .B(n[164]), .Z(n[292]) );
  GTECH_AND2 C845 ( .A(b[6]), .B(n[164]), .Z(n[419]) );
  GTECH_AND2 C846 ( .A(a[6]), .B(n[165]), .Z(n[293]) );
  GTECH_AND2 C847 ( .A(b[6]), .B(n[165]), .Z(n[420]) );
  GTECH_AND2 C848 ( .A(a[6]), .B(n[166]), .Z(n[294]) );
  GTECH_AND2 C849 ( .A(b[6]), .B(n[166]), .Z(n[421]) );
  GTECH_AND2 C850 ( .A(a[6]), .B(n[167]), .Z(n[295]) );
  GTECH_AND2 C851 ( .A(b[6]), .B(n[167]), .Z(n[422]) );
  GTECH_AND2 C852 ( .A(a[6]), .B(n[168]), .Z(n[296]) );
  GTECH_AND2 C853 ( .A(b[6]), .B(n[168]), .Z(n[423]) );
  GTECH_AND2 C854 ( .A(a[6]), .B(n[169]), .Z(n[297]) );
  GTECH_AND2 C855 ( .A(b[6]), .B(n[169]), .Z(n[424]) );
  GTECH_AND2 C856 ( .A(a[6]), .B(n[170]), .Z(n[298]) );
  GTECH_AND2 C857 ( .A(b[6]), .B(n[170]), .Z(n[425]) );
  GTECH_AND2 C858 ( .A(a[6]), .B(n[171]), .Z(n[299]) );
  GTECH_AND2 C859 ( .A(b[6]), .B(n[171]), .Z(n[426]) );
  GTECH_AND2 C860 ( .A(a[6]), .B(n[172]), .Z(n[300]) );
  GTECH_AND2 C861 ( .A(b[6]), .B(n[172]), .Z(n[427]) );
  GTECH_AND2 C862 ( .A(a[6]), .B(n[173]), .Z(n[301]) );
  GTECH_AND2 C863 ( .A(b[6]), .B(n[173]), .Z(n[428]) );
  GTECH_AND2 C864 ( .A(a[6]), .B(n[174]), .Z(n[302]) );
  GTECH_AND2 C865 ( .A(b[6]), .B(n[174]), .Z(n[429]) );
  GTECH_AND2 C866 ( .A(a[6]), .B(n[175]), .Z(n[303]) );
  GTECH_AND2 C867 ( .A(b[6]), .B(n[175]), .Z(n[430]) );
  GTECH_AND2 C868 ( .A(a[6]), .B(n[176]), .Z(n[304]) );
  GTECH_AND2 C869 ( .A(b[6]), .B(n[176]), .Z(n[431]) );
  GTECH_AND2 C870 ( .A(a[6]), .B(n[177]), .Z(n[305]) );
  GTECH_AND2 C871 ( .A(b[6]), .B(n[177]), .Z(n[432]) );
  GTECH_AND2 C872 ( .A(a[6]), .B(n[178]), .Z(n[306]) );
  GTECH_AND2 C873 ( .A(b[6]), .B(n[178]), .Z(n[433]) );
  GTECH_AND2 C874 ( .A(a[6]), .B(n[179]), .Z(n[307]) );
  GTECH_AND2 C875 ( .A(b[6]), .B(n[179]), .Z(n[434]) );
  GTECH_AND2 C876 ( .A(a[6]), .B(n[180]), .Z(n[308]) );
  GTECH_AND2 C877 ( .A(b[6]), .B(n[180]), .Z(n[435]) );
  GTECH_AND2 C878 ( .A(a[6]), .B(n[181]), .Z(n[309]) );
  GTECH_AND2 C879 ( .A(b[6]), .B(n[181]), .Z(n[436]) );
  GTECH_AND2 C880 ( .A(a[6]), .B(n[182]), .Z(n[310]) );
  GTECH_AND2 C881 ( .A(b[6]), .B(n[182]), .Z(n[437]) );
  GTECH_AND2 C882 ( .A(a[6]), .B(n[183]), .Z(n[311]) );
  GTECH_AND2 C883 ( .A(b[6]), .B(n[183]), .Z(n[438]) );
  GTECH_AND2 C884 ( .A(a[6]), .B(n[184]), .Z(n[312]) );
  GTECH_AND2 C885 ( .A(b[6]), .B(n[184]), .Z(n[439]) );
  GTECH_AND2 C886 ( .A(a[6]), .B(n[185]), .Z(n[313]) );
  GTECH_AND2 C887 ( .A(b[6]), .B(n[185]), .Z(n[440]) );
  GTECH_AND2 C888 ( .A(a[6]), .B(n[186]), .Z(n[314]) );
  GTECH_AND2 C889 ( .A(b[6]), .B(n[186]), .Z(n[441]) );
  GTECH_AND2 C890 ( .A(a[6]), .B(n[187]), .Z(n[315]) );
  GTECH_AND2 C891 ( .A(b[6]), .B(n[187]), .Z(n[442]) );
  GTECH_AND2 C892 ( .A(a[6]), .B(n[188]), .Z(n[316]) );
  GTECH_AND2 C893 ( .A(b[6]), .B(n[188]), .Z(n[443]) );
  GTECH_AND2 C894 ( .A(a[6]), .B(n[189]), .Z(n[317]) );
  GTECH_AND2 C895 ( .A(b[6]), .B(n[189]), .Z(n[444]) );
  GTECH_AND2 C896 ( .A(a[6]), .B(n[190]), .Z(n[318]) );
  GTECH_AND2 C897 ( .A(b[6]), .B(n[190]), .Z(n[445]) );
  GTECH_AND2 C898 ( .A(a[6]), .B(n[191]), .Z(n[319]) );
  GTECH_AND2 C899 ( .A(b[6]), .B(n[191]), .Z(n[446]) );
  GTECH_AND2 C900 ( .A(a[6]), .B(n[192]), .Z(n[320]) );
  GTECH_AND2 C901 ( .A(b[6]), .B(n[192]), .Z(n[447]) );
  GTECH_AND2 C902 ( .A(a[6]), .B(n[193]), .Z(n[321]) );
  GTECH_AND2 C903 ( .A(b[6]), .B(n[193]), .Z(n[448]) );
  GTECH_AND2 C904 ( .A(a[6]), .B(n[194]), .Z(n[322]) );
  GTECH_AND2 C905 ( .A(b[6]), .B(n[194]), .Z(n[449]) );
  GTECH_AND2 C906 ( .A(a[6]), .B(n[195]), .Z(n[323]) );
  GTECH_AND2 C907 ( .A(b[6]), .B(n[195]), .Z(n[450]) );
  GTECH_AND2 C908 ( .A(a[6]), .B(n[196]), .Z(n[324]) );
  GTECH_AND2 C909 ( .A(b[6]), .B(n[196]), .Z(n[451]) );
  GTECH_AND2 C910 ( .A(a[6]), .B(n[197]), .Z(n[325]) );
  GTECH_AND2 C911 ( .A(b[6]), .B(n[197]), .Z(n[452]) );
  GTECH_AND2 C912 ( .A(a[6]), .B(n[198]), .Z(n[326]) );
  GTECH_AND2 C913 ( .A(b[6]), .B(n[198]), .Z(n[453]) );
  GTECH_AND2 C914 ( .A(a[6]), .B(n[199]), .Z(n[327]) );
  GTECH_AND2 C915 ( .A(b[6]), .B(n[199]), .Z(n[454]) );
  GTECH_AND2 C916 ( .A(a[6]), .B(n[200]), .Z(n[328]) );
  GTECH_AND2 C917 ( .A(b[6]), .B(n[200]), .Z(n[455]) );
  GTECH_AND2 C918 ( .A(a[6]), .B(n[201]), .Z(n[329]) );
  GTECH_AND2 C919 ( .A(b[6]), .B(n[201]), .Z(n[456]) );
  GTECH_AND2 C920 ( .A(a[6]), .B(n[202]), .Z(n[330]) );
  GTECH_AND2 C921 ( .A(b[6]), .B(n[202]), .Z(n[457]) );
  GTECH_AND2 C922 ( .A(a[6]), .B(n[203]), .Z(n[331]) );
  GTECH_AND2 C923 ( .A(b[6]), .B(n[203]), .Z(n[458]) );
  GTECH_AND2 C924 ( .A(a[6]), .B(n[204]), .Z(n[332]) );
  GTECH_AND2 C925 ( .A(b[6]), .B(n[204]), .Z(n[459]) );
  GTECH_AND2 C926 ( .A(a[6]), .B(n[205]), .Z(n[333]) );
  GTECH_AND2 C927 ( .A(b[6]), .B(n[205]), .Z(n[460]) );
  GTECH_AND2 C928 ( .A(a[6]), .B(n[206]), .Z(n[334]) );
  GTECH_AND2 C929 ( .A(b[6]), .B(n[206]), .Z(n[461]) );
  GTECH_AND2 C930 ( .A(a[6]), .B(n[207]), .Z(n[335]) );
  GTECH_AND2 C931 ( .A(b[6]), .B(n[207]), .Z(n[462]) );
  GTECH_AND2 C932 ( .A(a[6]), .B(n[208]), .Z(n[336]) );
  GTECH_AND2 C933 ( .A(b[6]), .B(n[208]), .Z(n[463]) );
  GTECH_AND2 C934 ( .A(a[6]), .B(n[209]), .Z(n[337]) );
  GTECH_AND2 C935 ( .A(b[6]), .B(n[209]), .Z(n[464]) );
  GTECH_AND2 C936 ( .A(a[6]), .B(n[210]), .Z(n[338]) );
  GTECH_AND2 C937 ( .A(b[6]), .B(n[210]), .Z(n[465]) );
  GTECH_AND2 C938 ( .A(a[6]), .B(n[211]), .Z(n[339]) );
  GTECH_AND2 C939 ( .A(b[6]), .B(n[211]), .Z(n[466]) );
  GTECH_AND2 C940 ( .A(a[6]), .B(n[212]), .Z(n[340]) );
  GTECH_AND2 C941 ( .A(b[6]), .B(n[212]), .Z(n[467]) );
  GTECH_AND2 C942 ( .A(a[6]), .B(n[213]), .Z(n[341]) );
  GTECH_AND2 C943 ( .A(b[6]), .B(n[213]), .Z(n[468]) );
  GTECH_AND2 C944 ( .A(a[6]), .B(n[214]), .Z(n[342]) );
  GTECH_AND2 C945 ( .A(b[6]), .B(n[214]), .Z(n[469]) );
  GTECH_AND2 C946 ( .A(a[6]), .B(n[215]), .Z(n[343]) );
  GTECH_AND2 C947 ( .A(b[6]), .B(n[215]), .Z(n[470]) );
  GTECH_AND2 C948 ( .A(a[6]), .B(n[216]), .Z(n[344]) );
  GTECH_AND2 C949 ( .A(b[6]), .B(n[216]), .Z(n[471]) );
  GTECH_AND2 C950 ( .A(a[6]), .B(n[217]), .Z(n[345]) );
  GTECH_AND2 C951 ( .A(b[6]), .B(n[217]), .Z(n[472]) );
  GTECH_AND2 C952 ( .A(a[6]), .B(n[218]), .Z(n[346]) );
  GTECH_AND2 C953 ( .A(b[6]), .B(n[218]), .Z(n[473]) );
  GTECH_AND2 C954 ( .A(a[6]), .B(n[219]), .Z(n[347]) );
  GTECH_AND2 C955 ( .A(b[6]), .B(n[219]), .Z(n[474]) );
  GTECH_AND2 C956 ( .A(a[6]), .B(n[220]), .Z(n[348]) );
  GTECH_AND2 C957 ( .A(b[6]), .B(n[220]), .Z(n[475]) );
  GTECH_AND2 C958 ( .A(a[6]), .B(n[221]), .Z(n[349]) );
  GTECH_AND2 C959 ( .A(b[6]), .B(n[221]), .Z(n[476]) );
  GTECH_AND2 C960 ( .A(a[6]), .B(n[222]), .Z(n[350]) );
  GTECH_AND2 C961 ( .A(b[6]), .B(n[222]), .Z(n[477]) );
  GTECH_AND2 C962 ( .A(a[6]), .B(n[223]), .Z(n[351]) );
  GTECH_AND2 C963 ( .A(b[6]), .B(n[223]), .Z(n[478]) );
  GTECH_AND2 C964 ( .A(a[6]), .B(n[224]), .Z(n[352]) );
  GTECH_AND2 C965 ( .A(b[6]), .B(n[224]), .Z(n[479]) );
  GTECH_AND2 C966 ( .A(a[6]), .B(n[225]), .Z(n[353]) );
  GTECH_AND2 C967 ( .A(b[6]), .B(n[225]), .Z(n[480]) );
  GTECH_AND2 C968 ( .A(a[6]), .B(n[226]), .Z(n[354]) );
  GTECH_AND2 C969 ( .A(b[6]), .B(n[226]), .Z(n[481]) );
  GTECH_AND2 C970 ( .A(a[6]), .B(n[227]), .Z(n[355]) );
  GTECH_AND2 C971 ( .A(b[6]), .B(n[227]), .Z(n[482]) );
  GTECH_AND2 C972 ( .A(a[6]), .B(n[228]), .Z(n[356]) );
  GTECH_AND2 C973 ( .A(b[6]), .B(n[228]), .Z(n[483]) );
  GTECH_AND2 C974 ( .A(a[6]), .B(n[229]), .Z(n[357]) );
  GTECH_AND2 C975 ( .A(b[6]), .B(n[229]), .Z(n[484]) );
  GTECH_AND2 C976 ( .A(a[6]), .B(n[230]), .Z(n[358]) );
  GTECH_AND2 C977 ( .A(b[6]), .B(n[230]), .Z(n[485]) );
  GTECH_AND2 C978 ( .A(a[6]), .B(n[231]), .Z(n[359]) );
  GTECH_AND2 C979 ( .A(b[6]), .B(n[231]), .Z(n[486]) );
  GTECH_AND2 C980 ( .A(a[6]), .B(n[232]), .Z(n[360]) );
  GTECH_AND2 C981 ( .A(b[6]), .B(n[232]), .Z(n[487]) );
  GTECH_AND2 C982 ( .A(a[6]), .B(n[233]), .Z(n[361]) );
  GTECH_AND2 C983 ( .A(b[6]), .B(n[233]), .Z(n[488]) );
  GTECH_AND2 C984 ( .A(a[6]), .B(n[234]), .Z(n[362]) );
  GTECH_AND2 C985 ( .A(b[6]), .B(n[234]), .Z(n[489]) );
  GTECH_AND2 C986 ( .A(a[6]), .B(n[235]), .Z(n[363]) );
  GTECH_AND2 C987 ( .A(b[6]), .B(n[235]), .Z(n[490]) );
  GTECH_AND2 C988 ( .A(a[6]), .B(n[236]), .Z(n[364]) );
  GTECH_AND2 C989 ( .A(b[6]), .B(n[236]), .Z(n[491]) );
  GTECH_AND2 C990 ( .A(a[6]), .B(n[237]), .Z(n[365]) );
  GTECH_AND2 C991 ( .A(b[6]), .B(n[237]), .Z(n[492]) );
  GTECH_AND2 C992 ( .A(a[6]), .B(n[238]), .Z(n[366]) );
  GTECH_AND2 C993 ( .A(b[6]), .B(n[238]), .Z(n[493]) );
  GTECH_AND2 C994 ( .A(a[6]), .B(n[239]), .Z(n[367]) );
  GTECH_AND2 C995 ( .A(b[6]), .B(n[239]), .Z(n[494]) );
  GTECH_AND2 C996 ( .A(a[6]), .B(n[240]), .Z(n[368]) );
  GTECH_AND2 C997 ( .A(b[6]), .B(n[240]), .Z(n[495]) );
  GTECH_AND2 C998 ( .A(a[6]), .B(n[241]), .Z(n[369]) );
  GTECH_AND2 C999 ( .A(b[6]), .B(n[241]), .Z(n[496]) );
  GTECH_AND2 C1000 ( .A(a[6]), .B(n[242]), .Z(n[370]) );
  GTECH_AND2 C1001 ( .A(b[6]), .B(n[242]), .Z(n[497]) );
  GTECH_AND2 C1002 ( .A(a[6]), .B(n[243]), .Z(n[371]) );
  GTECH_AND2 C1003 ( .A(b[6]), .B(n[243]), .Z(n[498]) );
  GTECH_AND2 C1004 ( .A(a[6]), .B(n[244]), .Z(n[372]) );
  GTECH_AND2 C1005 ( .A(b[6]), .B(n[244]), .Z(n[499]) );
  GTECH_AND2 C1006 ( .A(a[6]), .B(n[245]), .Z(n[373]) );
  GTECH_AND2 C1007 ( .A(b[6]), .B(n[245]), .Z(n[500]) );
endmodule


module adder_cpe ( a, b, code );
  input [6:0] a;
  input [6:0] b;
  output [14:0] code;

  wire   [500:0] nonlin;
  wire   [7:0] sum;

  gen_nonlinear_part NONLIN_ADDER ( .a(a), .b(b), .c(1'b0), .n(nonlin) );
  gen_linear_part LIN_ADDER ( .a(a), .b(b), .c_in(1'b0), .n(nonlin), .s(sum)
         );
  generator CPE ( .i(sum[6:0]), .c(code) );
endmodule

