module pearson();

endmodule
