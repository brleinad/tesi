library verilog;
use verilog.vl_types.all;
entity tb_RM is
end tb_RM;
