
module cla_adder ( a, b, s, cin, cout );
  input [511:0] a;
  input [511:0] b;
  output [511:0] s;
  input cin;
  output cout;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242,
         N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253,
         N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264,
         N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374,
         N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N385,
         N386, N387, N388, N389, N390, N391, N392, N393, N394, N395, N396,
         N397, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440,
         N441, N442, N443, N444, N445, N446, N447, N448, N449, N450, N451,
         N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, N462,
         N463, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N496, N497, N498, N499, N500, N501, N502, N503, N504, N505, N506,
         N507, N508, N509, N510;
  wire   [510:0] g;
  wire   [511:0] p;
  wire   [511:1] c;

  XOR2D0 C4610 ( .A1(p[0]), .A2(cin), .Z(s[0]) );
  XOR2D0 C4609 ( .A1(p[1]), .A2(c[1]), .Z(s[1]) );
  XOR2D0 C4608 ( .A1(p[2]), .A2(c[2]), .Z(s[2]) );
  XOR2D0 C4607 ( .A1(p[3]), .A2(c[3]), .Z(s[3]) );
  XOR2D0 C4606 ( .A1(p[4]), .A2(c[4]), .Z(s[4]) );
  XOR2D0 C4605 ( .A1(p[5]), .A2(c[5]), .Z(s[5]) );
  XOR2D0 C4604 ( .A1(p[6]), .A2(c[6]), .Z(s[6]) );
  XOR2D0 C4603 ( .A1(p[7]), .A2(c[7]), .Z(s[7]) );
  XOR2D0 C4602 ( .A1(p[8]), .A2(c[8]), .Z(s[8]) );
  XOR2D0 C4601 ( .A1(p[9]), .A2(c[9]), .Z(s[9]) );
  XOR2D0 C4600 ( .A1(p[10]), .A2(c[10]), .Z(s[10]) );
  XOR2D0 C4599 ( .A1(p[11]), .A2(c[11]), .Z(s[11]) );
  XOR2D0 C4598 ( .A1(p[12]), .A2(c[12]), .Z(s[12]) );
  XOR2D0 C4597 ( .A1(p[13]), .A2(c[13]), .Z(s[13]) );
  XOR2D0 C4596 ( .A1(p[14]), .A2(c[14]), .Z(s[14]) );
  XOR2D0 C4595 ( .A1(p[15]), .A2(c[15]), .Z(s[15]) );
  XOR2D0 C4594 ( .A1(p[16]), .A2(c[16]), .Z(s[16]) );
  XOR2D0 C4593 ( .A1(p[17]), .A2(c[17]), .Z(s[17]) );
  XOR2D0 C4592 ( .A1(p[18]), .A2(c[18]), .Z(s[18]) );
  XOR2D0 C4591 ( .A1(p[19]), .A2(c[19]), .Z(s[19]) );
  XOR2D0 C4590 ( .A1(p[20]), .A2(c[20]), .Z(s[20]) );
  XOR2D0 C4589 ( .A1(p[21]), .A2(c[21]), .Z(s[21]) );
  XOR2D0 C4588 ( .A1(p[22]), .A2(c[22]), .Z(s[22]) );
  XOR2D0 C4587 ( .A1(p[23]), .A2(c[23]), .Z(s[23]) );
  XOR2D0 C4586 ( .A1(p[24]), .A2(c[24]), .Z(s[24]) );
  XOR2D0 C4585 ( .A1(p[25]), .A2(c[25]), .Z(s[25]) );
  XOR2D0 C4584 ( .A1(p[26]), .A2(c[26]), .Z(s[26]) );
  XOR2D0 C4583 ( .A1(p[27]), .A2(c[27]), .Z(s[27]) );
  XOR2D0 C4582 ( .A1(p[28]), .A2(c[28]), .Z(s[28]) );
  XOR2D0 C4581 ( .A1(p[29]), .A2(c[29]), .Z(s[29]) );
  XOR2D0 C4580 ( .A1(p[30]), .A2(c[30]), .Z(s[30]) );
  XOR2D0 C4579 ( .A1(p[31]), .A2(c[31]), .Z(s[31]) );
  XOR2D0 C4578 ( .A1(p[32]), .A2(c[32]), .Z(s[32]) );
  XOR2D0 C4577 ( .A1(p[33]), .A2(c[33]), .Z(s[33]) );
  XOR2D0 C4576 ( .A1(p[34]), .A2(c[34]), .Z(s[34]) );
  XOR2D0 C4575 ( .A1(p[35]), .A2(c[35]), .Z(s[35]) );
  XOR2D0 C4574 ( .A1(p[36]), .A2(c[36]), .Z(s[36]) );
  XOR2D0 C4573 ( .A1(p[37]), .A2(c[37]), .Z(s[37]) );
  XOR2D0 C4572 ( .A1(p[38]), .A2(c[38]), .Z(s[38]) );
  XOR2D0 C4571 ( .A1(p[39]), .A2(c[39]), .Z(s[39]) );
  XOR2D0 C4570 ( .A1(p[40]), .A2(c[40]), .Z(s[40]) );
  XOR2D0 C4569 ( .A1(p[41]), .A2(c[41]), .Z(s[41]) );
  XOR2D0 C4568 ( .A1(p[42]), .A2(c[42]), .Z(s[42]) );
  XOR2D0 C4567 ( .A1(p[43]), .A2(c[43]), .Z(s[43]) );
  XOR2D0 C4566 ( .A1(p[44]), .A2(c[44]), .Z(s[44]) );
  XOR2D0 C4565 ( .A1(p[45]), .A2(c[45]), .Z(s[45]) );
  XOR2D0 C4564 ( .A1(p[46]), .A2(c[46]), .Z(s[46]) );
  XOR2D0 C4563 ( .A1(p[47]), .A2(c[47]), .Z(s[47]) );
  XOR2D0 C4562 ( .A1(p[48]), .A2(c[48]), .Z(s[48]) );
  XOR2D0 C4561 ( .A1(p[49]), .A2(c[49]), .Z(s[49]) );
  XOR2D0 C4560 ( .A1(p[50]), .A2(c[50]), .Z(s[50]) );
  XOR2D0 C4559 ( .A1(p[51]), .A2(c[51]), .Z(s[51]) );
  XOR2D0 C4558 ( .A1(p[52]), .A2(c[52]), .Z(s[52]) );
  XOR2D0 C4557 ( .A1(p[53]), .A2(c[53]), .Z(s[53]) );
  XOR2D0 C4556 ( .A1(p[54]), .A2(c[54]), .Z(s[54]) );
  XOR2D0 C4555 ( .A1(p[55]), .A2(c[55]), .Z(s[55]) );
  XOR2D0 C4554 ( .A1(p[56]), .A2(c[56]), .Z(s[56]) );
  XOR2D0 C4553 ( .A1(p[57]), .A2(c[57]), .Z(s[57]) );
  XOR2D0 C4552 ( .A1(p[58]), .A2(c[58]), .Z(s[58]) );
  XOR2D0 C4551 ( .A1(p[59]), .A2(c[59]), .Z(s[59]) );
  XOR2D0 C4550 ( .A1(p[60]), .A2(c[60]), .Z(s[60]) );
  XOR2D0 C4549 ( .A1(p[61]), .A2(c[61]), .Z(s[61]) );
  XOR2D0 C4548 ( .A1(p[62]), .A2(c[62]), .Z(s[62]) );
  XOR2D0 C4547 ( .A1(p[63]), .A2(c[63]), .Z(s[63]) );
  XOR2D0 C4546 ( .A1(p[64]), .A2(c[64]), .Z(s[64]) );
  XOR2D0 C4545 ( .A1(p[65]), .A2(c[65]), .Z(s[65]) );
  XOR2D0 C4544 ( .A1(p[66]), .A2(c[66]), .Z(s[66]) );
  XOR2D0 C4543 ( .A1(p[67]), .A2(c[67]), .Z(s[67]) );
  XOR2D0 C4542 ( .A1(p[68]), .A2(c[68]), .Z(s[68]) );
  XOR2D0 C4541 ( .A1(p[69]), .A2(c[69]), .Z(s[69]) );
  XOR2D0 C4540 ( .A1(p[70]), .A2(c[70]), .Z(s[70]) );
  XOR2D0 C4539 ( .A1(p[71]), .A2(c[71]), .Z(s[71]) );
  XOR2D0 C4538 ( .A1(p[72]), .A2(c[72]), .Z(s[72]) );
  XOR2D0 C4537 ( .A1(p[73]), .A2(c[73]), .Z(s[73]) );
  XOR2D0 C4536 ( .A1(p[74]), .A2(c[74]), .Z(s[74]) );
  XOR2D0 C4535 ( .A1(p[75]), .A2(c[75]), .Z(s[75]) );
  XOR2D0 C4534 ( .A1(p[76]), .A2(c[76]), .Z(s[76]) );
  XOR2D0 C4533 ( .A1(p[77]), .A2(c[77]), .Z(s[77]) );
  XOR2D0 C4532 ( .A1(p[78]), .A2(c[78]), .Z(s[78]) );
  XOR2D0 C4531 ( .A1(p[79]), .A2(c[79]), .Z(s[79]) );
  XOR2D0 C4530 ( .A1(p[80]), .A2(c[80]), .Z(s[80]) );
  XOR2D0 C4529 ( .A1(p[81]), .A2(c[81]), .Z(s[81]) );
  XOR2D0 C4528 ( .A1(p[82]), .A2(c[82]), .Z(s[82]) );
  XOR2D0 C4527 ( .A1(p[83]), .A2(c[83]), .Z(s[83]) );
  XOR2D0 C4526 ( .A1(p[84]), .A2(c[84]), .Z(s[84]) );
  XOR2D0 C4525 ( .A1(p[85]), .A2(c[85]), .Z(s[85]) );
  XOR2D0 C4524 ( .A1(p[86]), .A2(c[86]), .Z(s[86]) );
  XOR2D0 C4523 ( .A1(p[87]), .A2(c[87]), .Z(s[87]) );
  XOR2D0 C4522 ( .A1(p[88]), .A2(c[88]), .Z(s[88]) );
  XOR2D0 C4521 ( .A1(p[89]), .A2(c[89]), .Z(s[89]) );
  XOR2D0 C4520 ( .A1(p[90]), .A2(c[90]), .Z(s[90]) );
  XOR2D0 C4519 ( .A1(p[91]), .A2(c[91]), .Z(s[91]) );
  XOR2D0 C4518 ( .A1(p[92]), .A2(c[92]), .Z(s[92]) );
  XOR2D0 C4517 ( .A1(p[93]), .A2(c[93]), .Z(s[93]) );
  XOR2D0 C4516 ( .A1(p[94]), .A2(c[94]), .Z(s[94]) );
  XOR2D0 C4515 ( .A1(p[95]), .A2(c[95]), .Z(s[95]) );
  XOR2D0 C4514 ( .A1(p[96]), .A2(c[96]), .Z(s[96]) );
  XOR2D0 C4513 ( .A1(p[97]), .A2(c[97]), .Z(s[97]) );
  XOR2D0 C4512 ( .A1(p[98]), .A2(c[98]), .Z(s[98]) );
  XOR2D0 C4511 ( .A1(p[99]), .A2(c[99]), .Z(s[99]) );
  XOR2D0 C4510 ( .A1(p[100]), .A2(c[100]), .Z(s[100]) );
  XOR2D0 C4509 ( .A1(p[101]), .A2(c[101]), .Z(s[101]) );
  XOR2D0 C4508 ( .A1(p[102]), .A2(c[102]), .Z(s[102]) );
  XOR2D0 C4507 ( .A1(p[103]), .A2(c[103]), .Z(s[103]) );
  XOR2D0 C4506 ( .A1(p[104]), .A2(c[104]), .Z(s[104]) );
  XOR2D0 C4505 ( .A1(p[105]), .A2(c[105]), .Z(s[105]) );
  XOR2D0 C4504 ( .A1(p[106]), .A2(c[106]), .Z(s[106]) );
  XOR2D0 C4503 ( .A1(p[107]), .A2(c[107]), .Z(s[107]) );
  XOR2D0 C4502 ( .A1(p[108]), .A2(c[108]), .Z(s[108]) );
  XOR2D0 C4501 ( .A1(p[109]), .A2(c[109]), .Z(s[109]) );
  XOR2D0 C4500 ( .A1(p[110]), .A2(c[110]), .Z(s[110]) );
  XOR2D0 C4499 ( .A1(p[111]), .A2(c[111]), .Z(s[111]) );
  XOR2D0 C4498 ( .A1(p[112]), .A2(c[112]), .Z(s[112]) );
  XOR2D0 C4497 ( .A1(p[113]), .A2(c[113]), .Z(s[113]) );
  XOR2D0 C4496 ( .A1(p[114]), .A2(c[114]), .Z(s[114]) );
  XOR2D0 C4495 ( .A1(p[115]), .A2(c[115]), .Z(s[115]) );
  XOR2D0 C4494 ( .A1(p[116]), .A2(c[116]), .Z(s[116]) );
  XOR2D0 C4493 ( .A1(p[117]), .A2(c[117]), .Z(s[117]) );
  XOR2D0 C4492 ( .A1(p[118]), .A2(c[118]), .Z(s[118]) );
  XOR2D0 C4491 ( .A1(p[119]), .A2(c[119]), .Z(s[119]) );
  XOR2D0 C4490 ( .A1(p[120]), .A2(c[120]), .Z(s[120]) );
  XOR2D0 C4489 ( .A1(p[121]), .A2(c[121]), .Z(s[121]) );
  XOR2D0 C4488 ( .A1(p[122]), .A2(c[122]), .Z(s[122]) );
  XOR2D0 C4487 ( .A1(p[123]), .A2(c[123]), .Z(s[123]) );
  XOR2D0 C4486 ( .A1(p[124]), .A2(c[124]), .Z(s[124]) );
  XOR2D0 C4485 ( .A1(p[125]), .A2(c[125]), .Z(s[125]) );
  XOR2D0 C4484 ( .A1(p[126]), .A2(c[126]), .Z(s[126]) );
  XOR2D0 C4483 ( .A1(p[127]), .A2(c[127]), .Z(s[127]) );
  XOR2D0 C4482 ( .A1(p[128]), .A2(c[128]), .Z(s[128]) );
  XOR2D0 C4481 ( .A1(p[129]), .A2(c[129]), .Z(s[129]) );
  XOR2D0 C4480 ( .A1(p[130]), .A2(c[130]), .Z(s[130]) );
  XOR2D0 C4479 ( .A1(p[131]), .A2(c[131]), .Z(s[131]) );
  XOR2D0 C4478 ( .A1(p[132]), .A2(c[132]), .Z(s[132]) );
  XOR2D0 C4477 ( .A1(p[133]), .A2(c[133]), .Z(s[133]) );
  XOR2D0 C4476 ( .A1(p[134]), .A2(c[134]), .Z(s[134]) );
  XOR2D0 C4475 ( .A1(p[135]), .A2(c[135]), .Z(s[135]) );
  XOR2D0 C4474 ( .A1(p[136]), .A2(c[136]), .Z(s[136]) );
  XOR2D0 C4473 ( .A1(p[137]), .A2(c[137]), .Z(s[137]) );
  XOR2D0 C4472 ( .A1(p[138]), .A2(c[138]), .Z(s[138]) );
  XOR2D0 C4471 ( .A1(p[139]), .A2(c[139]), .Z(s[139]) );
  XOR2D0 C4470 ( .A1(p[140]), .A2(c[140]), .Z(s[140]) );
  XOR2D0 C4469 ( .A1(p[141]), .A2(c[141]), .Z(s[141]) );
  XOR2D0 C4468 ( .A1(p[142]), .A2(c[142]), .Z(s[142]) );
  XOR2D0 C4467 ( .A1(p[143]), .A2(c[143]), .Z(s[143]) );
  XOR2D0 C4466 ( .A1(p[144]), .A2(c[144]), .Z(s[144]) );
  XOR2D0 C4465 ( .A1(p[145]), .A2(c[145]), .Z(s[145]) );
  XOR2D0 C4464 ( .A1(p[146]), .A2(c[146]), .Z(s[146]) );
  XOR2D0 C4463 ( .A1(p[147]), .A2(c[147]), .Z(s[147]) );
  XOR2D0 C4462 ( .A1(p[148]), .A2(c[148]), .Z(s[148]) );
  XOR2D0 C4461 ( .A1(p[149]), .A2(c[149]), .Z(s[149]) );
  XOR2D0 C4460 ( .A1(p[150]), .A2(c[150]), .Z(s[150]) );
  XOR2D0 C4459 ( .A1(p[151]), .A2(c[151]), .Z(s[151]) );
  XOR2D0 C4458 ( .A1(p[152]), .A2(c[152]), .Z(s[152]) );
  XOR2D0 C4457 ( .A1(p[153]), .A2(c[153]), .Z(s[153]) );
  XOR2D0 C4456 ( .A1(p[154]), .A2(c[154]), .Z(s[154]) );
  XOR2D0 C4455 ( .A1(p[155]), .A2(c[155]), .Z(s[155]) );
  XOR2D0 C4454 ( .A1(p[156]), .A2(c[156]), .Z(s[156]) );
  XOR2D0 C4453 ( .A1(p[157]), .A2(c[157]), .Z(s[157]) );
  XOR2D0 C4452 ( .A1(p[158]), .A2(c[158]), .Z(s[158]) );
  XOR2D0 C4451 ( .A1(p[159]), .A2(c[159]), .Z(s[159]) );
  XOR2D0 C4450 ( .A1(p[160]), .A2(c[160]), .Z(s[160]) );
  XOR2D0 C4449 ( .A1(p[161]), .A2(c[161]), .Z(s[161]) );
  XOR2D0 C4448 ( .A1(p[162]), .A2(c[162]), .Z(s[162]) );
  XOR2D0 C4447 ( .A1(p[163]), .A2(c[163]), .Z(s[163]) );
  XOR2D0 C4446 ( .A1(p[164]), .A2(c[164]), .Z(s[164]) );
  XOR2D0 C4445 ( .A1(p[165]), .A2(c[165]), .Z(s[165]) );
  XOR2D0 C4444 ( .A1(p[166]), .A2(c[166]), .Z(s[166]) );
  XOR2D0 C4443 ( .A1(p[167]), .A2(c[167]), .Z(s[167]) );
  XOR2D0 C4442 ( .A1(p[168]), .A2(c[168]), .Z(s[168]) );
  XOR2D0 C4441 ( .A1(p[169]), .A2(c[169]), .Z(s[169]) );
  XOR2D0 C4440 ( .A1(p[170]), .A2(c[170]), .Z(s[170]) );
  XOR2D0 C4439 ( .A1(p[171]), .A2(c[171]), .Z(s[171]) );
  XOR2D0 C4438 ( .A1(p[172]), .A2(c[172]), .Z(s[172]) );
  XOR2D0 C4437 ( .A1(p[173]), .A2(c[173]), .Z(s[173]) );
  XOR2D0 C4436 ( .A1(p[174]), .A2(c[174]), .Z(s[174]) );
  XOR2D0 C4435 ( .A1(p[175]), .A2(c[175]), .Z(s[175]) );
  XOR2D0 C4434 ( .A1(p[176]), .A2(c[176]), .Z(s[176]) );
  XOR2D0 C4433 ( .A1(p[177]), .A2(c[177]), .Z(s[177]) );
  XOR2D0 C4432 ( .A1(p[178]), .A2(c[178]), .Z(s[178]) );
  XOR2D0 C4431 ( .A1(p[179]), .A2(c[179]), .Z(s[179]) );
  XOR2D0 C4430 ( .A1(p[180]), .A2(c[180]), .Z(s[180]) );
  XOR2D0 C4429 ( .A1(p[181]), .A2(c[181]), .Z(s[181]) );
  XOR2D0 C4428 ( .A1(p[182]), .A2(c[182]), .Z(s[182]) );
  XOR2D0 C4427 ( .A1(p[183]), .A2(c[183]), .Z(s[183]) );
  XOR2D0 C4426 ( .A1(p[184]), .A2(c[184]), .Z(s[184]) );
  XOR2D0 C4425 ( .A1(p[185]), .A2(c[185]), .Z(s[185]) );
  XOR2D0 C4424 ( .A1(p[186]), .A2(c[186]), .Z(s[186]) );
  XOR2D0 C4423 ( .A1(p[187]), .A2(c[187]), .Z(s[187]) );
  XOR2D0 C4422 ( .A1(p[188]), .A2(c[188]), .Z(s[188]) );
  XOR2D0 C4421 ( .A1(p[189]), .A2(c[189]), .Z(s[189]) );
  XOR2D0 C4420 ( .A1(p[190]), .A2(c[190]), .Z(s[190]) );
  XOR2D0 C4419 ( .A1(p[191]), .A2(c[191]), .Z(s[191]) );
  XOR2D0 C4418 ( .A1(p[192]), .A2(c[192]), .Z(s[192]) );
  XOR2D0 C4417 ( .A1(p[193]), .A2(c[193]), .Z(s[193]) );
  XOR2D0 C4416 ( .A1(p[194]), .A2(c[194]), .Z(s[194]) );
  XOR2D0 C4415 ( .A1(p[195]), .A2(c[195]), .Z(s[195]) );
  XOR2D0 C4414 ( .A1(p[196]), .A2(c[196]), .Z(s[196]) );
  XOR2D0 C4413 ( .A1(p[197]), .A2(c[197]), .Z(s[197]) );
  XOR2D0 C4412 ( .A1(p[198]), .A2(c[198]), .Z(s[198]) );
  XOR2D0 C4411 ( .A1(p[199]), .A2(c[199]), .Z(s[199]) );
  XOR2D0 C4410 ( .A1(p[200]), .A2(c[200]), .Z(s[200]) );
  XOR2D0 C4409 ( .A1(p[201]), .A2(c[201]), .Z(s[201]) );
  XOR2D0 C4408 ( .A1(p[202]), .A2(c[202]), .Z(s[202]) );
  XOR2D0 C4407 ( .A1(p[203]), .A2(c[203]), .Z(s[203]) );
  XOR2D0 C4406 ( .A1(p[204]), .A2(c[204]), .Z(s[204]) );
  XOR2D0 C4405 ( .A1(p[205]), .A2(c[205]), .Z(s[205]) );
  XOR2D0 C4404 ( .A1(p[206]), .A2(c[206]), .Z(s[206]) );
  XOR2D0 C4403 ( .A1(p[207]), .A2(c[207]), .Z(s[207]) );
  XOR2D0 C4402 ( .A1(p[208]), .A2(c[208]), .Z(s[208]) );
  XOR2D0 C4401 ( .A1(p[209]), .A2(c[209]), .Z(s[209]) );
  XOR2D0 C4400 ( .A1(p[210]), .A2(c[210]), .Z(s[210]) );
  XOR2D0 C4399 ( .A1(p[211]), .A2(c[211]), .Z(s[211]) );
  XOR2D0 C4398 ( .A1(p[212]), .A2(c[212]), .Z(s[212]) );
  XOR2D0 C4397 ( .A1(p[213]), .A2(c[213]), .Z(s[213]) );
  XOR2D0 C4396 ( .A1(p[214]), .A2(c[214]), .Z(s[214]) );
  XOR2D0 C4395 ( .A1(p[215]), .A2(c[215]), .Z(s[215]) );
  XOR2D0 C4394 ( .A1(p[216]), .A2(c[216]), .Z(s[216]) );
  XOR2D0 C4393 ( .A1(p[217]), .A2(c[217]), .Z(s[217]) );
  XOR2D0 C4392 ( .A1(p[218]), .A2(c[218]), .Z(s[218]) );
  XOR2D0 C4391 ( .A1(p[219]), .A2(c[219]), .Z(s[219]) );
  XOR2D0 C4390 ( .A1(p[220]), .A2(c[220]), .Z(s[220]) );
  XOR2D0 C4389 ( .A1(p[221]), .A2(c[221]), .Z(s[221]) );
  XOR2D0 C4388 ( .A1(p[222]), .A2(c[222]), .Z(s[222]) );
  XOR2D0 C4387 ( .A1(p[223]), .A2(c[223]), .Z(s[223]) );
  XOR2D0 C4386 ( .A1(p[224]), .A2(c[224]), .Z(s[224]) );
  XOR2D0 C4385 ( .A1(p[225]), .A2(c[225]), .Z(s[225]) );
  XOR2D0 C4384 ( .A1(p[226]), .A2(c[226]), .Z(s[226]) );
  XOR2D0 C4383 ( .A1(p[227]), .A2(c[227]), .Z(s[227]) );
  XOR2D0 C4382 ( .A1(p[228]), .A2(c[228]), .Z(s[228]) );
  XOR2D0 C4381 ( .A1(p[229]), .A2(c[229]), .Z(s[229]) );
  XOR2D0 C4380 ( .A1(p[230]), .A2(c[230]), .Z(s[230]) );
  XOR2D0 C4379 ( .A1(p[231]), .A2(c[231]), .Z(s[231]) );
  XOR2D0 C4378 ( .A1(p[232]), .A2(c[232]), .Z(s[232]) );
  XOR2D0 C4377 ( .A1(p[233]), .A2(c[233]), .Z(s[233]) );
  XOR2D0 C4376 ( .A1(p[234]), .A2(c[234]), .Z(s[234]) );
  XOR2D0 C4375 ( .A1(p[235]), .A2(c[235]), .Z(s[235]) );
  XOR2D0 C4374 ( .A1(p[236]), .A2(c[236]), .Z(s[236]) );
  XOR2D0 C4373 ( .A1(p[237]), .A2(c[237]), .Z(s[237]) );
  XOR2D0 C4372 ( .A1(p[238]), .A2(c[238]), .Z(s[238]) );
  XOR2D0 C4371 ( .A1(p[239]), .A2(c[239]), .Z(s[239]) );
  XOR2D0 C4370 ( .A1(p[240]), .A2(c[240]), .Z(s[240]) );
  XOR2D0 C4369 ( .A1(p[241]), .A2(c[241]), .Z(s[241]) );
  XOR2D0 C4368 ( .A1(p[242]), .A2(c[242]), .Z(s[242]) );
  XOR2D0 C4367 ( .A1(p[243]), .A2(c[243]), .Z(s[243]) );
  XOR2D0 C4366 ( .A1(p[244]), .A2(c[244]), .Z(s[244]) );
  XOR2D0 C4365 ( .A1(p[245]), .A2(c[245]), .Z(s[245]) );
  XOR2D0 C4364 ( .A1(p[246]), .A2(c[246]), .Z(s[246]) );
  XOR2D0 C4363 ( .A1(p[247]), .A2(c[247]), .Z(s[247]) );
  XOR2D0 C4362 ( .A1(p[248]), .A2(c[248]), .Z(s[248]) );
  XOR2D0 C4361 ( .A1(p[249]), .A2(c[249]), .Z(s[249]) );
  XOR2D0 C4360 ( .A1(p[250]), .A2(c[250]), .Z(s[250]) );
  XOR2D0 C4359 ( .A1(p[251]), .A2(c[251]), .Z(s[251]) );
  XOR2D0 C4358 ( .A1(p[252]), .A2(c[252]), .Z(s[252]) );
  XOR2D0 C4357 ( .A1(p[253]), .A2(c[253]), .Z(s[253]) );
  XOR2D0 C4356 ( .A1(p[254]), .A2(c[254]), .Z(s[254]) );
  XOR2D0 C4355 ( .A1(p[255]), .A2(c[255]), .Z(s[255]) );
  XOR2D0 C4354 ( .A1(p[256]), .A2(c[256]), .Z(s[256]) );
  XOR2D0 C4353 ( .A1(p[257]), .A2(c[257]), .Z(s[257]) );
  XOR2D0 C4352 ( .A1(p[258]), .A2(c[258]), .Z(s[258]) );
  XOR2D0 C4351 ( .A1(p[259]), .A2(c[259]), .Z(s[259]) );
  XOR2D0 C4350 ( .A1(p[260]), .A2(c[260]), .Z(s[260]) );
  XOR2D0 C4349 ( .A1(p[261]), .A2(c[261]), .Z(s[261]) );
  XOR2D0 C4348 ( .A1(p[262]), .A2(c[262]), .Z(s[262]) );
  XOR2D0 C4347 ( .A1(p[263]), .A2(c[263]), .Z(s[263]) );
  XOR2D0 C4346 ( .A1(p[264]), .A2(c[264]), .Z(s[264]) );
  XOR2D0 C4345 ( .A1(p[265]), .A2(c[265]), .Z(s[265]) );
  XOR2D0 C4344 ( .A1(p[266]), .A2(c[266]), .Z(s[266]) );
  XOR2D0 C4343 ( .A1(p[267]), .A2(c[267]), .Z(s[267]) );
  XOR2D0 C4342 ( .A1(p[268]), .A2(c[268]), .Z(s[268]) );
  XOR2D0 C4341 ( .A1(p[269]), .A2(c[269]), .Z(s[269]) );
  XOR2D0 C4340 ( .A1(p[270]), .A2(c[270]), .Z(s[270]) );
  XOR2D0 C4339 ( .A1(p[271]), .A2(c[271]), .Z(s[271]) );
  XOR2D0 C4338 ( .A1(p[272]), .A2(c[272]), .Z(s[272]) );
  XOR2D0 C4337 ( .A1(p[273]), .A2(c[273]), .Z(s[273]) );
  XOR2D0 C4336 ( .A1(p[274]), .A2(c[274]), .Z(s[274]) );
  XOR2D0 C4335 ( .A1(p[275]), .A2(c[275]), .Z(s[275]) );
  XOR2D0 C4334 ( .A1(p[276]), .A2(c[276]), .Z(s[276]) );
  XOR2D0 C4333 ( .A1(p[277]), .A2(c[277]), .Z(s[277]) );
  XOR2D0 C4332 ( .A1(p[278]), .A2(c[278]), .Z(s[278]) );
  XOR2D0 C4331 ( .A1(p[279]), .A2(c[279]), .Z(s[279]) );
  XOR2D0 C4330 ( .A1(p[280]), .A2(c[280]), .Z(s[280]) );
  XOR2D0 C4329 ( .A1(p[281]), .A2(c[281]), .Z(s[281]) );
  XOR2D0 C4328 ( .A1(p[282]), .A2(c[282]), .Z(s[282]) );
  XOR2D0 C4327 ( .A1(p[283]), .A2(c[283]), .Z(s[283]) );
  XOR2D0 C4326 ( .A1(p[284]), .A2(c[284]), .Z(s[284]) );
  XOR2D0 C4325 ( .A1(p[285]), .A2(c[285]), .Z(s[285]) );
  XOR2D0 C4324 ( .A1(p[286]), .A2(c[286]), .Z(s[286]) );
  XOR2D0 C4323 ( .A1(p[287]), .A2(c[287]), .Z(s[287]) );
  XOR2D0 C4322 ( .A1(p[288]), .A2(c[288]), .Z(s[288]) );
  XOR2D0 C4321 ( .A1(p[289]), .A2(c[289]), .Z(s[289]) );
  XOR2D0 C4320 ( .A1(p[290]), .A2(c[290]), .Z(s[290]) );
  XOR2D0 C4319 ( .A1(p[291]), .A2(c[291]), .Z(s[291]) );
  XOR2D0 C4318 ( .A1(p[292]), .A2(c[292]), .Z(s[292]) );
  XOR2D0 C4317 ( .A1(p[293]), .A2(c[293]), .Z(s[293]) );
  XOR2D0 C4316 ( .A1(p[294]), .A2(c[294]), .Z(s[294]) );
  XOR2D0 C4315 ( .A1(p[295]), .A2(c[295]), .Z(s[295]) );
  XOR2D0 C4314 ( .A1(p[296]), .A2(c[296]), .Z(s[296]) );
  XOR2D0 C4313 ( .A1(p[297]), .A2(c[297]), .Z(s[297]) );
  XOR2D0 C4312 ( .A1(p[298]), .A2(c[298]), .Z(s[298]) );
  XOR2D0 C4311 ( .A1(p[299]), .A2(c[299]), .Z(s[299]) );
  XOR2D0 C4310 ( .A1(p[300]), .A2(c[300]), .Z(s[300]) );
  XOR2D0 C4309 ( .A1(p[301]), .A2(c[301]), .Z(s[301]) );
  XOR2D0 C4308 ( .A1(p[302]), .A2(c[302]), .Z(s[302]) );
  XOR2D0 C4307 ( .A1(p[303]), .A2(c[303]), .Z(s[303]) );
  XOR2D0 C4306 ( .A1(p[304]), .A2(c[304]), .Z(s[304]) );
  XOR2D0 C4305 ( .A1(p[305]), .A2(c[305]), .Z(s[305]) );
  XOR2D0 C4304 ( .A1(p[306]), .A2(c[306]), .Z(s[306]) );
  XOR2D0 C4303 ( .A1(p[307]), .A2(c[307]), .Z(s[307]) );
  XOR2D0 C4302 ( .A1(p[308]), .A2(c[308]), .Z(s[308]) );
  XOR2D0 C4301 ( .A1(p[309]), .A2(c[309]), .Z(s[309]) );
  XOR2D0 C4300 ( .A1(p[310]), .A2(c[310]), .Z(s[310]) );
  XOR2D0 C4299 ( .A1(p[311]), .A2(c[311]), .Z(s[311]) );
  XOR2D0 C4298 ( .A1(p[312]), .A2(c[312]), .Z(s[312]) );
  XOR2D0 C4297 ( .A1(p[313]), .A2(c[313]), .Z(s[313]) );
  XOR2D0 C4296 ( .A1(p[314]), .A2(c[314]), .Z(s[314]) );
  XOR2D0 C4295 ( .A1(p[315]), .A2(c[315]), .Z(s[315]) );
  XOR2D0 C4294 ( .A1(p[316]), .A2(c[316]), .Z(s[316]) );
  XOR2D0 C4293 ( .A1(p[317]), .A2(c[317]), .Z(s[317]) );
  XOR2D0 C4292 ( .A1(p[318]), .A2(c[318]), .Z(s[318]) );
  XOR2D0 C4291 ( .A1(p[319]), .A2(c[319]), .Z(s[319]) );
  XOR2D0 C4290 ( .A1(p[320]), .A2(c[320]), .Z(s[320]) );
  XOR2D0 C4289 ( .A1(p[321]), .A2(c[321]), .Z(s[321]) );
  XOR2D0 C4288 ( .A1(p[322]), .A2(c[322]), .Z(s[322]) );
  XOR2D0 C4287 ( .A1(p[323]), .A2(c[323]), .Z(s[323]) );
  XOR2D0 C4286 ( .A1(p[324]), .A2(c[324]), .Z(s[324]) );
  XOR2D0 C4285 ( .A1(p[325]), .A2(c[325]), .Z(s[325]) );
  XOR2D0 C4284 ( .A1(p[326]), .A2(c[326]), .Z(s[326]) );
  XOR2D0 C4283 ( .A1(p[327]), .A2(c[327]), .Z(s[327]) );
  XOR2D0 C4282 ( .A1(p[328]), .A2(c[328]), .Z(s[328]) );
  XOR2D0 C4281 ( .A1(p[329]), .A2(c[329]), .Z(s[329]) );
  XOR2D0 C4280 ( .A1(p[330]), .A2(c[330]), .Z(s[330]) );
  XOR2D0 C4279 ( .A1(p[331]), .A2(c[331]), .Z(s[331]) );
  XOR2D0 C4278 ( .A1(p[332]), .A2(c[332]), .Z(s[332]) );
  XOR2D0 C4277 ( .A1(p[333]), .A2(c[333]), .Z(s[333]) );
  XOR2D0 C4276 ( .A1(p[334]), .A2(c[334]), .Z(s[334]) );
  XOR2D0 C4275 ( .A1(p[335]), .A2(c[335]), .Z(s[335]) );
  XOR2D0 C4274 ( .A1(p[336]), .A2(c[336]), .Z(s[336]) );
  XOR2D0 C4273 ( .A1(p[337]), .A2(c[337]), .Z(s[337]) );
  XOR2D0 C4272 ( .A1(p[338]), .A2(c[338]), .Z(s[338]) );
  XOR2D0 C4271 ( .A1(p[339]), .A2(c[339]), .Z(s[339]) );
  XOR2D0 C4270 ( .A1(p[340]), .A2(c[340]), .Z(s[340]) );
  XOR2D0 C4269 ( .A1(p[341]), .A2(c[341]), .Z(s[341]) );
  XOR2D0 C4268 ( .A1(p[342]), .A2(c[342]), .Z(s[342]) );
  XOR2D0 C4267 ( .A1(p[343]), .A2(c[343]), .Z(s[343]) );
  XOR2D0 C4266 ( .A1(p[344]), .A2(c[344]), .Z(s[344]) );
  XOR2D0 C4265 ( .A1(p[345]), .A2(c[345]), .Z(s[345]) );
  XOR2D0 C4264 ( .A1(p[346]), .A2(c[346]), .Z(s[346]) );
  XOR2D0 C4263 ( .A1(p[347]), .A2(c[347]), .Z(s[347]) );
  XOR2D0 C4262 ( .A1(p[348]), .A2(c[348]), .Z(s[348]) );
  XOR2D0 C4261 ( .A1(p[349]), .A2(c[349]), .Z(s[349]) );
  XOR2D0 C4260 ( .A1(p[350]), .A2(c[350]), .Z(s[350]) );
  XOR2D0 C4259 ( .A1(p[351]), .A2(c[351]), .Z(s[351]) );
  XOR2D0 C4258 ( .A1(p[352]), .A2(c[352]), .Z(s[352]) );
  XOR2D0 C4257 ( .A1(p[353]), .A2(c[353]), .Z(s[353]) );
  XOR2D0 C4256 ( .A1(p[354]), .A2(c[354]), .Z(s[354]) );
  XOR2D0 C4255 ( .A1(p[355]), .A2(c[355]), .Z(s[355]) );
  XOR2D0 C4254 ( .A1(p[356]), .A2(c[356]), .Z(s[356]) );
  XOR2D0 C4253 ( .A1(p[357]), .A2(c[357]), .Z(s[357]) );
  XOR2D0 C4252 ( .A1(p[358]), .A2(c[358]), .Z(s[358]) );
  XOR2D0 C4251 ( .A1(p[359]), .A2(c[359]), .Z(s[359]) );
  XOR2D0 C4250 ( .A1(p[360]), .A2(c[360]), .Z(s[360]) );
  XOR2D0 C4249 ( .A1(p[361]), .A2(c[361]), .Z(s[361]) );
  XOR2D0 C4248 ( .A1(p[362]), .A2(c[362]), .Z(s[362]) );
  XOR2D0 C4247 ( .A1(p[363]), .A2(c[363]), .Z(s[363]) );
  XOR2D0 C4246 ( .A1(p[364]), .A2(c[364]), .Z(s[364]) );
  XOR2D0 C4245 ( .A1(p[365]), .A2(c[365]), .Z(s[365]) );
  XOR2D0 C4244 ( .A1(p[366]), .A2(c[366]), .Z(s[366]) );
  XOR2D0 C4243 ( .A1(p[367]), .A2(c[367]), .Z(s[367]) );
  XOR2D0 C4242 ( .A1(p[368]), .A2(c[368]), .Z(s[368]) );
  XOR2D0 C4241 ( .A1(p[369]), .A2(c[369]), .Z(s[369]) );
  XOR2D0 C4240 ( .A1(p[370]), .A2(c[370]), .Z(s[370]) );
  XOR2D0 C4239 ( .A1(p[371]), .A2(c[371]), .Z(s[371]) );
  XOR2D0 C4238 ( .A1(p[372]), .A2(c[372]), .Z(s[372]) );
  XOR2D0 C4237 ( .A1(p[373]), .A2(c[373]), .Z(s[373]) );
  XOR2D0 C4236 ( .A1(p[374]), .A2(c[374]), .Z(s[374]) );
  XOR2D0 C4235 ( .A1(p[375]), .A2(c[375]), .Z(s[375]) );
  XOR2D0 C4234 ( .A1(p[376]), .A2(c[376]), .Z(s[376]) );
  XOR2D0 C4233 ( .A1(p[377]), .A2(c[377]), .Z(s[377]) );
  XOR2D0 C4232 ( .A1(p[378]), .A2(c[378]), .Z(s[378]) );
  XOR2D0 C4231 ( .A1(p[379]), .A2(c[379]), .Z(s[379]) );
  XOR2D0 C4230 ( .A1(p[380]), .A2(c[380]), .Z(s[380]) );
  XOR2D0 C4229 ( .A1(p[381]), .A2(c[381]), .Z(s[381]) );
  XOR2D0 C4228 ( .A1(p[382]), .A2(c[382]), .Z(s[382]) );
  XOR2D0 C4227 ( .A1(p[383]), .A2(c[383]), .Z(s[383]) );
  XOR2D0 C4226 ( .A1(p[384]), .A2(c[384]), .Z(s[384]) );
  XOR2D0 C4225 ( .A1(p[385]), .A2(c[385]), .Z(s[385]) );
  XOR2D0 C4224 ( .A1(p[386]), .A2(c[386]), .Z(s[386]) );
  XOR2D0 C4223 ( .A1(p[387]), .A2(c[387]), .Z(s[387]) );
  XOR2D0 C4222 ( .A1(p[388]), .A2(c[388]), .Z(s[388]) );
  XOR2D0 C4221 ( .A1(p[389]), .A2(c[389]), .Z(s[389]) );
  XOR2D0 C4220 ( .A1(p[390]), .A2(c[390]), .Z(s[390]) );
  XOR2D0 C4219 ( .A1(p[391]), .A2(c[391]), .Z(s[391]) );
  XOR2D0 C4218 ( .A1(p[392]), .A2(c[392]), .Z(s[392]) );
  XOR2D0 C4217 ( .A1(p[393]), .A2(c[393]), .Z(s[393]) );
  XOR2D0 C4216 ( .A1(p[394]), .A2(c[394]), .Z(s[394]) );
  XOR2D0 C4215 ( .A1(p[395]), .A2(c[395]), .Z(s[395]) );
  XOR2D0 C4214 ( .A1(p[396]), .A2(c[396]), .Z(s[396]) );
  XOR2D0 C4213 ( .A1(p[397]), .A2(c[397]), .Z(s[397]) );
  XOR2D0 C4212 ( .A1(p[398]), .A2(c[398]), .Z(s[398]) );
  XOR2D0 C4211 ( .A1(p[399]), .A2(c[399]), .Z(s[399]) );
  XOR2D0 C4210 ( .A1(p[400]), .A2(c[400]), .Z(s[400]) );
  XOR2D0 C4209 ( .A1(p[401]), .A2(c[401]), .Z(s[401]) );
  XOR2D0 C4208 ( .A1(p[402]), .A2(c[402]), .Z(s[402]) );
  XOR2D0 C4207 ( .A1(p[403]), .A2(c[403]), .Z(s[403]) );
  XOR2D0 C4206 ( .A1(p[404]), .A2(c[404]), .Z(s[404]) );
  XOR2D0 C4205 ( .A1(p[405]), .A2(c[405]), .Z(s[405]) );
  XOR2D0 C4204 ( .A1(p[406]), .A2(c[406]), .Z(s[406]) );
  XOR2D0 C4203 ( .A1(p[407]), .A2(c[407]), .Z(s[407]) );
  XOR2D0 C4202 ( .A1(p[408]), .A2(c[408]), .Z(s[408]) );
  XOR2D0 C4201 ( .A1(p[409]), .A2(c[409]), .Z(s[409]) );
  XOR2D0 C4200 ( .A1(p[410]), .A2(c[410]), .Z(s[410]) );
  XOR2D0 C4199 ( .A1(p[411]), .A2(c[411]), .Z(s[411]) );
  XOR2D0 C4198 ( .A1(p[412]), .A2(c[412]), .Z(s[412]) );
  XOR2D0 C4197 ( .A1(p[413]), .A2(c[413]), .Z(s[413]) );
  XOR2D0 C4196 ( .A1(p[414]), .A2(c[414]), .Z(s[414]) );
  XOR2D0 C4195 ( .A1(p[415]), .A2(c[415]), .Z(s[415]) );
  XOR2D0 C4194 ( .A1(p[416]), .A2(c[416]), .Z(s[416]) );
  XOR2D0 C4193 ( .A1(p[417]), .A2(c[417]), .Z(s[417]) );
  XOR2D0 C4192 ( .A1(p[418]), .A2(c[418]), .Z(s[418]) );
  XOR2D0 C4191 ( .A1(p[419]), .A2(c[419]), .Z(s[419]) );
  XOR2D0 C4190 ( .A1(p[420]), .A2(c[420]), .Z(s[420]) );
  XOR2D0 C4189 ( .A1(p[421]), .A2(c[421]), .Z(s[421]) );
  XOR2D0 C4188 ( .A1(p[422]), .A2(c[422]), .Z(s[422]) );
  XOR2D0 C4187 ( .A1(p[423]), .A2(c[423]), .Z(s[423]) );
  XOR2D0 C4186 ( .A1(p[424]), .A2(c[424]), .Z(s[424]) );
  XOR2D0 C4185 ( .A1(p[425]), .A2(c[425]), .Z(s[425]) );
  XOR2D0 C4184 ( .A1(p[426]), .A2(c[426]), .Z(s[426]) );
  XOR2D0 C4183 ( .A1(p[427]), .A2(c[427]), .Z(s[427]) );
  XOR2D0 C4182 ( .A1(p[428]), .A2(c[428]), .Z(s[428]) );
  XOR2D0 C4181 ( .A1(p[429]), .A2(c[429]), .Z(s[429]) );
  XOR2D0 C4180 ( .A1(p[430]), .A2(c[430]), .Z(s[430]) );
  XOR2D0 C4179 ( .A1(p[431]), .A2(c[431]), .Z(s[431]) );
  XOR2D0 C4178 ( .A1(p[432]), .A2(c[432]), .Z(s[432]) );
  XOR2D0 C4177 ( .A1(p[433]), .A2(c[433]), .Z(s[433]) );
  XOR2D0 C4176 ( .A1(p[434]), .A2(c[434]), .Z(s[434]) );
  XOR2D0 C4175 ( .A1(p[435]), .A2(c[435]), .Z(s[435]) );
  XOR2D0 C4174 ( .A1(p[436]), .A2(c[436]), .Z(s[436]) );
  XOR2D0 C4173 ( .A1(p[437]), .A2(c[437]), .Z(s[437]) );
  XOR2D0 C4172 ( .A1(p[438]), .A2(c[438]), .Z(s[438]) );
  XOR2D0 C4171 ( .A1(p[439]), .A2(c[439]), .Z(s[439]) );
  XOR2D0 C4170 ( .A1(p[440]), .A2(c[440]), .Z(s[440]) );
  XOR2D0 C4169 ( .A1(p[441]), .A2(c[441]), .Z(s[441]) );
  XOR2D0 C4168 ( .A1(p[442]), .A2(c[442]), .Z(s[442]) );
  XOR2D0 C4167 ( .A1(p[443]), .A2(c[443]), .Z(s[443]) );
  XOR2D0 C4166 ( .A1(p[444]), .A2(c[444]), .Z(s[444]) );
  XOR2D0 C4165 ( .A1(p[445]), .A2(c[445]), .Z(s[445]) );
  XOR2D0 C4164 ( .A1(p[446]), .A2(c[446]), .Z(s[446]) );
  XOR2D0 C4163 ( .A1(p[447]), .A2(c[447]), .Z(s[447]) );
  XOR2D0 C4162 ( .A1(p[448]), .A2(c[448]), .Z(s[448]) );
  XOR2D0 C4161 ( .A1(p[449]), .A2(c[449]), .Z(s[449]) );
  XOR2D0 C4160 ( .A1(p[450]), .A2(c[450]), .Z(s[450]) );
  XOR2D0 C4159 ( .A1(p[451]), .A2(c[451]), .Z(s[451]) );
  XOR2D0 C4158 ( .A1(p[452]), .A2(c[452]), .Z(s[452]) );
  XOR2D0 C4157 ( .A1(p[453]), .A2(c[453]), .Z(s[453]) );
  XOR2D0 C4156 ( .A1(p[454]), .A2(c[454]), .Z(s[454]) );
  XOR2D0 C4155 ( .A1(p[455]), .A2(c[455]), .Z(s[455]) );
  XOR2D0 C4154 ( .A1(p[456]), .A2(c[456]), .Z(s[456]) );
  XOR2D0 C4153 ( .A1(p[457]), .A2(c[457]), .Z(s[457]) );
  XOR2D0 C4152 ( .A1(p[458]), .A2(c[458]), .Z(s[458]) );
  XOR2D0 C4151 ( .A1(p[459]), .A2(c[459]), .Z(s[459]) );
  XOR2D0 C4150 ( .A1(p[460]), .A2(c[460]), .Z(s[460]) );
  XOR2D0 C4149 ( .A1(p[461]), .A2(c[461]), .Z(s[461]) );
  XOR2D0 C4148 ( .A1(p[462]), .A2(c[462]), .Z(s[462]) );
  XOR2D0 C4147 ( .A1(p[463]), .A2(c[463]), .Z(s[463]) );
  XOR2D0 C4146 ( .A1(p[464]), .A2(c[464]), .Z(s[464]) );
  XOR2D0 C4145 ( .A1(p[465]), .A2(c[465]), .Z(s[465]) );
  XOR2D0 C4144 ( .A1(p[466]), .A2(c[466]), .Z(s[466]) );
  XOR2D0 C4143 ( .A1(p[467]), .A2(c[467]), .Z(s[467]) );
  XOR2D0 C4142 ( .A1(p[468]), .A2(c[468]), .Z(s[468]) );
  XOR2D0 C4141 ( .A1(p[469]), .A2(c[469]), .Z(s[469]) );
  XOR2D0 C4140 ( .A1(p[470]), .A2(c[470]), .Z(s[470]) );
  XOR2D0 C4139 ( .A1(p[471]), .A2(c[471]), .Z(s[471]) );
  XOR2D0 C4138 ( .A1(p[472]), .A2(c[472]), .Z(s[472]) );
  XOR2D0 C4137 ( .A1(p[473]), .A2(c[473]), .Z(s[473]) );
  XOR2D0 C4136 ( .A1(p[474]), .A2(c[474]), .Z(s[474]) );
  XOR2D0 C4135 ( .A1(p[475]), .A2(c[475]), .Z(s[475]) );
  XOR2D0 C4134 ( .A1(p[476]), .A2(c[476]), .Z(s[476]) );
  XOR2D0 C4133 ( .A1(p[477]), .A2(c[477]), .Z(s[477]) );
  XOR2D0 C4132 ( .A1(p[478]), .A2(c[478]), .Z(s[478]) );
  XOR2D0 C4131 ( .A1(p[479]), .A2(c[479]), .Z(s[479]) );
  XOR2D0 C4130 ( .A1(p[480]), .A2(c[480]), .Z(s[480]) );
  XOR2D0 C4129 ( .A1(p[481]), .A2(c[481]), .Z(s[481]) );
  XOR2D0 C4128 ( .A1(p[482]), .A2(c[482]), .Z(s[482]) );
  XOR2D0 C4127 ( .A1(p[483]), .A2(c[483]), .Z(s[483]) );
  XOR2D0 C4126 ( .A1(p[484]), .A2(c[484]), .Z(s[484]) );
  XOR2D0 C4125 ( .A1(p[485]), .A2(c[485]), .Z(s[485]) );
  XOR2D0 C4124 ( .A1(p[486]), .A2(c[486]), .Z(s[486]) );
  XOR2D0 C4123 ( .A1(p[487]), .A2(c[487]), .Z(s[487]) );
  XOR2D0 C4122 ( .A1(p[488]), .A2(c[488]), .Z(s[488]) );
  XOR2D0 C4121 ( .A1(p[489]), .A2(c[489]), .Z(s[489]) );
  XOR2D0 C4120 ( .A1(p[490]), .A2(c[490]), .Z(s[490]) );
  XOR2D0 C4119 ( .A1(p[491]), .A2(c[491]), .Z(s[491]) );
  XOR2D0 C4118 ( .A1(p[492]), .A2(c[492]), .Z(s[492]) );
  XOR2D0 C4117 ( .A1(p[493]), .A2(c[493]), .Z(s[493]) );
  XOR2D0 C4116 ( .A1(p[494]), .A2(c[494]), .Z(s[494]) );
  XOR2D0 C4115 ( .A1(p[495]), .A2(c[495]), .Z(s[495]) );
  XOR2D0 C4114 ( .A1(p[496]), .A2(c[496]), .Z(s[496]) );
  XOR2D0 C4113 ( .A1(p[497]), .A2(c[497]), .Z(s[497]) );
  XOR2D0 C4112 ( .A1(p[498]), .A2(c[498]), .Z(s[498]) );
  XOR2D0 C4111 ( .A1(p[499]), .A2(c[499]), .Z(s[499]) );
  XOR2D0 C4110 ( .A1(p[500]), .A2(c[500]), .Z(s[500]) );
  XOR2D0 C4109 ( .A1(p[501]), .A2(c[501]), .Z(s[501]) );
  XOR2D0 C4108 ( .A1(p[502]), .A2(c[502]), .Z(s[502]) );
  XOR2D0 C4107 ( .A1(p[503]), .A2(c[503]), .Z(s[503]) );
  XOR2D0 C4106 ( .A1(p[504]), .A2(c[504]), .Z(s[504]) );
  XOR2D0 C4105 ( .A1(p[505]), .A2(c[505]), .Z(s[505]) );
  XOR2D0 C4104 ( .A1(p[506]), .A2(c[506]), .Z(s[506]) );
  XOR2D0 C4103 ( .A1(p[507]), .A2(c[507]), .Z(s[507]) );
  XOR2D0 C4102 ( .A1(p[508]), .A2(c[508]), .Z(s[508]) );
  XOR2D0 C4101 ( .A1(p[509]), .A2(c[509]), .Z(s[509]) );
  XOR2D0 C4100 ( .A1(p[510]), .A2(c[510]), .Z(s[510]) );
  XOR2D0 C4099 ( .A1(p[511]), .A2(c[511]), .Z(s[511]) );
  AN2D0 C4098 ( .A1(p[510]), .A2(c[510]), .Z(N510) );
  OR2D0 C4097 ( .A1(g[510]), .A2(N510), .Z(c[511]) );
  AN2D0 C4096 ( .A1(p[509]), .A2(c[509]), .Z(N509) );
  OR2D0 C4095 ( .A1(g[509]), .A2(N509), .Z(c[510]) );
  AN2D0 C4094 ( .A1(p[508]), .A2(c[508]), .Z(N508) );
  OR2D0 C4093 ( .A1(g[508]), .A2(N508), .Z(c[509]) );
  AN2D0 C4092 ( .A1(p[507]), .A2(c[507]), .Z(N507) );
  OR2D0 C4091 ( .A1(g[507]), .A2(N507), .Z(c[508]) );
  AN2D0 C4090 ( .A1(p[506]), .A2(c[506]), .Z(N506) );
  OR2D0 C4089 ( .A1(g[506]), .A2(N506), .Z(c[507]) );
  AN2D0 C4088 ( .A1(p[505]), .A2(c[505]), .Z(N505) );
  OR2D0 C4087 ( .A1(g[505]), .A2(N505), .Z(c[506]) );
  AN2D0 C4086 ( .A1(p[504]), .A2(c[504]), .Z(N504) );
  OR2D0 C4085 ( .A1(g[504]), .A2(N504), .Z(c[505]) );
  AN2D0 C4084 ( .A1(p[503]), .A2(c[503]), .Z(N503) );
  OR2D0 C4083 ( .A1(g[503]), .A2(N503), .Z(c[504]) );
  AN2D0 C4082 ( .A1(p[502]), .A2(c[502]), .Z(N502) );
  OR2D0 C4081 ( .A1(g[502]), .A2(N502), .Z(c[503]) );
  AN2D0 C4080 ( .A1(p[501]), .A2(c[501]), .Z(N501) );
  OR2D0 C4079 ( .A1(g[501]), .A2(N501), .Z(c[502]) );
  AN2D0 C4078 ( .A1(p[500]), .A2(c[500]), .Z(N500) );
  OR2D0 C4077 ( .A1(g[500]), .A2(N500), .Z(c[501]) );
  AN2D0 C4076 ( .A1(p[499]), .A2(c[499]), .Z(N499) );
  OR2D0 C4075 ( .A1(g[499]), .A2(N499), .Z(c[500]) );
  AN2D0 C4074 ( .A1(p[498]), .A2(c[498]), .Z(N498) );
  OR2D0 C4073 ( .A1(g[498]), .A2(N498), .Z(c[499]) );
  AN2D0 C4072 ( .A1(p[497]), .A2(c[497]), .Z(N497) );
  OR2D0 C4071 ( .A1(g[497]), .A2(N497), .Z(c[498]) );
  AN2D0 C4070 ( .A1(p[496]), .A2(c[496]), .Z(N496) );
  OR2D0 C4069 ( .A1(g[496]), .A2(N496), .Z(c[497]) );
  AN2D0 C4068 ( .A1(p[495]), .A2(c[495]), .Z(N495) );
  OR2D0 C4067 ( .A1(g[495]), .A2(N495), .Z(c[496]) );
  AN2D0 C4066 ( .A1(p[494]), .A2(c[494]), .Z(N494) );
  OR2D0 C4065 ( .A1(g[494]), .A2(N494), .Z(c[495]) );
  AN2D0 C4064 ( .A1(p[493]), .A2(c[493]), .Z(N493) );
  OR2D0 C4063 ( .A1(g[493]), .A2(N493), .Z(c[494]) );
  AN2D0 C4062 ( .A1(p[492]), .A2(c[492]), .Z(N492) );
  OR2D0 C4061 ( .A1(g[492]), .A2(N492), .Z(c[493]) );
  AN2D0 C4060 ( .A1(p[491]), .A2(c[491]), .Z(N491) );
  OR2D0 C4059 ( .A1(g[491]), .A2(N491), .Z(c[492]) );
  AN2D0 C4058 ( .A1(p[490]), .A2(c[490]), .Z(N490) );
  OR2D0 C4057 ( .A1(g[490]), .A2(N490), .Z(c[491]) );
  AN2D0 C4056 ( .A1(p[489]), .A2(c[489]), .Z(N489) );
  OR2D0 C4055 ( .A1(g[489]), .A2(N489), .Z(c[490]) );
  AN2D0 C4054 ( .A1(p[488]), .A2(c[488]), .Z(N488) );
  OR2D0 C4053 ( .A1(g[488]), .A2(N488), .Z(c[489]) );
  AN2D0 C4052 ( .A1(p[487]), .A2(c[487]), .Z(N487) );
  OR2D0 C4051 ( .A1(g[487]), .A2(N487), .Z(c[488]) );
  AN2D0 C4050 ( .A1(p[486]), .A2(c[486]), .Z(N486) );
  OR2D0 C4049 ( .A1(g[486]), .A2(N486), .Z(c[487]) );
  AN2D0 C4048 ( .A1(p[485]), .A2(c[485]), .Z(N485) );
  OR2D0 C4047 ( .A1(g[485]), .A2(N485), .Z(c[486]) );
  AN2D0 C4046 ( .A1(p[484]), .A2(c[484]), .Z(N484) );
  OR2D0 C4045 ( .A1(g[484]), .A2(N484), .Z(c[485]) );
  AN2D0 C4044 ( .A1(p[483]), .A2(c[483]), .Z(N483) );
  OR2D0 C4043 ( .A1(g[483]), .A2(N483), .Z(c[484]) );
  AN2D0 C4042 ( .A1(p[482]), .A2(c[482]), .Z(N482) );
  OR2D0 C4041 ( .A1(g[482]), .A2(N482), .Z(c[483]) );
  AN2D0 C4040 ( .A1(p[481]), .A2(c[481]), .Z(N481) );
  OR2D0 C4039 ( .A1(g[481]), .A2(N481), .Z(c[482]) );
  AN2D0 C4038 ( .A1(p[480]), .A2(c[480]), .Z(N480) );
  OR2D0 C4037 ( .A1(g[480]), .A2(N480), .Z(c[481]) );
  AN2D0 C4036 ( .A1(p[479]), .A2(c[479]), .Z(N479) );
  OR2D0 C4035 ( .A1(g[479]), .A2(N479), .Z(c[480]) );
  AN2D0 C4034 ( .A1(p[478]), .A2(c[478]), .Z(N478) );
  OR2D0 C4033 ( .A1(g[478]), .A2(N478), .Z(c[479]) );
  AN2D0 C4032 ( .A1(p[477]), .A2(c[477]), .Z(N477) );
  OR2D0 C4031 ( .A1(g[477]), .A2(N477), .Z(c[478]) );
  AN2D0 C4030 ( .A1(p[476]), .A2(c[476]), .Z(N476) );
  OR2D0 C4029 ( .A1(g[476]), .A2(N476), .Z(c[477]) );
  AN2D0 C4028 ( .A1(p[475]), .A2(c[475]), .Z(N475) );
  OR2D0 C4027 ( .A1(g[475]), .A2(N475), .Z(c[476]) );
  AN2D0 C4026 ( .A1(p[474]), .A2(c[474]), .Z(N474) );
  OR2D0 C4025 ( .A1(g[474]), .A2(N474), .Z(c[475]) );
  AN2D0 C4024 ( .A1(p[473]), .A2(c[473]), .Z(N473) );
  OR2D0 C4023 ( .A1(g[473]), .A2(N473), .Z(c[474]) );
  AN2D0 C4022 ( .A1(p[472]), .A2(c[472]), .Z(N472) );
  OR2D0 C4021 ( .A1(g[472]), .A2(N472), .Z(c[473]) );
  AN2D0 C4020 ( .A1(p[471]), .A2(c[471]), .Z(N471) );
  OR2D0 C4019 ( .A1(g[471]), .A2(N471), .Z(c[472]) );
  AN2D0 C4018 ( .A1(p[470]), .A2(c[470]), .Z(N470) );
  OR2D0 C4017 ( .A1(g[470]), .A2(N470), .Z(c[471]) );
  AN2D0 C4016 ( .A1(p[469]), .A2(c[469]), .Z(N469) );
  OR2D0 C4015 ( .A1(g[469]), .A2(N469), .Z(c[470]) );
  AN2D0 C4014 ( .A1(p[468]), .A2(c[468]), .Z(N468) );
  OR2D0 C4013 ( .A1(g[468]), .A2(N468), .Z(c[469]) );
  AN2D0 C4012 ( .A1(p[467]), .A2(c[467]), .Z(N467) );
  OR2D0 C4011 ( .A1(g[467]), .A2(N467), .Z(c[468]) );
  AN2D0 C4010 ( .A1(p[466]), .A2(c[466]), .Z(N466) );
  OR2D0 C4009 ( .A1(g[466]), .A2(N466), .Z(c[467]) );
  AN2D0 C4008 ( .A1(p[465]), .A2(c[465]), .Z(N465) );
  OR2D0 C4007 ( .A1(g[465]), .A2(N465), .Z(c[466]) );
  AN2D0 C4006 ( .A1(p[464]), .A2(c[464]), .Z(N464) );
  OR2D0 C4005 ( .A1(g[464]), .A2(N464), .Z(c[465]) );
  AN2D0 C4004 ( .A1(p[463]), .A2(c[463]), .Z(N463) );
  OR2D0 C4003 ( .A1(g[463]), .A2(N463), .Z(c[464]) );
  AN2D0 C4002 ( .A1(p[462]), .A2(c[462]), .Z(N462) );
  OR2D0 C4001 ( .A1(g[462]), .A2(N462), .Z(c[463]) );
  AN2D0 C4000 ( .A1(p[461]), .A2(c[461]), .Z(N461) );
  OR2D0 C3999 ( .A1(g[461]), .A2(N461), .Z(c[462]) );
  AN2D0 C3998 ( .A1(p[460]), .A2(c[460]), .Z(N460) );
  OR2D0 C3997 ( .A1(g[460]), .A2(N460), .Z(c[461]) );
  AN2D0 C3996 ( .A1(p[459]), .A2(c[459]), .Z(N459) );
  OR2D0 C3995 ( .A1(g[459]), .A2(N459), .Z(c[460]) );
  AN2D0 C3994 ( .A1(p[458]), .A2(c[458]), .Z(N458) );
  OR2D0 C3993 ( .A1(g[458]), .A2(N458), .Z(c[459]) );
  AN2D0 C3992 ( .A1(p[457]), .A2(c[457]), .Z(N457) );
  OR2D0 C3991 ( .A1(g[457]), .A2(N457), .Z(c[458]) );
  AN2D0 C3990 ( .A1(p[456]), .A2(c[456]), .Z(N456) );
  OR2D0 C3989 ( .A1(g[456]), .A2(N456), .Z(c[457]) );
  AN2D0 C3988 ( .A1(p[455]), .A2(c[455]), .Z(N455) );
  OR2D0 C3987 ( .A1(g[455]), .A2(N455), .Z(c[456]) );
  AN2D0 C3986 ( .A1(p[454]), .A2(c[454]), .Z(N454) );
  OR2D0 C3985 ( .A1(g[454]), .A2(N454), .Z(c[455]) );
  AN2D0 C3984 ( .A1(p[453]), .A2(c[453]), .Z(N453) );
  OR2D0 C3983 ( .A1(g[453]), .A2(N453), .Z(c[454]) );
  AN2D0 C3982 ( .A1(p[452]), .A2(c[452]), .Z(N452) );
  OR2D0 C3981 ( .A1(g[452]), .A2(N452), .Z(c[453]) );
  AN2D0 C3980 ( .A1(p[451]), .A2(c[451]), .Z(N451) );
  OR2D0 C3979 ( .A1(g[451]), .A2(N451), .Z(c[452]) );
  AN2D0 C3978 ( .A1(p[450]), .A2(c[450]), .Z(N450) );
  OR2D0 C3977 ( .A1(g[450]), .A2(N450), .Z(c[451]) );
  AN2D0 C3976 ( .A1(p[449]), .A2(c[449]), .Z(N449) );
  OR2D0 C3975 ( .A1(g[449]), .A2(N449), .Z(c[450]) );
  AN2D0 C3974 ( .A1(p[448]), .A2(c[448]), .Z(N448) );
  OR2D0 C3973 ( .A1(g[448]), .A2(N448), .Z(c[449]) );
  AN2D0 C3972 ( .A1(p[447]), .A2(c[447]), .Z(N447) );
  OR2D0 C3971 ( .A1(g[447]), .A2(N447), .Z(c[448]) );
  AN2D0 C3970 ( .A1(p[446]), .A2(c[446]), .Z(N446) );
  OR2D0 C3969 ( .A1(g[446]), .A2(N446), .Z(c[447]) );
  AN2D0 C3968 ( .A1(p[445]), .A2(c[445]), .Z(N445) );
  OR2D0 C3967 ( .A1(g[445]), .A2(N445), .Z(c[446]) );
  AN2D0 C3966 ( .A1(p[444]), .A2(c[444]), .Z(N444) );
  OR2D0 C3965 ( .A1(g[444]), .A2(N444), .Z(c[445]) );
  AN2D0 C3964 ( .A1(p[443]), .A2(c[443]), .Z(N443) );
  OR2D0 C3963 ( .A1(g[443]), .A2(N443), .Z(c[444]) );
  AN2D0 C3962 ( .A1(p[442]), .A2(c[442]), .Z(N442) );
  OR2D0 C3961 ( .A1(g[442]), .A2(N442), .Z(c[443]) );
  AN2D0 C3960 ( .A1(p[441]), .A2(c[441]), .Z(N441) );
  OR2D0 C3959 ( .A1(g[441]), .A2(N441), .Z(c[442]) );
  AN2D0 C3958 ( .A1(p[440]), .A2(c[440]), .Z(N440) );
  OR2D0 C3957 ( .A1(g[440]), .A2(N440), .Z(c[441]) );
  AN2D0 C3956 ( .A1(p[439]), .A2(c[439]), .Z(N439) );
  OR2D0 C3955 ( .A1(g[439]), .A2(N439), .Z(c[440]) );
  AN2D0 C3954 ( .A1(p[438]), .A2(c[438]), .Z(N438) );
  OR2D0 C3953 ( .A1(g[438]), .A2(N438), .Z(c[439]) );
  AN2D0 C3952 ( .A1(p[437]), .A2(c[437]), .Z(N437) );
  OR2D0 C3951 ( .A1(g[437]), .A2(N437), .Z(c[438]) );
  AN2D0 C3950 ( .A1(p[436]), .A2(c[436]), .Z(N436) );
  OR2D0 C3949 ( .A1(g[436]), .A2(N436), .Z(c[437]) );
  AN2D0 C3948 ( .A1(p[435]), .A2(c[435]), .Z(N435) );
  OR2D0 C3947 ( .A1(g[435]), .A2(N435), .Z(c[436]) );
  AN2D0 C3946 ( .A1(p[434]), .A2(c[434]), .Z(N434) );
  OR2D0 C3945 ( .A1(g[434]), .A2(N434), .Z(c[435]) );
  AN2D0 C3944 ( .A1(p[433]), .A2(c[433]), .Z(N433) );
  OR2D0 C3943 ( .A1(g[433]), .A2(N433), .Z(c[434]) );
  AN2D0 C3942 ( .A1(p[432]), .A2(c[432]), .Z(N432) );
  OR2D0 C3941 ( .A1(g[432]), .A2(N432), .Z(c[433]) );
  AN2D0 C3940 ( .A1(p[431]), .A2(c[431]), .Z(N431) );
  OR2D0 C3939 ( .A1(g[431]), .A2(N431), .Z(c[432]) );
  AN2D0 C3938 ( .A1(p[430]), .A2(c[430]), .Z(N430) );
  OR2D0 C3937 ( .A1(g[430]), .A2(N430), .Z(c[431]) );
  AN2D0 C3936 ( .A1(p[429]), .A2(c[429]), .Z(N429) );
  OR2D0 C3935 ( .A1(g[429]), .A2(N429), .Z(c[430]) );
  AN2D0 C3934 ( .A1(p[428]), .A2(c[428]), .Z(N428) );
  OR2D0 C3933 ( .A1(g[428]), .A2(N428), .Z(c[429]) );
  AN2D0 C3932 ( .A1(p[427]), .A2(c[427]), .Z(N427) );
  OR2D0 C3931 ( .A1(g[427]), .A2(N427), .Z(c[428]) );
  AN2D0 C3930 ( .A1(p[426]), .A2(c[426]), .Z(N426) );
  OR2D0 C3929 ( .A1(g[426]), .A2(N426), .Z(c[427]) );
  AN2D0 C3928 ( .A1(p[425]), .A2(c[425]), .Z(N425) );
  OR2D0 C3927 ( .A1(g[425]), .A2(N425), .Z(c[426]) );
  AN2D0 C3926 ( .A1(p[424]), .A2(c[424]), .Z(N424) );
  OR2D0 C3925 ( .A1(g[424]), .A2(N424), .Z(c[425]) );
  AN2D0 C3924 ( .A1(p[423]), .A2(c[423]), .Z(N423) );
  OR2D0 C3923 ( .A1(g[423]), .A2(N423), .Z(c[424]) );
  AN2D0 C3922 ( .A1(p[422]), .A2(c[422]), .Z(N422) );
  OR2D0 C3921 ( .A1(g[422]), .A2(N422), .Z(c[423]) );
  AN2D0 C3920 ( .A1(p[421]), .A2(c[421]), .Z(N421) );
  OR2D0 C3919 ( .A1(g[421]), .A2(N421), .Z(c[422]) );
  AN2D0 C3918 ( .A1(p[420]), .A2(c[420]), .Z(N420) );
  OR2D0 C3917 ( .A1(g[420]), .A2(N420), .Z(c[421]) );
  AN2D0 C3916 ( .A1(p[419]), .A2(c[419]), .Z(N419) );
  OR2D0 C3915 ( .A1(g[419]), .A2(N419), .Z(c[420]) );
  AN2D0 C3914 ( .A1(p[418]), .A2(c[418]), .Z(N418) );
  OR2D0 C3913 ( .A1(g[418]), .A2(N418), .Z(c[419]) );
  AN2D0 C3912 ( .A1(p[417]), .A2(c[417]), .Z(N417) );
  OR2D0 C3911 ( .A1(g[417]), .A2(N417), .Z(c[418]) );
  AN2D0 C3910 ( .A1(p[416]), .A2(c[416]), .Z(N416) );
  OR2D0 C3909 ( .A1(g[416]), .A2(N416), .Z(c[417]) );
  AN2D0 C3908 ( .A1(p[415]), .A2(c[415]), .Z(N415) );
  OR2D0 C3907 ( .A1(g[415]), .A2(N415), .Z(c[416]) );
  AN2D0 C3906 ( .A1(p[414]), .A2(c[414]), .Z(N414) );
  OR2D0 C3905 ( .A1(g[414]), .A2(N414), .Z(c[415]) );
  AN2D0 C3904 ( .A1(p[413]), .A2(c[413]), .Z(N413) );
  OR2D0 C3903 ( .A1(g[413]), .A2(N413), .Z(c[414]) );
  AN2D0 C3902 ( .A1(p[412]), .A2(c[412]), .Z(N412) );
  OR2D0 C3901 ( .A1(g[412]), .A2(N412), .Z(c[413]) );
  AN2D0 C3900 ( .A1(p[411]), .A2(c[411]), .Z(N411) );
  OR2D0 C3899 ( .A1(g[411]), .A2(N411), .Z(c[412]) );
  AN2D0 C3898 ( .A1(p[410]), .A2(c[410]), .Z(N410) );
  OR2D0 C3897 ( .A1(g[410]), .A2(N410), .Z(c[411]) );
  AN2D0 C3896 ( .A1(p[409]), .A2(c[409]), .Z(N409) );
  OR2D0 C3895 ( .A1(g[409]), .A2(N409), .Z(c[410]) );
  AN2D0 C3894 ( .A1(p[408]), .A2(c[408]), .Z(N408) );
  OR2D0 C3893 ( .A1(g[408]), .A2(N408), .Z(c[409]) );
  AN2D0 C3892 ( .A1(p[407]), .A2(c[407]), .Z(N407) );
  OR2D0 C3891 ( .A1(g[407]), .A2(N407), .Z(c[408]) );
  AN2D0 C3890 ( .A1(p[406]), .A2(c[406]), .Z(N406) );
  OR2D0 C3889 ( .A1(g[406]), .A2(N406), .Z(c[407]) );
  AN2D0 C3888 ( .A1(p[405]), .A2(c[405]), .Z(N405) );
  OR2D0 C3887 ( .A1(g[405]), .A2(N405), .Z(c[406]) );
  AN2D0 C3886 ( .A1(p[404]), .A2(c[404]), .Z(N404) );
  OR2D0 C3885 ( .A1(g[404]), .A2(N404), .Z(c[405]) );
  AN2D0 C3884 ( .A1(p[403]), .A2(c[403]), .Z(N403) );
  OR2D0 C3883 ( .A1(g[403]), .A2(N403), .Z(c[404]) );
  AN2D0 C3882 ( .A1(p[402]), .A2(c[402]), .Z(N402) );
  OR2D0 C3881 ( .A1(g[402]), .A2(N402), .Z(c[403]) );
  AN2D0 C3880 ( .A1(p[401]), .A2(c[401]), .Z(N401) );
  OR2D0 C3879 ( .A1(g[401]), .A2(N401), .Z(c[402]) );
  AN2D0 C3878 ( .A1(p[400]), .A2(c[400]), .Z(N400) );
  OR2D0 C3877 ( .A1(g[400]), .A2(N400), .Z(c[401]) );
  AN2D0 C3876 ( .A1(p[399]), .A2(c[399]), .Z(N399) );
  OR2D0 C3875 ( .A1(g[399]), .A2(N399), .Z(c[400]) );
  AN2D0 C3874 ( .A1(p[398]), .A2(c[398]), .Z(N398) );
  OR2D0 C3873 ( .A1(g[398]), .A2(N398), .Z(c[399]) );
  AN2D0 C3872 ( .A1(p[397]), .A2(c[397]), .Z(N397) );
  OR2D0 C3871 ( .A1(g[397]), .A2(N397), .Z(c[398]) );
  AN2D0 C3870 ( .A1(p[396]), .A2(c[396]), .Z(N396) );
  OR2D0 C3869 ( .A1(g[396]), .A2(N396), .Z(c[397]) );
  AN2D0 C3868 ( .A1(p[395]), .A2(c[395]), .Z(N395) );
  OR2D0 C3867 ( .A1(g[395]), .A2(N395), .Z(c[396]) );
  AN2D0 C3866 ( .A1(p[394]), .A2(c[394]), .Z(N394) );
  OR2D0 C3865 ( .A1(g[394]), .A2(N394), .Z(c[395]) );
  AN2D0 C3864 ( .A1(p[393]), .A2(c[393]), .Z(N393) );
  OR2D0 C3863 ( .A1(g[393]), .A2(N393), .Z(c[394]) );
  AN2D0 C3862 ( .A1(p[392]), .A2(c[392]), .Z(N392) );
  OR2D0 C3861 ( .A1(g[392]), .A2(N392), .Z(c[393]) );
  AN2D0 C3860 ( .A1(p[391]), .A2(c[391]), .Z(N391) );
  OR2D0 C3859 ( .A1(g[391]), .A2(N391), .Z(c[392]) );
  AN2D0 C3858 ( .A1(p[390]), .A2(c[390]), .Z(N390) );
  OR2D0 C3857 ( .A1(g[390]), .A2(N390), .Z(c[391]) );
  AN2D0 C3856 ( .A1(p[389]), .A2(c[389]), .Z(N389) );
  OR2D0 C3855 ( .A1(g[389]), .A2(N389), .Z(c[390]) );
  AN2D0 C3854 ( .A1(p[388]), .A2(c[388]), .Z(N388) );
  OR2D0 C3853 ( .A1(g[388]), .A2(N388), .Z(c[389]) );
  AN2D0 C3852 ( .A1(p[387]), .A2(c[387]), .Z(N387) );
  OR2D0 C3851 ( .A1(g[387]), .A2(N387), .Z(c[388]) );
  AN2D0 C3850 ( .A1(p[386]), .A2(c[386]), .Z(N386) );
  OR2D0 C3849 ( .A1(g[386]), .A2(N386), .Z(c[387]) );
  AN2D0 C3848 ( .A1(p[385]), .A2(c[385]), .Z(N385) );
  OR2D0 C3847 ( .A1(g[385]), .A2(N385), .Z(c[386]) );
  AN2D0 C3846 ( .A1(p[384]), .A2(c[384]), .Z(N384) );
  OR2D0 C3845 ( .A1(g[384]), .A2(N384), .Z(c[385]) );
  AN2D0 C3844 ( .A1(p[383]), .A2(c[383]), .Z(N383) );
  OR2D0 C3843 ( .A1(g[383]), .A2(N383), .Z(c[384]) );
  AN2D0 C3842 ( .A1(p[382]), .A2(c[382]), .Z(N382) );
  OR2D0 C3841 ( .A1(g[382]), .A2(N382), .Z(c[383]) );
  AN2D0 C3840 ( .A1(p[381]), .A2(c[381]), .Z(N381) );
  OR2D0 C3839 ( .A1(g[381]), .A2(N381), .Z(c[382]) );
  AN2D0 C3838 ( .A1(p[380]), .A2(c[380]), .Z(N380) );
  OR2D0 C3837 ( .A1(g[380]), .A2(N380), .Z(c[381]) );
  AN2D0 C3836 ( .A1(p[379]), .A2(c[379]), .Z(N379) );
  OR2D0 C3835 ( .A1(g[379]), .A2(N379), .Z(c[380]) );
  AN2D0 C3834 ( .A1(p[378]), .A2(c[378]), .Z(N378) );
  OR2D0 C3833 ( .A1(g[378]), .A2(N378), .Z(c[379]) );
  AN2D0 C3832 ( .A1(p[377]), .A2(c[377]), .Z(N377) );
  OR2D0 C3831 ( .A1(g[377]), .A2(N377), .Z(c[378]) );
  AN2D0 C3830 ( .A1(p[376]), .A2(c[376]), .Z(N376) );
  OR2D0 C3829 ( .A1(g[376]), .A2(N376), .Z(c[377]) );
  AN2D0 C3828 ( .A1(p[375]), .A2(c[375]), .Z(N375) );
  OR2D0 C3827 ( .A1(g[375]), .A2(N375), .Z(c[376]) );
  AN2D0 C3826 ( .A1(p[374]), .A2(c[374]), .Z(N374) );
  OR2D0 C3825 ( .A1(g[374]), .A2(N374), .Z(c[375]) );
  AN2D0 C3824 ( .A1(p[373]), .A2(c[373]), .Z(N373) );
  OR2D0 C3823 ( .A1(g[373]), .A2(N373), .Z(c[374]) );
  AN2D0 C3822 ( .A1(p[372]), .A2(c[372]), .Z(N372) );
  OR2D0 C3821 ( .A1(g[372]), .A2(N372), .Z(c[373]) );
  AN2D0 C3820 ( .A1(p[371]), .A2(c[371]), .Z(N371) );
  OR2D0 C3819 ( .A1(g[371]), .A2(N371), .Z(c[372]) );
  AN2D0 C3818 ( .A1(p[370]), .A2(c[370]), .Z(N370) );
  OR2D0 C3817 ( .A1(g[370]), .A2(N370), .Z(c[371]) );
  AN2D0 C3816 ( .A1(p[369]), .A2(c[369]), .Z(N369) );
  OR2D0 C3815 ( .A1(g[369]), .A2(N369), .Z(c[370]) );
  AN2D0 C3814 ( .A1(p[368]), .A2(c[368]), .Z(N368) );
  OR2D0 C3813 ( .A1(g[368]), .A2(N368), .Z(c[369]) );
  AN2D0 C3812 ( .A1(p[367]), .A2(c[367]), .Z(N367) );
  OR2D0 C3811 ( .A1(g[367]), .A2(N367), .Z(c[368]) );
  AN2D0 C3810 ( .A1(p[366]), .A2(c[366]), .Z(N366) );
  OR2D0 C3809 ( .A1(g[366]), .A2(N366), .Z(c[367]) );
  AN2D0 C3808 ( .A1(p[365]), .A2(c[365]), .Z(N365) );
  OR2D0 C3807 ( .A1(g[365]), .A2(N365), .Z(c[366]) );
  AN2D0 C3806 ( .A1(p[364]), .A2(c[364]), .Z(N364) );
  OR2D0 C3805 ( .A1(g[364]), .A2(N364), .Z(c[365]) );
  AN2D0 C3804 ( .A1(p[363]), .A2(c[363]), .Z(N363) );
  OR2D0 C3803 ( .A1(g[363]), .A2(N363), .Z(c[364]) );
  AN2D0 C3802 ( .A1(p[362]), .A2(c[362]), .Z(N362) );
  OR2D0 C3801 ( .A1(g[362]), .A2(N362), .Z(c[363]) );
  AN2D0 C3800 ( .A1(p[361]), .A2(c[361]), .Z(N361) );
  OR2D0 C3799 ( .A1(g[361]), .A2(N361), .Z(c[362]) );
  AN2D0 C3798 ( .A1(p[360]), .A2(c[360]), .Z(N360) );
  OR2D0 C3797 ( .A1(g[360]), .A2(N360), .Z(c[361]) );
  AN2D0 C3796 ( .A1(p[359]), .A2(c[359]), .Z(N359) );
  OR2D0 C3795 ( .A1(g[359]), .A2(N359), .Z(c[360]) );
  AN2D0 C3794 ( .A1(p[358]), .A2(c[358]), .Z(N358) );
  OR2D0 C3793 ( .A1(g[358]), .A2(N358), .Z(c[359]) );
  AN2D0 C3792 ( .A1(p[357]), .A2(c[357]), .Z(N357) );
  OR2D0 C3791 ( .A1(g[357]), .A2(N357), .Z(c[358]) );
  AN2D0 C3790 ( .A1(p[356]), .A2(c[356]), .Z(N356) );
  OR2D0 C3789 ( .A1(g[356]), .A2(N356), .Z(c[357]) );
  AN2D0 C3788 ( .A1(p[355]), .A2(c[355]), .Z(N355) );
  OR2D0 C3787 ( .A1(g[355]), .A2(N355), .Z(c[356]) );
  AN2D0 C3786 ( .A1(p[354]), .A2(c[354]), .Z(N354) );
  OR2D0 C3785 ( .A1(g[354]), .A2(N354), .Z(c[355]) );
  AN2D0 C3784 ( .A1(p[353]), .A2(c[353]), .Z(N353) );
  OR2D0 C3783 ( .A1(g[353]), .A2(N353), .Z(c[354]) );
  AN2D0 C3782 ( .A1(p[352]), .A2(c[352]), .Z(N352) );
  OR2D0 C3781 ( .A1(g[352]), .A2(N352), .Z(c[353]) );
  AN2D0 C3780 ( .A1(p[351]), .A2(c[351]), .Z(N351) );
  OR2D0 C3779 ( .A1(g[351]), .A2(N351), .Z(c[352]) );
  AN2D0 C3778 ( .A1(p[350]), .A2(c[350]), .Z(N350) );
  OR2D0 C3777 ( .A1(g[350]), .A2(N350), .Z(c[351]) );
  AN2D0 C3776 ( .A1(p[349]), .A2(c[349]), .Z(N349) );
  OR2D0 C3775 ( .A1(g[349]), .A2(N349), .Z(c[350]) );
  AN2D0 C3774 ( .A1(p[348]), .A2(c[348]), .Z(N348) );
  OR2D0 C3773 ( .A1(g[348]), .A2(N348), .Z(c[349]) );
  AN2D0 C3772 ( .A1(p[347]), .A2(c[347]), .Z(N347) );
  OR2D0 C3771 ( .A1(g[347]), .A2(N347), .Z(c[348]) );
  AN2D0 C3770 ( .A1(p[346]), .A2(c[346]), .Z(N346) );
  OR2D0 C3769 ( .A1(g[346]), .A2(N346), .Z(c[347]) );
  AN2D0 C3768 ( .A1(p[345]), .A2(c[345]), .Z(N345) );
  OR2D0 C3767 ( .A1(g[345]), .A2(N345), .Z(c[346]) );
  AN2D0 C3766 ( .A1(p[344]), .A2(c[344]), .Z(N344) );
  OR2D0 C3765 ( .A1(g[344]), .A2(N344), .Z(c[345]) );
  AN2D0 C3764 ( .A1(p[343]), .A2(c[343]), .Z(N343) );
  OR2D0 C3763 ( .A1(g[343]), .A2(N343), .Z(c[344]) );
  AN2D0 C3762 ( .A1(p[342]), .A2(c[342]), .Z(N342) );
  OR2D0 C3761 ( .A1(g[342]), .A2(N342), .Z(c[343]) );
  AN2D0 C3760 ( .A1(p[341]), .A2(c[341]), .Z(N341) );
  OR2D0 C3759 ( .A1(g[341]), .A2(N341), .Z(c[342]) );
  AN2D0 C3758 ( .A1(p[340]), .A2(c[340]), .Z(N340) );
  OR2D0 C3757 ( .A1(g[340]), .A2(N340), .Z(c[341]) );
  AN2D0 C3756 ( .A1(p[339]), .A2(c[339]), .Z(N339) );
  OR2D0 C3755 ( .A1(g[339]), .A2(N339), .Z(c[340]) );
  AN2D0 C3754 ( .A1(p[338]), .A2(c[338]), .Z(N338) );
  OR2D0 C3753 ( .A1(g[338]), .A2(N338), .Z(c[339]) );
  AN2D0 C3752 ( .A1(p[337]), .A2(c[337]), .Z(N337) );
  OR2D0 C3751 ( .A1(g[337]), .A2(N337), .Z(c[338]) );
  AN2D0 C3750 ( .A1(p[336]), .A2(c[336]), .Z(N336) );
  OR2D0 C3749 ( .A1(g[336]), .A2(N336), .Z(c[337]) );
  AN2D0 C3748 ( .A1(p[335]), .A2(c[335]), .Z(N335) );
  OR2D0 C3747 ( .A1(g[335]), .A2(N335), .Z(c[336]) );
  AN2D0 C3746 ( .A1(p[334]), .A2(c[334]), .Z(N334) );
  OR2D0 C3745 ( .A1(g[334]), .A2(N334), .Z(c[335]) );
  AN2D0 C3744 ( .A1(p[333]), .A2(c[333]), .Z(N333) );
  OR2D0 C3743 ( .A1(g[333]), .A2(N333), .Z(c[334]) );
  AN2D0 C3742 ( .A1(p[332]), .A2(c[332]), .Z(N332) );
  OR2D0 C3741 ( .A1(g[332]), .A2(N332), .Z(c[333]) );
  AN2D0 C3740 ( .A1(p[331]), .A2(c[331]), .Z(N331) );
  OR2D0 C3739 ( .A1(g[331]), .A2(N331), .Z(c[332]) );
  AN2D0 C3738 ( .A1(p[330]), .A2(c[330]), .Z(N330) );
  OR2D0 C3737 ( .A1(g[330]), .A2(N330), .Z(c[331]) );
  AN2D0 C3736 ( .A1(p[329]), .A2(c[329]), .Z(N329) );
  OR2D0 C3735 ( .A1(g[329]), .A2(N329), .Z(c[330]) );
  AN2D0 C3734 ( .A1(p[328]), .A2(c[328]), .Z(N328) );
  OR2D0 C3733 ( .A1(g[328]), .A2(N328), .Z(c[329]) );
  AN2D0 C3732 ( .A1(p[327]), .A2(c[327]), .Z(N327) );
  OR2D0 C3731 ( .A1(g[327]), .A2(N327), .Z(c[328]) );
  AN2D0 C3730 ( .A1(p[326]), .A2(c[326]), .Z(N326) );
  OR2D0 C3729 ( .A1(g[326]), .A2(N326), .Z(c[327]) );
  AN2D0 C3728 ( .A1(p[325]), .A2(c[325]), .Z(N325) );
  OR2D0 C3727 ( .A1(g[325]), .A2(N325), .Z(c[326]) );
  AN2D0 C3726 ( .A1(p[324]), .A2(c[324]), .Z(N324) );
  OR2D0 C3725 ( .A1(g[324]), .A2(N324), .Z(c[325]) );
  AN2D0 C3724 ( .A1(p[323]), .A2(c[323]), .Z(N323) );
  OR2D0 C3723 ( .A1(g[323]), .A2(N323), .Z(c[324]) );
  AN2D0 C3722 ( .A1(p[322]), .A2(c[322]), .Z(N322) );
  OR2D0 C3721 ( .A1(g[322]), .A2(N322), .Z(c[323]) );
  AN2D0 C3720 ( .A1(p[321]), .A2(c[321]), .Z(N321) );
  OR2D0 C3719 ( .A1(g[321]), .A2(N321), .Z(c[322]) );
  AN2D0 C3718 ( .A1(p[320]), .A2(c[320]), .Z(N320) );
  OR2D0 C3717 ( .A1(g[320]), .A2(N320), .Z(c[321]) );
  AN2D0 C3716 ( .A1(p[319]), .A2(c[319]), .Z(N319) );
  OR2D0 C3715 ( .A1(g[319]), .A2(N319), .Z(c[320]) );
  AN2D0 C3714 ( .A1(p[318]), .A2(c[318]), .Z(N318) );
  OR2D0 C3713 ( .A1(g[318]), .A2(N318), .Z(c[319]) );
  AN2D0 C3712 ( .A1(p[317]), .A2(c[317]), .Z(N317) );
  OR2D0 C3711 ( .A1(g[317]), .A2(N317), .Z(c[318]) );
  AN2D0 C3710 ( .A1(p[316]), .A2(c[316]), .Z(N316) );
  OR2D0 C3709 ( .A1(g[316]), .A2(N316), .Z(c[317]) );
  AN2D0 C3708 ( .A1(p[315]), .A2(c[315]), .Z(N315) );
  OR2D0 C3707 ( .A1(g[315]), .A2(N315), .Z(c[316]) );
  AN2D0 C3706 ( .A1(p[314]), .A2(c[314]), .Z(N314) );
  OR2D0 C3705 ( .A1(g[314]), .A2(N314), .Z(c[315]) );
  AN2D0 C3704 ( .A1(p[313]), .A2(c[313]), .Z(N313) );
  OR2D0 C3703 ( .A1(g[313]), .A2(N313), .Z(c[314]) );
  AN2D0 C3702 ( .A1(p[312]), .A2(c[312]), .Z(N312) );
  OR2D0 C3701 ( .A1(g[312]), .A2(N312), .Z(c[313]) );
  AN2D0 C3700 ( .A1(p[311]), .A2(c[311]), .Z(N311) );
  OR2D0 C3699 ( .A1(g[311]), .A2(N311), .Z(c[312]) );
  AN2D0 C3698 ( .A1(p[310]), .A2(c[310]), .Z(N310) );
  OR2D0 C3697 ( .A1(g[310]), .A2(N310), .Z(c[311]) );
  AN2D0 C3696 ( .A1(p[309]), .A2(c[309]), .Z(N309) );
  OR2D0 C3695 ( .A1(g[309]), .A2(N309), .Z(c[310]) );
  AN2D0 C3694 ( .A1(p[308]), .A2(c[308]), .Z(N308) );
  OR2D0 C3693 ( .A1(g[308]), .A2(N308), .Z(c[309]) );
  AN2D0 C3692 ( .A1(p[307]), .A2(c[307]), .Z(N307) );
  OR2D0 C3691 ( .A1(g[307]), .A2(N307), .Z(c[308]) );
  AN2D0 C3690 ( .A1(p[306]), .A2(c[306]), .Z(N306) );
  OR2D0 C3689 ( .A1(g[306]), .A2(N306), .Z(c[307]) );
  AN2D0 C3688 ( .A1(p[305]), .A2(c[305]), .Z(N305) );
  OR2D0 C3687 ( .A1(g[305]), .A2(N305), .Z(c[306]) );
  AN2D0 C3686 ( .A1(p[304]), .A2(c[304]), .Z(N304) );
  OR2D0 C3685 ( .A1(g[304]), .A2(N304), .Z(c[305]) );
  AN2D0 C3684 ( .A1(p[303]), .A2(c[303]), .Z(N303) );
  OR2D0 C3683 ( .A1(g[303]), .A2(N303), .Z(c[304]) );
  AN2D0 C3682 ( .A1(p[302]), .A2(c[302]), .Z(N302) );
  OR2D0 C3681 ( .A1(g[302]), .A2(N302), .Z(c[303]) );
  AN2D0 C3680 ( .A1(p[301]), .A2(c[301]), .Z(N301) );
  OR2D0 C3679 ( .A1(g[301]), .A2(N301), .Z(c[302]) );
  AN2D0 C3678 ( .A1(p[300]), .A2(c[300]), .Z(N300) );
  OR2D0 C3677 ( .A1(g[300]), .A2(N300), .Z(c[301]) );
  AN2D0 C3676 ( .A1(p[299]), .A2(c[299]), .Z(N299) );
  OR2D0 C3675 ( .A1(g[299]), .A2(N299), .Z(c[300]) );
  AN2D0 C3674 ( .A1(p[298]), .A2(c[298]), .Z(N298) );
  OR2D0 C3673 ( .A1(g[298]), .A2(N298), .Z(c[299]) );
  AN2D0 C3672 ( .A1(p[297]), .A2(c[297]), .Z(N297) );
  OR2D0 C3671 ( .A1(g[297]), .A2(N297), .Z(c[298]) );
  AN2D0 C3670 ( .A1(p[296]), .A2(c[296]), .Z(N296) );
  OR2D0 C3669 ( .A1(g[296]), .A2(N296), .Z(c[297]) );
  AN2D0 C3668 ( .A1(p[295]), .A2(c[295]), .Z(N295) );
  OR2D0 C3667 ( .A1(g[295]), .A2(N295), .Z(c[296]) );
  AN2D0 C3666 ( .A1(p[294]), .A2(c[294]), .Z(N294) );
  OR2D0 C3665 ( .A1(g[294]), .A2(N294), .Z(c[295]) );
  AN2D0 C3664 ( .A1(p[293]), .A2(c[293]), .Z(N293) );
  OR2D0 C3663 ( .A1(g[293]), .A2(N293), .Z(c[294]) );
  AN2D0 C3662 ( .A1(p[292]), .A2(c[292]), .Z(N292) );
  OR2D0 C3661 ( .A1(g[292]), .A2(N292), .Z(c[293]) );
  AN2D0 C3660 ( .A1(p[291]), .A2(c[291]), .Z(N291) );
  OR2D0 C3659 ( .A1(g[291]), .A2(N291), .Z(c[292]) );
  AN2D0 C3658 ( .A1(p[290]), .A2(c[290]), .Z(N290) );
  OR2D0 C3657 ( .A1(g[290]), .A2(N290), .Z(c[291]) );
  AN2D0 C3656 ( .A1(p[289]), .A2(c[289]), .Z(N289) );
  OR2D0 C3655 ( .A1(g[289]), .A2(N289), .Z(c[290]) );
  AN2D0 C3654 ( .A1(p[288]), .A2(c[288]), .Z(N288) );
  OR2D0 C3653 ( .A1(g[288]), .A2(N288), .Z(c[289]) );
  AN2D0 C3652 ( .A1(p[287]), .A2(c[287]), .Z(N287) );
  OR2D0 C3651 ( .A1(g[287]), .A2(N287), .Z(c[288]) );
  AN2D0 C3650 ( .A1(p[286]), .A2(c[286]), .Z(N286) );
  OR2D0 C3649 ( .A1(g[286]), .A2(N286), .Z(c[287]) );
  AN2D0 C3648 ( .A1(p[285]), .A2(c[285]), .Z(N285) );
  OR2D0 C3647 ( .A1(g[285]), .A2(N285), .Z(c[286]) );
  AN2D0 C3646 ( .A1(p[284]), .A2(c[284]), .Z(N284) );
  OR2D0 C3645 ( .A1(g[284]), .A2(N284), .Z(c[285]) );
  AN2D0 C3644 ( .A1(p[283]), .A2(c[283]), .Z(N283) );
  OR2D0 C3643 ( .A1(g[283]), .A2(N283), .Z(c[284]) );
  AN2D0 C3642 ( .A1(p[282]), .A2(c[282]), .Z(N282) );
  OR2D0 C3641 ( .A1(g[282]), .A2(N282), .Z(c[283]) );
  AN2D0 C3640 ( .A1(p[281]), .A2(c[281]), .Z(N281) );
  OR2D0 C3639 ( .A1(g[281]), .A2(N281), .Z(c[282]) );
  AN2D0 C3638 ( .A1(p[280]), .A2(c[280]), .Z(N280) );
  OR2D0 C3637 ( .A1(g[280]), .A2(N280), .Z(c[281]) );
  AN2D0 C3636 ( .A1(p[279]), .A2(c[279]), .Z(N279) );
  OR2D0 C3635 ( .A1(g[279]), .A2(N279), .Z(c[280]) );
  AN2D0 C3634 ( .A1(p[278]), .A2(c[278]), .Z(N278) );
  OR2D0 C3633 ( .A1(g[278]), .A2(N278), .Z(c[279]) );
  AN2D0 C3632 ( .A1(p[277]), .A2(c[277]), .Z(N277) );
  OR2D0 C3631 ( .A1(g[277]), .A2(N277), .Z(c[278]) );
  AN2D0 C3630 ( .A1(p[276]), .A2(c[276]), .Z(N276) );
  OR2D0 C3629 ( .A1(g[276]), .A2(N276), .Z(c[277]) );
  AN2D0 C3628 ( .A1(p[275]), .A2(c[275]), .Z(N275) );
  OR2D0 C3627 ( .A1(g[275]), .A2(N275), .Z(c[276]) );
  AN2D0 C3626 ( .A1(p[274]), .A2(c[274]), .Z(N274) );
  OR2D0 C3625 ( .A1(g[274]), .A2(N274), .Z(c[275]) );
  AN2D0 C3624 ( .A1(p[273]), .A2(c[273]), .Z(N273) );
  OR2D0 C3623 ( .A1(g[273]), .A2(N273), .Z(c[274]) );
  AN2D0 C3622 ( .A1(p[272]), .A2(c[272]), .Z(N272) );
  OR2D0 C3621 ( .A1(g[272]), .A2(N272), .Z(c[273]) );
  AN2D0 C3620 ( .A1(p[271]), .A2(c[271]), .Z(N271) );
  OR2D0 C3619 ( .A1(g[271]), .A2(N271), .Z(c[272]) );
  AN2D0 C3618 ( .A1(p[270]), .A2(c[270]), .Z(N270) );
  OR2D0 C3617 ( .A1(g[270]), .A2(N270), .Z(c[271]) );
  AN2D0 C3616 ( .A1(p[269]), .A2(c[269]), .Z(N269) );
  OR2D0 C3615 ( .A1(g[269]), .A2(N269), .Z(c[270]) );
  AN2D0 C3614 ( .A1(p[268]), .A2(c[268]), .Z(N268) );
  OR2D0 C3613 ( .A1(g[268]), .A2(N268), .Z(c[269]) );
  AN2D0 C3612 ( .A1(p[267]), .A2(c[267]), .Z(N267) );
  OR2D0 C3611 ( .A1(g[267]), .A2(N267), .Z(c[268]) );
  AN2D0 C3610 ( .A1(p[266]), .A2(c[266]), .Z(N266) );
  OR2D0 C3609 ( .A1(g[266]), .A2(N266), .Z(c[267]) );
  AN2D0 C3608 ( .A1(p[265]), .A2(c[265]), .Z(N265) );
  OR2D0 C3607 ( .A1(g[265]), .A2(N265), .Z(c[266]) );
  AN2D0 C3606 ( .A1(p[264]), .A2(c[264]), .Z(N264) );
  OR2D0 C3605 ( .A1(g[264]), .A2(N264), .Z(c[265]) );
  AN2D0 C3604 ( .A1(p[263]), .A2(c[263]), .Z(N263) );
  OR2D0 C3603 ( .A1(g[263]), .A2(N263), .Z(c[264]) );
  AN2D0 C3602 ( .A1(p[262]), .A2(c[262]), .Z(N262) );
  OR2D0 C3601 ( .A1(g[262]), .A2(N262), .Z(c[263]) );
  AN2D0 C3600 ( .A1(p[261]), .A2(c[261]), .Z(N261) );
  OR2D0 C3599 ( .A1(g[261]), .A2(N261), .Z(c[262]) );
  AN2D0 C3598 ( .A1(p[260]), .A2(c[260]), .Z(N260) );
  OR2D0 C3597 ( .A1(g[260]), .A2(N260), .Z(c[261]) );
  AN2D0 C3596 ( .A1(p[259]), .A2(c[259]), .Z(N259) );
  OR2D0 C3595 ( .A1(g[259]), .A2(N259), .Z(c[260]) );
  AN2D0 C3594 ( .A1(p[258]), .A2(c[258]), .Z(N258) );
  OR2D0 C3593 ( .A1(g[258]), .A2(N258), .Z(c[259]) );
  AN2D0 C3592 ( .A1(p[257]), .A2(c[257]), .Z(N257) );
  OR2D0 C3591 ( .A1(g[257]), .A2(N257), .Z(c[258]) );
  AN2D0 C3590 ( .A1(p[256]), .A2(c[256]), .Z(N256) );
  OR2D0 C3589 ( .A1(g[256]), .A2(N256), .Z(c[257]) );
  AN2D0 C3588 ( .A1(p[255]), .A2(c[255]), .Z(N255) );
  OR2D0 C3587 ( .A1(g[255]), .A2(N255), .Z(c[256]) );
  AN2D0 C3586 ( .A1(p[254]), .A2(c[254]), .Z(N254) );
  OR2D0 C3585 ( .A1(g[254]), .A2(N254), .Z(c[255]) );
  AN2D0 C3584 ( .A1(p[253]), .A2(c[253]), .Z(N253) );
  OR2D0 C3583 ( .A1(g[253]), .A2(N253), .Z(c[254]) );
  AN2D0 C3582 ( .A1(p[252]), .A2(c[252]), .Z(N252) );
  OR2D0 C3581 ( .A1(g[252]), .A2(N252), .Z(c[253]) );
  AN2D0 C3580 ( .A1(p[251]), .A2(c[251]), .Z(N251) );
  OR2D0 C3579 ( .A1(g[251]), .A2(N251), .Z(c[252]) );
  AN2D0 C3578 ( .A1(p[250]), .A2(c[250]), .Z(N250) );
  OR2D0 C3577 ( .A1(g[250]), .A2(N250), .Z(c[251]) );
  AN2D0 C3576 ( .A1(p[249]), .A2(c[249]), .Z(N249) );
  OR2D0 C3575 ( .A1(g[249]), .A2(N249), .Z(c[250]) );
  AN2D0 C3574 ( .A1(p[248]), .A2(c[248]), .Z(N248) );
  OR2D0 C3573 ( .A1(g[248]), .A2(N248), .Z(c[249]) );
  AN2D0 C3572 ( .A1(p[247]), .A2(c[247]), .Z(N247) );
  OR2D0 C3571 ( .A1(g[247]), .A2(N247), .Z(c[248]) );
  AN2D0 C3570 ( .A1(p[246]), .A2(c[246]), .Z(N246) );
  OR2D0 C3569 ( .A1(g[246]), .A2(N246), .Z(c[247]) );
  AN2D0 C3568 ( .A1(p[245]), .A2(c[245]), .Z(N245) );
  OR2D0 C3567 ( .A1(g[245]), .A2(N245), .Z(c[246]) );
  AN2D0 C3566 ( .A1(p[244]), .A2(c[244]), .Z(N244) );
  OR2D0 C3565 ( .A1(g[244]), .A2(N244), .Z(c[245]) );
  AN2D0 C3564 ( .A1(p[243]), .A2(c[243]), .Z(N243) );
  OR2D0 C3563 ( .A1(g[243]), .A2(N243), .Z(c[244]) );
  AN2D0 C3562 ( .A1(p[242]), .A2(c[242]), .Z(N242) );
  OR2D0 C3561 ( .A1(g[242]), .A2(N242), .Z(c[243]) );
  AN2D0 C3560 ( .A1(p[241]), .A2(c[241]), .Z(N241) );
  OR2D0 C3559 ( .A1(g[241]), .A2(N241), .Z(c[242]) );
  AN2D0 C3558 ( .A1(p[240]), .A2(c[240]), .Z(N240) );
  OR2D0 C3557 ( .A1(g[240]), .A2(N240), .Z(c[241]) );
  AN2D0 C3556 ( .A1(p[239]), .A2(c[239]), .Z(N239) );
  OR2D0 C3555 ( .A1(g[239]), .A2(N239), .Z(c[240]) );
  AN2D0 C3554 ( .A1(p[238]), .A2(c[238]), .Z(N238) );
  OR2D0 C3553 ( .A1(g[238]), .A2(N238), .Z(c[239]) );
  AN2D0 C3552 ( .A1(p[237]), .A2(c[237]), .Z(N237) );
  OR2D0 C3551 ( .A1(g[237]), .A2(N237), .Z(c[238]) );
  AN2D0 C3550 ( .A1(p[236]), .A2(c[236]), .Z(N236) );
  OR2D0 C3549 ( .A1(g[236]), .A2(N236), .Z(c[237]) );
  AN2D0 C3548 ( .A1(p[235]), .A2(c[235]), .Z(N235) );
  OR2D0 C3547 ( .A1(g[235]), .A2(N235), .Z(c[236]) );
  AN2D0 C3546 ( .A1(p[234]), .A2(c[234]), .Z(N234) );
  OR2D0 C3545 ( .A1(g[234]), .A2(N234), .Z(c[235]) );
  AN2D0 C3544 ( .A1(p[233]), .A2(c[233]), .Z(N233) );
  OR2D0 C3543 ( .A1(g[233]), .A2(N233), .Z(c[234]) );
  AN2D0 C3542 ( .A1(p[232]), .A2(c[232]), .Z(N232) );
  OR2D0 C3541 ( .A1(g[232]), .A2(N232), .Z(c[233]) );
  AN2D0 C3540 ( .A1(p[231]), .A2(c[231]), .Z(N231) );
  OR2D0 C3539 ( .A1(g[231]), .A2(N231), .Z(c[232]) );
  AN2D0 C3538 ( .A1(p[230]), .A2(c[230]), .Z(N230) );
  OR2D0 C3537 ( .A1(g[230]), .A2(N230), .Z(c[231]) );
  AN2D0 C3536 ( .A1(p[229]), .A2(c[229]), .Z(N229) );
  OR2D0 C3535 ( .A1(g[229]), .A2(N229), .Z(c[230]) );
  AN2D0 C3534 ( .A1(p[228]), .A2(c[228]), .Z(N228) );
  OR2D0 C3533 ( .A1(g[228]), .A2(N228), .Z(c[229]) );
  AN2D0 C3532 ( .A1(p[227]), .A2(c[227]), .Z(N227) );
  OR2D0 C3531 ( .A1(g[227]), .A2(N227), .Z(c[228]) );
  AN2D0 C3530 ( .A1(p[226]), .A2(c[226]), .Z(N226) );
  OR2D0 C3529 ( .A1(g[226]), .A2(N226), .Z(c[227]) );
  AN2D0 C3528 ( .A1(p[225]), .A2(c[225]), .Z(N225) );
  OR2D0 C3527 ( .A1(g[225]), .A2(N225), .Z(c[226]) );
  AN2D0 C3526 ( .A1(p[224]), .A2(c[224]), .Z(N224) );
  OR2D0 C3525 ( .A1(g[224]), .A2(N224), .Z(c[225]) );
  AN2D0 C3524 ( .A1(p[223]), .A2(c[223]), .Z(N223) );
  OR2D0 C3523 ( .A1(g[223]), .A2(N223), .Z(c[224]) );
  AN2D0 C3522 ( .A1(p[222]), .A2(c[222]), .Z(N222) );
  OR2D0 C3521 ( .A1(g[222]), .A2(N222), .Z(c[223]) );
  AN2D0 C3520 ( .A1(p[221]), .A2(c[221]), .Z(N221) );
  OR2D0 C3519 ( .A1(g[221]), .A2(N221), .Z(c[222]) );
  AN2D0 C3518 ( .A1(p[220]), .A2(c[220]), .Z(N220) );
  OR2D0 C3517 ( .A1(g[220]), .A2(N220), .Z(c[221]) );
  AN2D0 C3516 ( .A1(p[219]), .A2(c[219]), .Z(N219) );
  OR2D0 C3515 ( .A1(g[219]), .A2(N219), .Z(c[220]) );
  AN2D0 C3514 ( .A1(p[218]), .A2(c[218]), .Z(N218) );
  OR2D0 C3513 ( .A1(g[218]), .A2(N218), .Z(c[219]) );
  AN2D0 C3512 ( .A1(p[217]), .A2(c[217]), .Z(N217) );
  OR2D0 C3511 ( .A1(g[217]), .A2(N217), .Z(c[218]) );
  AN2D0 C3510 ( .A1(p[216]), .A2(c[216]), .Z(N216) );
  OR2D0 C3509 ( .A1(g[216]), .A2(N216), .Z(c[217]) );
  AN2D0 C3508 ( .A1(p[215]), .A2(c[215]), .Z(N215) );
  OR2D0 C3507 ( .A1(g[215]), .A2(N215), .Z(c[216]) );
  AN2D0 C3506 ( .A1(p[214]), .A2(c[214]), .Z(N214) );
  OR2D0 C3505 ( .A1(g[214]), .A2(N214), .Z(c[215]) );
  AN2D0 C3504 ( .A1(p[213]), .A2(c[213]), .Z(N213) );
  OR2D0 C3503 ( .A1(g[213]), .A2(N213), .Z(c[214]) );
  AN2D0 C3502 ( .A1(p[212]), .A2(c[212]), .Z(N212) );
  OR2D0 C3501 ( .A1(g[212]), .A2(N212), .Z(c[213]) );
  AN2D0 C3500 ( .A1(p[211]), .A2(c[211]), .Z(N211) );
  OR2D0 C3499 ( .A1(g[211]), .A2(N211), .Z(c[212]) );
  AN2D0 C3498 ( .A1(p[210]), .A2(c[210]), .Z(N210) );
  OR2D0 C3497 ( .A1(g[210]), .A2(N210), .Z(c[211]) );
  AN2D0 C3496 ( .A1(p[209]), .A2(c[209]), .Z(N209) );
  OR2D0 C3495 ( .A1(g[209]), .A2(N209), .Z(c[210]) );
  AN2D0 C3494 ( .A1(p[208]), .A2(c[208]), .Z(N208) );
  OR2D0 C3493 ( .A1(g[208]), .A2(N208), .Z(c[209]) );
  AN2D0 C3492 ( .A1(p[207]), .A2(c[207]), .Z(N207) );
  OR2D0 C3491 ( .A1(g[207]), .A2(N207), .Z(c[208]) );
  AN2D0 C3490 ( .A1(p[206]), .A2(c[206]), .Z(N206) );
  OR2D0 C3489 ( .A1(g[206]), .A2(N206), .Z(c[207]) );
  AN2D0 C3488 ( .A1(p[205]), .A2(c[205]), .Z(N205) );
  OR2D0 C3487 ( .A1(g[205]), .A2(N205), .Z(c[206]) );
  AN2D0 C3486 ( .A1(p[204]), .A2(c[204]), .Z(N204) );
  OR2D0 C3485 ( .A1(g[204]), .A2(N204), .Z(c[205]) );
  AN2D0 C3484 ( .A1(p[203]), .A2(c[203]), .Z(N203) );
  OR2D0 C3483 ( .A1(g[203]), .A2(N203), .Z(c[204]) );
  AN2D0 C3482 ( .A1(p[202]), .A2(c[202]), .Z(N202) );
  OR2D0 C3481 ( .A1(g[202]), .A2(N202), .Z(c[203]) );
  AN2D0 C3480 ( .A1(p[201]), .A2(c[201]), .Z(N201) );
  OR2D0 C3479 ( .A1(g[201]), .A2(N201), .Z(c[202]) );
  AN2D0 C3478 ( .A1(p[200]), .A2(c[200]), .Z(N200) );
  OR2D0 C3477 ( .A1(g[200]), .A2(N200), .Z(c[201]) );
  AN2D0 C3476 ( .A1(p[199]), .A2(c[199]), .Z(N199) );
  OR2D0 C3475 ( .A1(g[199]), .A2(N199), .Z(c[200]) );
  AN2D0 C3474 ( .A1(p[198]), .A2(c[198]), .Z(N198) );
  OR2D0 C3473 ( .A1(g[198]), .A2(N198), .Z(c[199]) );
  AN2D0 C3472 ( .A1(p[197]), .A2(c[197]), .Z(N197) );
  OR2D0 C3471 ( .A1(g[197]), .A2(N197), .Z(c[198]) );
  AN2D0 C3470 ( .A1(p[196]), .A2(c[196]), .Z(N196) );
  OR2D0 C3469 ( .A1(g[196]), .A2(N196), .Z(c[197]) );
  AN2D0 C3468 ( .A1(p[195]), .A2(c[195]), .Z(N195) );
  OR2D0 C3467 ( .A1(g[195]), .A2(N195), .Z(c[196]) );
  AN2D0 C3466 ( .A1(p[194]), .A2(c[194]), .Z(N194) );
  OR2D0 C3465 ( .A1(g[194]), .A2(N194), .Z(c[195]) );
  AN2D0 C3464 ( .A1(p[193]), .A2(c[193]), .Z(N193) );
  OR2D0 C3463 ( .A1(g[193]), .A2(N193), .Z(c[194]) );
  AN2D0 C3462 ( .A1(p[192]), .A2(c[192]), .Z(N192) );
  OR2D0 C3461 ( .A1(g[192]), .A2(N192), .Z(c[193]) );
  AN2D0 C3460 ( .A1(p[191]), .A2(c[191]), .Z(N191) );
  OR2D0 C3459 ( .A1(g[191]), .A2(N191), .Z(c[192]) );
  AN2D0 C3458 ( .A1(p[190]), .A2(c[190]), .Z(N190) );
  OR2D0 C3457 ( .A1(g[190]), .A2(N190), .Z(c[191]) );
  AN2D0 C3456 ( .A1(p[189]), .A2(c[189]), .Z(N189) );
  OR2D0 C3455 ( .A1(g[189]), .A2(N189), .Z(c[190]) );
  AN2D0 C3454 ( .A1(p[188]), .A2(c[188]), .Z(N188) );
  OR2D0 C3453 ( .A1(g[188]), .A2(N188), .Z(c[189]) );
  AN2D0 C3452 ( .A1(p[187]), .A2(c[187]), .Z(N187) );
  OR2D0 C3451 ( .A1(g[187]), .A2(N187), .Z(c[188]) );
  AN2D0 C3450 ( .A1(p[186]), .A2(c[186]), .Z(N186) );
  OR2D0 C3449 ( .A1(g[186]), .A2(N186), .Z(c[187]) );
  AN2D0 C3448 ( .A1(p[185]), .A2(c[185]), .Z(N185) );
  OR2D0 C3447 ( .A1(g[185]), .A2(N185), .Z(c[186]) );
  AN2D0 C3446 ( .A1(p[184]), .A2(c[184]), .Z(N184) );
  OR2D0 C3445 ( .A1(g[184]), .A2(N184), .Z(c[185]) );
  AN2D0 C3444 ( .A1(p[183]), .A2(c[183]), .Z(N183) );
  OR2D0 C3443 ( .A1(g[183]), .A2(N183), .Z(c[184]) );
  AN2D0 C3442 ( .A1(p[182]), .A2(c[182]), .Z(N182) );
  OR2D0 C3441 ( .A1(g[182]), .A2(N182), .Z(c[183]) );
  AN2D0 C3440 ( .A1(p[181]), .A2(c[181]), .Z(N181) );
  OR2D0 C3439 ( .A1(g[181]), .A2(N181), .Z(c[182]) );
  AN2D0 C3438 ( .A1(p[180]), .A2(c[180]), .Z(N180) );
  OR2D0 C3437 ( .A1(g[180]), .A2(N180), .Z(c[181]) );
  AN2D0 C3436 ( .A1(p[179]), .A2(c[179]), .Z(N179) );
  OR2D0 C3435 ( .A1(g[179]), .A2(N179), .Z(c[180]) );
  AN2D0 C3434 ( .A1(p[178]), .A2(c[178]), .Z(N178) );
  OR2D0 C3433 ( .A1(g[178]), .A2(N178), .Z(c[179]) );
  AN2D0 C3432 ( .A1(p[177]), .A2(c[177]), .Z(N177) );
  OR2D0 C3431 ( .A1(g[177]), .A2(N177), .Z(c[178]) );
  AN2D0 C3430 ( .A1(p[176]), .A2(c[176]), .Z(N176) );
  OR2D0 C3429 ( .A1(g[176]), .A2(N176), .Z(c[177]) );
  AN2D0 C3428 ( .A1(p[175]), .A2(c[175]), .Z(N175) );
  OR2D0 C3427 ( .A1(g[175]), .A2(N175), .Z(c[176]) );
  AN2D0 C3426 ( .A1(p[174]), .A2(c[174]), .Z(N174) );
  OR2D0 C3425 ( .A1(g[174]), .A2(N174), .Z(c[175]) );
  AN2D0 C3424 ( .A1(p[173]), .A2(c[173]), .Z(N173) );
  OR2D0 C3423 ( .A1(g[173]), .A2(N173), .Z(c[174]) );
  AN2D0 C3422 ( .A1(p[172]), .A2(c[172]), .Z(N172) );
  OR2D0 C3421 ( .A1(g[172]), .A2(N172), .Z(c[173]) );
  AN2D0 C3420 ( .A1(p[171]), .A2(c[171]), .Z(N171) );
  OR2D0 C3419 ( .A1(g[171]), .A2(N171), .Z(c[172]) );
  AN2D0 C3418 ( .A1(p[170]), .A2(c[170]), .Z(N170) );
  OR2D0 C3417 ( .A1(g[170]), .A2(N170), .Z(c[171]) );
  AN2D0 C3416 ( .A1(p[169]), .A2(c[169]), .Z(N169) );
  OR2D0 C3415 ( .A1(g[169]), .A2(N169), .Z(c[170]) );
  AN2D0 C3414 ( .A1(p[168]), .A2(c[168]), .Z(N168) );
  OR2D0 C3413 ( .A1(g[168]), .A2(N168), .Z(c[169]) );
  AN2D0 C3412 ( .A1(p[167]), .A2(c[167]), .Z(N167) );
  OR2D0 C3411 ( .A1(g[167]), .A2(N167), .Z(c[168]) );
  AN2D0 C3410 ( .A1(p[166]), .A2(c[166]), .Z(N166) );
  OR2D0 C3409 ( .A1(g[166]), .A2(N166), .Z(c[167]) );
  AN2D0 C3408 ( .A1(p[165]), .A2(c[165]), .Z(N165) );
  OR2D0 C3407 ( .A1(g[165]), .A2(N165), .Z(c[166]) );
  AN2D0 C3406 ( .A1(p[164]), .A2(c[164]), .Z(N164) );
  OR2D0 C3405 ( .A1(g[164]), .A2(N164), .Z(c[165]) );
  AN2D0 C3404 ( .A1(p[163]), .A2(c[163]), .Z(N163) );
  OR2D0 C3403 ( .A1(g[163]), .A2(N163), .Z(c[164]) );
  AN2D0 C3402 ( .A1(p[162]), .A2(c[162]), .Z(N162) );
  OR2D0 C3401 ( .A1(g[162]), .A2(N162), .Z(c[163]) );
  AN2D0 C3400 ( .A1(p[161]), .A2(c[161]), .Z(N161) );
  OR2D0 C3399 ( .A1(g[161]), .A2(N161), .Z(c[162]) );
  AN2D0 C3398 ( .A1(p[160]), .A2(c[160]), .Z(N160) );
  OR2D0 C3397 ( .A1(g[160]), .A2(N160), .Z(c[161]) );
  AN2D0 C3396 ( .A1(p[159]), .A2(c[159]), .Z(N159) );
  OR2D0 C3395 ( .A1(g[159]), .A2(N159), .Z(c[160]) );
  AN2D0 C3394 ( .A1(p[158]), .A2(c[158]), .Z(N158) );
  OR2D0 C3393 ( .A1(g[158]), .A2(N158), .Z(c[159]) );
  AN2D0 C3392 ( .A1(p[157]), .A2(c[157]), .Z(N157) );
  OR2D0 C3391 ( .A1(g[157]), .A2(N157), .Z(c[158]) );
  AN2D0 C3390 ( .A1(p[156]), .A2(c[156]), .Z(N156) );
  OR2D0 C3389 ( .A1(g[156]), .A2(N156), .Z(c[157]) );
  AN2D0 C3388 ( .A1(p[155]), .A2(c[155]), .Z(N155) );
  OR2D0 C3387 ( .A1(g[155]), .A2(N155), .Z(c[156]) );
  AN2D0 C3386 ( .A1(p[154]), .A2(c[154]), .Z(N154) );
  OR2D0 C3385 ( .A1(g[154]), .A2(N154), .Z(c[155]) );
  AN2D0 C3384 ( .A1(p[153]), .A2(c[153]), .Z(N153) );
  OR2D0 C3383 ( .A1(g[153]), .A2(N153), .Z(c[154]) );
  AN2D0 C3382 ( .A1(p[152]), .A2(c[152]), .Z(N152) );
  OR2D0 C3381 ( .A1(g[152]), .A2(N152), .Z(c[153]) );
  AN2D0 C3380 ( .A1(p[151]), .A2(c[151]), .Z(N151) );
  OR2D0 C3379 ( .A1(g[151]), .A2(N151), .Z(c[152]) );
  AN2D0 C3378 ( .A1(p[150]), .A2(c[150]), .Z(N150) );
  OR2D0 C3377 ( .A1(g[150]), .A2(N150), .Z(c[151]) );
  AN2D0 C3376 ( .A1(p[149]), .A2(c[149]), .Z(N149) );
  OR2D0 C3375 ( .A1(g[149]), .A2(N149), .Z(c[150]) );
  AN2D0 C3374 ( .A1(p[148]), .A2(c[148]), .Z(N148) );
  OR2D0 C3373 ( .A1(g[148]), .A2(N148), .Z(c[149]) );
  AN2D0 C3372 ( .A1(p[147]), .A2(c[147]), .Z(N147) );
  OR2D0 C3371 ( .A1(g[147]), .A2(N147), .Z(c[148]) );
  AN2D0 C3370 ( .A1(p[146]), .A2(c[146]), .Z(N146) );
  OR2D0 C3369 ( .A1(g[146]), .A2(N146), .Z(c[147]) );
  AN2D0 C3368 ( .A1(p[145]), .A2(c[145]), .Z(N145) );
  OR2D0 C3367 ( .A1(g[145]), .A2(N145), .Z(c[146]) );
  AN2D0 C3366 ( .A1(p[144]), .A2(c[144]), .Z(N144) );
  OR2D0 C3365 ( .A1(g[144]), .A2(N144), .Z(c[145]) );
  AN2D0 C3364 ( .A1(p[143]), .A2(c[143]), .Z(N143) );
  OR2D0 C3363 ( .A1(g[143]), .A2(N143), .Z(c[144]) );
  AN2D0 C3362 ( .A1(p[142]), .A2(c[142]), .Z(N142) );
  OR2D0 C3361 ( .A1(g[142]), .A2(N142), .Z(c[143]) );
  AN2D0 C3360 ( .A1(p[141]), .A2(c[141]), .Z(N141) );
  OR2D0 C3359 ( .A1(g[141]), .A2(N141), .Z(c[142]) );
  AN2D0 C3358 ( .A1(p[140]), .A2(c[140]), .Z(N140) );
  OR2D0 C3357 ( .A1(g[140]), .A2(N140), .Z(c[141]) );
  AN2D0 C3356 ( .A1(p[139]), .A2(c[139]), .Z(N139) );
  OR2D0 C3355 ( .A1(g[139]), .A2(N139), .Z(c[140]) );
  AN2D0 C3354 ( .A1(p[138]), .A2(c[138]), .Z(N138) );
  OR2D0 C3353 ( .A1(g[138]), .A2(N138), .Z(c[139]) );
  AN2D0 C3352 ( .A1(p[137]), .A2(c[137]), .Z(N137) );
  OR2D0 C3351 ( .A1(g[137]), .A2(N137), .Z(c[138]) );
  AN2D0 C3350 ( .A1(p[136]), .A2(c[136]), .Z(N136) );
  OR2D0 C3349 ( .A1(g[136]), .A2(N136), .Z(c[137]) );
  AN2D0 C3348 ( .A1(p[135]), .A2(c[135]), .Z(N135) );
  OR2D0 C3347 ( .A1(g[135]), .A2(N135), .Z(c[136]) );
  AN2D0 C3346 ( .A1(p[134]), .A2(c[134]), .Z(N134) );
  OR2D0 C3345 ( .A1(g[134]), .A2(N134), .Z(c[135]) );
  AN2D0 C3344 ( .A1(p[133]), .A2(c[133]), .Z(N133) );
  OR2D0 C3343 ( .A1(g[133]), .A2(N133), .Z(c[134]) );
  AN2D0 C3342 ( .A1(p[132]), .A2(c[132]), .Z(N132) );
  OR2D0 C3341 ( .A1(g[132]), .A2(N132), .Z(c[133]) );
  AN2D0 C3340 ( .A1(p[131]), .A2(c[131]), .Z(N131) );
  OR2D0 C3339 ( .A1(g[131]), .A2(N131), .Z(c[132]) );
  AN2D0 C3338 ( .A1(p[130]), .A2(c[130]), .Z(N130) );
  OR2D0 C3337 ( .A1(g[130]), .A2(N130), .Z(c[131]) );
  AN2D0 C3336 ( .A1(p[129]), .A2(c[129]), .Z(N129) );
  OR2D0 C3335 ( .A1(g[129]), .A2(N129), .Z(c[130]) );
  AN2D0 C3334 ( .A1(p[128]), .A2(c[128]), .Z(N128) );
  OR2D0 C3333 ( .A1(g[128]), .A2(N128), .Z(c[129]) );
  AN2D0 C3332 ( .A1(p[127]), .A2(c[127]), .Z(N127) );
  OR2D0 C3331 ( .A1(g[127]), .A2(N127), .Z(c[128]) );
  AN2D0 C3330 ( .A1(p[126]), .A2(c[126]), .Z(N126) );
  OR2D0 C3329 ( .A1(g[126]), .A2(N126), .Z(c[127]) );
  AN2D0 C3328 ( .A1(p[125]), .A2(c[125]), .Z(N125) );
  OR2D0 C3327 ( .A1(g[125]), .A2(N125), .Z(c[126]) );
  AN2D0 C3326 ( .A1(p[124]), .A2(c[124]), .Z(N124) );
  OR2D0 C3325 ( .A1(g[124]), .A2(N124), .Z(c[125]) );
  AN2D0 C3324 ( .A1(p[123]), .A2(c[123]), .Z(N123) );
  OR2D0 C3323 ( .A1(g[123]), .A2(N123), .Z(c[124]) );
  AN2D0 C3322 ( .A1(p[122]), .A2(c[122]), .Z(N122) );
  OR2D0 C3321 ( .A1(g[122]), .A2(N122), .Z(c[123]) );
  AN2D0 C3320 ( .A1(p[121]), .A2(c[121]), .Z(N121) );
  OR2D0 C3319 ( .A1(g[121]), .A2(N121), .Z(c[122]) );
  AN2D0 C3318 ( .A1(p[120]), .A2(c[120]), .Z(N120) );
  OR2D0 C3317 ( .A1(g[120]), .A2(N120), .Z(c[121]) );
  AN2D0 C3316 ( .A1(p[119]), .A2(c[119]), .Z(N119) );
  OR2D0 C3315 ( .A1(g[119]), .A2(N119), .Z(c[120]) );
  AN2D0 C3314 ( .A1(p[118]), .A2(c[118]), .Z(N118) );
  OR2D0 C3313 ( .A1(g[118]), .A2(N118), .Z(c[119]) );
  AN2D0 C3312 ( .A1(p[117]), .A2(c[117]), .Z(N117) );
  OR2D0 C3311 ( .A1(g[117]), .A2(N117), .Z(c[118]) );
  AN2D0 C3310 ( .A1(p[116]), .A2(c[116]), .Z(N116) );
  OR2D0 C3309 ( .A1(g[116]), .A2(N116), .Z(c[117]) );
  AN2D0 C3308 ( .A1(p[115]), .A2(c[115]), .Z(N115) );
  OR2D0 C3307 ( .A1(g[115]), .A2(N115), .Z(c[116]) );
  AN2D0 C3306 ( .A1(p[114]), .A2(c[114]), .Z(N114) );
  OR2D0 C3305 ( .A1(g[114]), .A2(N114), .Z(c[115]) );
  AN2D0 C3304 ( .A1(p[113]), .A2(c[113]), .Z(N113) );
  OR2D0 C3303 ( .A1(g[113]), .A2(N113), .Z(c[114]) );
  AN2D0 C3302 ( .A1(p[112]), .A2(c[112]), .Z(N112) );
  OR2D0 C3301 ( .A1(g[112]), .A2(N112), .Z(c[113]) );
  AN2D0 C3300 ( .A1(p[111]), .A2(c[111]), .Z(N111) );
  OR2D0 C3299 ( .A1(g[111]), .A2(N111), .Z(c[112]) );
  AN2D0 C3298 ( .A1(p[110]), .A2(c[110]), .Z(N110) );
  OR2D0 C3297 ( .A1(g[110]), .A2(N110), .Z(c[111]) );
  AN2D0 C3296 ( .A1(p[109]), .A2(c[109]), .Z(N109) );
  OR2D0 C3295 ( .A1(g[109]), .A2(N109), .Z(c[110]) );
  AN2D0 C3294 ( .A1(p[108]), .A2(c[108]), .Z(N108) );
  OR2D0 C3293 ( .A1(g[108]), .A2(N108), .Z(c[109]) );
  AN2D0 C3292 ( .A1(p[107]), .A2(c[107]), .Z(N107) );
  OR2D0 C3291 ( .A1(g[107]), .A2(N107), .Z(c[108]) );
  AN2D0 C3290 ( .A1(p[106]), .A2(c[106]), .Z(N106) );
  OR2D0 C3289 ( .A1(g[106]), .A2(N106), .Z(c[107]) );
  AN2D0 C3288 ( .A1(p[105]), .A2(c[105]), .Z(N105) );
  OR2D0 C3287 ( .A1(g[105]), .A2(N105), .Z(c[106]) );
  AN2D0 C3286 ( .A1(p[104]), .A2(c[104]), .Z(N104) );
  OR2D0 C3285 ( .A1(g[104]), .A2(N104), .Z(c[105]) );
  AN2D0 C3284 ( .A1(p[103]), .A2(c[103]), .Z(N103) );
  OR2D0 C3283 ( .A1(g[103]), .A2(N103), .Z(c[104]) );
  AN2D0 C3282 ( .A1(p[102]), .A2(c[102]), .Z(N102) );
  OR2D0 C3281 ( .A1(g[102]), .A2(N102), .Z(c[103]) );
  AN2D0 C3280 ( .A1(p[101]), .A2(c[101]), .Z(N101) );
  OR2D0 C3279 ( .A1(g[101]), .A2(N101), .Z(c[102]) );
  AN2D0 C3278 ( .A1(p[100]), .A2(c[100]), .Z(N100) );
  OR2D0 C3277 ( .A1(g[100]), .A2(N100), .Z(c[101]) );
  AN2D0 C3276 ( .A1(p[99]), .A2(c[99]), .Z(N99) );
  OR2D0 C3275 ( .A1(g[99]), .A2(N99), .Z(c[100]) );
  AN2D0 C3274 ( .A1(p[98]), .A2(c[98]), .Z(N98) );
  OR2D0 C3273 ( .A1(g[98]), .A2(N98), .Z(c[99]) );
  AN2D0 C3272 ( .A1(p[97]), .A2(c[97]), .Z(N97) );
  OR2D0 C3271 ( .A1(g[97]), .A2(N97), .Z(c[98]) );
  AN2D0 C3270 ( .A1(p[96]), .A2(c[96]), .Z(N96) );
  OR2D0 C3269 ( .A1(g[96]), .A2(N96), .Z(c[97]) );
  AN2D0 C3268 ( .A1(p[95]), .A2(c[95]), .Z(N95) );
  OR2D0 C3267 ( .A1(g[95]), .A2(N95), .Z(c[96]) );
  AN2D0 C3266 ( .A1(p[94]), .A2(c[94]), .Z(N94) );
  OR2D0 C3265 ( .A1(g[94]), .A2(N94), .Z(c[95]) );
  AN2D0 C3264 ( .A1(p[93]), .A2(c[93]), .Z(N93) );
  OR2D0 C3263 ( .A1(g[93]), .A2(N93), .Z(c[94]) );
  AN2D0 C3262 ( .A1(p[92]), .A2(c[92]), .Z(N92) );
  OR2D0 C3261 ( .A1(g[92]), .A2(N92), .Z(c[93]) );
  AN2D0 C3260 ( .A1(p[91]), .A2(c[91]), .Z(N91) );
  OR2D0 C3259 ( .A1(g[91]), .A2(N91), .Z(c[92]) );
  AN2D0 C3258 ( .A1(p[90]), .A2(c[90]), .Z(N90) );
  OR2D0 C3257 ( .A1(g[90]), .A2(N90), .Z(c[91]) );
  AN2D0 C3256 ( .A1(p[89]), .A2(c[89]), .Z(N89) );
  OR2D0 C3255 ( .A1(g[89]), .A2(N89), .Z(c[90]) );
  AN2D0 C3254 ( .A1(p[88]), .A2(c[88]), .Z(N88) );
  OR2D0 C3253 ( .A1(g[88]), .A2(N88), .Z(c[89]) );
  AN2D0 C3252 ( .A1(p[87]), .A2(c[87]), .Z(N87) );
  OR2D0 C3251 ( .A1(g[87]), .A2(N87), .Z(c[88]) );
  AN2D0 C3250 ( .A1(p[86]), .A2(c[86]), .Z(N86) );
  OR2D0 C3249 ( .A1(g[86]), .A2(N86), .Z(c[87]) );
  AN2D0 C3248 ( .A1(p[85]), .A2(c[85]), .Z(N85) );
  OR2D0 C3247 ( .A1(g[85]), .A2(N85), .Z(c[86]) );
  AN2D0 C3246 ( .A1(p[84]), .A2(c[84]), .Z(N84) );
  OR2D0 C3245 ( .A1(g[84]), .A2(N84), .Z(c[85]) );
  AN2D0 C3244 ( .A1(p[83]), .A2(c[83]), .Z(N83) );
  OR2D0 C3243 ( .A1(g[83]), .A2(N83), .Z(c[84]) );
  AN2D0 C3242 ( .A1(p[82]), .A2(c[82]), .Z(N82) );
  OR2D0 C3241 ( .A1(g[82]), .A2(N82), .Z(c[83]) );
  AN2D0 C3240 ( .A1(p[81]), .A2(c[81]), .Z(N81) );
  OR2D0 C3239 ( .A1(g[81]), .A2(N81), .Z(c[82]) );
  AN2D0 C3238 ( .A1(p[80]), .A2(c[80]), .Z(N80) );
  OR2D0 C3237 ( .A1(g[80]), .A2(N80), .Z(c[81]) );
  AN2D0 C3236 ( .A1(p[79]), .A2(c[79]), .Z(N79) );
  OR2D0 C3235 ( .A1(g[79]), .A2(N79), .Z(c[80]) );
  AN2D0 C3234 ( .A1(p[78]), .A2(c[78]), .Z(N78) );
  OR2D0 C3233 ( .A1(g[78]), .A2(N78), .Z(c[79]) );
  AN2D0 C3232 ( .A1(p[77]), .A2(c[77]), .Z(N77) );
  OR2D0 C3231 ( .A1(g[77]), .A2(N77), .Z(c[78]) );
  AN2D0 C3230 ( .A1(p[76]), .A2(c[76]), .Z(N76) );
  OR2D0 C3229 ( .A1(g[76]), .A2(N76), .Z(c[77]) );
  AN2D0 C3228 ( .A1(p[75]), .A2(c[75]), .Z(N75) );
  OR2D0 C3227 ( .A1(g[75]), .A2(N75), .Z(c[76]) );
  AN2D0 C3226 ( .A1(p[74]), .A2(c[74]), .Z(N74) );
  OR2D0 C3225 ( .A1(g[74]), .A2(N74), .Z(c[75]) );
  AN2D0 C3224 ( .A1(p[73]), .A2(c[73]), .Z(N73) );
  OR2D0 C3223 ( .A1(g[73]), .A2(N73), .Z(c[74]) );
  AN2D0 C3222 ( .A1(p[72]), .A2(c[72]), .Z(N72) );
  OR2D0 C3221 ( .A1(g[72]), .A2(N72), .Z(c[73]) );
  AN2D0 C3220 ( .A1(p[71]), .A2(c[71]), .Z(N71) );
  OR2D0 C3219 ( .A1(g[71]), .A2(N71), .Z(c[72]) );
  AN2D0 C3218 ( .A1(p[70]), .A2(c[70]), .Z(N70) );
  OR2D0 C3217 ( .A1(g[70]), .A2(N70), .Z(c[71]) );
  AN2D0 C3216 ( .A1(p[69]), .A2(c[69]), .Z(N69) );
  OR2D0 C3215 ( .A1(g[69]), .A2(N69), .Z(c[70]) );
  AN2D0 C3214 ( .A1(p[68]), .A2(c[68]), .Z(N68) );
  OR2D0 C3213 ( .A1(g[68]), .A2(N68), .Z(c[69]) );
  AN2D0 C3212 ( .A1(p[67]), .A2(c[67]), .Z(N67) );
  OR2D0 C3211 ( .A1(g[67]), .A2(N67), .Z(c[68]) );
  AN2D0 C3210 ( .A1(p[66]), .A2(c[66]), .Z(N66) );
  OR2D0 C3209 ( .A1(g[66]), .A2(N66), .Z(c[67]) );
  AN2D0 C3208 ( .A1(p[65]), .A2(c[65]), .Z(N65) );
  OR2D0 C3207 ( .A1(g[65]), .A2(N65), .Z(c[66]) );
  AN2D0 C3206 ( .A1(p[64]), .A2(c[64]), .Z(N64) );
  OR2D0 C3205 ( .A1(g[64]), .A2(N64), .Z(c[65]) );
  AN2D0 C3204 ( .A1(p[63]), .A2(c[63]), .Z(N63) );
  OR2D0 C3203 ( .A1(g[63]), .A2(N63), .Z(c[64]) );
  AN2D0 C3202 ( .A1(p[62]), .A2(c[62]), .Z(N62) );
  OR2D0 C3201 ( .A1(g[62]), .A2(N62), .Z(c[63]) );
  AN2D0 C3200 ( .A1(p[61]), .A2(c[61]), .Z(N61) );
  OR2D0 C3199 ( .A1(g[61]), .A2(N61), .Z(c[62]) );
  AN2D0 C3198 ( .A1(p[60]), .A2(c[60]), .Z(N60) );
  OR2D0 C3197 ( .A1(g[60]), .A2(N60), .Z(c[61]) );
  AN2D0 C3196 ( .A1(p[59]), .A2(c[59]), .Z(N59) );
  OR2D0 C3195 ( .A1(g[59]), .A2(N59), .Z(c[60]) );
  AN2D0 C3194 ( .A1(p[58]), .A2(c[58]), .Z(N58) );
  OR2D0 C3193 ( .A1(g[58]), .A2(N58), .Z(c[59]) );
  AN2D0 C3192 ( .A1(p[57]), .A2(c[57]), .Z(N57) );
  OR2D0 C3191 ( .A1(g[57]), .A2(N57), .Z(c[58]) );
  AN2D0 C3190 ( .A1(p[56]), .A2(c[56]), .Z(N56) );
  OR2D0 C3189 ( .A1(g[56]), .A2(N56), .Z(c[57]) );
  AN2D0 C3188 ( .A1(p[55]), .A2(c[55]), .Z(N55) );
  OR2D0 C3187 ( .A1(g[55]), .A2(N55), .Z(c[56]) );
  AN2D0 C3186 ( .A1(p[54]), .A2(c[54]), .Z(N54) );
  OR2D0 C3185 ( .A1(g[54]), .A2(N54), .Z(c[55]) );
  AN2D0 C3184 ( .A1(p[53]), .A2(c[53]), .Z(N53) );
  OR2D0 C3183 ( .A1(g[53]), .A2(N53), .Z(c[54]) );
  AN2D0 C3182 ( .A1(p[52]), .A2(c[52]), .Z(N52) );
  OR2D0 C3181 ( .A1(g[52]), .A2(N52), .Z(c[53]) );
  AN2D0 C3180 ( .A1(p[51]), .A2(c[51]), .Z(N51) );
  OR2D0 C3179 ( .A1(g[51]), .A2(N51), .Z(c[52]) );
  AN2D0 C3178 ( .A1(p[50]), .A2(c[50]), .Z(N50) );
  OR2D0 C3177 ( .A1(g[50]), .A2(N50), .Z(c[51]) );
  AN2D0 C3176 ( .A1(p[49]), .A2(c[49]), .Z(N49) );
  OR2D0 C3175 ( .A1(g[49]), .A2(N49), .Z(c[50]) );
  AN2D0 C3174 ( .A1(p[48]), .A2(c[48]), .Z(N48) );
  OR2D0 C3173 ( .A1(g[48]), .A2(N48), .Z(c[49]) );
  AN2D0 C3172 ( .A1(p[47]), .A2(c[47]), .Z(N47) );
  OR2D0 C3171 ( .A1(g[47]), .A2(N47), .Z(c[48]) );
  AN2D0 C3170 ( .A1(p[46]), .A2(c[46]), .Z(N46) );
  OR2D0 C3169 ( .A1(g[46]), .A2(N46), .Z(c[47]) );
  AN2D0 C3168 ( .A1(p[45]), .A2(c[45]), .Z(N45) );
  OR2D0 C3167 ( .A1(g[45]), .A2(N45), .Z(c[46]) );
  AN2D0 C3166 ( .A1(p[44]), .A2(c[44]), .Z(N44) );
  OR2D0 C3165 ( .A1(g[44]), .A2(N44), .Z(c[45]) );
  AN2D0 C3164 ( .A1(p[43]), .A2(c[43]), .Z(N43) );
  OR2D0 C3163 ( .A1(g[43]), .A2(N43), .Z(c[44]) );
  AN2D0 C3162 ( .A1(p[42]), .A2(c[42]), .Z(N42) );
  OR2D0 C3161 ( .A1(g[42]), .A2(N42), .Z(c[43]) );
  AN2D0 C3160 ( .A1(p[41]), .A2(c[41]), .Z(N41) );
  OR2D0 C3159 ( .A1(g[41]), .A2(N41), .Z(c[42]) );
  AN2D0 C3158 ( .A1(p[40]), .A2(c[40]), .Z(N40) );
  OR2D0 C3157 ( .A1(g[40]), .A2(N40), .Z(c[41]) );
  AN2D0 C3156 ( .A1(p[39]), .A2(c[39]), .Z(N39) );
  OR2D0 C3155 ( .A1(g[39]), .A2(N39), .Z(c[40]) );
  AN2D0 C3154 ( .A1(p[38]), .A2(c[38]), .Z(N38) );
  OR2D0 C3153 ( .A1(g[38]), .A2(N38), .Z(c[39]) );
  AN2D0 C3152 ( .A1(p[37]), .A2(c[37]), .Z(N37) );
  OR2D0 C3151 ( .A1(g[37]), .A2(N37), .Z(c[38]) );
  AN2D0 C3150 ( .A1(p[36]), .A2(c[36]), .Z(N36) );
  OR2D0 C3149 ( .A1(g[36]), .A2(N36), .Z(c[37]) );
  AN2D0 C3148 ( .A1(p[35]), .A2(c[35]), .Z(N35) );
  OR2D0 C3147 ( .A1(g[35]), .A2(N35), .Z(c[36]) );
  AN2D0 C3146 ( .A1(p[34]), .A2(c[34]), .Z(N34) );
  OR2D0 C3145 ( .A1(g[34]), .A2(N34), .Z(c[35]) );
  AN2D0 C3144 ( .A1(p[33]), .A2(c[33]), .Z(N33) );
  OR2D0 C3143 ( .A1(g[33]), .A2(N33), .Z(c[34]) );
  AN2D0 C3142 ( .A1(p[32]), .A2(c[32]), .Z(N32) );
  OR2D0 C3141 ( .A1(g[32]), .A2(N32), .Z(c[33]) );
  AN2D0 C3140 ( .A1(p[31]), .A2(c[31]), .Z(N31) );
  OR2D0 C3139 ( .A1(g[31]), .A2(N31), .Z(c[32]) );
  AN2D0 C3138 ( .A1(p[30]), .A2(c[30]), .Z(N30) );
  OR2D0 C3137 ( .A1(g[30]), .A2(N30), .Z(c[31]) );
  AN2D0 C3136 ( .A1(p[29]), .A2(c[29]), .Z(N29) );
  OR2D0 C3135 ( .A1(g[29]), .A2(N29), .Z(c[30]) );
  AN2D0 C3134 ( .A1(p[28]), .A2(c[28]), .Z(N28) );
  OR2D0 C3133 ( .A1(g[28]), .A2(N28), .Z(c[29]) );
  AN2D0 C3132 ( .A1(p[27]), .A2(c[27]), .Z(N27) );
  OR2D0 C3131 ( .A1(g[27]), .A2(N27), .Z(c[28]) );
  AN2D0 C3130 ( .A1(p[26]), .A2(c[26]), .Z(N26) );
  OR2D0 C3129 ( .A1(g[26]), .A2(N26), .Z(c[27]) );
  AN2D0 C3128 ( .A1(p[25]), .A2(c[25]), .Z(N25) );
  OR2D0 C3127 ( .A1(g[25]), .A2(N25), .Z(c[26]) );
  AN2D0 C3126 ( .A1(p[24]), .A2(c[24]), .Z(N24) );
  OR2D0 C3125 ( .A1(g[24]), .A2(N24), .Z(c[25]) );
  AN2D0 C3124 ( .A1(p[23]), .A2(c[23]), .Z(N23) );
  OR2D0 C3123 ( .A1(g[23]), .A2(N23), .Z(c[24]) );
  AN2D0 C3122 ( .A1(p[22]), .A2(c[22]), .Z(N22) );
  OR2D0 C3121 ( .A1(g[22]), .A2(N22), .Z(c[23]) );
  AN2D0 C3120 ( .A1(p[21]), .A2(c[21]), .Z(N21) );
  OR2D0 C3119 ( .A1(g[21]), .A2(N21), .Z(c[22]) );
  AN2D0 C3118 ( .A1(p[20]), .A2(c[20]), .Z(N20) );
  OR2D0 C3117 ( .A1(g[20]), .A2(N20), .Z(c[21]) );
  AN2D0 C3116 ( .A1(p[19]), .A2(c[19]), .Z(N19) );
  OR2D0 C3115 ( .A1(g[19]), .A2(N19), .Z(c[20]) );
  AN2D0 C3114 ( .A1(p[18]), .A2(c[18]), .Z(N18) );
  OR2D0 C3113 ( .A1(g[18]), .A2(N18), .Z(c[19]) );
  AN2D0 C3112 ( .A1(p[17]), .A2(c[17]), .Z(N17) );
  OR2D0 C3111 ( .A1(g[17]), .A2(N17), .Z(c[18]) );
  AN2D0 C3110 ( .A1(p[16]), .A2(c[16]), .Z(N16) );
  OR2D0 C3109 ( .A1(g[16]), .A2(N16), .Z(c[17]) );
  AN2D0 C3108 ( .A1(p[15]), .A2(c[15]), .Z(N15) );
  OR2D0 C3107 ( .A1(g[15]), .A2(N15), .Z(c[16]) );
  AN2D0 C3106 ( .A1(p[14]), .A2(c[14]), .Z(N14) );
  OR2D0 C3105 ( .A1(g[14]), .A2(N14), .Z(c[15]) );
  AN2D0 C3104 ( .A1(p[13]), .A2(c[13]), .Z(N13) );
  OR2D0 C3103 ( .A1(g[13]), .A2(N13), .Z(c[14]) );
  AN2D0 C3102 ( .A1(p[12]), .A2(c[12]), .Z(N12) );
  OR2D0 C3101 ( .A1(g[12]), .A2(N12), .Z(c[13]) );
  AN2D0 C3100 ( .A1(p[11]), .A2(c[11]), .Z(N11) );
  OR2D0 C3099 ( .A1(g[11]), .A2(N11), .Z(c[12]) );
  AN2D0 C3098 ( .A1(p[10]), .A2(c[10]), .Z(N10) );
  OR2D0 C3097 ( .A1(g[10]), .A2(N10), .Z(c[11]) );
  AN2D0 C3096 ( .A1(p[9]), .A2(c[9]), .Z(N9) );
  OR2D0 C3095 ( .A1(g[9]), .A2(N9), .Z(c[10]) );
  AN2D0 C3094 ( .A1(p[8]), .A2(c[8]), .Z(N8) );
  OR2D0 C3093 ( .A1(g[8]), .A2(N8), .Z(c[9]) );
  AN2D0 C3092 ( .A1(p[7]), .A2(c[7]), .Z(N7) );
  OR2D0 C3091 ( .A1(g[7]), .A2(N7), .Z(c[8]) );
  AN2D0 C3090 ( .A1(p[6]), .A2(c[6]), .Z(N6) );
  OR2D0 C3089 ( .A1(g[6]), .A2(N6), .Z(c[7]) );
  AN2D0 C3088 ( .A1(p[5]), .A2(c[5]), .Z(N5) );
  OR2D0 C3087 ( .A1(g[5]), .A2(N5), .Z(c[6]) );
  AN2D0 C3086 ( .A1(p[4]), .A2(c[4]), .Z(N4) );
  OR2D0 C3085 ( .A1(g[4]), .A2(N4), .Z(c[5]) );
  AN2D0 C3084 ( .A1(p[3]), .A2(c[3]), .Z(N3) );
  OR2D0 C3083 ( .A1(g[3]), .A2(N3), .Z(c[4]) );
  AN2D0 C3082 ( .A1(p[2]), .A2(c[2]), .Z(N2) );
  OR2D0 C3081 ( .A1(g[2]), .A2(N2), .Z(c[3]) );
  AN2D0 C3080 ( .A1(p[1]), .A2(c[1]), .Z(N1) );
  OR2D0 C3079 ( .A1(g[1]), .A2(N1), .Z(c[2]) );
  AN2D0 C3078 ( .A1(p[0]), .A2(cin), .Z(N0) );
  OR2D0 C3077 ( .A1(g[0]), .A2(N0), .Z(c[1]) );
  XOR2D0 C3076 ( .A1(a[0]), .A2(b[0]), .Z(p[0]) );
  XOR2D0 C3075 ( .A1(a[1]), .A2(b[1]), .Z(p[1]) );
  XOR2D0 C3074 ( .A1(a[2]), .A2(b[2]), .Z(p[2]) );
  XOR2D0 C3073 ( .A1(a[3]), .A2(b[3]), .Z(p[3]) );
  XOR2D0 C3072 ( .A1(a[4]), .A2(b[4]), .Z(p[4]) );
  XOR2D0 C3071 ( .A1(a[5]), .A2(b[5]), .Z(p[5]) );
  XOR2D0 C3070 ( .A1(a[6]), .A2(b[6]), .Z(p[6]) );
  XOR2D0 C3069 ( .A1(a[7]), .A2(b[7]), .Z(p[7]) );
  XOR2D0 C3068 ( .A1(a[8]), .A2(b[8]), .Z(p[8]) );
  XOR2D0 C3067 ( .A1(a[9]), .A2(b[9]), .Z(p[9]) );
  XOR2D0 C3066 ( .A1(a[10]), .A2(b[10]), .Z(p[10]) );
  XOR2D0 C3065 ( .A1(a[11]), .A2(b[11]), .Z(p[11]) );
  XOR2D0 C3064 ( .A1(a[12]), .A2(b[12]), .Z(p[12]) );
  XOR2D0 C3063 ( .A1(a[13]), .A2(b[13]), .Z(p[13]) );
  XOR2D0 C3062 ( .A1(a[14]), .A2(b[14]), .Z(p[14]) );
  XOR2D0 C3061 ( .A1(a[15]), .A2(b[15]), .Z(p[15]) );
  XOR2D0 C3060 ( .A1(a[16]), .A2(b[16]), .Z(p[16]) );
  XOR2D0 C3059 ( .A1(a[17]), .A2(b[17]), .Z(p[17]) );
  XOR2D0 C3058 ( .A1(a[18]), .A2(b[18]), .Z(p[18]) );
  XOR2D0 C3057 ( .A1(a[19]), .A2(b[19]), .Z(p[19]) );
  XOR2D0 C3056 ( .A1(a[20]), .A2(b[20]), .Z(p[20]) );
  XOR2D0 C3055 ( .A1(a[21]), .A2(b[21]), .Z(p[21]) );
  XOR2D0 C3054 ( .A1(a[22]), .A2(b[22]), .Z(p[22]) );
  XOR2D0 C3053 ( .A1(a[23]), .A2(b[23]), .Z(p[23]) );
  XOR2D0 C3052 ( .A1(a[24]), .A2(b[24]), .Z(p[24]) );
  XOR2D0 C3051 ( .A1(a[25]), .A2(b[25]), .Z(p[25]) );
  XOR2D0 C3050 ( .A1(a[26]), .A2(b[26]), .Z(p[26]) );
  XOR2D0 C3049 ( .A1(a[27]), .A2(b[27]), .Z(p[27]) );
  XOR2D0 C3048 ( .A1(a[28]), .A2(b[28]), .Z(p[28]) );
  XOR2D0 C3047 ( .A1(a[29]), .A2(b[29]), .Z(p[29]) );
  XOR2D0 C3046 ( .A1(a[30]), .A2(b[30]), .Z(p[30]) );
  XOR2D0 C3045 ( .A1(a[31]), .A2(b[31]), .Z(p[31]) );
  XOR2D0 C3044 ( .A1(a[32]), .A2(b[32]), .Z(p[32]) );
  XOR2D0 C3043 ( .A1(a[33]), .A2(b[33]), .Z(p[33]) );
  XOR2D0 C3042 ( .A1(a[34]), .A2(b[34]), .Z(p[34]) );
  XOR2D0 C3041 ( .A1(a[35]), .A2(b[35]), .Z(p[35]) );
  XOR2D0 C3040 ( .A1(a[36]), .A2(b[36]), .Z(p[36]) );
  XOR2D0 C3039 ( .A1(a[37]), .A2(b[37]), .Z(p[37]) );
  XOR2D0 C3038 ( .A1(a[38]), .A2(b[38]), .Z(p[38]) );
  XOR2D0 C3037 ( .A1(a[39]), .A2(b[39]), .Z(p[39]) );
  XOR2D0 C3036 ( .A1(a[40]), .A2(b[40]), .Z(p[40]) );
  XOR2D0 C3035 ( .A1(a[41]), .A2(b[41]), .Z(p[41]) );
  XOR2D0 C3034 ( .A1(a[42]), .A2(b[42]), .Z(p[42]) );
  XOR2D0 C3033 ( .A1(a[43]), .A2(b[43]), .Z(p[43]) );
  XOR2D0 C3032 ( .A1(a[44]), .A2(b[44]), .Z(p[44]) );
  XOR2D0 C3031 ( .A1(a[45]), .A2(b[45]), .Z(p[45]) );
  XOR2D0 C3030 ( .A1(a[46]), .A2(b[46]), .Z(p[46]) );
  XOR2D0 C3029 ( .A1(a[47]), .A2(b[47]), .Z(p[47]) );
  XOR2D0 C3028 ( .A1(a[48]), .A2(b[48]), .Z(p[48]) );
  XOR2D0 C3027 ( .A1(a[49]), .A2(b[49]), .Z(p[49]) );
  XOR2D0 C3026 ( .A1(a[50]), .A2(b[50]), .Z(p[50]) );
  XOR2D0 C3025 ( .A1(a[51]), .A2(b[51]), .Z(p[51]) );
  XOR2D0 C3024 ( .A1(a[52]), .A2(b[52]), .Z(p[52]) );
  XOR2D0 C3023 ( .A1(a[53]), .A2(b[53]), .Z(p[53]) );
  XOR2D0 C3022 ( .A1(a[54]), .A2(b[54]), .Z(p[54]) );
  XOR2D0 C3021 ( .A1(a[55]), .A2(b[55]), .Z(p[55]) );
  XOR2D0 C3020 ( .A1(a[56]), .A2(b[56]), .Z(p[56]) );
  XOR2D0 C3019 ( .A1(a[57]), .A2(b[57]), .Z(p[57]) );
  XOR2D0 C3018 ( .A1(a[58]), .A2(b[58]), .Z(p[58]) );
  XOR2D0 C3017 ( .A1(a[59]), .A2(b[59]), .Z(p[59]) );
  XOR2D0 C3016 ( .A1(a[60]), .A2(b[60]), .Z(p[60]) );
  XOR2D0 C3015 ( .A1(a[61]), .A2(b[61]), .Z(p[61]) );
  XOR2D0 C3014 ( .A1(a[62]), .A2(b[62]), .Z(p[62]) );
  XOR2D0 C3013 ( .A1(a[63]), .A2(b[63]), .Z(p[63]) );
  XOR2D0 C3012 ( .A1(a[64]), .A2(b[64]), .Z(p[64]) );
  XOR2D0 C3011 ( .A1(a[65]), .A2(b[65]), .Z(p[65]) );
  XOR2D0 C3010 ( .A1(a[66]), .A2(b[66]), .Z(p[66]) );
  XOR2D0 C3009 ( .A1(a[67]), .A2(b[67]), .Z(p[67]) );
  XOR2D0 C3008 ( .A1(a[68]), .A2(b[68]), .Z(p[68]) );
  XOR2D0 C3007 ( .A1(a[69]), .A2(b[69]), .Z(p[69]) );
  XOR2D0 C3006 ( .A1(a[70]), .A2(b[70]), .Z(p[70]) );
  XOR2D0 C3005 ( .A1(a[71]), .A2(b[71]), .Z(p[71]) );
  XOR2D0 C3004 ( .A1(a[72]), .A2(b[72]), .Z(p[72]) );
  XOR2D0 C3003 ( .A1(a[73]), .A2(b[73]), .Z(p[73]) );
  XOR2D0 C3002 ( .A1(a[74]), .A2(b[74]), .Z(p[74]) );
  XOR2D0 C3001 ( .A1(a[75]), .A2(b[75]), .Z(p[75]) );
  XOR2D0 C3000 ( .A1(a[76]), .A2(b[76]), .Z(p[76]) );
  XOR2D0 C2999 ( .A1(a[77]), .A2(b[77]), .Z(p[77]) );
  XOR2D0 C2998 ( .A1(a[78]), .A2(b[78]), .Z(p[78]) );
  XOR2D0 C2997 ( .A1(a[79]), .A2(b[79]), .Z(p[79]) );
  XOR2D0 C2996 ( .A1(a[80]), .A2(b[80]), .Z(p[80]) );
  XOR2D0 C2995 ( .A1(a[81]), .A2(b[81]), .Z(p[81]) );
  XOR2D0 C2994 ( .A1(a[82]), .A2(b[82]), .Z(p[82]) );
  XOR2D0 C2993 ( .A1(a[83]), .A2(b[83]), .Z(p[83]) );
  XOR2D0 C2992 ( .A1(a[84]), .A2(b[84]), .Z(p[84]) );
  XOR2D0 C2991 ( .A1(a[85]), .A2(b[85]), .Z(p[85]) );
  XOR2D0 C2990 ( .A1(a[86]), .A2(b[86]), .Z(p[86]) );
  XOR2D0 C2989 ( .A1(a[87]), .A2(b[87]), .Z(p[87]) );
  XOR2D0 C2988 ( .A1(a[88]), .A2(b[88]), .Z(p[88]) );
  XOR2D0 C2987 ( .A1(a[89]), .A2(b[89]), .Z(p[89]) );
  XOR2D0 C2986 ( .A1(a[90]), .A2(b[90]), .Z(p[90]) );
  XOR2D0 C2985 ( .A1(a[91]), .A2(b[91]), .Z(p[91]) );
  XOR2D0 C2984 ( .A1(a[92]), .A2(b[92]), .Z(p[92]) );
  XOR2D0 C2983 ( .A1(a[93]), .A2(b[93]), .Z(p[93]) );
  XOR2D0 C2982 ( .A1(a[94]), .A2(b[94]), .Z(p[94]) );
  XOR2D0 C2981 ( .A1(a[95]), .A2(b[95]), .Z(p[95]) );
  XOR2D0 C2980 ( .A1(a[96]), .A2(b[96]), .Z(p[96]) );
  XOR2D0 C2979 ( .A1(a[97]), .A2(b[97]), .Z(p[97]) );
  XOR2D0 C2978 ( .A1(a[98]), .A2(b[98]), .Z(p[98]) );
  XOR2D0 C2977 ( .A1(a[99]), .A2(b[99]), .Z(p[99]) );
  XOR2D0 C2976 ( .A1(a[100]), .A2(b[100]), .Z(p[100]) );
  XOR2D0 C2975 ( .A1(a[101]), .A2(b[101]), .Z(p[101]) );
  XOR2D0 C2974 ( .A1(a[102]), .A2(b[102]), .Z(p[102]) );
  XOR2D0 C2973 ( .A1(a[103]), .A2(b[103]), .Z(p[103]) );
  XOR2D0 C2972 ( .A1(a[104]), .A2(b[104]), .Z(p[104]) );
  XOR2D0 C2971 ( .A1(a[105]), .A2(b[105]), .Z(p[105]) );
  XOR2D0 C2970 ( .A1(a[106]), .A2(b[106]), .Z(p[106]) );
  XOR2D0 C2969 ( .A1(a[107]), .A2(b[107]), .Z(p[107]) );
  XOR2D0 C2968 ( .A1(a[108]), .A2(b[108]), .Z(p[108]) );
  XOR2D0 C2967 ( .A1(a[109]), .A2(b[109]), .Z(p[109]) );
  XOR2D0 C2966 ( .A1(a[110]), .A2(b[110]), .Z(p[110]) );
  XOR2D0 C2965 ( .A1(a[111]), .A2(b[111]), .Z(p[111]) );
  XOR2D0 C2964 ( .A1(a[112]), .A2(b[112]), .Z(p[112]) );
  XOR2D0 C2963 ( .A1(a[113]), .A2(b[113]), .Z(p[113]) );
  XOR2D0 C2962 ( .A1(a[114]), .A2(b[114]), .Z(p[114]) );
  XOR2D0 C2961 ( .A1(a[115]), .A2(b[115]), .Z(p[115]) );
  XOR2D0 C2960 ( .A1(a[116]), .A2(b[116]), .Z(p[116]) );
  XOR2D0 C2959 ( .A1(a[117]), .A2(b[117]), .Z(p[117]) );
  XOR2D0 C2958 ( .A1(a[118]), .A2(b[118]), .Z(p[118]) );
  XOR2D0 C2957 ( .A1(a[119]), .A2(b[119]), .Z(p[119]) );
  XOR2D0 C2956 ( .A1(a[120]), .A2(b[120]), .Z(p[120]) );
  XOR2D0 C2955 ( .A1(a[121]), .A2(b[121]), .Z(p[121]) );
  XOR2D0 C2954 ( .A1(a[122]), .A2(b[122]), .Z(p[122]) );
  XOR2D0 C2953 ( .A1(a[123]), .A2(b[123]), .Z(p[123]) );
  XOR2D0 C2952 ( .A1(a[124]), .A2(b[124]), .Z(p[124]) );
  XOR2D0 C2951 ( .A1(a[125]), .A2(b[125]), .Z(p[125]) );
  XOR2D0 C2950 ( .A1(a[126]), .A2(b[126]), .Z(p[126]) );
  XOR2D0 C2949 ( .A1(a[127]), .A2(b[127]), .Z(p[127]) );
  XOR2D0 C2948 ( .A1(a[128]), .A2(b[128]), .Z(p[128]) );
  XOR2D0 C2947 ( .A1(a[129]), .A2(b[129]), .Z(p[129]) );
  XOR2D0 C2946 ( .A1(a[130]), .A2(b[130]), .Z(p[130]) );
  XOR2D0 C2945 ( .A1(a[131]), .A2(b[131]), .Z(p[131]) );
  XOR2D0 C2944 ( .A1(a[132]), .A2(b[132]), .Z(p[132]) );
  XOR2D0 C2943 ( .A1(a[133]), .A2(b[133]), .Z(p[133]) );
  XOR2D0 C2942 ( .A1(a[134]), .A2(b[134]), .Z(p[134]) );
  XOR2D0 C2941 ( .A1(a[135]), .A2(b[135]), .Z(p[135]) );
  XOR2D0 C2940 ( .A1(a[136]), .A2(b[136]), .Z(p[136]) );
  XOR2D0 C2939 ( .A1(a[137]), .A2(b[137]), .Z(p[137]) );
  XOR2D0 C2938 ( .A1(a[138]), .A2(b[138]), .Z(p[138]) );
  XOR2D0 C2937 ( .A1(a[139]), .A2(b[139]), .Z(p[139]) );
  XOR2D0 C2936 ( .A1(a[140]), .A2(b[140]), .Z(p[140]) );
  XOR2D0 C2935 ( .A1(a[141]), .A2(b[141]), .Z(p[141]) );
  XOR2D0 C2934 ( .A1(a[142]), .A2(b[142]), .Z(p[142]) );
  XOR2D0 C2933 ( .A1(a[143]), .A2(b[143]), .Z(p[143]) );
  XOR2D0 C2932 ( .A1(a[144]), .A2(b[144]), .Z(p[144]) );
  XOR2D0 C2931 ( .A1(a[145]), .A2(b[145]), .Z(p[145]) );
  XOR2D0 C2930 ( .A1(a[146]), .A2(b[146]), .Z(p[146]) );
  XOR2D0 C2929 ( .A1(a[147]), .A2(b[147]), .Z(p[147]) );
  XOR2D0 C2928 ( .A1(a[148]), .A2(b[148]), .Z(p[148]) );
  XOR2D0 C2927 ( .A1(a[149]), .A2(b[149]), .Z(p[149]) );
  XOR2D0 C2926 ( .A1(a[150]), .A2(b[150]), .Z(p[150]) );
  XOR2D0 C2925 ( .A1(a[151]), .A2(b[151]), .Z(p[151]) );
  XOR2D0 C2924 ( .A1(a[152]), .A2(b[152]), .Z(p[152]) );
  XOR2D0 C2923 ( .A1(a[153]), .A2(b[153]), .Z(p[153]) );
  XOR2D0 C2922 ( .A1(a[154]), .A2(b[154]), .Z(p[154]) );
  XOR2D0 C2921 ( .A1(a[155]), .A2(b[155]), .Z(p[155]) );
  XOR2D0 C2920 ( .A1(a[156]), .A2(b[156]), .Z(p[156]) );
  XOR2D0 C2919 ( .A1(a[157]), .A2(b[157]), .Z(p[157]) );
  XOR2D0 C2918 ( .A1(a[158]), .A2(b[158]), .Z(p[158]) );
  XOR2D0 C2917 ( .A1(a[159]), .A2(b[159]), .Z(p[159]) );
  XOR2D0 C2916 ( .A1(a[160]), .A2(b[160]), .Z(p[160]) );
  XOR2D0 C2915 ( .A1(a[161]), .A2(b[161]), .Z(p[161]) );
  XOR2D0 C2914 ( .A1(a[162]), .A2(b[162]), .Z(p[162]) );
  XOR2D0 C2913 ( .A1(a[163]), .A2(b[163]), .Z(p[163]) );
  XOR2D0 C2912 ( .A1(a[164]), .A2(b[164]), .Z(p[164]) );
  XOR2D0 C2911 ( .A1(a[165]), .A2(b[165]), .Z(p[165]) );
  XOR2D0 C2910 ( .A1(a[166]), .A2(b[166]), .Z(p[166]) );
  XOR2D0 C2909 ( .A1(a[167]), .A2(b[167]), .Z(p[167]) );
  XOR2D0 C2908 ( .A1(a[168]), .A2(b[168]), .Z(p[168]) );
  XOR2D0 C2907 ( .A1(a[169]), .A2(b[169]), .Z(p[169]) );
  XOR2D0 C2906 ( .A1(a[170]), .A2(b[170]), .Z(p[170]) );
  XOR2D0 C2905 ( .A1(a[171]), .A2(b[171]), .Z(p[171]) );
  XOR2D0 C2904 ( .A1(a[172]), .A2(b[172]), .Z(p[172]) );
  XOR2D0 C2903 ( .A1(a[173]), .A2(b[173]), .Z(p[173]) );
  XOR2D0 C2902 ( .A1(a[174]), .A2(b[174]), .Z(p[174]) );
  XOR2D0 C2901 ( .A1(a[175]), .A2(b[175]), .Z(p[175]) );
  XOR2D0 C2900 ( .A1(a[176]), .A2(b[176]), .Z(p[176]) );
  XOR2D0 C2899 ( .A1(a[177]), .A2(b[177]), .Z(p[177]) );
  XOR2D0 C2898 ( .A1(a[178]), .A2(b[178]), .Z(p[178]) );
  XOR2D0 C2897 ( .A1(a[179]), .A2(b[179]), .Z(p[179]) );
  XOR2D0 C2896 ( .A1(a[180]), .A2(b[180]), .Z(p[180]) );
  XOR2D0 C2895 ( .A1(a[181]), .A2(b[181]), .Z(p[181]) );
  XOR2D0 C2894 ( .A1(a[182]), .A2(b[182]), .Z(p[182]) );
  XOR2D0 C2893 ( .A1(a[183]), .A2(b[183]), .Z(p[183]) );
  XOR2D0 C2892 ( .A1(a[184]), .A2(b[184]), .Z(p[184]) );
  XOR2D0 C2891 ( .A1(a[185]), .A2(b[185]), .Z(p[185]) );
  XOR2D0 C2890 ( .A1(a[186]), .A2(b[186]), .Z(p[186]) );
  XOR2D0 C2889 ( .A1(a[187]), .A2(b[187]), .Z(p[187]) );
  XOR2D0 C2888 ( .A1(a[188]), .A2(b[188]), .Z(p[188]) );
  XOR2D0 C2887 ( .A1(a[189]), .A2(b[189]), .Z(p[189]) );
  XOR2D0 C2886 ( .A1(a[190]), .A2(b[190]), .Z(p[190]) );
  XOR2D0 C2885 ( .A1(a[191]), .A2(b[191]), .Z(p[191]) );
  XOR2D0 C2884 ( .A1(a[192]), .A2(b[192]), .Z(p[192]) );
  XOR2D0 C2883 ( .A1(a[193]), .A2(b[193]), .Z(p[193]) );
  XOR2D0 C2882 ( .A1(a[194]), .A2(b[194]), .Z(p[194]) );
  XOR2D0 C2881 ( .A1(a[195]), .A2(b[195]), .Z(p[195]) );
  XOR2D0 C2880 ( .A1(a[196]), .A2(b[196]), .Z(p[196]) );
  XOR2D0 C2879 ( .A1(a[197]), .A2(b[197]), .Z(p[197]) );
  XOR2D0 C2878 ( .A1(a[198]), .A2(b[198]), .Z(p[198]) );
  XOR2D0 C2877 ( .A1(a[199]), .A2(b[199]), .Z(p[199]) );
  XOR2D0 C2876 ( .A1(a[200]), .A2(b[200]), .Z(p[200]) );
  XOR2D0 C2875 ( .A1(a[201]), .A2(b[201]), .Z(p[201]) );
  XOR2D0 C2874 ( .A1(a[202]), .A2(b[202]), .Z(p[202]) );
  XOR2D0 C2873 ( .A1(a[203]), .A2(b[203]), .Z(p[203]) );
  XOR2D0 C2872 ( .A1(a[204]), .A2(b[204]), .Z(p[204]) );
  XOR2D0 C2871 ( .A1(a[205]), .A2(b[205]), .Z(p[205]) );
  XOR2D0 C2870 ( .A1(a[206]), .A2(b[206]), .Z(p[206]) );
  XOR2D0 C2869 ( .A1(a[207]), .A2(b[207]), .Z(p[207]) );
  XOR2D0 C2868 ( .A1(a[208]), .A2(b[208]), .Z(p[208]) );
  XOR2D0 C2867 ( .A1(a[209]), .A2(b[209]), .Z(p[209]) );
  XOR2D0 C2866 ( .A1(a[210]), .A2(b[210]), .Z(p[210]) );
  XOR2D0 C2865 ( .A1(a[211]), .A2(b[211]), .Z(p[211]) );
  XOR2D0 C2864 ( .A1(a[212]), .A2(b[212]), .Z(p[212]) );
  XOR2D0 C2863 ( .A1(a[213]), .A2(b[213]), .Z(p[213]) );
  XOR2D0 C2862 ( .A1(a[214]), .A2(b[214]), .Z(p[214]) );
  XOR2D0 C2861 ( .A1(a[215]), .A2(b[215]), .Z(p[215]) );
  XOR2D0 C2860 ( .A1(a[216]), .A2(b[216]), .Z(p[216]) );
  XOR2D0 C2859 ( .A1(a[217]), .A2(b[217]), .Z(p[217]) );
  XOR2D0 C2858 ( .A1(a[218]), .A2(b[218]), .Z(p[218]) );
  XOR2D0 C2857 ( .A1(a[219]), .A2(b[219]), .Z(p[219]) );
  XOR2D0 C2856 ( .A1(a[220]), .A2(b[220]), .Z(p[220]) );
  XOR2D0 C2855 ( .A1(a[221]), .A2(b[221]), .Z(p[221]) );
  XOR2D0 C2854 ( .A1(a[222]), .A2(b[222]), .Z(p[222]) );
  XOR2D0 C2853 ( .A1(a[223]), .A2(b[223]), .Z(p[223]) );
  XOR2D0 C2852 ( .A1(a[224]), .A2(b[224]), .Z(p[224]) );
  XOR2D0 C2851 ( .A1(a[225]), .A2(b[225]), .Z(p[225]) );
  XOR2D0 C2850 ( .A1(a[226]), .A2(b[226]), .Z(p[226]) );
  XOR2D0 C2849 ( .A1(a[227]), .A2(b[227]), .Z(p[227]) );
  XOR2D0 C2848 ( .A1(a[228]), .A2(b[228]), .Z(p[228]) );
  XOR2D0 C2847 ( .A1(a[229]), .A2(b[229]), .Z(p[229]) );
  XOR2D0 C2846 ( .A1(a[230]), .A2(b[230]), .Z(p[230]) );
  XOR2D0 C2845 ( .A1(a[231]), .A2(b[231]), .Z(p[231]) );
  XOR2D0 C2844 ( .A1(a[232]), .A2(b[232]), .Z(p[232]) );
  XOR2D0 C2843 ( .A1(a[233]), .A2(b[233]), .Z(p[233]) );
  XOR2D0 C2842 ( .A1(a[234]), .A2(b[234]), .Z(p[234]) );
  XOR2D0 C2841 ( .A1(a[235]), .A2(b[235]), .Z(p[235]) );
  XOR2D0 C2840 ( .A1(a[236]), .A2(b[236]), .Z(p[236]) );
  XOR2D0 C2839 ( .A1(a[237]), .A2(b[237]), .Z(p[237]) );
  XOR2D0 C2838 ( .A1(a[238]), .A2(b[238]), .Z(p[238]) );
  XOR2D0 C2837 ( .A1(a[239]), .A2(b[239]), .Z(p[239]) );
  XOR2D0 C2836 ( .A1(a[240]), .A2(b[240]), .Z(p[240]) );
  XOR2D0 C2835 ( .A1(a[241]), .A2(b[241]), .Z(p[241]) );
  XOR2D0 C2834 ( .A1(a[242]), .A2(b[242]), .Z(p[242]) );
  XOR2D0 C2833 ( .A1(a[243]), .A2(b[243]), .Z(p[243]) );
  XOR2D0 C2832 ( .A1(a[244]), .A2(b[244]), .Z(p[244]) );
  XOR2D0 C2831 ( .A1(a[245]), .A2(b[245]), .Z(p[245]) );
  XOR2D0 C2830 ( .A1(a[246]), .A2(b[246]), .Z(p[246]) );
  XOR2D0 C2829 ( .A1(a[247]), .A2(b[247]), .Z(p[247]) );
  XOR2D0 C2828 ( .A1(a[248]), .A2(b[248]), .Z(p[248]) );
  XOR2D0 C2827 ( .A1(a[249]), .A2(b[249]), .Z(p[249]) );
  XOR2D0 C2826 ( .A1(a[250]), .A2(b[250]), .Z(p[250]) );
  XOR2D0 C2825 ( .A1(a[251]), .A2(b[251]), .Z(p[251]) );
  XOR2D0 C2824 ( .A1(a[252]), .A2(b[252]), .Z(p[252]) );
  XOR2D0 C2823 ( .A1(a[253]), .A2(b[253]), .Z(p[253]) );
  XOR2D0 C2822 ( .A1(a[254]), .A2(b[254]), .Z(p[254]) );
  XOR2D0 C2821 ( .A1(a[255]), .A2(b[255]), .Z(p[255]) );
  XOR2D0 C2820 ( .A1(a[256]), .A2(b[256]), .Z(p[256]) );
  XOR2D0 C2819 ( .A1(a[257]), .A2(b[257]), .Z(p[257]) );
  XOR2D0 C2818 ( .A1(a[258]), .A2(b[258]), .Z(p[258]) );
  XOR2D0 C2817 ( .A1(a[259]), .A2(b[259]), .Z(p[259]) );
  XOR2D0 C2816 ( .A1(a[260]), .A2(b[260]), .Z(p[260]) );
  XOR2D0 C2815 ( .A1(a[261]), .A2(b[261]), .Z(p[261]) );
  XOR2D0 C2814 ( .A1(a[262]), .A2(b[262]), .Z(p[262]) );
  XOR2D0 C2813 ( .A1(a[263]), .A2(b[263]), .Z(p[263]) );
  XOR2D0 C2812 ( .A1(a[264]), .A2(b[264]), .Z(p[264]) );
  XOR2D0 C2811 ( .A1(a[265]), .A2(b[265]), .Z(p[265]) );
  XOR2D0 C2810 ( .A1(a[266]), .A2(b[266]), .Z(p[266]) );
  XOR2D0 C2809 ( .A1(a[267]), .A2(b[267]), .Z(p[267]) );
  XOR2D0 C2808 ( .A1(a[268]), .A2(b[268]), .Z(p[268]) );
  XOR2D0 C2807 ( .A1(a[269]), .A2(b[269]), .Z(p[269]) );
  XOR2D0 C2806 ( .A1(a[270]), .A2(b[270]), .Z(p[270]) );
  XOR2D0 C2805 ( .A1(a[271]), .A2(b[271]), .Z(p[271]) );
  XOR2D0 C2804 ( .A1(a[272]), .A2(b[272]), .Z(p[272]) );
  XOR2D0 C2803 ( .A1(a[273]), .A2(b[273]), .Z(p[273]) );
  XOR2D0 C2802 ( .A1(a[274]), .A2(b[274]), .Z(p[274]) );
  XOR2D0 C2801 ( .A1(a[275]), .A2(b[275]), .Z(p[275]) );
  XOR2D0 C2800 ( .A1(a[276]), .A2(b[276]), .Z(p[276]) );
  XOR2D0 C2799 ( .A1(a[277]), .A2(b[277]), .Z(p[277]) );
  XOR2D0 C2798 ( .A1(a[278]), .A2(b[278]), .Z(p[278]) );
  XOR2D0 C2797 ( .A1(a[279]), .A2(b[279]), .Z(p[279]) );
  XOR2D0 C2796 ( .A1(a[280]), .A2(b[280]), .Z(p[280]) );
  XOR2D0 C2795 ( .A1(a[281]), .A2(b[281]), .Z(p[281]) );
  XOR2D0 C2794 ( .A1(a[282]), .A2(b[282]), .Z(p[282]) );
  XOR2D0 C2793 ( .A1(a[283]), .A2(b[283]), .Z(p[283]) );
  XOR2D0 C2792 ( .A1(a[284]), .A2(b[284]), .Z(p[284]) );
  XOR2D0 C2791 ( .A1(a[285]), .A2(b[285]), .Z(p[285]) );
  XOR2D0 C2790 ( .A1(a[286]), .A2(b[286]), .Z(p[286]) );
  XOR2D0 C2789 ( .A1(a[287]), .A2(b[287]), .Z(p[287]) );
  XOR2D0 C2788 ( .A1(a[288]), .A2(b[288]), .Z(p[288]) );
  XOR2D0 C2787 ( .A1(a[289]), .A2(b[289]), .Z(p[289]) );
  XOR2D0 C2786 ( .A1(a[290]), .A2(b[290]), .Z(p[290]) );
  XOR2D0 C2785 ( .A1(a[291]), .A2(b[291]), .Z(p[291]) );
  XOR2D0 C2784 ( .A1(a[292]), .A2(b[292]), .Z(p[292]) );
  XOR2D0 C2783 ( .A1(a[293]), .A2(b[293]), .Z(p[293]) );
  XOR2D0 C2782 ( .A1(a[294]), .A2(b[294]), .Z(p[294]) );
  XOR2D0 C2781 ( .A1(a[295]), .A2(b[295]), .Z(p[295]) );
  XOR2D0 C2780 ( .A1(a[296]), .A2(b[296]), .Z(p[296]) );
  XOR2D0 C2779 ( .A1(a[297]), .A2(b[297]), .Z(p[297]) );
  XOR2D0 C2778 ( .A1(a[298]), .A2(b[298]), .Z(p[298]) );
  XOR2D0 C2777 ( .A1(a[299]), .A2(b[299]), .Z(p[299]) );
  XOR2D0 C2776 ( .A1(a[300]), .A2(b[300]), .Z(p[300]) );
  XOR2D0 C2775 ( .A1(a[301]), .A2(b[301]), .Z(p[301]) );
  XOR2D0 C2774 ( .A1(a[302]), .A2(b[302]), .Z(p[302]) );
  XOR2D0 C2773 ( .A1(a[303]), .A2(b[303]), .Z(p[303]) );
  XOR2D0 C2772 ( .A1(a[304]), .A2(b[304]), .Z(p[304]) );
  XOR2D0 C2771 ( .A1(a[305]), .A2(b[305]), .Z(p[305]) );
  XOR2D0 C2770 ( .A1(a[306]), .A2(b[306]), .Z(p[306]) );
  XOR2D0 C2769 ( .A1(a[307]), .A2(b[307]), .Z(p[307]) );
  XOR2D0 C2768 ( .A1(a[308]), .A2(b[308]), .Z(p[308]) );
  XOR2D0 C2767 ( .A1(a[309]), .A2(b[309]), .Z(p[309]) );
  XOR2D0 C2766 ( .A1(a[310]), .A2(b[310]), .Z(p[310]) );
  XOR2D0 C2765 ( .A1(a[311]), .A2(b[311]), .Z(p[311]) );
  XOR2D0 C2764 ( .A1(a[312]), .A2(b[312]), .Z(p[312]) );
  XOR2D0 C2763 ( .A1(a[313]), .A2(b[313]), .Z(p[313]) );
  XOR2D0 C2762 ( .A1(a[314]), .A2(b[314]), .Z(p[314]) );
  XOR2D0 C2761 ( .A1(a[315]), .A2(b[315]), .Z(p[315]) );
  XOR2D0 C2760 ( .A1(a[316]), .A2(b[316]), .Z(p[316]) );
  XOR2D0 C2759 ( .A1(a[317]), .A2(b[317]), .Z(p[317]) );
  XOR2D0 C2758 ( .A1(a[318]), .A2(b[318]), .Z(p[318]) );
  XOR2D0 C2757 ( .A1(a[319]), .A2(b[319]), .Z(p[319]) );
  XOR2D0 C2756 ( .A1(a[320]), .A2(b[320]), .Z(p[320]) );
  XOR2D0 C2755 ( .A1(a[321]), .A2(b[321]), .Z(p[321]) );
  XOR2D0 C2754 ( .A1(a[322]), .A2(b[322]), .Z(p[322]) );
  XOR2D0 C2753 ( .A1(a[323]), .A2(b[323]), .Z(p[323]) );
  XOR2D0 C2752 ( .A1(a[324]), .A2(b[324]), .Z(p[324]) );
  XOR2D0 C2751 ( .A1(a[325]), .A2(b[325]), .Z(p[325]) );
  XOR2D0 C2750 ( .A1(a[326]), .A2(b[326]), .Z(p[326]) );
  XOR2D0 C2749 ( .A1(a[327]), .A2(b[327]), .Z(p[327]) );
  XOR2D0 C2748 ( .A1(a[328]), .A2(b[328]), .Z(p[328]) );
  XOR2D0 C2747 ( .A1(a[329]), .A2(b[329]), .Z(p[329]) );
  XOR2D0 C2746 ( .A1(a[330]), .A2(b[330]), .Z(p[330]) );
  XOR2D0 C2745 ( .A1(a[331]), .A2(b[331]), .Z(p[331]) );
  XOR2D0 C2744 ( .A1(a[332]), .A2(b[332]), .Z(p[332]) );
  XOR2D0 C2743 ( .A1(a[333]), .A2(b[333]), .Z(p[333]) );
  XOR2D0 C2742 ( .A1(a[334]), .A2(b[334]), .Z(p[334]) );
  XOR2D0 C2741 ( .A1(a[335]), .A2(b[335]), .Z(p[335]) );
  XOR2D0 C2740 ( .A1(a[336]), .A2(b[336]), .Z(p[336]) );
  XOR2D0 C2739 ( .A1(a[337]), .A2(b[337]), .Z(p[337]) );
  XOR2D0 C2738 ( .A1(a[338]), .A2(b[338]), .Z(p[338]) );
  XOR2D0 C2737 ( .A1(a[339]), .A2(b[339]), .Z(p[339]) );
  XOR2D0 C2736 ( .A1(a[340]), .A2(b[340]), .Z(p[340]) );
  XOR2D0 C2735 ( .A1(a[341]), .A2(b[341]), .Z(p[341]) );
  XOR2D0 C2734 ( .A1(a[342]), .A2(b[342]), .Z(p[342]) );
  XOR2D0 C2733 ( .A1(a[343]), .A2(b[343]), .Z(p[343]) );
  XOR2D0 C2732 ( .A1(a[344]), .A2(b[344]), .Z(p[344]) );
  XOR2D0 C2731 ( .A1(a[345]), .A2(b[345]), .Z(p[345]) );
  XOR2D0 C2730 ( .A1(a[346]), .A2(b[346]), .Z(p[346]) );
  XOR2D0 C2729 ( .A1(a[347]), .A2(b[347]), .Z(p[347]) );
  XOR2D0 C2728 ( .A1(a[348]), .A2(b[348]), .Z(p[348]) );
  XOR2D0 C2727 ( .A1(a[349]), .A2(b[349]), .Z(p[349]) );
  XOR2D0 C2726 ( .A1(a[350]), .A2(b[350]), .Z(p[350]) );
  XOR2D0 C2725 ( .A1(a[351]), .A2(b[351]), .Z(p[351]) );
  XOR2D0 C2724 ( .A1(a[352]), .A2(b[352]), .Z(p[352]) );
  XOR2D0 C2723 ( .A1(a[353]), .A2(b[353]), .Z(p[353]) );
  XOR2D0 C2722 ( .A1(a[354]), .A2(b[354]), .Z(p[354]) );
  XOR2D0 C2721 ( .A1(a[355]), .A2(b[355]), .Z(p[355]) );
  XOR2D0 C2720 ( .A1(a[356]), .A2(b[356]), .Z(p[356]) );
  XOR2D0 C2719 ( .A1(a[357]), .A2(b[357]), .Z(p[357]) );
  XOR2D0 C2718 ( .A1(a[358]), .A2(b[358]), .Z(p[358]) );
  XOR2D0 C2717 ( .A1(a[359]), .A2(b[359]), .Z(p[359]) );
  XOR2D0 C2716 ( .A1(a[360]), .A2(b[360]), .Z(p[360]) );
  XOR2D0 C2715 ( .A1(a[361]), .A2(b[361]), .Z(p[361]) );
  XOR2D0 C2714 ( .A1(a[362]), .A2(b[362]), .Z(p[362]) );
  XOR2D0 C2713 ( .A1(a[363]), .A2(b[363]), .Z(p[363]) );
  XOR2D0 C2712 ( .A1(a[364]), .A2(b[364]), .Z(p[364]) );
  XOR2D0 C2711 ( .A1(a[365]), .A2(b[365]), .Z(p[365]) );
  XOR2D0 C2710 ( .A1(a[366]), .A2(b[366]), .Z(p[366]) );
  XOR2D0 C2709 ( .A1(a[367]), .A2(b[367]), .Z(p[367]) );
  XOR2D0 C2708 ( .A1(a[368]), .A2(b[368]), .Z(p[368]) );
  XOR2D0 C2707 ( .A1(a[369]), .A2(b[369]), .Z(p[369]) );
  XOR2D0 C2706 ( .A1(a[370]), .A2(b[370]), .Z(p[370]) );
  XOR2D0 C2705 ( .A1(a[371]), .A2(b[371]), .Z(p[371]) );
  XOR2D0 C2704 ( .A1(a[372]), .A2(b[372]), .Z(p[372]) );
  XOR2D0 C2703 ( .A1(a[373]), .A2(b[373]), .Z(p[373]) );
  XOR2D0 C2702 ( .A1(a[374]), .A2(b[374]), .Z(p[374]) );
  XOR2D0 C2701 ( .A1(a[375]), .A2(b[375]), .Z(p[375]) );
  XOR2D0 C2700 ( .A1(a[376]), .A2(b[376]), .Z(p[376]) );
  XOR2D0 C2699 ( .A1(a[377]), .A2(b[377]), .Z(p[377]) );
  XOR2D0 C2698 ( .A1(a[378]), .A2(b[378]), .Z(p[378]) );
  XOR2D0 C2697 ( .A1(a[379]), .A2(b[379]), .Z(p[379]) );
  XOR2D0 C2696 ( .A1(a[380]), .A2(b[380]), .Z(p[380]) );
  XOR2D0 C2695 ( .A1(a[381]), .A2(b[381]), .Z(p[381]) );
  XOR2D0 C2694 ( .A1(a[382]), .A2(b[382]), .Z(p[382]) );
  XOR2D0 C2693 ( .A1(a[383]), .A2(b[383]), .Z(p[383]) );
  XOR2D0 C2692 ( .A1(a[384]), .A2(b[384]), .Z(p[384]) );
  XOR2D0 C2691 ( .A1(a[385]), .A2(b[385]), .Z(p[385]) );
  XOR2D0 C2690 ( .A1(a[386]), .A2(b[386]), .Z(p[386]) );
  XOR2D0 C2689 ( .A1(a[387]), .A2(b[387]), .Z(p[387]) );
  XOR2D0 C2688 ( .A1(a[388]), .A2(b[388]), .Z(p[388]) );
  XOR2D0 C2687 ( .A1(a[389]), .A2(b[389]), .Z(p[389]) );
  XOR2D0 C2686 ( .A1(a[390]), .A2(b[390]), .Z(p[390]) );
  XOR2D0 C2685 ( .A1(a[391]), .A2(b[391]), .Z(p[391]) );
  XOR2D0 C2684 ( .A1(a[392]), .A2(b[392]), .Z(p[392]) );
  XOR2D0 C2683 ( .A1(a[393]), .A2(b[393]), .Z(p[393]) );
  XOR2D0 C2682 ( .A1(a[394]), .A2(b[394]), .Z(p[394]) );
  XOR2D0 C2681 ( .A1(a[395]), .A2(b[395]), .Z(p[395]) );
  XOR2D0 C2680 ( .A1(a[396]), .A2(b[396]), .Z(p[396]) );
  XOR2D0 C2679 ( .A1(a[397]), .A2(b[397]), .Z(p[397]) );
  XOR2D0 C2678 ( .A1(a[398]), .A2(b[398]), .Z(p[398]) );
  XOR2D0 C2677 ( .A1(a[399]), .A2(b[399]), .Z(p[399]) );
  XOR2D0 C2676 ( .A1(a[400]), .A2(b[400]), .Z(p[400]) );
  XOR2D0 C2675 ( .A1(a[401]), .A2(b[401]), .Z(p[401]) );
  XOR2D0 C2674 ( .A1(a[402]), .A2(b[402]), .Z(p[402]) );
  XOR2D0 C2673 ( .A1(a[403]), .A2(b[403]), .Z(p[403]) );
  XOR2D0 C2672 ( .A1(a[404]), .A2(b[404]), .Z(p[404]) );
  XOR2D0 C2671 ( .A1(a[405]), .A2(b[405]), .Z(p[405]) );
  XOR2D0 C2670 ( .A1(a[406]), .A2(b[406]), .Z(p[406]) );
  XOR2D0 C2669 ( .A1(a[407]), .A2(b[407]), .Z(p[407]) );
  XOR2D0 C2668 ( .A1(a[408]), .A2(b[408]), .Z(p[408]) );
  XOR2D0 C2667 ( .A1(a[409]), .A2(b[409]), .Z(p[409]) );
  XOR2D0 C2666 ( .A1(a[410]), .A2(b[410]), .Z(p[410]) );
  XOR2D0 C2665 ( .A1(a[411]), .A2(b[411]), .Z(p[411]) );
  XOR2D0 C2664 ( .A1(a[412]), .A2(b[412]), .Z(p[412]) );
  XOR2D0 C2663 ( .A1(a[413]), .A2(b[413]), .Z(p[413]) );
  XOR2D0 C2662 ( .A1(a[414]), .A2(b[414]), .Z(p[414]) );
  XOR2D0 C2661 ( .A1(a[415]), .A2(b[415]), .Z(p[415]) );
  XOR2D0 C2660 ( .A1(a[416]), .A2(b[416]), .Z(p[416]) );
  XOR2D0 C2659 ( .A1(a[417]), .A2(b[417]), .Z(p[417]) );
  XOR2D0 C2658 ( .A1(a[418]), .A2(b[418]), .Z(p[418]) );
  XOR2D0 C2657 ( .A1(a[419]), .A2(b[419]), .Z(p[419]) );
  XOR2D0 C2656 ( .A1(a[420]), .A2(b[420]), .Z(p[420]) );
  XOR2D0 C2655 ( .A1(a[421]), .A2(b[421]), .Z(p[421]) );
  XOR2D0 C2654 ( .A1(a[422]), .A2(b[422]), .Z(p[422]) );
  XOR2D0 C2653 ( .A1(a[423]), .A2(b[423]), .Z(p[423]) );
  XOR2D0 C2652 ( .A1(a[424]), .A2(b[424]), .Z(p[424]) );
  XOR2D0 C2651 ( .A1(a[425]), .A2(b[425]), .Z(p[425]) );
  XOR2D0 C2650 ( .A1(a[426]), .A2(b[426]), .Z(p[426]) );
  XOR2D0 C2649 ( .A1(a[427]), .A2(b[427]), .Z(p[427]) );
  XOR2D0 C2648 ( .A1(a[428]), .A2(b[428]), .Z(p[428]) );
  XOR2D0 C2647 ( .A1(a[429]), .A2(b[429]), .Z(p[429]) );
  XOR2D0 C2646 ( .A1(a[430]), .A2(b[430]), .Z(p[430]) );
  XOR2D0 C2645 ( .A1(a[431]), .A2(b[431]), .Z(p[431]) );
  XOR2D0 C2644 ( .A1(a[432]), .A2(b[432]), .Z(p[432]) );
  XOR2D0 C2643 ( .A1(a[433]), .A2(b[433]), .Z(p[433]) );
  XOR2D0 C2642 ( .A1(a[434]), .A2(b[434]), .Z(p[434]) );
  XOR2D0 C2641 ( .A1(a[435]), .A2(b[435]), .Z(p[435]) );
  XOR2D0 C2640 ( .A1(a[436]), .A2(b[436]), .Z(p[436]) );
  XOR2D0 C2639 ( .A1(a[437]), .A2(b[437]), .Z(p[437]) );
  XOR2D0 C2638 ( .A1(a[438]), .A2(b[438]), .Z(p[438]) );
  XOR2D0 C2637 ( .A1(a[439]), .A2(b[439]), .Z(p[439]) );
  XOR2D0 C2636 ( .A1(a[440]), .A2(b[440]), .Z(p[440]) );
  XOR2D0 C2635 ( .A1(a[441]), .A2(b[441]), .Z(p[441]) );
  XOR2D0 C2634 ( .A1(a[442]), .A2(b[442]), .Z(p[442]) );
  XOR2D0 C2633 ( .A1(a[443]), .A2(b[443]), .Z(p[443]) );
  XOR2D0 C2632 ( .A1(a[444]), .A2(b[444]), .Z(p[444]) );
  XOR2D0 C2631 ( .A1(a[445]), .A2(b[445]), .Z(p[445]) );
  XOR2D0 C2630 ( .A1(a[446]), .A2(b[446]), .Z(p[446]) );
  XOR2D0 C2629 ( .A1(a[447]), .A2(b[447]), .Z(p[447]) );
  XOR2D0 C2628 ( .A1(a[448]), .A2(b[448]), .Z(p[448]) );
  XOR2D0 C2627 ( .A1(a[449]), .A2(b[449]), .Z(p[449]) );
  XOR2D0 C2626 ( .A1(a[450]), .A2(b[450]), .Z(p[450]) );
  XOR2D0 C2625 ( .A1(a[451]), .A2(b[451]), .Z(p[451]) );
  XOR2D0 C2624 ( .A1(a[452]), .A2(b[452]), .Z(p[452]) );
  XOR2D0 C2623 ( .A1(a[453]), .A2(b[453]), .Z(p[453]) );
  XOR2D0 C2622 ( .A1(a[454]), .A2(b[454]), .Z(p[454]) );
  XOR2D0 C2621 ( .A1(a[455]), .A2(b[455]), .Z(p[455]) );
  XOR2D0 C2620 ( .A1(a[456]), .A2(b[456]), .Z(p[456]) );
  XOR2D0 C2619 ( .A1(a[457]), .A2(b[457]), .Z(p[457]) );
  XOR2D0 C2618 ( .A1(a[458]), .A2(b[458]), .Z(p[458]) );
  XOR2D0 C2617 ( .A1(a[459]), .A2(b[459]), .Z(p[459]) );
  XOR2D0 C2616 ( .A1(a[460]), .A2(b[460]), .Z(p[460]) );
  XOR2D0 C2615 ( .A1(a[461]), .A2(b[461]), .Z(p[461]) );
  XOR2D0 C2614 ( .A1(a[462]), .A2(b[462]), .Z(p[462]) );
  XOR2D0 C2613 ( .A1(a[463]), .A2(b[463]), .Z(p[463]) );
  XOR2D0 C2612 ( .A1(a[464]), .A2(b[464]), .Z(p[464]) );
  XOR2D0 C2611 ( .A1(a[465]), .A2(b[465]), .Z(p[465]) );
  XOR2D0 C2610 ( .A1(a[466]), .A2(b[466]), .Z(p[466]) );
  XOR2D0 C2609 ( .A1(a[467]), .A2(b[467]), .Z(p[467]) );
  XOR2D0 C2608 ( .A1(a[468]), .A2(b[468]), .Z(p[468]) );
  XOR2D0 C2607 ( .A1(a[469]), .A2(b[469]), .Z(p[469]) );
  XOR2D0 C2606 ( .A1(a[470]), .A2(b[470]), .Z(p[470]) );
  XOR2D0 C2605 ( .A1(a[471]), .A2(b[471]), .Z(p[471]) );
  XOR2D0 C2604 ( .A1(a[472]), .A2(b[472]), .Z(p[472]) );
  XOR2D0 C2603 ( .A1(a[473]), .A2(b[473]), .Z(p[473]) );
  XOR2D0 C2602 ( .A1(a[474]), .A2(b[474]), .Z(p[474]) );
  XOR2D0 C2601 ( .A1(a[475]), .A2(b[475]), .Z(p[475]) );
  XOR2D0 C2600 ( .A1(a[476]), .A2(b[476]), .Z(p[476]) );
  XOR2D0 C2599 ( .A1(a[477]), .A2(b[477]), .Z(p[477]) );
  XOR2D0 C2598 ( .A1(a[478]), .A2(b[478]), .Z(p[478]) );
  XOR2D0 C2597 ( .A1(a[479]), .A2(b[479]), .Z(p[479]) );
  XOR2D0 C2596 ( .A1(a[480]), .A2(b[480]), .Z(p[480]) );
  XOR2D0 C2595 ( .A1(a[481]), .A2(b[481]), .Z(p[481]) );
  XOR2D0 C2594 ( .A1(a[482]), .A2(b[482]), .Z(p[482]) );
  XOR2D0 C2593 ( .A1(a[483]), .A2(b[483]), .Z(p[483]) );
  XOR2D0 C2592 ( .A1(a[484]), .A2(b[484]), .Z(p[484]) );
  XOR2D0 C2591 ( .A1(a[485]), .A2(b[485]), .Z(p[485]) );
  XOR2D0 C2590 ( .A1(a[486]), .A2(b[486]), .Z(p[486]) );
  XOR2D0 C2589 ( .A1(a[487]), .A2(b[487]), .Z(p[487]) );
  XOR2D0 C2588 ( .A1(a[488]), .A2(b[488]), .Z(p[488]) );
  XOR2D0 C2587 ( .A1(a[489]), .A2(b[489]), .Z(p[489]) );
  XOR2D0 C2586 ( .A1(a[490]), .A2(b[490]), .Z(p[490]) );
  XOR2D0 C2585 ( .A1(a[491]), .A2(b[491]), .Z(p[491]) );
  XOR2D0 C2584 ( .A1(a[492]), .A2(b[492]), .Z(p[492]) );
  XOR2D0 C2583 ( .A1(a[493]), .A2(b[493]), .Z(p[493]) );
  XOR2D0 C2582 ( .A1(a[494]), .A2(b[494]), .Z(p[494]) );
  XOR2D0 C2581 ( .A1(a[495]), .A2(b[495]), .Z(p[495]) );
  XOR2D0 C2580 ( .A1(a[496]), .A2(b[496]), .Z(p[496]) );
  XOR2D0 C2579 ( .A1(a[497]), .A2(b[497]), .Z(p[497]) );
  XOR2D0 C2578 ( .A1(a[498]), .A2(b[498]), .Z(p[498]) );
  XOR2D0 C2577 ( .A1(a[499]), .A2(b[499]), .Z(p[499]) );
  XOR2D0 C2576 ( .A1(a[500]), .A2(b[500]), .Z(p[500]) );
  XOR2D0 C2575 ( .A1(a[501]), .A2(b[501]), .Z(p[501]) );
  XOR2D0 C2574 ( .A1(a[502]), .A2(b[502]), .Z(p[502]) );
  XOR2D0 C2573 ( .A1(a[503]), .A2(b[503]), .Z(p[503]) );
  XOR2D0 C2572 ( .A1(a[504]), .A2(b[504]), .Z(p[504]) );
  XOR2D0 C2571 ( .A1(a[505]), .A2(b[505]), .Z(p[505]) );
  XOR2D0 C2570 ( .A1(a[506]), .A2(b[506]), .Z(p[506]) );
  XOR2D0 C2569 ( .A1(a[507]), .A2(b[507]), .Z(p[507]) );
  XOR2D0 C2568 ( .A1(a[508]), .A2(b[508]), .Z(p[508]) );
  XOR2D0 C2567 ( .A1(a[509]), .A2(b[509]), .Z(p[509]) );
  XOR2D0 C2566 ( .A1(a[510]), .A2(b[510]), .Z(p[510]) );
  XOR2D0 C2565 ( .A1(a[511]), .A2(b[511]), .Z(p[511]) );
  AN2D0 C2564 ( .A1(a[0]), .A2(b[0]), .Z(g[0]) );
  AN2D0 C2563 ( .A1(a[1]), .A2(b[1]), .Z(g[1]) );
  AN2D0 C2562 ( .A1(a[2]), .A2(b[2]), .Z(g[2]) );
  AN2D0 C2561 ( .A1(a[3]), .A2(b[3]), .Z(g[3]) );
  AN2D0 C2560 ( .A1(a[4]), .A2(b[4]), .Z(g[4]) );
  AN2D0 C2559 ( .A1(a[5]), .A2(b[5]), .Z(g[5]) );
  AN2D0 C2558 ( .A1(a[6]), .A2(b[6]), .Z(g[6]) );
  AN2D0 C2557 ( .A1(a[7]), .A2(b[7]), .Z(g[7]) );
  AN2D0 C2556 ( .A1(a[8]), .A2(b[8]), .Z(g[8]) );
  AN2D0 C2555 ( .A1(a[9]), .A2(b[9]), .Z(g[9]) );
  AN2D0 C2554 ( .A1(a[10]), .A2(b[10]), .Z(g[10]) );
  AN2D0 C2553 ( .A1(a[11]), .A2(b[11]), .Z(g[11]) );
  AN2D0 C2552 ( .A1(a[12]), .A2(b[12]), .Z(g[12]) );
  AN2D0 C2551 ( .A1(a[13]), .A2(b[13]), .Z(g[13]) );
  AN2D0 C2550 ( .A1(a[14]), .A2(b[14]), .Z(g[14]) );
  AN2D0 C2549 ( .A1(a[15]), .A2(b[15]), .Z(g[15]) );
  AN2D0 C2548 ( .A1(a[16]), .A2(b[16]), .Z(g[16]) );
  AN2D0 C2547 ( .A1(a[17]), .A2(b[17]), .Z(g[17]) );
  AN2D0 C2546 ( .A1(a[18]), .A2(b[18]), .Z(g[18]) );
  AN2D0 C2545 ( .A1(a[19]), .A2(b[19]), .Z(g[19]) );
  AN2D0 C2544 ( .A1(a[20]), .A2(b[20]), .Z(g[20]) );
  AN2D0 C2543 ( .A1(a[21]), .A2(b[21]), .Z(g[21]) );
  AN2D0 C2542 ( .A1(a[22]), .A2(b[22]), .Z(g[22]) );
  AN2D0 C2541 ( .A1(a[23]), .A2(b[23]), .Z(g[23]) );
  AN2D0 C2540 ( .A1(a[24]), .A2(b[24]), .Z(g[24]) );
  AN2D0 C2539 ( .A1(a[25]), .A2(b[25]), .Z(g[25]) );
  AN2D0 C2538 ( .A1(a[26]), .A2(b[26]), .Z(g[26]) );
  AN2D0 C2537 ( .A1(a[27]), .A2(b[27]), .Z(g[27]) );
  AN2D0 C2536 ( .A1(a[28]), .A2(b[28]), .Z(g[28]) );
  AN2D0 C2535 ( .A1(a[29]), .A2(b[29]), .Z(g[29]) );
  AN2D0 C2534 ( .A1(a[30]), .A2(b[30]), .Z(g[30]) );
  AN2D0 C2533 ( .A1(a[31]), .A2(b[31]), .Z(g[31]) );
  AN2D0 C2532 ( .A1(a[32]), .A2(b[32]), .Z(g[32]) );
  AN2D0 C2531 ( .A1(a[33]), .A2(b[33]), .Z(g[33]) );
  AN2D0 C2530 ( .A1(a[34]), .A2(b[34]), .Z(g[34]) );
  AN2D0 C2529 ( .A1(a[35]), .A2(b[35]), .Z(g[35]) );
  AN2D0 C2528 ( .A1(a[36]), .A2(b[36]), .Z(g[36]) );
  AN2D0 C2527 ( .A1(a[37]), .A2(b[37]), .Z(g[37]) );
  AN2D0 C2526 ( .A1(a[38]), .A2(b[38]), .Z(g[38]) );
  AN2D0 C2525 ( .A1(a[39]), .A2(b[39]), .Z(g[39]) );
  AN2D0 C2524 ( .A1(a[40]), .A2(b[40]), .Z(g[40]) );
  AN2D0 C2523 ( .A1(a[41]), .A2(b[41]), .Z(g[41]) );
  AN2D0 C2522 ( .A1(a[42]), .A2(b[42]), .Z(g[42]) );
  AN2D0 C2521 ( .A1(a[43]), .A2(b[43]), .Z(g[43]) );
  AN2D0 C2520 ( .A1(a[44]), .A2(b[44]), .Z(g[44]) );
  AN2D0 C2519 ( .A1(a[45]), .A2(b[45]), .Z(g[45]) );
  AN2D0 C2518 ( .A1(a[46]), .A2(b[46]), .Z(g[46]) );
  AN2D0 C2517 ( .A1(a[47]), .A2(b[47]), .Z(g[47]) );
  AN2D0 C2516 ( .A1(a[48]), .A2(b[48]), .Z(g[48]) );
  AN2D0 C2515 ( .A1(a[49]), .A2(b[49]), .Z(g[49]) );
  AN2D0 C2514 ( .A1(a[50]), .A2(b[50]), .Z(g[50]) );
  AN2D0 C2513 ( .A1(a[51]), .A2(b[51]), .Z(g[51]) );
  AN2D0 C2512 ( .A1(a[52]), .A2(b[52]), .Z(g[52]) );
  AN2D0 C2511 ( .A1(a[53]), .A2(b[53]), .Z(g[53]) );
  AN2D0 C2510 ( .A1(a[54]), .A2(b[54]), .Z(g[54]) );
  AN2D0 C2509 ( .A1(a[55]), .A2(b[55]), .Z(g[55]) );
  AN2D0 C2508 ( .A1(a[56]), .A2(b[56]), .Z(g[56]) );
  AN2D0 C2507 ( .A1(a[57]), .A2(b[57]), .Z(g[57]) );
  AN2D0 C2506 ( .A1(a[58]), .A2(b[58]), .Z(g[58]) );
  AN2D0 C2505 ( .A1(a[59]), .A2(b[59]), .Z(g[59]) );
  AN2D0 C2504 ( .A1(a[60]), .A2(b[60]), .Z(g[60]) );
  AN2D0 C2503 ( .A1(a[61]), .A2(b[61]), .Z(g[61]) );
  AN2D0 C2502 ( .A1(a[62]), .A2(b[62]), .Z(g[62]) );
  AN2D0 C2501 ( .A1(a[63]), .A2(b[63]), .Z(g[63]) );
  AN2D0 C2500 ( .A1(a[64]), .A2(b[64]), .Z(g[64]) );
  AN2D0 C2499 ( .A1(a[65]), .A2(b[65]), .Z(g[65]) );
  AN2D0 C2498 ( .A1(a[66]), .A2(b[66]), .Z(g[66]) );
  AN2D0 C2497 ( .A1(a[67]), .A2(b[67]), .Z(g[67]) );
  AN2D0 C2496 ( .A1(a[68]), .A2(b[68]), .Z(g[68]) );
  AN2D0 C2495 ( .A1(a[69]), .A2(b[69]), .Z(g[69]) );
  AN2D0 C2494 ( .A1(a[70]), .A2(b[70]), .Z(g[70]) );
  AN2D0 C2493 ( .A1(a[71]), .A2(b[71]), .Z(g[71]) );
  AN2D0 C2492 ( .A1(a[72]), .A2(b[72]), .Z(g[72]) );
  AN2D0 C2491 ( .A1(a[73]), .A2(b[73]), .Z(g[73]) );
  AN2D0 C2490 ( .A1(a[74]), .A2(b[74]), .Z(g[74]) );
  AN2D0 C2489 ( .A1(a[75]), .A2(b[75]), .Z(g[75]) );
  AN2D0 C2488 ( .A1(a[76]), .A2(b[76]), .Z(g[76]) );
  AN2D0 C2487 ( .A1(a[77]), .A2(b[77]), .Z(g[77]) );
  AN2D0 C2486 ( .A1(a[78]), .A2(b[78]), .Z(g[78]) );
  AN2D0 C2485 ( .A1(a[79]), .A2(b[79]), .Z(g[79]) );
  AN2D0 C2484 ( .A1(a[80]), .A2(b[80]), .Z(g[80]) );
  AN2D0 C2483 ( .A1(a[81]), .A2(b[81]), .Z(g[81]) );
  AN2D0 C2482 ( .A1(a[82]), .A2(b[82]), .Z(g[82]) );
  AN2D0 C2481 ( .A1(a[83]), .A2(b[83]), .Z(g[83]) );
  AN2D0 C2480 ( .A1(a[84]), .A2(b[84]), .Z(g[84]) );
  AN2D0 C2479 ( .A1(a[85]), .A2(b[85]), .Z(g[85]) );
  AN2D0 C2478 ( .A1(a[86]), .A2(b[86]), .Z(g[86]) );
  AN2D0 C2477 ( .A1(a[87]), .A2(b[87]), .Z(g[87]) );
  AN2D0 C2476 ( .A1(a[88]), .A2(b[88]), .Z(g[88]) );
  AN2D0 C2475 ( .A1(a[89]), .A2(b[89]), .Z(g[89]) );
  AN2D0 C2474 ( .A1(a[90]), .A2(b[90]), .Z(g[90]) );
  AN2D0 C2473 ( .A1(a[91]), .A2(b[91]), .Z(g[91]) );
  AN2D0 C2472 ( .A1(a[92]), .A2(b[92]), .Z(g[92]) );
  AN2D0 C2471 ( .A1(a[93]), .A2(b[93]), .Z(g[93]) );
  AN2D0 C2470 ( .A1(a[94]), .A2(b[94]), .Z(g[94]) );
  AN2D0 C2469 ( .A1(a[95]), .A2(b[95]), .Z(g[95]) );
  AN2D0 C2468 ( .A1(a[96]), .A2(b[96]), .Z(g[96]) );
  AN2D0 C2467 ( .A1(a[97]), .A2(b[97]), .Z(g[97]) );
  AN2D0 C2466 ( .A1(a[98]), .A2(b[98]), .Z(g[98]) );
  AN2D0 C2465 ( .A1(a[99]), .A2(b[99]), .Z(g[99]) );
  AN2D0 C2464 ( .A1(a[100]), .A2(b[100]), .Z(g[100]) );
  AN2D0 C2463 ( .A1(a[101]), .A2(b[101]), .Z(g[101]) );
  AN2D0 C2462 ( .A1(a[102]), .A2(b[102]), .Z(g[102]) );
  AN2D0 C2461 ( .A1(a[103]), .A2(b[103]), .Z(g[103]) );
  AN2D0 C2460 ( .A1(a[104]), .A2(b[104]), .Z(g[104]) );
  AN2D0 C2459 ( .A1(a[105]), .A2(b[105]), .Z(g[105]) );
  AN2D0 C2458 ( .A1(a[106]), .A2(b[106]), .Z(g[106]) );
  AN2D0 C2457 ( .A1(a[107]), .A2(b[107]), .Z(g[107]) );
  AN2D0 C2456 ( .A1(a[108]), .A2(b[108]), .Z(g[108]) );
  AN2D0 C2455 ( .A1(a[109]), .A2(b[109]), .Z(g[109]) );
  AN2D0 C2454 ( .A1(a[110]), .A2(b[110]), .Z(g[110]) );
  AN2D0 C2453 ( .A1(a[111]), .A2(b[111]), .Z(g[111]) );
  AN2D0 C2452 ( .A1(a[112]), .A2(b[112]), .Z(g[112]) );
  AN2D0 C2451 ( .A1(a[113]), .A2(b[113]), .Z(g[113]) );
  AN2D0 C2450 ( .A1(a[114]), .A2(b[114]), .Z(g[114]) );
  AN2D0 C2449 ( .A1(a[115]), .A2(b[115]), .Z(g[115]) );
  AN2D0 C2448 ( .A1(a[116]), .A2(b[116]), .Z(g[116]) );
  AN2D0 C2447 ( .A1(a[117]), .A2(b[117]), .Z(g[117]) );
  AN2D0 C2446 ( .A1(a[118]), .A2(b[118]), .Z(g[118]) );
  AN2D0 C2445 ( .A1(a[119]), .A2(b[119]), .Z(g[119]) );
  AN2D0 C2444 ( .A1(a[120]), .A2(b[120]), .Z(g[120]) );
  AN2D0 C2443 ( .A1(a[121]), .A2(b[121]), .Z(g[121]) );
  AN2D0 C2442 ( .A1(a[122]), .A2(b[122]), .Z(g[122]) );
  AN2D0 C2441 ( .A1(a[123]), .A2(b[123]), .Z(g[123]) );
  AN2D0 C2440 ( .A1(a[124]), .A2(b[124]), .Z(g[124]) );
  AN2D0 C2439 ( .A1(a[125]), .A2(b[125]), .Z(g[125]) );
  AN2D0 C2438 ( .A1(a[126]), .A2(b[126]), .Z(g[126]) );
  AN2D0 C2437 ( .A1(a[127]), .A2(b[127]), .Z(g[127]) );
  AN2D0 C2436 ( .A1(a[128]), .A2(b[128]), .Z(g[128]) );
  AN2D0 C2435 ( .A1(a[129]), .A2(b[129]), .Z(g[129]) );
  AN2D0 C2434 ( .A1(a[130]), .A2(b[130]), .Z(g[130]) );
  AN2D0 C2433 ( .A1(a[131]), .A2(b[131]), .Z(g[131]) );
  AN2D0 C2432 ( .A1(a[132]), .A2(b[132]), .Z(g[132]) );
  AN2D0 C2431 ( .A1(a[133]), .A2(b[133]), .Z(g[133]) );
  AN2D0 C2430 ( .A1(a[134]), .A2(b[134]), .Z(g[134]) );
  AN2D0 C2429 ( .A1(a[135]), .A2(b[135]), .Z(g[135]) );
  AN2D0 C2428 ( .A1(a[136]), .A2(b[136]), .Z(g[136]) );
  AN2D0 C2427 ( .A1(a[137]), .A2(b[137]), .Z(g[137]) );
  AN2D0 C2426 ( .A1(a[138]), .A2(b[138]), .Z(g[138]) );
  AN2D0 C2425 ( .A1(a[139]), .A2(b[139]), .Z(g[139]) );
  AN2D0 C2424 ( .A1(a[140]), .A2(b[140]), .Z(g[140]) );
  AN2D0 C2423 ( .A1(a[141]), .A2(b[141]), .Z(g[141]) );
  AN2D0 C2422 ( .A1(a[142]), .A2(b[142]), .Z(g[142]) );
  AN2D0 C2421 ( .A1(a[143]), .A2(b[143]), .Z(g[143]) );
  AN2D0 C2420 ( .A1(a[144]), .A2(b[144]), .Z(g[144]) );
  AN2D0 C2419 ( .A1(a[145]), .A2(b[145]), .Z(g[145]) );
  AN2D0 C2418 ( .A1(a[146]), .A2(b[146]), .Z(g[146]) );
  AN2D0 C2417 ( .A1(a[147]), .A2(b[147]), .Z(g[147]) );
  AN2D0 C2416 ( .A1(a[148]), .A2(b[148]), .Z(g[148]) );
  AN2D0 C2415 ( .A1(a[149]), .A2(b[149]), .Z(g[149]) );
  AN2D0 C2414 ( .A1(a[150]), .A2(b[150]), .Z(g[150]) );
  AN2D0 C2413 ( .A1(a[151]), .A2(b[151]), .Z(g[151]) );
  AN2D0 C2412 ( .A1(a[152]), .A2(b[152]), .Z(g[152]) );
  AN2D0 C2411 ( .A1(a[153]), .A2(b[153]), .Z(g[153]) );
  AN2D0 C2410 ( .A1(a[154]), .A2(b[154]), .Z(g[154]) );
  AN2D0 C2409 ( .A1(a[155]), .A2(b[155]), .Z(g[155]) );
  AN2D0 C2408 ( .A1(a[156]), .A2(b[156]), .Z(g[156]) );
  AN2D0 C2407 ( .A1(a[157]), .A2(b[157]), .Z(g[157]) );
  AN2D0 C2406 ( .A1(a[158]), .A2(b[158]), .Z(g[158]) );
  AN2D0 C2405 ( .A1(a[159]), .A2(b[159]), .Z(g[159]) );
  AN2D0 C2404 ( .A1(a[160]), .A2(b[160]), .Z(g[160]) );
  AN2D0 C2403 ( .A1(a[161]), .A2(b[161]), .Z(g[161]) );
  AN2D0 C2402 ( .A1(a[162]), .A2(b[162]), .Z(g[162]) );
  AN2D0 C2401 ( .A1(a[163]), .A2(b[163]), .Z(g[163]) );
  AN2D0 C2400 ( .A1(a[164]), .A2(b[164]), .Z(g[164]) );
  AN2D0 C2399 ( .A1(a[165]), .A2(b[165]), .Z(g[165]) );
  AN2D0 C2398 ( .A1(a[166]), .A2(b[166]), .Z(g[166]) );
  AN2D0 C2397 ( .A1(a[167]), .A2(b[167]), .Z(g[167]) );
  AN2D0 C2396 ( .A1(a[168]), .A2(b[168]), .Z(g[168]) );
  AN2D0 C2395 ( .A1(a[169]), .A2(b[169]), .Z(g[169]) );
  AN2D0 C2394 ( .A1(a[170]), .A2(b[170]), .Z(g[170]) );
  AN2D0 C2393 ( .A1(a[171]), .A2(b[171]), .Z(g[171]) );
  AN2D0 C2392 ( .A1(a[172]), .A2(b[172]), .Z(g[172]) );
  AN2D0 C2391 ( .A1(a[173]), .A2(b[173]), .Z(g[173]) );
  AN2D0 C2390 ( .A1(a[174]), .A2(b[174]), .Z(g[174]) );
  AN2D0 C2389 ( .A1(a[175]), .A2(b[175]), .Z(g[175]) );
  AN2D0 C2388 ( .A1(a[176]), .A2(b[176]), .Z(g[176]) );
  AN2D0 C2387 ( .A1(a[177]), .A2(b[177]), .Z(g[177]) );
  AN2D0 C2386 ( .A1(a[178]), .A2(b[178]), .Z(g[178]) );
  AN2D0 C2385 ( .A1(a[179]), .A2(b[179]), .Z(g[179]) );
  AN2D0 C2384 ( .A1(a[180]), .A2(b[180]), .Z(g[180]) );
  AN2D0 C2383 ( .A1(a[181]), .A2(b[181]), .Z(g[181]) );
  AN2D0 C2382 ( .A1(a[182]), .A2(b[182]), .Z(g[182]) );
  AN2D0 C2381 ( .A1(a[183]), .A2(b[183]), .Z(g[183]) );
  AN2D0 C2380 ( .A1(a[184]), .A2(b[184]), .Z(g[184]) );
  AN2D0 C2379 ( .A1(a[185]), .A2(b[185]), .Z(g[185]) );
  AN2D0 C2378 ( .A1(a[186]), .A2(b[186]), .Z(g[186]) );
  AN2D0 C2377 ( .A1(a[187]), .A2(b[187]), .Z(g[187]) );
  AN2D0 C2376 ( .A1(a[188]), .A2(b[188]), .Z(g[188]) );
  AN2D0 C2375 ( .A1(a[189]), .A2(b[189]), .Z(g[189]) );
  AN2D0 C2374 ( .A1(a[190]), .A2(b[190]), .Z(g[190]) );
  AN2D0 C2373 ( .A1(a[191]), .A2(b[191]), .Z(g[191]) );
  AN2D0 C2372 ( .A1(a[192]), .A2(b[192]), .Z(g[192]) );
  AN2D0 C2371 ( .A1(a[193]), .A2(b[193]), .Z(g[193]) );
  AN2D0 C2370 ( .A1(a[194]), .A2(b[194]), .Z(g[194]) );
  AN2D0 C2369 ( .A1(a[195]), .A2(b[195]), .Z(g[195]) );
  AN2D0 C2368 ( .A1(a[196]), .A2(b[196]), .Z(g[196]) );
  AN2D0 C2367 ( .A1(a[197]), .A2(b[197]), .Z(g[197]) );
  AN2D0 C2366 ( .A1(a[198]), .A2(b[198]), .Z(g[198]) );
  AN2D0 C2365 ( .A1(a[199]), .A2(b[199]), .Z(g[199]) );
  AN2D0 C2364 ( .A1(a[200]), .A2(b[200]), .Z(g[200]) );
  AN2D0 C2363 ( .A1(a[201]), .A2(b[201]), .Z(g[201]) );
  AN2D0 C2362 ( .A1(a[202]), .A2(b[202]), .Z(g[202]) );
  AN2D0 C2361 ( .A1(a[203]), .A2(b[203]), .Z(g[203]) );
  AN2D0 C2360 ( .A1(a[204]), .A2(b[204]), .Z(g[204]) );
  AN2D0 C2359 ( .A1(a[205]), .A2(b[205]), .Z(g[205]) );
  AN2D0 C2358 ( .A1(a[206]), .A2(b[206]), .Z(g[206]) );
  AN2D0 C2357 ( .A1(a[207]), .A2(b[207]), .Z(g[207]) );
  AN2D0 C2356 ( .A1(a[208]), .A2(b[208]), .Z(g[208]) );
  AN2D0 C2355 ( .A1(a[209]), .A2(b[209]), .Z(g[209]) );
  AN2D0 C2354 ( .A1(a[210]), .A2(b[210]), .Z(g[210]) );
  AN2D0 C2353 ( .A1(a[211]), .A2(b[211]), .Z(g[211]) );
  AN2D0 C2352 ( .A1(a[212]), .A2(b[212]), .Z(g[212]) );
  AN2D0 C2351 ( .A1(a[213]), .A2(b[213]), .Z(g[213]) );
  AN2D0 C2350 ( .A1(a[214]), .A2(b[214]), .Z(g[214]) );
  AN2D0 C2349 ( .A1(a[215]), .A2(b[215]), .Z(g[215]) );
  AN2D0 C2348 ( .A1(a[216]), .A2(b[216]), .Z(g[216]) );
  AN2D0 C2347 ( .A1(a[217]), .A2(b[217]), .Z(g[217]) );
  AN2D0 C2346 ( .A1(a[218]), .A2(b[218]), .Z(g[218]) );
  AN2D0 C2345 ( .A1(a[219]), .A2(b[219]), .Z(g[219]) );
  AN2D0 C2344 ( .A1(a[220]), .A2(b[220]), .Z(g[220]) );
  AN2D0 C2343 ( .A1(a[221]), .A2(b[221]), .Z(g[221]) );
  AN2D0 C2342 ( .A1(a[222]), .A2(b[222]), .Z(g[222]) );
  AN2D0 C2341 ( .A1(a[223]), .A2(b[223]), .Z(g[223]) );
  AN2D0 C2340 ( .A1(a[224]), .A2(b[224]), .Z(g[224]) );
  AN2D0 C2339 ( .A1(a[225]), .A2(b[225]), .Z(g[225]) );
  AN2D0 C2338 ( .A1(a[226]), .A2(b[226]), .Z(g[226]) );
  AN2D0 C2337 ( .A1(a[227]), .A2(b[227]), .Z(g[227]) );
  AN2D0 C2336 ( .A1(a[228]), .A2(b[228]), .Z(g[228]) );
  AN2D0 C2335 ( .A1(a[229]), .A2(b[229]), .Z(g[229]) );
  AN2D0 C2334 ( .A1(a[230]), .A2(b[230]), .Z(g[230]) );
  AN2D0 C2333 ( .A1(a[231]), .A2(b[231]), .Z(g[231]) );
  AN2D0 C2332 ( .A1(a[232]), .A2(b[232]), .Z(g[232]) );
  AN2D0 C2331 ( .A1(a[233]), .A2(b[233]), .Z(g[233]) );
  AN2D0 C2330 ( .A1(a[234]), .A2(b[234]), .Z(g[234]) );
  AN2D0 C2329 ( .A1(a[235]), .A2(b[235]), .Z(g[235]) );
  AN2D0 C2328 ( .A1(a[236]), .A2(b[236]), .Z(g[236]) );
  AN2D0 C2327 ( .A1(a[237]), .A2(b[237]), .Z(g[237]) );
  AN2D0 C2326 ( .A1(a[238]), .A2(b[238]), .Z(g[238]) );
  AN2D0 C2325 ( .A1(a[239]), .A2(b[239]), .Z(g[239]) );
  AN2D0 C2324 ( .A1(a[240]), .A2(b[240]), .Z(g[240]) );
  AN2D0 C2323 ( .A1(a[241]), .A2(b[241]), .Z(g[241]) );
  AN2D0 C2322 ( .A1(a[242]), .A2(b[242]), .Z(g[242]) );
  AN2D0 C2321 ( .A1(a[243]), .A2(b[243]), .Z(g[243]) );
  AN2D0 C2320 ( .A1(a[244]), .A2(b[244]), .Z(g[244]) );
  AN2D0 C2319 ( .A1(a[245]), .A2(b[245]), .Z(g[245]) );
  AN2D0 C2318 ( .A1(a[246]), .A2(b[246]), .Z(g[246]) );
  AN2D0 C2317 ( .A1(a[247]), .A2(b[247]), .Z(g[247]) );
  AN2D0 C2316 ( .A1(a[248]), .A2(b[248]), .Z(g[248]) );
  AN2D0 C2315 ( .A1(a[249]), .A2(b[249]), .Z(g[249]) );
  AN2D0 C2314 ( .A1(a[250]), .A2(b[250]), .Z(g[250]) );
  AN2D0 C2313 ( .A1(a[251]), .A2(b[251]), .Z(g[251]) );
  AN2D0 C2312 ( .A1(a[252]), .A2(b[252]), .Z(g[252]) );
  AN2D0 C2311 ( .A1(a[253]), .A2(b[253]), .Z(g[253]) );
  AN2D0 C2310 ( .A1(a[254]), .A2(b[254]), .Z(g[254]) );
  AN2D0 C2309 ( .A1(a[255]), .A2(b[255]), .Z(g[255]) );
  AN2D0 C2308 ( .A1(a[256]), .A2(b[256]), .Z(g[256]) );
  AN2D0 C2307 ( .A1(a[257]), .A2(b[257]), .Z(g[257]) );
  AN2D0 C2306 ( .A1(a[258]), .A2(b[258]), .Z(g[258]) );
  AN2D0 C2305 ( .A1(a[259]), .A2(b[259]), .Z(g[259]) );
  AN2D0 C2304 ( .A1(a[260]), .A2(b[260]), .Z(g[260]) );
  AN2D0 C2303 ( .A1(a[261]), .A2(b[261]), .Z(g[261]) );
  AN2D0 C2302 ( .A1(a[262]), .A2(b[262]), .Z(g[262]) );
  AN2D0 C2301 ( .A1(a[263]), .A2(b[263]), .Z(g[263]) );
  AN2D0 C2300 ( .A1(a[264]), .A2(b[264]), .Z(g[264]) );
  AN2D0 C2299 ( .A1(a[265]), .A2(b[265]), .Z(g[265]) );
  AN2D0 C2298 ( .A1(a[266]), .A2(b[266]), .Z(g[266]) );
  AN2D0 C2297 ( .A1(a[267]), .A2(b[267]), .Z(g[267]) );
  AN2D0 C2296 ( .A1(a[268]), .A2(b[268]), .Z(g[268]) );
  AN2D0 C2295 ( .A1(a[269]), .A2(b[269]), .Z(g[269]) );
  AN2D0 C2294 ( .A1(a[270]), .A2(b[270]), .Z(g[270]) );
  AN2D0 C2293 ( .A1(a[271]), .A2(b[271]), .Z(g[271]) );
  AN2D0 C2292 ( .A1(a[272]), .A2(b[272]), .Z(g[272]) );
  AN2D0 C2291 ( .A1(a[273]), .A2(b[273]), .Z(g[273]) );
  AN2D0 C2290 ( .A1(a[274]), .A2(b[274]), .Z(g[274]) );
  AN2D0 C2289 ( .A1(a[275]), .A2(b[275]), .Z(g[275]) );
  AN2D0 C2288 ( .A1(a[276]), .A2(b[276]), .Z(g[276]) );
  AN2D0 C2287 ( .A1(a[277]), .A2(b[277]), .Z(g[277]) );
  AN2D0 C2286 ( .A1(a[278]), .A2(b[278]), .Z(g[278]) );
  AN2D0 C2285 ( .A1(a[279]), .A2(b[279]), .Z(g[279]) );
  AN2D0 C2284 ( .A1(a[280]), .A2(b[280]), .Z(g[280]) );
  AN2D0 C2283 ( .A1(a[281]), .A2(b[281]), .Z(g[281]) );
  AN2D0 C2282 ( .A1(a[282]), .A2(b[282]), .Z(g[282]) );
  AN2D0 C2281 ( .A1(a[283]), .A2(b[283]), .Z(g[283]) );
  AN2D0 C2280 ( .A1(a[284]), .A2(b[284]), .Z(g[284]) );
  AN2D0 C2279 ( .A1(a[285]), .A2(b[285]), .Z(g[285]) );
  AN2D0 C2278 ( .A1(a[286]), .A2(b[286]), .Z(g[286]) );
  AN2D0 C2277 ( .A1(a[287]), .A2(b[287]), .Z(g[287]) );
  AN2D0 C2276 ( .A1(a[288]), .A2(b[288]), .Z(g[288]) );
  AN2D0 C2275 ( .A1(a[289]), .A2(b[289]), .Z(g[289]) );
  AN2D0 C2274 ( .A1(a[290]), .A2(b[290]), .Z(g[290]) );
  AN2D0 C2273 ( .A1(a[291]), .A2(b[291]), .Z(g[291]) );
  AN2D0 C2272 ( .A1(a[292]), .A2(b[292]), .Z(g[292]) );
  AN2D0 C2271 ( .A1(a[293]), .A2(b[293]), .Z(g[293]) );
  AN2D0 C2270 ( .A1(a[294]), .A2(b[294]), .Z(g[294]) );
  AN2D0 C2269 ( .A1(a[295]), .A2(b[295]), .Z(g[295]) );
  AN2D0 C2268 ( .A1(a[296]), .A2(b[296]), .Z(g[296]) );
  AN2D0 C2267 ( .A1(a[297]), .A2(b[297]), .Z(g[297]) );
  AN2D0 C2266 ( .A1(a[298]), .A2(b[298]), .Z(g[298]) );
  AN2D0 C2265 ( .A1(a[299]), .A2(b[299]), .Z(g[299]) );
  AN2D0 C2264 ( .A1(a[300]), .A2(b[300]), .Z(g[300]) );
  AN2D0 C2263 ( .A1(a[301]), .A2(b[301]), .Z(g[301]) );
  AN2D0 C2262 ( .A1(a[302]), .A2(b[302]), .Z(g[302]) );
  AN2D0 C2261 ( .A1(a[303]), .A2(b[303]), .Z(g[303]) );
  AN2D0 C2260 ( .A1(a[304]), .A2(b[304]), .Z(g[304]) );
  AN2D0 C2259 ( .A1(a[305]), .A2(b[305]), .Z(g[305]) );
  AN2D0 C2258 ( .A1(a[306]), .A2(b[306]), .Z(g[306]) );
  AN2D0 C2257 ( .A1(a[307]), .A2(b[307]), .Z(g[307]) );
  AN2D0 C2256 ( .A1(a[308]), .A2(b[308]), .Z(g[308]) );
  AN2D0 C2255 ( .A1(a[309]), .A2(b[309]), .Z(g[309]) );
  AN2D0 C2254 ( .A1(a[310]), .A2(b[310]), .Z(g[310]) );
  AN2D0 C2253 ( .A1(a[311]), .A2(b[311]), .Z(g[311]) );
  AN2D0 C2252 ( .A1(a[312]), .A2(b[312]), .Z(g[312]) );
  AN2D0 C2251 ( .A1(a[313]), .A2(b[313]), .Z(g[313]) );
  AN2D0 C2250 ( .A1(a[314]), .A2(b[314]), .Z(g[314]) );
  AN2D0 C2249 ( .A1(a[315]), .A2(b[315]), .Z(g[315]) );
  AN2D0 C2248 ( .A1(a[316]), .A2(b[316]), .Z(g[316]) );
  AN2D0 C2247 ( .A1(a[317]), .A2(b[317]), .Z(g[317]) );
  AN2D0 C2246 ( .A1(a[318]), .A2(b[318]), .Z(g[318]) );
  AN2D0 C2245 ( .A1(a[319]), .A2(b[319]), .Z(g[319]) );
  AN2D0 C2244 ( .A1(a[320]), .A2(b[320]), .Z(g[320]) );
  AN2D0 C2243 ( .A1(a[321]), .A2(b[321]), .Z(g[321]) );
  AN2D0 C2242 ( .A1(a[322]), .A2(b[322]), .Z(g[322]) );
  AN2D0 C2241 ( .A1(a[323]), .A2(b[323]), .Z(g[323]) );
  AN2D0 C2240 ( .A1(a[324]), .A2(b[324]), .Z(g[324]) );
  AN2D0 C2239 ( .A1(a[325]), .A2(b[325]), .Z(g[325]) );
  AN2D0 C2238 ( .A1(a[326]), .A2(b[326]), .Z(g[326]) );
  AN2D0 C2237 ( .A1(a[327]), .A2(b[327]), .Z(g[327]) );
  AN2D0 C2236 ( .A1(a[328]), .A2(b[328]), .Z(g[328]) );
  AN2D0 C2235 ( .A1(a[329]), .A2(b[329]), .Z(g[329]) );
  AN2D0 C2234 ( .A1(a[330]), .A2(b[330]), .Z(g[330]) );
  AN2D0 C2233 ( .A1(a[331]), .A2(b[331]), .Z(g[331]) );
  AN2D0 C2232 ( .A1(a[332]), .A2(b[332]), .Z(g[332]) );
  AN2D0 C2231 ( .A1(a[333]), .A2(b[333]), .Z(g[333]) );
  AN2D0 C2230 ( .A1(a[334]), .A2(b[334]), .Z(g[334]) );
  AN2D0 C2229 ( .A1(a[335]), .A2(b[335]), .Z(g[335]) );
  AN2D0 C2228 ( .A1(a[336]), .A2(b[336]), .Z(g[336]) );
  AN2D0 C2227 ( .A1(a[337]), .A2(b[337]), .Z(g[337]) );
  AN2D0 C2226 ( .A1(a[338]), .A2(b[338]), .Z(g[338]) );
  AN2D0 C2225 ( .A1(a[339]), .A2(b[339]), .Z(g[339]) );
  AN2D0 C2224 ( .A1(a[340]), .A2(b[340]), .Z(g[340]) );
  AN2D0 C2223 ( .A1(a[341]), .A2(b[341]), .Z(g[341]) );
  AN2D0 C2222 ( .A1(a[342]), .A2(b[342]), .Z(g[342]) );
  AN2D0 C2221 ( .A1(a[343]), .A2(b[343]), .Z(g[343]) );
  AN2D0 C2220 ( .A1(a[344]), .A2(b[344]), .Z(g[344]) );
  AN2D0 C2219 ( .A1(a[345]), .A2(b[345]), .Z(g[345]) );
  AN2D0 C2218 ( .A1(a[346]), .A2(b[346]), .Z(g[346]) );
  AN2D0 C2217 ( .A1(a[347]), .A2(b[347]), .Z(g[347]) );
  AN2D0 C2216 ( .A1(a[348]), .A2(b[348]), .Z(g[348]) );
  AN2D0 C2215 ( .A1(a[349]), .A2(b[349]), .Z(g[349]) );
  AN2D0 C2214 ( .A1(a[350]), .A2(b[350]), .Z(g[350]) );
  AN2D0 C2213 ( .A1(a[351]), .A2(b[351]), .Z(g[351]) );
  AN2D0 C2212 ( .A1(a[352]), .A2(b[352]), .Z(g[352]) );
  AN2D0 C2211 ( .A1(a[353]), .A2(b[353]), .Z(g[353]) );
  AN2D0 C2210 ( .A1(a[354]), .A2(b[354]), .Z(g[354]) );
  AN2D0 C2209 ( .A1(a[355]), .A2(b[355]), .Z(g[355]) );
  AN2D0 C2208 ( .A1(a[356]), .A2(b[356]), .Z(g[356]) );
  AN2D0 C2207 ( .A1(a[357]), .A2(b[357]), .Z(g[357]) );
  AN2D0 C2206 ( .A1(a[358]), .A2(b[358]), .Z(g[358]) );
  AN2D0 C2205 ( .A1(a[359]), .A2(b[359]), .Z(g[359]) );
  AN2D0 C2204 ( .A1(a[360]), .A2(b[360]), .Z(g[360]) );
  AN2D0 C2203 ( .A1(a[361]), .A2(b[361]), .Z(g[361]) );
  AN2D0 C2202 ( .A1(a[362]), .A2(b[362]), .Z(g[362]) );
  AN2D0 C2201 ( .A1(a[363]), .A2(b[363]), .Z(g[363]) );
  AN2D0 C2200 ( .A1(a[364]), .A2(b[364]), .Z(g[364]) );
  AN2D0 C2199 ( .A1(a[365]), .A2(b[365]), .Z(g[365]) );
  AN2D0 C2198 ( .A1(a[366]), .A2(b[366]), .Z(g[366]) );
  AN2D0 C2197 ( .A1(a[367]), .A2(b[367]), .Z(g[367]) );
  AN2D0 C2196 ( .A1(a[368]), .A2(b[368]), .Z(g[368]) );
  AN2D0 C2195 ( .A1(a[369]), .A2(b[369]), .Z(g[369]) );
  AN2D0 C2194 ( .A1(a[370]), .A2(b[370]), .Z(g[370]) );
  AN2D0 C2193 ( .A1(a[371]), .A2(b[371]), .Z(g[371]) );
  AN2D0 C2192 ( .A1(a[372]), .A2(b[372]), .Z(g[372]) );
  AN2D0 C2191 ( .A1(a[373]), .A2(b[373]), .Z(g[373]) );
  AN2D0 C2190 ( .A1(a[374]), .A2(b[374]), .Z(g[374]) );
  AN2D0 C2189 ( .A1(a[375]), .A2(b[375]), .Z(g[375]) );
  AN2D0 C2188 ( .A1(a[376]), .A2(b[376]), .Z(g[376]) );
  AN2D0 C2187 ( .A1(a[377]), .A2(b[377]), .Z(g[377]) );
  AN2D0 C2186 ( .A1(a[378]), .A2(b[378]), .Z(g[378]) );
  AN2D0 C2185 ( .A1(a[379]), .A2(b[379]), .Z(g[379]) );
  AN2D0 C2184 ( .A1(a[380]), .A2(b[380]), .Z(g[380]) );
  AN2D0 C2183 ( .A1(a[381]), .A2(b[381]), .Z(g[381]) );
  AN2D0 C2182 ( .A1(a[382]), .A2(b[382]), .Z(g[382]) );
  AN2D0 C2181 ( .A1(a[383]), .A2(b[383]), .Z(g[383]) );
  AN2D0 C2180 ( .A1(a[384]), .A2(b[384]), .Z(g[384]) );
  AN2D0 C2179 ( .A1(a[385]), .A2(b[385]), .Z(g[385]) );
  AN2D0 C2178 ( .A1(a[386]), .A2(b[386]), .Z(g[386]) );
  AN2D0 C2177 ( .A1(a[387]), .A2(b[387]), .Z(g[387]) );
  AN2D0 C2176 ( .A1(a[388]), .A2(b[388]), .Z(g[388]) );
  AN2D0 C2175 ( .A1(a[389]), .A2(b[389]), .Z(g[389]) );
  AN2D0 C2174 ( .A1(a[390]), .A2(b[390]), .Z(g[390]) );
  AN2D0 C2173 ( .A1(a[391]), .A2(b[391]), .Z(g[391]) );
  AN2D0 C2172 ( .A1(a[392]), .A2(b[392]), .Z(g[392]) );
  AN2D0 C2171 ( .A1(a[393]), .A2(b[393]), .Z(g[393]) );
  AN2D0 C2170 ( .A1(a[394]), .A2(b[394]), .Z(g[394]) );
  AN2D0 C2169 ( .A1(a[395]), .A2(b[395]), .Z(g[395]) );
  AN2D0 C2168 ( .A1(a[396]), .A2(b[396]), .Z(g[396]) );
  AN2D0 C2167 ( .A1(a[397]), .A2(b[397]), .Z(g[397]) );
  AN2D0 C2166 ( .A1(a[398]), .A2(b[398]), .Z(g[398]) );
  AN2D0 C2165 ( .A1(a[399]), .A2(b[399]), .Z(g[399]) );
  AN2D0 C2164 ( .A1(a[400]), .A2(b[400]), .Z(g[400]) );
  AN2D0 C2163 ( .A1(a[401]), .A2(b[401]), .Z(g[401]) );
  AN2D0 C2162 ( .A1(a[402]), .A2(b[402]), .Z(g[402]) );
  AN2D0 C2161 ( .A1(a[403]), .A2(b[403]), .Z(g[403]) );
  AN2D0 C2160 ( .A1(a[404]), .A2(b[404]), .Z(g[404]) );
  AN2D0 C2159 ( .A1(a[405]), .A2(b[405]), .Z(g[405]) );
  AN2D0 C2158 ( .A1(a[406]), .A2(b[406]), .Z(g[406]) );
  AN2D0 C2157 ( .A1(a[407]), .A2(b[407]), .Z(g[407]) );
  AN2D0 C2156 ( .A1(a[408]), .A2(b[408]), .Z(g[408]) );
  AN2D0 C2155 ( .A1(a[409]), .A2(b[409]), .Z(g[409]) );
  AN2D0 C2154 ( .A1(a[410]), .A2(b[410]), .Z(g[410]) );
  AN2D0 C2153 ( .A1(a[411]), .A2(b[411]), .Z(g[411]) );
  AN2D0 C2152 ( .A1(a[412]), .A2(b[412]), .Z(g[412]) );
  AN2D0 C2151 ( .A1(a[413]), .A2(b[413]), .Z(g[413]) );
  AN2D0 C2150 ( .A1(a[414]), .A2(b[414]), .Z(g[414]) );
  AN2D0 C2149 ( .A1(a[415]), .A2(b[415]), .Z(g[415]) );
  AN2D0 C2148 ( .A1(a[416]), .A2(b[416]), .Z(g[416]) );
  AN2D0 C2147 ( .A1(a[417]), .A2(b[417]), .Z(g[417]) );
  AN2D0 C2146 ( .A1(a[418]), .A2(b[418]), .Z(g[418]) );
  AN2D0 C2145 ( .A1(a[419]), .A2(b[419]), .Z(g[419]) );
  AN2D0 C2144 ( .A1(a[420]), .A2(b[420]), .Z(g[420]) );
  AN2D0 C2143 ( .A1(a[421]), .A2(b[421]), .Z(g[421]) );
  AN2D0 C2142 ( .A1(a[422]), .A2(b[422]), .Z(g[422]) );
  AN2D0 C2141 ( .A1(a[423]), .A2(b[423]), .Z(g[423]) );
  AN2D0 C2140 ( .A1(a[424]), .A2(b[424]), .Z(g[424]) );
  AN2D0 C2139 ( .A1(a[425]), .A2(b[425]), .Z(g[425]) );
  AN2D0 C2138 ( .A1(a[426]), .A2(b[426]), .Z(g[426]) );
  AN2D0 C2137 ( .A1(a[427]), .A2(b[427]), .Z(g[427]) );
  AN2D0 C2136 ( .A1(a[428]), .A2(b[428]), .Z(g[428]) );
  AN2D0 C2135 ( .A1(a[429]), .A2(b[429]), .Z(g[429]) );
  AN2D0 C2134 ( .A1(a[430]), .A2(b[430]), .Z(g[430]) );
  AN2D0 C2133 ( .A1(a[431]), .A2(b[431]), .Z(g[431]) );
  AN2D0 C2132 ( .A1(a[432]), .A2(b[432]), .Z(g[432]) );
  AN2D0 C2131 ( .A1(a[433]), .A2(b[433]), .Z(g[433]) );
  AN2D0 C2130 ( .A1(a[434]), .A2(b[434]), .Z(g[434]) );
  AN2D0 C2129 ( .A1(a[435]), .A2(b[435]), .Z(g[435]) );
  AN2D0 C2128 ( .A1(a[436]), .A2(b[436]), .Z(g[436]) );
  AN2D0 C2127 ( .A1(a[437]), .A2(b[437]), .Z(g[437]) );
  AN2D0 C2126 ( .A1(a[438]), .A2(b[438]), .Z(g[438]) );
  AN2D0 C2125 ( .A1(a[439]), .A2(b[439]), .Z(g[439]) );
  AN2D0 C2124 ( .A1(a[440]), .A2(b[440]), .Z(g[440]) );
  AN2D0 C2123 ( .A1(a[441]), .A2(b[441]), .Z(g[441]) );
  AN2D0 C2122 ( .A1(a[442]), .A2(b[442]), .Z(g[442]) );
  AN2D0 C2121 ( .A1(a[443]), .A2(b[443]), .Z(g[443]) );
  AN2D0 C2120 ( .A1(a[444]), .A2(b[444]), .Z(g[444]) );
  AN2D0 C2119 ( .A1(a[445]), .A2(b[445]), .Z(g[445]) );
  AN2D0 C2118 ( .A1(a[446]), .A2(b[446]), .Z(g[446]) );
  AN2D0 C2117 ( .A1(a[447]), .A2(b[447]), .Z(g[447]) );
  AN2D0 C2116 ( .A1(a[448]), .A2(b[448]), .Z(g[448]) );
  AN2D0 C2115 ( .A1(a[449]), .A2(b[449]), .Z(g[449]) );
  AN2D0 C2114 ( .A1(a[450]), .A2(b[450]), .Z(g[450]) );
  AN2D0 C2113 ( .A1(a[451]), .A2(b[451]), .Z(g[451]) );
  AN2D0 C2112 ( .A1(a[452]), .A2(b[452]), .Z(g[452]) );
  AN2D0 C2111 ( .A1(a[453]), .A2(b[453]), .Z(g[453]) );
  AN2D0 C2110 ( .A1(a[454]), .A2(b[454]), .Z(g[454]) );
  AN2D0 C2109 ( .A1(a[455]), .A2(b[455]), .Z(g[455]) );
  AN2D0 C2108 ( .A1(a[456]), .A2(b[456]), .Z(g[456]) );
  AN2D0 C2107 ( .A1(a[457]), .A2(b[457]), .Z(g[457]) );
  AN2D0 C2106 ( .A1(a[458]), .A2(b[458]), .Z(g[458]) );
  AN2D0 C2105 ( .A1(a[459]), .A2(b[459]), .Z(g[459]) );
  AN2D0 C2104 ( .A1(a[460]), .A2(b[460]), .Z(g[460]) );
  AN2D0 C2103 ( .A1(a[461]), .A2(b[461]), .Z(g[461]) );
  AN2D0 C2102 ( .A1(a[462]), .A2(b[462]), .Z(g[462]) );
  AN2D0 C2101 ( .A1(a[463]), .A2(b[463]), .Z(g[463]) );
  AN2D0 C2100 ( .A1(a[464]), .A2(b[464]), .Z(g[464]) );
  AN2D0 C2099 ( .A1(a[465]), .A2(b[465]), .Z(g[465]) );
  AN2D0 C2098 ( .A1(a[466]), .A2(b[466]), .Z(g[466]) );
  AN2D0 C2097 ( .A1(a[467]), .A2(b[467]), .Z(g[467]) );
  AN2D0 C2096 ( .A1(a[468]), .A2(b[468]), .Z(g[468]) );
  AN2D0 C2095 ( .A1(a[469]), .A2(b[469]), .Z(g[469]) );
  AN2D0 C2094 ( .A1(a[470]), .A2(b[470]), .Z(g[470]) );
  AN2D0 C2093 ( .A1(a[471]), .A2(b[471]), .Z(g[471]) );
  AN2D0 C2092 ( .A1(a[472]), .A2(b[472]), .Z(g[472]) );
  AN2D0 C2091 ( .A1(a[473]), .A2(b[473]), .Z(g[473]) );
  AN2D0 C2090 ( .A1(a[474]), .A2(b[474]), .Z(g[474]) );
  AN2D0 C2089 ( .A1(a[475]), .A2(b[475]), .Z(g[475]) );
  AN2D0 C2088 ( .A1(a[476]), .A2(b[476]), .Z(g[476]) );
  AN2D0 C2087 ( .A1(a[477]), .A2(b[477]), .Z(g[477]) );
  AN2D0 C2086 ( .A1(a[478]), .A2(b[478]), .Z(g[478]) );
  AN2D0 C2085 ( .A1(a[479]), .A2(b[479]), .Z(g[479]) );
  AN2D0 C2084 ( .A1(a[480]), .A2(b[480]), .Z(g[480]) );
  AN2D0 C2083 ( .A1(a[481]), .A2(b[481]), .Z(g[481]) );
  AN2D0 C2082 ( .A1(a[482]), .A2(b[482]), .Z(g[482]) );
  AN2D0 C2081 ( .A1(a[483]), .A2(b[483]), .Z(g[483]) );
  AN2D0 C2080 ( .A1(a[484]), .A2(b[484]), .Z(g[484]) );
  AN2D0 C2079 ( .A1(a[485]), .A2(b[485]), .Z(g[485]) );
  AN2D0 C2078 ( .A1(a[486]), .A2(b[486]), .Z(g[486]) );
  AN2D0 C2077 ( .A1(a[487]), .A2(b[487]), .Z(g[487]) );
  AN2D0 C2076 ( .A1(a[488]), .A2(b[488]), .Z(g[488]) );
  AN2D0 C2075 ( .A1(a[489]), .A2(b[489]), .Z(g[489]) );
  AN2D0 C2074 ( .A1(a[490]), .A2(b[490]), .Z(g[490]) );
  AN2D0 C2073 ( .A1(a[491]), .A2(b[491]), .Z(g[491]) );
  AN2D0 C2072 ( .A1(a[492]), .A2(b[492]), .Z(g[492]) );
  AN2D0 C2071 ( .A1(a[493]), .A2(b[493]), .Z(g[493]) );
  AN2D0 C2070 ( .A1(a[494]), .A2(b[494]), .Z(g[494]) );
  AN2D0 C2069 ( .A1(a[495]), .A2(b[495]), .Z(g[495]) );
  AN2D0 C2068 ( .A1(a[496]), .A2(b[496]), .Z(g[496]) );
  AN2D0 C2067 ( .A1(a[497]), .A2(b[497]), .Z(g[497]) );
  AN2D0 C2066 ( .A1(a[498]), .A2(b[498]), .Z(g[498]) );
  AN2D0 C2065 ( .A1(a[499]), .A2(b[499]), .Z(g[499]) );
  AN2D0 C2064 ( .A1(a[500]), .A2(b[500]), .Z(g[500]) );
  AN2D0 C2063 ( .A1(a[501]), .A2(b[501]), .Z(g[501]) );
  AN2D0 C2062 ( .A1(a[502]), .A2(b[502]), .Z(g[502]) );
  AN2D0 C2061 ( .A1(a[503]), .A2(b[503]), .Z(g[503]) );
  AN2D0 C2060 ( .A1(a[504]), .A2(b[504]), .Z(g[504]) );
  AN2D0 C2059 ( .A1(a[505]), .A2(b[505]), .Z(g[505]) );
  AN2D0 C2058 ( .A1(a[506]), .A2(b[506]), .Z(g[506]) );
  AN2D0 C2057 ( .A1(a[507]), .A2(b[507]), .Z(g[507]) );
  AN2D0 C2056 ( .A1(a[508]), .A2(b[508]), .Z(g[508]) );
  AN2D0 C2055 ( .A1(a[509]), .A2(b[509]), .Z(g[509]) );
  AN2D0 C2054 ( .A1(a[510]), .A2(b[510]), .Z(g[510]) );
endmodule

