
module cla_adder ( a, b, s, cin, cout );
  input [1023:0] a;
  input [1023:0] b;
  output [1023:0] s;
  input cin;
  output cout;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242,
         N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253,
         N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264,
         N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374,
         N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N385,
         N386, N387, N388, N389, N390, N391, N392, N393, N394, N395, N396,
         N397, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440,
         N441, N442, N443, N444, N445, N446, N447, N448, N449, N450, N451,
         N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, N462,
         N463, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N496, N497, N498, N499, N500, N501, N502, N503, N504, N505, N506,
         N507, N508, N509, N510, N511, N512, N513, N514, N515, N516, N517,
         N518, N519, N520, N521, N522, N523, N524, N525, N526, N527, N528,
         N529, N530, N531, N532, N533, N534, N535, N536, N537, N538, N539,
         N540, N541, N542, N543, N544, N545, N546, N547, N548, N549, N550,
         N551, N552, N553, N554, N555, N556, N557, N558, N559, N560, N561,
         N562, N563, N564, N565, N566, N567, N568, N569, N570, N571, N572,
         N573, N574, N575, N576, N577, N578, N579, N580, N581, N582, N583,
         N584, N585, N586, N587, N588, N589, N590, N591, N592, N593, N594,
         N595, N596, N597, N598, N599, N600, N601, N602, N603, N604, N605,
         N606, N607, N608, N609, N610, N611, N612, N613, N614, N615, N616,
         N617, N618, N619, N620, N621, N622, N623, N624, N625, N626, N627,
         N628, N629, N630, N631, N632, N633, N634, N635, N636, N637, N638,
         N639, N640, N641, N642, N643, N644, N645, N646, N647, N648, N649,
         N650, N651, N652, N653, N654, N655, N656, N657, N658, N659, N660,
         N661, N662, N663, N664, N665, N666, N667, N668, N669, N670, N671,
         N672, N673, N674, N675, N676, N677, N678, N679, N680, N681, N682,
         N683, N684, N685, N686, N687, N688, N689, N690, N691, N692, N693,
         N694, N695, N696, N697, N698, N699, N700, N701, N702, N703, N704,
         N705, N706, N707, N708, N709, N710, N711, N712, N713, N714, N715,
         N716, N717, N718, N719, N720, N721, N722, N723, N724, N725, N726,
         N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737,
         N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748,
         N749, N750, N751, N752, N753, N754, N755, N756, N757, N758, N759,
         N760, N761, N762, N763, N764, N765, N766, N767, N768, N769, N770,
         N771, N772, N773, N774, N775, N776, N777, N778, N779, N780, N781,
         N782, N783, N784, N785, N786, N787, N788, N789, N790, N791, N792,
         N793, N794, N795, N796, N797, N798, N799, N800, N801, N802, N803,
         N804, N805, N806, N807, N808, N809, N810, N811, N812, N813, N814,
         N815, N816, N817, N818, N819, N820, N821, N822, N823, N824, N825,
         N826, N827, N828, N829, N830, N831, N832, N833, N834, N835, N836,
         N837, N838, N839, N840, N841, N842, N843, N844, N845, N846, N847,
         N848, N849, N850, N851, N852, N853, N854, N855, N856, N857, N858,
         N859, N860, N861, N862, N863, N864, N865, N866, N867, N868, N869,
         N870, N871, N872, N873, N874, N875, N876, N877, N878, N879, N880,
         N881, N882, N883, N884, N885, N886, N887, N888, N889, N890, N891,
         N892, N893, N894, N895, N896, N897, N898, N899, N900, N901, N902,
         N903, N904, N905, N906, N907, N908, N909, N910, N911, N912, N913,
         N914, N915, N916, N917, N918, N919, N920, N921, N922, N923, N924,
         N925, N926, N927, N928, N929, N930, N931, N932, N933, N934, N935,
         N936, N937, N938, N939, N940, N941, N942, N943, N944, N945, N946,
         N947, N948, N949, N950, N951, N952, N953, N954, N955, N956, N957,
         N958, N959, N960, N961, N962, N963, N964, N965, N966, N967, N968,
         N969, N970, N971, N972, N973, N974, N975, N976, N977, N978, N979,
         N980, N981, N982, N983, N984, N985, N986, N987, N988, N989, N990,
         N991, N992, N993, N994, N995, N996, N997, N998, N999, N1000, N1001,
         N1002, N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011,
         N1012, N1013, N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021,
         N1022;
  wire   [1022:0] g;
  wire   [1023:0] p;
  wire   [1023:1] c;

  XOR2D0 C9218 ( .A1(p[0]), .A2(cin), .Z(s[0]) );
  XOR2D0 C9217 ( .A1(p[1]), .A2(c[1]), .Z(s[1]) );
  XOR2D0 C9216 ( .A1(p[2]), .A2(c[2]), .Z(s[2]) );
  XOR2D0 C9215 ( .A1(p[3]), .A2(c[3]), .Z(s[3]) );
  XOR2D0 C9214 ( .A1(p[4]), .A2(c[4]), .Z(s[4]) );
  XOR2D0 C9213 ( .A1(p[5]), .A2(c[5]), .Z(s[5]) );
  XOR2D0 C9212 ( .A1(p[6]), .A2(c[6]), .Z(s[6]) );
  XOR2D0 C9211 ( .A1(p[7]), .A2(c[7]), .Z(s[7]) );
  XOR2D0 C9210 ( .A1(p[8]), .A2(c[8]), .Z(s[8]) );
  XOR2D0 C9209 ( .A1(p[9]), .A2(c[9]), .Z(s[9]) );
  XOR2D0 C9208 ( .A1(p[10]), .A2(c[10]), .Z(s[10]) );
  XOR2D0 C9207 ( .A1(p[11]), .A2(c[11]), .Z(s[11]) );
  XOR2D0 C9206 ( .A1(p[12]), .A2(c[12]), .Z(s[12]) );
  XOR2D0 C9205 ( .A1(p[13]), .A2(c[13]), .Z(s[13]) );
  XOR2D0 C9204 ( .A1(p[14]), .A2(c[14]), .Z(s[14]) );
  XOR2D0 C9203 ( .A1(p[15]), .A2(c[15]), .Z(s[15]) );
  XOR2D0 C9202 ( .A1(p[16]), .A2(c[16]), .Z(s[16]) );
  XOR2D0 C9201 ( .A1(p[17]), .A2(c[17]), .Z(s[17]) );
  XOR2D0 C9200 ( .A1(p[18]), .A2(c[18]), .Z(s[18]) );
  XOR2D0 C9199 ( .A1(p[19]), .A2(c[19]), .Z(s[19]) );
  XOR2D0 C9198 ( .A1(p[20]), .A2(c[20]), .Z(s[20]) );
  XOR2D0 C9197 ( .A1(p[21]), .A2(c[21]), .Z(s[21]) );
  XOR2D0 C9196 ( .A1(p[22]), .A2(c[22]), .Z(s[22]) );
  XOR2D0 C9195 ( .A1(p[23]), .A2(c[23]), .Z(s[23]) );
  XOR2D0 C9194 ( .A1(p[24]), .A2(c[24]), .Z(s[24]) );
  XOR2D0 C9193 ( .A1(p[25]), .A2(c[25]), .Z(s[25]) );
  XOR2D0 C9192 ( .A1(p[26]), .A2(c[26]), .Z(s[26]) );
  XOR2D0 C9191 ( .A1(p[27]), .A2(c[27]), .Z(s[27]) );
  XOR2D0 C9190 ( .A1(p[28]), .A2(c[28]), .Z(s[28]) );
  XOR2D0 C9189 ( .A1(p[29]), .A2(c[29]), .Z(s[29]) );
  XOR2D0 C9188 ( .A1(p[30]), .A2(c[30]), .Z(s[30]) );
  XOR2D0 C9187 ( .A1(p[31]), .A2(c[31]), .Z(s[31]) );
  XOR2D0 C9186 ( .A1(p[32]), .A2(c[32]), .Z(s[32]) );
  XOR2D0 C9185 ( .A1(p[33]), .A2(c[33]), .Z(s[33]) );
  XOR2D0 C9184 ( .A1(p[34]), .A2(c[34]), .Z(s[34]) );
  XOR2D0 C9183 ( .A1(p[35]), .A2(c[35]), .Z(s[35]) );
  XOR2D0 C9182 ( .A1(p[36]), .A2(c[36]), .Z(s[36]) );
  XOR2D0 C9181 ( .A1(p[37]), .A2(c[37]), .Z(s[37]) );
  XOR2D0 C9180 ( .A1(p[38]), .A2(c[38]), .Z(s[38]) );
  XOR2D0 C9179 ( .A1(p[39]), .A2(c[39]), .Z(s[39]) );
  XOR2D0 C9178 ( .A1(p[40]), .A2(c[40]), .Z(s[40]) );
  XOR2D0 C9177 ( .A1(p[41]), .A2(c[41]), .Z(s[41]) );
  XOR2D0 C9176 ( .A1(p[42]), .A2(c[42]), .Z(s[42]) );
  XOR2D0 C9175 ( .A1(p[43]), .A2(c[43]), .Z(s[43]) );
  XOR2D0 C9174 ( .A1(p[44]), .A2(c[44]), .Z(s[44]) );
  XOR2D0 C9173 ( .A1(p[45]), .A2(c[45]), .Z(s[45]) );
  XOR2D0 C9172 ( .A1(p[46]), .A2(c[46]), .Z(s[46]) );
  XOR2D0 C9171 ( .A1(p[47]), .A2(c[47]), .Z(s[47]) );
  XOR2D0 C9170 ( .A1(p[48]), .A2(c[48]), .Z(s[48]) );
  XOR2D0 C9169 ( .A1(p[49]), .A2(c[49]), .Z(s[49]) );
  XOR2D0 C9168 ( .A1(p[50]), .A2(c[50]), .Z(s[50]) );
  XOR2D0 C9167 ( .A1(p[51]), .A2(c[51]), .Z(s[51]) );
  XOR2D0 C9166 ( .A1(p[52]), .A2(c[52]), .Z(s[52]) );
  XOR2D0 C9165 ( .A1(p[53]), .A2(c[53]), .Z(s[53]) );
  XOR2D0 C9164 ( .A1(p[54]), .A2(c[54]), .Z(s[54]) );
  XOR2D0 C9163 ( .A1(p[55]), .A2(c[55]), .Z(s[55]) );
  XOR2D0 C9162 ( .A1(p[56]), .A2(c[56]), .Z(s[56]) );
  XOR2D0 C9161 ( .A1(p[57]), .A2(c[57]), .Z(s[57]) );
  XOR2D0 C9160 ( .A1(p[58]), .A2(c[58]), .Z(s[58]) );
  XOR2D0 C9159 ( .A1(p[59]), .A2(c[59]), .Z(s[59]) );
  XOR2D0 C9158 ( .A1(p[60]), .A2(c[60]), .Z(s[60]) );
  XOR2D0 C9157 ( .A1(p[61]), .A2(c[61]), .Z(s[61]) );
  XOR2D0 C9156 ( .A1(p[62]), .A2(c[62]), .Z(s[62]) );
  XOR2D0 C9155 ( .A1(p[63]), .A2(c[63]), .Z(s[63]) );
  XOR2D0 C9154 ( .A1(p[64]), .A2(c[64]), .Z(s[64]) );
  XOR2D0 C9153 ( .A1(p[65]), .A2(c[65]), .Z(s[65]) );
  XOR2D0 C9152 ( .A1(p[66]), .A2(c[66]), .Z(s[66]) );
  XOR2D0 C9151 ( .A1(p[67]), .A2(c[67]), .Z(s[67]) );
  XOR2D0 C9150 ( .A1(p[68]), .A2(c[68]), .Z(s[68]) );
  XOR2D0 C9149 ( .A1(p[69]), .A2(c[69]), .Z(s[69]) );
  XOR2D0 C9148 ( .A1(p[70]), .A2(c[70]), .Z(s[70]) );
  XOR2D0 C9147 ( .A1(p[71]), .A2(c[71]), .Z(s[71]) );
  XOR2D0 C9146 ( .A1(p[72]), .A2(c[72]), .Z(s[72]) );
  XOR2D0 C9145 ( .A1(p[73]), .A2(c[73]), .Z(s[73]) );
  XOR2D0 C9144 ( .A1(p[74]), .A2(c[74]), .Z(s[74]) );
  XOR2D0 C9143 ( .A1(p[75]), .A2(c[75]), .Z(s[75]) );
  XOR2D0 C9142 ( .A1(p[76]), .A2(c[76]), .Z(s[76]) );
  XOR2D0 C9141 ( .A1(p[77]), .A2(c[77]), .Z(s[77]) );
  XOR2D0 C9140 ( .A1(p[78]), .A2(c[78]), .Z(s[78]) );
  XOR2D0 C9139 ( .A1(p[79]), .A2(c[79]), .Z(s[79]) );
  XOR2D0 C9138 ( .A1(p[80]), .A2(c[80]), .Z(s[80]) );
  XOR2D0 C9137 ( .A1(p[81]), .A2(c[81]), .Z(s[81]) );
  XOR2D0 C9136 ( .A1(p[82]), .A2(c[82]), .Z(s[82]) );
  XOR2D0 C9135 ( .A1(p[83]), .A2(c[83]), .Z(s[83]) );
  XOR2D0 C9134 ( .A1(p[84]), .A2(c[84]), .Z(s[84]) );
  XOR2D0 C9133 ( .A1(p[85]), .A2(c[85]), .Z(s[85]) );
  XOR2D0 C9132 ( .A1(p[86]), .A2(c[86]), .Z(s[86]) );
  XOR2D0 C9131 ( .A1(p[87]), .A2(c[87]), .Z(s[87]) );
  XOR2D0 C9130 ( .A1(p[88]), .A2(c[88]), .Z(s[88]) );
  XOR2D0 C9129 ( .A1(p[89]), .A2(c[89]), .Z(s[89]) );
  XOR2D0 C9128 ( .A1(p[90]), .A2(c[90]), .Z(s[90]) );
  XOR2D0 C9127 ( .A1(p[91]), .A2(c[91]), .Z(s[91]) );
  XOR2D0 C9126 ( .A1(p[92]), .A2(c[92]), .Z(s[92]) );
  XOR2D0 C9125 ( .A1(p[93]), .A2(c[93]), .Z(s[93]) );
  XOR2D0 C9124 ( .A1(p[94]), .A2(c[94]), .Z(s[94]) );
  XOR2D0 C9123 ( .A1(p[95]), .A2(c[95]), .Z(s[95]) );
  XOR2D0 C9122 ( .A1(p[96]), .A2(c[96]), .Z(s[96]) );
  XOR2D0 C9121 ( .A1(p[97]), .A2(c[97]), .Z(s[97]) );
  XOR2D0 C9120 ( .A1(p[98]), .A2(c[98]), .Z(s[98]) );
  XOR2D0 C9119 ( .A1(p[99]), .A2(c[99]), .Z(s[99]) );
  XOR2D0 C9118 ( .A1(p[100]), .A2(c[100]), .Z(s[100]) );
  XOR2D0 C9117 ( .A1(p[101]), .A2(c[101]), .Z(s[101]) );
  XOR2D0 C9116 ( .A1(p[102]), .A2(c[102]), .Z(s[102]) );
  XOR2D0 C9115 ( .A1(p[103]), .A2(c[103]), .Z(s[103]) );
  XOR2D0 C9114 ( .A1(p[104]), .A2(c[104]), .Z(s[104]) );
  XOR2D0 C9113 ( .A1(p[105]), .A2(c[105]), .Z(s[105]) );
  XOR2D0 C9112 ( .A1(p[106]), .A2(c[106]), .Z(s[106]) );
  XOR2D0 C9111 ( .A1(p[107]), .A2(c[107]), .Z(s[107]) );
  XOR2D0 C9110 ( .A1(p[108]), .A2(c[108]), .Z(s[108]) );
  XOR2D0 C9109 ( .A1(p[109]), .A2(c[109]), .Z(s[109]) );
  XOR2D0 C9108 ( .A1(p[110]), .A2(c[110]), .Z(s[110]) );
  XOR2D0 C9107 ( .A1(p[111]), .A2(c[111]), .Z(s[111]) );
  XOR2D0 C9106 ( .A1(p[112]), .A2(c[112]), .Z(s[112]) );
  XOR2D0 C9105 ( .A1(p[113]), .A2(c[113]), .Z(s[113]) );
  XOR2D0 C9104 ( .A1(p[114]), .A2(c[114]), .Z(s[114]) );
  XOR2D0 C9103 ( .A1(p[115]), .A2(c[115]), .Z(s[115]) );
  XOR2D0 C9102 ( .A1(p[116]), .A2(c[116]), .Z(s[116]) );
  XOR2D0 C9101 ( .A1(p[117]), .A2(c[117]), .Z(s[117]) );
  XOR2D0 C9100 ( .A1(p[118]), .A2(c[118]), .Z(s[118]) );
  XOR2D0 C9099 ( .A1(p[119]), .A2(c[119]), .Z(s[119]) );
  XOR2D0 C9098 ( .A1(p[120]), .A2(c[120]), .Z(s[120]) );
  XOR2D0 C9097 ( .A1(p[121]), .A2(c[121]), .Z(s[121]) );
  XOR2D0 C9096 ( .A1(p[122]), .A2(c[122]), .Z(s[122]) );
  XOR2D0 C9095 ( .A1(p[123]), .A2(c[123]), .Z(s[123]) );
  XOR2D0 C9094 ( .A1(p[124]), .A2(c[124]), .Z(s[124]) );
  XOR2D0 C9093 ( .A1(p[125]), .A2(c[125]), .Z(s[125]) );
  XOR2D0 C9092 ( .A1(p[126]), .A2(c[126]), .Z(s[126]) );
  XOR2D0 C9091 ( .A1(p[127]), .A2(c[127]), .Z(s[127]) );
  XOR2D0 C9090 ( .A1(p[128]), .A2(c[128]), .Z(s[128]) );
  XOR2D0 C9089 ( .A1(p[129]), .A2(c[129]), .Z(s[129]) );
  XOR2D0 C9088 ( .A1(p[130]), .A2(c[130]), .Z(s[130]) );
  XOR2D0 C9087 ( .A1(p[131]), .A2(c[131]), .Z(s[131]) );
  XOR2D0 C9086 ( .A1(p[132]), .A2(c[132]), .Z(s[132]) );
  XOR2D0 C9085 ( .A1(p[133]), .A2(c[133]), .Z(s[133]) );
  XOR2D0 C9084 ( .A1(p[134]), .A2(c[134]), .Z(s[134]) );
  XOR2D0 C9083 ( .A1(p[135]), .A2(c[135]), .Z(s[135]) );
  XOR2D0 C9082 ( .A1(p[136]), .A2(c[136]), .Z(s[136]) );
  XOR2D0 C9081 ( .A1(p[137]), .A2(c[137]), .Z(s[137]) );
  XOR2D0 C9080 ( .A1(p[138]), .A2(c[138]), .Z(s[138]) );
  XOR2D0 C9079 ( .A1(p[139]), .A2(c[139]), .Z(s[139]) );
  XOR2D0 C9078 ( .A1(p[140]), .A2(c[140]), .Z(s[140]) );
  XOR2D0 C9077 ( .A1(p[141]), .A2(c[141]), .Z(s[141]) );
  XOR2D0 C9076 ( .A1(p[142]), .A2(c[142]), .Z(s[142]) );
  XOR2D0 C9075 ( .A1(p[143]), .A2(c[143]), .Z(s[143]) );
  XOR2D0 C9074 ( .A1(p[144]), .A2(c[144]), .Z(s[144]) );
  XOR2D0 C9073 ( .A1(p[145]), .A2(c[145]), .Z(s[145]) );
  XOR2D0 C9072 ( .A1(p[146]), .A2(c[146]), .Z(s[146]) );
  XOR2D0 C9071 ( .A1(p[147]), .A2(c[147]), .Z(s[147]) );
  XOR2D0 C9070 ( .A1(p[148]), .A2(c[148]), .Z(s[148]) );
  XOR2D0 C9069 ( .A1(p[149]), .A2(c[149]), .Z(s[149]) );
  XOR2D0 C9068 ( .A1(p[150]), .A2(c[150]), .Z(s[150]) );
  XOR2D0 C9067 ( .A1(p[151]), .A2(c[151]), .Z(s[151]) );
  XOR2D0 C9066 ( .A1(p[152]), .A2(c[152]), .Z(s[152]) );
  XOR2D0 C9065 ( .A1(p[153]), .A2(c[153]), .Z(s[153]) );
  XOR2D0 C9064 ( .A1(p[154]), .A2(c[154]), .Z(s[154]) );
  XOR2D0 C9063 ( .A1(p[155]), .A2(c[155]), .Z(s[155]) );
  XOR2D0 C9062 ( .A1(p[156]), .A2(c[156]), .Z(s[156]) );
  XOR2D0 C9061 ( .A1(p[157]), .A2(c[157]), .Z(s[157]) );
  XOR2D0 C9060 ( .A1(p[158]), .A2(c[158]), .Z(s[158]) );
  XOR2D0 C9059 ( .A1(p[159]), .A2(c[159]), .Z(s[159]) );
  XOR2D0 C9058 ( .A1(p[160]), .A2(c[160]), .Z(s[160]) );
  XOR2D0 C9057 ( .A1(p[161]), .A2(c[161]), .Z(s[161]) );
  XOR2D0 C9056 ( .A1(p[162]), .A2(c[162]), .Z(s[162]) );
  XOR2D0 C9055 ( .A1(p[163]), .A2(c[163]), .Z(s[163]) );
  XOR2D0 C9054 ( .A1(p[164]), .A2(c[164]), .Z(s[164]) );
  XOR2D0 C9053 ( .A1(p[165]), .A2(c[165]), .Z(s[165]) );
  XOR2D0 C9052 ( .A1(p[166]), .A2(c[166]), .Z(s[166]) );
  XOR2D0 C9051 ( .A1(p[167]), .A2(c[167]), .Z(s[167]) );
  XOR2D0 C9050 ( .A1(p[168]), .A2(c[168]), .Z(s[168]) );
  XOR2D0 C9049 ( .A1(p[169]), .A2(c[169]), .Z(s[169]) );
  XOR2D0 C9048 ( .A1(p[170]), .A2(c[170]), .Z(s[170]) );
  XOR2D0 C9047 ( .A1(p[171]), .A2(c[171]), .Z(s[171]) );
  XOR2D0 C9046 ( .A1(p[172]), .A2(c[172]), .Z(s[172]) );
  XOR2D0 C9045 ( .A1(p[173]), .A2(c[173]), .Z(s[173]) );
  XOR2D0 C9044 ( .A1(p[174]), .A2(c[174]), .Z(s[174]) );
  XOR2D0 C9043 ( .A1(p[175]), .A2(c[175]), .Z(s[175]) );
  XOR2D0 C9042 ( .A1(p[176]), .A2(c[176]), .Z(s[176]) );
  XOR2D0 C9041 ( .A1(p[177]), .A2(c[177]), .Z(s[177]) );
  XOR2D0 C9040 ( .A1(p[178]), .A2(c[178]), .Z(s[178]) );
  XOR2D0 C9039 ( .A1(p[179]), .A2(c[179]), .Z(s[179]) );
  XOR2D0 C9038 ( .A1(p[180]), .A2(c[180]), .Z(s[180]) );
  XOR2D0 C9037 ( .A1(p[181]), .A2(c[181]), .Z(s[181]) );
  XOR2D0 C9036 ( .A1(p[182]), .A2(c[182]), .Z(s[182]) );
  XOR2D0 C9035 ( .A1(p[183]), .A2(c[183]), .Z(s[183]) );
  XOR2D0 C9034 ( .A1(p[184]), .A2(c[184]), .Z(s[184]) );
  XOR2D0 C9033 ( .A1(p[185]), .A2(c[185]), .Z(s[185]) );
  XOR2D0 C9032 ( .A1(p[186]), .A2(c[186]), .Z(s[186]) );
  XOR2D0 C9031 ( .A1(p[187]), .A2(c[187]), .Z(s[187]) );
  XOR2D0 C9030 ( .A1(p[188]), .A2(c[188]), .Z(s[188]) );
  XOR2D0 C9029 ( .A1(p[189]), .A2(c[189]), .Z(s[189]) );
  XOR2D0 C9028 ( .A1(p[190]), .A2(c[190]), .Z(s[190]) );
  XOR2D0 C9027 ( .A1(p[191]), .A2(c[191]), .Z(s[191]) );
  XOR2D0 C9026 ( .A1(p[192]), .A2(c[192]), .Z(s[192]) );
  XOR2D0 C9025 ( .A1(p[193]), .A2(c[193]), .Z(s[193]) );
  XOR2D0 C9024 ( .A1(p[194]), .A2(c[194]), .Z(s[194]) );
  XOR2D0 C9023 ( .A1(p[195]), .A2(c[195]), .Z(s[195]) );
  XOR2D0 C9022 ( .A1(p[196]), .A2(c[196]), .Z(s[196]) );
  XOR2D0 C9021 ( .A1(p[197]), .A2(c[197]), .Z(s[197]) );
  XOR2D0 C9020 ( .A1(p[198]), .A2(c[198]), .Z(s[198]) );
  XOR2D0 C9019 ( .A1(p[199]), .A2(c[199]), .Z(s[199]) );
  XOR2D0 C9018 ( .A1(p[200]), .A2(c[200]), .Z(s[200]) );
  XOR2D0 C9017 ( .A1(p[201]), .A2(c[201]), .Z(s[201]) );
  XOR2D0 C9016 ( .A1(p[202]), .A2(c[202]), .Z(s[202]) );
  XOR2D0 C9015 ( .A1(p[203]), .A2(c[203]), .Z(s[203]) );
  XOR2D0 C9014 ( .A1(p[204]), .A2(c[204]), .Z(s[204]) );
  XOR2D0 C9013 ( .A1(p[205]), .A2(c[205]), .Z(s[205]) );
  XOR2D0 C9012 ( .A1(p[206]), .A2(c[206]), .Z(s[206]) );
  XOR2D0 C9011 ( .A1(p[207]), .A2(c[207]), .Z(s[207]) );
  XOR2D0 C9010 ( .A1(p[208]), .A2(c[208]), .Z(s[208]) );
  XOR2D0 C9009 ( .A1(p[209]), .A2(c[209]), .Z(s[209]) );
  XOR2D0 C9008 ( .A1(p[210]), .A2(c[210]), .Z(s[210]) );
  XOR2D0 C9007 ( .A1(p[211]), .A2(c[211]), .Z(s[211]) );
  XOR2D0 C9006 ( .A1(p[212]), .A2(c[212]), .Z(s[212]) );
  XOR2D0 C9005 ( .A1(p[213]), .A2(c[213]), .Z(s[213]) );
  XOR2D0 C9004 ( .A1(p[214]), .A2(c[214]), .Z(s[214]) );
  XOR2D0 C9003 ( .A1(p[215]), .A2(c[215]), .Z(s[215]) );
  XOR2D0 C9002 ( .A1(p[216]), .A2(c[216]), .Z(s[216]) );
  XOR2D0 C9001 ( .A1(p[217]), .A2(c[217]), .Z(s[217]) );
  XOR2D0 C9000 ( .A1(p[218]), .A2(c[218]), .Z(s[218]) );
  XOR2D0 C8999 ( .A1(p[219]), .A2(c[219]), .Z(s[219]) );
  XOR2D0 C8998 ( .A1(p[220]), .A2(c[220]), .Z(s[220]) );
  XOR2D0 C8997 ( .A1(p[221]), .A2(c[221]), .Z(s[221]) );
  XOR2D0 C8996 ( .A1(p[222]), .A2(c[222]), .Z(s[222]) );
  XOR2D0 C8995 ( .A1(p[223]), .A2(c[223]), .Z(s[223]) );
  XOR2D0 C8994 ( .A1(p[224]), .A2(c[224]), .Z(s[224]) );
  XOR2D0 C8993 ( .A1(p[225]), .A2(c[225]), .Z(s[225]) );
  XOR2D0 C8992 ( .A1(p[226]), .A2(c[226]), .Z(s[226]) );
  XOR2D0 C8991 ( .A1(p[227]), .A2(c[227]), .Z(s[227]) );
  XOR2D0 C8990 ( .A1(p[228]), .A2(c[228]), .Z(s[228]) );
  XOR2D0 C8989 ( .A1(p[229]), .A2(c[229]), .Z(s[229]) );
  XOR2D0 C8988 ( .A1(p[230]), .A2(c[230]), .Z(s[230]) );
  XOR2D0 C8987 ( .A1(p[231]), .A2(c[231]), .Z(s[231]) );
  XOR2D0 C8986 ( .A1(p[232]), .A2(c[232]), .Z(s[232]) );
  XOR2D0 C8985 ( .A1(p[233]), .A2(c[233]), .Z(s[233]) );
  XOR2D0 C8984 ( .A1(p[234]), .A2(c[234]), .Z(s[234]) );
  XOR2D0 C8983 ( .A1(p[235]), .A2(c[235]), .Z(s[235]) );
  XOR2D0 C8982 ( .A1(p[236]), .A2(c[236]), .Z(s[236]) );
  XOR2D0 C8981 ( .A1(p[237]), .A2(c[237]), .Z(s[237]) );
  XOR2D0 C8980 ( .A1(p[238]), .A2(c[238]), .Z(s[238]) );
  XOR2D0 C8979 ( .A1(p[239]), .A2(c[239]), .Z(s[239]) );
  XOR2D0 C8978 ( .A1(p[240]), .A2(c[240]), .Z(s[240]) );
  XOR2D0 C8977 ( .A1(p[241]), .A2(c[241]), .Z(s[241]) );
  XOR2D0 C8976 ( .A1(p[242]), .A2(c[242]), .Z(s[242]) );
  XOR2D0 C8975 ( .A1(p[243]), .A2(c[243]), .Z(s[243]) );
  XOR2D0 C8974 ( .A1(p[244]), .A2(c[244]), .Z(s[244]) );
  XOR2D0 C8973 ( .A1(p[245]), .A2(c[245]), .Z(s[245]) );
  XOR2D0 C8972 ( .A1(p[246]), .A2(c[246]), .Z(s[246]) );
  XOR2D0 C8971 ( .A1(p[247]), .A2(c[247]), .Z(s[247]) );
  XOR2D0 C8970 ( .A1(p[248]), .A2(c[248]), .Z(s[248]) );
  XOR2D0 C8969 ( .A1(p[249]), .A2(c[249]), .Z(s[249]) );
  XOR2D0 C8968 ( .A1(p[250]), .A2(c[250]), .Z(s[250]) );
  XOR2D0 C8967 ( .A1(p[251]), .A2(c[251]), .Z(s[251]) );
  XOR2D0 C8966 ( .A1(p[252]), .A2(c[252]), .Z(s[252]) );
  XOR2D0 C8965 ( .A1(p[253]), .A2(c[253]), .Z(s[253]) );
  XOR2D0 C8964 ( .A1(p[254]), .A2(c[254]), .Z(s[254]) );
  XOR2D0 C8963 ( .A1(p[255]), .A2(c[255]), .Z(s[255]) );
  XOR2D0 C8962 ( .A1(p[256]), .A2(c[256]), .Z(s[256]) );
  XOR2D0 C8961 ( .A1(p[257]), .A2(c[257]), .Z(s[257]) );
  XOR2D0 C8960 ( .A1(p[258]), .A2(c[258]), .Z(s[258]) );
  XOR2D0 C8959 ( .A1(p[259]), .A2(c[259]), .Z(s[259]) );
  XOR2D0 C8958 ( .A1(p[260]), .A2(c[260]), .Z(s[260]) );
  XOR2D0 C8957 ( .A1(p[261]), .A2(c[261]), .Z(s[261]) );
  XOR2D0 C8956 ( .A1(p[262]), .A2(c[262]), .Z(s[262]) );
  XOR2D0 C8955 ( .A1(p[263]), .A2(c[263]), .Z(s[263]) );
  XOR2D0 C8954 ( .A1(p[264]), .A2(c[264]), .Z(s[264]) );
  XOR2D0 C8953 ( .A1(p[265]), .A2(c[265]), .Z(s[265]) );
  XOR2D0 C8952 ( .A1(p[266]), .A2(c[266]), .Z(s[266]) );
  XOR2D0 C8951 ( .A1(p[267]), .A2(c[267]), .Z(s[267]) );
  XOR2D0 C8950 ( .A1(p[268]), .A2(c[268]), .Z(s[268]) );
  XOR2D0 C8949 ( .A1(p[269]), .A2(c[269]), .Z(s[269]) );
  XOR2D0 C8948 ( .A1(p[270]), .A2(c[270]), .Z(s[270]) );
  XOR2D0 C8947 ( .A1(p[271]), .A2(c[271]), .Z(s[271]) );
  XOR2D0 C8946 ( .A1(p[272]), .A2(c[272]), .Z(s[272]) );
  XOR2D0 C8945 ( .A1(p[273]), .A2(c[273]), .Z(s[273]) );
  XOR2D0 C8944 ( .A1(p[274]), .A2(c[274]), .Z(s[274]) );
  XOR2D0 C8943 ( .A1(p[275]), .A2(c[275]), .Z(s[275]) );
  XOR2D0 C8942 ( .A1(p[276]), .A2(c[276]), .Z(s[276]) );
  XOR2D0 C8941 ( .A1(p[277]), .A2(c[277]), .Z(s[277]) );
  XOR2D0 C8940 ( .A1(p[278]), .A2(c[278]), .Z(s[278]) );
  XOR2D0 C8939 ( .A1(p[279]), .A2(c[279]), .Z(s[279]) );
  XOR2D0 C8938 ( .A1(p[280]), .A2(c[280]), .Z(s[280]) );
  XOR2D0 C8937 ( .A1(p[281]), .A2(c[281]), .Z(s[281]) );
  XOR2D0 C8936 ( .A1(p[282]), .A2(c[282]), .Z(s[282]) );
  XOR2D0 C8935 ( .A1(p[283]), .A2(c[283]), .Z(s[283]) );
  XOR2D0 C8934 ( .A1(p[284]), .A2(c[284]), .Z(s[284]) );
  XOR2D0 C8933 ( .A1(p[285]), .A2(c[285]), .Z(s[285]) );
  XOR2D0 C8932 ( .A1(p[286]), .A2(c[286]), .Z(s[286]) );
  XOR2D0 C8931 ( .A1(p[287]), .A2(c[287]), .Z(s[287]) );
  XOR2D0 C8930 ( .A1(p[288]), .A2(c[288]), .Z(s[288]) );
  XOR2D0 C8929 ( .A1(p[289]), .A2(c[289]), .Z(s[289]) );
  XOR2D0 C8928 ( .A1(p[290]), .A2(c[290]), .Z(s[290]) );
  XOR2D0 C8927 ( .A1(p[291]), .A2(c[291]), .Z(s[291]) );
  XOR2D0 C8926 ( .A1(p[292]), .A2(c[292]), .Z(s[292]) );
  XOR2D0 C8925 ( .A1(p[293]), .A2(c[293]), .Z(s[293]) );
  XOR2D0 C8924 ( .A1(p[294]), .A2(c[294]), .Z(s[294]) );
  XOR2D0 C8923 ( .A1(p[295]), .A2(c[295]), .Z(s[295]) );
  XOR2D0 C8922 ( .A1(p[296]), .A2(c[296]), .Z(s[296]) );
  XOR2D0 C8921 ( .A1(p[297]), .A2(c[297]), .Z(s[297]) );
  XOR2D0 C8920 ( .A1(p[298]), .A2(c[298]), .Z(s[298]) );
  XOR2D0 C8919 ( .A1(p[299]), .A2(c[299]), .Z(s[299]) );
  XOR2D0 C8918 ( .A1(p[300]), .A2(c[300]), .Z(s[300]) );
  XOR2D0 C8917 ( .A1(p[301]), .A2(c[301]), .Z(s[301]) );
  XOR2D0 C8916 ( .A1(p[302]), .A2(c[302]), .Z(s[302]) );
  XOR2D0 C8915 ( .A1(p[303]), .A2(c[303]), .Z(s[303]) );
  XOR2D0 C8914 ( .A1(p[304]), .A2(c[304]), .Z(s[304]) );
  XOR2D0 C8913 ( .A1(p[305]), .A2(c[305]), .Z(s[305]) );
  XOR2D0 C8912 ( .A1(p[306]), .A2(c[306]), .Z(s[306]) );
  XOR2D0 C8911 ( .A1(p[307]), .A2(c[307]), .Z(s[307]) );
  XOR2D0 C8910 ( .A1(p[308]), .A2(c[308]), .Z(s[308]) );
  XOR2D0 C8909 ( .A1(p[309]), .A2(c[309]), .Z(s[309]) );
  XOR2D0 C8908 ( .A1(p[310]), .A2(c[310]), .Z(s[310]) );
  XOR2D0 C8907 ( .A1(p[311]), .A2(c[311]), .Z(s[311]) );
  XOR2D0 C8906 ( .A1(p[312]), .A2(c[312]), .Z(s[312]) );
  XOR2D0 C8905 ( .A1(p[313]), .A2(c[313]), .Z(s[313]) );
  XOR2D0 C8904 ( .A1(p[314]), .A2(c[314]), .Z(s[314]) );
  XOR2D0 C8903 ( .A1(p[315]), .A2(c[315]), .Z(s[315]) );
  XOR2D0 C8902 ( .A1(p[316]), .A2(c[316]), .Z(s[316]) );
  XOR2D0 C8901 ( .A1(p[317]), .A2(c[317]), .Z(s[317]) );
  XOR2D0 C8900 ( .A1(p[318]), .A2(c[318]), .Z(s[318]) );
  XOR2D0 C8899 ( .A1(p[319]), .A2(c[319]), .Z(s[319]) );
  XOR2D0 C8898 ( .A1(p[320]), .A2(c[320]), .Z(s[320]) );
  XOR2D0 C8897 ( .A1(p[321]), .A2(c[321]), .Z(s[321]) );
  XOR2D0 C8896 ( .A1(p[322]), .A2(c[322]), .Z(s[322]) );
  XOR2D0 C8895 ( .A1(p[323]), .A2(c[323]), .Z(s[323]) );
  XOR2D0 C8894 ( .A1(p[324]), .A2(c[324]), .Z(s[324]) );
  XOR2D0 C8893 ( .A1(p[325]), .A2(c[325]), .Z(s[325]) );
  XOR2D0 C8892 ( .A1(p[326]), .A2(c[326]), .Z(s[326]) );
  XOR2D0 C8891 ( .A1(p[327]), .A2(c[327]), .Z(s[327]) );
  XOR2D0 C8890 ( .A1(p[328]), .A2(c[328]), .Z(s[328]) );
  XOR2D0 C8889 ( .A1(p[329]), .A2(c[329]), .Z(s[329]) );
  XOR2D0 C8888 ( .A1(p[330]), .A2(c[330]), .Z(s[330]) );
  XOR2D0 C8887 ( .A1(p[331]), .A2(c[331]), .Z(s[331]) );
  XOR2D0 C8886 ( .A1(p[332]), .A2(c[332]), .Z(s[332]) );
  XOR2D0 C8885 ( .A1(p[333]), .A2(c[333]), .Z(s[333]) );
  XOR2D0 C8884 ( .A1(p[334]), .A2(c[334]), .Z(s[334]) );
  XOR2D0 C8883 ( .A1(p[335]), .A2(c[335]), .Z(s[335]) );
  XOR2D0 C8882 ( .A1(p[336]), .A2(c[336]), .Z(s[336]) );
  XOR2D0 C8881 ( .A1(p[337]), .A2(c[337]), .Z(s[337]) );
  XOR2D0 C8880 ( .A1(p[338]), .A2(c[338]), .Z(s[338]) );
  XOR2D0 C8879 ( .A1(p[339]), .A2(c[339]), .Z(s[339]) );
  XOR2D0 C8878 ( .A1(p[340]), .A2(c[340]), .Z(s[340]) );
  XOR2D0 C8877 ( .A1(p[341]), .A2(c[341]), .Z(s[341]) );
  XOR2D0 C8876 ( .A1(p[342]), .A2(c[342]), .Z(s[342]) );
  XOR2D0 C8875 ( .A1(p[343]), .A2(c[343]), .Z(s[343]) );
  XOR2D0 C8874 ( .A1(p[344]), .A2(c[344]), .Z(s[344]) );
  XOR2D0 C8873 ( .A1(p[345]), .A2(c[345]), .Z(s[345]) );
  XOR2D0 C8872 ( .A1(p[346]), .A2(c[346]), .Z(s[346]) );
  XOR2D0 C8871 ( .A1(p[347]), .A2(c[347]), .Z(s[347]) );
  XOR2D0 C8870 ( .A1(p[348]), .A2(c[348]), .Z(s[348]) );
  XOR2D0 C8869 ( .A1(p[349]), .A2(c[349]), .Z(s[349]) );
  XOR2D0 C8868 ( .A1(p[350]), .A2(c[350]), .Z(s[350]) );
  XOR2D0 C8867 ( .A1(p[351]), .A2(c[351]), .Z(s[351]) );
  XOR2D0 C8866 ( .A1(p[352]), .A2(c[352]), .Z(s[352]) );
  XOR2D0 C8865 ( .A1(p[353]), .A2(c[353]), .Z(s[353]) );
  XOR2D0 C8864 ( .A1(p[354]), .A2(c[354]), .Z(s[354]) );
  XOR2D0 C8863 ( .A1(p[355]), .A2(c[355]), .Z(s[355]) );
  XOR2D0 C8862 ( .A1(p[356]), .A2(c[356]), .Z(s[356]) );
  XOR2D0 C8861 ( .A1(p[357]), .A2(c[357]), .Z(s[357]) );
  XOR2D0 C8860 ( .A1(p[358]), .A2(c[358]), .Z(s[358]) );
  XOR2D0 C8859 ( .A1(p[359]), .A2(c[359]), .Z(s[359]) );
  XOR2D0 C8858 ( .A1(p[360]), .A2(c[360]), .Z(s[360]) );
  XOR2D0 C8857 ( .A1(p[361]), .A2(c[361]), .Z(s[361]) );
  XOR2D0 C8856 ( .A1(p[362]), .A2(c[362]), .Z(s[362]) );
  XOR2D0 C8855 ( .A1(p[363]), .A2(c[363]), .Z(s[363]) );
  XOR2D0 C8854 ( .A1(p[364]), .A2(c[364]), .Z(s[364]) );
  XOR2D0 C8853 ( .A1(p[365]), .A2(c[365]), .Z(s[365]) );
  XOR2D0 C8852 ( .A1(p[366]), .A2(c[366]), .Z(s[366]) );
  XOR2D0 C8851 ( .A1(p[367]), .A2(c[367]), .Z(s[367]) );
  XOR2D0 C8850 ( .A1(p[368]), .A2(c[368]), .Z(s[368]) );
  XOR2D0 C8849 ( .A1(p[369]), .A2(c[369]), .Z(s[369]) );
  XOR2D0 C8848 ( .A1(p[370]), .A2(c[370]), .Z(s[370]) );
  XOR2D0 C8847 ( .A1(p[371]), .A2(c[371]), .Z(s[371]) );
  XOR2D0 C8846 ( .A1(p[372]), .A2(c[372]), .Z(s[372]) );
  XOR2D0 C8845 ( .A1(p[373]), .A2(c[373]), .Z(s[373]) );
  XOR2D0 C8844 ( .A1(p[374]), .A2(c[374]), .Z(s[374]) );
  XOR2D0 C8843 ( .A1(p[375]), .A2(c[375]), .Z(s[375]) );
  XOR2D0 C8842 ( .A1(p[376]), .A2(c[376]), .Z(s[376]) );
  XOR2D0 C8841 ( .A1(p[377]), .A2(c[377]), .Z(s[377]) );
  XOR2D0 C8840 ( .A1(p[378]), .A2(c[378]), .Z(s[378]) );
  XOR2D0 C8839 ( .A1(p[379]), .A2(c[379]), .Z(s[379]) );
  XOR2D0 C8838 ( .A1(p[380]), .A2(c[380]), .Z(s[380]) );
  XOR2D0 C8837 ( .A1(p[381]), .A2(c[381]), .Z(s[381]) );
  XOR2D0 C8836 ( .A1(p[382]), .A2(c[382]), .Z(s[382]) );
  XOR2D0 C8835 ( .A1(p[383]), .A2(c[383]), .Z(s[383]) );
  XOR2D0 C8834 ( .A1(p[384]), .A2(c[384]), .Z(s[384]) );
  XOR2D0 C8833 ( .A1(p[385]), .A2(c[385]), .Z(s[385]) );
  XOR2D0 C8832 ( .A1(p[386]), .A2(c[386]), .Z(s[386]) );
  XOR2D0 C8831 ( .A1(p[387]), .A2(c[387]), .Z(s[387]) );
  XOR2D0 C8830 ( .A1(p[388]), .A2(c[388]), .Z(s[388]) );
  XOR2D0 C8829 ( .A1(p[389]), .A2(c[389]), .Z(s[389]) );
  XOR2D0 C8828 ( .A1(p[390]), .A2(c[390]), .Z(s[390]) );
  XOR2D0 C8827 ( .A1(p[391]), .A2(c[391]), .Z(s[391]) );
  XOR2D0 C8826 ( .A1(p[392]), .A2(c[392]), .Z(s[392]) );
  XOR2D0 C8825 ( .A1(p[393]), .A2(c[393]), .Z(s[393]) );
  XOR2D0 C8824 ( .A1(p[394]), .A2(c[394]), .Z(s[394]) );
  XOR2D0 C8823 ( .A1(p[395]), .A2(c[395]), .Z(s[395]) );
  XOR2D0 C8822 ( .A1(p[396]), .A2(c[396]), .Z(s[396]) );
  XOR2D0 C8821 ( .A1(p[397]), .A2(c[397]), .Z(s[397]) );
  XOR2D0 C8820 ( .A1(p[398]), .A2(c[398]), .Z(s[398]) );
  XOR2D0 C8819 ( .A1(p[399]), .A2(c[399]), .Z(s[399]) );
  XOR2D0 C8818 ( .A1(p[400]), .A2(c[400]), .Z(s[400]) );
  XOR2D0 C8817 ( .A1(p[401]), .A2(c[401]), .Z(s[401]) );
  XOR2D0 C8816 ( .A1(p[402]), .A2(c[402]), .Z(s[402]) );
  XOR2D0 C8815 ( .A1(p[403]), .A2(c[403]), .Z(s[403]) );
  XOR2D0 C8814 ( .A1(p[404]), .A2(c[404]), .Z(s[404]) );
  XOR2D0 C8813 ( .A1(p[405]), .A2(c[405]), .Z(s[405]) );
  XOR2D0 C8812 ( .A1(p[406]), .A2(c[406]), .Z(s[406]) );
  XOR2D0 C8811 ( .A1(p[407]), .A2(c[407]), .Z(s[407]) );
  XOR2D0 C8810 ( .A1(p[408]), .A2(c[408]), .Z(s[408]) );
  XOR2D0 C8809 ( .A1(p[409]), .A2(c[409]), .Z(s[409]) );
  XOR2D0 C8808 ( .A1(p[410]), .A2(c[410]), .Z(s[410]) );
  XOR2D0 C8807 ( .A1(p[411]), .A2(c[411]), .Z(s[411]) );
  XOR2D0 C8806 ( .A1(p[412]), .A2(c[412]), .Z(s[412]) );
  XOR2D0 C8805 ( .A1(p[413]), .A2(c[413]), .Z(s[413]) );
  XOR2D0 C8804 ( .A1(p[414]), .A2(c[414]), .Z(s[414]) );
  XOR2D0 C8803 ( .A1(p[415]), .A2(c[415]), .Z(s[415]) );
  XOR2D0 C8802 ( .A1(p[416]), .A2(c[416]), .Z(s[416]) );
  XOR2D0 C8801 ( .A1(p[417]), .A2(c[417]), .Z(s[417]) );
  XOR2D0 C8800 ( .A1(p[418]), .A2(c[418]), .Z(s[418]) );
  XOR2D0 C8799 ( .A1(p[419]), .A2(c[419]), .Z(s[419]) );
  XOR2D0 C8798 ( .A1(p[420]), .A2(c[420]), .Z(s[420]) );
  XOR2D0 C8797 ( .A1(p[421]), .A2(c[421]), .Z(s[421]) );
  XOR2D0 C8796 ( .A1(p[422]), .A2(c[422]), .Z(s[422]) );
  XOR2D0 C8795 ( .A1(p[423]), .A2(c[423]), .Z(s[423]) );
  XOR2D0 C8794 ( .A1(p[424]), .A2(c[424]), .Z(s[424]) );
  XOR2D0 C8793 ( .A1(p[425]), .A2(c[425]), .Z(s[425]) );
  XOR2D0 C8792 ( .A1(p[426]), .A2(c[426]), .Z(s[426]) );
  XOR2D0 C8791 ( .A1(p[427]), .A2(c[427]), .Z(s[427]) );
  XOR2D0 C8790 ( .A1(p[428]), .A2(c[428]), .Z(s[428]) );
  XOR2D0 C8789 ( .A1(p[429]), .A2(c[429]), .Z(s[429]) );
  XOR2D0 C8788 ( .A1(p[430]), .A2(c[430]), .Z(s[430]) );
  XOR2D0 C8787 ( .A1(p[431]), .A2(c[431]), .Z(s[431]) );
  XOR2D0 C8786 ( .A1(p[432]), .A2(c[432]), .Z(s[432]) );
  XOR2D0 C8785 ( .A1(p[433]), .A2(c[433]), .Z(s[433]) );
  XOR2D0 C8784 ( .A1(p[434]), .A2(c[434]), .Z(s[434]) );
  XOR2D0 C8783 ( .A1(p[435]), .A2(c[435]), .Z(s[435]) );
  XOR2D0 C8782 ( .A1(p[436]), .A2(c[436]), .Z(s[436]) );
  XOR2D0 C8781 ( .A1(p[437]), .A2(c[437]), .Z(s[437]) );
  XOR2D0 C8780 ( .A1(p[438]), .A2(c[438]), .Z(s[438]) );
  XOR2D0 C8779 ( .A1(p[439]), .A2(c[439]), .Z(s[439]) );
  XOR2D0 C8778 ( .A1(p[440]), .A2(c[440]), .Z(s[440]) );
  XOR2D0 C8777 ( .A1(p[441]), .A2(c[441]), .Z(s[441]) );
  XOR2D0 C8776 ( .A1(p[442]), .A2(c[442]), .Z(s[442]) );
  XOR2D0 C8775 ( .A1(p[443]), .A2(c[443]), .Z(s[443]) );
  XOR2D0 C8774 ( .A1(p[444]), .A2(c[444]), .Z(s[444]) );
  XOR2D0 C8773 ( .A1(p[445]), .A2(c[445]), .Z(s[445]) );
  XOR2D0 C8772 ( .A1(p[446]), .A2(c[446]), .Z(s[446]) );
  XOR2D0 C8771 ( .A1(p[447]), .A2(c[447]), .Z(s[447]) );
  XOR2D0 C8770 ( .A1(p[448]), .A2(c[448]), .Z(s[448]) );
  XOR2D0 C8769 ( .A1(p[449]), .A2(c[449]), .Z(s[449]) );
  XOR2D0 C8768 ( .A1(p[450]), .A2(c[450]), .Z(s[450]) );
  XOR2D0 C8767 ( .A1(p[451]), .A2(c[451]), .Z(s[451]) );
  XOR2D0 C8766 ( .A1(p[452]), .A2(c[452]), .Z(s[452]) );
  XOR2D0 C8765 ( .A1(p[453]), .A2(c[453]), .Z(s[453]) );
  XOR2D0 C8764 ( .A1(p[454]), .A2(c[454]), .Z(s[454]) );
  XOR2D0 C8763 ( .A1(p[455]), .A2(c[455]), .Z(s[455]) );
  XOR2D0 C8762 ( .A1(p[456]), .A2(c[456]), .Z(s[456]) );
  XOR2D0 C8761 ( .A1(p[457]), .A2(c[457]), .Z(s[457]) );
  XOR2D0 C8760 ( .A1(p[458]), .A2(c[458]), .Z(s[458]) );
  XOR2D0 C8759 ( .A1(p[459]), .A2(c[459]), .Z(s[459]) );
  XOR2D0 C8758 ( .A1(p[460]), .A2(c[460]), .Z(s[460]) );
  XOR2D0 C8757 ( .A1(p[461]), .A2(c[461]), .Z(s[461]) );
  XOR2D0 C8756 ( .A1(p[462]), .A2(c[462]), .Z(s[462]) );
  XOR2D0 C8755 ( .A1(p[463]), .A2(c[463]), .Z(s[463]) );
  XOR2D0 C8754 ( .A1(p[464]), .A2(c[464]), .Z(s[464]) );
  XOR2D0 C8753 ( .A1(p[465]), .A2(c[465]), .Z(s[465]) );
  XOR2D0 C8752 ( .A1(p[466]), .A2(c[466]), .Z(s[466]) );
  XOR2D0 C8751 ( .A1(p[467]), .A2(c[467]), .Z(s[467]) );
  XOR2D0 C8750 ( .A1(p[468]), .A2(c[468]), .Z(s[468]) );
  XOR2D0 C8749 ( .A1(p[469]), .A2(c[469]), .Z(s[469]) );
  XOR2D0 C8748 ( .A1(p[470]), .A2(c[470]), .Z(s[470]) );
  XOR2D0 C8747 ( .A1(p[471]), .A2(c[471]), .Z(s[471]) );
  XOR2D0 C8746 ( .A1(p[472]), .A2(c[472]), .Z(s[472]) );
  XOR2D0 C8745 ( .A1(p[473]), .A2(c[473]), .Z(s[473]) );
  XOR2D0 C8744 ( .A1(p[474]), .A2(c[474]), .Z(s[474]) );
  XOR2D0 C8743 ( .A1(p[475]), .A2(c[475]), .Z(s[475]) );
  XOR2D0 C8742 ( .A1(p[476]), .A2(c[476]), .Z(s[476]) );
  XOR2D0 C8741 ( .A1(p[477]), .A2(c[477]), .Z(s[477]) );
  XOR2D0 C8740 ( .A1(p[478]), .A2(c[478]), .Z(s[478]) );
  XOR2D0 C8739 ( .A1(p[479]), .A2(c[479]), .Z(s[479]) );
  XOR2D0 C8738 ( .A1(p[480]), .A2(c[480]), .Z(s[480]) );
  XOR2D0 C8737 ( .A1(p[481]), .A2(c[481]), .Z(s[481]) );
  XOR2D0 C8736 ( .A1(p[482]), .A2(c[482]), .Z(s[482]) );
  XOR2D0 C8735 ( .A1(p[483]), .A2(c[483]), .Z(s[483]) );
  XOR2D0 C8734 ( .A1(p[484]), .A2(c[484]), .Z(s[484]) );
  XOR2D0 C8733 ( .A1(p[485]), .A2(c[485]), .Z(s[485]) );
  XOR2D0 C8732 ( .A1(p[486]), .A2(c[486]), .Z(s[486]) );
  XOR2D0 C8731 ( .A1(p[487]), .A2(c[487]), .Z(s[487]) );
  XOR2D0 C8730 ( .A1(p[488]), .A2(c[488]), .Z(s[488]) );
  XOR2D0 C8729 ( .A1(p[489]), .A2(c[489]), .Z(s[489]) );
  XOR2D0 C8728 ( .A1(p[490]), .A2(c[490]), .Z(s[490]) );
  XOR2D0 C8727 ( .A1(p[491]), .A2(c[491]), .Z(s[491]) );
  XOR2D0 C8726 ( .A1(p[492]), .A2(c[492]), .Z(s[492]) );
  XOR2D0 C8725 ( .A1(p[493]), .A2(c[493]), .Z(s[493]) );
  XOR2D0 C8724 ( .A1(p[494]), .A2(c[494]), .Z(s[494]) );
  XOR2D0 C8723 ( .A1(p[495]), .A2(c[495]), .Z(s[495]) );
  XOR2D0 C8722 ( .A1(p[496]), .A2(c[496]), .Z(s[496]) );
  XOR2D0 C8721 ( .A1(p[497]), .A2(c[497]), .Z(s[497]) );
  XOR2D0 C8720 ( .A1(p[498]), .A2(c[498]), .Z(s[498]) );
  XOR2D0 C8719 ( .A1(p[499]), .A2(c[499]), .Z(s[499]) );
  XOR2D0 C8718 ( .A1(p[500]), .A2(c[500]), .Z(s[500]) );
  XOR2D0 C8717 ( .A1(p[501]), .A2(c[501]), .Z(s[501]) );
  XOR2D0 C8716 ( .A1(p[502]), .A2(c[502]), .Z(s[502]) );
  XOR2D0 C8715 ( .A1(p[503]), .A2(c[503]), .Z(s[503]) );
  XOR2D0 C8714 ( .A1(p[504]), .A2(c[504]), .Z(s[504]) );
  XOR2D0 C8713 ( .A1(p[505]), .A2(c[505]), .Z(s[505]) );
  XOR2D0 C8712 ( .A1(p[506]), .A2(c[506]), .Z(s[506]) );
  XOR2D0 C8711 ( .A1(p[507]), .A2(c[507]), .Z(s[507]) );
  XOR2D0 C8710 ( .A1(p[508]), .A2(c[508]), .Z(s[508]) );
  XOR2D0 C8709 ( .A1(p[509]), .A2(c[509]), .Z(s[509]) );
  XOR2D0 C8708 ( .A1(p[510]), .A2(c[510]), .Z(s[510]) );
  XOR2D0 C8707 ( .A1(p[511]), .A2(c[511]), .Z(s[511]) );
  XOR2D0 C8706 ( .A1(p[512]), .A2(c[512]), .Z(s[512]) );
  XOR2D0 C8705 ( .A1(p[513]), .A2(c[513]), .Z(s[513]) );
  XOR2D0 C8704 ( .A1(p[514]), .A2(c[514]), .Z(s[514]) );
  XOR2D0 C8703 ( .A1(p[515]), .A2(c[515]), .Z(s[515]) );
  XOR2D0 C8702 ( .A1(p[516]), .A2(c[516]), .Z(s[516]) );
  XOR2D0 C8701 ( .A1(p[517]), .A2(c[517]), .Z(s[517]) );
  XOR2D0 C8700 ( .A1(p[518]), .A2(c[518]), .Z(s[518]) );
  XOR2D0 C8699 ( .A1(p[519]), .A2(c[519]), .Z(s[519]) );
  XOR2D0 C8698 ( .A1(p[520]), .A2(c[520]), .Z(s[520]) );
  XOR2D0 C8697 ( .A1(p[521]), .A2(c[521]), .Z(s[521]) );
  XOR2D0 C8696 ( .A1(p[522]), .A2(c[522]), .Z(s[522]) );
  XOR2D0 C8695 ( .A1(p[523]), .A2(c[523]), .Z(s[523]) );
  XOR2D0 C8694 ( .A1(p[524]), .A2(c[524]), .Z(s[524]) );
  XOR2D0 C8693 ( .A1(p[525]), .A2(c[525]), .Z(s[525]) );
  XOR2D0 C8692 ( .A1(p[526]), .A2(c[526]), .Z(s[526]) );
  XOR2D0 C8691 ( .A1(p[527]), .A2(c[527]), .Z(s[527]) );
  XOR2D0 C8690 ( .A1(p[528]), .A2(c[528]), .Z(s[528]) );
  XOR2D0 C8689 ( .A1(p[529]), .A2(c[529]), .Z(s[529]) );
  XOR2D0 C8688 ( .A1(p[530]), .A2(c[530]), .Z(s[530]) );
  XOR2D0 C8687 ( .A1(p[531]), .A2(c[531]), .Z(s[531]) );
  XOR2D0 C8686 ( .A1(p[532]), .A2(c[532]), .Z(s[532]) );
  XOR2D0 C8685 ( .A1(p[533]), .A2(c[533]), .Z(s[533]) );
  XOR2D0 C8684 ( .A1(p[534]), .A2(c[534]), .Z(s[534]) );
  XOR2D0 C8683 ( .A1(p[535]), .A2(c[535]), .Z(s[535]) );
  XOR2D0 C8682 ( .A1(p[536]), .A2(c[536]), .Z(s[536]) );
  XOR2D0 C8681 ( .A1(p[537]), .A2(c[537]), .Z(s[537]) );
  XOR2D0 C8680 ( .A1(p[538]), .A2(c[538]), .Z(s[538]) );
  XOR2D0 C8679 ( .A1(p[539]), .A2(c[539]), .Z(s[539]) );
  XOR2D0 C8678 ( .A1(p[540]), .A2(c[540]), .Z(s[540]) );
  XOR2D0 C8677 ( .A1(p[541]), .A2(c[541]), .Z(s[541]) );
  XOR2D0 C8676 ( .A1(p[542]), .A2(c[542]), .Z(s[542]) );
  XOR2D0 C8675 ( .A1(p[543]), .A2(c[543]), .Z(s[543]) );
  XOR2D0 C8674 ( .A1(p[544]), .A2(c[544]), .Z(s[544]) );
  XOR2D0 C8673 ( .A1(p[545]), .A2(c[545]), .Z(s[545]) );
  XOR2D0 C8672 ( .A1(p[546]), .A2(c[546]), .Z(s[546]) );
  XOR2D0 C8671 ( .A1(p[547]), .A2(c[547]), .Z(s[547]) );
  XOR2D0 C8670 ( .A1(p[548]), .A2(c[548]), .Z(s[548]) );
  XOR2D0 C8669 ( .A1(p[549]), .A2(c[549]), .Z(s[549]) );
  XOR2D0 C8668 ( .A1(p[550]), .A2(c[550]), .Z(s[550]) );
  XOR2D0 C8667 ( .A1(p[551]), .A2(c[551]), .Z(s[551]) );
  XOR2D0 C8666 ( .A1(p[552]), .A2(c[552]), .Z(s[552]) );
  XOR2D0 C8665 ( .A1(p[553]), .A2(c[553]), .Z(s[553]) );
  XOR2D0 C8664 ( .A1(p[554]), .A2(c[554]), .Z(s[554]) );
  XOR2D0 C8663 ( .A1(p[555]), .A2(c[555]), .Z(s[555]) );
  XOR2D0 C8662 ( .A1(p[556]), .A2(c[556]), .Z(s[556]) );
  XOR2D0 C8661 ( .A1(p[557]), .A2(c[557]), .Z(s[557]) );
  XOR2D0 C8660 ( .A1(p[558]), .A2(c[558]), .Z(s[558]) );
  XOR2D0 C8659 ( .A1(p[559]), .A2(c[559]), .Z(s[559]) );
  XOR2D0 C8658 ( .A1(p[560]), .A2(c[560]), .Z(s[560]) );
  XOR2D0 C8657 ( .A1(p[561]), .A2(c[561]), .Z(s[561]) );
  XOR2D0 C8656 ( .A1(p[562]), .A2(c[562]), .Z(s[562]) );
  XOR2D0 C8655 ( .A1(p[563]), .A2(c[563]), .Z(s[563]) );
  XOR2D0 C8654 ( .A1(p[564]), .A2(c[564]), .Z(s[564]) );
  XOR2D0 C8653 ( .A1(p[565]), .A2(c[565]), .Z(s[565]) );
  XOR2D0 C8652 ( .A1(p[566]), .A2(c[566]), .Z(s[566]) );
  XOR2D0 C8651 ( .A1(p[567]), .A2(c[567]), .Z(s[567]) );
  XOR2D0 C8650 ( .A1(p[568]), .A2(c[568]), .Z(s[568]) );
  XOR2D0 C8649 ( .A1(p[569]), .A2(c[569]), .Z(s[569]) );
  XOR2D0 C8648 ( .A1(p[570]), .A2(c[570]), .Z(s[570]) );
  XOR2D0 C8647 ( .A1(p[571]), .A2(c[571]), .Z(s[571]) );
  XOR2D0 C8646 ( .A1(p[572]), .A2(c[572]), .Z(s[572]) );
  XOR2D0 C8645 ( .A1(p[573]), .A2(c[573]), .Z(s[573]) );
  XOR2D0 C8644 ( .A1(p[574]), .A2(c[574]), .Z(s[574]) );
  XOR2D0 C8643 ( .A1(p[575]), .A2(c[575]), .Z(s[575]) );
  XOR2D0 C8642 ( .A1(p[576]), .A2(c[576]), .Z(s[576]) );
  XOR2D0 C8641 ( .A1(p[577]), .A2(c[577]), .Z(s[577]) );
  XOR2D0 C8640 ( .A1(p[578]), .A2(c[578]), .Z(s[578]) );
  XOR2D0 C8639 ( .A1(p[579]), .A2(c[579]), .Z(s[579]) );
  XOR2D0 C8638 ( .A1(p[580]), .A2(c[580]), .Z(s[580]) );
  XOR2D0 C8637 ( .A1(p[581]), .A2(c[581]), .Z(s[581]) );
  XOR2D0 C8636 ( .A1(p[582]), .A2(c[582]), .Z(s[582]) );
  XOR2D0 C8635 ( .A1(p[583]), .A2(c[583]), .Z(s[583]) );
  XOR2D0 C8634 ( .A1(p[584]), .A2(c[584]), .Z(s[584]) );
  XOR2D0 C8633 ( .A1(p[585]), .A2(c[585]), .Z(s[585]) );
  XOR2D0 C8632 ( .A1(p[586]), .A2(c[586]), .Z(s[586]) );
  XOR2D0 C8631 ( .A1(p[587]), .A2(c[587]), .Z(s[587]) );
  XOR2D0 C8630 ( .A1(p[588]), .A2(c[588]), .Z(s[588]) );
  XOR2D0 C8629 ( .A1(p[589]), .A2(c[589]), .Z(s[589]) );
  XOR2D0 C8628 ( .A1(p[590]), .A2(c[590]), .Z(s[590]) );
  XOR2D0 C8627 ( .A1(p[591]), .A2(c[591]), .Z(s[591]) );
  XOR2D0 C8626 ( .A1(p[592]), .A2(c[592]), .Z(s[592]) );
  XOR2D0 C8625 ( .A1(p[593]), .A2(c[593]), .Z(s[593]) );
  XOR2D0 C8624 ( .A1(p[594]), .A2(c[594]), .Z(s[594]) );
  XOR2D0 C8623 ( .A1(p[595]), .A2(c[595]), .Z(s[595]) );
  XOR2D0 C8622 ( .A1(p[596]), .A2(c[596]), .Z(s[596]) );
  XOR2D0 C8621 ( .A1(p[597]), .A2(c[597]), .Z(s[597]) );
  XOR2D0 C8620 ( .A1(p[598]), .A2(c[598]), .Z(s[598]) );
  XOR2D0 C8619 ( .A1(p[599]), .A2(c[599]), .Z(s[599]) );
  XOR2D0 C8618 ( .A1(p[600]), .A2(c[600]), .Z(s[600]) );
  XOR2D0 C8617 ( .A1(p[601]), .A2(c[601]), .Z(s[601]) );
  XOR2D0 C8616 ( .A1(p[602]), .A2(c[602]), .Z(s[602]) );
  XOR2D0 C8615 ( .A1(p[603]), .A2(c[603]), .Z(s[603]) );
  XOR2D0 C8614 ( .A1(p[604]), .A2(c[604]), .Z(s[604]) );
  XOR2D0 C8613 ( .A1(p[605]), .A2(c[605]), .Z(s[605]) );
  XOR2D0 C8612 ( .A1(p[606]), .A2(c[606]), .Z(s[606]) );
  XOR2D0 C8611 ( .A1(p[607]), .A2(c[607]), .Z(s[607]) );
  XOR2D0 C8610 ( .A1(p[608]), .A2(c[608]), .Z(s[608]) );
  XOR2D0 C8609 ( .A1(p[609]), .A2(c[609]), .Z(s[609]) );
  XOR2D0 C8608 ( .A1(p[610]), .A2(c[610]), .Z(s[610]) );
  XOR2D0 C8607 ( .A1(p[611]), .A2(c[611]), .Z(s[611]) );
  XOR2D0 C8606 ( .A1(p[612]), .A2(c[612]), .Z(s[612]) );
  XOR2D0 C8605 ( .A1(p[613]), .A2(c[613]), .Z(s[613]) );
  XOR2D0 C8604 ( .A1(p[614]), .A2(c[614]), .Z(s[614]) );
  XOR2D0 C8603 ( .A1(p[615]), .A2(c[615]), .Z(s[615]) );
  XOR2D0 C8602 ( .A1(p[616]), .A2(c[616]), .Z(s[616]) );
  XOR2D0 C8601 ( .A1(p[617]), .A2(c[617]), .Z(s[617]) );
  XOR2D0 C8600 ( .A1(p[618]), .A2(c[618]), .Z(s[618]) );
  XOR2D0 C8599 ( .A1(p[619]), .A2(c[619]), .Z(s[619]) );
  XOR2D0 C8598 ( .A1(p[620]), .A2(c[620]), .Z(s[620]) );
  XOR2D0 C8597 ( .A1(p[621]), .A2(c[621]), .Z(s[621]) );
  XOR2D0 C8596 ( .A1(p[622]), .A2(c[622]), .Z(s[622]) );
  XOR2D0 C8595 ( .A1(p[623]), .A2(c[623]), .Z(s[623]) );
  XOR2D0 C8594 ( .A1(p[624]), .A2(c[624]), .Z(s[624]) );
  XOR2D0 C8593 ( .A1(p[625]), .A2(c[625]), .Z(s[625]) );
  XOR2D0 C8592 ( .A1(p[626]), .A2(c[626]), .Z(s[626]) );
  XOR2D0 C8591 ( .A1(p[627]), .A2(c[627]), .Z(s[627]) );
  XOR2D0 C8590 ( .A1(p[628]), .A2(c[628]), .Z(s[628]) );
  XOR2D0 C8589 ( .A1(p[629]), .A2(c[629]), .Z(s[629]) );
  XOR2D0 C8588 ( .A1(p[630]), .A2(c[630]), .Z(s[630]) );
  XOR2D0 C8587 ( .A1(p[631]), .A2(c[631]), .Z(s[631]) );
  XOR2D0 C8586 ( .A1(p[632]), .A2(c[632]), .Z(s[632]) );
  XOR2D0 C8585 ( .A1(p[633]), .A2(c[633]), .Z(s[633]) );
  XOR2D0 C8584 ( .A1(p[634]), .A2(c[634]), .Z(s[634]) );
  XOR2D0 C8583 ( .A1(p[635]), .A2(c[635]), .Z(s[635]) );
  XOR2D0 C8582 ( .A1(p[636]), .A2(c[636]), .Z(s[636]) );
  XOR2D0 C8581 ( .A1(p[637]), .A2(c[637]), .Z(s[637]) );
  XOR2D0 C8580 ( .A1(p[638]), .A2(c[638]), .Z(s[638]) );
  XOR2D0 C8579 ( .A1(p[639]), .A2(c[639]), .Z(s[639]) );
  XOR2D0 C8578 ( .A1(p[640]), .A2(c[640]), .Z(s[640]) );
  XOR2D0 C8577 ( .A1(p[641]), .A2(c[641]), .Z(s[641]) );
  XOR2D0 C8576 ( .A1(p[642]), .A2(c[642]), .Z(s[642]) );
  XOR2D0 C8575 ( .A1(p[643]), .A2(c[643]), .Z(s[643]) );
  XOR2D0 C8574 ( .A1(p[644]), .A2(c[644]), .Z(s[644]) );
  XOR2D0 C8573 ( .A1(p[645]), .A2(c[645]), .Z(s[645]) );
  XOR2D0 C8572 ( .A1(p[646]), .A2(c[646]), .Z(s[646]) );
  XOR2D0 C8571 ( .A1(p[647]), .A2(c[647]), .Z(s[647]) );
  XOR2D0 C8570 ( .A1(p[648]), .A2(c[648]), .Z(s[648]) );
  XOR2D0 C8569 ( .A1(p[649]), .A2(c[649]), .Z(s[649]) );
  XOR2D0 C8568 ( .A1(p[650]), .A2(c[650]), .Z(s[650]) );
  XOR2D0 C8567 ( .A1(p[651]), .A2(c[651]), .Z(s[651]) );
  XOR2D0 C8566 ( .A1(p[652]), .A2(c[652]), .Z(s[652]) );
  XOR2D0 C8565 ( .A1(p[653]), .A2(c[653]), .Z(s[653]) );
  XOR2D0 C8564 ( .A1(p[654]), .A2(c[654]), .Z(s[654]) );
  XOR2D0 C8563 ( .A1(p[655]), .A2(c[655]), .Z(s[655]) );
  XOR2D0 C8562 ( .A1(p[656]), .A2(c[656]), .Z(s[656]) );
  XOR2D0 C8561 ( .A1(p[657]), .A2(c[657]), .Z(s[657]) );
  XOR2D0 C8560 ( .A1(p[658]), .A2(c[658]), .Z(s[658]) );
  XOR2D0 C8559 ( .A1(p[659]), .A2(c[659]), .Z(s[659]) );
  XOR2D0 C8558 ( .A1(p[660]), .A2(c[660]), .Z(s[660]) );
  XOR2D0 C8557 ( .A1(p[661]), .A2(c[661]), .Z(s[661]) );
  XOR2D0 C8556 ( .A1(p[662]), .A2(c[662]), .Z(s[662]) );
  XOR2D0 C8555 ( .A1(p[663]), .A2(c[663]), .Z(s[663]) );
  XOR2D0 C8554 ( .A1(p[664]), .A2(c[664]), .Z(s[664]) );
  XOR2D0 C8553 ( .A1(p[665]), .A2(c[665]), .Z(s[665]) );
  XOR2D0 C8552 ( .A1(p[666]), .A2(c[666]), .Z(s[666]) );
  XOR2D0 C8551 ( .A1(p[667]), .A2(c[667]), .Z(s[667]) );
  XOR2D0 C8550 ( .A1(p[668]), .A2(c[668]), .Z(s[668]) );
  XOR2D0 C8549 ( .A1(p[669]), .A2(c[669]), .Z(s[669]) );
  XOR2D0 C8548 ( .A1(p[670]), .A2(c[670]), .Z(s[670]) );
  XOR2D0 C8547 ( .A1(p[671]), .A2(c[671]), .Z(s[671]) );
  XOR2D0 C8546 ( .A1(p[672]), .A2(c[672]), .Z(s[672]) );
  XOR2D0 C8545 ( .A1(p[673]), .A2(c[673]), .Z(s[673]) );
  XOR2D0 C8544 ( .A1(p[674]), .A2(c[674]), .Z(s[674]) );
  XOR2D0 C8543 ( .A1(p[675]), .A2(c[675]), .Z(s[675]) );
  XOR2D0 C8542 ( .A1(p[676]), .A2(c[676]), .Z(s[676]) );
  XOR2D0 C8541 ( .A1(p[677]), .A2(c[677]), .Z(s[677]) );
  XOR2D0 C8540 ( .A1(p[678]), .A2(c[678]), .Z(s[678]) );
  XOR2D0 C8539 ( .A1(p[679]), .A2(c[679]), .Z(s[679]) );
  XOR2D0 C8538 ( .A1(p[680]), .A2(c[680]), .Z(s[680]) );
  XOR2D0 C8537 ( .A1(p[681]), .A2(c[681]), .Z(s[681]) );
  XOR2D0 C8536 ( .A1(p[682]), .A2(c[682]), .Z(s[682]) );
  XOR2D0 C8535 ( .A1(p[683]), .A2(c[683]), .Z(s[683]) );
  XOR2D0 C8534 ( .A1(p[684]), .A2(c[684]), .Z(s[684]) );
  XOR2D0 C8533 ( .A1(p[685]), .A2(c[685]), .Z(s[685]) );
  XOR2D0 C8532 ( .A1(p[686]), .A2(c[686]), .Z(s[686]) );
  XOR2D0 C8531 ( .A1(p[687]), .A2(c[687]), .Z(s[687]) );
  XOR2D0 C8530 ( .A1(p[688]), .A2(c[688]), .Z(s[688]) );
  XOR2D0 C8529 ( .A1(p[689]), .A2(c[689]), .Z(s[689]) );
  XOR2D0 C8528 ( .A1(p[690]), .A2(c[690]), .Z(s[690]) );
  XOR2D0 C8527 ( .A1(p[691]), .A2(c[691]), .Z(s[691]) );
  XOR2D0 C8526 ( .A1(p[692]), .A2(c[692]), .Z(s[692]) );
  XOR2D0 C8525 ( .A1(p[693]), .A2(c[693]), .Z(s[693]) );
  XOR2D0 C8524 ( .A1(p[694]), .A2(c[694]), .Z(s[694]) );
  XOR2D0 C8523 ( .A1(p[695]), .A2(c[695]), .Z(s[695]) );
  XOR2D0 C8522 ( .A1(p[696]), .A2(c[696]), .Z(s[696]) );
  XOR2D0 C8521 ( .A1(p[697]), .A2(c[697]), .Z(s[697]) );
  XOR2D0 C8520 ( .A1(p[698]), .A2(c[698]), .Z(s[698]) );
  XOR2D0 C8519 ( .A1(p[699]), .A2(c[699]), .Z(s[699]) );
  XOR2D0 C8518 ( .A1(p[700]), .A2(c[700]), .Z(s[700]) );
  XOR2D0 C8517 ( .A1(p[701]), .A2(c[701]), .Z(s[701]) );
  XOR2D0 C8516 ( .A1(p[702]), .A2(c[702]), .Z(s[702]) );
  XOR2D0 C8515 ( .A1(p[703]), .A2(c[703]), .Z(s[703]) );
  XOR2D0 C8514 ( .A1(p[704]), .A2(c[704]), .Z(s[704]) );
  XOR2D0 C8513 ( .A1(p[705]), .A2(c[705]), .Z(s[705]) );
  XOR2D0 C8512 ( .A1(p[706]), .A2(c[706]), .Z(s[706]) );
  XOR2D0 C8511 ( .A1(p[707]), .A2(c[707]), .Z(s[707]) );
  XOR2D0 C8510 ( .A1(p[708]), .A2(c[708]), .Z(s[708]) );
  XOR2D0 C8509 ( .A1(p[709]), .A2(c[709]), .Z(s[709]) );
  XOR2D0 C8508 ( .A1(p[710]), .A2(c[710]), .Z(s[710]) );
  XOR2D0 C8507 ( .A1(p[711]), .A2(c[711]), .Z(s[711]) );
  XOR2D0 C8506 ( .A1(p[712]), .A2(c[712]), .Z(s[712]) );
  XOR2D0 C8505 ( .A1(p[713]), .A2(c[713]), .Z(s[713]) );
  XOR2D0 C8504 ( .A1(p[714]), .A2(c[714]), .Z(s[714]) );
  XOR2D0 C8503 ( .A1(p[715]), .A2(c[715]), .Z(s[715]) );
  XOR2D0 C8502 ( .A1(p[716]), .A2(c[716]), .Z(s[716]) );
  XOR2D0 C8501 ( .A1(p[717]), .A2(c[717]), .Z(s[717]) );
  XOR2D0 C8500 ( .A1(p[718]), .A2(c[718]), .Z(s[718]) );
  XOR2D0 C8499 ( .A1(p[719]), .A2(c[719]), .Z(s[719]) );
  XOR2D0 C8498 ( .A1(p[720]), .A2(c[720]), .Z(s[720]) );
  XOR2D0 C8497 ( .A1(p[721]), .A2(c[721]), .Z(s[721]) );
  XOR2D0 C8496 ( .A1(p[722]), .A2(c[722]), .Z(s[722]) );
  XOR2D0 C8495 ( .A1(p[723]), .A2(c[723]), .Z(s[723]) );
  XOR2D0 C8494 ( .A1(p[724]), .A2(c[724]), .Z(s[724]) );
  XOR2D0 C8493 ( .A1(p[725]), .A2(c[725]), .Z(s[725]) );
  XOR2D0 C8492 ( .A1(p[726]), .A2(c[726]), .Z(s[726]) );
  XOR2D0 C8491 ( .A1(p[727]), .A2(c[727]), .Z(s[727]) );
  XOR2D0 C8490 ( .A1(p[728]), .A2(c[728]), .Z(s[728]) );
  XOR2D0 C8489 ( .A1(p[729]), .A2(c[729]), .Z(s[729]) );
  XOR2D0 C8488 ( .A1(p[730]), .A2(c[730]), .Z(s[730]) );
  XOR2D0 C8487 ( .A1(p[731]), .A2(c[731]), .Z(s[731]) );
  XOR2D0 C8486 ( .A1(p[732]), .A2(c[732]), .Z(s[732]) );
  XOR2D0 C8485 ( .A1(p[733]), .A2(c[733]), .Z(s[733]) );
  XOR2D0 C8484 ( .A1(p[734]), .A2(c[734]), .Z(s[734]) );
  XOR2D0 C8483 ( .A1(p[735]), .A2(c[735]), .Z(s[735]) );
  XOR2D0 C8482 ( .A1(p[736]), .A2(c[736]), .Z(s[736]) );
  XOR2D0 C8481 ( .A1(p[737]), .A2(c[737]), .Z(s[737]) );
  XOR2D0 C8480 ( .A1(p[738]), .A2(c[738]), .Z(s[738]) );
  XOR2D0 C8479 ( .A1(p[739]), .A2(c[739]), .Z(s[739]) );
  XOR2D0 C8478 ( .A1(p[740]), .A2(c[740]), .Z(s[740]) );
  XOR2D0 C8477 ( .A1(p[741]), .A2(c[741]), .Z(s[741]) );
  XOR2D0 C8476 ( .A1(p[742]), .A2(c[742]), .Z(s[742]) );
  XOR2D0 C8475 ( .A1(p[743]), .A2(c[743]), .Z(s[743]) );
  XOR2D0 C8474 ( .A1(p[744]), .A2(c[744]), .Z(s[744]) );
  XOR2D0 C8473 ( .A1(p[745]), .A2(c[745]), .Z(s[745]) );
  XOR2D0 C8472 ( .A1(p[746]), .A2(c[746]), .Z(s[746]) );
  XOR2D0 C8471 ( .A1(p[747]), .A2(c[747]), .Z(s[747]) );
  XOR2D0 C8470 ( .A1(p[748]), .A2(c[748]), .Z(s[748]) );
  XOR2D0 C8469 ( .A1(p[749]), .A2(c[749]), .Z(s[749]) );
  XOR2D0 C8468 ( .A1(p[750]), .A2(c[750]), .Z(s[750]) );
  XOR2D0 C8467 ( .A1(p[751]), .A2(c[751]), .Z(s[751]) );
  XOR2D0 C8466 ( .A1(p[752]), .A2(c[752]), .Z(s[752]) );
  XOR2D0 C8465 ( .A1(p[753]), .A2(c[753]), .Z(s[753]) );
  XOR2D0 C8464 ( .A1(p[754]), .A2(c[754]), .Z(s[754]) );
  XOR2D0 C8463 ( .A1(p[755]), .A2(c[755]), .Z(s[755]) );
  XOR2D0 C8462 ( .A1(p[756]), .A2(c[756]), .Z(s[756]) );
  XOR2D0 C8461 ( .A1(p[757]), .A2(c[757]), .Z(s[757]) );
  XOR2D0 C8460 ( .A1(p[758]), .A2(c[758]), .Z(s[758]) );
  XOR2D0 C8459 ( .A1(p[759]), .A2(c[759]), .Z(s[759]) );
  XOR2D0 C8458 ( .A1(p[760]), .A2(c[760]), .Z(s[760]) );
  XOR2D0 C8457 ( .A1(p[761]), .A2(c[761]), .Z(s[761]) );
  XOR2D0 C8456 ( .A1(p[762]), .A2(c[762]), .Z(s[762]) );
  XOR2D0 C8455 ( .A1(p[763]), .A2(c[763]), .Z(s[763]) );
  XOR2D0 C8454 ( .A1(p[764]), .A2(c[764]), .Z(s[764]) );
  XOR2D0 C8453 ( .A1(p[765]), .A2(c[765]), .Z(s[765]) );
  XOR2D0 C8452 ( .A1(p[766]), .A2(c[766]), .Z(s[766]) );
  XOR2D0 C8451 ( .A1(p[767]), .A2(c[767]), .Z(s[767]) );
  XOR2D0 C8450 ( .A1(p[768]), .A2(c[768]), .Z(s[768]) );
  XOR2D0 C8449 ( .A1(p[769]), .A2(c[769]), .Z(s[769]) );
  XOR2D0 C8448 ( .A1(p[770]), .A2(c[770]), .Z(s[770]) );
  XOR2D0 C8447 ( .A1(p[771]), .A2(c[771]), .Z(s[771]) );
  XOR2D0 C8446 ( .A1(p[772]), .A2(c[772]), .Z(s[772]) );
  XOR2D0 C8445 ( .A1(p[773]), .A2(c[773]), .Z(s[773]) );
  XOR2D0 C8444 ( .A1(p[774]), .A2(c[774]), .Z(s[774]) );
  XOR2D0 C8443 ( .A1(p[775]), .A2(c[775]), .Z(s[775]) );
  XOR2D0 C8442 ( .A1(p[776]), .A2(c[776]), .Z(s[776]) );
  XOR2D0 C8441 ( .A1(p[777]), .A2(c[777]), .Z(s[777]) );
  XOR2D0 C8440 ( .A1(p[778]), .A2(c[778]), .Z(s[778]) );
  XOR2D0 C8439 ( .A1(p[779]), .A2(c[779]), .Z(s[779]) );
  XOR2D0 C8438 ( .A1(p[780]), .A2(c[780]), .Z(s[780]) );
  XOR2D0 C8437 ( .A1(p[781]), .A2(c[781]), .Z(s[781]) );
  XOR2D0 C8436 ( .A1(p[782]), .A2(c[782]), .Z(s[782]) );
  XOR2D0 C8435 ( .A1(p[783]), .A2(c[783]), .Z(s[783]) );
  XOR2D0 C8434 ( .A1(p[784]), .A2(c[784]), .Z(s[784]) );
  XOR2D0 C8433 ( .A1(p[785]), .A2(c[785]), .Z(s[785]) );
  XOR2D0 C8432 ( .A1(p[786]), .A2(c[786]), .Z(s[786]) );
  XOR2D0 C8431 ( .A1(p[787]), .A2(c[787]), .Z(s[787]) );
  XOR2D0 C8430 ( .A1(p[788]), .A2(c[788]), .Z(s[788]) );
  XOR2D0 C8429 ( .A1(p[789]), .A2(c[789]), .Z(s[789]) );
  XOR2D0 C8428 ( .A1(p[790]), .A2(c[790]), .Z(s[790]) );
  XOR2D0 C8427 ( .A1(p[791]), .A2(c[791]), .Z(s[791]) );
  XOR2D0 C8426 ( .A1(p[792]), .A2(c[792]), .Z(s[792]) );
  XOR2D0 C8425 ( .A1(p[793]), .A2(c[793]), .Z(s[793]) );
  XOR2D0 C8424 ( .A1(p[794]), .A2(c[794]), .Z(s[794]) );
  XOR2D0 C8423 ( .A1(p[795]), .A2(c[795]), .Z(s[795]) );
  XOR2D0 C8422 ( .A1(p[796]), .A2(c[796]), .Z(s[796]) );
  XOR2D0 C8421 ( .A1(p[797]), .A2(c[797]), .Z(s[797]) );
  XOR2D0 C8420 ( .A1(p[798]), .A2(c[798]), .Z(s[798]) );
  XOR2D0 C8419 ( .A1(p[799]), .A2(c[799]), .Z(s[799]) );
  XOR2D0 C8418 ( .A1(p[800]), .A2(c[800]), .Z(s[800]) );
  XOR2D0 C8417 ( .A1(p[801]), .A2(c[801]), .Z(s[801]) );
  XOR2D0 C8416 ( .A1(p[802]), .A2(c[802]), .Z(s[802]) );
  XOR2D0 C8415 ( .A1(p[803]), .A2(c[803]), .Z(s[803]) );
  XOR2D0 C8414 ( .A1(p[804]), .A2(c[804]), .Z(s[804]) );
  XOR2D0 C8413 ( .A1(p[805]), .A2(c[805]), .Z(s[805]) );
  XOR2D0 C8412 ( .A1(p[806]), .A2(c[806]), .Z(s[806]) );
  XOR2D0 C8411 ( .A1(p[807]), .A2(c[807]), .Z(s[807]) );
  XOR2D0 C8410 ( .A1(p[808]), .A2(c[808]), .Z(s[808]) );
  XOR2D0 C8409 ( .A1(p[809]), .A2(c[809]), .Z(s[809]) );
  XOR2D0 C8408 ( .A1(p[810]), .A2(c[810]), .Z(s[810]) );
  XOR2D0 C8407 ( .A1(p[811]), .A2(c[811]), .Z(s[811]) );
  XOR2D0 C8406 ( .A1(p[812]), .A2(c[812]), .Z(s[812]) );
  XOR2D0 C8405 ( .A1(p[813]), .A2(c[813]), .Z(s[813]) );
  XOR2D0 C8404 ( .A1(p[814]), .A2(c[814]), .Z(s[814]) );
  XOR2D0 C8403 ( .A1(p[815]), .A2(c[815]), .Z(s[815]) );
  XOR2D0 C8402 ( .A1(p[816]), .A2(c[816]), .Z(s[816]) );
  XOR2D0 C8401 ( .A1(p[817]), .A2(c[817]), .Z(s[817]) );
  XOR2D0 C8400 ( .A1(p[818]), .A2(c[818]), .Z(s[818]) );
  XOR2D0 C8399 ( .A1(p[819]), .A2(c[819]), .Z(s[819]) );
  XOR2D0 C8398 ( .A1(p[820]), .A2(c[820]), .Z(s[820]) );
  XOR2D0 C8397 ( .A1(p[821]), .A2(c[821]), .Z(s[821]) );
  XOR2D0 C8396 ( .A1(p[822]), .A2(c[822]), .Z(s[822]) );
  XOR2D0 C8395 ( .A1(p[823]), .A2(c[823]), .Z(s[823]) );
  XOR2D0 C8394 ( .A1(p[824]), .A2(c[824]), .Z(s[824]) );
  XOR2D0 C8393 ( .A1(p[825]), .A2(c[825]), .Z(s[825]) );
  XOR2D0 C8392 ( .A1(p[826]), .A2(c[826]), .Z(s[826]) );
  XOR2D0 C8391 ( .A1(p[827]), .A2(c[827]), .Z(s[827]) );
  XOR2D0 C8390 ( .A1(p[828]), .A2(c[828]), .Z(s[828]) );
  XOR2D0 C8389 ( .A1(p[829]), .A2(c[829]), .Z(s[829]) );
  XOR2D0 C8388 ( .A1(p[830]), .A2(c[830]), .Z(s[830]) );
  XOR2D0 C8387 ( .A1(p[831]), .A2(c[831]), .Z(s[831]) );
  XOR2D0 C8386 ( .A1(p[832]), .A2(c[832]), .Z(s[832]) );
  XOR2D0 C8385 ( .A1(p[833]), .A2(c[833]), .Z(s[833]) );
  XOR2D0 C8384 ( .A1(p[834]), .A2(c[834]), .Z(s[834]) );
  XOR2D0 C8383 ( .A1(p[835]), .A2(c[835]), .Z(s[835]) );
  XOR2D0 C8382 ( .A1(p[836]), .A2(c[836]), .Z(s[836]) );
  XOR2D0 C8381 ( .A1(p[837]), .A2(c[837]), .Z(s[837]) );
  XOR2D0 C8380 ( .A1(p[838]), .A2(c[838]), .Z(s[838]) );
  XOR2D0 C8379 ( .A1(p[839]), .A2(c[839]), .Z(s[839]) );
  XOR2D0 C8378 ( .A1(p[840]), .A2(c[840]), .Z(s[840]) );
  XOR2D0 C8377 ( .A1(p[841]), .A2(c[841]), .Z(s[841]) );
  XOR2D0 C8376 ( .A1(p[842]), .A2(c[842]), .Z(s[842]) );
  XOR2D0 C8375 ( .A1(p[843]), .A2(c[843]), .Z(s[843]) );
  XOR2D0 C8374 ( .A1(p[844]), .A2(c[844]), .Z(s[844]) );
  XOR2D0 C8373 ( .A1(p[845]), .A2(c[845]), .Z(s[845]) );
  XOR2D0 C8372 ( .A1(p[846]), .A2(c[846]), .Z(s[846]) );
  XOR2D0 C8371 ( .A1(p[847]), .A2(c[847]), .Z(s[847]) );
  XOR2D0 C8370 ( .A1(p[848]), .A2(c[848]), .Z(s[848]) );
  XOR2D0 C8369 ( .A1(p[849]), .A2(c[849]), .Z(s[849]) );
  XOR2D0 C8368 ( .A1(p[850]), .A2(c[850]), .Z(s[850]) );
  XOR2D0 C8367 ( .A1(p[851]), .A2(c[851]), .Z(s[851]) );
  XOR2D0 C8366 ( .A1(p[852]), .A2(c[852]), .Z(s[852]) );
  XOR2D0 C8365 ( .A1(p[853]), .A2(c[853]), .Z(s[853]) );
  XOR2D0 C8364 ( .A1(p[854]), .A2(c[854]), .Z(s[854]) );
  XOR2D0 C8363 ( .A1(p[855]), .A2(c[855]), .Z(s[855]) );
  XOR2D0 C8362 ( .A1(p[856]), .A2(c[856]), .Z(s[856]) );
  XOR2D0 C8361 ( .A1(p[857]), .A2(c[857]), .Z(s[857]) );
  XOR2D0 C8360 ( .A1(p[858]), .A2(c[858]), .Z(s[858]) );
  XOR2D0 C8359 ( .A1(p[859]), .A2(c[859]), .Z(s[859]) );
  XOR2D0 C8358 ( .A1(p[860]), .A2(c[860]), .Z(s[860]) );
  XOR2D0 C8357 ( .A1(p[861]), .A2(c[861]), .Z(s[861]) );
  XOR2D0 C8356 ( .A1(p[862]), .A2(c[862]), .Z(s[862]) );
  XOR2D0 C8355 ( .A1(p[863]), .A2(c[863]), .Z(s[863]) );
  XOR2D0 C8354 ( .A1(p[864]), .A2(c[864]), .Z(s[864]) );
  XOR2D0 C8353 ( .A1(p[865]), .A2(c[865]), .Z(s[865]) );
  XOR2D0 C8352 ( .A1(p[866]), .A2(c[866]), .Z(s[866]) );
  XOR2D0 C8351 ( .A1(p[867]), .A2(c[867]), .Z(s[867]) );
  XOR2D0 C8350 ( .A1(p[868]), .A2(c[868]), .Z(s[868]) );
  XOR2D0 C8349 ( .A1(p[869]), .A2(c[869]), .Z(s[869]) );
  XOR2D0 C8348 ( .A1(p[870]), .A2(c[870]), .Z(s[870]) );
  XOR2D0 C8347 ( .A1(p[871]), .A2(c[871]), .Z(s[871]) );
  XOR2D0 C8346 ( .A1(p[872]), .A2(c[872]), .Z(s[872]) );
  XOR2D0 C8345 ( .A1(p[873]), .A2(c[873]), .Z(s[873]) );
  XOR2D0 C8344 ( .A1(p[874]), .A2(c[874]), .Z(s[874]) );
  XOR2D0 C8343 ( .A1(p[875]), .A2(c[875]), .Z(s[875]) );
  XOR2D0 C8342 ( .A1(p[876]), .A2(c[876]), .Z(s[876]) );
  XOR2D0 C8341 ( .A1(p[877]), .A2(c[877]), .Z(s[877]) );
  XOR2D0 C8340 ( .A1(p[878]), .A2(c[878]), .Z(s[878]) );
  XOR2D0 C8339 ( .A1(p[879]), .A2(c[879]), .Z(s[879]) );
  XOR2D0 C8338 ( .A1(p[880]), .A2(c[880]), .Z(s[880]) );
  XOR2D0 C8337 ( .A1(p[881]), .A2(c[881]), .Z(s[881]) );
  XOR2D0 C8336 ( .A1(p[882]), .A2(c[882]), .Z(s[882]) );
  XOR2D0 C8335 ( .A1(p[883]), .A2(c[883]), .Z(s[883]) );
  XOR2D0 C8334 ( .A1(p[884]), .A2(c[884]), .Z(s[884]) );
  XOR2D0 C8333 ( .A1(p[885]), .A2(c[885]), .Z(s[885]) );
  XOR2D0 C8332 ( .A1(p[886]), .A2(c[886]), .Z(s[886]) );
  XOR2D0 C8331 ( .A1(p[887]), .A2(c[887]), .Z(s[887]) );
  XOR2D0 C8330 ( .A1(p[888]), .A2(c[888]), .Z(s[888]) );
  XOR2D0 C8329 ( .A1(p[889]), .A2(c[889]), .Z(s[889]) );
  XOR2D0 C8328 ( .A1(p[890]), .A2(c[890]), .Z(s[890]) );
  XOR2D0 C8327 ( .A1(p[891]), .A2(c[891]), .Z(s[891]) );
  XOR2D0 C8326 ( .A1(p[892]), .A2(c[892]), .Z(s[892]) );
  XOR2D0 C8325 ( .A1(p[893]), .A2(c[893]), .Z(s[893]) );
  XOR2D0 C8324 ( .A1(p[894]), .A2(c[894]), .Z(s[894]) );
  XOR2D0 C8323 ( .A1(p[895]), .A2(c[895]), .Z(s[895]) );
  XOR2D0 C8322 ( .A1(p[896]), .A2(c[896]), .Z(s[896]) );
  XOR2D0 C8321 ( .A1(p[897]), .A2(c[897]), .Z(s[897]) );
  XOR2D0 C8320 ( .A1(p[898]), .A2(c[898]), .Z(s[898]) );
  XOR2D0 C8319 ( .A1(p[899]), .A2(c[899]), .Z(s[899]) );
  XOR2D0 C8318 ( .A1(p[900]), .A2(c[900]), .Z(s[900]) );
  XOR2D0 C8317 ( .A1(p[901]), .A2(c[901]), .Z(s[901]) );
  XOR2D0 C8316 ( .A1(p[902]), .A2(c[902]), .Z(s[902]) );
  XOR2D0 C8315 ( .A1(p[903]), .A2(c[903]), .Z(s[903]) );
  XOR2D0 C8314 ( .A1(p[904]), .A2(c[904]), .Z(s[904]) );
  XOR2D0 C8313 ( .A1(p[905]), .A2(c[905]), .Z(s[905]) );
  XOR2D0 C8312 ( .A1(p[906]), .A2(c[906]), .Z(s[906]) );
  XOR2D0 C8311 ( .A1(p[907]), .A2(c[907]), .Z(s[907]) );
  XOR2D0 C8310 ( .A1(p[908]), .A2(c[908]), .Z(s[908]) );
  XOR2D0 C8309 ( .A1(p[909]), .A2(c[909]), .Z(s[909]) );
  XOR2D0 C8308 ( .A1(p[910]), .A2(c[910]), .Z(s[910]) );
  XOR2D0 C8307 ( .A1(p[911]), .A2(c[911]), .Z(s[911]) );
  XOR2D0 C8306 ( .A1(p[912]), .A2(c[912]), .Z(s[912]) );
  XOR2D0 C8305 ( .A1(p[913]), .A2(c[913]), .Z(s[913]) );
  XOR2D0 C8304 ( .A1(p[914]), .A2(c[914]), .Z(s[914]) );
  XOR2D0 C8303 ( .A1(p[915]), .A2(c[915]), .Z(s[915]) );
  XOR2D0 C8302 ( .A1(p[916]), .A2(c[916]), .Z(s[916]) );
  XOR2D0 C8301 ( .A1(p[917]), .A2(c[917]), .Z(s[917]) );
  XOR2D0 C8300 ( .A1(p[918]), .A2(c[918]), .Z(s[918]) );
  XOR2D0 C8299 ( .A1(p[919]), .A2(c[919]), .Z(s[919]) );
  XOR2D0 C8298 ( .A1(p[920]), .A2(c[920]), .Z(s[920]) );
  XOR2D0 C8297 ( .A1(p[921]), .A2(c[921]), .Z(s[921]) );
  XOR2D0 C8296 ( .A1(p[922]), .A2(c[922]), .Z(s[922]) );
  XOR2D0 C8295 ( .A1(p[923]), .A2(c[923]), .Z(s[923]) );
  XOR2D0 C8294 ( .A1(p[924]), .A2(c[924]), .Z(s[924]) );
  XOR2D0 C8293 ( .A1(p[925]), .A2(c[925]), .Z(s[925]) );
  XOR2D0 C8292 ( .A1(p[926]), .A2(c[926]), .Z(s[926]) );
  XOR2D0 C8291 ( .A1(p[927]), .A2(c[927]), .Z(s[927]) );
  XOR2D0 C8290 ( .A1(p[928]), .A2(c[928]), .Z(s[928]) );
  XOR2D0 C8289 ( .A1(p[929]), .A2(c[929]), .Z(s[929]) );
  XOR2D0 C8288 ( .A1(p[930]), .A2(c[930]), .Z(s[930]) );
  XOR2D0 C8287 ( .A1(p[931]), .A2(c[931]), .Z(s[931]) );
  XOR2D0 C8286 ( .A1(p[932]), .A2(c[932]), .Z(s[932]) );
  XOR2D0 C8285 ( .A1(p[933]), .A2(c[933]), .Z(s[933]) );
  XOR2D0 C8284 ( .A1(p[934]), .A2(c[934]), .Z(s[934]) );
  XOR2D0 C8283 ( .A1(p[935]), .A2(c[935]), .Z(s[935]) );
  XOR2D0 C8282 ( .A1(p[936]), .A2(c[936]), .Z(s[936]) );
  XOR2D0 C8281 ( .A1(p[937]), .A2(c[937]), .Z(s[937]) );
  XOR2D0 C8280 ( .A1(p[938]), .A2(c[938]), .Z(s[938]) );
  XOR2D0 C8279 ( .A1(p[939]), .A2(c[939]), .Z(s[939]) );
  XOR2D0 C8278 ( .A1(p[940]), .A2(c[940]), .Z(s[940]) );
  XOR2D0 C8277 ( .A1(p[941]), .A2(c[941]), .Z(s[941]) );
  XOR2D0 C8276 ( .A1(p[942]), .A2(c[942]), .Z(s[942]) );
  XOR2D0 C8275 ( .A1(p[943]), .A2(c[943]), .Z(s[943]) );
  XOR2D0 C8274 ( .A1(p[944]), .A2(c[944]), .Z(s[944]) );
  XOR2D0 C8273 ( .A1(p[945]), .A2(c[945]), .Z(s[945]) );
  XOR2D0 C8272 ( .A1(p[946]), .A2(c[946]), .Z(s[946]) );
  XOR2D0 C8271 ( .A1(p[947]), .A2(c[947]), .Z(s[947]) );
  XOR2D0 C8270 ( .A1(p[948]), .A2(c[948]), .Z(s[948]) );
  XOR2D0 C8269 ( .A1(p[949]), .A2(c[949]), .Z(s[949]) );
  XOR2D0 C8268 ( .A1(p[950]), .A2(c[950]), .Z(s[950]) );
  XOR2D0 C8267 ( .A1(p[951]), .A2(c[951]), .Z(s[951]) );
  XOR2D0 C8266 ( .A1(p[952]), .A2(c[952]), .Z(s[952]) );
  XOR2D0 C8265 ( .A1(p[953]), .A2(c[953]), .Z(s[953]) );
  XOR2D0 C8264 ( .A1(p[954]), .A2(c[954]), .Z(s[954]) );
  XOR2D0 C8263 ( .A1(p[955]), .A2(c[955]), .Z(s[955]) );
  XOR2D0 C8262 ( .A1(p[956]), .A2(c[956]), .Z(s[956]) );
  XOR2D0 C8261 ( .A1(p[957]), .A2(c[957]), .Z(s[957]) );
  XOR2D0 C8260 ( .A1(p[958]), .A2(c[958]), .Z(s[958]) );
  XOR2D0 C8259 ( .A1(p[959]), .A2(c[959]), .Z(s[959]) );
  XOR2D0 C8258 ( .A1(p[960]), .A2(c[960]), .Z(s[960]) );
  XOR2D0 C8257 ( .A1(p[961]), .A2(c[961]), .Z(s[961]) );
  XOR2D0 C8256 ( .A1(p[962]), .A2(c[962]), .Z(s[962]) );
  XOR2D0 C8255 ( .A1(p[963]), .A2(c[963]), .Z(s[963]) );
  XOR2D0 C8254 ( .A1(p[964]), .A2(c[964]), .Z(s[964]) );
  XOR2D0 C8253 ( .A1(p[965]), .A2(c[965]), .Z(s[965]) );
  XOR2D0 C8252 ( .A1(p[966]), .A2(c[966]), .Z(s[966]) );
  XOR2D0 C8251 ( .A1(p[967]), .A2(c[967]), .Z(s[967]) );
  XOR2D0 C8250 ( .A1(p[968]), .A2(c[968]), .Z(s[968]) );
  XOR2D0 C8249 ( .A1(p[969]), .A2(c[969]), .Z(s[969]) );
  XOR2D0 C8248 ( .A1(p[970]), .A2(c[970]), .Z(s[970]) );
  XOR2D0 C8247 ( .A1(p[971]), .A2(c[971]), .Z(s[971]) );
  XOR2D0 C8246 ( .A1(p[972]), .A2(c[972]), .Z(s[972]) );
  XOR2D0 C8245 ( .A1(p[973]), .A2(c[973]), .Z(s[973]) );
  XOR2D0 C8244 ( .A1(p[974]), .A2(c[974]), .Z(s[974]) );
  XOR2D0 C8243 ( .A1(p[975]), .A2(c[975]), .Z(s[975]) );
  XOR2D0 C8242 ( .A1(p[976]), .A2(c[976]), .Z(s[976]) );
  XOR2D0 C8241 ( .A1(p[977]), .A2(c[977]), .Z(s[977]) );
  XOR2D0 C8240 ( .A1(p[978]), .A2(c[978]), .Z(s[978]) );
  XOR2D0 C8239 ( .A1(p[979]), .A2(c[979]), .Z(s[979]) );
  XOR2D0 C8238 ( .A1(p[980]), .A2(c[980]), .Z(s[980]) );
  XOR2D0 C8237 ( .A1(p[981]), .A2(c[981]), .Z(s[981]) );
  XOR2D0 C8236 ( .A1(p[982]), .A2(c[982]), .Z(s[982]) );
  XOR2D0 C8235 ( .A1(p[983]), .A2(c[983]), .Z(s[983]) );
  XOR2D0 C8234 ( .A1(p[984]), .A2(c[984]), .Z(s[984]) );
  XOR2D0 C8233 ( .A1(p[985]), .A2(c[985]), .Z(s[985]) );
  XOR2D0 C8232 ( .A1(p[986]), .A2(c[986]), .Z(s[986]) );
  XOR2D0 C8231 ( .A1(p[987]), .A2(c[987]), .Z(s[987]) );
  XOR2D0 C8230 ( .A1(p[988]), .A2(c[988]), .Z(s[988]) );
  XOR2D0 C8229 ( .A1(p[989]), .A2(c[989]), .Z(s[989]) );
  XOR2D0 C8228 ( .A1(p[990]), .A2(c[990]), .Z(s[990]) );
  XOR2D0 C8227 ( .A1(p[991]), .A2(c[991]), .Z(s[991]) );
  XOR2D0 C8226 ( .A1(p[992]), .A2(c[992]), .Z(s[992]) );
  XOR2D0 C8225 ( .A1(p[993]), .A2(c[993]), .Z(s[993]) );
  XOR2D0 C8224 ( .A1(p[994]), .A2(c[994]), .Z(s[994]) );
  XOR2D0 C8223 ( .A1(p[995]), .A2(c[995]), .Z(s[995]) );
  XOR2D0 C8222 ( .A1(p[996]), .A2(c[996]), .Z(s[996]) );
  XOR2D0 C8221 ( .A1(p[997]), .A2(c[997]), .Z(s[997]) );
  XOR2D0 C8220 ( .A1(p[998]), .A2(c[998]), .Z(s[998]) );
  XOR2D0 C8219 ( .A1(p[999]), .A2(c[999]), .Z(s[999]) );
  XOR2D0 C8218 ( .A1(p[1000]), .A2(c[1000]), .Z(s[1000]) );
  XOR2D0 C8217 ( .A1(p[1001]), .A2(c[1001]), .Z(s[1001]) );
  XOR2D0 C8216 ( .A1(p[1002]), .A2(c[1002]), .Z(s[1002]) );
  XOR2D0 C8215 ( .A1(p[1003]), .A2(c[1003]), .Z(s[1003]) );
  XOR2D0 C8214 ( .A1(p[1004]), .A2(c[1004]), .Z(s[1004]) );
  XOR2D0 C8213 ( .A1(p[1005]), .A2(c[1005]), .Z(s[1005]) );
  XOR2D0 C8212 ( .A1(p[1006]), .A2(c[1006]), .Z(s[1006]) );
  XOR2D0 C8211 ( .A1(p[1007]), .A2(c[1007]), .Z(s[1007]) );
  XOR2D0 C8210 ( .A1(p[1008]), .A2(c[1008]), .Z(s[1008]) );
  XOR2D0 C8209 ( .A1(p[1009]), .A2(c[1009]), .Z(s[1009]) );
  XOR2D0 C8208 ( .A1(p[1010]), .A2(c[1010]), .Z(s[1010]) );
  XOR2D0 C8207 ( .A1(p[1011]), .A2(c[1011]), .Z(s[1011]) );
  XOR2D0 C8206 ( .A1(p[1012]), .A2(c[1012]), .Z(s[1012]) );
  XOR2D0 C8205 ( .A1(p[1013]), .A2(c[1013]), .Z(s[1013]) );
  XOR2D0 C8204 ( .A1(p[1014]), .A2(c[1014]), .Z(s[1014]) );
  XOR2D0 C8203 ( .A1(p[1015]), .A2(c[1015]), .Z(s[1015]) );
  XOR2D0 C8202 ( .A1(p[1016]), .A2(c[1016]), .Z(s[1016]) );
  XOR2D0 C8201 ( .A1(p[1017]), .A2(c[1017]), .Z(s[1017]) );
  XOR2D0 C8200 ( .A1(p[1018]), .A2(c[1018]), .Z(s[1018]) );
  XOR2D0 C8199 ( .A1(p[1019]), .A2(c[1019]), .Z(s[1019]) );
  XOR2D0 C8198 ( .A1(p[1020]), .A2(c[1020]), .Z(s[1020]) );
  XOR2D0 C8197 ( .A1(p[1021]), .A2(c[1021]), .Z(s[1021]) );
  XOR2D0 C8196 ( .A1(p[1022]), .A2(c[1022]), .Z(s[1022]) );
  XOR2D0 C8195 ( .A1(p[1023]), .A2(c[1023]), .Z(s[1023]) );
  AN2D0 C8194 ( .A1(p[1022]), .A2(c[1022]), .Z(N1022) );
  OR2D0 C8193 ( .A1(g[1022]), .A2(N1022), .Z(c[1023]) );
  AN2D0 C8192 ( .A1(p[1021]), .A2(c[1021]), .Z(N1021) );
  OR2D0 C8191 ( .A1(g[1021]), .A2(N1021), .Z(c[1022]) );
  AN2D0 C8190 ( .A1(p[1020]), .A2(c[1020]), .Z(N1020) );
  OR2D0 C8189 ( .A1(g[1020]), .A2(N1020), .Z(c[1021]) );
  AN2D0 C8188 ( .A1(p[1019]), .A2(c[1019]), .Z(N1019) );
  OR2D0 C8187 ( .A1(g[1019]), .A2(N1019), .Z(c[1020]) );
  AN2D0 C8186 ( .A1(p[1018]), .A2(c[1018]), .Z(N1018) );
  OR2D0 C8185 ( .A1(g[1018]), .A2(N1018), .Z(c[1019]) );
  AN2D0 C8184 ( .A1(p[1017]), .A2(c[1017]), .Z(N1017) );
  OR2D0 C8183 ( .A1(g[1017]), .A2(N1017), .Z(c[1018]) );
  AN2D0 C8182 ( .A1(p[1016]), .A2(c[1016]), .Z(N1016) );
  OR2D0 C8181 ( .A1(g[1016]), .A2(N1016), .Z(c[1017]) );
  AN2D0 C8180 ( .A1(p[1015]), .A2(c[1015]), .Z(N1015) );
  OR2D0 C8179 ( .A1(g[1015]), .A2(N1015), .Z(c[1016]) );
  AN2D0 C8178 ( .A1(p[1014]), .A2(c[1014]), .Z(N1014) );
  OR2D0 C8177 ( .A1(g[1014]), .A2(N1014), .Z(c[1015]) );
  AN2D0 C8176 ( .A1(p[1013]), .A2(c[1013]), .Z(N1013) );
  OR2D0 C8175 ( .A1(g[1013]), .A2(N1013), .Z(c[1014]) );
  AN2D0 C8174 ( .A1(p[1012]), .A2(c[1012]), .Z(N1012) );
  OR2D0 C8173 ( .A1(g[1012]), .A2(N1012), .Z(c[1013]) );
  AN2D0 C8172 ( .A1(p[1011]), .A2(c[1011]), .Z(N1011) );
  OR2D0 C8171 ( .A1(g[1011]), .A2(N1011), .Z(c[1012]) );
  AN2D0 C8170 ( .A1(p[1010]), .A2(c[1010]), .Z(N1010) );
  OR2D0 C8169 ( .A1(g[1010]), .A2(N1010), .Z(c[1011]) );
  AN2D0 C8168 ( .A1(p[1009]), .A2(c[1009]), .Z(N1009) );
  OR2D0 C8167 ( .A1(g[1009]), .A2(N1009), .Z(c[1010]) );
  AN2D0 C8166 ( .A1(p[1008]), .A2(c[1008]), .Z(N1008) );
  OR2D0 C8165 ( .A1(g[1008]), .A2(N1008), .Z(c[1009]) );
  AN2D0 C8164 ( .A1(p[1007]), .A2(c[1007]), .Z(N1007) );
  OR2D0 C8163 ( .A1(g[1007]), .A2(N1007), .Z(c[1008]) );
  AN2D0 C8162 ( .A1(p[1006]), .A2(c[1006]), .Z(N1006) );
  OR2D0 C8161 ( .A1(g[1006]), .A2(N1006), .Z(c[1007]) );
  AN2D0 C8160 ( .A1(p[1005]), .A2(c[1005]), .Z(N1005) );
  OR2D0 C8159 ( .A1(g[1005]), .A2(N1005), .Z(c[1006]) );
  AN2D0 C8158 ( .A1(p[1004]), .A2(c[1004]), .Z(N1004) );
  OR2D0 C8157 ( .A1(g[1004]), .A2(N1004), .Z(c[1005]) );
  AN2D0 C8156 ( .A1(p[1003]), .A2(c[1003]), .Z(N1003) );
  OR2D0 C8155 ( .A1(g[1003]), .A2(N1003), .Z(c[1004]) );
  AN2D0 C8154 ( .A1(p[1002]), .A2(c[1002]), .Z(N1002) );
  OR2D0 C8153 ( .A1(g[1002]), .A2(N1002), .Z(c[1003]) );
  AN2D0 C8152 ( .A1(p[1001]), .A2(c[1001]), .Z(N1001) );
  OR2D0 C8151 ( .A1(g[1001]), .A2(N1001), .Z(c[1002]) );
  AN2D0 C8150 ( .A1(p[1000]), .A2(c[1000]), .Z(N1000) );
  OR2D0 C8149 ( .A1(g[1000]), .A2(N1000), .Z(c[1001]) );
  AN2D0 C8148 ( .A1(p[999]), .A2(c[999]), .Z(N999) );
  OR2D0 C8147 ( .A1(g[999]), .A2(N999), .Z(c[1000]) );
  AN2D0 C8146 ( .A1(p[998]), .A2(c[998]), .Z(N998) );
  OR2D0 C8145 ( .A1(g[998]), .A2(N998), .Z(c[999]) );
  AN2D0 C8144 ( .A1(p[997]), .A2(c[997]), .Z(N997) );
  OR2D0 C8143 ( .A1(g[997]), .A2(N997), .Z(c[998]) );
  AN2D0 C8142 ( .A1(p[996]), .A2(c[996]), .Z(N996) );
  OR2D0 C8141 ( .A1(g[996]), .A2(N996), .Z(c[997]) );
  AN2D0 C8140 ( .A1(p[995]), .A2(c[995]), .Z(N995) );
  OR2D0 C8139 ( .A1(g[995]), .A2(N995), .Z(c[996]) );
  AN2D0 C8138 ( .A1(p[994]), .A2(c[994]), .Z(N994) );
  OR2D0 C8137 ( .A1(g[994]), .A2(N994), .Z(c[995]) );
  AN2D0 C8136 ( .A1(p[993]), .A2(c[993]), .Z(N993) );
  OR2D0 C8135 ( .A1(g[993]), .A2(N993), .Z(c[994]) );
  AN2D0 C8134 ( .A1(p[992]), .A2(c[992]), .Z(N992) );
  OR2D0 C8133 ( .A1(g[992]), .A2(N992), .Z(c[993]) );
  AN2D0 C8132 ( .A1(p[991]), .A2(c[991]), .Z(N991) );
  OR2D0 C8131 ( .A1(g[991]), .A2(N991), .Z(c[992]) );
  AN2D0 C8130 ( .A1(p[990]), .A2(c[990]), .Z(N990) );
  OR2D0 C8129 ( .A1(g[990]), .A2(N990), .Z(c[991]) );
  AN2D0 C8128 ( .A1(p[989]), .A2(c[989]), .Z(N989) );
  OR2D0 C8127 ( .A1(g[989]), .A2(N989), .Z(c[990]) );
  AN2D0 C8126 ( .A1(p[988]), .A2(c[988]), .Z(N988) );
  OR2D0 C8125 ( .A1(g[988]), .A2(N988), .Z(c[989]) );
  AN2D0 C8124 ( .A1(p[987]), .A2(c[987]), .Z(N987) );
  OR2D0 C8123 ( .A1(g[987]), .A2(N987), .Z(c[988]) );
  AN2D0 C8122 ( .A1(p[986]), .A2(c[986]), .Z(N986) );
  OR2D0 C8121 ( .A1(g[986]), .A2(N986), .Z(c[987]) );
  AN2D0 C8120 ( .A1(p[985]), .A2(c[985]), .Z(N985) );
  OR2D0 C8119 ( .A1(g[985]), .A2(N985), .Z(c[986]) );
  AN2D0 C8118 ( .A1(p[984]), .A2(c[984]), .Z(N984) );
  OR2D0 C8117 ( .A1(g[984]), .A2(N984), .Z(c[985]) );
  AN2D0 C8116 ( .A1(p[983]), .A2(c[983]), .Z(N983) );
  OR2D0 C8115 ( .A1(g[983]), .A2(N983), .Z(c[984]) );
  AN2D0 C8114 ( .A1(p[982]), .A2(c[982]), .Z(N982) );
  OR2D0 C8113 ( .A1(g[982]), .A2(N982), .Z(c[983]) );
  AN2D0 C8112 ( .A1(p[981]), .A2(c[981]), .Z(N981) );
  OR2D0 C8111 ( .A1(g[981]), .A2(N981), .Z(c[982]) );
  AN2D0 C8110 ( .A1(p[980]), .A2(c[980]), .Z(N980) );
  OR2D0 C8109 ( .A1(g[980]), .A2(N980), .Z(c[981]) );
  AN2D0 C8108 ( .A1(p[979]), .A2(c[979]), .Z(N979) );
  OR2D0 C8107 ( .A1(g[979]), .A2(N979), .Z(c[980]) );
  AN2D0 C8106 ( .A1(p[978]), .A2(c[978]), .Z(N978) );
  OR2D0 C8105 ( .A1(g[978]), .A2(N978), .Z(c[979]) );
  AN2D0 C8104 ( .A1(p[977]), .A2(c[977]), .Z(N977) );
  OR2D0 C8103 ( .A1(g[977]), .A2(N977), .Z(c[978]) );
  AN2D0 C8102 ( .A1(p[976]), .A2(c[976]), .Z(N976) );
  OR2D0 C8101 ( .A1(g[976]), .A2(N976), .Z(c[977]) );
  AN2D0 C8100 ( .A1(p[975]), .A2(c[975]), .Z(N975) );
  OR2D0 C8099 ( .A1(g[975]), .A2(N975), .Z(c[976]) );
  AN2D0 C8098 ( .A1(p[974]), .A2(c[974]), .Z(N974) );
  OR2D0 C8097 ( .A1(g[974]), .A2(N974), .Z(c[975]) );
  AN2D0 C8096 ( .A1(p[973]), .A2(c[973]), .Z(N973) );
  OR2D0 C8095 ( .A1(g[973]), .A2(N973), .Z(c[974]) );
  AN2D0 C8094 ( .A1(p[972]), .A2(c[972]), .Z(N972) );
  OR2D0 C8093 ( .A1(g[972]), .A2(N972), .Z(c[973]) );
  AN2D0 C8092 ( .A1(p[971]), .A2(c[971]), .Z(N971) );
  OR2D0 C8091 ( .A1(g[971]), .A2(N971), .Z(c[972]) );
  AN2D0 C8090 ( .A1(p[970]), .A2(c[970]), .Z(N970) );
  OR2D0 C8089 ( .A1(g[970]), .A2(N970), .Z(c[971]) );
  AN2D0 C8088 ( .A1(p[969]), .A2(c[969]), .Z(N969) );
  OR2D0 C8087 ( .A1(g[969]), .A2(N969), .Z(c[970]) );
  AN2D0 C8086 ( .A1(p[968]), .A2(c[968]), .Z(N968) );
  OR2D0 C8085 ( .A1(g[968]), .A2(N968), .Z(c[969]) );
  AN2D0 C8084 ( .A1(p[967]), .A2(c[967]), .Z(N967) );
  OR2D0 C8083 ( .A1(g[967]), .A2(N967), .Z(c[968]) );
  AN2D0 C8082 ( .A1(p[966]), .A2(c[966]), .Z(N966) );
  OR2D0 C8081 ( .A1(g[966]), .A2(N966), .Z(c[967]) );
  AN2D0 C8080 ( .A1(p[965]), .A2(c[965]), .Z(N965) );
  OR2D0 C8079 ( .A1(g[965]), .A2(N965), .Z(c[966]) );
  AN2D0 C8078 ( .A1(p[964]), .A2(c[964]), .Z(N964) );
  OR2D0 C8077 ( .A1(g[964]), .A2(N964), .Z(c[965]) );
  AN2D0 C8076 ( .A1(p[963]), .A2(c[963]), .Z(N963) );
  OR2D0 C8075 ( .A1(g[963]), .A2(N963), .Z(c[964]) );
  AN2D0 C8074 ( .A1(p[962]), .A2(c[962]), .Z(N962) );
  OR2D0 C8073 ( .A1(g[962]), .A2(N962), .Z(c[963]) );
  AN2D0 C8072 ( .A1(p[961]), .A2(c[961]), .Z(N961) );
  OR2D0 C8071 ( .A1(g[961]), .A2(N961), .Z(c[962]) );
  AN2D0 C8070 ( .A1(p[960]), .A2(c[960]), .Z(N960) );
  OR2D0 C8069 ( .A1(g[960]), .A2(N960), .Z(c[961]) );
  AN2D0 C8068 ( .A1(p[959]), .A2(c[959]), .Z(N959) );
  OR2D0 C8067 ( .A1(g[959]), .A2(N959), .Z(c[960]) );
  AN2D0 C8066 ( .A1(p[958]), .A2(c[958]), .Z(N958) );
  OR2D0 C8065 ( .A1(g[958]), .A2(N958), .Z(c[959]) );
  AN2D0 C8064 ( .A1(p[957]), .A2(c[957]), .Z(N957) );
  OR2D0 C8063 ( .A1(g[957]), .A2(N957), .Z(c[958]) );
  AN2D0 C8062 ( .A1(p[956]), .A2(c[956]), .Z(N956) );
  OR2D0 C8061 ( .A1(g[956]), .A2(N956), .Z(c[957]) );
  AN2D0 C8060 ( .A1(p[955]), .A2(c[955]), .Z(N955) );
  OR2D0 C8059 ( .A1(g[955]), .A2(N955), .Z(c[956]) );
  AN2D0 C8058 ( .A1(p[954]), .A2(c[954]), .Z(N954) );
  OR2D0 C8057 ( .A1(g[954]), .A2(N954), .Z(c[955]) );
  AN2D0 C8056 ( .A1(p[953]), .A2(c[953]), .Z(N953) );
  OR2D0 C8055 ( .A1(g[953]), .A2(N953), .Z(c[954]) );
  AN2D0 C8054 ( .A1(p[952]), .A2(c[952]), .Z(N952) );
  OR2D0 C8053 ( .A1(g[952]), .A2(N952), .Z(c[953]) );
  AN2D0 C8052 ( .A1(p[951]), .A2(c[951]), .Z(N951) );
  OR2D0 C8051 ( .A1(g[951]), .A2(N951), .Z(c[952]) );
  AN2D0 C8050 ( .A1(p[950]), .A2(c[950]), .Z(N950) );
  OR2D0 C8049 ( .A1(g[950]), .A2(N950), .Z(c[951]) );
  AN2D0 C8048 ( .A1(p[949]), .A2(c[949]), .Z(N949) );
  OR2D0 C8047 ( .A1(g[949]), .A2(N949), .Z(c[950]) );
  AN2D0 C8046 ( .A1(p[948]), .A2(c[948]), .Z(N948) );
  OR2D0 C8045 ( .A1(g[948]), .A2(N948), .Z(c[949]) );
  AN2D0 C8044 ( .A1(p[947]), .A2(c[947]), .Z(N947) );
  OR2D0 C8043 ( .A1(g[947]), .A2(N947), .Z(c[948]) );
  AN2D0 C8042 ( .A1(p[946]), .A2(c[946]), .Z(N946) );
  OR2D0 C8041 ( .A1(g[946]), .A2(N946), .Z(c[947]) );
  AN2D0 C8040 ( .A1(p[945]), .A2(c[945]), .Z(N945) );
  OR2D0 C8039 ( .A1(g[945]), .A2(N945), .Z(c[946]) );
  AN2D0 C8038 ( .A1(p[944]), .A2(c[944]), .Z(N944) );
  OR2D0 C8037 ( .A1(g[944]), .A2(N944), .Z(c[945]) );
  AN2D0 C8036 ( .A1(p[943]), .A2(c[943]), .Z(N943) );
  OR2D0 C8035 ( .A1(g[943]), .A2(N943), .Z(c[944]) );
  AN2D0 C8034 ( .A1(p[942]), .A2(c[942]), .Z(N942) );
  OR2D0 C8033 ( .A1(g[942]), .A2(N942), .Z(c[943]) );
  AN2D0 C8032 ( .A1(p[941]), .A2(c[941]), .Z(N941) );
  OR2D0 C8031 ( .A1(g[941]), .A2(N941), .Z(c[942]) );
  AN2D0 C8030 ( .A1(p[940]), .A2(c[940]), .Z(N940) );
  OR2D0 C8029 ( .A1(g[940]), .A2(N940), .Z(c[941]) );
  AN2D0 C8028 ( .A1(p[939]), .A2(c[939]), .Z(N939) );
  OR2D0 C8027 ( .A1(g[939]), .A2(N939), .Z(c[940]) );
  AN2D0 C8026 ( .A1(p[938]), .A2(c[938]), .Z(N938) );
  OR2D0 C8025 ( .A1(g[938]), .A2(N938), .Z(c[939]) );
  AN2D0 C8024 ( .A1(p[937]), .A2(c[937]), .Z(N937) );
  OR2D0 C8023 ( .A1(g[937]), .A2(N937), .Z(c[938]) );
  AN2D0 C8022 ( .A1(p[936]), .A2(c[936]), .Z(N936) );
  OR2D0 C8021 ( .A1(g[936]), .A2(N936), .Z(c[937]) );
  AN2D0 C8020 ( .A1(p[935]), .A2(c[935]), .Z(N935) );
  OR2D0 C8019 ( .A1(g[935]), .A2(N935), .Z(c[936]) );
  AN2D0 C8018 ( .A1(p[934]), .A2(c[934]), .Z(N934) );
  OR2D0 C8017 ( .A1(g[934]), .A2(N934), .Z(c[935]) );
  AN2D0 C8016 ( .A1(p[933]), .A2(c[933]), .Z(N933) );
  OR2D0 C8015 ( .A1(g[933]), .A2(N933), .Z(c[934]) );
  AN2D0 C8014 ( .A1(p[932]), .A2(c[932]), .Z(N932) );
  OR2D0 C8013 ( .A1(g[932]), .A2(N932), .Z(c[933]) );
  AN2D0 C8012 ( .A1(p[931]), .A2(c[931]), .Z(N931) );
  OR2D0 C8011 ( .A1(g[931]), .A2(N931), .Z(c[932]) );
  AN2D0 C8010 ( .A1(p[930]), .A2(c[930]), .Z(N930) );
  OR2D0 C8009 ( .A1(g[930]), .A2(N930), .Z(c[931]) );
  AN2D0 C8008 ( .A1(p[929]), .A2(c[929]), .Z(N929) );
  OR2D0 C8007 ( .A1(g[929]), .A2(N929), .Z(c[930]) );
  AN2D0 C8006 ( .A1(p[928]), .A2(c[928]), .Z(N928) );
  OR2D0 C8005 ( .A1(g[928]), .A2(N928), .Z(c[929]) );
  AN2D0 C8004 ( .A1(p[927]), .A2(c[927]), .Z(N927) );
  OR2D0 C8003 ( .A1(g[927]), .A2(N927), .Z(c[928]) );
  AN2D0 C8002 ( .A1(p[926]), .A2(c[926]), .Z(N926) );
  OR2D0 C8001 ( .A1(g[926]), .A2(N926), .Z(c[927]) );
  AN2D0 C8000 ( .A1(p[925]), .A2(c[925]), .Z(N925) );
  OR2D0 C7999 ( .A1(g[925]), .A2(N925), .Z(c[926]) );
  AN2D0 C7998 ( .A1(p[924]), .A2(c[924]), .Z(N924) );
  OR2D0 C7997 ( .A1(g[924]), .A2(N924), .Z(c[925]) );
  AN2D0 C7996 ( .A1(p[923]), .A2(c[923]), .Z(N923) );
  OR2D0 C7995 ( .A1(g[923]), .A2(N923), .Z(c[924]) );
  AN2D0 C7994 ( .A1(p[922]), .A2(c[922]), .Z(N922) );
  OR2D0 C7993 ( .A1(g[922]), .A2(N922), .Z(c[923]) );
  AN2D0 C7992 ( .A1(p[921]), .A2(c[921]), .Z(N921) );
  OR2D0 C7991 ( .A1(g[921]), .A2(N921), .Z(c[922]) );
  AN2D0 C7990 ( .A1(p[920]), .A2(c[920]), .Z(N920) );
  OR2D0 C7989 ( .A1(g[920]), .A2(N920), .Z(c[921]) );
  AN2D0 C7988 ( .A1(p[919]), .A2(c[919]), .Z(N919) );
  OR2D0 C7987 ( .A1(g[919]), .A2(N919), .Z(c[920]) );
  AN2D0 C7986 ( .A1(p[918]), .A2(c[918]), .Z(N918) );
  OR2D0 C7985 ( .A1(g[918]), .A2(N918), .Z(c[919]) );
  AN2D0 C7984 ( .A1(p[917]), .A2(c[917]), .Z(N917) );
  OR2D0 C7983 ( .A1(g[917]), .A2(N917), .Z(c[918]) );
  AN2D0 C7982 ( .A1(p[916]), .A2(c[916]), .Z(N916) );
  OR2D0 C7981 ( .A1(g[916]), .A2(N916), .Z(c[917]) );
  AN2D0 C7980 ( .A1(p[915]), .A2(c[915]), .Z(N915) );
  OR2D0 C7979 ( .A1(g[915]), .A2(N915), .Z(c[916]) );
  AN2D0 C7978 ( .A1(p[914]), .A2(c[914]), .Z(N914) );
  OR2D0 C7977 ( .A1(g[914]), .A2(N914), .Z(c[915]) );
  AN2D0 C7976 ( .A1(p[913]), .A2(c[913]), .Z(N913) );
  OR2D0 C7975 ( .A1(g[913]), .A2(N913), .Z(c[914]) );
  AN2D0 C7974 ( .A1(p[912]), .A2(c[912]), .Z(N912) );
  OR2D0 C7973 ( .A1(g[912]), .A2(N912), .Z(c[913]) );
  AN2D0 C7972 ( .A1(p[911]), .A2(c[911]), .Z(N911) );
  OR2D0 C7971 ( .A1(g[911]), .A2(N911), .Z(c[912]) );
  AN2D0 C7970 ( .A1(p[910]), .A2(c[910]), .Z(N910) );
  OR2D0 C7969 ( .A1(g[910]), .A2(N910), .Z(c[911]) );
  AN2D0 C7968 ( .A1(p[909]), .A2(c[909]), .Z(N909) );
  OR2D0 C7967 ( .A1(g[909]), .A2(N909), .Z(c[910]) );
  AN2D0 C7966 ( .A1(p[908]), .A2(c[908]), .Z(N908) );
  OR2D0 C7965 ( .A1(g[908]), .A2(N908), .Z(c[909]) );
  AN2D0 C7964 ( .A1(p[907]), .A2(c[907]), .Z(N907) );
  OR2D0 C7963 ( .A1(g[907]), .A2(N907), .Z(c[908]) );
  AN2D0 C7962 ( .A1(p[906]), .A2(c[906]), .Z(N906) );
  OR2D0 C7961 ( .A1(g[906]), .A2(N906), .Z(c[907]) );
  AN2D0 C7960 ( .A1(p[905]), .A2(c[905]), .Z(N905) );
  OR2D0 C7959 ( .A1(g[905]), .A2(N905), .Z(c[906]) );
  AN2D0 C7958 ( .A1(p[904]), .A2(c[904]), .Z(N904) );
  OR2D0 C7957 ( .A1(g[904]), .A2(N904), .Z(c[905]) );
  AN2D0 C7956 ( .A1(p[903]), .A2(c[903]), .Z(N903) );
  OR2D0 C7955 ( .A1(g[903]), .A2(N903), .Z(c[904]) );
  AN2D0 C7954 ( .A1(p[902]), .A2(c[902]), .Z(N902) );
  OR2D0 C7953 ( .A1(g[902]), .A2(N902), .Z(c[903]) );
  AN2D0 C7952 ( .A1(p[901]), .A2(c[901]), .Z(N901) );
  OR2D0 C7951 ( .A1(g[901]), .A2(N901), .Z(c[902]) );
  AN2D0 C7950 ( .A1(p[900]), .A2(c[900]), .Z(N900) );
  OR2D0 C7949 ( .A1(g[900]), .A2(N900), .Z(c[901]) );
  AN2D0 C7948 ( .A1(p[899]), .A2(c[899]), .Z(N899) );
  OR2D0 C7947 ( .A1(g[899]), .A2(N899), .Z(c[900]) );
  AN2D0 C7946 ( .A1(p[898]), .A2(c[898]), .Z(N898) );
  OR2D0 C7945 ( .A1(g[898]), .A2(N898), .Z(c[899]) );
  AN2D0 C7944 ( .A1(p[897]), .A2(c[897]), .Z(N897) );
  OR2D0 C7943 ( .A1(g[897]), .A2(N897), .Z(c[898]) );
  AN2D0 C7942 ( .A1(p[896]), .A2(c[896]), .Z(N896) );
  OR2D0 C7941 ( .A1(g[896]), .A2(N896), .Z(c[897]) );
  AN2D0 C7940 ( .A1(p[895]), .A2(c[895]), .Z(N895) );
  OR2D0 C7939 ( .A1(g[895]), .A2(N895), .Z(c[896]) );
  AN2D0 C7938 ( .A1(p[894]), .A2(c[894]), .Z(N894) );
  OR2D0 C7937 ( .A1(g[894]), .A2(N894), .Z(c[895]) );
  AN2D0 C7936 ( .A1(p[893]), .A2(c[893]), .Z(N893) );
  OR2D0 C7935 ( .A1(g[893]), .A2(N893), .Z(c[894]) );
  AN2D0 C7934 ( .A1(p[892]), .A2(c[892]), .Z(N892) );
  OR2D0 C7933 ( .A1(g[892]), .A2(N892), .Z(c[893]) );
  AN2D0 C7932 ( .A1(p[891]), .A2(c[891]), .Z(N891) );
  OR2D0 C7931 ( .A1(g[891]), .A2(N891), .Z(c[892]) );
  AN2D0 C7930 ( .A1(p[890]), .A2(c[890]), .Z(N890) );
  OR2D0 C7929 ( .A1(g[890]), .A2(N890), .Z(c[891]) );
  AN2D0 C7928 ( .A1(p[889]), .A2(c[889]), .Z(N889) );
  OR2D0 C7927 ( .A1(g[889]), .A2(N889), .Z(c[890]) );
  AN2D0 C7926 ( .A1(p[888]), .A2(c[888]), .Z(N888) );
  OR2D0 C7925 ( .A1(g[888]), .A2(N888), .Z(c[889]) );
  AN2D0 C7924 ( .A1(p[887]), .A2(c[887]), .Z(N887) );
  OR2D0 C7923 ( .A1(g[887]), .A2(N887), .Z(c[888]) );
  AN2D0 C7922 ( .A1(p[886]), .A2(c[886]), .Z(N886) );
  OR2D0 C7921 ( .A1(g[886]), .A2(N886), .Z(c[887]) );
  AN2D0 C7920 ( .A1(p[885]), .A2(c[885]), .Z(N885) );
  OR2D0 C7919 ( .A1(g[885]), .A2(N885), .Z(c[886]) );
  AN2D0 C7918 ( .A1(p[884]), .A2(c[884]), .Z(N884) );
  OR2D0 C7917 ( .A1(g[884]), .A2(N884), .Z(c[885]) );
  AN2D0 C7916 ( .A1(p[883]), .A2(c[883]), .Z(N883) );
  OR2D0 C7915 ( .A1(g[883]), .A2(N883), .Z(c[884]) );
  AN2D0 C7914 ( .A1(p[882]), .A2(c[882]), .Z(N882) );
  OR2D0 C7913 ( .A1(g[882]), .A2(N882), .Z(c[883]) );
  AN2D0 C7912 ( .A1(p[881]), .A2(c[881]), .Z(N881) );
  OR2D0 C7911 ( .A1(g[881]), .A2(N881), .Z(c[882]) );
  AN2D0 C7910 ( .A1(p[880]), .A2(c[880]), .Z(N880) );
  OR2D0 C7909 ( .A1(g[880]), .A2(N880), .Z(c[881]) );
  AN2D0 C7908 ( .A1(p[879]), .A2(c[879]), .Z(N879) );
  OR2D0 C7907 ( .A1(g[879]), .A2(N879), .Z(c[880]) );
  AN2D0 C7906 ( .A1(p[878]), .A2(c[878]), .Z(N878) );
  OR2D0 C7905 ( .A1(g[878]), .A2(N878), .Z(c[879]) );
  AN2D0 C7904 ( .A1(p[877]), .A2(c[877]), .Z(N877) );
  OR2D0 C7903 ( .A1(g[877]), .A2(N877), .Z(c[878]) );
  AN2D0 C7902 ( .A1(p[876]), .A2(c[876]), .Z(N876) );
  OR2D0 C7901 ( .A1(g[876]), .A2(N876), .Z(c[877]) );
  AN2D0 C7900 ( .A1(p[875]), .A2(c[875]), .Z(N875) );
  OR2D0 C7899 ( .A1(g[875]), .A2(N875), .Z(c[876]) );
  AN2D0 C7898 ( .A1(p[874]), .A2(c[874]), .Z(N874) );
  OR2D0 C7897 ( .A1(g[874]), .A2(N874), .Z(c[875]) );
  AN2D0 C7896 ( .A1(p[873]), .A2(c[873]), .Z(N873) );
  OR2D0 C7895 ( .A1(g[873]), .A2(N873), .Z(c[874]) );
  AN2D0 C7894 ( .A1(p[872]), .A2(c[872]), .Z(N872) );
  OR2D0 C7893 ( .A1(g[872]), .A2(N872), .Z(c[873]) );
  AN2D0 C7892 ( .A1(p[871]), .A2(c[871]), .Z(N871) );
  OR2D0 C7891 ( .A1(g[871]), .A2(N871), .Z(c[872]) );
  AN2D0 C7890 ( .A1(p[870]), .A2(c[870]), .Z(N870) );
  OR2D0 C7889 ( .A1(g[870]), .A2(N870), .Z(c[871]) );
  AN2D0 C7888 ( .A1(p[869]), .A2(c[869]), .Z(N869) );
  OR2D0 C7887 ( .A1(g[869]), .A2(N869), .Z(c[870]) );
  AN2D0 C7886 ( .A1(p[868]), .A2(c[868]), .Z(N868) );
  OR2D0 C7885 ( .A1(g[868]), .A2(N868), .Z(c[869]) );
  AN2D0 C7884 ( .A1(p[867]), .A2(c[867]), .Z(N867) );
  OR2D0 C7883 ( .A1(g[867]), .A2(N867), .Z(c[868]) );
  AN2D0 C7882 ( .A1(p[866]), .A2(c[866]), .Z(N866) );
  OR2D0 C7881 ( .A1(g[866]), .A2(N866), .Z(c[867]) );
  AN2D0 C7880 ( .A1(p[865]), .A2(c[865]), .Z(N865) );
  OR2D0 C7879 ( .A1(g[865]), .A2(N865), .Z(c[866]) );
  AN2D0 C7878 ( .A1(p[864]), .A2(c[864]), .Z(N864) );
  OR2D0 C7877 ( .A1(g[864]), .A2(N864), .Z(c[865]) );
  AN2D0 C7876 ( .A1(p[863]), .A2(c[863]), .Z(N863) );
  OR2D0 C7875 ( .A1(g[863]), .A2(N863), .Z(c[864]) );
  AN2D0 C7874 ( .A1(p[862]), .A2(c[862]), .Z(N862) );
  OR2D0 C7873 ( .A1(g[862]), .A2(N862), .Z(c[863]) );
  AN2D0 C7872 ( .A1(p[861]), .A2(c[861]), .Z(N861) );
  OR2D0 C7871 ( .A1(g[861]), .A2(N861), .Z(c[862]) );
  AN2D0 C7870 ( .A1(p[860]), .A2(c[860]), .Z(N860) );
  OR2D0 C7869 ( .A1(g[860]), .A2(N860), .Z(c[861]) );
  AN2D0 C7868 ( .A1(p[859]), .A2(c[859]), .Z(N859) );
  OR2D0 C7867 ( .A1(g[859]), .A2(N859), .Z(c[860]) );
  AN2D0 C7866 ( .A1(p[858]), .A2(c[858]), .Z(N858) );
  OR2D0 C7865 ( .A1(g[858]), .A2(N858), .Z(c[859]) );
  AN2D0 C7864 ( .A1(p[857]), .A2(c[857]), .Z(N857) );
  OR2D0 C7863 ( .A1(g[857]), .A2(N857), .Z(c[858]) );
  AN2D0 C7862 ( .A1(p[856]), .A2(c[856]), .Z(N856) );
  OR2D0 C7861 ( .A1(g[856]), .A2(N856), .Z(c[857]) );
  AN2D0 C7860 ( .A1(p[855]), .A2(c[855]), .Z(N855) );
  OR2D0 C7859 ( .A1(g[855]), .A2(N855), .Z(c[856]) );
  AN2D0 C7858 ( .A1(p[854]), .A2(c[854]), .Z(N854) );
  OR2D0 C7857 ( .A1(g[854]), .A2(N854), .Z(c[855]) );
  AN2D0 C7856 ( .A1(p[853]), .A2(c[853]), .Z(N853) );
  OR2D0 C7855 ( .A1(g[853]), .A2(N853), .Z(c[854]) );
  AN2D0 C7854 ( .A1(p[852]), .A2(c[852]), .Z(N852) );
  OR2D0 C7853 ( .A1(g[852]), .A2(N852), .Z(c[853]) );
  AN2D0 C7852 ( .A1(p[851]), .A2(c[851]), .Z(N851) );
  OR2D0 C7851 ( .A1(g[851]), .A2(N851), .Z(c[852]) );
  AN2D0 C7850 ( .A1(p[850]), .A2(c[850]), .Z(N850) );
  OR2D0 C7849 ( .A1(g[850]), .A2(N850), .Z(c[851]) );
  AN2D0 C7848 ( .A1(p[849]), .A2(c[849]), .Z(N849) );
  OR2D0 C7847 ( .A1(g[849]), .A2(N849), .Z(c[850]) );
  AN2D0 C7846 ( .A1(p[848]), .A2(c[848]), .Z(N848) );
  OR2D0 C7845 ( .A1(g[848]), .A2(N848), .Z(c[849]) );
  AN2D0 C7844 ( .A1(p[847]), .A2(c[847]), .Z(N847) );
  OR2D0 C7843 ( .A1(g[847]), .A2(N847), .Z(c[848]) );
  AN2D0 C7842 ( .A1(p[846]), .A2(c[846]), .Z(N846) );
  OR2D0 C7841 ( .A1(g[846]), .A2(N846), .Z(c[847]) );
  AN2D0 C7840 ( .A1(p[845]), .A2(c[845]), .Z(N845) );
  OR2D0 C7839 ( .A1(g[845]), .A2(N845), .Z(c[846]) );
  AN2D0 C7838 ( .A1(p[844]), .A2(c[844]), .Z(N844) );
  OR2D0 C7837 ( .A1(g[844]), .A2(N844), .Z(c[845]) );
  AN2D0 C7836 ( .A1(p[843]), .A2(c[843]), .Z(N843) );
  OR2D0 C7835 ( .A1(g[843]), .A2(N843), .Z(c[844]) );
  AN2D0 C7834 ( .A1(p[842]), .A2(c[842]), .Z(N842) );
  OR2D0 C7833 ( .A1(g[842]), .A2(N842), .Z(c[843]) );
  AN2D0 C7832 ( .A1(p[841]), .A2(c[841]), .Z(N841) );
  OR2D0 C7831 ( .A1(g[841]), .A2(N841), .Z(c[842]) );
  AN2D0 C7830 ( .A1(p[840]), .A2(c[840]), .Z(N840) );
  OR2D0 C7829 ( .A1(g[840]), .A2(N840), .Z(c[841]) );
  AN2D0 C7828 ( .A1(p[839]), .A2(c[839]), .Z(N839) );
  OR2D0 C7827 ( .A1(g[839]), .A2(N839), .Z(c[840]) );
  AN2D0 C7826 ( .A1(p[838]), .A2(c[838]), .Z(N838) );
  OR2D0 C7825 ( .A1(g[838]), .A2(N838), .Z(c[839]) );
  AN2D0 C7824 ( .A1(p[837]), .A2(c[837]), .Z(N837) );
  OR2D0 C7823 ( .A1(g[837]), .A2(N837), .Z(c[838]) );
  AN2D0 C7822 ( .A1(p[836]), .A2(c[836]), .Z(N836) );
  OR2D0 C7821 ( .A1(g[836]), .A2(N836), .Z(c[837]) );
  AN2D0 C7820 ( .A1(p[835]), .A2(c[835]), .Z(N835) );
  OR2D0 C7819 ( .A1(g[835]), .A2(N835), .Z(c[836]) );
  AN2D0 C7818 ( .A1(p[834]), .A2(c[834]), .Z(N834) );
  OR2D0 C7817 ( .A1(g[834]), .A2(N834), .Z(c[835]) );
  AN2D0 C7816 ( .A1(p[833]), .A2(c[833]), .Z(N833) );
  OR2D0 C7815 ( .A1(g[833]), .A2(N833), .Z(c[834]) );
  AN2D0 C7814 ( .A1(p[832]), .A2(c[832]), .Z(N832) );
  OR2D0 C7813 ( .A1(g[832]), .A2(N832), .Z(c[833]) );
  AN2D0 C7812 ( .A1(p[831]), .A2(c[831]), .Z(N831) );
  OR2D0 C7811 ( .A1(g[831]), .A2(N831), .Z(c[832]) );
  AN2D0 C7810 ( .A1(p[830]), .A2(c[830]), .Z(N830) );
  OR2D0 C7809 ( .A1(g[830]), .A2(N830), .Z(c[831]) );
  AN2D0 C7808 ( .A1(p[829]), .A2(c[829]), .Z(N829) );
  OR2D0 C7807 ( .A1(g[829]), .A2(N829), .Z(c[830]) );
  AN2D0 C7806 ( .A1(p[828]), .A2(c[828]), .Z(N828) );
  OR2D0 C7805 ( .A1(g[828]), .A2(N828), .Z(c[829]) );
  AN2D0 C7804 ( .A1(p[827]), .A2(c[827]), .Z(N827) );
  OR2D0 C7803 ( .A1(g[827]), .A2(N827), .Z(c[828]) );
  AN2D0 C7802 ( .A1(p[826]), .A2(c[826]), .Z(N826) );
  OR2D0 C7801 ( .A1(g[826]), .A2(N826), .Z(c[827]) );
  AN2D0 C7800 ( .A1(p[825]), .A2(c[825]), .Z(N825) );
  OR2D0 C7799 ( .A1(g[825]), .A2(N825), .Z(c[826]) );
  AN2D0 C7798 ( .A1(p[824]), .A2(c[824]), .Z(N824) );
  OR2D0 C7797 ( .A1(g[824]), .A2(N824), .Z(c[825]) );
  AN2D0 C7796 ( .A1(p[823]), .A2(c[823]), .Z(N823) );
  OR2D0 C7795 ( .A1(g[823]), .A2(N823), .Z(c[824]) );
  AN2D0 C7794 ( .A1(p[822]), .A2(c[822]), .Z(N822) );
  OR2D0 C7793 ( .A1(g[822]), .A2(N822), .Z(c[823]) );
  AN2D0 C7792 ( .A1(p[821]), .A2(c[821]), .Z(N821) );
  OR2D0 C7791 ( .A1(g[821]), .A2(N821), .Z(c[822]) );
  AN2D0 C7790 ( .A1(p[820]), .A2(c[820]), .Z(N820) );
  OR2D0 C7789 ( .A1(g[820]), .A2(N820), .Z(c[821]) );
  AN2D0 C7788 ( .A1(p[819]), .A2(c[819]), .Z(N819) );
  OR2D0 C7787 ( .A1(g[819]), .A2(N819), .Z(c[820]) );
  AN2D0 C7786 ( .A1(p[818]), .A2(c[818]), .Z(N818) );
  OR2D0 C7785 ( .A1(g[818]), .A2(N818), .Z(c[819]) );
  AN2D0 C7784 ( .A1(p[817]), .A2(c[817]), .Z(N817) );
  OR2D0 C7783 ( .A1(g[817]), .A2(N817), .Z(c[818]) );
  AN2D0 C7782 ( .A1(p[816]), .A2(c[816]), .Z(N816) );
  OR2D0 C7781 ( .A1(g[816]), .A2(N816), .Z(c[817]) );
  AN2D0 C7780 ( .A1(p[815]), .A2(c[815]), .Z(N815) );
  OR2D0 C7779 ( .A1(g[815]), .A2(N815), .Z(c[816]) );
  AN2D0 C7778 ( .A1(p[814]), .A2(c[814]), .Z(N814) );
  OR2D0 C7777 ( .A1(g[814]), .A2(N814), .Z(c[815]) );
  AN2D0 C7776 ( .A1(p[813]), .A2(c[813]), .Z(N813) );
  OR2D0 C7775 ( .A1(g[813]), .A2(N813), .Z(c[814]) );
  AN2D0 C7774 ( .A1(p[812]), .A2(c[812]), .Z(N812) );
  OR2D0 C7773 ( .A1(g[812]), .A2(N812), .Z(c[813]) );
  AN2D0 C7772 ( .A1(p[811]), .A2(c[811]), .Z(N811) );
  OR2D0 C7771 ( .A1(g[811]), .A2(N811), .Z(c[812]) );
  AN2D0 C7770 ( .A1(p[810]), .A2(c[810]), .Z(N810) );
  OR2D0 C7769 ( .A1(g[810]), .A2(N810), .Z(c[811]) );
  AN2D0 C7768 ( .A1(p[809]), .A2(c[809]), .Z(N809) );
  OR2D0 C7767 ( .A1(g[809]), .A2(N809), .Z(c[810]) );
  AN2D0 C7766 ( .A1(p[808]), .A2(c[808]), .Z(N808) );
  OR2D0 C7765 ( .A1(g[808]), .A2(N808), .Z(c[809]) );
  AN2D0 C7764 ( .A1(p[807]), .A2(c[807]), .Z(N807) );
  OR2D0 C7763 ( .A1(g[807]), .A2(N807), .Z(c[808]) );
  AN2D0 C7762 ( .A1(p[806]), .A2(c[806]), .Z(N806) );
  OR2D0 C7761 ( .A1(g[806]), .A2(N806), .Z(c[807]) );
  AN2D0 C7760 ( .A1(p[805]), .A2(c[805]), .Z(N805) );
  OR2D0 C7759 ( .A1(g[805]), .A2(N805), .Z(c[806]) );
  AN2D0 C7758 ( .A1(p[804]), .A2(c[804]), .Z(N804) );
  OR2D0 C7757 ( .A1(g[804]), .A2(N804), .Z(c[805]) );
  AN2D0 C7756 ( .A1(p[803]), .A2(c[803]), .Z(N803) );
  OR2D0 C7755 ( .A1(g[803]), .A2(N803), .Z(c[804]) );
  AN2D0 C7754 ( .A1(p[802]), .A2(c[802]), .Z(N802) );
  OR2D0 C7753 ( .A1(g[802]), .A2(N802), .Z(c[803]) );
  AN2D0 C7752 ( .A1(p[801]), .A2(c[801]), .Z(N801) );
  OR2D0 C7751 ( .A1(g[801]), .A2(N801), .Z(c[802]) );
  AN2D0 C7750 ( .A1(p[800]), .A2(c[800]), .Z(N800) );
  OR2D0 C7749 ( .A1(g[800]), .A2(N800), .Z(c[801]) );
  AN2D0 C7748 ( .A1(p[799]), .A2(c[799]), .Z(N799) );
  OR2D0 C7747 ( .A1(g[799]), .A2(N799), .Z(c[800]) );
  AN2D0 C7746 ( .A1(p[798]), .A2(c[798]), .Z(N798) );
  OR2D0 C7745 ( .A1(g[798]), .A2(N798), .Z(c[799]) );
  AN2D0 C7744 ( .A1(p[797]), .A2(c[797]), .Z(N797) );
  OR2D0 C7743 ( .A1(g[797]), .A2(N797), .Z(c[798]) );
  AN2D0 C7742 ( .A1(p[796]), .A2(c[796]), .Z(N796) );
  OR2D0 C7741 ( .A1(g[796]), .A2(N796), .Z(c[797]) );
  AN2D0 C7740 ( .A1(p[795]), .A2(c[795]), .Z(N795) );
  OR2D0 C7739 ( .A1(g[795]), .A2(N795), .Z(c[796]) );
  AN2D0 C7738 ( .A1(p[794]), .A2(c[794]), .Z(N794) );
  OR2D0 C7737 ( .A1(g[794]), .A2(N794), .Z(c[795]) );
  AN2D0 C7736 ( .A1(p[793]), .A2(c[793]), .Z(N793) );
  OR2D0 C7735 ( .A1(g[793]), .A2(N793), .Z(c[794]) );
  AN2D0 C7734 ( .A1(p[792]), .A2(c[792]), .Z(N792) );
  OR2D0 C7733 ( .A1(g[792]), .A2(N792), .Z(c[793]) );
  AN2D0 C7732 ( .A1(p[791]), .A2(c[791]), .Z(N791) );
  OR2D0 C7731 ( .A1(g[791]), .A2(N791), .Z(c[792]) );
  AN2D0 C7730 ( .A1(p[790]), .A2(c[790]), .Z(N790) );
  OR2D0 C7729 ( .A1(g[790]), .A2(N790), .Z(c[791]) );
  AN2D0 C7728 ( .A1(p[789]), .A2(c[789]), .Z(N789) );
  OR2D0 C7727 ( .A1(g[789]), .A2(N789), .Z(c[790]) );
  AN2D0 C7726 ( .A1(p[788]), .A2(c[788]), .Z(N788) );
  OR2D0 C7725 ( .A1(g[788]), .A2(N788), .Z(c[789]) );
  AN2D0 C7724 ( .A1(p[787]), .A2(c[787]), .Z(N787) );
  OR2D0 C7723 ( .A1(g[787]), .A2(N787), .Z(c[788]) );
  AN2D0 C7722 ( .A1(p[786]), .A2(c[786]), .Z(N786) );
  OR2D0 C7721 ( .A1(g[786]), .A2(N786), .Z(c[787]) );
  AN2D0 C7720 ( .A1(p[785]), .A2(c[785]), .Z(N785) );
  OR2D0 C7719 ( .A1(g[785]), .A2(N785), .Z(c[786]) );
  AN2D0 C7718 ( .A1(p[784]), .A2(c[784]), .Z(N784) );
  OR2D0 C7717 ( .A1(g[784]), .A2(N784), .Z(c[785]) );
  AN2D0 C7716 ( .A1(p[783]), .A2(c[783]), .Z(N783) );
  OR2D0 C7715 ( .A1(g[783]), .A2(N783), .Z(c[784]) );
  AN2D0 C7714 ( .A1(p[782]), .A2(c[782]), .Z(N782) );
  OR2D0 C7713 ( .A1(g[782]), .A2(N782), .Z(c[783]) );
  AN2D0 C7712 ( .A1(p[781]), .A2(c[781]), .Z(N781) );
  OR2D0 C7711 ( .A1(g[781]), .A2(N781), .Z(c[782]) );
  AN2D0 C7710 ( .A1(p[780]), .A2(c[780]), .Z(N780) );
  OR2D0 C7709 ( .A1(g[780]), .A2(N780), .Z(c[781]) );
  AN2D0 C7708 ( .A1(p[779]), .A2(c[779]), .Z(N779) );
  OR2D0 C7707 ( .A1(g[779]), .A2(N779), .Z(c[780]) );
  AN2D0 C7706 ( .A1(p[778]), .A2(c[778]), .Z(N778) );
  OR2D0 C7705 ( .A1(g[778]), .A2(N778), .Z(c[779]) );
  AN2D0 C7704 ( .A1(p[777]), .A2(c[777]), .Z(N777) );
  OR2D0 C7703 ( .A1(g[777]), .A2(N777), .Z(c[778]) );
  AN2D0 C7702 ( .A1(p[776]), .A2(c[776]), .Z(N776) );
  OR2D0 C7701 ( .A1(g[776]), .A2(N776), .Z(c[777]) );
  AN2D0 C7700 ( .A1(p[775]), .A2(c[775]), .Z(N775) );
  OR2D0 C7699 ( .A1(g[775]), .A2(N775), .Z(c[776]) );
  AN2D0 C7698 ( .A1(p[774]), .A2(c[774]), .Z(N774) );
  OR2D0 C7697 ( .A1(g[774]), .A2(N774), .Z(c[775]) );
  AN2D0 C7696 ( .A1(p[773]), .A2(c[773]), .Z(N773) );
  OR2D0 C7695 ( .A1(g[773]), .A2(N773), .Z(c[774]) );
  AN2D0 C7694 ( .A1(p[772]), .A2(c[772]), .Z(N772) );
  OR2D0 C7693 ( .A1(g[772]), .A2(N772), .Z(c[773]) );
  AN2D0 C7692 ( .A1(p[771]), .A2(c[771]), .Z(N771) );
  OR2D0 C7691 ( .A1(g[771]), .A2(N771), .Z(c[772]) );
  AN2D0 C7690 ( .A1(p[770]), .A2(c[770]), .Z(N770) );
  OR2D0 C7689 ( .A1(g[770]), .A2(N770), .Z(c[771]) );
  AN2D0 C7688 ( .A1(p[769]), .A2(c[769]), .Z(N769) );
  OR2D0 C7687 ( .A1(g[769]), .A2(N769), .Z(c[770]) );
  AN2D0 C7686 ( .A1(p[768]), .A2(c[768]), .Z(N768) );
  OR2D0 C7685 ( .A1(g[768]), .A2(N768), .Z(c[769]) );
  AN2D0 C7684 ( .A1(p[767]), .A2(c[767]), .Z(N767) );
  OR2D0 C7683 ( .A1(g[767]), .A2(N767), .Z(c[768]) );
  AN2D0 C7682 ( .A1(p[766]), .A2(c[766]), .Z(N766) );
  OR2D0 C7681 ( .A1(g[766]), .A2(N766), .Z(c[767]) );
  AN2D0 C7680 ( .A1(p[765]), .A2(c[765]), .Z(N765) );
  OR2D0 C7679 ( .A1(g[765]), .A2(N765), .Z(c[766]) );
  AN2D0 C7678 ( .A1(p[764]), .A2(c[764]), .Z(N764) );
  OR2D0 C7677 ( .A1(g[764]), .A2(N764), .Z(c[765]) );
  AN2D0 C7676 ( .A1(p[763]), .A2(c[763]), .Z(N763) );
  OR2D0 C7675 ( .A1(g[763]), .A2(N763), .Z(c[764]) );
  AN2D0 C7674 ( .A1(p[762]), .A2(c[762]), .Z(N762) );
  OR2D0 C7673 ( .A1(g[762]), .A2(N762), .Z(c[763]) );
  AN2D0 C7672 ( .A1(p[761]), .A2(c[761]), .Z(N761) );
  OR2D0 C7671 ( .A1(g[761]), .A2(N761), .Z(c[762]) );
  AN2D0 C7670 ( .A1(p[760]), .A2(c[760]), .Z(N760) );
  OR2D0 C7669 ( .A1(g[760]), .A2(N760), .Z(c[761]) );
  AN2D0 C7668 ( .A1(p[759]), .A2(c[759]), .Z(N759) );
  OR2D0 C7667 ( .A1(g[759]), .A2(N759), .Z(c[760]) );
  AN2D0 C7666 ( .A1(p[758]), .A2(c[758]), .Z(N758) );
  OR2D0 C7665 ( .A1(g[758]), .A2(N758), .Z(c[759]) );
  AN2D0 C7664 ( .A1(p[757]), .A2(c[757]), .Z(N757) );
  OR2D0 C7663 ( .A1(g[757]), .A2(N757), .Z(c[758]) );
  AN2D0 C7662 ( .A1(p[756]), .A2(c[756]), .Z(N756) );
  OR2D0 C7661 ( .A1(g[756]), .A2(N756), .Z(c[757]) );
  AN2D0 C7660 ( .A1(p[755]), .A2(c[755]), .Z(N755) );
  OR2D0 C7659 ( .A1(g[755]), .A2(N755), .Z(c[756]) );
  AN2D0 C7658 ( .A1(p[754]), .A2(c[754]), .Z(N754) );
  OR2D0 C7657 ( .A1(g[754]), .A2(N754), .Z(c[755]) );
  AN2D0 C7656 ( .A1(p[753]), .A2(c[753]), .Z(N753) );
  OR2D0 C7655 ( .A1(g[753]), .A2(N753), .Z(c[754]) );
  AN2D0 C7654 ( .A1(p[752]), .A2(c[752]), .Z(N752) );
  OR2D0 C7653 ( .A1(g[752]), .A2(N752), .Z(c[753]) );
  AN2D0 C7652 ( .A1(p[751]), .A2(c[751]), .Z(N751) );
  OR2D0 C7651 ( .A1(g[751]), .A2(N751), .Z(c[752]) );
  AN2D0 C7650 ( .A1(p[750]), .A2(c[750]), .Z(N750) );
  OR2D0 C7649 ( .A1(g[750]), .A2(N750), .Z(c[751]) );
  AN2D0 C7648 ( .A1(p[749]), .A2(c[749]), .Z(N749) );
  OR2D0 C7647 ( .A1(g[749]), .A2(N749), .Z(c[750]) );
  AN2D0 C7646 ( .A1(p[748]), .A2(c[748]), .Z(N748) );
  OR2D0 C7645 ( .A1(g[748]), .A2(N748), .Z(c[749]) );
  AN2D0 C7644 ( .A1(p[747]), .A2(c[747]), .Z(N747) );
  OR2D0 C7643 ( .A1(g[747]), .A2(N747), .Z(c[748]) );
  AN2D0 C7642 ( .A1(p[746]), .A2(c[746]), .Z(N746) );
  OR2D0 C7641 ( .A1(g[746]), .A2(N746), .Z(c[747]) );
  AN2D0 C7640 ( .A1(p[745]), .A2(c[745]), .Z(N745) );
  OR2D0 C7639 ( .A1(g[745]), .A2(N745), .Z(c[746]) );
  AN2D0 C7638 ( .A1(p[744]), .A2(c[744]), .Z(N744) );
  OR2D0 C7637 ( .A1(g[744]), .A2(N744), .Z(c[745]) );
  AN2D0 C7636 ( .A1(p[743]), .A2(c[743]), .Z(N743) );
  OR2D0 C7635 ( .A1(g[743]), .A2(N743), .Z(c[744]) );
  AN2D0 C7634 ( .A1(p[742]), .A2(c[742]), .Z(N742) );
  OR2D0 C7633 ( .A1(g[742]), .A2(N742), .Z(c[743]) );
  AN2D0 C7632 ( .A1(p[741]), .A2(c[741]), .Z(N741) );
  OR2D0 C7631 ( .A1(g[741]), .A2(N741), .Z(c[742]) );
  AN2D0 C7630 ( .A1(p[740]), .A2(c[740]), .Z(N740) );
  OR2D0 C7629 ( .A1(g[740]), .A2(N740), .Z(c[741]) );
  AN2D0 C7628 ( .A1(p[739]), .A2(c[739]), .Z(N739) );
  OR2D0 C7627 ( .A1(g[739]), .A2(N739), .Z(c[740]) );
  AN2D0 C7626 ( .A1(p[738]), .A2(c[738]), .Z(N738) );
  OR2D0 C7625 ( .A1(g[738]), .A2(N738), .Z(c[739]) );
  AN2D0 C7624 ( .A1(p[737]), .A2(c[737]), .Z(N737) );
  OR2D0 C7623 ( .A1(g[737]), .A2(N737), .Z(c[738]) );
  AN2D0 C7622 ( .A1(p[736]), .A2(c[736]), .Z(N736) );
  OR2D0 C7621 ( .A1(g[736]), .A2(N736), .Z(c[737]) );
  AN2D0 C7620 ( .A1(p[735]), .A2(c[735]), .Z(N735) );
  OR2D0 C7619 ( .A1(g[735]), .A2(N735), .Z(c[736]) );
  AN2D0 C7618 ( .A1(p[734]), .A2(c[734]), .Z(N734) );
  OR2D0 C7617 ( .A1(g[734]), .A2(N734), .Z(c[735]) );
  AN2D0 C7616 ( .A1(p[733]), .A2(c[733]), .Z(N733) );
  OR2D0 C7615 ( .A1(g[733]), .A2(N733), .Z(c[734]) );
  AN2D0 C7614 ( .A1(p[732]), .A2(c[732]), .Z(N732) );
  OR2D0 C7613 ( .A1(g[732]), .A2(N732), .Z(c[733]) );
  AN2D0 C7612 ( .A1(p[731]), .A2(c[731]), .Z(N731) );
  OR2D0 C7611 ( .A1(g[731]), .A2(N731), .Z(c[732]) );
  AN2D0 C7610 ( .A1(p[730]), .A2(c[730]), .Z(N730) );
  OR2D0 C7609 ( .A1(g[730]), .A2(N730), .Z(c[731]) );
  AN2D0 C7608 ( .A1(p[729]), .A2(c[729]), .Z(N729) );
  OR2D0 C7607 ( .A1(g[729]), .A2(N729), .Z(c[730]) );
  AN2D0 C7606 ( .A1(p[728]), .A2(c[728]), .Z(N728) );
  OR2D0 C7605 ( .A1(g[728]), .A2(N728), .Z(c[729]) );
  AN2D0 C7604 ( .A1(p[727]), .A2(c[727]), .Z(N727) );
  OR2D0 C7603 ( .A1(g[727]), .A2(N727), .Z(c[728]) );
  AN2D0 C7602 ( .A1(p[726]), .A2(c[726]), .Z(N726) );
  OR2D0 C7601 ( .A1(g[726]), .A2(N726), .Z(c[727]) );
  AN2D0 C7600 ( .A1(p[725]), .A2(c[725]), .Z(N725) );
  OR2D0 C7599 ( .A1(g[725]), .A2(N725), .Z(c[726]) );
  AN2D0 C7598 ( .A1(p[724]), .A2(c[724]), .Z(N724) );
  OR2D0 C7597 ( .A1(g[724]), .A2(N724), .Z(c[725]) );
  AN2D0 C7596 ( .A1(p[723]), .A2(c[723]), .Z(N723) );
  OR2D0 C7595 ( .A1(g[723]), .A2(N723), .Z(c[724]) );
  AN2D0 C7594 ( .A1(p[722]), .A2(c[722]), .Z(N722) );
  OR2D0 C7593 ( .A1(g[722]), .A2(N722), .Z(c[723]) );
  AN2D0 C7592 ( .A1(p[721]), .A2(c[721]), .Z(N721) );
  OR2D0 C7591 ( .A1(g[721]), .A2(N721), .Z(c[722]) );
  AN2D0 C7590 ( .A1(p[720]), .A2(c[720]), .Z(N720) );
  OR2D0 C7589 ( .A1(g[720]), .A2(N720), .Z(c[721]) );
  AN2D0 C7588 ( .A1(p[719]), .A2(c[719]), .Z(N719) );
  OR2D0 C7587 ( .A1(g[719]), .A2(N719), .Z(c[720]) );
  AN2D0 C7586 ( .A1(p[718]), .A2(c[718]), .Z(N718) );
  OR2D0 C7585 ( .A1(g[718]), .A2(N718), .Z(c[719]) );
  AN2D0 C7584 ( .A1(p[717]), .A2(c[717]), .Z(N717) );
  OR2D0 C7583 ( .A1(g[717]), .A2(N717), .Z(c[718]) );
  AN2D0 C7582 ( .A1(p[716]), .A2(c[716]), .Z(N716) );
  OR2D0 C7581 ( .A1(g[716]), .A2(N716), .Z(c[717]) );
  AN2D0 C7580 ( .A1(p[715]), .A2(c[715]), .Z(N715) );
  OR2D0 C7579 ( .A1(g[715]), .A2(N715), .Z(c[716]) );
  AN2D0 C7578 ( .A1(p[714]), .A2(c[714]), .Z(N714) );
  OR2D0 C7577 ( .A1(g[714]), .A2(N714), .Z(c[715]) );
  AN2D0 C7576 ( .A1(p[713]), .A2(c[713]), .Z(N713) );
  OR2D0 C7575 ( .A1(g[713]), .A2(N713), .Z(c[714]) );
  AN2D0 C7574 ( .A1(p[712]), .A2(c[712]), .Z(N712) );
  OR2D0 C7573 ( .A1(g[712]), .A2(N712), .Z(c[713]) );
  AN2D0 C7572 ( .A1(p[711]), .A2(c[711]), .Z(N711) );
  OR2D0 C7571 ( .A1(g[711]), .A2(N711), .Z(c[712]) );
  AN2D0 C7570 ( .A1(p[710]), .A2(c[710]), .Z(N710) );
  OR2D0 C7569 ( .A1(g[710]), .A2(N710), .Z(c[711]) );
  AN2D0 C7568 ( .A1(p[709]), .A2(c[709]), .Z(N709) );
  OR2D0 C7567 ( .A1(g[709]), .A2(N709), .Z(c[710]) );
  AN2D0 C7566 ( .A1(p[708]), .A2(c[708]), .Z(N708) );
  OR2D0 C7565 ( .A1(g[708]), .A2(N708), .Z(c[709]) );
  AN2D0 C7564 ( .A1(p[707]), .A2(c[707]), .Z(N707) );
  OR2D0 C7563 ( .A1(g[707]), .A2(N707), .Z(c[708]) );
  AN2D0 C7562 ( .A1(p[706]), .A2(c[706]), .Z(N706) );
  OR2D0 C7561 ( .A1(g[706]), .A2(N706), .Z(c[707]) );
  AN2D0 C7560 ( .A1(p[705]), .A2(c[705]), .Z(N705) );
  OR2D0 C7559 ( .A1(g[705]), .A2(N705), .Z(c[706]) );
  AN2D0 C7558 ( .A1(p[704]), .A2(c[704]), .Z(N704) );
  OR2D0 C7557 ( .A1(g[704]), .A2(N704), .Z(c[705]) );
  AN2D0 C7556 ( .A1(p[703]), .A2(c[703]), .Z(N703) );
  OR2D0 C7555 ( .A1(g[703]), .A2(N703), .Z(c[704]) );
  AN2D0 C7554 ( .A1(p[702]), .A2(c[702]), .Z(N702) );
  OR2D0 C7553 ( .A1(g[702]), .A2(N702), .Z(c[703]) );
  AN2D0 C7552 ( .A1(p[701]), .A2(c[701]), .Z(N701) );
  OR2D0 C7551 ( .A1(g[701]), .A2(N701), .Z(c[702]) );
  AN2D0 C7550 ( .A1(p[700]), .A2(c[700]), .Z(N700) );
  OR2D0 C7549 ( .A1(g[700]), .A2(N700), .Z(c[701]) );
  AN2D0 C7548 ( .A1(p[699]), .A2(c[699]), .Z(N699) );
  OR2D0 C7547 ( .A1(g[699]), .A2(N699), .Z(c[700]) );
  AN2D0 C7546 ( .A1(p[698]), .A2(c[698]), .Z(N698) );
  OR2D0 C7545 ( .A1(g[698]), .A2(N698), .Z(c[699]) );
  AN2D0 C7544 ( .A1(p[697]), .A2(c[697]), .Z(N697) );
  OR2D0 C7543 ( .A1(g[697]), .A2(N697), .Z(c[698]) );
  AN2D0 C7542 ( .A1(p[696]), .A2(c[696]), .Z(N696) );
  OR2D0 C7541 ( .A1(g[696]), .A2(N696), .Z(c[697]) );
  AN2D0 C7540 ( .A1(p[695]), .A2(c[695]), .Z(N695) );
  OR2D0 C7539 ( .A1(g[695]), .A2(N695), .Z(c[696]) );
  AN2D0 C7538 ( .A1(p[694]), .A2(c[694]), .Z(N694) );
  OR2D0 C7537 ( .A1(g[694]), .A2(N694), .Z(c[695]) );
  AN2D0 C7536 ( .A1(p[693]), .A2(c[693]), .Z(N693) );
  OR2D0 C7535 ( .A1(g[693]), .A2(N693), .Z(c[694]) );
  AN2D0 C7534 ( .A1(p[692]), .A2(c[692]), .Z(N692) );
  OR2D0 C7533 ( .A1(g[692]), .A2(N692), .Z(c[693]) );
  AN2D0 C7532 ( .A1(p[691]), .A2(c[691]), .Z(N691) );
  OR2D0 C7531 ( .A1(g[691]), .A2(N691), .Z(c[692]) );
  AN2D0 C7530 ( .A1(p[690]), .A2(c[690]), .Z(N690) );
  OR2D0 C7529 ( .A1(g[690]), .A2(N690), .Z(c[691]) );
  AN2D0 C7528 ( .A1(p[689]), .A2(c[689]), .Z(N689) );
  OR2D0 C7527 ( .A1(g[689]), .A2(N689), .Z(c[690]) );
  AN2D0 C7526 ( .A1(p[688]), .A2(c[688]), .Z(N688) );
  OR2D0 C7525 ( .A1(g[688]), .A2(N688), .Z(c[689]) );
  AN2D0 C7524 ( .A1(p[687]), .A2(c[687]), .Z(N687) );
  OR2D0 C7523 ( .A1(g[687]), .A2(N687), .Z(c[688]) );
  AN2D0 C7522 ( .A1(p[686]), .A2(c[686]), .Z(N686) );
  OR2D0 C7521 ( .A1(g[686]), .A2(N686), .Z(c[687]) );
  AN2D0 C7520 ( .A1(p[685]), .A2(c[685]), .Z(N685) );
  OR2D0 C7519 ( .A1(g[685]), .A2(N685), .Z(c[686]) );
  AN2D0 C7518 ( .A1(p[684]), .A2(c[684]), .Z(N684) );
  OR2D0 C7517 ( .A1(g[684]), .A2(N684), .Z(c[685]) );
  AN2D0 C7516 ( .A1(p[683]), .A2(c[683]), .Z(N683) );
  OR2D0 C7515 ( .A1(g[683]), .A2(N683), .Z(c[684]) );
  AN2D0 C7514 ( .A1(p[682]), .A2(c[682]), .Z(N682) );
  OR2D0 C7513 ( .A1(g[682]), .A2(N682), .Z(c[683]) );
  AN2D0 C7512 ( .A1(p[681]), .A2(c[681]), .Z(N681) );
  OR2D0 C7511 ( .A1(g[681]), .A2(N681), .Z(c[682]) );
  AN2D0 C7510 ( .A1(p[680]), .A2(c[680]), .Z(N680) );
  OR2D0 C7509 ( .A1(g[680]), .A2(N680), .Z(c[681]) );
  AN2D0 C7508 ( .A1(p[679]), .A2(c[679]), .Z(N679) );
  OR2D0 C7507 ( .A1(g[679]), .A2(N679), .Z(c[680]) );
  AN2D0 C7506 ( .A1(p[678]), .A2(c[678]), .Z(N678) );
  OR2D0 C7505 ( .A1(g[678]), .A2(N678), .Z(c[679]) );
  AN2D0 C7504 ( .A1(p[677]), .A2(c[677]), .Z(N677) );
  OR2D0 C7503 ( .A1(g[677]), .A2(N677), .Z(c[678]) );
  AN2D0 C7502 ( .A1(p[676]), .A2(c[676]), .Z(N676) );
  OR2D0 C7501 ( .A1(g[676]), .A2(N676), .Z(c[677]) );
  AN2D0 C7500 ( .A1(p[675]), .A2(c[675]), .Z(N675) );
  OR2D0 C7499 ( .A1(g[675]), .A2(N675), .Z(c[676]) );
  AN2D0 C7498 ( .A1(p[674]), .A2(c[674]), .Z(N674) );
  OR2D0 C7497 ( .A1(g[674]), .A2(N674), .Z(c[675]) );
  AN2D0 C7496 ( .A1(p[673]), .A2(c[673]), .Z(N673) );
  OR2D0 C7495 ( .A1(g[673]), .A2(N673), .Z(c[674]) );
  AN2D0 C7494 ( .A1(p[672]), .A2(c[672]), .Z(N672) );
  OR2D0 C7493 ( .A1(g[672]), .A2(N672), .Z(c[673]) );
  AN2D0 C7492 ( .A1(p[671]), .A2(c[671]), .Z(N671) );
  OR2D0 C7491 ( .A1(g[671]), .A2(N671), .Z(c[672]) );
  AN2D0 C7490 ( .A1(p[670]), .A2(c[670]), .Z(N670) );
  OR2D0 C7489 ( .A1(g[670]), .A2(N670), .Z(c[671]) );
  AN2D0 C7488 ( .A1(p[669]), .A2(c[669]), .Z(N669) );
  OR2D0 C7487 ( .A1(g[669]), .A2(N669), .Z(c[670]) );
  AN2D0 C7486 ( .A1(p[668]), .A2(c[668]), .Z(N668) );
  OR2D0 C7485 ( .A1(g[668]), .A2(N668), .Z(c[669]) );
  AN2D0 C7484 ( .A1(p[667]), .A2(c[667]), .Z(N667) );
  OR2D0 C7483 ( .A1(g[667]), .A2(N667), .Z(c[668]) );
  AN2D0 C7482 ( .A1(p[666]), .A2(c[666]), .Z(N666) );
  OR2D0 C7481 ( .A1(g[666]), .A2(N666), .Z(c[667]) );
  AN2D0 C7480 ( .A1(p[665]), .A2(c[665]), .Z(N665) );
  OR2D0 C7479 ( .A1(g[665]), .A2(N665), .Z(c[666]) );
  AN2D0 C7478 ( .A1(p[664]), .A2(c[664]), .Z(N664) );
  OR2D0 C7477 ( .A1(g[664]), .A2(N664), .Z(c[665]) );
  AN2D0 C7476 ( .A1(p[663]), .A2(c[663]), .Z(N663) );
  OR2D0 C7475 ( .A1(g[663]), .A2(N663), .Z(c[664]) );
  AN2D0 C7474 ( .A1(p[662]), .A2(c[662]), .Z(N662) );
  OR2D0 C7473 ( .A1(g[662]), .A2(N662), .Z(c[663]) );
  AN2D0 C7472 ( .A1(p[661]), .A2(c[661]), .Z(N661) );
  OR2D0 C7471 ( .A1(g[661]), .A2(N661), .Z(c[662]) );
  AN2D0 C7470 ( .A1(p[660]), .A2(c[660]), .Z(N660) );
  OR2D0 C7469 ( .A1(g[660]), .A2(N660), .Z(c[661]) );
  AN2D0 C7468 ( .A1(p[659]), .A2(c[659]), .Z(N659) );
  OR2D0 C7467 ( .A1(g[659]), .A2(N659), .Z(c[660]) );
  AN2D0 C7466 ( .A1(p[658]), .A2(c[658]), .Z(N658) );
  OR2D0 C7465 ( .A1(g[658]), .A2(N658), .Z(c[659]) );
  AN2D0 C7464 ( .A1(p[657]), .A2(c[657]), .Z(N657) );
  OR2D0 C7463 ( .A1(g[657]), .A2(N657), .Z(c[658]) );
  AN2D0 C7462 ( .A1(p[656]), .A2(c[656]), .Z(N656) );
  OR2D0 C7461 ( .A1(g[656]), .A2(N656), .Z(c[657]) );
  AN2D0 C7460 ( .A1(p[655]), .A2(c[655]), .Z(N655) );
  OR2D0 C7459 ( .A1(g[655]), .A2(N655), .Z(c[656]) );
  AN2D0 C7458 ( .A1(p[654]), .A2(c[654]), .Z(N654) );
  OR2D0 C7457 ( .A1(g[654]), .A2(N654), .Z(c[655]) );
  AN2D0 C7456 ( .A1(p[653]), .A2(c[653]), .Z(N653) );
  OR2D0 C7455 ( .A1(g[653]), .A2(N653), .Z(c[654]) );
  AN2D0 C7454 ( .A1(p[652]), .A2(c[652]), .Z(N652) );
  OR2D0 C7453 ( .A1(g[652]), .A2(N652), .Z(c[653]) );
  AN2D0 C7452 ( .A1(p[651]), .A2(c[651]), .Z(N651) );
  OR2D0 C7451 ( .A1(g[651]), .A2(N651), .Z(c[652]) );
  AN2D0 C7450 ( .A1(p[650]), .A2(c[650]), .Z(N650) );
  OR2D0 C7449 ( .A1(g[650]), .A2(N650), .Z(c[651]) );
  AN2D0 C7448 ( .A1(p[649]), .A2(c[649]), .Z(N649) );
  OR2D0 C7447 ( .A1(g[649]), .A2(N649), .Z(c[650]) );
  AN2D0 C7446 ( .A1(p[648]), .A2(c[648]), .Z(N648) );
  OR2D0 C7445 ( .A1(g[648]), .A2(N648), .Z(c[649]) );
  AN2D0 C7444 ( .A1(p[647]), .A2(c[647]), .Z(N647) );
  OR2D0 C7443 ( .A1(g[647]), .A2(N647), .Z(c[648]) );
  AN2D0 C7442 ( .A1(p[646]), .A2(c[646]), .Z(N646) );
  OR2D0 C7441 ( .A1(g[646]), .A2(N646), .Z(c[647]) );
  AN2D0 C7440 ( .A1(p[645]), .A2(c[645]), .Z(N645) );
  OR2D0 C7439 ( .A1(g[645]), .A2(N645), .Z(c[646]) );
  AN2D0 C7438 ( .A1(p[644]), .A2(c[644]), .Z(N644) );
  OR2D0 C7437 ( .A1(g[644]), .A2(N644), .Z(c[645]) );
  AN2D0 C7436 ( .A1(p[643]), .A2(c[643]), .Z(N643) );
  OR2D0 C7435 ( .A1(g[643]), .A2(N643), .Z(c[644]) );
  AN2D0 C7434 ( .A1(p[642]), .A2(c[642]), .Z(N642) );
  OR2D0 C7433 ( .A1(g[642]), .A2(N642), .Z(c[643]) );
  AN2D0 C7432 ( .A1(p[641]), .A2(c[641]), .Z(N641) );
  OR2D0 C7431 ( .A1(g[641]), .A2(N641), .Z(c[642]) );
  AN2D0 C7430 ( .A1(p[640]), .A2(c[640]), .Z(N640) );
  OR2D0 C7429 ( .A1(g[640]), .A2(N640), .Z(c[641]) );
  AN2D0 C7428 ( .A1(p[639]), .A2(c[639]), .Z(N639) );
  OR2D0 C7427 ( .A1(g[639]), .A2(N639), .Z(c[640]) );
  AN2D0 C7426 ( .A1(p[638]), .A2(c[638]), .Z(N638) );
  OR2D0 C7425 ( .A1(g[638]), .A2(N638), .Z(c[639]) );
  AN2D0 C7424 ( .A1(p[637]), .A2(c[637]), .Z(N637) );
  OR2D0 C7423 ( .A1(g[637]), .A2(N637), .Z(c[638]) );
  AN2D0 C7422 ( .A1(p[636]), .A2(c[636]), .Z(N636) );
  OR2D0 C7421 ( .A1(g[636]), .A2(N636), .Z(c[637]) );
  AN2D0 C7420 ( .A1(p[635]), .A2(c[635]), .Z(N635) );
  OR2D0 C7419 ( .A1(g[635]), .A2(N635), .Z(c[636]) );
  AN2D0 C7418 ( .A1(p[634]), .A2(c[634]), .Z(N634) );
  OR2D0 C7417 ( .A1(g[634]), .A2(N634), .Z(c[635]) );
  AN2D0 C7416 ( .A1(p[633]), .A2(c[633]), .Z(N633) );
  OR2D0 C7415 ( .A1(g[633]), .A2(N633), .Z(c[634]) );
  AN2D0 C7414 ( .A1(p[632]), .A2(c[632]), .Z(N632) );
  OR2D0 C7413 ( .A1(g[632]), .A2(N632), .Z(c[633]) );
  AN2D0 C7412 ( .A1(p[631]), .A2(c[631]), .Z(N631) );
  OR2D0 C7411 ( .A1(g[631]), .A2(N631), .Z(c[632]) );
  AN2D0 C7410 ( .A1(p[630]), .A2(c[630]), .Z(N630) );
  OR2D0 C7409 ( .A1(g[630]), .A2(N630), .Z(c[631]) );
  AN2D0 C7408 ( .A1(p[629]), .A2(c[629]), .Z(N629) );
  OR2D0 C7407 ( .A1(g[629]), .A2(N629), .Z(c[630]) );
  AN2D0 C7406 ( .A1(p[628]), .A2(c[628]), .Z(N628) );
  OR2D0 C7405 ( .A1(g[628]), .A2(N628), .Z(c[629]) );
  AN2D0 C7404 ( .A1(p[627]), .A2(c[627]), .Z(N627) );
  OR2D0 C7403 ( .A1(g[627]), .A2(N627), .Z(c[628]) );
  AN2D0 C7402 ( .A1(p[626]), .A2(c[626]), .Z(N626) );
  OR2D0 C7401 ( .A1(g[626]), .A2(N626), .Z(c[627]) );
  AN2D0 C7400 ( .A1(p[625]), .A2(c[625]), .Z(N625) );
  OR2D0 C7399 ( .A1(g[625]), .A2(N625), .Z(c[626]) );
  AN2D0 C7398 ( .A1(p[624]), .A2(c[624]), .Z(N624) );
  OR2D0 C7397 ( .A1(g[624]), .A2(N624), .Z(c[625]) );
  AN2D0 C7396 ( .A1(p[623]), .A2(c[623]), .Z(N623) );
  OR2D0 C7395 ( .A1(g[623]), .A2(N623), .Z(c[624]) );
  AN2D0 C7394 ( .A1(p[622]), .A2(c[622]), .Z(N622) );
  OR2D0 C7393 ( .A1(g[622]), .A2(N622), .Z(c[623]) );
  AN2D0 C7392 ( .A1(p[621]), .A2(c[621]), .Z(N621) );
  OR2D0 C7391 ( .A1(g[621]), .A2(N621), .Z(c[622]) );
  AN2D0 C7390 ( .A1(p[620]), .A2(c[620]), .Z(N620) );
  OR2D0 C7389 ( .A1(g[620]), .A2(N620), .Z(c[621]) );
  AN2D0 C7388 ( .A1(p[619]), .A2(c[619]), .Z(N619) );
  OR2D0 C7387 ( .A1(g[619]), .A2(N619), .Z(c[620]) );
  AN2D0 C7386 ( .A1(p[618]), .A2(c[618]), .Z(N618) );
  OR2D0 C7385 ( .A1(g[618]), .A2(N618), .Z(c[619]) );
  AN2D0 C7384 ( .A1(p[617]), .A2(c[617]), .Z(N617) );
  OR2D0 C7383 ( .A1(g[617]), .A2(N617), .Z(c[618]) );
  AN2D0 C7382 ( .A1(p[616]), .A2(c[616]), .Z(N616) );
  OR2D0 C7381 ( .A1(g[616]), .A2(N616), .Z(c[617]) );
  AN2D0 C7380 ( .A1(p[615]), .A2(c[615]), .Z(N615) );
  OR2D0 C7379 ( .A1(g[615]), .A2(N615), .Z(c[616]) );
  AN2D0 C7378 ( .A1(p[614]), .A2(c[614]), .Z(N614) );
  OR2D0 C7377 ( .A1(g[614]), .A2(N614), .Z(c[615]) );
  AN2D0 C7376 ( .A1(p[613]), .A2(c[613]), .Z(N613) );
  OR2D0 C7375 ( .A1(g[613]), .A2(N613), .Z(c[614]) );
  AN2D0 C7374 ( .A1(p[612]), .A2(c[612]), .Z(N612) );
  OR2D0 C7373 ( .A1(g[612]), .A2(N612), .Z(c[613]) );
  AN2D0 C7372 ( .A1(p[611]), .A2(c[611]), .Z(N611) );
  OR2D0 C7371 ( .A1(g[611]), .A2(N611), .Z(c[612]) );
  AN2D0 C7370 ( .A1(p[610]), .A2(c[610]), .Z(N610) );
  OR2D0 C7369 ( .A1(g[610]), .A2(N610), .Z(c[611]) );
  AN2D0 C7368 ( .A1(p[609]), .A2(c[609]), .Z(N609) );
  OR2D0 C7367 ( .A1(g[609]), .A2(N609), .Z(c[610]) );
  AN2D0 C7366 ( .A1(p[608]), .A2(c[608]), .Z(N608) );
  OR2D0 C7365 ( .A1(g[608]), .A2(N608), .Z(c[609]) );
  AN2D0 C7364 ( .A1(p[607]), .A2(c[607]), .Z(N607) );
  OR2D0 C7363 ( .A1(g[607]), .A2(N607), .Z(c[608]) );
  AN2D0 C7362 ( .A1(p[606]), .A2(c[606]), .Z(N606) );
  OR2D0 C7361 ( .A1(g[606]), .A2(N606), .Z(c[607]) );
  AN2D0 C7360 ( .A1(p[605]), .A2(c[605]), .Z(N605) );
  OR2D0 C7359 ( .A1(g[605]), .A2(N605), .Z(c[606]) );
  AN2D0 C7358 ( .A1(p[604]), .A2(c[604]), .Z(N604) );
  OR2D0 C7357 ( .A1(g[604]), .A2(N604), .Z(c[605]) );
  AN2D0 C7356 ( .A1(p[603]), .A2(c[603]), .Z(N603) );
  OR2D0 C7355 ( .A1(g[603]), .A2(N603), .Z(c[604]) );
  AN2D0 C7354 ( .A1(p[602]), .A2(c[602]), .Z(N602) );
  OR2D0 C7353 ( .A1(g[602]), .A2(N602), .Z(c[603]) );
  AN2D0 C7352 ( .A1(p[601]), .A2(c[601]), .Z(N601) );
  OR2D0 C7351 ( .A1(g[601]), .A2(N601), .Z(c[602]) );
  AN2D0 C7350 ( .A1(p[600]), .A2(c[600]), .Z(N600) );
  OR2D0 C7349 ( .A1(g[600]), .A2(N600), .Z(c[601]) );
  AN2D0 C7348 ( .A1(p[599]), .A2(c[599]), .Z(N599) );
  OR2D0 C7347 ( .A1(g[599]), .A2(N599), .Z(c[600]) );
  AN2D0 C7346 ( .A1(p[598]), .A2(c[598]), .Z(N598) );
  OR2D0 C7345 ( .A1(g[598]), .A2(N598), .Z(c[599]) );
  AN2D0 C7344 ( .A1(p[597]), .A2(c[597]), .Z(N597) );
  OR2D0 C7343 ( .A1(g[597]), .A2(N597), .Z(c[598]) );
  AN2D0 C7342 ( .A1(p[596]), .A2(c[596]), .Z(N596) );
  OR2D0 C7341 ( .A1(g[596]), .A2(N596), .Z(c[597]) );
  AN2D0 C7340 ( .A1(p[595]), .A2(c[595]), .Z(N595) );
  OR2D0 C7339 ( .A1(g[595]), .A2(N595), .Z(c[596]) );
  AN2D0 C7338 ( .A1(p[594]), .A2(c[594]), .Z(N594) );
  OR2D0 C7337 ( .A1(g[594]), .A2(N594), .Z(c[595]) );
  AN2D0 C7336 ( .A1(p[593]), .A2(c[593]), .Z(N593) );
  OR2D0 C7335 ( .A1(g[593]), .A2(N593), .Z(c[594]) );
  AN2D0 C7334 ( .A1(p[592]), .A2(c[592]), .Z(N592) );
  OR2D0 C7333 ( .A1(g[592]), .A2(N592), .Z(c[593]) );
  AN2D0 C7332 ( .A1(p[591]), .A2(c[591]), .Z(N591) );
  OR2D0 C7331 ( .A1(g[591]), .A2(N591), .Z(c[592]) );
  AN2D0 C7330 ( .A1(p[590]), .A2(c[590]), .Z(N590) );
  OR2D0 C7329 ( .A1(g[590]), .A2(N590), .Z(c[591]) );
  AN2D0 C7328 ( .A1(p[589]), .A2(c[589]), .Z(N589) );
  OR2D0 C7327 ( .A1(g[589]), .A2(N589), .Z(c[590]) );
  AN2D0 C7326 ( .A1(p[588]), .A2(c[588]), .Z(N588) );
  OR2D0 C7325 ( .A1(g[588]), .A2(N588), .Z(c[589]) );
  AN2D0 C7324 ( .A1(p[587]), .A2(c[587]), .Z(N587) );
  OR2D0 C7323 ( .A1(g[587]), .A2(N587), .Z(c[588]) );
  AN2D0 C7322 ( .A1(p[586]), .A2(c[586]), .Z(N586) );
  OR2D0 C7321 ( .A1(g[586]), .A2(N586), .Z(c[587]) );
  AN2D0 C7320 ( .A1(p[585]), .A2(c[585]), .Z(N585) );
  OR2D0 C7319 ( .A1(g[585]), .A2(N585), .Z(c[586]) );
  AN2D0 C7318 ( .A1(p[584]), .A2(c[584]), .Z(N584) );
  OR2D0 C7317 ( .A1(g[584]), .A2(N584), .Z(c[585]) );
  AN2D0 C7316 ( .A1(p[583]), .A2(c[583]), .Z(N583) );
  OR2D0 C7315 ( .A1(g[583]), .A2(N583), .Z(c[584]) );
  AN2D0 C7314 ( .A1(p[582]), .A2(c[582]), .Z(N582) );
  OR2D0 C7313 ( .A1(g[582]), .A2(N582), .Z(c[583]) );
  AN2D0 C7312 ( .A1(p[581]), .A2(c[581]), .Z(N581) );
  OR2D0 C7311 ( .A1(g[581]), .A2(N581), .Z(c[582]) );
  AN2D0 C7310 ( .A1(p[580]), .A2(c[580]), .Z(N580) );
  OR2D0 C7309 ( .A1(g[580]), .A2(N580), .Z(c[581]) );
  AN2D0 C7308 ( .A1(p[579]), .A2(c[579]), .Z(N579) );
  OR2D0 C7307 ( .A1(g[579]), .A2(N579), .Z(c[580]) );
  AN2D0 C7306 ( .A1(p[578]), .A2(c[578]), .Z(N578) );
  OR2D0 C7305 ( .A1(g[578]), .A2(N578), .Z(c[579]) );
  AN2D0 C7304 ( .A1(p[577]), .A2(c[577]), .Z(N577) );
  OR2D0 C7303 ( .A1(g[577]), .A2(N577), .Z(c[578]) );
  AN2D0 C7302 ( .A1(p[576]), .A2(c[576]), .Z(N576) );
  OR2D0 C7301 ( .A1(g[576]), .A2(N576), .Z(c[577]) );
  AN2D0 C7300 ( .A1(p[575]), .A2(c[575]), .Z(N575) );
  OR2D0 C7299 ( .A1(g[575]), .A2(N575), .Z(c[576]) );
  AN2D0 C7298 ( .A1(p[574]), .A2(c[574]), .Z(N574) );
  OR2D0 C7297 ( .A1(g[574]), .A2(N574), .Z(c[575]) );
  AN2D0 C7296 ( .A1(p[573]), .A2(c[573]), .Z(N573) );
  OR2D0 C7295 ( .A1(g[573]), .A2(N573), .Z(c[574]) );
  AN2D0 C7294 ( .A1(p[572]), .A2(c[572]), .Z(N572) );
  OR2D0 C7293 ( .A1(g[572]), .A2(N572), .Z(c[573]) );
  AN2D0 C7292 ( .A1(p[571]), .A2(c[571]), .Z(N571) );
  OR2D0 C7291 ( .A1(g[571]), .A2(N571), .Z(c[572]) );
  AN2D0 C7290 ( .A1(p[570]), .A2(c[570]), .Z(N570) );
  OR2D0 C7289 ( .A1(g[570]), .A2(N570), .Z(c[571]) );
  AN2D0 C7288 ( .A1(p[569]), .A2(c[569]), .Z(N569) );
  OR2D0 C7287 ( .A1(g[569]), .A2(N569), .Z(c[570]) );
  AN2D0 C7286 ( .A1(p[568]), .A2(c[568]), .Z(N568) );
  OR2D0 C7285 ( .A1(g[568]), .A2(N568), .Z(c[569]) );
  AN2D0 C7284 ( .A1(p[567]), .A2(c[567]), .Z(N567) );
  OR2D0 C7283 ( .A1(g[567]), .A2(N567), .Z(c[568]) );
  AN2D0 C7282 ( .A1(p[566]), .A2(c[566]), .Z(N566) );
  OR2D0 C7281 ( .A1(g[566]), .A2(N566), .Z(c[567]) );
  AN2D0 C7280 ( .A1(p[565]), .A2(c[565]), .Z(N565) );
  OR2D0 C7279 ( .A1(g[565]), .A2(N565), .Z(c[566]) );
  AN2D0 C7278 ( .A1(p[564]), .A2(c[564]), .Z(N564) );
  OR2D0 C7277 ( .A1(g[564]), .A2(N564), .Z(c[565]) );
  AN2D0 C7276 ( .A1(p[563]), .A2(c[563]), .Z(N563) );
  OR2D0 C7275 ( .A1(g[563]), .A2(N563), .Z(c[564]) );
  AN2D0 C7274 ( .A1(p[562]), .A2(c[562]), .Z(N562) );
  OR2D0 C7273 ( .A1(g[562]), .A2(N562), .Z(c[563]) );
  AN2D0 C7272 ( .A1(p[561]), .A2(c[561]), .Z(N561) );
  OR2D0 C7271 ( .A1(g[561]), .A2(N561), .Z(c[562]) );
  AN2D0 C7270 ( .A1(p[560]), .A2(c[560]), .Z(N560) );
  OR2D0 C7269 ( .A1(g[560]), .A2(N560), .Z(c[561]) );
  AN2D0 C7268 ( .A1(p[559]), .A2(c[559]), .Z(N559) );
  OR2D0 C7267 ( .A1(g[559]), .A2(N559), .Z(c[560]) );
  AN2D0 C7266 ( .A1(p[558]), .A2(c[558]), .Z(N558) );
  OR2D0 C7265 ( .A1(g[558]), .A2(N558), .Z(c[559]) );
  AN2D0 C7264 ( .A1(p[557]), .A2(c[557]), .Z(N557) );
  OR2D0 C7263 ( .A1(g[557]), .A2(N557), .Z(c[558]) );
  AN2D0 C7262 ( .A1(p[556]), .A2(c[556]), .Z(N556) );
  OR2D0 C7261 ( .A1(g[556]), .A2(N556), .Z(c[557]) );
  AN2D0 C7260 ( .A1(p[555]), .A2(c[555]), .Z(N555) );
  OR2D0 C7259 ( .A1(g[555]), .A2(N555), .Z(c[556]) );
  AN2D0 C7258 ( .A1(p[554]), .A2(c[554]), .Z(N554) );
  OR2D0 C7257 ( .A1(g[554]), .A2(N554), .Z(c[555]) );
  AN2D0 C7256 ( .A1(p[553]), .A2(c[553]), .Z(N553) );
  OR2D0 C7255 ( .A1(g[553]), .A2(N553), .Z(c[554]) );
  AN2D0 C7254 ( .A1(p[552]), .A2(c[552]), .Z(N552) );
  OR2D0 C7253 ( .A1(g[552]), .A2(N552), .Z(c[553]) );
  AN2D0 C7252 ( .A1(p[551]), .A2(c[551]), .Z(N551) );
  OR2D0 C7251 ( .A1(g[551]), .A2(N551), .Z(c[552]) );
  AN2D0 C7250 ( .A1(p[550]), .A2(c[550]), .Z(N550) );
  OR2D0 C7249 ( .A1(g[550]), .A2(N550), .Z(c[551]) );
  AN2D0 C7248 ( .A1(p[549]), .A2(c[549]), .Z(N549) );
  OR2D0 C7247 ( .A1(g[549]), .A2(N549), .Z(c[550]) );
  AN2D0 C7246 ( .A1(p[548]), .A2(c[548]), .Z(N548) );
  OR2D0 C7245 ( .A1(g[548]), .A2(N548), .Z(c[549]) );
  AN2D0 C7244 ( .A1(p[547]), .A2(c[547]), .Z(N547) );
  OR2D0 C7243 ( .A1(g[547]), .A2(N547), .Z(c[548]) );
  AN2D0 C7242 ( .A1(p[546]), .A2(c[546]), .Z(N546) );
  OR2D0 C7241 ( .A1(g[546]), .A2(N546), .Z(c[547]) );
  AN2D0 C7240 ( .A1(p[545]), .A2(c[545]), .Z(N545) );
  OR2D0 C7239 ( .A1(g[545]), .A2(N545), .Z(c[546]) );
  AN2D0 C7238 ( .A1(p[544]), .A2(c[544]), .Z(N544) );
  OR2D0 C7237 ( .A1(g[544]), .A2(N544), .Z(c[545]) );
  AN2D0 C7236 ( .A1(p[543]), .A2(c[543]), .Z(N543) );
  OR2D0 C7235 ( .A1(g[543]), .A2(N543), .Z(c[544]) );
  AN2D0 C7234 ( .A1(p[542]), .A2(c[542]), .Z(N542) );
  OR2D0 C7233 ( .A1(g[542]), .A2(N542), .Z(c[543]) );
  AN2D0 C7232 ( .A1(p[541]), .A2(c[541]), .Z(N541) );
  OR2D0 C7231 ( .A1(g[541]), .A2(N541), .Z(c[542]) );
  AN2D0 C7230 ( .A1(p[540]), .A2(c[540]), .Z(N540) );
  OR2D0 C7229 ( .A1(g[540]), .A2(N540), .Z(c[541]) );
  AN2D0 C7228 ( .A1(p[539]), .A2(c[539]), .Z(N539) );
  OR2D0 C7227 ( .A1(g[539]), .A2(N539), .Z(c[540]) );
  AN2D0 C7226 ( .A1(p[538]), .A2(c[538]), .Z(N538) );
  OR2D0 C7225 ( .A1(g[538]), .A2(N538), .Z(c[539]) );
  AN2D0 C7224 ( .A1(p[537]), .A2(c[537]), .Z(N537) );
  OR2D0 C7223 ( .A1(g[537]), .A2(N537), .Z(c[538]) );
  AN2D0 C7222 ( .A1(p[536]), .A2(c[536]), .Z(N536) );
  OR2D0 C7221 ( .A1(g[536]), .A2(N536), .Z(c[537]) );
  AN2D0 C7220 ( .A1(p[535]), .A2(c[535]), .Z(N535) );
  OR2D0 C7219 ( .A1(g[535]), .A2(N535), .Z(c[536]) );
  AN2D0 C7218 ( .A1(p[534]), .A2(c[534]), .Z(N534) );
  OR2D0 C7217 ( .A1(g[534]), .A2(N534), .Z(c[535]) );
  AN2D0 C7216 ( .A1(p[533]), .A2(c[533]), .Z(N533) );
  OR2D0 C7215 ( .A1(g[533]), .A2(N533), .Z(c[534]) );
  AN2D0 C7214 ( .A1(p[532]), .A2(c[532]), .Z(N532) );
  OR2D0 C7213 ( .A1(g[532]), .A2(N532), .Z(c[533]) );
  AN2D0 C7212 ( .A1(p[531]), .A2(c[531]), .Z(N531) );
  OR2D0 C7211 ( .A1(g[531]), .A2(N531), .Z(c[532]) );
  AN2D0 C7210 ( .A1(p[530]), .A2(c[530]), .Z(N530) );
  OR2D0 C7209 ( .A1(g[530]), .A2(N530), .Z(c[531]) );
  AN2D0 C7208 ( .A1(p[529]), .A2(c[529]), .Z(N529) );
  OR2D0 C7207 ( .A1(g[529]), .A2(N529), .Z(c[530]) );
  AN2D0 C7206 ( .A1(p[528]), .A2(c[528]), .Z(N528) );
  OR2D0 C7205 ( .A1(g[528]), .A2(N528), .Z(c[529]) );
  AN2D0 C7204 ( .A1(p[527]), .A2(c[527]), .Z(N527) );
  OR2D0 C7203 ( .A1(g[527]), .A2(N527), .Z(c[528]) );
  AN2D0 C7202 ( .A1(p[526]), .A2(c[526]), .Z(N526) );
  OR2D0 C7201 ( .A1(g[526]), .A2(N526), .Z(c[527]) );
  AN2D0 C7200 ( .A1(p[525]), .A2(c[525]), .Z(N525) );
  OR2D0 C7199 ( .A1(g[525]), .A2(N525), .Z(c[526]) );
  AN2D0 C7198 ( .A1(p[524]), .A2(c[524]), .Z(N524) );
  OR2D0 C7197 ( .A1(g[524]), .A2(N524), .Z(c[525]) );
  AN2D0 C7196 ( .A1(p[523]), .A2(c[523]), .Z(N523) );
  OR2D0 C7195 ( .A1(g[523]), .A2(N523), .Z(c[524]) );
  AN2D0 C7194 ( .A1(p[522]), .A2(c[522]), .Z(N522) );
  OR2D0 C7193 ( .A1(g[522]), .A2(N522), .Z(c[523]) );
  AN2D0 C7192 ( .A1(p[521]), .A2(c[521]), .Z(N521) );
  OR2D0 C7191 ( .A1(g[521]), .A2(N521), .Z(c[522]) );
  AN2D0 C7190 ( .A1(p[520]), .A2(c[520]), .Z(N520) );
  OR2D0 C7189 ( .A1(g[520]), .A2(N520), .Z(c[521]) );
  AN2D0 C7188 ( .A1(p[519]), .A2(c[519]), .Z(N519) );
  OR2D0 C7187 ( .A1(g[519]), .A2(N519), .Z(c[520]) );
  AN2D0 C7186 ( .A1(p[518]), .A2(c[518]), .Z(N518) );
  OR2D0 C7185 ( .A1(g[518]), .A2(N518), .Z(c[519]) );
  AN2D0 C7184 ( .A1(p[517]), .A2(c[517]), .Z(N517) );
  OR2D0 C7183 ( .A1(g[517]), .A2(N517), .Z(c[518]) );
  AN2D0 C7182 ( .A1(p[516]), .A2(c[516]), .Z(N516) );
  OR2D0 C7181 ( .A1(g[516]), .A2(N516), .Z(c[517]) );
  AN2D0 C7180 ( .A1(p[515]), .A2(c[515]), .Z(N515) );
  OR2D0 C7179 ( .A1(g[515]), .A2(N515), .Z(c[516]) );
  AN2D0 C7178 ( .A1(p[514]), .A2(c[514]), .Z(N514) );
  OR2D0 C7177 ( .A1(g[514]), .A2(N514), .Z(c[515]) );
  AN2D0 C7176 ( .A1(p[513]), .A2(c[513]), .Z(N513) );
  OR2D0 C7175 ( .A1(g[513]), .A2(N513), .Z(c[514]) );
  AN2D0 C7174 ( .A1(p[512]), .A2(c[512]), .Z(N512) );
  OR2D0 C7173 ( .A1(g[512]), .A2(N512), .Z(c[513]) );
  AN2D0 C7172 ( .A1(p[511]), .A2(c[511]), .Z(N511) );
  OR2D0 C7171 ( .A1(g[511]), .A2(N511), .Z(c[512]) );
  AN2D0 C7170 ( .A1(p[510]), .A2(c[510]), .Z(N510) );
  OR2D0 C7169 ( .A1(g[510]), .A2(N510), .Z(c[511]) );
  AN2D0 C7168 ( .A1(p[509]), .A2(c[509]), .Z(N509) );
  OR2D0 C7167 ( .A1(g[509]), .A2(N509), .Z(c[510]) );
  AN2D0 C7166 ( .A1(p[508]), .A2(c[508]), .Z(N508) );
  OR2D0 C7165 ( .A1(g[508]), .A2(N508), .Z(c[509]) );
  AN2D0 C7164 ( .A1(p[507]), .A2(c[507]), .Z(N507) );
  OR2D0 C7163 ( .A1(g[507]), .A2(N507), .Z(c[508]) );
  AN2D0 C7162 ( .A1(p[506]), .A2(c[506]), .Z(N506) );
  OR2D0 C7161 ( .A1(g[506]), .A2(N506), .Z(c[507]) );
  AN2D0 C7160 ( .A1(p[505]), .A2(c[505]), .Z(N505) );
  OR2D0 C7159 ( .A1(g[505]), .A2(N505), .Z(c[506]) );
  AN2D0 C7158 ( .A1(p[504]), .A2(c[504]), .Z(N504) );
  OR2D0 C7157 ( .A1(g[504]), .A2(N504), .Z(c[505]) );
  AN2D0 C7156 ( .A1(p[503]), .A2(c[503]), .Z(N503) );
  OR2D0 C7155 ( .A1(g[503]), .A2(N503), .Z(c[504]) );
  AN2D0 C7154 ( .A1(p[502]), .A2(c[502]), .Z(N502) );
  OR2D0 C7153 ( .A1(g[502]), .A2(N502), .Z(c[503]) );
  AN2D0 C7152 ( .A1(p[501]), .A2(c[501]), .Z(N501) );
  OR2D0 C7151 ( .A1(g[501]), .A2(N501), .Z(c[502]) );
  AN2D0 C7150 ( .A1(p[500]), .A2(c[500]), .Z(N500) );
  OR2D0 C7149 ( .A1(g[500]), .A2(N500), .Z(c[501]) );
  AN2D0 C7148 ( .A1(p[499]), .A2(c[499]), .Z(N499) );
  OR2D0 C7147 ( .A1(g[499]), .A2(N499), .Z(c[500]) );
  AN2D0 C7146 ( .A1(p[498]), .A2(c[498]), .Z(N498) );
  OR2D0 C7145 ( .A1(g[498]), .A2(N498), .Z(c[499]) );
  AN2D0 C7144 ( .A1(p[497]), .A2(c[497]), .Z(N497) );
  OR2D0 C7143 ( .A1(g[497]), .A2(N497), .Z(c[498]) );
  AN2D0 C7142 ( .A1(p[496]), .A2(c[496]), .Z(N496) );
  OR2D0 C7141 ( .A1(g[496]), .A2(N496), .Z(c[497]) );
  AN2D0 C7140 ( .A1(p[495]), .A2(c[495]), .Z(N495) );
  OR2D0 C7139 ( .A1(g[495]), .A2(N495), .Z(c[496]) );
  AN2D0 C7138 ( .A1(p[494]), .A2(c[494]), .Z(N494) );
  OR2D0 C7137 ( .A1(g[494]), .A2(N494), .Z(c[495]) );
  AN2D0 C7136 ( .A1(p[493]), .A2(c[493]), .Z(N493) );
  OR2D0 C7135 ( .A1(g[493]), .A2(N493), .Z(c[494]) );
  AN2D0 C7134 ( .A1(p[492]), .A2(c[492]), .Z(N492) );
  OR2D0 C7133 ( .A1(g[492]), .A2(N492), .Z(c[493]) );
  AN2D0 C7132 ( .A1(p[491]), .A2(c[491]), .Z(N491) );
  OR2D0 C7131 ( .A1(g[491]), .A2(N491), .Z(c[492]) );
  AN2D0 C7130 ( .A1(p[490]), .A2(c[490]), .Z(N490) );
  OR2D0 C7129 ( .A1(g[490]), .A2(N490), .Z(c[491]) );
  AN2D0 C7128 ( .A1(p[489]), .A2(c[489]), .Z(N489) );
  OR2D0 C7127 ( .A1(g[489]), .A2(N489), .Z(c[490]) );
  AN2D0 C7126 ( .A1(p[488]), .A2(c[488]), .Z(N488) );
  OR2D0 C7125 ( .A1(g[488]), .A2(N488), .Z(c[489]) );
  AN2D0 C7124 ( .A1(p[487]), .A2(c[487]), .Z(N487) );
  OR2D0 C7123 ( .A1(g[487]), .A2(N487), .Z(c[488]) );
  AN2D0 C7122 ( .A1(p[486]), .A2(c[486]), .Z(N486) );
  OR2D0 C7121 ( .A1(g[486]), .A2(N486), .Z(c[487]) );
  AN2D0 C7120 ( .A1(p[485]), .A2(c[485]), .Z(N485) );
  OR2D0 C7119 ( .A1(g[485]), .A2(N485), .Z(c[486]) );
  AN2D0 C7118 ( .A1(p[484]), .A2(c[484]), .Z(N484) );
  OR2D0 C7117 ( .A1(g[484]), .A2(N484), .Z(c[485]) );
  AN2D0 C7116 ( .A1(p[483]), .A2(c[483]), .Z(N483) );
  OR2D0 C7115 ( .A1(g[483]), .A2(N483), .Z(c[484]) );
  AN2D0 C7114 ( .A1(p[482]), .A2(c[482]), .Z(N482) );
  OR2D0 C7113 ( .A1(g[482]), .A2(N482), .Z(c[483]) );
  AN2D0 C7112 ( .A1(p[481]), .A2(c[481]), .Z(N481) );
  OR2D0 C7111 ( .A1(g[481]), .A2(N481), .Z(c[482]) );
  AN2D0 C7110 ( .A1(p[480]), .A2(c[480]), .Z(N480) );
  OR2D0 C7109 ( .A1(g[480]), .A2(N480), .Z(c[481]) );
  AN2D0 C7108 ( .A1(p[479]), .A2(c[479]), .Z(N479) );
  OR2D0 C7107 ( .A1(g[479]), .A2(N479), .Z(c[480]) );
  AN2D0 C7106 ( .A1(p[478]), .A2(c[478]), .Z(N478) );
  OR2D0 C7105 ( .A1(g[478]), .A2(N478), .Z(c[479]) );
  AN2D0 C7104 ( .A1(p[477]), .A2(c[477]), .Z(N477) );
  OR2D0 C7103 ( .A1(g[477]), .A2(N477), .Z(c[478]) );
  AN2D0 C7102 ( .A1(p[476]), .A2(c[476]), .Z(N476) );
  OR2D0 C7101 ( .A1(g[476]), .A2(N476), .Z(c[477]) );
  AN2D0 C7100 ( .A1(p[475]), .A2(c[475]), .Z(N475) );
  OR2D0 C7099 ( .A1(g[475]), .A2(N475), .Z(c[476]) );
  AN2D0 C7098 ( .A1(p[474]), .A2(c[474]), .Z(N474) );
  OR2D0 C7097 ( .A1(g[474]), .A2(N474), .Z(c[475]) );
  AN2D0 C7096 ( .A1(p[473]), .A2(c[473]), .Z(N473) );
  OR2D0 C7095 ( .A1(g[473]), .A2(N473), .Z(c[474]) );
  AN2D0 C7094 ( .A1(p[472]), .A2(c[472]), .Z(N472) );
  OR2D0 C7093 ( .A1(g[472]), .A2(N472), .Z(c[473]) );
  AN2D0 C7092 ( .A1(p[471]), .A2(c[471]), .Z(N471) );
  OR2D0 C7091 ( .A1(g[471]), .A2(N471), .Z(c[472]) );
  AN2D0 C7090 ( .A1(p[470]), .A2(c[470]), .Z(N470) );
  OR2D0 C7089 ( .A1(g[470]), .A2(N470), .Z(c[471]) );
  AN2D0 C7088 ( .A1(p[469]), .A2(c[469]), .Z(N469) );
  OR2D0 C7087 ( .A1(g[469]), .A2(N469), .Z(c[470]) );
  AN2D0 C7086 ( .A1(p[468]), .A2(c[468]), .Z(N468) );
  OR2D0 C7085 ( .A1(g[468]), .A2(N468), .Z(c[469]) );
  AN2D0 C7084 ( .A1(p[467]), .A2(c[467]), .Z(N467) );
  OR2D0 C7083 ( .A1(g[467]), .A2(N467), .Z(c[468]) );
  AN2D0 C7082 ( .A1(p[466]), .A2(c[466]), .Z(N466) );
  OR2D0 C7081 ( .A1(g[466]), .A2(N466), .Z(c[467]) );
  AN2D0 C7080 ( .A1(p[465]), .A2(c[465]), .Z(N465) );
  OR2D0 C7079 ( .A1(g[465]), .A2(N465), .Z(c[466]) );
  AN2D0 C7078 ( .A1(p[464]), .A2(c[464]), .Z(N464) );
  OR2D0 C7077 ( .A1(g[464]), .A2(N464), .Z(c[465]) );
  AN2D0 C7076 ( .A1(p[463]), .A2(c[463]), .Z(N463) );
  OR2D0 C7075 ( .A1(g[463]), .A2(N463), .Z(c[464]) );
  AN2D0 C7074 ( .A1(p[462]), .A2(c[462]), .Z(N462) );
  OR2D0 C7073 ( .A1(g[462]), .A2(N462), .Z(c[463]) );
  AN2D0 C7072 ( .A1(p[461]), .A2(c[461]), .Z(N461) );
  OR2D0 C7071 ( .A1(g[461]), .A2(N461), .Z(c[462]) );
  AN2D0 C7070 ( .A1(p[460]), .A2(c[460]), .Z(N460) );
  OR2D0 C7069 ( .A1(g[460]), .A2(N460), .Z(c[461]) );
  AN2D0 C7068 ( .A1(p[459]), .A2(c[459]), .Z(N459) );
  OR2D0 C7067 ( .A1(g[459]), .A2(N459), .Z(c[460]) );
  AN2D0 C7066 ( .A1(p[458]), .A2(c[458]), .Z(N458) );
  OR2D0 C7065 ( .A1(g[458]), .A2(N458), .Z(c[459]) );
  AN2D0 C7064 ( .A1(p[457]), .A2(c[457]), .Z(N457) );
  OR2D0 C7063 ( .A1(g[457]), .A2(N457), .Z(c[458]) );
  AN2D0 C7062 ( .A1(p[456]), .A2(c[456]), .Z(N456) );
  OR2D0 C7061 ( .A1(g[456]), .A2(N456), .Z(c[457]) );
  AN2D0 C7060 ( .A1(p[455]), .A2(c[455]), .Z(N455) );
  OR2D0 C7059 ( .A1(g[455]), .A2(N455), .Z(c[456]) );
  AN2D0 C7058 ( .A1(p[454]), .A2(c[454]), .Z(N454) );
  OR2D0 C7057 ( .A1(g[454]), .A2(N454), .Z(c[455]) );
  AN2D0 C7056 ( .A1(p[453]), .A2(c[453]), .Z(N453) );
  OR2D0 C7055 ( .A1(g[453]), .A2(N453), .Z(c[454]) );
  AN2D0 C7054 ( .A1(p[452]), .A2(c[452]), .Z(N452) );
  OR2D0 C7053 ( .A1(g[452]), .A2(N452), .Z(c[453]) );
  AN2D0 C7052 ( .A1(p[451]), .A2(c[451]), .Z(N451) );
  OR2D0 C7051 ( .A1(g[451]), .A2(N451), .Z(c[452]) );
  AN2D0 C7050 ( .A1(p[450]), .A2(c[450]), .Z(N450) );
  OR2D0 C7049 ( .A1(g[450]), .A2(N450), .Z(c[451]) );
  AN2D0 C7048 ( .A1(p[449]), .A2(c[449]), .Z(N449) );
  OR2D0 C7047 ( .A1(g[449]), .A2(N449), .Z(c[450]) );
  AN2D0 C7046 ( .A1(p[448]), .A2(c[448]), .Z(N448) );
  OR2D0 C7045 ( .A1(g[448]), .A2(N448), .Z(c[449]) );
  AN2D0 C7044 ( .A1(p[447]), .A2(c[447]), .Z(N447) );
  OR2D0 C7043 ( .A1(g[447]), .A2(N447), .Z(c[448]) );
  AN2D0 C7042 ( .A1(p[446]), .A2(c[446]), .Z(N446) );
  OR2D0 C7041 ( .A1(g[446]), .A2(N446), .Z(c[447]) );
  AN2D0 C7040 ( .A1(p[445]), .A2(c[445]), .Z(N445) );
  OR2D0 C7039 ( .A1(g[445]), .A2(N445), .Z(c[446]) );
  AN2D0 C7038 ( .A1(p[444]), .A2(c[444]), .Z(N444) );
  OR2D0 C7037 ( .A1(g[444]), .A2(N444), .Z(c[445]) );
  AN2D0 C7036 ( .A1(p[443]), .A2(c[443]), .Z(N443) );
  OR2D0 C7035 ( .A1(g[443]), .A2(N443), .Z(c[444]) );
  AN2D0 C7034 ( .A1(p[442]), .A2(c[442]), .Z(N442) );
  OR2D0 C7033 ( .A1(g[442]), .A2(N442), .Z(c[443]) );
  AN2D0 C7032 ( .A1(p[441]), .A2(c[441]), .Z(N441) );
  OR2D0 C7031 ( .A1(g[441]), .A2(N441), .Z(c[442]) );
  AN2D0 C7030 ( .A1(p[440]), .A2(c[440]), .Z(N440) );
  OR2D0 C7029 ( .A1(g[440]), .A2(N440), .Z(c[441]) );
  AN2D0 C7028 ( .A1(p[439]), .A2(c[439]), .Z(N439) );
  OR2D0 C7027 ( .A1(g[439]), .A2(N439), .Z(c[440]) );
  AN2D0 C7026 ( .A1(p[438]), .A2(c[438]), .Z(N438) );
  OR2D0 C7025 ( .A1(g[438]), .A2(N438), .Z(c[439]) );
  AN2D0 C7024 ( .A1(p[437]), .A2(c[437]), .Z(N437) );
  OR2D0 C7023 ( .A1(g[437]), .A2(N437), .Z(c[438]) );
  AN2D0 C7022 ( .A1(p[436]), .A2(c[436]), .Z(N436) );
  OR2D0 C7021 ( .A1(g[436]), .A2(N436), .Z(c[437]) );
  AN2D0 C7020 ( .A1(p[435]), .A2(c[435]), .Z(N435) );
  OR2D0 C7019 ( .A1(g[435]), .A2(N435), .Z(c[436]) );
  AN2D0 C7018 ( .A1(p[434]), .A2(c[434]), .Z(N434) );
  OR2D0 C7017 ( .A1(g[434]), .A2(N434), .Z(c[435]) );
  AN2D0 C7016 ( .A1(p[433]), .A2(c[433]), .Z(N433) );
  OR2D0 C7015 ( .A1(g[433]), .A2(N433), .Z(c[434]) );
  AN2D0 C7014 ( .A1(p[432]), .A2(c[432]), .Z(N432) );
  OR2D0 C7013 ( .A1(g[432]), .A2(N432), .Z(c[433]) );
  AN2D0 C7012 ( .A1(p[431]), .A2(c[431]), .Z(N431) );
  OR2D0 C7011 ( .A1(g[431]), .A2(N431), .Z(c[432]) );
  AN2D0 C7010 ( .A1(p[430]), .A2(c[430]), .Z(N430) );
  OR2D0 C7009 ( .A1(g[430]), .A2(N430), .Z(c[431]) );
  AN2D0 C7008 ( .A1(p[429]), .A2(c[429]), .Z(N429) );
  OR2D0 C7007 ( .A1(g[429]), .A2(N429), .Z(c[430]) );
  AN2D0 C7006 ( .A1(p[428]), .A2(c[428]), .Z(N428) );
  OR2D0 C7005 ( .A1(g[428]), .A2(N428), .Z(c[429]) );
  AN2D0 C7004 ( .A1(p[427]), .A2(c[427]), .Z(N427) );
  OR2D0 C7003 ( .A1(g[427]), .A2(N427), .Z(c[428]) );
  AN2D0 C7002 ( .A1(p[426]), .A2(c[426]), .Z(N426) );
  OR2D0 C7001 ( .A1(g[426]), .A2(N426), .Z(c[427]) );
  AN2D0 C7000 ( .A1(p[425]), .A2(c[425]), .Z(N425) );
  OR2D0 C6999 ( .A1(g[425]), .A2(N425), .Z(c[426]) );
  AN2D0 C6998 ( .A1(p[424]), .A2(c[424]), .Z(N424) );
  OR2D0 C6997 ( .A1(g[424]), .A2(N424), .Z(c[425]) );
  AN2D0 C6996 ( .A1(p[423]), .A2(c[423]), .Z(N423) );
  OR2D0 C6995 ( .A1(g[423]), .A2(N423), .Z(c[424]) );
  AN2D0 C6994 ( .A1(p[422]), .A2(c[422]), .Z(N422) );
  OR2D0 C6993 ( .A1(g[422]), .A2(N422), .Z(c[423]) );
  AN2D0 C6992 ( .A1(p[421]), .A2(c[421]), .Z(N421) );
  OR2D0 C6991 ( .A1(g[421]), .A2(N421), .Z(c[422]) );
  AN2D0 C6990 ( .A1(p[420]), .A2(c[420]), .Z(N420) );
  OR2D0 C6989 ( .A1(g[420]), .A2(N420), .Z(c[421]) );
  AN2D0 C6988 ( .A1(p[419]), .A2(c[419]), .Z(N419) );
  OR2D0 C6987 ( .A1(g[419]), .A2(N419), .Z(c[420]) );
  AN2D0 C6986 ( .A1(p[418]), .A2(c[418]), .Z(N418) );
  OR2D0 C6985 ( .A1(g[418]), .A2(N418), .Z(c[419]) );
  AN2D0 C6984 ( .A1(p[417]), .A2(c[417]), .Z(N417) );
  OR2D0 C6983 ( .A1(g[417]), .A2(N417), .Z(c[418]) );
  AN2D0 C6982 ( .A1(p[416]), .A2(c[416]), .Z(N416) );
  OR2D0 C6981 ( .A1(g[416]), .A2(N416), .Z(c[417]) );
  AN2D0 C6980 ( .A1(p[415]), .A2(c[415]), .Z(N415) );
  OR2D0 C6979 ( .A1(g[415]), .A2(N415), .Z(c[416]) );
  AN2D0 C6978 ( .A1(p[414]), .A2(c[414]), .Z(N414) );
  OR2D0 C6977 ( .A1(g[414]), .A2(N414), .Z(c[415]) );
  AN2D0 C6976 ( .A1(p[413]), .A2(c[413]), .Z(N413) );
  OR2D0 C6975 ( .A1(g[413]), .A2(N413), .Z(c[414]) );
  AN2D0 C6974 ( .A1(p[412]), .A2(c[412]), .Z(N412) );
  OR2D0 C6973 ( .A1(g[412]), .A2(N412), .Z(c[413]) );
  AN2D0 C6972 ( .A1(p[411]), .A2(c[411]), .Z(N411) );
  OR2D0 C6971 ( .A1(g[411]), .A2(N411), .Z(c[412]) );
  AN2D0 C6970 ( .A1(p[410]), .A2(c[410]), .Z(N410) );
  OR2D0 C6969 ( .A1(g[410]), .A2(N410), .Z(c[411]) );
  AN2D0 C6968 ( .A1(p[409]), .A2(c[409]), .Z(N409) );
  OR2D0 C6967 ( .A1(g[409]), .A2(N409), .Z(c[410]) );
  AN2D0 C6966 ( .A1(p[408]), .A2(c[408]), .Z(N408) );
  OR2D0 C6965 ( .A1(g[408]), .A2(N408), .Z(c[409]) );
  AN2D0 C6964 ( .A1(p[407]), .A2(c[407]), .Z(N407) );
  OR2D0 C6963 ( .A1(g[407]), .A2(N407), .Z(c[408]) );
  AN2D0 C6962 ( .A1(p[406]), .A2(c[406]), .Z(N406) );
  OR2D0 C6961 ( .A1(g[406]), .A2(N406), .Z(c[407]) );
  AN2D0 C6960 ( .A1(p[405]), .A2(c[405]), .Z(N405) );
  OR2D0 C6959 ( .A1(g[405]), .A2(N405), .Z(c[406]) );
  AN2D0 C6958 ( .A1(p[404]), .A2(c[404]), .Z(N404) );
  OR2D0 C6957 ( .A1(g[404]), .A2(N404), .Z(c[405]) );
  AN2D0 C6956 ( .A1(p[403]), .A2(c[403]), .Z(N403) );
  OR2D0 C6955 ( .A1(g[403]), .A2(N403), .Z(c[404]) );
  AN2D0 C6954 ( .A1(p[402]), .A2(c[402]), .Z(N402) );
  OR2D0 C6953 ( .A1(g[402]), .A2(N402), .Z(c[403]) );
  AN2D0 C6952 ( .A1(p[401]), .A2(c[401]), .Z(N401) );
  OR2D0 C6951 ( .A1(g[401]), .A2(N401), .Z(c[402]) );
  AN2D0 C6950 ( .A1(p[400]), .A2(c[400]), .Z(N400) );
  OR2D0 C6949 ( .A1(g[400]), .A2(N400), .Z(c[401]) );
  AN2D0 C6948 ( .A1(p[399]), .A2(c[399]), .Z(N399) );
  OR2D0 C6947 ( .A1(g[399]), .A2(N399), .Z(c[400]) );
  AN2D0 C6946 ( .A1(p[398]), .A2(c[398]), .Z(N398) );
  OR2D0 C6945 ( .A1(g[398]), .A2(N398), .Z(c[399]) );
  AN2D0 C6944 ( .A1(p[397]), .A2(c[397]), .Z(N397) );
  OR2D0 C6943 ( .A1(g[397]), .A2(N397), .Z(c[398]) );
  AN2D0 C6942 ( .A1(p[396]), .A2(c[396]), .Z(N396) );
  OR2D0 C6941 ( .A1(g[396]), .A2(N396), .Z(c[397]) );
  AN2D0 C6940 ( .A1(p[395]), .A2(c[395]), .Z(N395) );
  OR2D0 C6939 ( .A1(g[395]), .A2(N395), .Z(c[396]) );
  AN2D0 C6938 ( .A1(p[394]), .A2(c[394]), .Z(N394) );
  OR2D0 C6937 ( .A1(g[394]), .A2(N394), .Z(c[395]) );
  AN2D0 C6936 ( .A1(p[393]), .A2(c[393]), .Z(N393) );
  OR2D0 C6935 ( .A1(g[393]), .A2(N393), .Z(c[394]) );
  AN2D0 C6934 ( .A1(p[392]), .A2(c[392]), .Z(N392) );
  OR2D0 C6933 ( .A1(g[392]), .A2(N392), .Z(c[393]) );
  AN2D0 C6932 ( .A1(p[391]), .A2(c[391]), .Z(N391) );
  OR2D0 C6931 ( .A1(g[391]), .A2(N391), .Z(c[392]) );
  AN2D0 C6930 ( .A1(p[390]), .A2(c[390]), .Z(N390) );
  OR2D0 C6929 ( .A1(g[390]), .A2(N390), .Z(c[391]) );
  AN2D0 C6928 ( .A1(p[389]), .A2(c[389]), .Z(N389) );
  OR2D0 C6927 ( .A1(g[389]), .A2(N389), .Z(c[390]) );
  AN2D0 C6926 ( .A1(p[388]), .A2(c[388]), .Z(N388) );
  OR2D0 C6925 ( .A1(g[388]), .A2(N388), .Z(c[389]) );
  AN2D0 C6924 ( .A1(p[387]), .A2(c[387]), .Z(N387) );
  OR2D0 C6923 ( .A1(g[387]), .A2(N387), .Z(c[388]) );
  AN2D0 C6922 ( .A1(p[386]), .A2(c[386]), .Z(N386) );
  OR2D0 C6921 ( .A1(g[386]), .A2(N386), .Z(c[387]) );
  AN2D0 C6920 ( .A1(p[385]), .A2(c[385]), .Z(N385) );
  OR2D0 C6919 ( .A1(g[385]), .A2(N385), .Z(c[386]) );
  AN2D0 C6918 ( .A1(p[384]), .A2(c[384]), .Z(N384) );
  OR2D0 C6917 ( .A1(g[384]), .A2(N384), .Z(c[385]) );
  AN2D0 C6916 ( .A1(p[383]), .A2(c[383]), .Z(N383) );
  OR2D0 C6915 ( .A1(g[383]), .A2(N383), .Z(c[384]) );
  AN2D0 C6914 ( .A1(p[382]), .A2(c[382]), .Z(N382) );
  OR2D0 C6913 ( .A1(g[382]), .A2(N382), .Z(c[383]) );
  AN2D0 C6912 ( .A1(p[381]), .A2(c[381]), .Z(N381) );
  OR2D0 C6911 ( .A1(g[381]), .A2(N381), .Z(c[382]) );
  AN2D0 C6910 ( .A1(p[380]), .A2(c[380]), .Z(N380) );
  OR2D0 C6909 ( .A1(g[380]), .A2(N380), .Z(c[381]) );
  AN2D0 C6908 ( .A1(p[379]), .A2(c[379]), .Z(N379) );
  OR2D0 C6907 ( .A1(g[379]), .A2(N379), .Z(c[380]) );
  AN2D0 C6906 ( .A1(p[378]), .A2(c[378]), .Z(N378) );
  OR2D0 C6905 ( .A1(g[378]), .A2(N378), .Z(c[379]) );
  AN2D0 C6904 ( .A1(p[377]), .A2(c[377]), .Z(N377) );
  OR2D0 C6903 ( .A1(g[377]), .A2(N377), .Z(c[378]) );
  AN2D0 C6902 ( .A1(p[376]), .A2(c[376]), .Z(N376) );
  OR2D0 C6901 ( .A1(g[376]), .A2(N376), .Z(c[377]) );
  AN2D0 C6900 ( .A1(p[375]), .A2(c[375]), .Z(N375) );
  OR2D0 C6899 ( .A1(g[375]), .A2(N375), .Z(c[376]) );
  AN2D0 C6898 ( .A1(p[374]), .A2(c[374]), .Z(N374) );
  OR2D0 C6897 ( .A1(g[374]), .A2(N374), .Z(c[375]) );
  AN2D0 C6896 ( .A1(p[373]), .A2(c[373]), .Z(N373) );
  OR2D0 C6895 ( .A1(g[373]), .A2(N373), .Z(c[374]) );
  AN2D0 C6894 ( .A1(p[372]), .A2(c[372]), .Z(N372) );
  OR2D0 C6893 ( .A1(g[372]), .A2(N372), .Z(c[373]) );
  AN2D0 C6892 ( .A1(p[371]), .A2(c[371]), .Z(N371) );
  OR2D0 C6891 ( .A1(g[371]), .A2(N371), .Z(c[372]) );
  AN2D0 C6890 ( .A1(p[370]), .A2(c[370]), .Z(N370) );
  OR2D0 C6889 ( .A1(g[370]), .A2(N370), .Z(c[371]) );
  AN2D0 C6888 ( .A1(p[369]), .A2(c[369]), .Z(N369) );
  OR2D0 C6887 ( .A1(g[369]), .A2(N369), .Z(c[370]) );
  AN2D0 C6886 ( .A1(p[368]), .A2(c[368]), .Z(N368) );
  OR2D0 C6885 ( .A1(g[368]), .A2(N368), .Z(c[369]) );
  AN2D0 C6884 ( .A1(p[367]), .A2(c[367]), .Z(N367) );
  OR2D0 C6883 ( .A1(g[367]), .A2(N367), .Z(c[368]) );
  AN2D0 C6882 ( .A1(p[366]), .A2(c[366]), .Z(N366) );
  OR2D0 C6881 ( .A1(g[366]), .A2(N366), .Z(c[367]) );
  AN2D0 C6880 ( .A1(p[365]), .A2(c[365]), .Z(N365) );
  OR2D0 C6879 ( .A1(g[365]), .A2(N365), .Z(c[366]) );
  AN2D0 C6878 ( .A1(p[364]), .A2(c[364]), .Z(N364) );
  OR2D0 C6877 ( .A1(g[364]), .A2(N364), .Z(c[365]) );
  AN2D0 C6876 ( .A1(p[363]), .A2(c[363]), .Z(N363) );
  OR2D0 C6875 ( .A1(g[363]), .A2(N363), .Z(c[364]) );
  AN2D0 C6874 ( .A1(p[362]), .A2(c[362]), .Z(N362) );
  OR2D0 C6873 ( .A1(g[362]), .A2(N362), .Z(c[363]) );
  AN2D0 C6872 ( .A1(p[361]), .A2(c[361]), .Z(N361) );
  OR2D0 C6871 ( .A1(g[361]), .A2(N361), .Z(c[362]) );
  AN2D0 C6870 ( .A1(p[360]), .A2(c[360]), .Z(N360) );
  OR2D0 C6869 ( .A1(g[360]), .A2(N360), .Z(c[361]) );
  AN2D0 C6868 ( .A1(p[359]), .A2(c[359]), .Z(N359) );
  OR2D0 C6867 ( .A1(g[359]), .A2(N359), .Z(c[360]) );
  AN2D0 C6866 ( .A1(p[358]), .A2(c[358]), .Z(N358) );
  OR2D0 C6865 ( .A1(g[358]), .A2(N358), .Z(c[359]) );
  AN2D0 C6864 ( .A1(p[357]), .A2(c[357]), .Z(N357) );
  OR2D0 C6863 ( .A1(g[357]), .A2(N357), .Z(c[358]) );
  AN2D0 C6862 ( .A1(p[356]), .A2(c[356]), .Z(N356) );
  OR2D0 C6861 ( .A1(g[356]), .A2(N356), .Z(c[357]) );
  AN2D0 C6860 ( .A1(p[355]), .A2(c[355]), .Z(N355) );
  OR2D0 C6859 ( .A1(g[355]), .A2(N355), .Z(c[356]) );
  AN2D0 C6858 ( .A1(p[354]), .A2(c[354]), .Z(N354) );
  OR2D0 C6857 ( .A1(g[354]), .A2(N354), .Z(c[355]) );
  AN2D0 C6856 ( .A1(p[353]), .A2(c[353]), .Z(N353) );
  OR2D0 C6855 ( .A1(g[353]), .A2(N353), .Z(c[354]) );
  AN2D0 C6854 ( .A1(p[352]), .A2(c[352]), .Z(N352) );
  OR2D0 C6853 ( .A1(g[352]), .A2(N352), .Z(c[353]) );
  AN2D0 C6852 ( .A1(p[351]), .A2(c[351]), .Z(N351) );
  OR2D0 C6851 ( .A1(g[351]), .A2(N351), .Z(c[352]) );
  AN2D0 C6850 ( .A1(p[350]), .A2(c[350]), .Z(N350) );
  OR2D0 C6849 ( .A1(g[350]), .A2(N350), .Z(c[351]) );
  AN2D0 C6848 ( .A1(p[349]), .A2(c[349]), .Z(N349) );
  OR2D0 C6847 ( .A1(g[349]), .A2(N349), .Z(c[350]) );
  AN2D0 C6846 ( .A1(p[348]), .A2(c[348]), .Z(N348) );
  OR2D0 C6845 ( .A1(g[348]), .A2(N348), .Z(c[349]) );
  AN2D0 C6844 ( .A1(p[347]), .A2(c[347]), .Z(N347) );
  OR2D0 C6843 ( .A1(g[347]), .A2(N347), .Z(c[348]) );
  AN2D0 C6842 ( .A1(p[346]), .A2(c[346]), .Z(N346) );
  OR2D0 C6841 ( .A1(g[346]), .A2(N346), .Z(c[347]) );
  AN2D0 C6840 ( .A1(p[345]), .A2(c[345]), .Z(N345) );
  OR2D0 C6839 ( .A1(g[345]), .A2(N345), .Z(c[346]) );
  AN2D0 C6838 ( .A1(p[344]), .A2(c[344]), .Z(N344) );
  OR2D0 C6837 ( .A1(g[344]), .A2(N344), .Z(c[345]) );
  AN2D0 C6836 ( .A1(p[343]), .A2(c[343]), .Z(N343) );
  OR2D0 C6835 ( .A1(g[343]), .A2(N343), .Z(c[344]) );
  AN2D0 C6834 ( .A1(p[342]), .A2(c[342]), .Z(N342) );
  OR2D0 C6833 ( .A1(g[342]), .A2(N342), .Z(c[343]) );
  AN2D0 C6832 ( .A1(p[341]), .A2(c[341]), .Z(N341) );
  OR2D0 C6831 ( .A1(g[341]), .A2(N341), .Z(c[342]) );
  AN2D0 C6830 ( .A1(p[340]), .A2(c[340]), .Z(N340) );
  OR2D0 C6829 ( .A1(g[340]), .A2(N340), .Z(c[341]) );
  AN2D0 C6828 ( .A1(p[339]), .A2(c[339]), .Z(N339) );
  OR2D0 C6827 ( .A1(g[339]), .A2(N339), .Z(c[340]) );
  AN2D0 C6826 ( .A1(p[338]), .A2(c[338]), .Z(N338) );
  OR2D0 C6825 ( .A1(g[338]), .A2(N338), .Z(c[339]) );
  AN2D0 C6824 ( .A1(p[337]), .A2(c[337]), .Z(N337) );
  OR2D0 C6823 ( .A1(g[337]), .A2(N337), .Z(c[338]) );
  AN2D0 C6822 ( .A1(p[336]), .A2(c[336]), .Z(N336) );
  OR2D0 C6821 ( .A1(g[336]), .A2(N336), .Z(c[337]) );
  AN2D0 C6820 ( .A1(p[335]), .A2(c[335]), .Z(N335) );
  OR2D0 C6819 ( .A1(g[335]), .A2(N335), .Z(c[336]) );
  AN2D0 C6818 ( .A1(p[334]), .A2(c[334]), .Z(N334) );
  OR2D0 C6817 ( .A1(g[334]), .A2(N334), .Z(c[335]) );
  AN2D0 C6816 ( .A1(p[333]), .A2(c[333]), .Z(N333) );
  OR2D0 C6815 ( .A1(g[333]), .A2(N333), .Z(c[334]) );
  AN2D0 C6814 ( .A1(p[332]), .A2(c[332]), .Z(N332) );
  OR2D0 C6813 ( .A1(g[332]), .A2(N332), .Z(c[333]) );
  AN2D0 C6812 ( .A1(p[331]), .A2(c[331]), .Z(N331) );
  OR2D0 C6811 ( .A1(g[331]), .A2(N331), .Z(c[332]) );
  AN2D0 C6810 ( .A1(p[330]), .A2(c[330]), .Z(N330) );
  OR2D0 C6809 ( .A1(g[330]), .A2(N330), .Z(c[331]) );
  AN2D0 C6808 ( .A1(p[329]), .A2(c[329]), .Z(N329) );
  OR2D0 C6807 ( .A1(g[329]), .A2(N329), .Z(c[330]) );
  AN2D0 C6806 ( .A1(p[328]), .A2(c[328]), .Z(N328) );
  OR2D0 C6805 ( .A1(g[328]), .A2(N328), .Z(c[329]) );
  AN2D0 C6804 ( .A1(p[327]), .A2(c[327]), .Z(N327) );
  OR2D0 C6803 ( .A1(g[327]), .A2(N327), .Z(c[328]) );
  AN2D0 C6802 ( .A1(p[326]), .A2(c[326]), .Z(N326) );
  OR2D0 C6801 ( .A1(g[326]), .A2(N326), .Z(c[327]) );
  AN2D0 C6800 ( .A1(p[325]), .A2(c[325]), .Z(N325) );
  OR2D0 C6799 ( .A1(g[325]), .A2(N325), .Z(c[326]) );
  AN2D0 C6798 ( .A1(p[324]), .A2(c[324]), .Z(N324) );
  OR2D0 C6797 ( .A1(g[324]), .A2(N324), .Z(c[325]) );
  AN2D0 C6796 ( .A1(p[323]), .A2(c[323]), .Z(N323) );
  OR2D0 C6795 ( .A1(g[323]), .A2(N323), .Z(c[324]) );
  AN2D0 C6794 ( .A1(p[322]), .A2(c[322]), .Z(N322) );
  OR2D0 C6793 ( .A1(g[322]), .A2(N322), .Z(c[323]) );
  AN2D0 C6792 ( .A1(p[321]), .A2(c[321]), .Z(N321) );
  OR2D0 C6791 ( .A1(g[321]), .A2(N321), .Z(c[322]) );
  AN2D0 C6790 ( .A1(p[320]), .A2(c[320]), .Z(N320) );
  OR2D0 C6789 ( .A1(g[320]), .A2(N320), .Z(c[321]) );
  AN2D0 C6788 ( .A1(p[319]), .A2(c[319]), .Z(N319) );
  OR2D0 C6787 ( .A1(g[319]), .A2(N319), .Z(c[320]) );
  AN2D0 C6786 ( .A1(p[318]), .A2(c[318]), .Z(N318) );
  OR2D0 C6785 ( .A1(g[318]), .A2(N318), .Z(c[319]) );
  AN2D0 C6784 ( .A1(p[317]), .A2(c[317]), .Z(N317) );
  OR2D0 C6783 ( .A1(g[317]), .A2(N317), .Z(c[318]) );
  AN2D0 C6782 ( .A1(p[316]), .A2(c[316]), .Z(N316) );
  OR2D0 C6781 ( .A1(g[316]), .A2(N316), .Z(c[317]) );
  AN2D0 C6780 ( .A1(p[315]), .A2(c[315]), .Z(N315) );
  OR2D0 C6779 ( .A1(g[315]), .A2(N315), .Z(c[316]) );
  AN2D0 C6778 ( .A1(p[314]), .A2(c[314]), .Z(N314) );
  OR2D0 C6777 ( .A1(g[314]), .A2(N314), .Z(c[315]) );
  AN2D0 C6776 ( .A1(p[313]), .A2(c[313]), .Z(N313) );
  OR2D0 C6775 ( .A1(g[313]), .A2(N313), .Z(c[314]) );
  AN2D0 C6774 ( .A1(p[312]), .A2(c[312]), .Z(N312) );
  OR2D0 C6773 ( .A1(g[312]), .A2(N312), .Z(c[313]) );
  AN2D0 C6772 ( .A1(p[311]), .A2(c[311]), .Z(N311) );
  OR2D0 C6771 ( .A1(g[311]), .A2(N311), .Z(c[312]) );
  AN2D0 C6770 ( .A1(p[310]), .A2(c[310]), .Z(N310) );
  OR2D0 C6769 ( .A1(g[310]), .A2(N310), .Z(c[311]) );
  AN2D0 C6768 ( .A1(p[309]), .A2(c[309]), .Z(N309) );
  OR2D0 C6767 ( .A1(g[309]), .A2(N309), .Z(c[310]) );
  AN2D0 C6766 ( .A1(p[308]), .A2(c[308]), .Z(N308) );
  OR2D0 C6765 ( .A1(g[308]), .A2(N308), .Z(c[309]) );
  AN2D0 C6764 ( .A1(p[307]), .A2(c[307]), .Z(N307) );
  OR2D0 C6763 ( .A1(g[307]), .A2(N307), .Z(c[308]) );
  AN2D0 C6762 ( .A1(p[306]), .A2(c[306]), .Z(N306) );
  OR2D0 C6761 ( .A1(g[306]), .A2(N306), .Z(c[307]) );
  AN2D0 C6760 ( .A1(p[305]), .A2(c[305]), .Z(N305) );
  OR2D0 C6759 ( .A1(g[305]), .A2(N305), .Z(c[306]) );
  AN2D0 C6758 ( .A1(p[304]), .A2(c[304]), .Z(N304) );
  OR2D0 C6757 ( .A1(g[304]), .A2(N304), .Z(c[305]) );
  AN2D0 C6756 ( .A1(p[303]), .A2(c[303]), .Z(N303) );
  OR2D0 C6755 ( .A1(g[303]), .A2(N303), .Z(c[304]) );
  AN2D0 C6754 ( .A1(p[302]), .A2(c[302]), .Z(N302) );
  OR2D0 C6753 ( .A1(g[302]), .A2(N302), .Z(c[303]) );
  AN2D0 C6752 ( .A1(p[301]), .A2(c[301]), .Z(N301) );
  OR2D0 C6751 ( .A1(g[301]), .A2(N301), .Z(c[302]) );
  AN2D0 C6750 ( .A1(p[300]), .A2(c[300]), .Z(N300) );
  OR2D0 C6749 ( .A1(g[300]), .A2(N300), .Z(c[301]) );
  AN2D0 C6748 ( .A1(p[299]), .A2(c[299]), .Z(N299) );
  OR2D0 C6747 ( .A1(g[299]), .A2(N299), .Z(c[300]) );
  AN2D0 C6746 ( .A1(p[298]), .A2(c[298]), .Z(N298) );
  OR2D0 C6745 ( .A1(g[298]), .A2(N298), .Z(c[299]) );
  AN2D0 C6744 ( .A1(p[297]), .A2(c[297]), .Z(N297) );
  OR2D0 C6743 ( .A1(g[297]), .A2(N297), .Z(c[298]) );
  AN2D0 C6742 ( .A1(p[296]), .A2(c[296]), .Z(N296) );
  OR2D0 C6741 ( .A1(g[296]), .A2(N296), .Z(c[297]) );
  AN2D0 C6740 ( .A1(p[295]), .A2(c[295]), .Z(N295) );
  OR2D0 C6739 ( .A1(g[295]), .A2(N295), .Z(c[296]) );
  AN2D0 C6738 ( .A1(p[294]), .A2(c[294]), .Z(N294) );
  OR2D0 C6737 ( .A1(g[294]), .A2(N294), .Z(c[295]) );
  AN2D0 C6736 ( .A1(p[293]), .A2(c[293]), .Z(N293) );
  OR2D0 C6735 ( .A1(g[293]), .A2(N293), .Z(c[294]) );
  AN2D0 C6734 ( .A1(p[292]), .A2(c[292]), .Z(N292) );
  OR2D0 C6733 ( .A1(g[292]), .A2(N292), .Z(c[293]) );
  AN2D0 C6732 ( .A1(p[291]), .A2(c[291]), .Z(N291) );
  OR2D0 C6731 ( .A1(g[291]), .A2(N291), .Z(c[292]) );
  AN2D0 C6730 ( .A1(p[290]), .A2(c[290]), .Z(N290) );
  OR2D0 C6729 ( .A1(g[290]), .A2(N290), .Z(c[291]) );
  AN2D0 C6728 ( .A1(p[289]), .A2(c[289]), .Z(N289) );
  OR2D0 C6727 ( .A1(g[289]), .A2(N289), .Z(c[290]) );
  AN2D0 C6726 ( .A1(p[288]), .A2(c[288]), .Z(N288) );
  OR2D0 C6725 ( .A1(g[288]), .A2(N288), .Z(c[289]) );
  AN2D0 C6724 ( .A1(p[287]), .A2(c[287]), .Z(N287) );
  OR2D0 C6723 ( .A1(g[287]), .A2(N287), .Z(c[288]) );
  AN2D0 C6722 ( .A1(p[286]), .A2(c[286]), .Z(N286) );
  OR2D0 C6721 ( .A1(g[286]), .A2(N286), .Z(c[287]) );
  AN2D0 C6720 ( .A1(p[285]), .A2(c[285]), .Z(N285) );
  OR2D0 C6719 ( .A1(g[285]), .A2(N285), .Z(c[286]) );
  AN2D0 C6718 ( .A1(p[284]), .A2(c[284]), .Z(N284) );
  OR2D0 C6717 ( .A1(g[284]), .A2(N284), .Z(c[285]) );
  AN2D0 C6716 ( .A1(p[283]), .A2(c[283]), .Z(N283) );
  OR2D0 C6715 ( .A1(g[283]), .A2(N283), .Z(c[284]) );
  AN2D0 C6714 ( .A1(p[282]), .A2(c[282]), .Z(N282) );
  OR2D0 C6713 ( .A1(g[282]), .A2(N282), .Z(c[283]) );
  AN2D0 C6712 ( .A1(p[281]), .A2(c[281]), .Z(N281) );
  OR2D0 C6711 ( .A1(g[281]), .A2(N281), .Z(c[282]) );
  AN2D0 C6710 ( .A1(p[280]), .A2(c[280]), .Z(N280) );
  OR2D0 C6709 ( .A1(g[280]), .A2(N280), .Z(c[281]) );
  AN2D0 C6708 ( .A1(p[279]), .A2(c[279]), .Z(N279) );
  OR2D0 C6707 ( .A1(g[279]), .A2(N279), .Z(c[280]) );
  AN2D0 C6706 ( .A1(p[278]), .A2(c[278]), .Z(N278) );
  OR2D0 C6705 ( .A1(g[278]), .A2(N278), .Z(c[279]) );
  AN2D0 C6704 ( .A1(p[277]), .A2(c[277]), .Z(N277) );
  OR2D0 C6703 ( .A1(g[277]), .A2(N277), .Z(c[278]) );
  AN2D0 C6702 ( .A1(p[276]), .A2(c[276]), .Z(N276) );
  OR2D0 C6701 ( .A1(g[276]), .A2(N276), .Z(c[277]) );
  AN2D0 C6700 ( .A1(p[275]), .A2(c[275]), .Z(N275) );
  OR2D0 C6699 ( .A1(g[275]), .A2(N275), .Z(c[276]) );
  AN2D0 C6698 ( .A1(p[274]), .A2(c[274]), .Z(N274) );
  OR2D0 C6697 ( .A1(g[274]), .A2(N274), .Z(c[275]) );
  AN2D0 C6696 ( .A1(p[273]), .A2(c[273]), .Z(N273) );
  OR2D0 C6695 ( .A1(g[273]), .A2(N273), .Z(c[274]) );
  AN2D0 C6694 ( .A1(p[272]), .A2(c[272]), .Z(N272) );
  OR2D0 C6693 ( .A1(g[272]), .A2(N272), .Z(c[273]) );
  AN2D0 C6692 ( .A1(p[271]), .A2(c[271]), .Z(N271) );
  OR2D0 C6691 ( .A1(g[271]), .A2(N271), .Z(c[272]) );
  AN2D0 C6690 ( .A1(p[270]), .A2(c[270]), .Z(N270) );
  OR2D0 C6689 ( .A1(g[270]), .A2(N270), .Z(c[271]) );
  AN2D0 C6688 ( .A1(p[269]), .A2(c[269]), .Z(N269) );
  OR2D0 C6687 ( .A1(g[269]), .A2(N269), .Z(c[270]) );
  AN2D0 C6686 ( .A1(p[268]), .A2(c[268]), .Z(N268) );
  OR2D0 C6685 ( .A1(g[268]), .A2(N268), .Z(c[269]) );
  AN2D0 C6684 ( .A1(p[267]), .A2(c[267]), .Z(N267) );
  OR2D0 C6683 ( .A1(g[267]), .A2(N267), .Z(c[268]) );
  AN2D0 C6682 ( .A1(p[266]), .A2(c[266]), .Z(N266) );
  OR2D0 C6681 ( .A1(g[266]), .A2(N266), .Z(c[267]) );
  AN2D0 C6680 ( .A1(p[265]), .A2(c[265]), .Z(N265) );
  OR2D0 C6679 ( .A1(g[265]), .A2(N265), .Z(c[266]) );
  AN2D0 C6678 ( .A1(p[264]), .A2(c[264]), .Z(N264) );
  OR2D0 C6677 ( .A1(g[264]), .A2(N264), .Z(c[265]) );
  AN2D0 C6676 ( .A1(p[263]), .A2(c[263]), .Z(N263) );
  OR2D0 C6675 ( .A1(g[263]), .A2(N263), .Z(c[264]) );
  AN2D0 C6674 ( .A1(p[262]), .A2(c[262]), .Z(N262) );
  OR2D0 C6673 ( .A1(g[262]), .A2(N262), .Z(c[263]) );
  AN2D0 C6672 ( .A1(p[261]), .A2(c[261]), .Z(N261) );
  OR2D0 C6671 ( .A1(g[261]), .A2(N261), .Z(c[262]) );
  AN2D0 C6670 ( .A1(p[260]), .A2(c[260]), .Z(N260) );
  OR2D0 C6669 ( .A1(g[260]), .A2(N260), .Z(c[261]) );
  AN2D0 C6668 ( .A1(p[259]), .A2(c[259]), .Z(N259) );
  OR2D0 C6667 ( .A1(g[259]), .A2(N259), .Z(c[260]) );
  AN2D0 C6666 ( .A1(p[258]), .A2(c[258]), .Z(N258) );
  OR2D0 C6665 ( .A1(g[258]), .A2(N258), .Z(c[259]) );
  AN2D0 C6664 ( .A1(p[257]), .A2(c[257]), .Z(N257) );
  OR2D0 C6663 ( .A1(g[257]), .A2(N257), .Z(c[258]) );
  AN2D0 C6662 ( .A1(p[256]), .A2(c[256]), .Z(N256) );
  OR2D0 C6661 ( .A1(g[256]), .A2(N256), .Z(c[257]) );
  AN2D0 C6660 ( .A1(p[255]), .A2(c[255]), .Z(N255) );
  OR2D0 C6659 ( .A1(g[255]), .A2(N255), .Z(c[256]) );
  AN2D0 C6658 ( .A1(p[254]), .A2(c[254]), .Z(N254) );
  OR2D0 C6657 ( .A1(g[254]), .A2(N254), .Z(c[255]) );
  AN2D0 C6656 ( .A1(p[253]), .A2(c[253]), .Z(N253) );
  OR2D0 C6655 ( .A1(g[253]), .A2(N253), .Z(c[254]) );
  AN2D0 C6654 ( .A1(p[252]), .A2(c[252]), .Z(N252) );
  OR2D0 C6653 ( .A1(g[252]), .A2(N252), .Z(c[253]) );
  AN2D0 C6652 ( .A1(p[251]), .A2(c[251]), .Z(N251) );
  OR2D0 C6651 ( .A1(g[251]), .A2(N251), .Z(c[252]) );
  AN2D0 C6650 ( .A1(p[250]), .A2(c[250]), .Z(N250) );
  OR2D0 C6649 ( .A1(g[250]), .A2(N250), .Z(c[251]) );
  AN2D0 C6648 ( .A1(p[249]), .A2(c[249]), .Z(N249) );
  OR2D0 C6647 ( .A1(g[249]), .A2(N249), .Z(c[250]) );
  AN2D0 C6646 ( .A1(p[248]), .A2(c[248]), .Z(N248) );
  OR2D0 C6645 ( .A1(g[248]), .A2(N248), .Z(c[249]) );
  AN2D0 C6644 ( .A1(p[247]), .A2(c[247]), .Z(N247) );
  OR2D0 C6643 ( .A1(g[247]), .A2(N247), .Z(c[248]) );
  AN2D0 C6642 ( .A1(p[246]), .A2(c[246]), .Z(N246) );
  OR2D0 C6641 ( .A1(g[246]), .A2(N246), .Z(c[247]) );
  AN2D0 C6640 ( .A1(p[245]), .A2(c[245]), .Z(N245) );
  OR2D0 C6639 ( .A1(g[245]), .A2(N245), .Z(c[246]) );
  AN2D0 C6638 ( .A1(p[244]), .A2(c[244]), .Z(N244) );
  OR2D0 C6637 ( .A1(g[244]), .A2(N244), .Z(c[245]) );
  AN2D0 C6636 ( .A1(p[243]), .A2(c[243]), .Z(N243) );
  OR2D0 C6635 ( .A1(g[243]), .A2(N243), .Z(c[244]) );
  AN2D0 C6634 ( .A1(p[242]), .A2(c[242]), .Z(N242) );
  OR2D0 C6633 ( .A1(g[242]), .A2(N242), .Z(c[243]) );
  AN2D0 C6632 ( .A1(p[241]), .A2(c[241]), .Z(N241) );
  OR2D0 C6631 ( .A1(g[241]), .A2(N241), .Z(c[242]) );
  AN2D0 C6630 ( .A1(p[240]), .A2(c[240]), .Z(N240) );
  OR2D0 C6629 ( .A1(g[240]), .A2(N240), .Z(c[241]) );
  AN2D0 C6628 ( .A1(p[239]), .A2(c[239]), .Z(N239) );
  OR2D0 C6627 ( .A1(g[239]), .A2(N239), .Z(c[240]) );
  AN2D0 C6626 ( .A1(p[238]), .A2(c[238]), .Z(N238) );
  OR2D0 C6625 ( .A1(g[238]), .A2(N238), .Z(c[239]) );
  AN2D0 C6624 ( .A1(p[237]), .A2(c[237]), .Z(N237) );
  OR2D0 C6623 ( .A1(g[237]), .A2(N237), .Z(c[238]) );
  AN2D0 C6622 ( .A1(p[236]), .A2(c[236]), .Z(N236) );
  OR2D0 C6621 ( .A1(g[236]), .A2(N236), .Z(c[237]) );
  AN2D0 C6620 ( .A1(p[235]), .A2(c[235]), .Z(N235) );
  OR2D0 C6619 ( .A1(g[235]), .A2(N235), .Z(c[236]) );
  AN2D0 C6618 ( .A1(p[234]), .A2(c[234]), .Z(N234) );
  OR2D0 C6617 ( .A1(g[234]), .A2(N234), .Z(c[235]) );
  AN2D0 C6616 ( .A1(p[233]), .A2(c[233]), .Z(N233) );
  OR2D0 C6615 ( .A1(g[233]), .A2(N233), .Z(c[234]) );
  AN2D0 C6614 ( .A1(p[232]), .A2(c[232]), .Z(N232) );
  OR2D0 C6613 ( .A1(g[232]), .A2(N232), .Z(c[233]) );
  AN2D0 C6612 ( .A1(p[231]), .A2(c[231]), .Z(N231) );
  OR2D0 C6611 ( .A1(g[231]), .A2(N231), .Z(c[232]) );
  AN2D0 C6610 ( .A1(p[230]), .A2(c[230]), .Z(N230) );
  OR2D0 C6609 ( .A1(g[230]), .A2(N230), .Z(c[231]) );
  AN2D0 C6608 ( .A1(p[229]), .A2(c[229]), .Z(N229) );
  OR2D0 C6607 ( .A1(g[229]), .A2(N229), .Z(c[230]) );
  AN2D0 C6606 ( .A1(p[228]), .A2(c[228]), .Z(N228) );
  OR2D0 C6605 ( .A1(g[228]), .A2(N228), .Z(c[229]) );
  AN2D0 C6604 ( .A1(p[227]), .A2(c[227]), .Z(N227) );
  OR2D0 C6603 ( .A1(g[227]), .A2(N227), .Z(c[228]) );
  AN2D0 C6602 ( .A1(p[226]), .A2(c[226]), .Z(N226) );
  OR2D0 C6601 ( .A1(g[226]), .A2(N226), .Z(c[227]) );
  AN2D0 C6600 ( .A1(p[225]), .A2(c[225]), .Z(N225) );
  OR2D0 C6599 ( .A1(g[225]), .A2(N225), .Z(c[226]) );
  AN2D0 C6598 ( .A1(p[224]), .A2(c[224]), .Z(N224) );
  OR2D0 C6597 ( .A1(g[224]), .A2(N224), .Z(c[225]) );
  AN2D0 C6596 ( .A1(p[223]), .A2(c[223]), .Z(N223) );
  OR2D0 C6595 ( .A1(g[223]), .A2(N223), .Z(c[224]) );
  AN2D0 C6594 ( .A1(p[222]), .A2(c[222]), .Z(N222) );
  OR2D0 C6593 ( .A1(g[222]), .A2(N222), .Z(c[223]) );
  AN2D0 C6592 ( .A1(p[221]), .A2(c[221]), .Z(N221) );
  OR2D0 C6591 ( .A1(g[221]), .A2(N221), .Z(c[222]) );
  AN2D0 C6590 ( .A1(p[220]), .A2(c[220]), .Z(N220) );
  OR2D0 C6589 ( .A1(g[220]), .A2(N220), .Z(c[221]) );
  AN2D0 C6588 ( .A1(p[219]), .A2(c[219]), .Z(N219) );
  OR2D0 C6587 ( .A1(g[219]), .A2(N219), .Z(c[220]) );
  AN2D0 C6586 ( .A1(p[218]), .A2(c[218]), .Z(N218) );
  OR2D0 C6585 ( .A1(g[218]), .A2(N218), .Z(c[219]) );
  AN2D0 C6584 ( .A1(p[217]), .A2(c[217]), .Z(N217) );
  OR2D0 C6583 ( .A1(g[217]), .A2(N217), .Z(c[218]) );
  AN2D0 C6582 ( .A1(p[216]), .A2(c[216]), .Z(N216) );
  OR2D0 C6581 ( .A1(g[216]), .A2(N216), .Z(c[217]) );
  AN2D0 C6580 ( .A1(p[215]), .A2(c[215]), .Z(N215) );
  OR2D0 C6579 ( .A1(g[215]), .A2(N215), .Z(c[216]) );
  AN2D0 C6578 ( .A1(p[214]), .A2(c[214]), .Z(N214) );
  OR2D0 C6577 ( .A1(g[214]), .A2(N214), .Z(c[215]) );
  AN2D0 C6576 ( .A1(p[213]), .A2(c[213]), .Z(N213) );
  OR2D0 C6575 ( .A1(g[213]), .A2(N213), .Z(c[214]) );
  AN2D0 C6574 ( .A1(p[212]), .A2(c[212]), .Z(N212) );
  OR2D0 C6573 ( .A1(g[212]), .A2(N212), .Z(c[213]) );
  AN2D0 C6572 ( .A1(p[211]), .A2(c[211]), .Z(N211) );
  OR2D0 C6571 ( .A1(g[211]), .A2(N211), .Z(c[212]) );
  AN2D0 C6570 ( .A1(p[210]), .A2(c[210]), .Z(N210) );
  OR2D0 C6569 ( .A1(g[210]), .A2(N210), .Z(c[211]) );
  AN2D0 C6568 ( .A1(p[209]), .A2(c[209]), .Z(N209) );
  OR2D0 C6567 ( .A1(g[209]), .A2(N209), .Z(c[210]) );
  AN2D0 C6566 ( .A1(p[208]), .A2(c[208]), .Z(N208) );
  OR2D0 C6565 ( .A1(g[208]), .A2(N208), .Z(c[209]) );
  AN2D0 C6564 ( .A1(p[207]), .A2(c[207]), .Z(N207) );
  OR2D0 C6563 ( .A1(g[207]), .A2(N207), .Z(c[208]) );
  AN2D0 C6562 ( .A1(p[206]), .A2(c[206]), .Z(N206) );
  OR2D0 C6561 ( .A1(g[206]), .A2(N206), .Z(c[207]) );
  AN2D0 C6560 ( .A1(p[205]), .A2(c[205]), .Z(N205) );
  OR2D0 C6559 ( .A1(g[205]), .A2(N205), .Z(c[206]) );
  AN2D0 C6558 ( .A1(p[204]), .A2(c[204]), .Z(N204) );
  OR2D0 C6557 ( .A1(g[204]), .A2(N204), .Z(c[205]) );
  AN2D0 C6556 ( .A1(p[203]), .A2(c[203]), .Z(N203) );
  OR2D0 C6555 ( .A1(g[203]), .A2(N203), .Z(c[204]) );
  AN2D0 C6554 ( .A1(p[202]), .A2(c[202]), .Z(N202) );
  OR2D0 C6553 ( .A1(g[202]), .A2(N202), .Z(c[203]) );
  AN2D0 C6552 ( .A1(p[201]), .A2(c[201]), .Z(N201) );
  OR2D0 C6551 ( .A1(g[201]), .A2(N201), .Z(c[202]) );
  AN2D0 C6550 ( .A1(p[200]), .A2(c[200]), .Z(N200) );
  OR2D0 C6549 ( .A1(g[200]), .A2(N200), .Z(c[201]) );
  AN2D0 C6548 ( .A1(p[199]), .A2(c[199]), .Z(N199) );
  OR2D0 C6547 ( .A1(g[199]), .A2(N199), .Z(c[200]) );
  AN2D0 C6546 ( .A1(p[198]), .A2(c[198]), .Z(N198) );
  OR2D0 C6545 ( .A1(g[198]), .A2(N198), .Z(c[199]) );
  AN2D0 C6544 ( .A1(p[197]), .A2(c[197]), .Z(N197) );
  OR2D0 C6543 ( .A1(g[197]), .A2(N197), .Z(c[198]) );
  AN2D0 C6542 ( .A1(p[196]), .A2(c[196]), .Z(N196) );
  OR2D0 C6541 ( .A1(g[196]), .A2(N196), .Z(c[197]) );
  AN2D0 C6540 ( .A1(p[195]), .A2(c[195]), .Z(N195) );
  OR2D0 C6539 ( .A1(g[195]), .A2(N195), .Z(c[196]) );
  AN2D0 C6538 ( .A1(p[194]), .A2(c[194]), .Z(N194) );
  OR2D0 C6537 ( .A1(g[194]), .A2(N194), .Z(c[195]) );
  AN2D0 C6536 ( .A1(p[193]), .A2(c[193]), .Z(N193) );
  OR2D0 C6535 ( .A1(g[193]), .A2(N193), .Z(c[194]) );
  AN2D0 C6534 ( .A1(p[192]), .A2(c[192]), .Z(N192) );
  OR2D0 C6533 ( .A1(g[192]), .A2(N192), .Z(c[193]) );
  AN2D0 C6532 ( .A1(p[191]), .A2(c[191]), .Z(N191) );
  OR2D0 C6531 ( .A1(g[191]), .A2(N191), .Z(c[192]) );
  AN2D0 C6530 ( .A1(p[190]), .A2(c[190]), .Z(N190) );
  OR2D0 C6529 ( .A1(g[190]), .A2(N190), .Z(c[191]) );
  AN2D0 C6528 ( .A1(p[189]), .A2(c[189]), .Z(N189) );
  OR2D0 C6527 ( .A1(g[189]), .A2(N189), .Z(c[190]) );
  AN2D0 C6526 ( .A1(p[188]), .A2(c[188]), .Z(N188) );
  OR2D0 C6525 ( .A1(g[188]), .A2(N188), .Z(c[189]) );
  AN2D0 C6524 ( .A1(p[187]), .A2(c[187]), .Z(N187) );
  OR2D0 C6523 ( .A1(g[187]), .A2(N187), .Z(c[188]) );
  AN2D0 C6522 ( .A1(p[186]), .A2(c[186]), .Z(N186) );
  OR2D0 C6521 ( .A1(g[186]), .A2(N186), .Z(c[187]) );
  AN2D0 C6520 ( .A1(p[185]), .A2(c[185]), .Z(N185) );
  OR2D0 C6519 ( .A1(g[185]), .A2(N185), .Z(c[186]) );
  AN2D0 C6518 ( .A1(p[184]), .A2(c[184]), .Z(N184) );
  OR2D0 C6517 ( .A1(g[184]), .A2(N184), .Z(c[185]) );
  AN2D0 C6516 ( .A1(p[183]), .A2(c[183]), .Z(N183) );
  OR2D0 C6515 ( .A1(g[183]), .A2(N183), .Z(c[184]) );
  AN2D0 C6514 ( .A1(p[182]), .A2(c[182]), .Z(N182) );
  OR2D0 C6513 ( .A1(g[182]), .A2(N182), .Z(c[183]) );
  AN2D0 C6512 ( .A1(p[181]), .A2(c[181]), .Z(N181) );
  OR2D0 C6511 ( .A1(g[181]), .A2(N181), .Z(c[182]) );
  AN2D0 C6510 ( .A1(p[180]), .A2(c[180]), .Z(N180) );
  OR2D0 C6509 ( .A1(g[180]), .A2(N180), .Z(c[181]) );
  AN2D0 C6508 ( .A1(p[179]), .A2(c[179]), .Z(N179) );
  OR2D0 C6507 ( .A1(g[179]), .A2(N179), .Z(c[180]) );
  AN2D0 C6506 ( .A1(p[178]), .A2(c[178]), .Z(N178) );
  OR2D0 C6505 ( .A1(g[178]), .A2(N178), .Z(c[179]) );
  AN2D0 C6504 ( .A1(p[177]), .A2(c[177]), .Z(N177) );
  OR2D0 C6503 ( .A1(g[177]), .A2(N177), .Z(c[178]) );
  AN2D0 C6502 ( .A1(p[176]), .A2(c[176]), .Z(N176) );
  OR2D0 C6501 ( .A1(g[176]), .A2(N176), .Z(c[177]) );
  AN2D0 C6500 ( .A1(p[175]), .A2(c[175]), .Z(N175) );
  OR2D0 C6499 ( .A1(g[175]), .A2(N175), .Z(c[176]) );
  AN2D0 C6498 ( .A1(p[174]), .A2(c[174]), .Z(N174) );
  OR2D0 C6497 ( .A1(g[174]), .A2(N174), .Z(c[175]) );
  AN2D0 C6496 ( .A1(p[173]), .A2(c[173]), .Z(N173) );
  OR2D0 C6495 ( .A1(g[173]), .A2(N173), .Z(c[174]) );
  AN2D0 C6494 ( .A1(p[172]), .A2(c[172]), .Z(N172) );
  OR2D0 C6493 ( .A1(g[172]), .A2(N172), .Z(c[173]) );
  AN2D0 C6492 ( .A1(p[171]), .A2(c[171]), .Z(N171) );
  OR2D0 C6491 ( .A1(g[171]), .A2(N171), .Z(c[172]) );
  AN2D0 C6490 ( .A1(p[170]), .A2(c[170]), .Z(N170) );
  OR2D0 C6489 ( .A1(g[170]), .A2(N170), .Z(c[171]) );
  AN2D0 C6488 ( .A1(p[169]), .A2(c[169]), .Z(N169) );
  OR2D0 C6487 ( .A1(g[169]), .A2(N169), .Z(c[170]) );
  AN2D0 C6486 ( .A1(p[168]), .A2(c[168]), .Z(N168) );
  OR2D0 C6485 ( .A1(g[168]), .A2(N168), .Z(c[169]) );
  AN2D0 C6484 ( .A1(p[167]), .A2(c[167]), .Z(N167) );
  OR2D0 C6483 ( .A1(g[167]), .A2(N167), .Z(c[168]) );
  AN2D0 C6482 ( .A1(p[166]), .A2(c[166]), .Z(N166) );
  OR2D0 C6481 ( .A1(g[166]), .A2(N166), .Z(c[167]) );
  AN2D0 C6480 ( .A1(p[165]), .A2(c[165]), .Z(N165) );
  OR2D0 C6479 ( .A1(g[165]), .A2(N165), .Z(c[166]) );
  AN2D0 C6478 ( .A1(p[164]), .A2(c[164]), .Z(N164) );
  OR2D0 C6477 ( .A1(g[164]), .A2(N164), .Z(c[165]) );
  AN2D0 C6476 ( .A1(p[163]), .A2(c[163]), .Z(N163) );
  OR2D0 C6475 ( .A1(g[163]), .A2(N163), .Z(c[164]) );
  AN2D0 C6474 ( .A1(p[162]), .A2(c[162]), .Z(N162) );
  OR2D0 C6473 ( .A1(g[162]), .A2(N162), .Z(c[163]) );
  AN2D0 C6472 ( .A1(p[161]), .A2(c[161]), .Z(N161) );
  OR2D0 C6471 ( .A1(g[161]), .A2(N161), .Z(c[162]) );
  AN2D0 C6470 ( .A1(p[160]), .A2(c[160]), .Z(N160) );
  OR2D0 C6469 ( .A1(g[160]), .A2(N160), .Z(c[161]) );
  AN2D0 C6468 ( .A1(p[159]), .A2(c[159]), .Z(N159) );
  OR2D0 C6467 ( .A1(g[159]), .A2(N159), .Z(c[160]) );
  AN2D0 C6466 ( .A1(p[158]), .A2(c[158]), .Z(N158) );
  OR2D0 C6465 ( .A1(g[158]), .A2(N158), .Z(c[159]) );
  AN2D0 C6464 ( .A1(p[157]), .A2(c[157]), .Z(N157) );
  OR2D0 C6463 ( .A1(g[157]), .A2(N157), .Z(c[158]) );
  AN2D0 C6462 ( .A1(p[156]), .A2(c[156]), .Z(N156) );
  OR2D0 C6461 ( .A1(g[156]), .A2(N156), .Z(c[157]) );
  AN2D0 C6460 ( .A1(p[155]), .A2(c[155]), .Z(N155) );
  OR2D0 C6459 ( .A1(g[155]), .A2(N155), .Z(c[156]) );
  AN2D0 C6458 ( .A1(p[154]), .A2(c[154]), .Z(N154) );
  OR2D0 C6457 ( .A1(g[154]), .A2(N154), .Z(c[155]) );
  AN2D0 C6456 ( .A1(p[153]), .A2(c[153]), .Z(N153) );
  OR2D0 C6455 ( .A1(g[153]), .A2(N153), .Z(c[154]) );
  AN2D0 C6454 ( .A1(p[152]), .A2(c[152]), .Z(N152) );
  OR2D0 C6453 ( .A1(g[152]), .A2(N152), .Z(c[153]) );
  AN2D0 C6452 ( .A1(p[151]), .A2(c[151]), .Z(N151) );
  OR2D0 C6451 ( .A1(g[151]), .A2(N151), .Z(c[152]) );
  AN2D0 C6450 ( .A1(p[150]), .A2(c[150]), .Z(N150) );
  OR2D0 C6449 ( .A1(g[150]), .A2(N150), .Z(c[151]) );
  AN2D0 C6448 ( .A1(p[149]), .A2(c[149]), .Z(N149) );
  OR2D0 C6447 ( .A1(g[149]), .A2(N149), .Z(c[150]) );
  AN2D0 C6446 ( .A1(p[148]), .A2(c[148]), .Z(N148) );
  OR2D0 C6445 ( .A1(g[148]), .A2(N148), .Z(c[149]) );
  AN2D0 C6444 ( .A1(p[147]), .A2(c[147]), .Z(N147) );
  OR2D0 C6443 ( .A1(g[147]), .A2(N147), .Z(c[148]) );
  AN2D0 C6442 ( .A1(p[146]), .A2(c[146]), .Z(N146) );
  OR2D0 C6441 ( .A1(g[146]), .A2(N146), .Z(c[147]) );
  AN2D0 C6440 ( .A1(p[145]), .A2(c[145]), .Z(N145) );
  OR2D0 C6439 ( .A1(g[145]), .A2(N145), .Z(c[146]) );
  AN2D0 C6438 ( .A1(p[144]), .A2(c[144]), .Z(N144) );
  OR2D0 C6437 ( .A1(g[144]), .A2(N144), .Z(c[145]) );
  AN2D0 C6436 ( .A1(p[143]), .A2(c[143]), .Z(N143) );
  OR2D0 C6435 ( .A1(g[143]), .A2(N143), .Z(c[144]) );
  AN2D0 C6434 ( .A1(p[142]), .A2(c[142]), .Z(N142) );
  OR2D0 C6433 ( .A1(g[142]), .A2(N142), .Z(c[143]) );
  AN2D0 C6432 ( .A1(p[141]), .A2(c[141]), .Z(N141) );
  OR2D0 C6431 ( .A1(g[141]), .A2(N141), .Z(c[142]) );
  AN2D0 C6430 ( .A1(p[140]), .A2(c[140]), .Z(N140) );
  OR2D0 C6429 ( .A1(g[140]), .A2(N140), .Z(c[141]) );
  AN2D0 C6428 ( .A1(p[139]), .A2(c[139]), .Z(N139) );
  OR2D0 C6427 ( .A1(g[139]), .A2(N139), .Z(c[140]) );
  AN2D0 C6426 ( .A1(p[138]), .A2(c[138]), .Z(N138) );
  OR2D0 C6425 ( .A1(g[138]), .A2(N138), .Z(c[139]) );
  AN2D0 C6424 ( .A1(p[137]), .A2(c[137]), .Z(N137) );
  OR2D0 C6423 ( .A1(g[137]), .A2(N137), .Z(c[138]) );
  AN2D0 C6422 ( .A1(p[136]), .A2(c[136]), .Z(N136) );
  OR2D0 C6421 ( .A1(g[136]), .A2(N136), .Z(c[137]) );
  AN2D0 C6420 ( .A1(p[135]), .A2(c[135]), .Z(N135) );
  OR2D0 C6419 ( .A1(g[135]), .A2(N135), .Z(c[136]) );
  AN2D0 C6418 ( .A1(p[134]), .A2(c[134]), .Z(N134) );
  OR2D0 C6417 ( .A1(g[134]), .A2(N134), .Z(c[135]) );
  AN2D0 C6416 ( .A1(p[133]), .A2(c[133]), .Z(N133) );
  OR2D0 C6415 ( .A1(g[133]), .A2(N133), .Z(c[134]) );
  AN2D0 C6414 ( .A1(p[132]), .A2(c[132]), .Z(N132) );
  OR2D0 C6413 ( .A1(g[132]), .A2(N132), .Z(c[133]) );
  AN2D0 C6412 ( .A1(p[131]), .A2(c[131]), .Z(N131) );
  OR2D0 C6411 ( .A1(g[131]), .A2(N131), .Z(c[132]) );
  AN2D0 C6410 ( .A1(p[130]), .A2(c[130]), .Z(N130) );
  OR2D0 C6409 ( .A1(g[130]), .A2(N130), .Z(c[131]) );
  AN2D0 C6408 ( .A1(p[129]), .A2(c[129]), .Z(N129) );
  OR2D0 C6407 ( .A1(g[129]), .A2(N129), .Z(c[130]) );
  AN2D0 C6406 ( .A1(p[128]), .A2(c[128]), .Z(N128) );
  OR2D0 C6405 ( .A1(g[128]), .A2(N128), .Z(c[129]) );
  AN2D0 C6404 ( .A1(p[127]), .A2(c[127]), .Z(N127) );
  OR2D0 C6403 ( .A1(g[127]), .A2(N127), .Z(c[128]) );
  AN2D0 C6402 ( .A1(p[126]), .A2(c[126]), .Z(N126) );
  OR2D0 C6401 ( .A1(g[126]), .A2(N126), .Z(c[127]) );
  AN2D0 C6400 ( .A1(p[125]), .A2(c[125]), .Z(N125) );
  OR2D0 C6399 ( .A1(g[125]), .A2(N125), .Z(c[126]) );
  AN2D0 C6398 ( .A1(p[124]), .A2(c[124]), .Z(N124) );
  OR2D0 C6397 ( .A1(g[124]), .A2(N124), .Z(c[125]) );
  AN2D0 C6396 ( .A1(p[123]), .A2(c[123]), .Z(N123) );
  OR2D0 C6395 ( .A1(g[123]), .A2(N123), .Z(c[124]) );
  AN2D0 C6394 ( .A1(p[122]), .A2(c[122]), .Z(N122) );
  OR2D0 C6393 ( .A1(g[122]), .A2(N122), .Z(c[123]) );
  AN2D0 C6392 ( .A1(p[121]), .A2(c[121]), .Z(N121) );
  OR2D0 C6391 ( .A1(g[121]), .A2(N121), .Z(c[122]) );
  AN2D0 C6390 ( .A1(p[120]), .A2(c[120]), .Z(N120) );
  OR2D0 C6389 ( .A1(g[120]), .A2(N120), .Z(c[121]) );
  AN2D0 C6388 ( .A1(p[119]), .A2(c[119]), .Z(N119) );
  OR2D0 C6387 ( .A1(g[119]), .A2(N119), .Z(c[120]) );
  AN2D0 C6386 ( .A1(p[118]), .A2(c[118]), .Z(N118) );
  OR2D0 C6385 ( .A1(g[118]), .A2(N118), .Z(c[119]) );
  AN2D0 C6384 ( .A1(p[117]), .A2(c[117]), .Z(N117) );
  OR2D0 C6383 ( .A1(g[117]), .A2(N117), .Z(c[118]) );
  AN2D0 C6382 ( .A1(p[116]), .A2(c[116]), .Z(N116) );
  OR2D0 C6381 ( .A1(g[116]), .A2(N116), .Z(c[117]) );
  AN2D0 C6380 ( .A1(p[115]), .A2(c[115]), .Z(N115) );
  OR2D0 C6379 ( .A1(g[115]), .A2(N115), .Z(c[116]) );
  AN2D0 C6378 ( .A1(p[114]), .A2(c[114]), .Z(N114) );
  OR2D0 C6377 ( .A1(g[114]), .A2(N114), .Z(c[115]) );
  AN2D0 C6376 ( .A1(p[113]), .A2(c[113]), .Z(N113) );
  OR2D0 C6375 ( .A1(g[113]), .A2(N113), .Z(c[114]) );
  AN2D0 C6374 ( .A1(p[112]), .A2(c[112]), .Z(N112) );
  OR2D0 C6373 ( .A1(g[112]), .A2(N112), .Z(c[113]) );
  AN2D0 C6372 ( .A1(p[111]), .A2(c[111]), .Z(N111) );
  OR2D0 C6371 ( .A1(g[111]), .A2(N111), .Z(c[112]) );
  AN2D0 C6370 ( .A1(p[110]), .A2(c[110]), .Z(N110) );
  OR2D0 C6369 ( .A1(g[110]), .A2(N110), .Z(c[111]) );
  AN2D0 C6368 ( .A1(p[109]), .A2(c[109]), .Z(N109) );
  OR2D0 C6367 ( .A1(g[109]), .A2(N109), .Z(c[110]) );
  AN2D0 C6366 ( .A1(p[108]), .A2(c[108]), .Z(N108) );
  OR2D0 C6365 ( .A1(g[108]), .A2(N108), .Z(c[109]) );
  AN2D0 C6364 ( .A1(p[107]), .A2(c[107]), .Z(N107) );
  OR2D0 C6363 ( .A1(g[107]), .A2(N107), .Z(c[108]) );
  AN2D0 C6362 ( .A1(p[106]), .A2(c[106]), .Z(N106) );
  OR2D0 C6361 ( .A1(g[106]), .A2(N106), .Z(c[107]) );
  AN2D0 C6360 ( .A1(p[105]), .A2(c[105]), .Z(N105) );
  OR2D0 C6359 ( .A1(g[105]), .A2(N105), .Z(c[106]) );
  AN2D0 C6358 ( .A1(p[104]), .A2(c[104]), .Z(N104) );
  OR2D0 C6357 ( .A1(g[104]), .A2(N104), .Z(c[105]) );
  AN2D0 C6356 ( .A1(p[103]), .A2(c[103]), .Z(N103) );
  OR2D0 C6355 ( .A1(g[103]), .A2(N103), .Z(c[104]) );
  AN2D0 C6354 ( .A1(p[102]), .A2(c[102]), .Z(N102) );
  OR2D0 C6353 ( .A1(g[102]), .A2(N102), .Z(c[103]) );
  AN2D0 C6352 ( .A1(p[101]), .A2(c[101]), .Z(N101) );
  OR2D0 C6351 ( .A1(g[101]), .A2(N101), .Z(c[102]) );
  AN2D0 C6350 ( .A1(p[100]), .A2(c[100]), .Z(N100) );
  OR2D0 C6349 ( .A1(g[100]), .A2(N100), .Z(c[101]) );
  AN2D0 C6348 ( .A1(p[99]), .A2(c[99]), .Z(N99) );
  OR2D0 C6347 ( .A1(g[99]), .A2(N99), .Z(c[100]) );
  AN2D0 C6346 ( .A1(p[98]), .A2(c[98]), .Z(N98) );
  OR2D0 C6345 ( .A1(g[98]), .A2(N98), .Z(c[99]) );
  AN2D0 C6344 ( .A1(p[97]), .A2(c[97]), .Z(N97) );
  OR2D0 C6343 ( .A1(g[97]), .A2(N97), .Z(c[98]) );
  AN2D0 C6342 ( .A1(p[96]), .A2(c[96]), .Z(N96) );
  OR2D0 C6341 ( .A1(g[96]), .A2(N96), .Z(c[97]) );
  AN2D0 C6340 ( .A1(p[95]), .A2(c[95]), .Z(N95) );
  OR2D0 C6339 ( .A1(g[95]), .A2(N95), .Z(c[96]) );
  AN2D0 C6338 ( .A1(p[94]), .A2(c[94]), .Z(N94) );
  OR2D0 C6337 ( .A1(g[94]), .A2(N94), .Z(c[95]) );
  AN2D0 C6336 ( .A1(p[93]), .A2(c[93]), .Z(N93) );
  OR2D0 C6335 ( .A1(g[93]), .A2(N93), .Z(c[94]) );
  AN2D0 C6334 ( .A1(p[92]), .A2(c[92]), .Z(N92) );
  OR2D0 C6333 ( .A1(g[92]), .A2(N92), .Z(c[93]) );
  AN2D0 C6332 ( .A1(p[91]), .A2(c[91]), .Z(N91) );
  OR2D0 C6331 ( .A1(g[91]), .A2(N91), .Z(c[92]) );
  AN2D0 C6330 ( .A1(p[90]), .A2(c[90]), .Z(N90) );
  OR2D0 C6329 ( .A1(g[90]), .A2(N90), .Z(c[91]) );
  AN2D0 C6328 ( .A1(p[89]), .A2(c[89]), .Z(N89) );
  OR2D0 C6327 ( .A1(g[89]), .A2(N89), .Z(c[90]) );
  AN2D0 C6326 ( .A1(p[88]), .A2(c[88]), .Z(N88) );
  OR2D0 C6325 ( .A1(g[88]), .A2(N88), .Z(c[89]) );
  AN2D0 C6324 ( .A1(p[87]), .A2(c[87]), .Z(N87) );
  OR2D0 C6323 ( .A1(g[87]), .A2(N87), .Z(c[88]) );
  AN2D0 C6322 ( .A1(p[86]), .A2(c[86]), .Z(N86) );
  OR2D0 C6321 ( .A1(g[86]), .A2(N86), .Z(c[87]) );
  AN2D0 C6320 ( .A1(p[85]), .A2(c[85]), .Z(N85) );
  OR2D0 C6319 ( .A1(g[85]), .A2(N85), .Z(c[86]) );
  AN2D0 C6318 ( .A1(p[84]), .A2(c[84]), .Z(N84) );
  OR2D0 C6317 ( .A1(g[84]), .A2(N84), .Z(c[85]) );
  AN2D0 C6316 ( .A1(p[83]), .A2(c[83]), .Z(N83) );
  OR2D0 C6315 ( .A1(g[83]), .A2(N83), .Z(c[84]) );
  AN2D0 C6314 ( .A1(p[82]), .A2(c[82]), .Z(N82) );
  OR2D0 C6313 ( .A1(g[82]), .A2(N82), .Z(c[83]) );
  AN2D0 C6312 ( .A1(p[81]), .A2(c[81]), .Z(N81) );
  OR2D0 C6311 ( .A1(g[81]), .A2(N81), .Z(c[82]) );
  AN2D0 C6310 ( .A1(p[80]), .A2(c[80]), .Z(N80) );
  OR2D0 C6309 ( .A1(g[80]), .A2(N80), .Z(c[81]) );
  AN2D0 C6308 ( .A1(p[79]), .A2(c[79]), .Z(N79) );
  OR2D0 C6307 ( .A1(g[79]), .A2(N79), .Z(c[80]) );
  AN2D0 C6306 ( .A1(p[78]), .A2(c[78]), .Z(N78) );
  OR2D0 C6305 ( .A1(g[78]), .A2(N78), .Z(c[79]) );
  AN2D0 C6304 ( .A1(p[77]), .A2(c[77]), .Z(N77) );
  OR2D0 C6303 ( .A1(g[77]), .A2(N77), .Z(c[78]) );
  AN2D0 C6302 ( .A1(p[76]), .A2(c[76]), .Z(N76) );
  OR2D0 C6301 ( .A1(g[76]), .A2(N76), .Z(c[77]) );
  AN2D0 C6300 ( .A1(p[75]), .A2(c[75]), .Z(N75) );
  OR2D0 C6299 ( .A1(g[75]), .A2(N75), .Z(c[76]) );
  AN2D0 C6298 ( .A1(p[74]), .A2(c[74]), .Z(N74) );
  OR2D0 C6297 ( .A1(g[74]), .A2(N74), .Z(c[75]) );
  AN2D0 C6296 ( .A1(p[73]), .A2(c[73]), .Z(N73) );
  OR2D0 C6295 ( .A1(g[73]), .A2(N73), .Z(c[74]) );
  AN2D0 C6294 ( .A1(p[72]), .A2(c[72]), .Z(N72) );
  OR2D0 C6293 ( .A1(g[72]), .A2(N72), .Z(c[73]) );
  AN2D0 C6292 ( .A1(p[71]), .A2(c[71]), .Z(N71) );
  OR2D0 C6291 ( .A1(g[71]), .A2(N71), .Z(c[72]) );
  AN2D0 C6290 ( .A1(p[70]), .A2(c[70]), .Z(N70) );
  OR2D0 C6289 ( .A1(g[70]), .A2(N70), .Z(c[71]) );
  AN2D0 C6288 ( .A1(p[69]), .A2(c[69]), .Z(N69) );
  OR2D0 C6287 ( .A1(g[69]), .A2(N69), .Z(c[70]) );
  AN2D0 C6286 ( .A1(p[68]), .A2(c[68]), .Z(N68) );
  OR2D0 C6285 ( .A1(g[68]), .A2(N68), .Z(c[69]) );
  AN2D0 C6284 ( .A1(p[67]), .A2(c[67]), .Z(N67) );
  OR2D0 C6283 ( .A1(g[67]), .A2(N67), .Z(c[68]) );
  AN2D0 C6282 ( .A1(p[66]), .A2(c[66]), .Z(N66) );
  OR2D0 C6281 ( .A1(g[66]), .A2(N66), .Z(c[67]) );
  AN2D0 C6280 ( .A1(p[65]), .A2(c[65]), .Z(N65) );
  OR2D0 C6279 ( .A1(g[65]), .A2(N65), .Z(c[66]) );
  AN2D0 C6278 ( .A1(p[64]), .A2(c[64]), .Z(N64) );
  OR2D0 C6277 ( .A1(g[64]), .A2(N64), .Z(c[65]) );
  AN2D0 C6276 ( .A1(p[63]), .A2(c[63]), .Z(N63) );
  OR2D0 C6275 ( .A1(g[63]), .A2(N63), .Z(c[64]) );
  AN2D0 C6274 ( .A1(p[62]), .A2(c[62]), .Z(N62) );
  OR2D0 C6273 ( .A1(g[62]), .A2(N62), .Z(c[63]) );
  AN2D0 C6272 ( .A1(p[61]), .A2(c[61]), .Z(N61) );
  OR2D0 C6271 ( .A1(g[61]), .A2(N61), .Z(c[62]) );
  AN2D0 C6270 ( .A1(p[60]), .A2(c[60]), .Z(N60) );
  OR2D0 C6269 ( .A1(g[60]), .A2(N60), .Z(c[61]) );
  AN2D0 C6268 ( .A1(p[59]), .A2(c[59]), .Z(N59) );
  OR2D0 C6267 ( .A1(g[59]), .A2(N59), .Z(c[60]) );
  AN2D0 C6266 ( .A1(p[58]), .A2(c[58]), .Z(N58) );
  OR2D0 C6265 ( .A1(g[58]), .A2(N58), .Z(c[59]) );
  AN2D0 C6264 ( .A1(p[57]), .A2(c[57]), .Z(N57) );
  OR2D0 C6263 ( .A1(g[57]), .A2(N57), .Z(c[58]) );
  AN2D0 C6262 ( .A1(p[56]), .A2(c[56]), .Z(N56) );
  OR2D0 C6261 ( .A1(g[56]), .A2(N56), .Z(c[57]) );
  AN2D0 C6260 ( .A1(p[55]), .A2(c[55]), .Z(N55) );
  OR2D0 C6259 ( .A1(g[55]), .A2(N55), .Z(c[56]) );
  AN2D0 C6258 ( .A1(p[54]), .A2(c[54]), .Z(N54) );
  OR2D0 C6257 ( .A1(g[54]), .A2(N54), .Z(c[55]) );
  AN2D0 C6256 ( .A1(p[53]), .A2(c[53]), .Z(N53) );
  OR2D0 C6255 ( .A1(g[53]), .A2(N53), .Z(c[54]) );
  AN2D0 C6254 ( .A1(p[52]), .A2(c[52]), .Z(N52) );
  OR2D0 C6253 ( .A1(g[52]), .A2(N52), .Z(c[53]) );
  AN2D0 C6252 ( .A1(p[51]), .A2(c[51]), .Z(N51) );
  OR2D0 C6251 ( .A1(g[51]), .A2(N51), .Z(c[52]) );
  AN2D0 C6250 ( .A1(p[50]), .A2(c[50]), .Z(N50) );
  OR2D0 C6249 ( .A1(g[50]), .A2(N50), .Z(c[51]) );
  AN2D0 C6248 ( .A1(p[49]), .A2(c[49]), .Z(N49) );
  OR2D0 C6247 ( .A1(g[49]), .A2(N49), .Z(c[50]) );
  AN2D0 C6246 ( .A1(p[48]), .A2(c[48]), .Z(N48) );
  OR2D0 C6245 ( .A1(g[48]), .A2(N48), .Z(c[49]) );
  AN2D0 C6244 ( .A1(p[47]), .A2(c[47]), .Z(N47) );
  OR2D0 C6243 ( .A1(g[47]), .A2(N47), .Z(c[48]) );
  AN2D0 C6242 ( .A1(p[46]), .A2(c[46]), .Z(N46) );
  OR2D0 C6241 ( .A1(g[46]), .A2(N46), .Z(c[47]) );
  AN2D0 C6240 ( .A1(p[45]), .A2(c[45]), .Z(N45) );
  OR2D0 C6239 ( .A1(g[45]), .A2(N45), .Z(c[46]) );
  AN2D0 C6238 ( .A1(p[44]), .A2(c[44]), .Z(N44) );
  OR2D0 C6237 ( .A1(g[44]), .A2(N44), .Z(c[45]) );
  AN2D0 C6236 ( .A1(p[43]), .A2(c[43]), .Z(N43) );
  OR2D0 C6235 ( .A1(g[43]), .A2(N43), .Z(c[44]) );
  AN2D0 C6234 ( .A1(p[42]), .A2(c[42]), .Z(N42) );
  OR2D0 C6233 ( .A1(g[42]), .A2(N42), .Z(c[43]) );
  AN2D0 C6232 ( .A1(p[41]), .A2(c[41]), .Z(N41) );
  OR2D0 C6231 ( .A1(g[41]), .A2(N41), .Z(c[42]) );
  AN2D0 C6230 ( .A1(p[40]), .A2(c[40]), .Z(N40) );
  OR2D0 C6229 ( .A1(g[40]), .A2(N40), .Z(c[41]) );
  AN2D0 C6228 ( .A1(p[39]), .A2(c[39]), .Z(N39) );
  OR2D0 C6227 ( .A1(g[39]), .A2(N39), .Z(c[40]) );
  AN2D0 C6226 ( .A1(p[38]), .A2(c[38]), .Z(N38) );
  OR2D0 C6225 ( .A1(g[38]), .A2(N38), .Z(c[39]) );
  AN2D0 C6224 ( .A1(p[37]), .A2(c[37]), .Z(N37) );
  OR2D0 C6223 ( .A1(g[37]), .A2(N37), .Z(c[38]) );
  AN2D0 C6222 ( .A1(p[36]), .A2(c[36]), .Z(N36) );
  OR2D0 C6221 ( .A1(g[36]), .A2(N36), .Z(c[37]) );
  AN2D0 C6220 ( .A1(p[35]), .A2(c[35]), .Z(N35) );
  OR2D0 C6219 ( .A1(g[35]), .A2(N35), .Z(c[36]) );
  AN2D0 C6218 ( .A1(p[34]), .A2(c[34]), .Z(N34) );
  OR2D0 C6217 ( .A1(g[34]), .A2(N34), .Z(c[35]) );
  AN2D0 C6216 ( .A1(p[33]), .A2(c[33]), .Z(N33) );
  OR2D0 C6215 ( .A1(g[33]), .A2(N33), .Z(c[34]) );
  AN2D0 C6214 ( .A1(p[32]), .A2(c[32]), .Z(N32) );
  OR2D0 C6213 ( .A1(g[32]), .A2(N32), .Z(c[33]) );
  AN2D0 C6212 ( .A1(p[31]), .A2(c[31]), .Z(N31) );
  OR2D0 C6211 ( .A1(g[31]), .A2(N31), .Z(c[32]) );
  AN2D0 C6210 ( .A1(p[30]), .A2(c[30]), .Z(N30) );
  OR2D0 C6209 ( .A1(g[30]), .A2(N30), .Z(c[31]) );
  AN2D0 C6208 ( .A1(p[29]), .A2(c[29]), .Z(N29) );
  OR2D0 C6207 ( .A1(g[29]), .A2(N29), .Z(c[30]) );
  AN2D0 C6206 ( .A1(p[28]), .A2(c[28]), .Z(N28) );
  OR2D0 C6205 ( .A1(g[28]), .A2(N28), .Z(c[29]) );
  AN2D0 C6204 ( .A1(p[27]), .A2(c[27]), .Z(N27) );
  OR2D0 C6203 ( .A1(g[27]), .A2(N27), .Z(c[28]) );
  AN2D0 C6202 ( .A1(p[26]), .A2(c[26]), .Z(N26) );
  OR2D0 C6201 ( .A1(g[26]), .A2(N26), .Z(c[27]) );
  AN2D0 C6200 ( .A1(p[25]), .A2(c[25]), .Z(N25) );
  OR2D0 C6199 ( .A1(g[25]), .A2(N25), .Z(c[26]) );
  AN2D0 C6198 ( .A1(p[24]), .A2(c[24]), .Z(N24) );
  OR2D0 C6197 ( .A1(g[24]), .A2(N24), .Z(c[25]) );
  AN2D0 C6196 ( .A1(p[23]), .A2(c[23]), .Z(N23) );
  OR2D0 C6195 ( .A1(g[23]), .A2(N23), .Z(c[24]) );
  AN2D0 C6194 ( .A1(p[22]), .A2(c[22]), .Z(N22) );
  OR2D0 C6193 ( .A1(g[22]), .A2(N22), .Z(c[23]) );
  AN2D0 C6192 ( .A1(p[21]), .A2(c[21]), .Z(N21) );
  OR2D0 C6191 ( .A1(g[21]), .A2(N21), .Z(c[22]) );
  AN2D0 C6190 ( .A1(p[20]), .A2(c[20]), .Z(N20) );
  OR2D0 C6189 ( .A1(g[20]), .A2(N20), .Z(c[21]) );
  AN2D0 C6188 ( .A1(p[19]), .A2(c[19]), .Z(N19) );
  OR2D0 C6187 ( .A1(g[19]), .A2(N19), .Z(c[20]) );
  AN2D0 C6186 ( .A1(p[18]), .A2(c[18]), .Z(N18) );
  OR2D0 C6185 ( .A1(g[18]), .A2(N18), .Z(c[19]) );
  AN2D0 C6184 ( .A1(p[17]), .A2(c[17]), .Z(N17) );
  OR2D0 C6183 ( .A1(g[17]), .A2(N17), .Z(c[18]) );
  AN2D0 C6182 ( .A1(p[16]), .A2(c[16]), .Z(N16) );
  OR2D0 C6181 ( .A1(g[16]), .A2(N16), .Z(c[17]) );
  AN2D0 C6180 ( .A1(p[15]), .A2(c[15]), .Z(N15) );
  OR2D0 C6179 ( .A1(g[15]), .A2(N15), .Z(c[16]) );
  AN2D0 C6178 ( .A1(p[14]), .A2(c[14]), .Z(N14) );
  OR2D0 C6177 ( .A1(g[14]), .A2(N14), .Z(c[15]) );
  AN2D0 C6176 ( .A1(p[13]), .A2(c[13]), .Z(N13) );
  OR2D0 C6175 ( .A1(g[13]), .A2(N13), .Z(c[14]) );
  AN2D0 C6174 ( .A1(p[12]), .A2(c[12]), .Z(N12) );
  OR2D0 C6173 ( .A1(g[12]), .A2(N12), .Z(c[13]) );
  AN2D0 C6172 ( .A1(p[11]), .A2(c[11]), .Z(N11) );
  OR2D0 C6171 ( .A1(g[11]), .A2(N11), .Z(c[12]) );
  AN2D0 C6170 ( .A1(p[10]), .A2(c[10]), .Z(N10) );
  OR2D0 C6169 ( .A1(g[10]), .A2(N10), .Z(c[11]) );
  AN2D0 C6168 ( .A1(p[9]), .A2(c[9]), .Z(N9) );
  OR2D0 C6167 ( .A1(g[9]), .A2(N9), .Z(c[10]) );
  AN2D0 C6166 ( .A1(p[8]), .A2(c[8]), .Z(N8) );
  OR2D0 C6165 ( .A1(g[8]), .A2(N8), .Z(c[9]) );
  AN2D0 C6164 ( .A1(p[7]), .A2(c[7]), .Z(N7) );
  OR2D0 C6163 ( .A1(g[7]), .A2(N7), .Z(c[8]) );
  AN2D0 C6162 ( .A1(p[6]), .A2(c[6]), .Z(N6) );
  OR2D0 C6161 ( .A1(g[6]), .A2(N6), .Z(c[7]) );
  AN2D0 C6160 ( .A1(p[5]), .A2(c[5]), .Z(N5) );
  OR2D0 C6159 ( .A1(g[5]), .A2(N5), .Z(c[6]) );
  AN2D0 C6158 ( .A1(p[4]), .A2(c[4]), .Z(N4) );
  OR2D0 C6157 ( .A1(g[4]), .A2(N4), .Z(c[5]) );
  AN2D0 C6156 ( .A1(p[3]), .A2(c[3]), .Z(N3) );
  OR2D0 C6155 ( .A1(g[3]), .A2(N3), .Z(c[4]) );
  AN2D0 C6154 ( .A1(p[2]), .A2(c[2]), .Z(N2) );
  OR2D0 C6153 ( .A1(g[2]), .A2(N2), .Z(c[3]) );
  AN2D0 C6152 ( .A1(p[1]), .A2(c[1]), .Z(N1) );
  OR2D0 C6151 ( .A1(g[1]), .A2(N1), .Z(c[2]) );
  AN2D0 C6150 ( .A1(p[0]), .A2(cin), .Z(N0) );
  OR2D0 C6149 ( .A1(g[0]), .A2(N0), .Z(c[1]) );
  XOR2D0 C6148 ( .A1(a[0]), .A2(b[0]), .Z(p[0]) );
  XOR2D0 C6147 ( .A1(a[1]), .A2(b[1]), .Z(p[1]) );
  XOR2D0 C6146 ( .A1(a[2]), .A2(b[2]), .Z(p[2]) );
  XOR2D0 C6145 ( .A1(a[3]), .A2(b[3]), .Z(p[3]) );
  XOR2D0 C6144 ( .A1(a[4]), .A2(b[4]), .Z(p[4]) );
  XOR2D0 C6143 ( .A1(a[5]), .A2(b[5]), .Z(p[5]) );
  XOR2D0 C6142 ( .A1(a[6]), .A2(b[6]), .Z(p[6]) );
  XOR2D0 C6141 ( .A1(a[7]), .A2(b[7]), .Z(p[7]) );
  XOR2D0 C6140 ( .A1(a[8]), .A2(b[8]), .Z(p[8]) );
  XOR2D0 C6139 ( .A1(a[9]), .A2(b[9]), .Z(p[9]) );
  XOR2D0 C6138 ( .A1(a[10]), .A2(b[10]), .Z(p[10]) );
  XOR2D0 C6137 ( .A1(a[11]), .A2(b[11]), .Z(p[11]) );
  XOR2D0 C6136 ( .A1(a[12]), .A2(b[12]), .Z(p[12]) );
  XOR2D0 C6135 ( .A1(a[13]), .A2(b[13]), .Z(p[13]) );
  XOR2D0 C6134 ( .A1(a[14]), .A2(b[14]), .Z(p[14]) );
  XOR2D0 C6133 ( .A1(a[15]), .A2(b[15]), .Z(p[15]) );
  XOR2D0 C6132 ( .A1(a[16]), .A2(b[16]), .Z(p[16]) );
  XOR2D0 C6131 ( .A1(a[17]), .A2(b[17]), .Z(p[17]) );
  XOR2D0 C6130 ( .A1(a[18]), .A2(b[18]), .Z(p[18]) );
  XOR2D0 C6129 ( .A1(a[19]), .A2(b[19]), .Z(p[19]) );
  XOR2D0 C6128 ( .A1(a[20]), .A2(b[20]), .Z(p[20]) );
  XOR2D0 C6127 ( .A1(a[21]), .A2(b[21]), .Z(p[21]) );
  XOR2D0 C6126 ( .A1(a[22]), .A2(b[22]), .Z(p[22]) );
  XOR2D0 C6125 ( .A1(a[23]), .A2(b[23]), .Z(p[23]) );
  XOR2D0 C6124 ( .A1(a[24]), .A2(b[24]), .Z(p[24]) );
  XOR2D0 C6123 ( .A1(a[25]), .A2(b[25]), .Z(p[25]) );
  XOR2D0 C6122 ( .A1(a[26]), .A2(b[26]), .Z(p[26]) );
  XOR2D0 C6121 ( .A1(a[27]), .A2(b[27]), .Z(p[27]) );
  XOR2D0 C6120 ( .A1(a[28]), .A2(b[28]), .Z(p[28]) );
  XOR2D0 C6119 ( .A1(a[29]), .A2(b[29]), .Z(p[29]) );
  XOR2D0 C6118 ( .A1(a[30]), .A2(b[30]), .Z(p[30]) );
  XOR2D0 C6117 ( .A1(a[31]), .A2(b[31]), .Z(p[31]) );
  XOR2D0 C6116 ( .A1(a[32]), .A2(b[32]), .Z(p[32]) );
  XOR2D0 C6115 ( .A1(a[33]), .A2(b[33]), .Z(p[33]) );
  XOR2D0 C6114 ( .A1(a[34]), .A2(b[34]), .Z(p[34]) );
  XOR2D0 C6113 ( .A1(a[35]), .A2(b[35]), .Z(p[35]) );
  XOR2D0 C6112 ( .A1(a[36]), .A2(b[36]), .Z(p[36]) );
  XOR2D0 C6111 ( .A1(a[37]), .A2(b[37]), .Z(p[37]) );
  XOR2D0 C6110 ( .A1(a[38]), .A2(b[38]), .Z(p[38]) );
  XOR2D0 C6109 ( .A1(a[39]), .A2(b[39]), .Z(p[39]) );
  XOR2D0 C6108 ( .A1(a[40]), .A2(b[40]), .Z(p[40]) );
  XOR2D0 C6107 ( .A1(a[41]), .A2(b[41]), .Z(p[41]) );
  XOR2D0 C6106 ( .A1(a[42]), .A2(b[42]), .Z(p[42]) );
  XOR2D0 C6105 ( .A1(a[43]), .A2(b[43]), .Z(p[43]) );
  XOR2D0 C6104 ( .A1(a[44]), .A2(b[44]), .Z(p[44]) );
  XOR2D0 C6103 ( .A1(a[45]), .A2(b[45]), .Z(p[45]) );
  XOR2D0 C6102 ( .A1(a[46]), .A2(b[46]), .Z(p[46]) );
  XOR2D0 C6101 ( .A1(a[47]), .A2(b[47]), .Z(p[47]) );
  XOR2D0 C6100 ( .A1(a[48]), .A2(b[48]), .Z(p[48]) );
  XOR2D0 C6099 ( .A1(a[49]), .A2(b[49]), .Z(p[49]) );
  XOR2D0 C6098 ( .A1(a[50]), .A2(b[50]), .Z(p[50]) );
  XOR2D0 C6097 ( .A1(a[51]), .A2(b[51]), .Z(p[51]) );
  XOR2D0 C6096 ( .A1(a[52]), .A2(b[52]), .Z(p[52]) );
  XOR2D0 C6095 ( .A1(a[53]), .A2(b[53]), .Z(p[53]) );
  XOR2D0 C6094 ( .A1(a[54]), .A2(b[54]), .Z(p[54]) );
  XOR2D0 C6093 ( .A1(a[55]), .A2(b[55]), .Z(p[55]) );
  XOR2D0 C6092 ( .A1(a[56]), .A2(b[56]), .Z(p[56]) );
  XOR2D0 C6091 ( .A1(a[57]), .A2(b[57]), .Z(p[57]) );
  XOR2D0 C6090 ( .A1(a[58]), .A2(b[58]), .Z(p[58]) );
  XOR2D0 C6089 ( .A1(a[59]), .A2(b[59]), .Z(p[59]) );
  XOR2D0 C6088 ( .A1(a[60]), .A2(b[60]), .Z(p[60]) );
  XOR2D0 C6087 ( .A1(a[61]), .A2(b[61]), .Z(p[61]) );
  XOR2D0 C6086 ( .A1(a[62]), .A2(b[62]), .Z(p[62]) );
  XOR2D0 C6085 ( .A1(a[63]), .A2(b[63]), .Z(p[63]) );
  XOR2D0 C6084 ( .A1(a[64]), .A2(b[64]), .Z(p[64]) );
  XOR2D0 C6083 ( .A1(a[65]), .A2(b[65]), .Z(p[65]) );
  XOR2D0 C6082 ( .A1(a[66]), .A2(b[66]), .Z(p[66]) );
  XOR2D0 C6081 ( .A1(a[67]), .A2(b[67]), .Z(p[67]) );
  XOR2D0 C6080 ( .A1(a[68]), .A2(b[68]), .Z(p[68]) );
  XOR2D0 C6079 ( .A1(a[69]), .A2(b[69]), .Z(p[69]) );
  XOR2D0 C6078 ( .A1(a[70]), .A2(b[70]), .Z(p[70]) );
  XOR2D0 C6077 ( .A1(a[71]), .A2(b[71]), .Z(p[71]) );
  XOR2D0 C6076 ( .A1(a[72]), .A2(b[72]), .Z(p[72]) );
  XOR2D0 C6075 ( .A1(a[73]), .A2(b[73]), .Z(p[73]) );
  XOR2D0 C6074 ( .A1(a[74]), .A2(b[74]), .Z(p[74]) );
  XOR2D0 C6073 ( .A1(a[75]), .A2(b[75]), .Z(p[75]) );
  XOR2D0 C6072 ( .A1(a[76]), .A2(b[76]), .Z(p[76]) );
  XOR2D0 C6071 ( .A1(a[77]), .A2(b[77]), .Z(p[77]) );
  XOR2D0 C6070 ( .A1(a[78]), .A2(b[78]), .Z(p[78]) );
  XOR2D0 C6069 ( .A1(a[79]), .A2(b[79]), .Z(p[79]) );
  XOR2D0 C6068 ( .A1(a[80]), .A2(b[80]), .Z(p[80]) );
  XOR2D0 C6067 ( .A1(a[81]), .A2(b[81]), .Z(p[81]) );
  XOR2D0 C6066 ( .A1(a[82]), .A2(b[82]), .Z(p[82]) );
  XOR2D0 C6065 ( .A1(a[83]), .A2(b[83]), .Z(p[83]) );
  XOR2D0 C6064 ( .A1(a[84]), .A2(b[84]), .Z(p[84]) );
  XOR2D0 C6063 ( .A1(a[85]), .A2(b[85]), .Z(p[85]) );
  XOR2D0 C6062 ( .A1(a[86]), .A2(b[86]), .Z(p[86]) );
  XOR2D0 C6061 ( .A1(a[87]), .A2(b[87]), .Z(p[87]) );
  XOR2D0 C6060 ( .A1(a[88]), .A2(b[88]), .Z(p[88]) );
  XOR2D0 C6059 ( .A1(a[89]), .A2(b[89]), .Z(p[89]) );
  XOR2D0 C6058 ( .A1(a[90]), .A2(b[90]), .Z(p[90]) );
  XOR2D0 C6057 ( .A1(a[91]), .A2(b[91]), .Z(p[91]) );
  XOR2D0 C6056 ( .A1(a[92]), .A2(b[92]), .Z(p[92]) );
  XOR2D0 C6055 ( .A1(a[93]), .A2(b[93]), .Z(p[93]) );
  XOR2D0 C6054 ( .A1(a[94]), .A2(b[94]), .Z(p[94]) );
  XOR2D0 C6053 ( .A1(a[95]), .A2(b[95]), .Z(p[95]) );
  XOR2D0 C6052 ( .A1(a[96]), .A2(b[96]), .Z(p[96]) );
  XOR2D0 C6051 ( .A1(a[97]), .A2(b[97]), .Z(p[97]) );
  XOR2D0 C6050 ( .A1(a[98]), .A2(b[98]), .Z(p[98]) );
  XOR2D0 C6049 ( .A1(a[99]), .A2(b[99]), .Z(p[99]) );
  XOR2D0 C6048 ( .A1(a[100]), .A2(b[100]), .Z(p[100]) );
  XOR2D0 C6047 ( .A1(a[101]), .A2(b[101]), .Z(p[101]) );
  XOR2D0 C6046 ( .A1(a[102]), .A2(b[102]), .Z(p[102]) );
  XOR2D0 C6045 ( .A1(a[103]), .A2(b[103]), .Z(p[103]) );
  XOR2D0 C6044 ( .A1(a[104]), .A2(b[104]), .Z(p[104]) );
  XOR2D0 C6043 ( .A1(a[105]), .A2(b[105]), .Z(p[105]) );
  XOR2D0 C6042 ( .A1(a[106]), .A2(b[106]), .Z(p[106]) );
  XOR2D0 C6041 ( .A1(a[107]), .A2(b[107]), .Z(p[107]) );
  XOR2D0 C6040 ( .A1(a[108]), .A2(b[108]), .Z(p[108]) );
  XOR2D0 C6039 ( .A1(a[109]), .A2(b[109]), .Z(p[109]) );
  XOR2D0 C6038 ( .A1(a[110]), .A2(b[110]), .Z(p[110]) );
  XOR2D0 C6037 ( .A1(a[111]), .A2(b[111]), .Z(p[111]) );
  XOR2D0 C6036 ( .A1(a[112]), .A2(b[112]), .Z(p[112]) );
  XOR2D0 C6035 ( .A1(a[113]), .A2(b[113]), .Z(p[113]) );
  XOR2D0 C6034 ( .A1(a[114]), .A2(b[114]), .Z(p[114]) );
  XOR2D0 C6033 ( .A1(a[115]), .A2(b[115]), .Z(p[115]) );
  XOR2D0 C6032 ( .A1(a[116]), .A2(b[116]), .Z(p[116]) );
  XOR2D0 C6031 ( .A1(a[117]), .A2(b[117]), .Z(p[117]) );
  XOR2D0 C6030 ( .A1(a[118]), .A2(b[118]), .Z(p[118]) );
  XOR2D0 C6029 ( .A1(a[119]), .A2(b[119]), .Z(p[119]) );
  XOR2D0 C6028 ( .A1(a[120]), .A2(b[120]), .Z(p[120]) );
  XOR2D0 C6027 ( .A1(a[121]), .A2(b[121]), .Z(p[121]) );
  XOR2D0 C6026 ( .A1(a[122]), .A2(b[122]), .Z(p[122]) );
  XOR2D0 C6025 ( .A1(a[123]), .A2(b[123]), .Z(p[123]) );
  XOR2D0 C6024 ( .A1(a[124]), .A2(b[124]), .Z(p[124]) );
  XOR2D0 C6023 ( .A1(a[125]), .A2(b[125]), .Z(p[125]) );
  XOR2D0 C6022 ( .A1(a[126]), .A2(b[126]), .Z(p[126]) );
  XOR2D0 C6021 ( .A1(a[127]), .A2(b[127]), .Z(p[127]) );
  XOR2D0 C6020 ( .A1(a[128]), .A2(b[128]), .Z(p[128]) );
  XOR2D0 C6019 ( .A1(a[129]), .A2(b[129]), .Z(p[129]) );
  XOR2D0 C6018 ( .A1(a[130]), .A2(b[130]), .Z(p[130]) );
  XOR2D0 C6017 ( .A1(a[131]), .A2(b[131]), .Z(p[131]) );
  XOR2D0 C6016 ( .A1(a[132]), .A2(b[132]), .Z(p[132]) );
  XOR2D0 C6015 ( .A1(a[133]), .A2(b[133]), .Z(p[133]) );
  XOR2D0 C6014 ( .A1(a[134]), .A2(b[134]), .Z(p[134]) );
  XOR2D0 C6013 ( .A1(a[135]), .A2(b[135]), .Z(p[135]) );
  XOR2D0 C6012 ( .A1(a[136]), .A2(b[136]), .Z(p[136]) );
  XOR2D0 C6011 ( .A1(a[137]), .A2(b[137]), .Z(p[137]) );
  XOR2D0 C6010 ( .A1(a[138]), .A2(b[138]), .Z(p[138]) );
  XOR2D0 C6009 ( .A1(a[139]), .A2(b[139]), .Z(p[139]) );
  XOR2D0 C6008 ( .A1(a[140]), .A2(b[140]), .Z(p[140]) );
  XOR2D0 C6007 ( .A1(a[141]), .A2(b[141]), .Z(p[141]) );
  XOR2D0 C6006 ( .A1(a[142]), .A2(b[142]), .Z(p[142]) );
  XOR2D0 C6005 ( .A1(a[143]), .A2(b[143]), .Z(p[143]) );
  XOR2D0 C6004 ( .A1(a[144]), .A2(b[144]), .Z(p[144]) );
  XOR2D0 C6003 ( .A1(a[145]), .A2(b[145]), .Z(p[145]) );
  XOR2D0 C6002 ( .A1(a[146]), .A2(b[146]), .Z(p[146]) );
  XOR2D0 C6001 ( .A1(a[147]), .A2(b[147]), .Z(p[147]) );
  XOR2D0 C6000 ( .A1(a[148]), .A2(b[148]), .Z(p[148]) );
  XOR2D0 C5999 ( .A1(a[149]), .A2(b[149]), .Z(p[149]) );
  XOR2D0 C5998 ( .A1(a[150]), .A2(b[150]), .Z(p[150]) );
  XOR2D0 C5997 ( .A1(a[151]), .A2(b[151]), .Z(p[151]) );
  XOR2D0 C5996 ( .A1(a[152]), .A2(b[152]), .Z(p[152]) );
  XOR2D0 C5995 ( .A1(a[153]), .A2(b[153]), .Z(p[153]) );
  XOR2D0 C5994 ( .A1(a[154]), .A2(b[154]), .Z(p[154]) );
  XOR2D0 C5993 ( .A1(a[155]), .A2(b[155]), .Z(p[155]) );
  XOR2D0 C5992 ( .A1(a[156]), .A2(b[156]), .Z(p[156]) );
  XOR2D0 C5991 ( .A1(a[157]), .A2(b[157]), .Z(p[157]) );
  XOR2D0 C5990 ( .A1(a[158]), .A2(b[158]), .Z(p[158]) );
  XOR2D0 C5989 ( .A1(a[159]), .A2(b[159]), .Z(p[159]) );
  XOR2D0 C5988 ( .A1(a[160]), .A2(b[160]), .Z(p[160]) );
  XOR2D0 C5987 ( .A1(a[161]), .A2(b[161]), .Z(p[161]) );
  XOR2D0 C5986 ( .A1(a[162]), .A2(b[162]), .Z(p[162]) );
  XOR2D0 C5985 ( .A1(a[163]), .A2(b[163]), .Z(p[163]) );
  XOR2D0 C5984 ( .A1(a[164]), .A2(b[164]), .Z(p[164]) );
  XOR2D0 C5983 ( .A1(a[165]), .A2(b[165]), .Z(p[165]) );
  XOR2D0 C5982 ( .A1(a[166]), .A2(b[166]), .Z(p[166]) );
  XOR2D0 C5981 ( .A1(a[167]), .A2(b[167]), .Z(p[167]) );
  XOR2D0 C5980 ( .A1(a[168]), .A2(b[168]), .Z(p[168]) );
  XOR2D0 C5979 ( .A1(a[169]), .A2(b[169]), .Z(p[169]) );
  XOR2D0 C5978 ( .A1(a[170]), .A2(b[170]), .Z(p[170]) );
  XOR2D0 C5977 ( .A1(a[171]), .A2(b[171]), .Z(p[171]) );
  XOR2D0 C5976 ( .A1(a[172]), .A2(b[172]), .Z(p[172]) );
  XOR2D0 C5975 ( .A1(a[173]), .A2(b[173]), .Z(p[173]) );
  XOR2D0 C5974 ( .A1(a[174]), .A2(b[174]), .Z(p[174]) );
  XOR2D0 C5973 ( .A1(a[175]), .A2(b[175]), .Z(p[175]) );
  XOR2D0 C5972 ( .A1(a[176]), .A2(b[176]), .Z(p[176]) );
  XOR2D0 C5971 ( .A1(a[177]), .A2(b[177]), .Z(p[177]) );
  XOR2D0 C5970 ( .A1(a[178]), .A2(b[178]), .Z(p[178]) );
  XOR2D0 C5969 ( .A1(a[179]), .A2(b[179]), .Z(p[179]) );
  XOR2D0 C5968 ( .A1(a[180]), .A2(b[180]), .Z(p[180]) );
  XOR2D0 C5967 ( .A1(a[181]), .A2(b[181]), .Z(p[181]) );
  XOR2D0 C5966 ( .A1(a[182]), .A2(b[182]), .Z(p[182]) );
  XOR2D0 C5965 ( .A1(a[183]), .A2(b[183]), .Z(p[183]) );
  XOR2D0 C5964 ( .A1(a[184]), .A2(b[184]), .Z(p[184]) );
  XOR2D0 C5963 ( .A1(a[185]), .A2(b[185]), .Z(p[185]) );
  XOR2D0 C5962 ( .A1(a[186]), .A2(b[186]), .Z(p[186]) );
  XOR2D0 C5961 ( .A1(a[187]), .A2(b[187]), .Z(p[187]) );
  XOR2D0 C5960 ( .A1(a[188]), .A2(b[188]), .Z(p[188]) );
  XOR2D0 C5959 ( .A1(a[189]), .A2(b[189]), .Z(p[189]) );
  XOR2D0 C5958 ( .A1(a[190]), .A2(b[190]), .Z(p[190]) );
  XOR2D0 C5957 ( .A1(a[191]), .A2(b[191]), .Z(p[191]) );
  XOR2D0 C5956 ( .A1(a[192]), .A2(b[192]), .Z(p[192]) );
  XOR2D0 C5955 ( .A1(a[193]), .A2(b[193]), .Z(p[193]) );
  XOR2D0 C5954 ( .A1(a[194]), .A2(b[194]), .Z(p[194]) );
  XOR2D0 C5953 ( .A1(a[195]), .A2(b[195]), .Z(p[195]) );
  XOR2D0 C5952 ( .A1(a[196]), .A2(b[196]), .Z(p[196]) );
  XOR2D0 C5951 ( .A1(a[197]), .A2(b[197]), .Z(p[197]) );
  XOR2D0 C5950 ( .A1(a[198]), .A2(b[198]), .Z(p[198]) );
  XOR2D0 C5949 ( .A1(a[199]), .A2(b[199]), .Z(p[199]) );
  XOR2D0 C5948 ( .A1(a[200]), .A2(b[200]), .Z(p[200]) );
  XOR2D0 C5947 ( .A1(a[201]), .A2(b[201]), .Z(p[201]) );
  XOR2D0 C5946 ( .A1(a[202]), .A2(b[202]), .Z(p[202]) );
  XOR2D0 C5945 ( .A1(a[203]), .A2(b[203]), .Z(p[203]) );
  XOR2D0 C5944 ( .A1(a[204]), .A2(b[204]), .Z(p[204]) );
  XOR2D0 C5943 ( .A1(a[205]), .A2(b[205]), .Z(p[205]) );
  XOR2D0 C5942 ( .A1(a[206]), .A2(b[206]), .Z(p[206]) );
  XOR2D0 C5941 ( .A1(a[207]), .A2(b[207]), .Z(p[207]) );
  XOR2D0 C5940 ( .A1(a[208]), .A2(b[208]), .Z(p[208]) );
  XOR2D0 C5939 ( .A1(a[209]), .A2(b[209]), .Z(p[209]) );
  XOR2D0 C5938 ( .A1(a[210]), .A2(b[210]), .Z(p[210]) );
  XOR2D0 C5937 ( .A1(a[211]), .A2(b[211]), .Z(p[211]) );
  XOR2D0 C5936 ( .A1(a[212]), .A2(b[212]), .Z(p[212]) );
  XOR2D0 C5935 ( .A1(a[213]), .A2(b[213]), .Z(p[213]) );
  XOR2D0 C5934 ( .A1(a[214]), .A2(b[214]), .Z(p[214]) );
  XOR2D0 C5933 ( .A1(a[215]), .A2(b[215]), .Z(p[215]) );
  XOR2D0 C5932 ( .A1(a[216]), .A2(b[216]), .Z(p[216]) );
  XOR2D0 C5931 ( .A1(a[217]), .A2(b[217]), .Z(p[217]) );
  XOR2D0 C5930 ( .A1(a[218]), .A2(b[218]), .Z(p[218]) );
  XOR2D0 C5929 ( .A1(a[219]), .A2(b[219]), .Z(p[219]) );
  XOR2D0 C5928 ( .A1(a[220]), .A2(b[220]), .Z(p[220]) );
  XOR2D0 C5927 ( .A1(a[221]), .A2(b[221]), .Z(p[221]) );
  XOR2D0 C5926 ( .A1(a[222]), .A2(b[222]), .Z(p[222]) );
  XOR2D0 C5925 ( .A1(a[223]), .A2(b[223]), .Z(p[223]) );
  XOR2D0 C5924 ( .A1(a[224]), .A2(b[224]), .Z(p[224]) );
  XOR2D0 C5923 ( .A1(a[225]), .A2(b[225]), .Z(p[225]) );
  XOR2D0 C5922 ( .A1(a[226]), .A2(b[226]), .Z(p[226]) );
  XOR2D0 C5921 ( .A1(a[227]), .A2(b[227]), .Z(p[227]) );
  XOR2D0 C5920 ( .A1(a[228]), .A2(b[228]), .Z(p[228]) );
  XOR2D0 C5919 ( .A1(a[229]), .A2(b[229]), .Z(p[229]) );
  XOR2D0 C5918 ( .A1(a[230]), .A2(b[230]), .Z(p[230]) );
  XOR2D0 C5917 ( .A1(a[231]), .A2(b[231]), .Z(p[231]) );
  XOR2D0 C5916 ( .A1(a[232]), .A2(b[232]), .Z(p[232]) );
  XOR2D0 C5915 ( .A1(a[233]), .A2(b[233]), .Z(p[233]) );
  XOR2D0 C5914 ( .A1(a[234]), .A2(b[234]), .Z(p[234]) );
  XOR2D0 C5913 ( .A1(a[235]), .A2(b[235]), .Z(p[235]) );
  XOR2D0 C5912 ( .A1(a[236]), .A2(b[236]), .Z(p[236]) );
  XOR2D0 C5911 ( .A1(a[237]), .A2(b[237]), .Z(p[237]) );
  XOR2D0 C5910 ( .A1(a[238]), .A2(b[238]), .Z(p[238]) );
  XOR2D0 C5909 ( .A1(a[239]), .A2(b[239]), .Z(p[239]) );
  XOR2D0 C5908 ( .A1(a[240]), .A2(b[240]), .Z(p[240]) );
  XOR2D0 C5907 ( .A1(a[241]), .A2(b[241]), .Z(p[241]) );
  XOR2D0 C5906 ( .A1(a[242]), .A2(b[242]), .Z(p[242]) );
  XOR2D0 C5905 ( .A1(a[243]), .A2(b[243]), .Z(p[243]) );
  XOR2D0 C5904 ( .A1(a[244]), .A2(b[244]), .Z(p[244]) );
  XOR2D0 C5903 ( .A1(a[245]), .A2(b[245]), .Z(p[245]) );
  XOR2D0 C5902 ( .A1(a[246]), .A2(b[246]), .Z(p[246]) );
  XOR2D0 C5901 ( .A1(a[247]), .A2(b[247]), .Z(p[247]) );
  XOR2D0 C5900 ( .A1(a[248]), .A2(b[248]), .Z(p[248]) );
  XOR2D0 C5899 ( .A1(a[249]), .A2(b[249]), .Z(p[249]) );
  XOR2D0 C5898 ( .A1(a[250]), .A2(b[250]), .Z(p[250]) );
  XOR2D0 C5897 ( .A1(a[251]), .A2(b[251]), .Z(p[251]) );
  XOR2D0 C5896 ( .A1(a[252]), .A2(b[252]), .Z(p[252]) );
  XOR2D0 C5895 ( .A1(a[253]), .A2(b[253]), .Z(p[253]) );
  XOR2D0 C5894 ( .A1(a[254]), .A2(b[254]), .Z(p[254]) );
  XOR2D0 C5893 ( .A1(a[255]), .A2(b[255]), .Z(p[255]) );
  XOR2D0 C5892 ( .A1(a[256]), .A2(b[256]), .Z(p[256]) );
  XOR2D0 C5891 ( .A1(a[257]), .A2(b[257]), .Z(p[257]) );
  XOR2D0 C5890 ( .A1(a[258]), .A2(b[258]), .Z(p[258]) );
  XOR2D0 C5889 ( .A1(a[259]), .A2(b[259]), .Z(p[259]) );
  XOR2D0 C5888 ( .A1(a[260]), .A2(b[260]), .Z(p[260]) );
  XOR2D0 C5887 ( .A1(a[261]), .A2(b[261]), .Z(p[261]) );
  XOR2D0 C5886 ( .A1(a[262]), .A2(b[262]), .Z(p[262]) );
  XOR2D0 C5885 ( .A1(a[263]), .A2(b[263]), .Z(p[263]) );
  XOR2D0 C5884 ( .A1(a[264]), .A2(b[264]), .Z(p[264]) );
  XOR2D0 C5883 ( .A1(a[265]), .A2(b[265]), .Z(p[265]) );
  XOR2D0 C5882 ( .A1(a[266]), .A2(b[266]), .Z(p[266]) );
  XOR2D0 C5881 ( .A1(a[267]), .A2(b[267]), .Z(p[267]) );
  XOR2D0 C5880 ( .A1(a[268]), .A2(b[268]), .Z(p[268]) );
  XOR2D0 C5879 ( .A1(a[269]), .A2(b[269]), .Z(p[269]) );
  XOR2D0 C5878 ( .A1(a[270]), .A2(b[270]), .Z(p[270]) );
  XOR2D0 C5877 ( .A1(a[271]), .A2(b[271]), .Z(p[271]) );
  XOR2D0 C5876 ( .A1(a[272]), .A2(b[272]), .Z(p[272]) );
  XOR2D0 C5875 ( .A1(a[273]), .A2(b[273]), .Z(p[273]) );
  XOR2D0 C5874 ( .A1(a[274]), .A2(b[274]), .Z(p[274]) );
  XOR2D0 C5873 ( .A1(a[275]), .A2(b[275]), .Z(p[275]) );
  XOR2D0 C5872 ( .A1(a[276]), .A2(b[276]), .Z(p[276]) );
  XOR2D0 C5871 ( .A1(a[277]), .A2(b[277]), .Z(p[277]) );
  XOR2D0 C5870 ( .A1(a[278]), .A2(b[278]), .Z(p[278]) );
  XOR2D0 C5869 ( .A1(a[279]), .A2(b[279]), .Z(p[279]) );
  XOR2D0 C5868 ( .A1(a[280]), .A2(b[280]), .Z(p[280]) );
  XOR2D0 C5867 ( .A1(a[281]), .A2(b[281]), .Z(p[281]) );
  XOR2D0 C5866 ( .A1(a[282]), .A2(b[282]), .Z(p[282]) );
  XOR2D0 C5865 ( .A1(a[283]), .A2(b[283]), .Z(p[283]) );
  XOR2D0 C5864 ( .A1(a[284]), .A2(b[284]), .Z(p[284]) );
  XOR2D0 C5863 ( .A1(a[285]), .A2(b[285]), .Z(p[285]) );
  XOR2D0 C5862 ( .A1(a[286]), .A2(b[286]), .Z(p[286]) );
  XOR2D0 C5861 ( .A1(a[287]), .A2(b[287]), .Z(p[287]) );
  XOR2D0 C5860 ( .A1(a[288]), .A2(b[288]), .Z(p[288]) );
  XOR2D0 C5859 ( .A1(a[289]), .A2(b[289]), .Z(p[289]) );
  XOR2D0 C5858 ( .A1(a[290]), .A2(b[290]), .Z(p[290]) );
  XOR2D0 C5857 ( .A1(a[291]), .A2(b[291]), .Z(p[291]) );
  XOR2D0 C5856 ( .A1(a[292]), .A2(b[292]), .Z(p[292]) );
  XOR2D0 C5855 ( .A1(a[293]), .A2(b[293]), .Z(p[293]) );
  XOR2D0 C5854 ( .A1(a[294]), .A2(b[294]), .Z(p[294]) );
  XOR2D0 C5853 ( .A1(a[295]), .A2(b[295]), .Z(p[295]) );
  XOR2D0 C5852 ( .A1(a[296]), .A2(b[296]), .Z(p[296]) );
  XOR2D0 C5851 ( .A1(a[297]), .A2(b[297]), .Z(p[297]) );
  XOR2D0 C5850 ( .A1(a[298]), .A2(b[298]), .Z(p[298]) );
  XOR2D0 C5849 ( .A1(a[299]), .A2(b[299]), .Z(p[299]) );
  XOR2D0 C5848 ( .A1(a[300]), .A2(b[300]), .Z(p[300]) );
  XOR2D0 C5847 ( .A1(a[301]), .A2(b[301]), .Z(p[301]) );
  XOR2D0 C5846 ( .A1(a[302]), .A2(b[302]), .Z(p[302]) );
  XOR2D0 C5845 ( .A1(a[303]), .A2(b[303]), .Z(p[303]) );
  XOR2D0 C5844 ( .A1(a[304]), .A2(b[304]), .Z(p[304]) );
  XOR2D0 C5843 ( .A1(a[305]), .A2(b[305]), .Z(p[305]) );
  XOR2D0 C5842 ( .A1(a[306]), .A2(b[306]), .Z(p[306]) );
  XOR2D0 C5841 ( .A1(a[307]), .A2(b[307]), .Z(p[307]) );
  XOR2D0 C5840 ( .A1(a[308]), .A2(b[308]), .Z(p[308]) );
  XOR2D0 C5839 ( .A1(a[309]), .A2(b[309]), .Z(p[309]) );
  XOR2D0 C5838 ( .A1(a[310]), .A2(b[310]), .Z(p[310]) );
  XOR2D0 C5837 ( .A1(a[311]), .A2(b[311]), .Z(p[311]) );
  XOR2D0 C5836 ( .A1(a[312]), .A2(b[312]), .Z(p[312]) );
  XOR2D0 C5835 ( .A1(a[313]), .A2(b[313]), .Z(p[313]) );
  XOR2D0 C5834 ( .A1(a[314]), .A2(b[314]), .Z(p[314]) );
  XOR2D0 C5833 ( .A1(a[315]), .A2(b[315]), .Z(p[315]) );
  XOR2D0 C5832 ( .A1(a[316]), .A2(b[316]), .Z(p[316]) );
  XOR2D0 C5831 ( .A1(a[317]), .A2(b[317]), .Z(p[317]) );
  XOR2D0 C5830 ( .A1(a[318]), .A2(b[318]), .Z(p[318]) );
  XOR2D0 C5829 ( .A1(a[319]), .A2(b[319]), .Z(p[319]) );
  XOR2D0 C5828 ( .A1(a[320]), .A2(b[320]), .Z(p[320]) );
  XOR2D0 C5827 ( .A1(a[321]), .A2(b[321]), .Z(p[321]) );
  XOR2D0 C5826 ( .A1(a[322]), .A2(b[322]), .Z(p[322]) );
  XOR2D0 C5825 ( .A1(a[323]), .A2(b[323]), .Z(p[323]) );
  XOR2D0 C5824 ( .A1(a[324]), .A2(b[324]), .Z(p[324]) );
  XOR2D0 C5823 ( .A1(a[325]), .A2(b[325]), .Z(p[325]) );
  XOR2D0 C5822 ( .A1(a[326]), .A2(b[326]), .Z(p[326]) );
  XOR2D0 C5821 ( .A1(a[327]), .A2(b[327]), .Z(p[327]) );
  XOR2D0 C5820 ( .A1(a[328]), .A2(b[328]), .Z(p[328]) );
  XOR2D0 C5819 ( .A1(a[329]), .A2(b[329]), .Z(p[329]) );
  XOR2D0 C5818 ( .A1(a[330]), .A2(b[330]), .Z(p[330]) );
  XOR2D0 C5817 ( .A1(a[331]), .A2(b[331]), .Z(p[331]) );
  XOR2D0 C5816 ( .A1(a[332]), .A2(b[332]), .Z(p[332]) );
  XOR2D0 C5815 ( .A1(a[333]), .A2(b[333]), .Z(p[333]) );
  XOR2D0 C5814 ( .A1(a[334]), .A2(b[334]), .Z(p[334]) );
  XOR2D0 C5813 ( .A1(a[335]), .A2(b[335]), .Z(p[335]) );
  XOR2D0 C5812 ( .A1(a[336]), .A2(b[336]), .Z(p[336]) );
  XOR2D0 C5811 ( .A1(a[337]), .A2(b[337]), .Z(p[337]) );
  XOR2D0 C5810 ( .A1(a[338]), .A2(b[338]), .Z(p[338]) );
  XOR2D0 C5809 ( .A1(a[339]), .A2(b[339]), .Z(p[339]) );
  XOR2D0 C5808 ( .A1(a[340]), .A2(b[340]), .Z(p[340]) );
  XOR2D0 C5807 ( .A1(a[341]), .A2(b[341]), .Z(p[341]) );
  XOR2D0 C5806 ( .A1(a[342]), .A2(b[342]), .Z(p[342]) );
  XOR2D0 C5805 ( .A1(a[343]), .A2(b[343]), .Z(p[343]) );
  XOR2D0 C5804 ( .A1(a[344]), .A2(b[344]), .Z(p[344]) );
  XOR2D0 C5803 ( .A1(a[345]), .A2(b[345]), .Z(p[345]) );
  XOR2D0 C5802 ( .A1(a[346]), .A2(b[346]), .Z(p[346]) );
  XOR2D0 C5801 ( .A1(a[347]), .A2(b[347]), .Z(p[347]) );
  XOR2D0 C5800 ( .A1(a[348]), .A2(b[348]), .Z(p[348]) );
  XOR2D0 C5799 ( .A1(a[349]), .A2(b[349]), .Z(p[349]) );
  XOR2D0 C5798 ( .A1(a[350]), .A2(b[350]), .Z(p[350]) );
  XOR2D0 C5797 ( .A1(a[351]), .A2(b[351]), .Z(p[351]) );
  XOR2D0 C5796 ( .A1(a[352]), .A2(b[352]), .Z(p[352]) );
  XOR2D0 C5795 ( .A1(a[353]), .A2(b[353]), .Z(p[353]) );
  XOR2D0 C5794 ( .A1(a[354]), .A2(b[354]), .Z(p[354]) );
  XOR2D0 C5793 ( .A1(a[355]), .A2(b[355]), .Z(p[355]) );
  XOR2D0 C5792 ( .A1(a[356]), .A2(b[356]), .Z(p[356]) );
  XOR2D0 C5791 ( .A1(a[357]), .A2(b[357]), .Z(p[357]) );
  XOR2D0 C5790 ( .A1(a[358]), .A2(b[358]), .Z(p[358]) );
  XOR2D0 C5789 ( .A1(a[359]), .A2(b[359]), .Z(p[359]) );
  XOR2D0 C5788 ( .A1(a[360]), .A2(b[360]), .Z(p[360]) );
  XOR2D0 C5787 ( .A1(a[361]), .A2(b[361]), .Z(p[361]) );
  XOR2D0 C5786 ( .A1(a[362]), .A2(b[362]), .Z(p[362]) );
  XOR2D0 C5785 ( .A1(a[363]), .A2(b[363]), .Z(p[363]) );
  XOR2D0 C5784 ( .A1(a[364]), .A2(b[364]), .Z(p[364]) );
  XOR2D0 C5783 ( .A1(a[365]), .A2(b[365]), .Z(p[365]) );
  XOR2D0 C5782 ( .A1(a[366]), .A2(b[366]), .Z(p[366]) );
  XOR2D0 C5781 ( .A1(a[367]), .A2(b[367]), .Z(p[367]) );
  XOR2D0 C5780 ( .A1(a[368]), .A2(b[368]), .Z(p[368]) );
  XOR2D0 C5779 ( .A1(a[369]), .A2(b[369]), .Z(p[369]) );
  XOR2D0 C5778 ( .A1(a[370]), .A2(b[370]), .Z(p[370]) );
  XOR2D0 C5777 ( .A1(a[371]), .A2(b[371]), .Z(p[371]) );
  XOR2D0 C5776 ( .A1(a[372]), .A2(b[372]), .Z(p[372]) );
  XOR2D0 C5775 ( .A1(a[373]), .A2(b[373]), .Z(p[373]) );
  XOR2D0 C5774 ( .A1(a[374]), .A2(b[374]), .Z(p[374]) );
  XOR2D0 C5773 ( .A1(a[375]), .A2(b[375]), .Z(p[375]) );
  XOR2D0 C5772 ( .A1(a[376]), .A2(b[376]), .Z(p[376]) );
  XOR2D0 C5771 ( .A1(a[377]), .A2(b[377]), .Z(p[377]) );
  XOR2D0 C5770 ( .A1(a[378]), .A2(b[378]), .Z(p[378]) );
  XOR2D0 C5769 ( .A1(a[379]), .A2(b[379]), .Z(p[379]) );
  XOR2D0 C5768 ( .A1(a[380]), .A2(b[380]), .Z(p[380]) );
  XOR2D0 C5767 ( .A1(a[381]), .A2(b[381]), .Z(p[381]) );
  XOR2D0 C5766 ( .A1(a[382]), .A2(b[382]), .Z(p[382]) );
  XOR2D0 C5765 ( .A1(a[383]), .A2(b[383]), .Z(p[383]) );
  XOR2D0 C5764 ( .A1(a[384]), .A2(b[384]), .Z(p[384]) );
  XOR2D0 C5763 ( .A1(a[385]), .A2(b[385]), .Z(p[385]) );
  XOR2D0 C5762 ( .A1(a[386]), .A2(b[386]), .Z(p[386]) );
  XOR2D0 C5761 ( .A1(a[387]), .A2(b[387]), .Z(p[387]) );
  XOR2D0 C5760 ( .A1(a[388]), .A2(b[388]), .Z(p[388]) );
  XOR2D0 C5759 ( .A1(a[389]), .A2(b[389]), .Z(p[389]) );
  XOR2D0 C5758 ( .A1(a[390]), .A2(b[390]), .Z(p[390]) );
  XOR2D0 C5757 ( .A1(a[391]), .A2(b[391]), .Z(p[391]) );
  XOR2D0 C5756 ( .A1(a[392]), .A2(b[392]), .Z(p[392]) );
  XOR2D0 C5755 ( .A1(a[393]), .A2(b[393]), .Z(p[393]) );
  XOR2D0 C5754 ( .A1(a[394]), .A2(b[394]), .Z(p[394]) );
  XOR2D0 C5753 ( .A1(a[395]), .A2(b[395]), .Z(p[395]) );
  XOR2D0 C5752 ( .A1(a[396]), .A2(b[396]), .Z(p[396]) );
  XOR2D0 C5751 ( .A1(a[397]), .A2(b[397]), .Z(p[397]) );
  XOR2D0 C5750 ( .A1(a[398]), .A2(b[398]), .Z(p[398]) );
  XOR2D0 C5749 ( .A1(a[399]), .A2(b[399]), .Z(p[399]) );
  XOR2D0 C5748 ( .A1(a[400]), .A2(b[400]), .Z(p[400]) );
  XOR2D0 C5747 ( .A1(a[401]), .A2(b[401]), .Z(p[401]) );
  XOR2D0 C5746 ( .A1(a[402]), .A2(b[402]), .Z(p[402]) );
  XOR2D0 C5745 ( .A1(a[403]), .A2(b[403]), .Z(p[403]) );
  XOR2D0 C5744 ( .A1(a[404]), .A2(b[404]), .Z(p[404]) );
  XOR2D0 C5743 ( .A1(a[405]), .A2(b[405]), .Z(p[405]) );
  XOR2D0 C5742 ( .A1(a[406]), .A2(b[406]), .Z(p[406]) );
  XOR2D0 C5741 ( .A1(a[407]), .A2(b[407]), .Z(p[407]) );
  XOR2D0 C5740 ( .A1(a[408]), .A2(b[408]), .Z(p[408]) );
  XOR2D0 C5739 ( .A1(a[409]), .A2(b[409]), .Z(p[409]) );
  XOR2D0 C5738 ( .A1(a[410]), .A2(b[410]), .Z(p[410]) );
  XOR2D0 C5737 ( .A1(a[411]), .A2(b[411]), .Z(p[411]) );
  XOR2D0 C5736 ( .A1(a[412]), .A2(b[412]), .Z(p[412]) );
  XOR2D0 C5735 ( .A1(a[413]), .A2(b[413]), .Z(p[413]) );
  XOR2D0 C5734 ( .A1(a[414]), .A2(b[414]), .Z(p[414]) );
  XOR2D0 C5733 ( .A1(a[415]), .A2(b[415]), .Z(p[415]) );
  XOR2D0 C5732 ( .A1(a[416]), .A2(b[416]), .Z(p[416]) );
  XOR2D0 C5731 ( .A1(a[417]), .A2(b[417]), .Z(p[417]) );
  XOR2D0 C5730 ( .A1(a[418]), .A2(b[418]), .Z(p[418]) );
  XOR2D0 C5729 ( .A1(a[419]), .A2(b[419]), .Z(p[419]) );
  XOR2D0 C5728 ( .A1(a[420]), .A2(b[420]), .Z(p[420]) );
  XOR2D0 C5727 ( .A1(a[421]), .A2(b[421]), .Z(p[421]) );
  XOR2D0 C5726 ( .A1(a[422]), .A2(b[422]), .Z(p[422]) );
  XOR2D0 C5725 ( .A1(a[423]), .A2(b[423]), .Z(p[423]) );
  XOR2D0 C5724 ( .A1(a[424]), .A2(b[424]), .Z(p[424]) );
  XOR2D0 C5723 ( .A1(a[425]), .A2(b[425]), .Z(p[425]) );
  XOR2D0 C5722 ( .A1(a[426]), .A2(b[426]), .Z(p[426]) );
  XOR2D0 C5721 ( .A1(a[427]), .A2(b[427]), .Z(p[427]) );
  XOR2D0 C5720 ( .A1(a[428]), .A2(b[428]), .Z(p[428]) );
  XOR2D0 C5719 ( .A1(a[429]), .A2(b[429]), .Z(p[429]) );
  XOR2D0 C5718 ( .A1(a[430]), .A2(b[430]), .Z(p[430]) );
  XOR2D0 C5717 ( .A1(a[431]), .A2(b[431]), .Z(p[431]) );
  XOR2D0 C5716 ( .A1(a[432]), .A2(b[432]), .Z(p[432]) );
  XOR2D0 C5715 ( .A1(a[433]), .A2(b[433]), .Z(p[433]) );
  XOR2D0 C5714 ( .A1(a[434]), .A2(b[434]), .Z(p[434]) );
  XOR2D0 C5713 ( .A1(a[435]), .A2(b[435]), .Z(p[435]) );
  XOR2D0 C5712 ( .A1(a[436]), .A2(b[436]), .Z(p[436]) );
  XOR2D0 C5711 ( .A1(a[437]), .A2(b[437]), .Z(p[437]) );
  XOR2D0 C5710 ( .A1(a[438]), .A2(b[438]), .Z(p[438]) );
  XOR2D0 C5709 ( .A1(a[439]), .A2(b[439]), .Z(p[439]) );
  XOR2D0 C5708 ( .A1(a[440]), .A2(b[440]), .Z(p[440]) );
  XOR2D0 C5707 ( .A1(a[441]), .A2(b[441]), .Z(p[441]) );
  XOR2D0 C5706 ( .A1(a[442]), .A2(b[442]), .Z(p[442]) );
  XOR2D0 C5705 ( .A1(a[443]), .A2(b[443]), .Z(p[443]) );
  XOR2D0 C5704 ( .A1(a[444]), .A2(b[444]), .Z(p[444]) );
  XOR2D0 C5703 ( .A1(a[445]), .A2(b[445]), .Z(p[445]) );
  XOR2D0 C5702 ( .A1(a[446]), .A2(b[446]), .Z(p[446]) );
  XOR2D0 C5701 ( .A1(a[447]), .A2(b[447]), .Z(p[447]) );
  XOR2D0 C5700 ( .A1(a[448]), .A2(b[448]), .Z(p[448]) );
  XOR2D0 C5699 ( .A1(a[449]), .A2(b[449]), .Z(p[449]) );
  XOR2D0 C5698 ( .A1(a[450]), .A2(b[450]), .Z(p[450]) );
  XOR2D0 C5697 ( .A1(a[451]), .A2(b[451]), .Z(p[451]) );
  XOR2D0 C5696 ( .A1(a[452]), .A2(b[452]), .Z(p[452]) );
  XOR2D0 C5695 ( .A1(a[453]), .A2(b[453]), .Z(p[453]) );
  XOR2D0 C5694 ( .A1(a[454]), .A2(b[454]), .Z(p[454]) );
  XOR2D0 C5693 ( .A1(a[455]), .A2(b[455]), .Z(p[455]) );
  XOR2D0 C5692 ( .A1(a[456]), .A2(b[456]), .Z(p[456]) );
  XOR2D0 C5691 ( .A1(a[457]), .A2(b[457]), .Z(p[457]) );
  XOR2D0 C5690 ( .A1(a[458]), .A2(b[458]), .Z(p[458]) );
  XOR2D0 C5689 ( .A1(a[459]), .A2(b[459]), .Z(p[459]) );
  XOR2D0 C5688 ( .A1(a[460]), .A2(b[460]), .Z(p[460]) );
  XOR2D0 C5687 ( .A1(a[461]), .A2(b[461]), .Z(p[461]) );
  XOR2D0 C5686 ( .A1(a[462]), .A2(b[462]), .Z(p[462]) );
  XOR2D0 C5685 ( .A1(a[463]), .A2(b[463]), .Z(p[463]) );
  XOR2D0 C5684 ( .A1(a[464]), .A2(b[464]), .Z(p[464]) );
  XOR2D0 C5683 ( .A1(a[465]), .A2(b[465]), .Z(p[465]) );
  XOR2D0 C5682 ( .A1(a[466]), .A2(b[466]), .Z(p[466]) );
  XOR2D0 C5681 ( .A1(a[467]), .A2(b[467]), .Z(p[467]) );
  XOR2D0 C5680 ( .A1(a[468]), .A2(b[468]), .Z(p[468]) );
  XOR2D0 C5679 ( .A1(a[469]), .A2(b[469]), .Z(p[469]) );
  XOR2D0 C5678 ( .A1(a[470]), .A2(b[470]), .Z(p[470]) );
  XOR2D0 C5677 ( .A1(a[471]), .A2(b[471]), .Z(p[471]) );
  XOR2D0 C5676 ( .A1(a[472]), .A2(b[472]), .Z(p[472]) );
  XOR2D0 C5675 ( .A1(a[473]), .A2(b[473]), .Z(p[473]) );
  XOR2D0 C5674 ( .A1(a[474]), .A2(b[474]), .Z(p[474]) );
  XOR2D0 C5673 ( .A1(a[475]), .A2(b[475]), .Z(p[475]) );
  XOR2D0 C5672 ( .A1(a[476]), .A2(b[476]), .Z(p[476]) );
  XOR2D0 C5671 ( .A1(a[477]), .A2(b[477]), .Z(p[477]) );
  XOR2D0 C5670 ( .A1(a[478]), .A2(b[478]), .Z(p[478]) );
  XOR2D0 C5669 ( .A1(a[479]), .A2(b[479]), .Z(p[479]) );
  XOR2D0 C5668 ( .A1(a[480]), .A2(b[480]), .Z(p[480]) );
  XOR2D0 C5667 ( .A1(a[481]), .A2(b[481]), .Z(p[481]) );
  XOR2D0 C5666 ( .A1(a[482]), .A2(b[482]), .Z(p[482]) );
  XOR2D0 C5665 ( .A1(a[483]), .A2(b[483]), .Z(p[483]) );
  XOR2D0 C5664 ( .A1(a[484]), .A2(b[484]), .Z(p[484]) );
  XOR2D0 C5663 ( .A1(a[485]), .A2(b[485]), .Z(p[485]) );
  XOR2D0 C5662 ( .A1(a[486]), .A2(b[486]), .Z(p[486]) );
  XOR2D0 C5661 ( .A1(a[487]), .A2(b[487]), .Z(p[487]) );
  XOR2D0 C5660 ( .A1(a[488]), .A2(b[488]), .Z(p[488]) );
  XOR2D0 C5659 ( .A1(a[489]), .A2(b[489]), .Z(p[489]) );
  XOR2D0 C5658 ( .A1(a[490]), .A2(b[490]), .Z(p[490]) );
  XOR2D0 C5657 ( .A1(a[491]), .A2(b[491]), .Z(p[491]) );
  XOR2D0 C5656 ( .A1(a[492]), .A2(b[492]), .Z(p[492]) );
  XOR2D0 C5655 ( .A1(a[493]), .A2(b[493]), .Z(p[493]) );
  XOR2D0 C5654 ( .A1(a[494]), .A2(b[494]), .Z(p[494]) );
  XOR2D0 C5653 ( .A1(a[495]), .A2(b[495]), .Z(p[495]) );
  XOR2D0 C5652 ( .A1(a[496]), .A2(b[496]), .Z(p[496]) );
  XOR2D0 C5651 ( .A1(a[497]), .A2(b[497]), .Z(p[497]) );
  XOR2D0 C5650 ( .A1(a[498]), .A2(b[498]), .Z(p[498]) );
  XOR2D0 C5649 ( .A1(a[499]), .A2(b[499]), .Z(p[499]) );
  XOR2D0 C5648 ( .A1(a[500]), .A2(b[500]), .Z(p[500]) );
  XOR2D0 C5647 ( .A1(a[501]), .A2(b[501]), .Z(p[501]) );
  XOR2D0 C5646 ( .A1(a[502]), .A2(b[502]), .Z(p[502]) );
  XOR2D0 C5645 ( .A1(a[503]), .A2(b[503]), .Z(p[503]) );
  XOR2D0 C5644 ( .A1(a[504]), .A2(b[504]), .Z(p[504]) );
  XOR2D0 C5643 ( .A1(a[505]), .A2(b[505]), .Z(p[505]) );
  XOR2D0 C5642 ( .A1(a[506]), .A2(b[506]), .Z(p[506]) );
  XOR2D0 C5641 ( .A1(a[507]), .A2(b[507]), .Z(p[507]) );
  XOR2D0 C5640 ( .A1(a[508]), .A2(b[508]), .Z(p[508]) );
  XOR2D0 C5639 ( .A1(a[509]), .A2(b[509]), .Z(p[509]) );
  XOR2D0 C5638 ( .A1(a[510]), .A2(b[510]), .Z(p[510]) );
  XOR2D0 C5637 ( .A1(a[511]), .A2(b[511]), .Z(p[511]) );
  XOR2D0 C5636 ( .A1(a[512]), .A2(b[512]), .Z(p[512]) );
  XOR2D0 C5635 ( .A1(a[513]), .A2(b[513]), .Z(p[513]) );
  XOR2D0 C5634 ( .A1(a[514]), .A2(b[514]), .Z(p[514]) );
  XOR2D0 C5633 ( .A1(a[515]), .A2(b[515]), .Z(p[515]) );
  XOR2D0 C5632 ( .A1(a[516]), .A2(b[516]), .Z(p[516]) );
  XOR2D0 C5631 ( .A1(a[517]), .A2(b[517]), .Z(p[517]) );
  XOR2D0 C5630 ( .A1(a[518]), .A2(b[518]), .Z(p[518]) );
  XOR2D0 C5629 ( .A1(a[519]), .A2(b[519]), .Z(p[519]) );
  XOR2D0 C5628 ( .A1(a[520]), .A2(b[520]), .Z(p[520]) );
  XOR2D0 C5627 ( .A1(a[521]), .A2(b[521]), .Z(p[521]) );
  XOR2D0 C5626 ( .A1(a[522]), .A2(b[522]), .Z(p[522]) );
  XOR2D0 C5625 ( .A1(a[523]), .A2(b[523]), .Z(p[523]) );
  XOR2D0 C5624 ( .A1(a[524]), .A2(b[524]), .Z(p[524]) );
  XOR2D0 C5623 ( .A1(a[525]), .A2(b[525]), .Z(p[525]) );
  XOR2D0 C5622 ( .A1(a[526]), .A2(b[526]), .Z(p[526]) );
  XOR2D0 C5621 ( .A1(a[527]), .A2(b[527]), .Z(p[527]) );
  XOR2D0 C5620 ( .A1(a[528]), .A2(b[528]), .Z(p[528]) );
  XOR2D0 C5619 ( .A1(a[529]), .A2(b[529]), .Z(p[529]) );
  XOR2D0 C5618 ( .A1(a[530]), .A2(b[530]), .Z(p[530]) );
  XOR2D0 C5617 ( .A1(a[531]), .A2(b[531]), .Z(p[531]) );
  XOR2D0 C5616 ( .A1(a[532]), .A2(b[532]), .Z(p[532]) );
  XOR2D0 C5615 ( .A1(a[533]), .A2(b[533]), .Z(p[533]) );
  XOR2D0 C5614 ( .A1(a[534]), .A2(b[534]), .Z(p[534]) );
  XOR2D0 C5613 ( .A1(a[535]), .A2(b[535]), .Z(p[535]) );
  XOR2D0 C5612 ( .A1(a[536]), .A2(b[536]), .Z(p[536]) );
  XOR2D0 C5611 ( .A1(a[537]), .A2(b[537]), .Z(p[537]) );
  XOR2D0 C5610 ( .A1(a[538]), .A2(b[538]), .Z(p[538]) );
  XOR2D0 C5609 ( .A1(a[539]), .A2(b[539]), .Z(p[539]) );
  XOR2D0 C5608 ( .A1(a[540]), .A2(b[540]), .Z(p[540]) );
  XOR2D0 C5607 ( .A1(a[541]), .A2(b[541]), .Z(p[541]) );
  XOR2D0 C5606 ( .A1(a[542]), .A2(b[542]), .Z(p[542]) );
  XOR2D0 C5605 ( .A1(a[543]), .A2(b[543]), .Z(p[543]) );
  XOR2D0 C5604 ( .A1(a[544]), .A2(b[544]), .Z(p[544]) );
  XOR2D0 C5603 ( .A1(a[545]), .A2(b[545]), .Z(p[545]) );
  XOR2D0 C5602 ( .A1(a[546]), .A2(b[546]), .Z(p[546]) );
  XOR2D0 C5601 ( .A1(a[547]), .A2(b[547]), .Z(p[547]) );
  XOR2D0 C5600 ( .A1(a[548]), .A2(b[548]), .Z(p[548]) );
  XOR2D0 C5599 ( .A1(a[549]), .A2(b[549]), .Z(p[549]) );
  XOR2D0 C5598 ( .A1(a[550]), .A2(b[550]), .Z(p[550]) );
  XOR2D0 C5597 ( .A1(a[551]), .A2(b[551]), .Z(p[551]) );
  XOR2D0 C5596 ( .A1(a[552]), .A2(b[552]), .Z(p[552]) );
  XOR2D0 C5595 ( .A1(a[553]), .A2(b[553]), .Z(p[553]) );
  XOR2D0 C5594 ( .A1(a[554]), .A2(b[554]), .Z(p[554]) );
  XOR2D0 C5593 ( .A1(a[555]), .A2(b[555]), .Z(p[555]) );
  XOR2D0 C5592 ( .A1(a[556]), .A2(b[556]), .Z(p[556]) );
  XOR2D0 C5591 ( .A1(a[557]), .A2(b[557]), .Z(p[557]) );
  XOR2D0 C5590 ( .A1(a[558]), .A2(b[558]), .Z(p[558]) );
  XOR2D0 C5589 ( .A1(a[559]), .A2(b[559]), .Z(p[559]) );
  XOR2D0 C5588 ( .A1(a[560]), .A2(b[560]), .Z(p[560]) );
  XOR2D0 C5587 ( .A1(a[561]), .A2(b[561]), .Z(p[561]) );
  XOR2D0 C5586 ( .A1(a[562]), .A2(b[562]), .Z(p[562]) );
  XOR2D0 C5585 ( .A1(a[563]), .A2(b[563]), .Z(p[563]) );
  XOR2D0 C5584 ( .A1(a[564]), .A2(b[564]), .Z(p[564]) );
  XOR2D0 C5583 ( .A1(a[565]), .A2(b[565]), .Z(p[565]) );
  XOR2D0 C5582 ( .A1(a[566]), .A2(b[566]), .Z(p[566]) );
  XOR2D0 C5581 ( .A1(a[567]), .A2(b[567]), .Z(p[567]) );
  XOR2D0 C5580 ( .A1(a[568]), .A2(b[568]), .Z(p[568]) );
  XOR2D0 C5579 ( .A1(a[569]), .A2(b[569]), .Z(p[569]) );
  XOR2D0 C5578 ( .A1(a[570]), .A2(b[570]), .Z(p[570]) );
  XOR2D0 C5577 ( .A1(a[571]), .A2(b[571]), .Z(p[571]) );
  XOR2D0 C5576 ( .A1(a[572]), .A2(b[572]), .Z(p[572]) );
  XOR2D0 C5575 ( .A1(a[573]), .A2(b[573]), .Z(p[573]) );
  XOR2D0 C5574 ( .A1(a[574]), .A2(b[574]), .Z(p[574]) );
  XOR2D0 C5573 ( .A1(a[575]), .A2(b[575]), .Z(p[575]) );
  XOR2D0 C5572 ( .A1(a[576]), .A2(b[576]), .Z(p[576]) );
  XOR2D0 C5571 ( .A1(a[577]), .A2(b[577]), .Z(p[577]) );
  XOR2D0 C5570 ( .A1(a[578]), .A2(b[578]), .Z(p[578]) );
  XOR2D0 C5569 ( .A1(a[579]), .A2(b[579]), .Z(p[579]) );
  XOR2D0 C5568 ( .A1(a[580]), .A2(b[580]), .Z(p[580]) );
  XOR2D0 C5567 ( .A1(a[581]), .A2(b[581]), .Z(p[581]) );
  XOR2D0 C5566 ( .A1(a[582]), .A2(b[582]), .Z(p[582]) );
  XOR2D0 C5565 ( .A1(a[583]), .A2(b[583]), .Z(p[583]) );
  XOR2D0 C5564 ( .A1(a[584]), .A2(b[584]), .Z(p[584]) );
  XOR2D0 C5563 ( .A1(a[585]), .A2(b[585]), .Z(p[585]) );
  XOR2D0 C5562 ( .A1(a[586]), .A2(b[586]), .Z(p[586]) );
  XOR2D0 C5561 ( .A1(a[587]), .A2(b[587]), .Z(p[587]) );
  XOR2D0 C5560 ( .A1(a[588]), .A2(b[588]), .Z(p[588]) );
  XOR2D0 C5559 ( .A1(a[589]), .A2(b[589]), .Z(p[589]) );
  XOR2D0 C5558 ( .A1(a[590]), .A2(b[590]), .Z(p[590]) );
  XOR2D0 C5557 ( .A1(a[591]), .A2(b[591]), .Z(p[591]) );
  XOR2D0 C5556 ( .A1(a[592]), .A2(b[592]), .Z(p[592]) );
  XOR2D0 C5555 ( .A1(a[593]), .A2(b[593]), .Z(p[593]) );
  XOR2D0 C5554 ( .A1(a[594]), .A2(b[594]), .Z(p[594]) );
  XOR2D0 C5553 ( .A1(a[595]), .A2(b[595]), .Z(p[595]) );
  XOR2D0 C5552 ( .A1(a[596]), .A2(b[596]), .Z(p[596]) );
  XOR2D0 C5551 ( .A1(a[597]), .A2(b[597]), .Z(p[597]) );
  XOR2D0 C5550 ( .A1(a[598]), .A2(b[598]), .Z(p[598]) );
  XOR2D0 C5549 ( .A1(a[599]), .A2(b[599]), .Z(p[599]) );
  XOR2D0 C5548 ( .A1(a[600]), .A2(b[600]), .Z(p[600]) );
  XOR2D0 C5547 ( .A1(a[601]), .A2(b[601]), .Z(p[601]) );
  XOR2D0 C5546 ( .A1(a[602]), .A2(b[602]), .Z(p[602]) );
  XOR2D0 C5545 ( .A1(a[603]), .A2(b[603]), .Z(p[603]) );
  XOR2D0 C5544 ( .A1(a[604]), .A2(b[604]), .Z(p[604]) );
  XOR2D0 C5543 ( .A1(a[605]), .A2(b[605]), .Z(p[605]) );
  XOR2D0 C5542 ( .A1(a[606]), .A2(b[606]), .Z(p[606]) );
  XOR2D0 C5541 ( .A1(a[607]), .A2(b[607]), .Z(p[607]) );
  XOR2D0 C5540 ( .A1(a[608]), .A2(b[608]), .Z(p[608]) );
  XOR2D0 C5539 ( .A1(a[609]), .A2(b[609]), .Z(p[609]) );
  XOR2D0 C5538 ( .A1(a[610]), .A2(b[610]), .Z(p[610]) );
  XOR2D0 C5537 ( .A1(a[611]), .A2(b[611]), .Z(p[611]) );
  XOR2D0 C5536 ( .A1(a[612]), .A2(b[612]), .Z(p[612]) );
  XOR2D0 C5535 ( .A1(a[613]), .A2(b[613]), .Z(p[613]) );
  XOR2D0 C5534 ( .A1(a[614]), .A2(b[614]), .Z(p[614]) );
  XOR2D0 C5533 ( .A1(a[615]), .A2(b[615]), .Z(p[615]) );
  XOR2D0 C5532 ( .A1(a[616]), .A2(b[616]), .Z(p[616]) );
  XOR2D0 C5531 ( .A1(a[617]), .A2(b[617]), .Z(p[617]) );
  XOR2D0 C5530 ( .A1(a[618]), .A2(b[618]), .Z(p[618]) );
  XOR2D0 C5529 ( .A1(a[619]), .A2(b[619]), .Z(p[619]) );
  XOR2D0 C5528 ( .A1(a[620]), .A2(b[620]), .Z(p[620]) );
  XOR2D0 C5527 ( .A1(a[621]), .A2(b[621]), .Z(p[621]) );
  XOR2D0 C5526 ( .A1(a[622]), .A2(b[622]), .Z(p[622]) );
  XOR2D0 C5525 ( .A1(a[623]), .A2(b[623]), .Z(p[623]) );
  XOR2D0 C5524 ( .A1(a[624]), .A2(b[624]), .Z(p[624]) );
  XOR2D0 C5523 ( .A1(a[625]), .A2(b[625]), .Z(p[625]) );
  XOR2D0 C5522 ( .A1(a[626]), .A2(b[626]), .Z(p[626]) );
  XOR2D0 C5521 ( .A1(a[627]), .A2(b[627]), .Z(p[627]) );
  XOR2D0 C5520 ( .A1(a[628]), .A2(b[628]), .Z(p[628]) );
  XOR2D0 C5519 ( .A1(a[629]), .A2(b[629]), .Z(p[629]) );
  XOR2D0 C5518 ( .A1(a[630]), .A2(b[630]), .Z(p[630]) );
  XOR2D0 C5517 ( .A1(a[631]), .A2(b[631]), .Z(p[631]) );
  XOR2D0 C5516 ( .A1(a[632]), .A2(b[632]), .Z(p[632]) );
  XOR2D0 C5515 ( .A1(a[633]), .A2(b[633]), .Z(p[633]) );
  XOR2D0 C5514 ( .A1(a[634]), .A2(b[634]), .Z(p[634]) );
  XOR2D0 C5513 ( .A1(a[635]), .A2(b[635]), .Z(p[635]) );
  XOR2D0 C5512 ( .A1(a[636]), .A2(b[636]), .Z(p[636]) );
  XOR2D0 C5511 ( .A1(a[637]), .A2(b[637]), .Z(p[637]) );
  XOR2D0 C5510 ( .A1(a[638]), .A2(b[638]), .Z(p[638]) );
  XOR2D0 C5509 ( .A1(a[639]), .A2(b[639]), .Z(p[639]) );
  XOR2D0 C5508 ( .A1(a[640]), .A2(b[640]), .Z(p[640]) );
  XOR2D0 C5507 ( .A1(a[641]), .A2(b[641]), .Z(p[641]) );
  XOR2D0 C5506 ( .A1(a[642]), .A2(b[642]), .Z(p[642]) );
  XOR2D0 C5505 ( .A1(a[643]), .A2(b[643]), .Z(p[643]) );
  XOR2D0 C5504 ( .A1(a[644]), .A2(b[644]), .Z(p[644]) );
  XOR2D0 C5503 ( .A1(a[645]), .A2(b[645]), .Z(p[645]) );
  XOR2D0 C5502 ( .A1(a[646]), .A2(b[646]), .Z(p[646]) );
  XOR2D0 C5501 ( .A1(a[647]), .A2(b[647]), .Z(p[647]) );
  XOR2D0 C5500 ( .A1(a[648]), .A2(b[648]), .Z(p[648]) );
  XOR2D0 C5499 ( .A1(a[649]), .A2(b[649]), .Z(p[649]) );
  XOR2D0 C5498 ( .A1(a[650]), .A2(b[650]), .Z(p[650]) );
  XOR2D0 C5497 ( .A1(a[651]), .A2(b[651]), .Z(p[651]) );
  XOR2D0 C5496 ( .A1(a[652]), .A2(b[652]), .Z(p[652]) );
  XOR2D0 C5495 ( .A1(a[653]), .A2(b[653]), .Z(p[653]) );
  XOR2D0 C5494 ( .A1(a[654]), .A2(b[654]), .Z(p[654]) );
  XOR2D0 C5493 ( .A1(a[655]), .A2(b[655]), .Z(p[655]) );
  XOR2D0 C5492 ( .A1(a[656]), .A2(b[656]), .Z(p[656]) );
  XOR2D0 C5491 ( .A1(a[657]), .A2(b[657]), .Z(p[657]) );
  XOR2D0 C5490 ( .A1(a[658]), .A2(b[658]), .Z(p[658]) );
  XOR2D0 C5489 ( .A1(a[659]), .A2(b[659]), .Z(p[659]) );
  XOR2D0 C5488 ( .A1(a[660]), .A2(b[660]), .Z(p[660]) );
  XOR2D0 C5487 ( .A1(a[661]), .A2(b[661]), .Z(p[661]) );
  XOR2D0 C5486 ( .A1(a[662]), .A2(b[662]), .Z(p[662]) );
  XOR2D0 C5485 ( .A1(a[663]), .A2(b[663]), .Z(p[663]) );
  XOR2D0 C5484 ( .A1(a[664]), .A2(b[664]), .Z(p[664]) );
  XOR2D0 C5483 ( .A1(a[665]), .A2(b[665]), .Z(p[665]) );
  XOR2D0 C5482 ( .A1(a[666]), .A2(b[666]), .Z(p[666]) );
  XOR2D0 C5481 ( .A1(a[667]), .A2(b[667]), .Z(p[667]) );
  XOR2D0 C5480 ( .A1(a[668]), .A2(b[668]), .Z(p[668]) );
  XOR2D0 C5479 ( .A1(a[669]), .A2(b[669]), .Z(p[669]) );
  XOR2D0 C5478 ( .A1(a[670]), .A2(b[670]), .Z(p[670]) );
  XOR2D0 C5477 ( .A1(a[671]), .A2(b[671]), .Z(p[671]) );
  XOR2D0 C5476 ( .A1(a[672]), .A2(b[672]), .Z(p[672]) );
  XOR2D0 C5475 ( .A1(a[673]), .A2(b[673]), .Z(p[673]) );
  XOR2D0 C5474 ( .A1(a[674]), .A2(b[674]), .Z(p[674]) );
  XOR2D0 C5473 ( .A1(a[675]), .A2(b[675]), .Z(p[675]) );
  XOR2D0 C5472 ( .A1(a[676]), .A2(b[676]), .Z(p[676]) );
  XOR2D0 C5471 ( .A1(a[677]), .A2(b[677]), .Z(p[677]) );
  XOR2D0 C5470 ( .A1(a[678]), .A2(b[678]), .Z(p[678]) );
  XOR2D0 C5469 ( .A1(a[679]), .A2(b[679]), .Z(p[679]) );
  XOR2D0 C5468 ( .A1(a[680]), .A2(b[680]), .Z(p[680]) );
  XOR2D0 C5467 ( .A1(a[681]), .A2(b[681]), .Z(p[681]) );
  XOR2D0 C5466 ( .A1(a[682]), .A2(b[682]), .Z(p[682]) );
  XOR2D0 C5465 ( .A1(a[683]), .A2(b[683]), .Z(p[683]) );
  XOR2D0 C5464 ( .A1(a[684]), .A2(b[684]), .Z(p[684]) );
  XOR2D0 C5463 ( .A1(a[685]), .A2(b[685]), .Z(p[685]) );
  XOR2D0 C5462 ( .A1(a[686]), .A2(b[686]), .Z(p[686]) );
  XOR2D0 C5461 ( .A1(a[687]), .A2(b[687]), .Z(p[687]) );
  XOR2D0 C5460 ( .A1(a[688]), .A2(b[688]), .Z(p[688]) );
  XOR2D0 C5459 ( .A1(a[689]), .A2(b[689]), .Z(p[689]) );
  XOR2D0 C5458 ( .A1(a[690]), .A2(b[690]), .Z(p[690]) );
  XOR2D0 C5457 ( .A1(a[691]), .A2(b[691]), .Z(p[691]) );
  XOR2D0 C5456 ( .A1(a[692]), .A2(b[692]), .Z(p[692]) );
  XOR2D0 C5455 ( .A1(a[693]), .A2(b[693]), .Z(p[693]) );
  XOR2D0 C5454 ( .A1(a[694]), .A2(b[694]), .Z(p[694]) );
  XOR2D0 C5453 ( .A1(a[695]), .A2(b[695]), .Z(p[695]) );
  XOR2D0 C5452 ( .A1(a[696]), .A2(b[696]), .Z(p[696]) );
  XOR2D0 C5451 ( .A1(a[697]), .A2(b[697]), .Z(p[697]) );
  XOR2D0 C5450 ( .A1(a[698]), .A2(b[698]), .Z(p[698]) );
  XOR2D0 C5449 ( .A1(a[699]), .A2(b[699]), .Z(p[699]) );
  XOR2D0 C5448 ( .A1(a[700]), .A2(b[700]), .Z(p[700]) );
  XOR2D0 C5447 ( .A1(a[701]), .A2(b[701]), .Z(p[701]) );
  XOR2D0 C5446 ( .A1(a[702]), .A2(b[702]), .Z(p[702]) );
  XOR2D0 C5445 ( .A1(a[703]), .A2(b[703]), .Z(p[703]) );
  XOR2D0 C5444 ( .A1(a[704]), .A2(b[704]), .Z(p[704]) );
  XOR2D0 C5443 ( .A1(a[705]), .A2(b[705]), .Z(p[705]) );
  XOR2D0 C5442 ( .A1(a[706]), .A2(b[706]), .Z(p[706]) );
  XOR2D0 C5441 ( .A1(a[707]), .A2(b[707]), .Z(p[707]) );
  XOR2D0 C5440 ( .A1(a[708]), .A2(b[708]), .Z(p[708]) );
  XOR2D0 C5439 ( .A1(a[709]), .A2(b[709]), .Z(p[709]) );
  XOR2D0 C5438 ( .A1(a[710]), .A2(b[710]), .Z(p[710]) );
  XOR2D0 C5437 ( .A1(a[711]), .A2(b[711]), .Z(p[711]) );
  XOR2D0 C5436 ( .A1(a[712]), .A2(b[712]), .Z(p[712]) );
  XOR2D0 C5435 ( .A1(a[713]), .A2(b[713]), .Z(p[713]) );
  XOR2D0 C5434 ( .A1(a[714]), .A2(b[714]), .Z(p[714]) );
  XOR2D0 C5433 ( .A1(a[715]), .A2(b[715]), .Z(p[715]) );
  XOR2D0 C5432 ( .A1(a[716]), .A2(b[716]), .Z(p[716]) );
  XOR2D0 C5431 ( .A1(a[717]), .A2(b[717]), .Z(p[717]) );
  XOR2D0 C5430 ( .A1(a[718]), .A2(b[718]), .Z(p[718]) );
  XOR2D0 C5429 ( .A1(a[719]), .A2(b[719]), .Z(p[719]) );
  XOR2D0 C5428 ( .A1(a[720]), .A2(b[720]), .Z(p[720]) );
  XOR2D0 C5427 ( .A1(a[721]), .A2(b[721]), .Z(p[721]) );
  XOR2D0 C5426 ( .A1(a[722]), .A2(b[722]), .Z(p[722]) );
  XOR2D0 C5425 ( .A1(a[723]), .A2(b[723]), .Z(p[723]) );
  XOR2D0 C5424 ( .A1(a[724]), .A2(b[724]), .Z(p[724]) );
  XOR2D0 C5423 ( .A1(a[725]), .A2(b[725]), .Z(p[725]) );
  XOR2D0 C5422 ( .A1(a[726]), .A2(b[726]), .Z(p[726]) );
  XOR2D0 C5421 ( .A1(a[727]), .A2(b[727]), .Z(p[727]) );
  XOR2D0 C5420 ( .A1(a[728]), .A2(b[728]), .Z(p[728]) );
  XOR2D0 C5419 ( .A1(a[729]), .A2(b[729]), .Z(p[729]) );
  XOR2D0 C5418 ( .A1(a[730]), .A2(b[730]), .Z(p[730]) );
  XOR2D0 C5417 ( .A1(a[731]), .A2(b[731]), .Z(p[731]) );
  XOR2D0 C5416 ( .A1(a[732]), .A2(b[732]), .Z(p[732]) );
  XOR2D0 C5415 ( .A1(a[733]), .A2(b[733]), .Z(p[733]) );
  XOR2D0 C5414 ( .A1(a[734]), .A2(b[734]), .Z(p[734]) );
  XOR2D0 C5413 ( .A1(a[735]), .A2(b[735]), .Z(p[735]) );
  XOR2D0 C5412 ( .A1(a[736]), .A2(b[736]), .Z(p[736]) );
  XOR2D0 C5411 ( .A1(a[737]), .A2(b[737]), .Z(p[737]) );
  XOR2D0 C5410 ( .A1(a[738]), .A2(b[738]), .Z(p[738]) );
  XOR2D0 C5409 ( .A1(a[739]), .A2(b[739]), .Z(p[739]) );
  XOR2D0 C5408 ( .A1(a[740]), .A2(b[740]), .Z(p[740]) );
  XOR2D0 C5407 ( .A1(a[741]), .A2(b[741]), .Z(p[741]) );
  XOR2D0 C5406 ( .A1(a[742]), .A2(b[742]), .Z(p[742]) );
  XOR2D0 C5405 ( .A1(a[743]), .A2(b[743]), .Z(p[743]) );
  XOR2D0 C5404 ( .A1(a[744]), .A2(b[744]), .Z(p[744]) );
  XOR2D0 C5403 ( .A1(a[745]), .A2(b[745]), .Z(p[745]) );
  XOR2D0 C5402 ( .A1(a[746]), .A2(b[746]), .Z(p[746]) );
  XOR2D0 C5401 ( .A1(a[747]), .A2(b[747]), .Z(p[747]) );
  XOR2D0 C5400 ( .A1(a[748]), .A2(b[748]), .Z(p[748]) );
  XOR2D0 C5399 ( .A1(a[749]), .A2(b[749]), .Z(p[749]) );
  XOR2D0 C5398 ( .A1(a[750]), .A2(b[750]), .Z(p[750]) );
  XOR2D0 C5397 ( .A1(a[751]), .A2(b[751]), .Z(p[751]) );
  XOR2D0 C5396 ( .A1(a[752]), .A2(b[752]), .Z(p[752]) );
  XOR2D0 C5395 ( .A1(a[753]), .A2(b[753]), .Z(p[753]) );
  XOR2D0 C5394 ( .A1(a[754]), .A2(b[754]), .Z(p[754]) );
  XOR2D0 C5393 ( .A1(a[755]), .A2(b[755]), .Z(p[755]) );
  XOR2D0 C5392 ( .A1(a[756]), .A2(b[756]), .Z(p[756]) );
  XOR2D0 C5391 ( .A1(a[757]), .A2(b[757]), .Z(p[757]) );
  XOR2D0 C5390 ( .A1(a[758]), .A2(b[758]), .Z(p[758]) );
  XOR2D0 C5389 ( .A1(a[759]), .A2(b[759]), .Z(p[759]) );
  XOR2D0 C5388 ( .A1(a[760]), .A2(b[760]), .Z(p[760]) );
  XOR2D0 C5387 ( .A1(a[761]), .A2(b[761]), .Z(p[761]) );
  XOR2D0 C5386 ( .A1(a[762]), .A2(b[762]), .Z(p[762]) );
  XOR2D0 C5385 ( .A1(a[763]), .A2(b[763]), .Z(p[763]) );
  XOR2D0 C5384 ( .A1(a[764]), .A2(b[764]), .Z(p[764]) );
  XOR2D0 C5383 ( .A1(a[765]), .A2(b[765]), .Z(p[765]) );
  XOR2D0 C5382 ( .A1(a[766]), .A2(b[766]), .Z(p[766]) );
  XOR2D0 C5381 ( .A1(a[767]), .A2(b[767]), .Z(p[767]) );
  XOR2D0 C5380 ( .A1(a[768]), .A2(b[768]), .Z(p[768]) );
  XOR2D0 C5379 ( .A1(a[769]), .A2(b[769]), .Z(p[769]) );
  XOR2D0 C5378 ( .A1(a[770]), .A2(b[770]), .Z(p[770]) );
  XOR2D0 C5377 ( .A1(a[771]), .A2(b[771]), .Z(p[771]) );
  XOR2D0 C5376 ( .A1(a[772]), .A2(b[772]), .Z(p[772]) );
  XOR2D0 C5375 ( .A1(a[773]), .A2(b[773]), .Z(p[773]) );
  XOR2D0 C5374 ( .A1(a[774]), .A2(b[774]), .Z(p[774]) );
  XOR2D0 C5373 ( .A1(a[775]), .A2(b[775]), .Z(p[775]) );
  XOR2D0 C5372 ( .A1(a[776]), .A2(b[776]), .Z(p[776]) );
  XOR2D0 C5371 ( .A1(a[777]), .A2(b[777]), .Z(p[777]) );
  XOR2D0 C5370 ( .A1(a[778]), .A2(b[778]), .Z(p[778]) );
  XOR2D0 C5369 ( .A1(a[779]), .A2(b[779]), .Z(p[779]) );
  XOR2D0 C5368 ( .A1(a[780]), .A2(b[780]), .Z(p[780]) );
  XOR2D0 C5367 ( .A1(a[781]), .A2(b[781]), .Z(p[781]) );
  XOR2D0 C5366 ( .A1(a[782]), .A2(b[782]), .Z(p[782]) );
  XOR2D0 C5365 ( .A1(a[783]), .A2(b[783]), .Z(p[783]) );
  XOR2D0 C5364 ( .A1(a[784]), .A2(b[784]), .Z(p[784]) );
  XOR2D0 C5363 ( .A1(a[785]), .A2(b[785]), .Z(p[785]) );
  XOR2D0 C5362 ( .A1(a[786]), .A2(b[786]), .Z(p[786]) );
  XOR2D0 C5361 ( .A1(a[787]), .A2(b[787]), .Z(p[787]) );
  XOR2D0 C5360 ( .A1(a[788]), .A2(b[788]), .Z(p[788]) );
  XOR2D0 C5359 ( .A1(a[789]), .A2(b[789]), .Z(p[789]) );
  XOR2D0 C5358 ( .A1(a[790]), .A2(b[790]), .Z(p[790]) );
  XOR2D0 C5357 ( .A1(a[791]), .A2(b[791]), .Z(p[791]) );
  XOR2D0 C5356 ( .A1(a[792]), .A2(b[792]), .Z(p[792]) );
  XOR2D0 C5355 ( .A1(a[793]), .A2(b[793]), .Z(p[793]) );
  XOR2D0 C5354 ( .A1(a[794]), .A2(b[794]), .Z(p[794]) );
  XOR2D0 C5353 ( .A1(a[795]), .A2(b[795]), .Z(p[795]) );
  XOR2D0 C5352 ( .A1(a[796]), .A2(b[796]), .Z(p[796]) );
  XOR2D0 C5351 ( .A1(a[797]), .A2(b[797]), .Z(p[797]) );
  XOR2D0 C5350 ( .A1(a[798]), .A2(b[798]), .Z(p[798]) );
  XOR2D0 C5349 ( .A1(a[799]), .A2(b[799]), .Z(p[799]) );
  XOR2D0 C5348 ( .A1(a[800]), .A2(b[800]), .Z(p[800]) );
  XOR2D0 C5347 ( .A1(a[801]), .A2(b[801]), .Z(p[801]) );
  XOR2D0 C5346 ( .A1(a[802]), .A2(b[802]), .Z(p[802]) );
  XOR2D0 C5345 ( .A1(a[803]), .A2(b[803]), .Z(p[803]) );
  XOR2D0 C5344 ( .A1(a[804]), .A2(b[804]), .Z(p[804]) );
  XOR2D0 C5343 ( .A1(a[805]), .A2(b[805]), .Z(p[805]) );
  XOR2D0 C5342 ( .A1(a[806]), .A2(b[806]), .Z(p[806]) );
  XOR2D0 C5341 ( .A1(a[807]), .A2(b[807]), .Z(p[807]) );
  XOR2D0 C5340 ( .A1(a[808]), .A2(b[808]), .Z(p[808]) );
  XOR2D0 C5339 ( .A1(a[809]), .A2(b[809]), .Z(p[809]) );
  XOR2D0 C5338 ( .A1(a[810]), .A2(b[810]), .Z(p[810]) );
  XOR2D0 C5337 ( .A1(a[811]), .A2(b[811]), .Z(p[811]) );
  XOR2D0 C5336 ( .A1(a[812]), .A2(b[812]), .Z(p[812]) );
  XOR2D0 C5335 ( .A1(a[813]), .A2(b[813]), .Z(p[813]) );
  XOR2D0 C5334 ( .A1(a[814]), .A2(b[814]), .Z(p[814]) );
  XOR2D0 C5333 ( .A1(a[815]), .A2(b[815]), .Z(p[815]) );
  XOR2D0 C5332 ( .A1(a[816]), .A2(b[816]), .Z(p[816]) );
  XOR2D0 C5331 ( .A1(a[817]), .A2(b[817]), .Z(p[817]) );
  XOR2D0 C5330 ( .A1(a[818]), .A2(b[818]), .Z(p[818]) );
  XOR2D0 C5329 ( .A1(a[819]), .A2(b[819]), .Z(p[819]) );
  XOR2D0 C5328 ( .A1(a[820]), .A2(b[820]), .Z(p[820]) );
  XOR2D0 C5327 ( .A1(a[821]), .A2(b[821]), .Z(p[821]) );
  XOR2D0 C5326 ( .A1(a[822]), .A2(b[822]), .Z(p[822]) );
  XOR2D0 C5325 ( .A1(a[823]), .A2(b[823]), .Z(p[823]) );
  XOR2D0 C5324 ( .A1(a[824]), .A2(b[824]), .Z(p[824]) );
  XOR2D0 C5323 ( .A1(a[825]), .A2(b[825]), .Z(p[825]) );
  XOR2D0 C5322 ( .A1(a[826]), .A2(b[826]), .Z(p[826]) );
  XOR2D0 C5321 ( .A1(a[827]), .A2(b[827]), .Z(p[827]) );
  XOR2D0 C5320 ( .A1(a[828]), .A2(b[828]), .Z(p[828]) );
  XOR2D0 C5319 ( .A1(a[829]), .A2(b[829]), .Z(p[829]) );
  XOR2D0 C5318 ( .A1(a[830]), .A2(b[830]), .Z(p[830]) );
  XOR2D0 C5317 ( .A1(a[831]), .A2(b[831]), .Z(p[831]) );
  XOR2D0 C5316 ( .A1(a[832]), .A2(b[832]), .Z(p[832]) );
  XOR2D0 C5315 ( .A1(a[833]), .A2(b[833]), .Z(p[833]) );
  XOR2D0 C5314 ( .A1(a[834]), .A2(b[834]), .Z(p[834]) );
  XOR2D0 C5313 ( .A1(a[835]), .A2(b[835]), .Z(p[835]) );
  XOR2D0 C5312 ( .A1(a[836]), .A2(b[836]), .Z(p[836]) );
  XOR2D0 C5311 ( .A1(a[837]), .A2(b[837]), .Z(p[837]) );
  XOR2D0 C5310 ( .A1(a[838]), .A2(b[838]), .Z(p[838]) );
  XOR2D0 C5309 ( .A1(a[839]), .A2(b[839]), .Z(p[839]) );
  XOR2D0 C5308 ( .A1(a[840]), .A2(b[840]), .Z(p[840]) );
  XOR2D0 C5307 ( .A1(a[841]), .A2(b[841]), .Z(p[841]) );
  XOR2D0 C5306 ( .A1(a[842]), .A2(b[842]), .Z(p[842]) );
  XOR2D0 C5305 ( .A1(a[843]), .A2(b[843]), .Z(p[843]) );
  XOR2D0 C5304 ( .A1(a[844]), .A2(b[844]), .Z(p[844]) );
  XOR2D0 C5303 ( .A1(a[845]), .A2(b[845]), .Z(p[845]) );
  XOR2D0 C5302 ( .A1(a[846]), .A2(b[846]), .Z(p[846]) );
  XOR2D0 C5301 ( .A1(a[847]), .A2(b[847]), .Z(p[847]) );
  XOR2D0 C5300 ( .A1(a[848]), .A2(b[848]), .Z(p[848]) );
  XOR2D0 C5299 ( .A1(a[849]), .A2(b[849]), .Z(p[849]) );
  XOR2D0 C5298 ( .A1(a[850]), .A2(b[850]), .Z(p[850]) );
  XOR2D0 C5297 ( .A1(a[851]), .A2(b[851]), .Z(p[851]) );
  XOR2D0 C5296 ( .A1(a[852]), .A2(b[852]), .Z(p[852]) );
  XOR2D0 C5295 ( .A1(a[853]), .A2(b[853]), .Z(p[853]) );
  XOR2D0 C5294 ( .A1(a[854]), .A2(b[854]), .Z(p[854]) );
  XOR2D0 C5293 ( .A1(a[855]), .A2(b[855]), .Z(p[855]) );
  XOR2D0 C5292 ( .A1(a[856]), .A2(b[856]), .Z(p[856]) );
  XOR2D0 C5291 ( .A1(a[857]), .A2(b[857]), .Z(p[857]) );
  XOR2D0 C5290 ( .A1(a[858]), .A2(b[858]), .Z(p[858]) );
  XOR2D0 C5289 ( .A1(a[859]), .A2(b[859]), .Z(p[859]) );
  XOR2D0 C5288 ( .A1(a[860]), .A2(b[860]), .Z(p[860]) );
  XOR2D0 C5287 ( .A1(a[861]), .A2(b[861]), .Z(p[861]) );
  XOR2D0 C5286 ( .A1(a[862]), .A2(b[862]), .Z(p[862]) );
  XOR2D0 C5285 ( .A1(a[863]), .A2(b[863]), .Z(p[863]) );
  XOR2D0 C5284 ( .A1(a[864]), .A2(b[864]), .Z(p[864]) );
  XOR2D0 C5283 ( .A1(a[865]), .A2(b[865]), .Z(p[865]) );
  XOR2D0 C5282 ( .A1(a[866]), .A2(b[866]), .Z(p[866]) );
  XOR2D0 C5281 ( .A1(a[867]), .A2(b[867]), .Z(p[867]) );
  XOR2D0 C5280 ( .A1(a[868]), .A2(b[868]), .Z(p[868]) );
  XOR2D0 C5279 ( .A1(a[869]), .A2(b[869]), .Z(p[869]) );
  XOR2D0 C5278 ( .A1(a[870]), .A2(b[870]), .Z(p[870]) );
  XOR2D0 C5277 ( .A1(a[871]), .A2(b[871]), .Z(p[871]) );
  XOR2D0 C5276 ( .A1(a[872]), .A2(b[872]), .Z(p[872]) );
  XOR2D0 C5275 ( .A1(a[873]), .A2(b[873]), .Z(p[873]) );
  XOR2D0 C5274 ( .A1(a[874]), .A2(b[874]), .Z(p[874]) );
  XOR2D0 C5273 ( .A1(a[875]), .A2(b[875]), .Z(p[875]) );
  XOR2D0 C5272 ( .A1(a[876]), .A2(b[876]), .Z(p[876]) );
  XOR2D0 C5271 ( .A1(a[877]), .A2(b[877]), .Z(p[877]) );
  XOR2D0 C5270 ( .A1(a[878]), .A2(b[878]), .Z(p[878]) );
  XOR2D0 C5269 ( .A1(a[879]), .A2(b[879]), .Z(p[879]) );
  XOR2D0 C5268 ( .A1(a[880]), .A2(b[880]), .Z(p[880]) );
  XOR2D0 C5267 ( .A1(a[881]), .A2(b[881]), .Z(p[881]) );
  XOR2D0 C5266 ( .A1(a[882]), .A2(b[882]), .Z(p[882]) );
  XOR2D0 C5265 ( .A1(a[883]), .A2(b[883]), .Z(p[883]) );
  XOR2D0 C5264 ( .A1(a[884]), .A2(b[884]), .Z(p[884]) );
  XOR2D0 C5263 ( .A1(a[885]), .A2(b[885]), .Z(p[885]) );
  XOR2D0 C5262 ( .A1(a[886]), .A2(b[886]), .Z(p[886]) );
  XOR2D0 C5261 ( .A1(a[887]), .A2(b[887]), .Z(p[887]) );
  XOR2D0 C5260 ( .A1(a[888]), .A2(b[888]), .Z(p[888]) );
  XOR2D0 C5259 ( .A1(a[889]), .A2(b[889]), .Z(p[889]) );
  XOR2D0 C5258 ( .A1(a[890]), .A2(b[890]), .Z(p[890]) );
  XOR2D0 C5257 ( .A1(a[891]), .A2(b[891]), .Z(p[891]) );
  XOR2D0 C5256 ( .A1(a[892]), .A2(b[892]), .Z(p[892]) );
  XOR2D0 C5255 ( .A1(a[893]), .A2(b[893]), .Z(p[893]) );
  XOR2D0 C5254 ( .A1(a[894]), .A2(b[894]), .Z(p[894]) );
  XOR2D0 C5253 ( .A1(a[895]), .A2(b[895]), .Z(p[895]) );
  XOR2D0 C5252 ( .A1(a[896]), .A2(b[896]), .Z(p[896]) );
  XOR2D0 C5251 ( .A1(a[897]), .A2(b[897]), .Z(p[897]) );
  XOR2D0 C5250 ( .A1(a[898]), .A2(b[898]), .Z(p[898]) );
  XOR2D0 C5249 ( .A1(a[899]), .A2(b[899]), .Z(p[899]) );
  XOR2D0 C5248 ( .A1(a[900]), .A2(b[900]), .Z(p[900]) );
  XOR2D0 C5247 ( .A1(a[901]), .A2(b[901]), .Z(p[901]) );
  XOR2D0 C5246 ( .A1(a[902]), .A2(b[902]), .Z(p[902]) );
  XOR2D0 C5245 ( .A1(a[903]), .A2(b[903]), .Z(p[903]) );
  XOR2D0 C5244 ( .A1(a[904]), .A2(b[904]), .Z(p[904]) );
  XOR2D0 C5243 ( .A1(a[905]), .A2(b[905]), .Z(p[905]) );
  XOR2D0 C5242 ( .A1(a[906]), .A2(b[906]), .Z(p[906]) );
  XOR2D0 C5241 ( .A1(a[907]), .A2(b[907]), .Z(p[907]) );
  XOR2D0 C5240 ( .A1(a[908]), .A2(b[908]), .Z(p[908]) );
  XOR2D0 C5239 ( .A1(a[909]), .A2(b[909]), .Z(p[909]) );
  XOR2D0 C5238 ( .A1(a[910]), .A2(b[910]), .Z(p[910]) );
  XOR2D0 C5237 ( .A1(a[911]), .A2(b[911]), .Z(p[911]) );
  XOR2D0 C5236 ( .A1(a[912]), .A2(b[912]), .Z(p[912]) );
  XOR2D0 C5235 ( .A1(a[913]), .A2(b[913]), .Z(p[913]) );
  XOR2D0 C5234 ( .A1(a[914]), .A2(b[914]), .Z(p[914]) );
  XOR2D0 C5233 ( .A1(a[915]), .A2(b[915]), .Z(p[915]) );
  XOR2D0 C5232 ( .A1(a[916]), .A2(b[916]), .Z(p[916]) );
  XOR2D0 C5231 ( .A1(a[917]), .A2(b[917]), .Z(p[917]) );
  XOR2D0 C5230 ( .A1(a[918]), .A2(b[918]), .Z(p[918]) );
  XOR2D0 C5229 ( .A1(a[919]), .A2(b[919]), .Z(p[919]) );
  XOR2D0 C5228 ( .A1(a[920]), .A2(b[920]), .Z(p[920]) );
  XOR2D0 C5227 ( .A1(a[921]), .A2(b[921]), .Z(p[921]) );
  XOR2D0 C5226 ( .A1(a[922]), .A2(b[922]), .Z(p[922]) );
  XOR2D0 C5225 ( .A1(a[923]), .A2(b[923]), .Z(p[923]) );
  XOR2D0 C5224 ( .A1(a[924]), .A2(b[924]), .Z(p[924]) );
  XOR2D0 C5223 ( .A1(a[925]), .A2(b[925]), .Z(p[925]) );
  XOR2D0 C5222 ( .A1(a[926]), .A2(b[926]), .Z(p[926]) );
  XOR2D0 C5221 ( .A1(a[927]), .A2(b[927]), .Z(p[927]) );
  XOR2D0 C5220 ( .A1(a[928]), .A2(b[928]), .Z(p[928]) );
  XOR2D0 C5219 ( .A1(a[929]), .A2(b[929]), .Z(p[929]) );
  XOR2D0 C5218 ( .A1(a[930]), .A2(b[930]), .Z(p[930]) );
  XOR2D0 C5217 ( .A1(a[931]), .A2(b[931]), .Z(p[931]) );
  XOR2D0 C5216 ( .A1(a[932]), .A2(b[932]), .Z(p[932]) );
  XOR2D0 C5215 ( .A1(a[933]), .A2(b[933]), .Z(p[933]) );
  XOR2D0 C5214 ( .A1(a[934]), .A2(b[934]), .Z(p[934]) );
  XOR2D0 C5213 ( .A1(a[935]), .A2(b[935]), .Z(p[935]) );
  XOR2D0 C5212 ( .A1(a[936]), .A2(b[936]), .Z(p[936]) );
  XOR2D0 C5211 ( .A1(a[937]), .A2(b[937]), .Z(p[937]) );
  XOR2D0 C5210 ( .A1(a[938]), .A2(b[938]), .Z(p[938]) );
  XOR2D0 C5209 ( .A1(a[939]), .A2(b[939]), .Z(p[939]) );
  XOR2D0 C5208 ( .A1(a[940]), .A2(b[940]), .Z(p[940]) );
  XOR2D0 C5207 ( .A1(a[941]), .A2(b[941]), .Z(p[941]) );
  XOR2D0 C5206 ( .A1(a[942]), .A2(b[942]), .Z(p[942]) );
  XOR2D0 C5205 ( .A1(a[943]), .A2(b[943]), .Z(p[943]) );
  XOR2D0 C5204 ( .A1(a[944]), .A2(b[944]), .Z(p[944]) );
  XOR2D0 C5203 ( .A1(a[945]), .A2(b[945]), .Z(p[945]) );
  XOR2D0 C5202 ( .A1(a[946]), .A2(b[946]), .Z(p[946]) );
  XOR2D0 C5201 ( .A1(a[947]), .A2(b[947]), .Z(p[947]) );
  XOR2D0 C5200 ( .A1(a[948]), .A2(b[948]), .Z(p[948]) );
  XOR2D0 C5199 ( .A1(a[949]), .A2(b[949]), .Z(p[949]) );
  XOR2D0 C5198 ( .A1(a[950]), .A2(b[950]), .Z(p[950]) );
  XOR2D0 C5197 ( .A1(a[951]), .A2(b[951]), .Z(p[951]) );
  XOR2D0 C5196 ( .A1(a[952]), .A2(b[952]), .Z(p[952]) );
  XOR2D0 C5195 ( .A1(a[953]), .A2(b[953]), .Z(p[953]) );
  XOR2D0 C5194 ( .A1(a[954]), .A2(b[954]), .Z(p[954]) );
  XOR2D0 C5193 ( .A1(a[955]), .A2(b[955]), .Z(p[955]) );
  XOR2D0 C5192 ( .A1(a[956]), .A2(b[956]), .Z(p[956]) );
  XOR2D0 C5191 ( .A1(a[957]), .A2(b[957]), .Z(p[957]) );
  XOR2D0 C5190 ( .A1(a[958]), .A2(b[958]), .Z(p[958]) );
  XOR2D0 C5189 ( .A1(a[959]), .A2(b[959]), .Z(p[959]) );
  XOR2D0 C5188 ( .A1(a[960]), .A2(b[960]), .Z(p[960]) );
  XOR2D0 C5187 ( .A1(a[961]), .A2(b[961]), .Z(p[961]) );
  XOR2D0 C5186 ( .A1(a[962]), .A2(b[962]), .Z(p[962]) );
  XOR2D0 C5185 ( .A1(a[963]), .A2(b[963]), .Z(p[963]) );
  XOR2D0 C5184 ( .A1(a[964]), .A2(b[964]), .Z(p[964]) );
  XOR2D0 C5183 ( .A1(a[965]), .A2(b[965]), .Z(p[965]) );
  XOR2D0 C5182 ( .A1(a[966]), .A2(b[966]), .Z(p[966]) );
  XOR2D0 C5181 ( .A1(a[967]), .A2(b[967]), .Z(p[967]) );
  XOR2D0 C5180 ( .A1(a[968]), .A2(b[968]), .Z(p[968]) );
  XOR2D0 C5179 ( .A1(a[969]), .A2(b[969]), .Z(p[969]) );
  XOR2D0 C5178 ( .A1(a[970]), .A2(b[970]), .Z(p[970]) );
  XOR2D0 C5177 ( .A1(a[971]), .A2(b[971]), .Z(p[971]) );
  XOR2D0 C5176 ( .A1(a[972]), .A2(b[972]), .Z(p[972]) );
  XOR2D0 C5175 ( .A1(a[973]), .A2(b[973]), .Z(p[973]) );
  XOR2D0 C5174 ( .A1(a[974]), .A2(b[974]), .Z(p[974]) );
  XOR2D0 C5173 ( .A1(a[975]), .A2(b[975]), .Z(p[975]) );
  XOR2D0 C5172 ( .A1(a[976]), .A2(b[976]), .Z(p[976]) );
  XOR2D0 C5171 ( .A1(a[977]), .A2(b[977]), .Z(p[977]) );
  XOR2D0 C5170 ( .A1(a[978]), .A2(b[978]), .Z(p[978]) );
  XOR2D0 C5169 ( .A1(a[979]), .A2(b[979]), .Z(p[979]) );
  XOR2D0 C5168 ( .A1(a[980]), .A2(b[980]), .Z(p[980]) );
  XOR2D0 C5167 ( .A1(a[981]), .A2(b[981]), .Z(p[981]) );
  XOR2D0 C5166 ( .A1(a[982]), .A2(b[982]), .Z(p[982]) );
  XOR2D0 C5165 ( .A1(a[983]), .A2(b[983]), .Z(p[983]) );
  XOR2D0 C5164 ( .A1(a[984]), .A2(b[984]), .Z(p[984]) );
  XOR2D0 C5163 ( .A1(a[985]), .A2(b[985]), .Z(p[985]) );
  XOR2D0 C5162 ( .A1(a[986]), .A2(b[986]), .Z(p[986]) );
  XOR2D0 C5161 ( .A1(a[987]), .A2(b[987]), .Z(p[987]) );
  XOR2D0 C5160 ( .A1(a[988]), .A2(b[988]), .Z(p[988]) );
  XOR2D0 C5159 ( .A1(a[989]), .A2(b[989]), .Z(p[989]) );
  XOR2D0 C5158 ( .A1(a[990]), .A2(b[990]), .Z(p[990]) );
  XOR2D0 C5157 ( .A1(a[991]), .A2(b[991]), .Z(p[991]) );
  XOR2D0 C5156 ( .A1(a[992]), .A2(b[992]), .Z(p[992]) );
  XOR2D0 C5155 ( .A1(a[993]), .A2(b[993]), .Z(p[993]) );
  XOR2D0 C5154 ( .A1(a[994]), .A2(b[994]), .Z(p[994]) );
  XOR2D0 C5153 ( .A1(a[995]), .A2(b[995]), .Z(p[995]) );
  XOR2D0 C5152 ( .A1(a[996]), .A2(b[996]), .Z(p[996]) );
  XOR2D0 C5151 ( .A1(a[997]), .A2(b[997]), .Z(p[997]) );
  XOR2D0 C5150 ( .A1(a[998]), .A2(b[998]), .Z(p[998]) );
  XOR2D0 C5149 ( .A1(a[999]), .A2(b[999]), .Z(p[999]) );
  XOR2D0 C5148 ( .A1(a[1000]), .A2(b[1000]), .Z(p[1000]) );
  XOR2D0 C5147 ( .A1(a[1001]), .A2(b[1001]), .Z(p[1001]) );
  XOR2D0 C5146 ( .A1(a[1002]), .A2(b[1002]), .Z(p[1002]) );
  XOR2D0 C5145 ( .A1(a[1003]), .A2(b[1003]), .Z(p[1003]) );
  XOR2D0 C5144 ( .A1(a[1004]), .A2(b[1004]), .Z(p[1004]) );
  XOR2D0 C5143 ( .A1(a[1005]), .A2(b[1005]), .Z(p[1005]) );
  XOR2D0 C5142 ( .A1(a[1006]), .A2(b[1006]), .Z(p[1006]) );
  XOR2D0 C5141 ( .A1(a[1007]), .A2(b[1007]), .Z(p[1007]) );
  XOR2D0 C5140 ( .A1(a[1008]), .A2(b[1008]), .Z(p[1008]) );
  XOR2D0 C5139 ( .A1(a[1009]), .A2(b[1009]), .Z(p[1009]) );
  XOR2D0 C5138 ( .A1(a[1010]), .A2(b[1010]), .Z(p[1010]) );
  XOR2D0 C5137 ( .A1(a[1011]), .A2(b[1011]), .Z(p[1011]) );
  XOR2D0 C5136 ( .A1(a[1012]), .A2(b[1012]), .Z(p[1012]) );
  XOR2D0 C5135 ( .A1(a[1013]), .A2(b[1013]), .Z(p[1013]) );
  XOR2D0 C5134 ( .A1(a[1014]), .A2(b[1014]), .Z(p[1014]) );
  XOR2D0 C5133 ( .A1(a[1015]), .A2(b[1015]), .Z(p[1015]) );
  XOR2D0 C5132 ( .A1(a[1016]), .A2(b[1016]), .Z(p[1016]) );
  XOR2D0 C5131 ( .A1(a[1017]), .A2(b[1017]), .Z(p[1017]) );
  XOR2D0 C5130 ( .A1(a[1018]), .A2(b[1018]), .Z(p[1018]) );
  XOR2D0 C5129 ( .A1(a[1019]), .A2(b[1019]), .Z(p[1019]) );
  XOR2D0 C5128 ( .A1(a[1020]), .A2(b[1020]), .Z(p[1020]) );
  XOR2D0 C5127 ( .A1(a[1021]), .A2(b[1021]), .Z(p[1021]) );
  XOR2D0 C5126 ( .A1(a[1022]), .A2(b[1022]), .Z(p[1022]) );
  XOR2D0 C5125 ( .A1(a[1023]), .A2(b[1023]), .Z(p[1023]) );
  AN2D0 C5124 ( .A1(a[0]), .A2(b[0]), .Z(g[0]) );
  AN2D0 C5123 ( .A1(a[1]), .A2(b[1]), .Z(g[1]) );
  AN2D0 C5122 ( .A1(a[2]), .A2(b[2]), .Z(g[2]) );
  AN2D0 C5121 ( .A1(a[3]), .A2(b[3]), .Z(g[3]) );
  AN2D0 C5120 ( .A1(a[4]), .A2(b[4]), .Z(g[4]) );
  AN2D0 C5119 ( .A1(a[5]), .A2(b[5]), .Z(g[5]) );
  AN2D0 C5118 ( .A1(a[6]), .A2(b[6]), .Z(g[6]) );
  AN2D0 C5117 ( .A1(a[7]), .A2(b[7]), .Z(g[7]) );
  AN2D0 C5116 ( .A1(a[8]), .A2(b[8]), .Z(g[8]) );
  AN2D0 C5115 ( .A1(a[9]), .A2(b[9]), .Z(g[9]) );
  AN2D0 C5114 ( .A1(a[10]), .A2(b[10]), .Z(g[10]) );
  AN2D0 C5113 ( .A1(a[11]), .A2(b[11]), .Z(g[11]) );
  AN2D0 C5112 ( .A1(a[12]), .A2(b[12]), .Z(g[12]) );
  AN2D0 C5111 ( .A1(a[13]), .A2(b[13]), .Z(g[13]) );
  AN2D0 C5110 ( .A1(a[14]), .A2(b[14]), .Z(g[14]) );
  AN2D0 C5109 ( .A1(a[15]), .A2(b[15]), .Z(g[15]) );
  AN2D0 C5108 ( .A1(a[16]), .A2(b[16]), .Z(g[16]) );
  AN2D0 C5107 ( .A1(a[17]), .A2(b[17]), .Z(g[17]) );
  AN2D0 C5106 ( .A1(a[18]), .A2(b[18]), .Z(g[18]) );
  AN2D0 C5105 ( .A1(a[19]), .A2(b[19]), .Z(g[19]) );
  AN2D0 C5104 ( .A1(a[20]), .A2(b[20]), .Z(g[20]) );
  AN2D0 C5103 ( .A1(a[21]), .A2(b[21]), .Z(g[21]) );
  AN2D0 C5102 ( .A1(a[22]), .A2(b[22]), .Z(g[22]) );
  AN2D0 C5101 ( .A1(a[23]), .A2(b[23]), .Z(g[23]) );
  AN2D0 C5100 ( .A1(a[24]), .A2(b[24]), .Z(g[24]) );
  AN2D0 C5099 ( .A1(a[25]), .A2(b[25]), .Z(g[25]) );
  AN2D0 C5098 ( .A1(a[26]), .A2(b[26]), .Z(g[26]) );
  AN2D0 C5097 ( .A1(a[27]), .A2(b[27]), .Z(g[27]) );
  AN2D0 C5096 ( .A1(a[28]), .A2(b[28]), .Z(g[28]) );
  AN2D0 C5095 ( .A1(a[29]), .A2(b[29]), .Z(g[29]) );
  AN2D0 C5094 ( .A1(a[30]), .A2(b[30]), .Z(g[30]) );
  AN2D0 C5093 ( .A1(a[31]), .A2(b[31]), .Z(g[31]) );
  AN2D0 C5092 ( .A1(a[32]), .A2(b[32]), .Z(g[32]) );
  AN2D0 C5091 ( .A1(a[33]), .A2(b[33]), .Z(g[33]) );
  AN2D0 C5090 ( .A1(a[34]), .A2(b[34]), .Z(g[34]) );
  AN2D0 C5089 ( .A1(a[35]), .A2(b[35]), .Z(g[35]) );
  AN2D0 C5088 ( .A1(a[36]), .A2(b[36]), .Z(g[36]) );
  AN2D0 C5087 ( .A1(a[37]), .A2(b[37]), .Z(g[37]) );
  AN2D0 C5086 ( .A1(a[38]), .A2(b[38]), .Z(g[38]) );
  AN2D0 C5085 ( .A1(a[39]), .A2(b[39]), .Z(g[39]) );
  AN2D0 C5084 ( .A1(a[40]), .A2(b[40]), .Z(g[40]) );
  AN2D0 C5083 ( .A1(a[41]), .A2(b[41]), .Z(g[41]) );
  AN2D0 C5082 ( .A1(a[42]), .A2(b[42]), .Z(g[42]) );
  AN2D0 C5081 ( .A1(a[43]), .A2(b[43]), .Z(g[43]) );
  AN2D0 C5080 ( .A1(a[44]), .A2(b[44]), .Z(g[44]) );
  AN2D0 C5079 ( .A1(a[45]), .A2(b[45]), .Z(g[45]) );
  AN2D0 C5078 ( .A1(a[46]), .A2(b[46]), .Z(g[46]) );
  AN2D0 C5077 ( .A1(a[47]), .A2(b[47]), .Z(g[47]) );
  AN2D0 C5076 ( .A1(a[48]), .A2(b[48]), .Z(g[48]) );
  AN2D0 C5075 ( .A1(a[49]), .A2(b[49]), .Z(g[49]) );
  AN2D0 C5074 ( .A1(a[50]), .A2(b[50]), .Z(g[50]) );
  AN2D0 C5073 ( .A1(a[51]), .A2(b[51]), .Z(g[51]) );
  AN2D0 C5072 ( .A1(a[52]), .A2(b[52]), .Z(g[52]) );
  AN2D0 C5071 ( .A1(a[53]), .A2(b[53]), .Z(g[53]) );
  AN2D0 C5070 ( .A1(a[54]), .A2(b[54]), .Z(g[54]) );
  AN2D0 C5069 ( .A1(a[55]), .A2(b[55]), .Z(g[55]) );
  AN2D0 C5068 ( .A1(a[56]), .A2(b[56]), .Z(g[56]) );
  AN2D0 C5067 ( .A1(a[57]), .A2(b[57]), .Z(g[57]) );
  AN2D0 C5066 ( .A1(a[58]), .A2(b[58]), .Z(g[58]) );
  AN2D0 C5065 ( .A1(a[59]), .A2(b[59]), .Z(g[59]) );
  AN2D0 C5064 ( .A1(a[60]), .A2(b[60]), .Z(g[60]) );
  AN2D0 C5063 ( .A1(a[61]), .A2(b[61]), .Z(g[61]) );
  AN2D0 C5062 ( .A1(a[62]), .A2(b[62]), .Z(g[62]) );
  AN2D0 C5061 ( .A1(a[63]), .A2(b[63]), .Z(g[63]) );
  AN2D0 C5060 ( .A1(a[64]), .A2(b[64]), .Z(g[64]) );
  AN2D0 C5059 ( .A1(a[65]), .A2(b[65]), .Z(g[65]) );
  AN2D0 C5058 ( .A1(a[66]), .A2(b[66]), .Z(g[66]) );
  AN2D0 C5057 ( .A1(a[67]), .A2(b[67]), .Z(g[67]) );
  AN2D0 C5056 ( .A1(a[68]), .A2(b[68]), .Z(g[68]) );
  AN2D0 C5055 ( .A1(a[69]), .A2(b[69]), .Z(g[69]) );
  AN2D0 C5054 ( .A1(a[70]), .A2(b[70]), .Z(g[70]) );
  AN2D0 C5053 ( .A1(a[71]), .A2(b[71]), .Z(g[71]) );
  AN2D0 C5052 ( .A1(a[72]), .A2(b[72]), .Z(g[72]) );
  AN2D0 C5051 ( .A1(a[73]), .A2(b[73]), .Z(g[73]) );
  AN2D0 C5050 ( .A1(a[74]), .A2(b[74]), .Z(g[74]) );
  AN2D0 C5049 ( .A1(a[75]), .A2(b[75]), .Z(g[75]) );
  AN2D0 C5048 ( .A1(a[76]), .A2(b[76]), .Z(g[76]) );
  AN2D0 C5047 ( .A1(a[77]), .A2(b[77]), .Z(g[77]) );
  AN2D0 C5046 ( .A1(a[78]), .A2(b[78]), .Z(g[78]) );
  AN2D0 C5045 ( .A1(a[79]), .A2(b[79]), .Z(g[79]) );
  AN2D0 C5044 ( .A1(a[80]), .A2(b[80]), .Z(g[80]) );
  AN2D0 C5043 ( .A1(a[81]), .A2(b[81]), .Z(g[81]) );
  AN2D0 C5042 ( .A1(a[82]), .A2(b[82]), .Z(g[82]) );
  AN2D0 C5041 ( .A1(a[83]), .A2(b[83]), .Z(g[83]) );
  AN2D0 C5040 ( .A1(a[84]), .A2(b[84]), .Z(g[84]) );
  AN2D0 C5039 ( .A1(a[85]), .A2(b[85]), .Z(g[85]) );
  AN2D0 C5038 ( .A1(a[86]), .A2(b[86]), .Z(g[86]) );
  AN2D0 C5037 ( .A1(a[87]), .A2(b[87]), .Z(g[87]) );
  AN2D0 C5036 ( .A1(a[88]), .A2(b[88]), .Z(g[88]) );
  AN2D0 C5035 ( .A1(a[89]), .A2(b[89]), .Z(g[89]) );
  AN2D0 C5034 ( .A1(a[90]), .A2(b[90]), .Z(g[90]) );
  AN2D0 C5033 ( .A1(a[91]), .A2(b[91]), .Z(g[91]) );
  AN2D0 C5032 ( .A1(a[92]), .A2(b[92]), .Z(g[92]) );
  AN2D0 C5031 ( .A1(a[93]), .A2(b[93]), .Z(g[93]) );
  AN2D0 C5030 ( .A1(a[94]), .A2(b[94]), .Z(g[94]) );
  AN2D0 C5029 ( .A1(a[95]), .A2(b[95]), .Z(g[95]) );
  AN2D0 C5028 ( .A1(a[96]), .A2(b[96]), .Z(g[96]) );
  AN2D0 C5027 ( .A1(a[97]), .A2(b[97]), .Z(g[97]) );
  AN2D0 C5026 ( .A1(a[98]), .A2(b[98]), .Z(g[98]) );
  AN2D0 C5025 ( .A1(a[99]), .A2(b[99]), .Z(g[99]) );
  AN2D0 C5024 ( .A1(a[100]), .A2(b[100]), .Z(g[100]) );
  AN2D0 C5023 ( .A1(a[101]), .A2(b[101]), .Z(g[101]) );
  AN2D0 C5022 ( .A1(a[102]), .A2(b[102]), .Z(g[102]) );
  AN2D0 C5021 ( .A1(a[103]), .A2(b[103]), .Z(g[103]) );
  AN2D0 C5020 ( .A1(a[104]), .A2(b[104]), .Z(g[104]) );
  AN2D0 C5019 ( .A1(a[105]), .A2(b[105]), .Z(g[105]) );
  AN2D0 C5018 ( .A1(a[106]), .A2(b[106]), .Z(g[106]) );
  AN2D0 C5017 ( .A1(a[107]), .A2(b[107]), .Z(g[107]) );
  AN2D0 C5016 ( .A1(a[108]), .A2(b[108]), .Z(g[108]) );
  AN2D0 C5015 ( .A1(a[109]), .A2(b[109]), .Z(g[109]) );
  AN2D0 C5014 ( .A1(a[110]), .A2(b[110]), .Z(g[110]) );
  AN2D0 C5013 ( .A1(a[111]), .A2(b[111]), .Z(g[111]) );
  AN2D0 C5012 ( .A1(a[112]), .A2(b[112]), .Z(g[112]) );
  AN2D0 C5011 ( .A1(a[113]), .A2(b[113]), .Z(g[113]) );
  AN2D0 C5010 ( .A1(a[114]), .A2(b[114]), .Z(g[114]) );
  AN2D0 C5009 ( .A1(a[115]), .A2(b[115]), .Z(g[115]) );
  AN2D0 C5008 ( .A1(a[116]), .A2(b[116]), .Z(g[116]) );
  AN2D0 C5007 ( .A1(a[117]), .A2(b[117]), .Z(g[117]) );
  AN2D0 C5006 ( .A1(a[118]), .A2(b[118]), .Z(g[118]) );
  AN2D0 C5005 ( .A1(a[119]), .A2(b[119]), .Z(g[119]) );
  AN2D0 C5004 ( .A1(a[120]), .A2(b[120]), .Z(g[120]) );
  AN2D0 C5003 ( .A1(a[121]), .A2(b[121]), .Z(g[121]) );
  AN2D0 C5002 ( .A1(a[122]), .A2(b[122]), .Z(g[122]) );
  AN2D0 C5001 ( .A1(a[123]), .A2(b[123]), .Z(g[123]) );
  AN2D0 C5000 ( .A1(a[124]), .A2(b[124]), .Z(g[124]) );
  AN2D0 C4999 ( .A1(a[125]), .A2(b[125]), .Z(g[125]) );
  AN2D0 C4998 ( .A1(a[126]), .A2(b[126]), .Z(g[126]) );
  AN2D0 C4997 ( .A1(a[127]), .A2(b[127]), .Z(g[127]) );
  AN2D0 C4996 ( .A1(a[128]), .A2(b[128]), .Z(g[128]) );
  AN2D0 C4995 ( .A1(a[129]), .A2(b[129]), .Z(g[129]) );
  AN2D0 C4994 ( .A1(a[130]), .A2(b[130]), .Z(g[130]) );
  AN2D0 C4993 ( .A1(a[131]), .A2(b[131]), .Z(g[131]) );
  AN2D0 C4992 ( .A1(a[132]), .A2(b[132]), .Z(g[132]) );
  AN2D0 C4991 ( .A1(a[133]), .A2(b[133]), .Z(g[133]) );
  AN2D0 C4990 ( .A1(a[134]), .A2(b[134]), .Z(g[134]) );
  AN2D0 C4989 ( .A1(a[135]), .A2(b[135]), .Z(g[135]) );
  AN2D0 C4988 ( .A1(a[136]), .A2(b[136]), .Z(g[136]) );
  AN2D0 C4987 ( .A1(a[137]), .A2(b[137]), .Z(g[137]) );
  AN2D0 C4986 ( .A1(a[138]), .A2(b[138]), .Z(g[138]) );
  AN2D0 C4985 ( .A1(a[139]), .A2(b[139]), .Z(g[139]) );
  AN2D0 C4984 ( .A1(a[140]), .A2(b[140]), .Z(g[140]) );
  AN2D0 C4983 ( .A1(a[141]), .A2(b[141]), .Z(g[141]) );
  AN2D0 C4982 ( .A1(a[142]), .A2(b[142]), .Z(g[142]) );
  AN2D0 C4981 ( .A1(a[143]), .A2(b[143]), .Z(g[143]) );
  AN2D0 C4980 ( .A1(a[144]), .A2(b[144]), .Z(g[144]) );
  AN2D0 C4979 ( .A1(a[145]), .A2(b[145]), .Z(g[145]) );
  AN2D0 C4978 ( .A1(a[146]), .A2(b[146]), .Z(g[146]) );
  AN2D0 C4977 ( .A1(a[147]), .A2(b[147]), .Z(g[147]) );
  AN2D0 C4976 ( .A1(a[148]), .A2(b[148]), .Z(g[148]) );
  AN2D0 C4975 ( .A1(a[149]), .A2(b[149]), .Z(g[149]) );
  AN2D0 C4974 ( .A1(a[150]), .A2(b[150]), .Z(g[150]) );
  AN2D0 C4973 ( .A1(a[151]), .A2(b[151]), .Z(g[151]) );
  AN2D0 C4972 ( .A1(a[152]), .A2(b[152]), .Z(g[152]) );
  AN2D0 C4971 ( .A1(a[153]), .A2(b[153]), .Z(g[153]) );
  AN2D0 C4970 ( .A1(a[154]), .A2(b[154]), .Z(g[154]) );
  AN2D0 C4969 ( .A1(a[155]), .A2(b[155]), .Z(g[155]) );
  AN2D0 C4968 ( .A1(a[156]), .A2(b[156]), .Z(g[156]) );
  AN2D0 C4967 ( .A1(a[157]), .A2(b[157]), .Z(g[157]) );
  AN2D0 C4966 ( .A1(a[158]), .A2(b[158]), .Z(g[158]) );
  AN2D0 C4965 ( .A1(a[159]), .A2(b[159]), .Z(g[159]) );
  AN2D0 C4964 ( .A1(a[160]), .A2(b[160]), .Z(g[160]) );
  AN2D0 C4963 ( .A1(a[161]), .A2(b[161]), .Z(g[161]) );
  AN2D0 C4962 ( .A1(a[162]), .A2(b[162]), .Z(g[162]) );
  AN2D0 C4961 ( .A1(a[163]), .A2(b[163]), .Z(g[163]) );
  AN2D0 C4960 ( .A1(a[164]), .A2(b[164]), .Z(g[164]) );
  AN2D0 C4959 ( .A1(a[165]), .A2(b[165]), .Z(g[165]) );
  AN2D0 C4958 ( .A1(a[166]), .A2(b[166]), .Z(g[166]) );
  AN2D0 C4957 ( .A1(a[167]), .A2(b[167]), .Z(g[167]) );
  AN2D0 C4956 ( .A1(a[168]), .A2(b[168]), .Z(g[168]) );
  AN2D0 C4955 ( .A1(a[169]), .A2(b[169]), .Z(g[169]) );
  AN2D0 C4954 ( .A1(a[170]), .A2(b[170]), .Z(g[170]) );
  AN2D0 C4953 ( .A1(a[171]), .A2(b[171]), .Z(g[171]) );
  AN2D0 C4952 ( .A1(a[172]), .A2(b[172]), .Z(g[172]) );
  AN2D0 C4951 ( .A1(a[173]), .A2(b[173]), .Z(g[173]) );
  AN2D0 C4950 ( .A1(a[174]), .A2(b[174]), .Z(g[174]) );
  AN2D0 C4949 ( .A1(a[175]), .A2(b[175]), .Z(g[175]) );
  AN2D0 C4948 ( .A1(a[176]), .A2(b[176]), .Z(g[176]) );
  AN2D0 C4947 ( .A1(a[177]), .A2(b[177]), .Z(g[177]) );
  AN2D0 C4946 ( .A1(a[178]), .A2(b[178]), .Z(g[178]) );
  AN2D0 C4945 ( .A1(a[179]), .A2(b[179]), .Z(g[179]) );
  AN2D0 C4944 ( .A1(a[180]), .A2(b[180]), .Z(g[180]) );
  AN2D0 C4943 ( .A1(a[181]), .A2(b[181]), .Z(g[181]) );
  AN2D0 C4942 ( .A1(a[182]), .A2(b[182]), .Z(g[182]) );
  AN2D0 C4941 ( .A1(a[183]), .A2(b[183]), .Z(g[183]) );
  AN2D0 C4940 ( .A1(a[184]), .A2(b[184]), .Z(g[184]) );
  AN2D0 C4939 ( .A1(a[185]), .A2(b[185]), .Z(g[185]) );
  AN2D0 C4938 ( .A1(a[186]), .A2(b[186]), .Z(g[186]) );
  AN2D0 C4937 ( .A1(a[187]), .A2(b[187]), .Z(g[187]) );
  AN2D0 C4936 ( .A1(a[188]), .A2(b[188]), .Z(g[188]) );
  AN2D0 C4935 ( .A1(a[189]), .A2(b[189]), .Z(g[189]) );
  AN2D0 C4934 ( .A1(a[190]), .A2(b[190]), .Z(g[190]) );
  AN2D0 C4933 ( .A1(a[191]), .A2(b[191]), .Z(g[191]) );
  AN2D0 C4932 ( .A1(a[192]), .A2(b[192]), .Z(g[192]) );
  AN2D0 C4931 ( .A1(a[193]), .A2(b[193]), .Z(g[193]) );
  AN2D0 C4930 ( .A1(a[194]), .A2(b[194]), .Z(g[194]) );
  AN2D0 C4929 ( .A1(a[195]), .A2(b[195]), .Z(g[195]) );
  AN2D0 C4928 ( .A1(a[196]), .A2(b[196]), .Z(g[196]) );
  AN2D0 C4927 ( .A1(a[197]), .A2(b[197]), .Z(g[197]) );
  AN2D0 C4926 ( .A1(a[198]), .A2(b[198]), .Z(g[198]) );
  AN2D0 C4925 ( .A1(a[199]), .A2(b[199]), .Z(g[199]) );
  AN2D0 C4924 ( .A1(a[200]), .A2(b[200]), .Z(g[200]) );
  AN2D0 C4923 ( .A1(a[201]), .A2(b[201]), .Z(g[201]) );
  AN2D0 C4922 ( .A1(a[202]), .A2(b[202]), .Z(g[202]) );
  AN2D0 C4921 ( .A1(a[203]), .A2(b[203]), .Z(g[203]) );
  AN2D0 C4920 ( .A1(a[204]), .A2(b[204]), .Z(g[204]) );
  AN2D0 C4919 ( .A1(a[205]), .A2(b[205]), .Z(g[205]) );
  AN2D0 C4918 ( .A1(a[206]), .A2(b[206]), .Z(g[206]) );
  AN2D0 C4917 ( .A1(a[207]), .A2(b[207]), .Z(g[207]) );
  AN2D0 C4916 ( .A1(a[208]), .A2(b[208]), .Z(g[208]) );
  AN2D0 C4915 ( .A1(a[209]), .A2(b[209]), .Z(g[209]) );
  AN2D0 C4914 ( .A1(a[210]), .A2(b[210]), .Z(g[210]) );
  AN2D0 C4913 ( .A1(a[211]), .A2(b[211]), .Z(g[211]) );
  AN2D0 C4912 ( .A1(a[212]), .A2(b[212]), .Z(g[212]) );
  AN2D0 C4911 ( .A1(a[213]), .A2(b[213]), .Z(g[213]) );
  AN2D0 C4910 ( .A1(a[214]), .A2(b[214]), .Z(g[214]) );
  AN2D0 C4909 ( .A1(a[215]), .A2(b[215]), .Z(g[215]) );
  AN2D0 C4908 ( .A1(a[216]), .A2(b[216]), .Z(g[216]) );
  AN2D0 C4907 ( .A1(a[217]), .A2(b[217]), .Z(g[217]) );
  AN2D0 C4906 ( .A1(a[218]), .A2(b[218]), .Z(g[218]) );
  AN2D0 C4905 ( .A1(a[219]), .A2(b[219]), .Z(g[219]) );
  AN2D0 C4904 ( .A1(a[220]), .A2(b[220]), .Z(g[220]) );
  AN2D0 C4903 ( .A1(a[221]), .A2(b[221]), .Z(g[221]) );
  AN2D0 C4902 ( .A1(a[222]), .A2(b[222]), .Z(g[222]) );
  AN2D0 C4901 ( .A1(a[223]), .A2(b[223]), .Z(g[223]) );
  AN2D0 C4900 ( .A1(a[224]), .A2(b[224]), .Z(g[224]) );
  AN2D0 C4899 ( .A1(a[225]), .A2(b[225]), .Z(g[225]) );
  AN2D0 C4898 ( .A1(a[226]), .A2(b[226]), .Z(g[226]) );
  AN2D0 C4897 ( .A1(a[227]), .A2(b[227]), .Z(g[227]) );
  AN2D0 C4896 ( .A1(a[228]), .A2(b[228]), .Z(g[228]) );
  AN2D0 C4895 ( .A1(a[229]), .A2(b[229]), .Z(g[229]) );
  AN2D0 C4894 ( .A1(a[230]), .A2(b[230]), .Z(g[230]) );
  AN2D0 C4893 ( .A1(a[231]), .A2(b[231]), .Z(g[231]) );
  AN2D0 C4892 ( .A1(a[232]), .A2(b[232]), .Z(g[232]) );
  AN2D0 C4891 ( .A1(a[233]), .A2(b[233]), .Z(g[233]) );
  AN2D0 C4890 ( .A1(a[234]), .A2(b[234]), .Z(g[234]) );
  AN2D0 C4889 ( .A1(a[235]), .A2(b[235]), .Z(g[235]) );
  AN2D0 C4888 ( .A1(a[236]), .A2(b[236]), .Z(g[236]) );
  AN2D0 C4887 ( .A1(a[237]), .A2(b[237]), .Z(g[237]) );
  AN2D0 C4886 ( .A1(a[238]), .A2(b[238]), .Z(g[238]) );
  AN2D0 C4885 ( .A1(a[239]), .A2(b[239]), .Z(g[239]) );
  AN2D0 C4884 ( .A1(a[240]), .A2(b[240]), .Z(g[240]) );
  AN2D0 C4883 ( .A1(a[241]), .A2(b[241]), .Z(g[241]) );
  AN2D0 C4882 ( .A1(a[242]), .A2(b[242]), .Z(g[242]) );
  AN2D0 C4881 ( .A1(a[243]), .A2(b[243]), .Z(g[243]) );
  AN2D0 C4880 ( .A1(a[244]), .A2(b[244]), .Z(g[244]) );
  AN2D0 C4879 ( .A1(a[245]), .A2(b[245]), .Z(g[245]) );
  AN2D0 C4878 ( .A1(a[246]), .A2(b[246]), .Z(g[246]) );
  AN2D0 C4877 ( .A1(a[247]), .A2(b[247]), .Z(g[247]) );
  AN2D0 C4876 ( .A1(a[248]), .A2(b[248]), .Z(g[248]) );
  AN2D0 C4875 ( .A1(a[249]), .A2(b[249]), .Z(g[249]) );
  AN2D0 C4874 ( .A1(a[250]), .A2(b[250]), .Z(g[250]) );
  AN2D0 C4873 ( .A1(a[251]), .A2(b[251]), .Z(g[251]) );
  AN2D0 C4872 ( .A1(a[252]), .A2(b[252]), .Z(g[252]) );
  AN2D0 C4871 ( .A1(a[253]), .A2(b[253]), .Z(g[253]) );
  AN2D0 C4870 ( .A1(a[254]), .A2(b[254]), .Z(g[254]) );
  AN2D0 C4869 ( .A1(a[255]), .A2(b[255]), .Z(g[255]) );
  AN2D0 C4868 ( .A1(a[256]), .A2(b[256]), .Z(g[256]) );
  AN2D0 C4867 ( .A1(a[257]), .A2(b[257]), .Z(g[257]) );
  AN2D0 C4866 ( .A1(a[258]), .A2(b[258]), .Z(g[258]) );
  AN2D0 C4865 ( .A1(a[259]), .A2(b[259]), .Z(g[259]) );
  AN2D0 C4864 ( .A1(a[260]), .A2(b[260]), .Z(g[260]) );
  AN2D0 C4863 ( .A1(a[261]), .A2(b[261]), .Z(g[261]) );
  AN2D0 C4862 ( .A1(a[262]), .A2(b[262]), .Z(g[262]) );
  AN2D0 C4861 ( .A1(a[263]), .A2(b[263]), .Z(g[263]) );
  AN2D0 C4860 ( .A1(a[264]), .A2(b[264]), .Z(g[264]) );
  AN2D0 C4859 ( .A1(a[265]), .A2(b[265]), .Z(g[265]) );
  AN2D0 C4858 ( .A1(a[266]), .A2(b[266]), .Z(g[266]) );
  AN2D0 C4857 ( .A1(a[267]), .A2(b[267]), .Z(g[267]) );
  AN2D0 C4856 ( .A1(a[268]), .A2(b[268]), .Z(g[268]) );
  AN2D0 C4855 ( .A1(a[269]), .A2(b[269]), .Z(g[269]) );
  AN2D0 C4854 ( .A1(a[270]), .A2(b[270]), .Z(g[270]) );
  AN2D0 C4853 ( .A1(a[271]), .A2(b[271]), .Z(g[271]) );
  AN2D0 C4852 ( .A1(a[272]), .A2(b[272]), .Z(g[272]) );
  AN2D0 C4851 ( .A1(a[273]), .A2(b[273]), .Z(g[273]) );
  AN2D0 C4850 ( .A1(a[274]), .A2(b[274]), .Z(g[274]) );
  AN2D0 C4849 ( .A1(a[275]), .A2(b[275]), .Z(g[275]) );
  AN2D0 C4848 ( .A1(a[276]), .A2(b[276]), .Z(g[276]) );
  AN2D0 C4847 ( .A1(a[277]), .A2(b[277]), .Z(g[277]) );
  AN2D0 C4846 ( .A1(a[278]), .A2(b[278]), .Z(g[278]) );
  AN2D0 C4845 ( .A1(a[279]), .A2(b[279]), .Z(g[279]) );
  AN2D0 C4844 ( .A1(a[280]), .A2(b[280]), .Z(g[280]) );
  AN2D0 C4843 ( .A1(a[281]), .A2(b[281]), .Z(g[281]) );
  AN2D0 C4842 ( .A1(a[282]), .A2(b[282]), .Z(g[282]) );
  AN2D0 C4841 ( .A1(a[283]), .A2(b[283]), .Z(g[283]) );
  AN2D0 C4840 ( .A1(a[284]), .A2(b[284]), .Z(g[284]) );
  AN2D0 C4839 ( .A1(a[285]), .A2(b[285]), .Z(g[285]) );
  AN2D0 C4838 ( .A1(a[286]), .A2(b[286]), .Z(g[286]) );
  AN2D0 C4837 ( .A1(a[287]), .A2(b[287]), .Z(g[287]) );
  AN2D0 C4836 ( .A1(a[288]), .A2(b[288]), .Z(g[288]) );
  AN2D0 C4835 ( .A1(a[289]), .A2(b[289]), .Z(g[289]) );
  AN2D0 C4834 ( .A1(a[290]), .A2(b[290]), .Z(g[290]) );
  AN2D0 C4833 ( .A1(a[291]), .A2(b[291]), .Z(g[291]) );
  AN2D0 C4832 ( .A1(a[292]), .A2(b[292]), .Z(g[292]) );
  AN2D0 C4831 ( .A1(a[293]), .A2(b[293]), .Z(g[293]) );
  AN2D0 C4830 ( .A1(a[294]), .A2(b[294]), .Z(g[294]) );
  AN2D0 C4829 ( .A1(a[295]), .A2(b[295]), .Z(g[295]) );
  AN2D0 C4828 ( .A1(a[296]), .A2(b[296]), .Z(g[296]) );
  AN2D0 C4827 ( .A1(a[297]), .A2(b[297]), .Z(g[297]) );
  AN2D0 C4826 ( .A1(a[298]), .A2(b[298]), .Z(g[298]) );
  AN2D0 C4825 ( .A1(a[299]), .A2(b[299]), .Z(g[299]) );
  AN2D0 C4824 ( .A1(a[300]), .A2(b[300]), .Z(g[300]) );
  AN2D0 C4823 ( .A1(a[301]), .A2(b[301]), .Z(g[301]) );
  AN2D0 C4822 ( .A1(a[302]), .A2(b[302]), .Z(g[302]) );
  AN2D0 C4821 ( .A1(a[303]), .A2(b[303]), .Z(g[303]) );
  AN2D0 C4820 ( .A1(a[304]), .A2(b[304]), .Z(g[304]) );
  AN2D0 C4819 ( .A1(a[305]), .A2(b[305]), .Z(g[305]) );
  AN2D0 C4818 ( .A1(a[306]), .A2(b[306]), .Z(g[306]) );
  AN2D0 C4817 ( .A1(a[307]), .A2(b[307]), .Z(g[307]) );
  AN2D0 C4816 ( .A1(a[308]), .A2(b[308]), .Z(g[308]) );
  AN2D0 C4815 ( .A1(a[309]), .A2(b[309]), .Z(g[309]) );
  AN2D0 C4814 ( .A1(a[310]), .A2(b[310]), .Z(g[310]) );
  AN2D0 C4813 ( .A1(a[311]), .A2(b[311]), .Z(g[311]) );
  AN2D0 C4812 ( .A1(a[312]), .A2(b[312]), .Z(g[312]) );
  AN2D0 C4811 ( .A1(a[313]), .A2(b[313]), .Z(g[313]) );
  AN2D0 C4810 ( .A1(a[314]), .A2(b[314]), .Z(g[314]) );
  AN2D0 C4809 ( .A1(a[315]), .A2(b[315]), .Z(g[315]) );
  AN2D0 C4808 ( .A1(a[316]), .A2(b[316]), .Z(g[316]) );
  AN2D0 C4807 ( .A1(a[317]), .A2(b[317]), .Z(g[317]) );
  AN2D0 C4806 ( .A1(a[318]), .A2(b[318]), .Z(g[318]) );
  AN2D0 C4805 ( .A1(a[319]), .A2(b[319]), .Z(g[319]) );
  AN2D0 C4804 ( .A1(a[320]), .A2(b[320]), .Z(g[320]) );
  AN2D0 C4803 ( .A1(a[321]), .A2(b[321]), .Z(g[321]) );
  AN2D0 C4802 ( .A1(a[322]), .A2(b[322]), .Z(g[322]) );
  AN2D0 C4801 ( .A1(a[323]), .A2(b[323]), .Z(g[323]) );
  AN2D0 C4800 ( .A1(a[324]), .A2(b[324]), .Z(g[324]) );
  AN2D0 C4799 ( .A1(a[325]), .A2(b[325]), .Z(g[325]) );
  AN2D0 C4798 ( .A1(a[326]), .A2(b[326]), .Z(g[326]) );
  AN2D0 C4797 ( .A1(a[327]), .A2(b[327]), .Z(g[327]) );
  AN2D0 C4796 ( .A1(a[328]), .A2(b[328]), .Z(g[328]) );
  AN2D0 C4795 ( .A1(a[329]), .A2(b[329]), .Z(g[329]) );
  AN2D0 C4794 ( .A1(a[330]), .A2(b[330]), .Z(g[330]) );
  AN2D0 C4793 ( .A1(a[331]), .A2(b[331]), .Z(g[331]) );
  AN2D0 C4792 ( .A1(a[332]), .A2(b[332]), .Z(g[332]) );
  AN2D0 C4791 ( .A1(a[333]), .A2(b[333]), .Z(g[333]) );
  AN2D0 C4790 ( .A1(a[334]), .A2(b[334]), .Z(g[334]) );
  AN2D0 C4789 ( .A1(a[335]), .A2(b[335]), .Z(g[335]) );
  AN2D0 C4788 ( .A1(a[336]), .A2(b[336]), .Z(g[336]) );
  AN2D0 C4787 ( .A1(a[337]), .A2(b[337]), .Z(g[337]) );
  AN2D0 C4786 ( .A1(a[338]), .A2(b[338]), .Z(g[338]) );
  AN2D0 C4785 ( .A1(a[339]), .A2(b[339]), .Z(g[339]) );
  AN2D0 C4784 ( .A1(a[340]), .A2(b[340]), .Z(g[340]) );
  AN2D0 C4783 ( .A1(a[341]), .A2(b[341]), .Z(g[341]) );
  AN2D0 C4782 ( .A1(a[342]), .A2(b[342]), .Z(g[342]) );
  AN2D0 C4781 ( .A1(a[343]), .A2(b[343]), .Z(g[343]) );
  AN2D0 C4780 ( .A1(a[344]), .A2(b[344]), .Z(g[344]) );
  AN2D0 C4779 ( .A1(a[345]), .A2(b[345]), .Z(g[345]) );
  AN2D0 C4778 ( .A1(a[346]), .A2(b[346]), .Z(g[346]) );
  AN2D0 C4777 ( .A1(a[347]), .A2(b[347]), .Z(g[347]) );
  AN2D0 C4776 ( .A1(a[348]), .A2(b[348]), .Z(g[348]) );
  AN2D0 C4775 ( .A1(a[349]), .A2(b[349]), .Z(g[349]) );
  AN2D0 C4774 ( .A1(a[350]), .A2(b[350]), .Z(g[350]) );
  AN2D0 C4773 ( .A1(a[351]), .A2(b[351]), .Z(g[351]) );
  AN2D0 C4772 ( .A1(a[352]), .A2(b[352]), .Z(g[352]) );
  AN2D0 C4771 ( .A1(a[353]), .A2(b[353]), .Z(g[353]) );
  AN2D0 C4770 ( .A1(a[354]), .A2(b[354]), .Z(g[354]) );
  AN2D0 C4769 ( .A1(a[355]), .A2(b[355]), .Z(g[355]) );
  AN2D0 C4768 ( .A1(a[356]), .A2(b[356]), .Z(g[356]) );
  AN2D0 C4767 ( .A1(a[357]), .A2(b[357]), .Z(g[357]) );
  AN2D0 C4766 ( .A1(a[358]), .A2(b[358]), .Z(g[358]) );
  AN2D0 C4765 ( .A1(a[359]), .A2(b[359]), .Z(g[359]) );
  AN2D0 C4764 ( .A1(a[360]), .A2(b[360]), .Z(g[360]) );
  AN2D0 C4763 ( .A1(a[361]), .A2(b[361]), .Z(g[361]) );
  AN2D0 C4762 ( .A1(a[362]), .A2(b[362]), .Z(g[362]) );
  AN2D0 C4761 ( .A1(a[363]), .A2(b[363]), .Z(g[363]) );
  AN2D0 C4760 ( .A1(a[364]), .A2(b[364]), .Z(g[364]) );
  AN2D0 C4759 ( .A1(a[365]), .A2(b[365]), .Z(g[365]) );
  AN2D0 C4758 ( .A1(a[366]), .A2(b[366]), .Z(g[366]) );
  AN2D0 C4757 ( .A1(a[367]), .A2(b[367]), .Z(g[367]) );
  AN2D0 C4756 ( .A1(a[368]), .A2(b[368]), .Z(g[368]) );
  AN2D0 C4755 ( .A1(a[369]), .A2(b[369]), .Z(g[369]) );
  AN2D0 C4754 ( .A1(a[370]), .A2(b[370]), .Z(g[370]) );
  AN2D0 C4753 ( .A1(a[371]), .A2(b[371]), .Z(g[371]) );
  AN2D0 C4752 ( .A1(a[372]), .A2(b[372]), .Z(g[372]) );
  AN2D0 C4751 ( .A1(a[373]), .A2(b[373]), .Z(g[373]) );
  AN2D0 C4750 ( .A1(a[374]), .A2(b[374]), .Z(g[374]) );
  AN2D0 C4749 ( .A1(a[375]), .A2(b[375]), .Z(g[375]) );
  AN2D0 C4748 ( .A1(a[376]), .A2(b[376]), .Z(g[376]) );
  AN2D0 C4747 ( .A1(a[377]), .A2(b[377]), .Z(g[377]) );
  AN2D0 C4746 ( .A1(a[378]), .A2(b[378]), .Z(g[378]) );
  AN2D0 C4745 ( .A1(a[379]), .A2(b[379]), .Z(g[379]) );
  AN2D0 C4744 ( .A1(a[380]), .A2(b[380]), .Z(g[380]) );
  AN2D0 C4743 ( .A1(a[381]), .A2(b[381]), .Z(g[381]) );
  AN2D0 C4742 ( .A1(a[382]), .A2(b[382]), .Z(g[382]) );
  AN2D0 C4741 ( .A1(a[383]), .A2(b[383]), .Z(g[383]) );
  AN2D0 C4740 ( .A1(a[384]), .A2(b[384]), .Z(g[384]) );
  AN2D0 C4739 ( .A1(a[385]), .A2(b[385]), .Z(g[385]) );
  AN2D0 C4738 ( .A1(a[386]), .A2(b[386]), .Z(g[386]) );
  AN2D0 C4737 ( .A1(a[387]), .A2(b[387]), .Z(g[387]) );
  AN2D0 C4736 ( .A1(a[388]), .A2(b[388]), .Z(g[388]) );
  AN2D0 C4735 ( .A1(a[389]), .A2(b[389]), .Z(g[389]) );
  AN2D0 C4734 ( .A1(a[390]), .A2(b[390]), .Z(g[390]) );
  AN2D0 C4733 ( .A1(a[391]), .A2(b[391]), .Z(g[391]) );
  AN2D0 C4732 ( .A1(a[392]), .A2(b[392]), .Z(g[392]) );
  AN2D0 C4731 ( .A1(a[393]), .A2(b[393]), .Z(g[393]) );
  AN2D0 C4730 ( .A1(a[394]), .A2(b[394]), .Z(g[394]) );
  AN2D0 C4729 ( .A1(a[395]), .A2(b[395]), .Z(g[395]) );
  AN2D0 C4728 ( .A1(a[396]), .A2(b[396]), .Z(g[396]) );
  AN2D0 C4727 ( .A1(a[397]), .A2(b[397]), .Z(g[397]) );
  AN2D0 C4726 ( .A1(a[398]), .A2(b[398]), .Z(g[398]) );
  AN2D0 C4725 ( .A1(a[399]), .A2(b[399]), .Z(g[399]) );
  AN2D0 C4724 ( .A1(a[400]), .A2(b[400]), .Z(g[400]) );
  AN2D0 C4723 ( .A1(a[401]), .A2(b[401]), .Z(g[401]) );
  AN2D0 C4722 ( .A1(a[402]), .A2(b[402]), .Z(g[402]) );
  AN2D0 C4721 ( .A1(a[403]), .A2(b[403]), .Z(g[403]) );
  AN2D0 C4720 ( .A1(a[404]), .A2(b[404]), .Z(g[404]) );
  AN2D0 C4719 ( .A1(a[405]), .A2(b[405]), .Z(g[405]) );
  AN2D0 C4718 ( .A1(a[406]), .A2(b[406]), .Z(g[406]) );
  AN2D0 C4717 ( .A1(a[407]), .A2(b[407]), .Z(g[407]) );
  AN2D0 C4716 ( .A1(a[408]), .A2(b[408]), .Z(g[408]) );
  AN2D0 C4715 ( .A1(a[409]), .A2(b[409]), .Z(g[409]) );
  AN2D0 C4714 ( .A1(a[410]), .A2(b[410]), .Z(g[410]) );
  AN2D0 C4713 ( .A1(a[411]), .A2(b[411]), .Z(g[411]) );
  AN2D0 C4712 ( .A1(a[412]), .A2(b[412]), .Z(g[412]) );
  AN2D0 C4711 ( .A1(a[413]), .A2(b[413]), .Z(g[413]) );
  AN2D0 C4710 ( .A1(a[414]), .A2(b[414]), .Z(g[414]) );
  AN2D0 C4709 ( .A1(a[415]), .A2(b[415]), .Z(g[415]) );
  AN2D0 C4708 ( .A1(a[416]), .A2(b[416]), .Z(g[416]) );
  AN2D0 C4707 ( .A1(a[417]), .A2(b[417]), .Z(g[417]) );
  AN2D0 C4706 ( .A1(a[418]), .A2(b[418]), .Z(g[418]) );
  AN2D0 C4705 ( .A1(a[419]), .A2(b[419]), .Z(g[419]) );
  AN2D0 C4704 ( .A1(a[420]), .A2(b[420]), .Z(g[420]) );
  AN2D0 C4703 ( .A1(a[421]), .A2(b[421]), .Z(g[421]) );
  AN2D0 C4702 ( .A1(a[422]), .A2(b[422]), .Z(g[422]) );
  AN2D0 C4701 ( .A1(a[423]), .A2(b[423]), .Z(g[423]) );
  AN2D0 C4700 ( .A1(a[424]), .A2(b[424]), .Z(g[424]) );
  AN2D0 C4699 ( .A1(a[425]), .A2(b[425]), .Z(g[425]) );
  AN2D0 C4698 ( .A1(a[426]), .A2(b[426]), .Z(g[426]) );
  AN2D0 C4697 ( .A1(a[427]), .A2(b[427]), .Z(g[427]) );
  AN2D0 C4696 ( .A1(a[428]), .A2(b[428]), .Z(g[428]) );
  AN2D0 C4695 ( .A1(a[429]), .A2(b[429]), .Z(g[429]) );
  AN2D0 C4694 ( .A1(a[430]), .A2(b[430]), .Z(g[430]) );
  AN2D0 C4693 ( .A1(a[431]), .A2(b[431]), .Z(g[431]) );
  AN2D0 C4692 ( .A1(a[432]), .A2(b[432]), .Z(g[432]) );
  AN2D0 C4691 ( .A1(a[433]), .A2(b[433]), .Z(g[433]) );
  AN2D0 C4690 ( .A1(a[434]), .A2(b[434]), .Z(g[434]) );
  AN2D0 C4689 ( .A1(a[435]), .A2(b[435]), .Z(g[435]) );
  AN2D0 C4688 ( .A1(a[436]), .A2(b[436]), .Z(g[436]) );
  AN2D0 C4687 ( .A1(a[437]), .A2(b[437]), .Z(g[437]) );
  AN2D0 C4686 ( .A1(a[438]), .A2(b[438]), .Z(g[438]) );
  AN2D0 C4685 ( .A1(a[439]), .A2(b[439]), .Z(g[439]) );
  AN2D0 C4684 ( .A1(a[440]), .A2(b[440]), .Z(g[440]) );
  AN2D0 C4683 ( .A1(a[441]), .A2(b[441]), .Z(g[441]) );
  AN2D0 C4682 ( .A1(a[442]), .A2(b[442]), .Z(g[442]) );
  AN2D0 C4681 ( .A1(a[443]), .A2(b[443]), .Z(g[443]) );
  AN2D0 C4680 ( .A1(a[444]), .A2(b[444]), .Z(g[444]) );
  AN2D0 C4679 ( .A1(a[445]), .A2(b[445]), .Z(g[445]) );
  AN2D0 C4678 ( .A1(a[446]), .A2(b[446]), .Z(g[446]) );
  AN2D0 C4677 ( .A1(a[447]), .A2(b[447]), .Z(g[447]) );
  AN2D0 C4676 ( .A1(a[448]), .A2(b[448]), .Z(g[448]) );
  AN2D0 C4675 ( .A1(a[449]), .A2(b[449]), .Z(g[449]) );
  AN2D0 C4674 ( .A1(a[450]), .A2(b[450]), .Z(g[450]) );
  AN2D0 C4673 ( .A1(a[451]), .A2(b[451]), .Z(g[451]) );
  AN2D0 C4672 ( .A1(a[452]), .A2(b[452]), .Z(g[452]) );
  AN2D0 C4671 ( .A1(a[453]), .A2(b[453]), .Z(g[453]) );
  AN2D0 C4670 ( .A1(a[454]), .A2(b[454]), .Z(g[454]) );
  AN2D0 C4669 ( .A1(a[455]), .A2(b[455]), .Z(g[455]) );
  AN2D0 C4668 ( .A1(a[456]), .A2(b[456]), .Z(g[456]) );
  AN2D0 C4667 ( .A1(a[457]), .A2(b[457]), .Z(g[457]) );
  AN2D0 C4666 ( .A1(a[458]), .A2(b[458]), .Z(g[458]) );
  AN2D0 C4665 ( .A1(a[459]), .A2(b[459]), .Z(g[459]) );
  AN2D0 C4664 ( .A1(a[460]), .A2(b[460]), .Z(g[460]) );
  AN2D0 C4663 ( .A1(a[461]), .A2(b[461]), .Z(g[461]) );
  AN2D0 C4662 ( .A1(a[462]), .A2(b[462]), .Z(g[462]) );
  AN2D0 C4661 ( .A1(a[463]), .A2(b[463]), .Z(g[463]) );
  AN2D0 C4660 ( .A1(a[464]), .A2(b[464]), .Z(g[464]) );
  AN2D0 C4659 ( .A1(a[465]), .A2(b[465]), .Z(g[465]) );
  AN2D0 C4658 ( .A1(a[466]), .A2(b[466]), .Z(g[466]) );
  AN2D0 C4657 ( .A1(a[467]), .A2(b[467]), .Z(g[467]) );
  AN2D0 C4656 ( .A1(a[468]), .A2(b[468]), .Z(g[468]) );
  AN2D0 C4655 ( .A1(a[469]), .A2(b[469]), .Z(g[469]) );
  AN2D0 C4654 ( .A1(a[470]), .A2(b[470]), .Z(g[470]) );
  AN2D0 C4653 ( .A1(a[471]), .A2(b[471]), .Z(g[471]) );
  AN2D0 C4652 ( .A1(a[472]), .A2(b[472]), .Z(g[472]) );
  AN2D0 C4651 ( .A1(a[473]), .A2(b[473]), .Z(g[473]) );
  AN2D0 C4650 ( .A1(a[474]), .A2(b[474]), .Z(g[474]) );
  AN2D0 C4649 ( .A1(a[475]), .A2(b[475]), .Z(g[475]) );
  AN2D0 C4648 ( .A1(a[476]), .A2(b[476]), .Z(g[476]) );
  AN2D0 C4647 ( .A1(a[477]), .A2(b[477]), .Z(g[477]) );
  AN2D0 C4646 ( .A1(a[478]), .A2(b[478]), .Z(g[478]) );
  AN2D0 C4645 ( .A1(a[479]), .A2(b[479]), .Z(g[479]) );
  AN2D0 C4644 ( .A1(a[480]), .A2(b[480]), .Z(g[480]) );
  AN2D0 C4643 ( .A1(a[481]), .A2(b[481]), .Z(g[481]) );
  AN2D0 C4642 ( .A1(a[482]), .A2(b[482]), .Z(g[482]) );
  AN2D0 C4641 ( .A1(a[483]), .A2(b[483]), .Z(g[483]) );
  AN2D0 C4640 ( .A1(a[484]), .A2(b[484]), .Z(g[484]) );
  AN2D0 C4639 ( .A1(a[485]), .A2(b[485]), .Z(g[485]) );
  AN2D0 C4638 ( .A1(a[486]), .A2(b[486]), .Z(g[486]) );
  AN2D0 C4637 ( .A1(a[487]), .A2(b[487]), .Z(g[487]) );
  AN2D0 C4636 ( .A1(a[488]), .A2(b[488]), .Z(g[488]) );
  AN2D0 C4635 ( .A1(a[489]), .A2(b[489]), .Z(g[489]) );
  AN2D0 C4634 ( .A1(a[490]), .A2(b[490]), .Z(g[490]) );
  AN2D0 C4633 ( .A1(a[491]), .A2(b[491]), .Z(g[491]) );
  AN2D0 C4632 ( .A1(a[492]), .A2(b[492]), .Z(g[492]) );
  AN2D0 C4631 ( .A1(a[493]), .A2(b[493]), .Z(g[493]) );
  AN2D0 C4630 ( .A1(a[494]), .A2(b[494]), .Z(g[494]) );
  AN2D0 C4629 ( .A1(a[495]), .A2(b[495]), .Z(g[495]) );
  AN2D0 C4628 ( .A1(a[496]), .A2(b[496]), .Z(g[496]) );
  AN2D0 C4627 ( .A1(a[497]), .A2(b[497]), .Z(g[497]) );
  AN2D0 C4626 ( .A1(a[498]), .A2(b[498]), .Z(g[498]) );
  AN2D0 C4625 ( .A1(a[499]), .A2(b[499]), .Z(g[499]) );
  AN2D0 C4624 ( .A1(a[500]), .A2(b[500]), .Z(g[500]) );
  AN2D0 C4623 ( .A1(a[501]), .A2(b[501]), .Z(g[501]) );
  AN2D0 C4622 ( .A1(a[502]), .A2(b[502]), .Z(g[502]) );
  AN2D0 C4621 ( .A1(a[503]), .A2(b[503]), .Z(g[503]) );
  AN2D0 C4620 ( .A1(a[504]), .A2(b[504]), .Z(g[504]) );
  AN2D0 C4619 ( .A1(a[505]), .A2(b[505]), .Z(g[505]) );
  AN2D0 C4618 ( .A1(a[506]), .A2(b[506]), .Z(g[506]) );
  AN2D0 C4617 ( .A1(a[507]), .A2(b[507]), .Z(g[507]) );
  AN2D0 C4616 ( .A1(a[508]), .A2(b[508]), .Z(g[508]) );
  AN2D0 C4615 ( .A1(a[509]), .A2(b[509]), .Z(g[509]) );
  AN2D0 C4614 ( .A1(a[510]), .A2(b[510]), .Z(g[510]) );
  AN2D0 C4613 ( .A1(a[511]), .A2(b[511]), .Z(g[511]) );
  AN2D0 C4612 ( .A1(a[512]), .A2(b[512]), .Z(g[512]) );
  AN2D0 C4611 ( .A1(a[513]), .A2(b[513]), .Z(g[513]) );
  AN2D0 C4610 ( .A1(a[514]), .A2(b[514]), .Z(g[514]) );
  AN2D0 C4609 ( .A1(a[515]), .A2(b[515]), .Z(g[515]) );
  AN2D0 C4608 ( .A1(a[516]), .A2(b[516]), .Z(g[516]) );
  AN2D0 C4607 ( .A1(a[517]), .A2(b[517]), .Z(g[517]) );
  AN2D0 C4606 ( .A1(a[518]), .A2(b[518]), .Z(g[518]) );
  AN2D0 C4605 ( .A1(a[519]), .A2(b[519]), .Z(g[519]) );
  AN2D0 C4604 ( .A1(a[520]), .A2(b[520]), .Z(g[520]) );
  AN2D0 C4603 ( .A1(a[521]), .A2(b[521]), .Z(g[521]) );
  AN2D0 C4602 ( .A1(a[522]), .A2(b[522]), .Z(g[522]) );
  AN2D0 C4601 ( .A1(a[523]), .A2(b[523]), .Z(g[523]) );
  AN2D0 C4600 ( .A1(a[524]), .A2(b[524]), .Z(g[524]) );
  AN2D0 C4599 ( .A1(a[525]), .A2(b[525]), .Z(g[525]) );
  AN2D0 C4598 ( .A1(a[526]), .A2(b[526]), .Z(g[526]) );
  AN2D0 C4597 ( .A1(a[527]), .A2(b[527]), .Z(g[527]) );
  AN2D0 C4596 ( .A1(a[528]), .A2(b[528]), .Z(g[528]) );
  AN2D0 C4595 ( .A1(a[529]), .A2(b[529]), .Z(g[529]) );
  AN2D0 C4594 ( .A1(a[530]), .A2(b[530]), .Z(g[530]) );
  AN2D0 C4593 ( .A1(a[531]), .A2(b[531]), .Z(g[531]) );
  AN2D0 C4592 ( .A1(a[532]), .A2(b[532]), .Z(g[532]) );
  AN2D0 C4591 ( .A1(a[533]), .A2(b[533]), .Z(g[533]) );
  AN2D0 C4590 ( .A1(a[534]), .A2(b[534]), .Z(g[534]) );
  AN2D0 C4589 ( .A1(a[535]), .A2(b[535]), .Z(g[535]) );
  AN2D0 C4588 ( .A1(a[536]), .A2(b[536]), .Z(g[536]) );
  AN2D0 C4587 ( .A1(a[537]), .A2(b[537]), .Z(g[537]) );
  AN2D0 C4586 ( .A1(a[538]), .A2(b[538]), .Z(g[538]) );
  AN2D0 C4585 ( .A1(a[539]), .A2(b[539]), .Z(g[539]) );
  AN2D0 C4584 ( .A1(a[540]), .A2(b[540]), .Z(g[540]) );
  AN2D0 C4583 ( .A1(a[541]), .A2(b[541]), .Z(g[541]) );
  AN2D0 C4582 ( .A1(a[542]), .A2(b[542]), .Z(g[542]) );
  AN2D0 C4581 ( .A1(a[543]), .A2(b[543]), .Z(g[543]) );
  AN2D0 C4580 ( .A1(a[544]), .A2(b[544]), .Z(g[544]) );
  AN2D0 C4579 ( .A1(a[545]), .A2(b[545]), .Z(g[545]) );
  AN2D0 C4578 ( .A1(a[546]), .A2(b[546]), .Z(g[546]) );
  AN2D0 C4577 ( .A1(a[547]), .A2(b[547]), .Z(g[547]) );
  AN2D0 C4576 ( .A1(a[548]), .A2(b[548]), .Z(g[548]) );
  AN2D0 C4575 ( .A1(a[549]), .A2(b[549]), .Z(g[549]) );
  AN2D0 C4574 ( .A1(a[550]), .A2(b[550]), .Z(g[550]) );
  AN2D0 C4573 ( .A1(a[551]), .A2(b[551]), .Z(g[551]) );
  AN2D0 C4572 ( .A1(a[552]), .A2(b[552]), .Z(g[552]) );
  AN2D0 C4571 ( .A1(a[553]), .A2(b[553]), .Z(g[553]) );
  AN2D0 C4570 ( .A1(a[554]), .A2(b[554]), .Z(g[554]) );
  AN2D0 C4569 ( .A1(a[555]), .A2(b[555]), .Z(g[555]) );
  AN2D0 C4568 ( .A1(a[556]), .A2(b[556]), .Z(g[556]) );
  AN2D0 C4567 ( .A1(a[557]), .A2(b[557]), .Z(g[557]) );
  AN2D0 C4566 ( .A1(a[558]), .A2(b[558]), .Z(g[558]) );
  AN2D0 C4565 ( .A1(a[559]), .A2(b[559]), .Z(g[559]) );
  AN2D0 C4564 ( .A1(a[560]), .A2(b[560]), .Z(g[560]) );
  AN2D0 C4563 ( .A1(a[561]), .A2(b[561]), .Z(g[561]) );
  AN2D0 C4562 ( .A1(a[562]), .A2(b[562]), .Z(g[562]) );
  AN2D0 C4561 ( .A1(a[563]), .A2(b[563]), .Z(g[563]) );
  AN2D0 C4560 ( .A1(a[564]), .A2(b[564]), .Z(g[564]) );
  AN2D0 C4559 ( .A1(a[565]), .A2(b[565]), .Z(g[565]) );
  AN2D0 C4558 ( .A1(a[566]), .A2(b[566]), .Z(g[566]) );
  AN2D0 C4557 ( .A1(a[567]), .A2(b[567]), .Z(g[567]) );
  AN2D0 C4556 ( .A1(a[568]), .A2(b[568]), .Z(g[568]) );
  AN2D0 C4555 ( .A1(a[569]), .A2(b[569]), .Z(g[569]) );
  AN2D0 C4554 ( .A1(a[570]), .A2(b[570]), .Z(g[570]) );
  AN2D0 C4553 ( .A1(a[571]), .A2(b[571]), .Z(g[571]) );
  AN2D0 C4552 ( .A1(a[572]), .A2(b[572]), .Z(g[572]) );
  AN2D0 C4551 ( .A1(a[573]), .A2(b[573]), .Z(g[573]) );
  AN2D0 C4550 ( .A1(a[574]), .A2(b[574]), .Z(g[574]) );
  AN2D0 C4549 ( .A1(a[575]), .A2(b[575]), .Z(g[575]) );
  AN2D0 C4548 ( .A1(a[576]), .A2(b[576]), .Z(g[576]) );
  AN2D0 C4547 ( .A1(a[577]), .A2(b[577]), .Z(g[577]) );
  AN2D0 C4546 ( .A1(a[578]), .A2(b[578]), .Z(g[578]) );
  AN2D0 C4545 ( .A1(a[579]), .A2(b[579]), .Z(g[579]) );
  AN2D0 C4544 ( .A1(a[580]), .A2(b[580]), .Z(g[580]) );
  AN2D0 C4543 ( .A1(a[581]), .A2(b[581]), .Z(g[581]) );
  AN2D0 C4542 ( .A1(a[582]), .A2(b[582]), .Z(g[582]) );
  AN2D0 C4541 ( .A1(a[583]), .A2(b[583]), .Z(g[583]) );
  AN2D0 C4540 ( .A1(a[584]), .A2(b[584]), .Z(g[584]) );
  AN2D0 C4539 ( .A1(a[585]), .A2(b[585]), .Z(g[585]) );
  AN2D0 C4538 ( .A1(a[586]), .A2(b[586]), .Z(g[586]) );
  AN2D0 C4537 ( .A1(a[587]), .A2(b[587]), .Z(g[587]) );
  AN2D0 C4536 ( .A1(a[588]), .A2(b[588]), .Z(g[588]) );
  AN2D0 C4535 ( .A1(a[589]), .A2(b[589]), .Z(g[589]) );
  AN2D0 C4534 ( .A1(a[590]), .A2(b[590]), .Z(g[590]) );
  AN2D0 C4533 ( .A1(a[591]), .A2(b[591]), .Z(g[591]) );
  AN2D0 C4532 ( .A1(a[592]), .A2(b[592]), .Z(g[592]) );
  AN2D0 C4531 ( .A1(a[593]), .A2(b[593]), .Z(g[593]) );
  AN2D0 C4530 ( .A1(a[594]), .A2(b[594]), .Z(g[594]) );
  AN2D0 C4529 ( .A1(a[595]), .A2(b[595]), .Z(g[595]) );
  AN2D0 C4528 ( .A1(a[596]), .A2(b[596]), .Z(g[596]) );
  AN2D0 C4527 ( .A1(a[597]), .A2(b[597]), .Z(g[597]) );
  AN2D0 C4526 ( .A1(a[598]), .A2(b[598]), .Z(g[598]) );
  AN2D0 C4525 ( .A1(a[599]), .A2(b[599]), .Z(g[599]) );
  AN2D0 C4524 ( .A1(a[600]), .A2(b[600]), .Z(g[600]) );
  AN2D0 C4523 ( .A1(a[601]), .A2(b[601]), .Z(g[601]) );
  AN2D0 C4522 ( .A1(a[602]), .A2(b[602]), .Z(g[602]) );
  AN2D0 C4521 ( .A1(a[603]), .A2(b[603]), .Z(g[603]) );
  AN2D0 C4520 ( .A1(a[604]), .A2(b[604]), .Z(g[604]) );
  AN2D0 C4519 ( .A1(a[605]), .A2(b[605]), .Z(g[605]) );
  AN2D0 C4518 ( .A1(a[606]), .A2(b[606]), .Z(g[606]) );
  AN2D0 C4517 ( .A1(a[607]), .A2(b[607]), .Z(g[607]) );
  AN2D0 C4516 ( .A1(a[608]), .A2(b[608]), .Z(g[608]) );
  AN2D0 C4515 ( .A1(a[609]), .A2(b[609]), .Z(g[609]) );
  AN2D0 C4514 ( .A1(a[610]), .A2(b[610]), .Z(g[610]) );
  AN2D0 C4513 ( .A1(a[611]), .A2(b[611]), .Z(g[611]) );
  AN2D0 C4512 ( .A1(a[612]), .A2(b[612]), .Z(g[612]) );
  AN2D0 C4511 ( .A1(a[613]), .A2(b[613]), .Z(g[613]) );
  AN2D0 C4510 ( .A1(a[614]), .A2(b[614]), .Z(g[614]) );
  AN2D0 C4509 ( .A1(a[615]), .A2(b[615]), .Z(g[615]) );
  AN2D0 C4508 ( .A1(a[616]), .A2(b[616]), .Z(g[616]) );
  AN2D0 C4507 ( .A1(a[617]), .A2(b[617]), .Z(g[617]) );
  AN2D0 C4506 ( .A1(a[618]), .A2(b[618]), .Z(g[618]) );
  AN2D0 C4505 ( .A1(a[619]), .A2(b[619]), .Z(g[619]) );
  AN2D0 C4504 ( .A1(a[620]), .A2(b[620]), .Z(g[620]) );
  AN2D0 C4503 ( .A1(a[621]), .A2(b[621]), .Z(g[621]) );
  AN2D0 C4502 ( .A1(a[622]), .A2(b[622]), .Z(g[622]) );
  AN2D0 C4501 ( .A1(a[623]), .A2(b[623]), .Z(g[623]) );
  AN2D0 C4500 ( .A1(a[624]), .A2(b[624]), .Z(g[624]) );
  AN2D0 C4499 ( .A1(a[625]), .A2(b[625]), .Z(g[625]) );
  AN2D0 C4498 ( .A1(a[626]), .A2(b[626]), .Z(g[626]) );
  AN2D0 C4497 ( .A1(a[627]), .A2(b[627]), .Z(g[627]) );
  AN2D0 C4496 ( .A1(a[628]), .A2(b[628]), .Z(g[628]) );
  AN2D0 C4495 ( .A1(a[629]), .A2(b[629]), .Z(g[629]) );
  AN2D0 C4494 ( .A1(a[630]), .A2(b[630]), .Z(g[630]) );
  AN2D0 C4493 ( .A1(a[631]), .A2(b[631]), .Z(g[631]) );
  AN2D0 C4492 ( .A1(a[632]), .A2(b[632]), .Z(g[632]) );
  AN2D0 C4491 ( .A1(a[633]), .A2(b[633]), .Z(g[633]) );
  AN2D0 C4490 ( .A1(a[634]), .A2(b[634]), .Z(g[634]) );
  AN2D0 C4489 ( .A1(a[635]), .A2(b[635]), .Z(g[635]) );
  AN2D0 C4488 ( .A1(a[636]), .A2(b[636]), .Z(g[636]) );
  AN2D0 C4487 ( .A1(a[637]), .A2(b[637]), .Z(g[637]) );
  AN2D0 C4486 ( .A1(a[638]), .A2(b[638]), .Z(g[638]) );
  AN2D0 C4485 ( .A1(a[639]), .A2(b[639]), .Z(g[639]) );
  AN2D0 C4484 ( .A1(a[640]), .A2(b[640]), .Z(g[640]) );
  AN2D0 C4483 ( .A1(a[641]), .A2(b[641]), .Z(g[641]) );
  AN2D0 C4482 ( .A1(a[642]), .A2(b[642]), .Z(g[642]) );
  AN2D0 C4481 ( .A1(a[643]), .A2(b[643]), .Z(g[643]) );
  AN2D0 C4480 ( .A1(a[644]), .A2(b[644]), .Z(g[644]) );
  AN2D0 C4479 ( .A1(a[645]), .A2(b[645]), .Z(g[645]) );
  AN2D0 C4478 ( .A1(a[646]), .A2(b[646]), .Z(g[646]) );
  AN2D0 C4477 ( .A1(a[647]), .A2(b[647]), .Z(g[647]) );
  AN2D0 C4476 ( .A1(a[648]), .A2(b[648]), .Z(g[648]) );
  AN2D0 C4475 ( .A1(a[649]), .A2(b[649]), .Z(g[649]) );
  AN2D0 C4474 ( .A1(a[650]), .A2(b[650]), .Z(g[650]) );
  AN2D0 C4473 ( .A1(a[651]), .A2(b[651]), .Z(g[651]) );
  AN2D0 C4472 ( .A1(a[652]), .A2(b[652]), .Z(g[652]) );
  AN2D0 C4471 ( .A1(a[653]), .A2(b[653]), .Z(g[653]) );
  AN2D0 C4470 ( .A1(a[654]), .A2(b[654]), .Z(g[654]) );
  AN2D0 C4469 ( .A1(a[655]), .A2(b[655]), .Z(g[655]) );
  AN2D0 C4468 ( .A1(a[656]), .A2(b[656]), .Z(g[656]) );
  AN2D0 C4467 ( .A1(a[657]), .A2(b[657]), .Z(g[657]) );
  AN2D0 C4466 ( .A1(a[658]), .A2(b[658]), .Z(g[658]) );
  AN2D0 C4465 ( .A1(a[659]), .A2(b[659]), .Z(g[659]) );
  AN2D0 C4464 ( .A1(a[660]), .A2(b[660]), .Z(g[660]) );
  AN2D0 C4463 ( .A1(a[661]), .A2(b[661]), .Z(g[661]) );
  AN2D0 C4462 ( .A1(a[662]), .A2(b[662]), .Z(g[662]) );
  AN2D0 C4461 ( .A1(a[663]), .A2(b[663]), .Z(g[663]) );
  AN2D0 C4460 ( .A1(a[664]), .A2(b[664]), .Z(g[664]) );
  AN2D0 C4459 ( .A1(a[665]), .A2(b[665]), .Z(g[665]) );
  AN2D0 C4458 ( .A1(a[666]), .A2(b[666]), .Z(g[666]) );
  AN2D0 C4457 ( .A1(a[667]), .A2(b[667]), .Z(g[667]) );
  AN2D0 C4456 ( .A1(a[668]), .A2(b[668]), .Z(g[668]) );
  AN2D0 C4455 ( .A1(a[669]), .A2(b[669]), .Z(g[669]) );
  AN2D0 C4454 ( .A1(a[670]), .A2(b[670]), .Z(g[670]) );
  AN2D0 C4453 ( .A1(a[671]), .A2(b[671]), .Z(g[671]) );
  AN2D0 C4452 ( .A1(a[672]), .A2(b[672]), .Z(g[672]) );
  AN2D0 C4451 ( .A1(a[673]), .A2(b[673]), .Z(g[673]) );
  AN2D0 C4450 ( .A1(a[674]), .A2(b[674]), .Z(g[674]) );
  AN2D0 C4449 ( .A1(a[675]), .A2(b[675]), .Z(g[675]) );
  AN2D0 C4448 ( .A1(a[676]), .A2(b[676]), .Z(g[676]) );
  AN2D0 C4447 ( .A1(a[677]), .A2(b[677]), .Z(g[677]) );
  AN2D0 C4446 ( .A1(a[678]), .A2(b[678]), .Z(g[678]) );
  AN2D0 C4445 ( .A1(a[679]), .A2(b[679]), .Z(g[679]) );
  AN2D0 C4444 ( .A1(a[680]), .A2(b[680]), .Z(g[680]) );
  AN2D0 C4443 ( .A1(a[681]), .A2(b[681]), .Z(g[681]) );
  AN2D0 C4442 ( .A1(a[682]), .A2(b[682]), .Z(g[682]) );
  AN2D0 C4441 ( .A1(a[683]), .A2(b[683]), .Z(g[683]) );
  AN2D0 C4440 ( .A1(a[684]), .A2(b[684]), .Z(g[684]) );
  AN2D0 C4439 ( .A1(a[685]), .A2(b[685]), .Z(g[685]) );
  AN2D0 C4438 ( .A1(a[686]), .A2(b[686]), .Z(g[686]) );
  AN2D0 C4437 ( .A1(a[687]), .A2(b[687]), .Z(g[687]) );
  AN2D0 C4436 ( .A1(a[688]), .A2(b[688]), .Z(g[688]) );
  AN2D0 C4435 ( .A1(a[689]), .A2(b[689]), .Z(g[689]) );
  AN2D0 C4434 ( .A1(a[690]), .A2(b[690]), .Z(g[690]) );
  AN2D0 C4433 ( .A1(a[691]), .A2(b[691]), .Z(g[691]) );
  AN2D0 C4432 ( .A1(a[692]), .A2(b[692]), .Z(g[692]) );
  AN2D0 C4431 ( .A1(a[693]), .A2(b[693]), .Z(g[693]) );
  AN2D0 C4430 ( .A1(a[694]), .A2(b[694]), .Z(g[694]) );
  AN2D0 C4429 ( .A1(a[695]), .A2(b[695]), .Z(g[695]) );
  AN2D0 C4428 ( .A1(a[696]), .A2(b[696]), .Z(g[696]) );
  AN2D0 C4427 ( .A1(a[697]), .A2(b[697]), .Z(g[697]) );
  AN2D0 C4426 ( .A1(a[698]), .A2(b[698]), .Z(g[698]) );
  AN2D0 C4425 ( .A1(a[699]), .A2(b[699]), .Z(g[699]) );
  AN2D0 C4424 ( .A1(a[700]), .A2(b[700]), .Z(g[700]) );
  AN2D0 C4423 ( .A1(a[701]), .A2(b[701]), .Z(g[701]) );
  AN2D0 C4422 ( .A1(a[702]), .A2(b[702]), .Z(g[702]) );
  AN2D0 C4421 ( .A1(a[703]), .A2(b[703]), .Z(g[703]) );
  AN2D0 C4420 ( .A1(a[704]), .A2(b[704]), .Z(g[704]) );
  AN2D0 C4419 ( .A1(a[705]), .A2(b[705]), .Z(g[705]) );
  AN2D0 C4418 ( .A1(a[706]), .A2(b[706]), .Z(g[706]) );
  AN2D0 C4417 ( .A1(a[707]), .A2(b[707]), .Z(g[707]) );
  AN2D0 C4416 ( .A1(a[708]), .A2(b[708]), .Z(g[708]) );
  AN2D0 C4415 ( .A1(a[709]), .A2(b[709]), .Z(g[709]) );
  AN2D0 C4414 ( .A1(a[710]), .A2(b[710]), .Z(g[710]) );
  AN2D0 C4413 ( .A1(a[711]), .A2(b[711]), .Z(g[711]) );
  AN2D0 C4412 ( .A1(a[712]), .A2(b[712]), .Z(g[712]) );
  AN2D0 C4411 ( .A1(a[713]), .A2(b[713]), .Z(g[713]) );
  AN2D0 C4410 ( .A1(a[714]), .A2(b[714]), .Z(g[714]) );
  AN2D0 C4409 ( .A1(a[715]), .A2(b[715]), .Z(g[715]) );
  AN2D0 C4408 ( .A1(a[716]), .A2(b[716]), .Z(g[716]) );
  AN2D0 C4407 ( .A1(a[717]), .A2(b[717]), .Z(g[717]) );
  AN2D0 C4406 ( .A1(a[718]), .A2(b[718]), .Z(g[718]) );
  AN2D0 C4405 ( .A1(a[719]), .A2(b[719]), .Z(g[719]) );
  AN2D0 C4404 ( .A1(a[720]), .A2(b[720]), .Z(g[720]) );
  AN2D0 C4403 ( .A1(a[721]), .A2(b[721]), .Z(g[721]) );
  AN2D0 C4402 ( .A1(a[722]), .A2(b[722]), .Z(g[722]) );
  AN2D0 C4401 ( .A1(a[723]), .A2(b[723]), .Z(g[723]) );
  AN2D0 C4400 ( .A1(a[724]), .A2(b[724]), .Z(g[724]) );
  AN2D0 C4399 ( .A1(a[725]), .A2(b[725]), .Z(g[725]) );
  AN2D0 C4398 ( .A1(a[726]), .A2(b[726]), .Z(g[726]) );
  AN2D0 C4397 ( .A1(a[727]), .A2(b[727]), .Z(g[727]) );
  AN2D0 C4396 ( .A1(a[728]), .A2(b[728]), .Z(g[728]) );
  AN2D0 C4395 ( .A1(a[729]), .A2(b[729]), .Z(g[729]) );
  AN2D0 C4394 ( .A1(a[730]), .A2(b[730]), .Z(g[730]) );
  AN2D0 C4393 ( .A1(a[731]), .A2(b[731]), .Z(g[731]) );
  AN2D0 C4392 ( .A1(a[732]), .A2(b[732]), .Z(g[732]) );
  AN2D0 C4391 ( .A1(a[733]), .A2(b[733]), .Z(g[733]) );
  AN2D0 C4390 ( .A1(a[734]), .A2(b[734]), .Z(g[734]) );
  AN2D0 C4389 ( .A1(a[735]), .A2(b[735]), .Z(g[735]) );
  AN2D0 C4388 ( .A1(a[736]), .A2(b[736]), .Z(g[736]) );
  AN2D0 C4387 ( .A1(a[737]), .A2(b[737]), .Z(g[737]) );
  AN2D0 C4386 ( .A1(a[738]), .A2(b[738]), .Z(g[738]) );
  AN2D0 C4385 ( .A1(a[739]), .A2(b[739]), .Z(g[739]) );
  AN2D0 C4384 ( .A1(a[740]), .A2(b[740]), .Z(g[740]) );
  AN2D0 C4383 ( .A1(a[741]), .A2(b[741]), .Z(g[741]) );
  AN2D0 C4382 ( .A1(a[742]), .A2(b[742]), .Z(g[742]) );
  AN2D0 C4381 ( .A1(a[743]), .A2(b[743]), .Z(g[743]) );
  AN2D0 C4380 ( .A1(a[744]), .A2(b[744]), .Z(g[744]) );
  AN2D0 C4379 ( .A1(a[745]), .A2(b[745]), .Z(g[745]) );
  AN2D0 C4378 ( .A1(a[746]), .A2(b[746]), .Z(g[746]) );
  AN2D0 C4377 ( .A1(a[747]), .A2(b[747]), .Z(g[747]) );
  AN2D0 C4376 ( .A1(a[748]), .A2(b[748]), .Z(g[748]) );
  AN2D0 C4375 ( .A1(a[749]), .A2(b[749]), .Z(g[749]) );
  AN2D0 C4374 ( .A1(a[750]), .A2(b[750]), .Z(g[750]) );
  AN2D0 C4373 ( .A1(a[751]), .A2(b[751]), .Z(g[751]) );
  AN2D0 C4372 ( .A1(a[752]), .A2(b[752]), .Z(g[752]) );
  AN2D0 C4371 ( .A1(a[753]), .A2(b[753]), .Z(g[753]) );
  AN2D0 C4370 ( .A1(a[754]), .A2(b[754]), .Z(g[754]) );
  AN2D0 C4369 ( .A1(a[755]), .A2(b[755]), .Z(g[755]) );
  AN2D0 C4368 ( .A1(a[756]), .A2(b[756]), .Z(g[756]) );
  AN2D0 C4367 ( .A1(a[757]), .A2(b[757]), .Z(g[757]) );
  AN2D0 C4366 ( .A1(a[758]), .A2(b[758]), .Z(g[758]) );
  AN2D0 C4365 ( .A1(a[759]), .A2(b[759]), .Z(g[759]) );
  AN2D0 C4364 ( .A1(a[760]), .A2(b[760]), .Z(g[760]) );
  AN2D0 C4363 ( .A1(a[761]), .A2(b[761]), .Z(g[761]) );
  AN2D0 C4362 ( .A1(a[762]), .A2(b[762]), .Z(g[762]) );
  AN2D0 C4361 ( .A1(a[763]), .A2(b[763]), .Z(g[763]) );
  AN2D0 C4360 ( .A1(a[764]), .A2(b[764]), .Z(g[764]) );
  AN2D0 C4359 ( .A1(a[765]), .A2(b[765]), .Z(g[765]) );
  AN2D0 C4358 ( .A1(a[766]), .A2(b[766]), .Z(g[766]) );
  AN2D0 C4357 ( .A1(a[767]), .A2(b[767]), .Z(g[767]) );
  AN2D0 C4356 ( .A1(a[768]), .A2(b[768]), .Z(g[768]) );
  AN2D0 C4355 ( .A1(a[769]), .A2(b[769]), .Z(g[769]) );
  AN2D0 C4354 ( .A1(a[770]), .A2(b[770]), .Z(g[770]) );
  AN2D0 C4353 ( .A1(a[771]), .A2(b[771]), .Z(g[771]) );
  AN2D0 C4352 ( .A1(a[772]), .A2(b[772]), .Z(g[772]) );
  AN2D0 C4351 ( .A1(a[773]), .A2(b[773]), .Z(g[773]) );
  AN2D0 C4350 ( .A1(a[774]), .A2(b[774]), .Z(g[774]) );
  AN2D0 C4349 ( .A1(a[775]), .A2(b[775]), .Z(g[775]) );
  AN2D0 C4348 ( .A1(a[776]), .A2(b[776]), .Z(g[776]) );
  AN2D0 C4347 ( .A1(a[777]), .A2(b[777]), .Z(g[777]) );
  AN2D0 C4346 ( .A1(a[778]), .A2(b[778]), .Z(g[778]) );
  AN2D0 C4345 ( .A1(a[779]), .A2(b[779]), .Z(g[779]) );
  AN2D0 C4344 ( .A1(a[780]), .A2(b[780]), .Z(g[780]) );
  AN2D0 C4343 ( .A1(a[781]), .A2(b[781]), .Z(g[781]) );
  AN2D0 C4342 ( .A1(a[782]), .A2(b[782]), .Z(g[782]) );
  AN2D0 C4341 ( .A1(a[783]), .A2(b[783]), .Z(g[783]) );
  AN2D0 C4340 ( .A1(a[784]), .A2(b[784]), .Z(g[784]) );
  AN2D0 C4339 ( .A1(a[785]), .A2(b[785]), .Z(g[785]) );
  AN2D0 C4338 ( .A1(a[786]), .A2(b[786]), .Z(g[786]) );
  AN2D0 C4337 ( .A1(a[787]), .A2(b[787]), .Z(g[787]) );
  AN2D0 C4336 ( .A1(a[788]), .A2(b[788]), .Z(g[788]) );
  AN2D0 C4335 ( .A1(a[789]), .A2(b[789]), .Z(g[789]) );
  AN2D0 C4334 ( .A1(a[790]), .A2(b[790]), .Z(g[790]) );
  AN2D0 C4333 ( .A1(a[791]), .A2(b[791]), .Z(g[791]) );
  AN2D0 C4332 ( .A1(a[792]), .A2(b[792]), .Z(g[792]) );
  AN2D0 C4331 ( .A1(a[793]), .A2(b[793]), .Z(g[793]) );
  AN2D0 C4330 ( .A1(a[794]), .A2(b[794]), .Z(g[794]) );
  AN2D0 C4329 ( .A1(a[795]), .A2(b[795]), .Z(g[795]) );
  AN2D0 C4328 ( .A1(a[796]), .A2(b[796]), .Z(g[796]) );
  AN2D0 C4327 ( .A1(a[797]), .A2(b[797]), .Z(g[797]) );
  AN2D0 C4326 ( .A1(a[798]), .A2(b[798]), .Z(g[798]) );
  AN2D0 C4325 ( .A1(a[799]), .A2(b[799]), .Z(g[799]) );
  AN2D0 C4324 ( .A1(a[800]), .A2(b[800]), .Z(g[800]) );
  AN2D0 C4323 ( .A1(a[801]), .A2(b[801]), .Z(g[801]) );
  AN2D0 C4322 ( .A1(a[802]), .A2(b[802]), .Z(g[802]) );
  AN2D0 C4321 ( .A1(a[803]), .A2(b[803]), .Z(g[803]) );
  AN2D0 C4320 ( .A1(a[804]), .A2(b[804]), .Z(g[804]) );
  AN2D0 C4319 ( .A1(a[805]), .A2(b[805]), .Z(g[805]) );
  AN2D0 C4318 ( .A1(a[806]), .A2(b[806]), .Z(g[806]) );
  AN2D0 C4317 ( .A1(a[807]), .A2(b[807]), .Z(g[807]) );
  AN2D0 C4316 ( .A1(a[808]), .A2(b[808]), .Z(g[808]) );
  AN2D0 C4315 ( .A1(a[809]), .A2(b[809]), .Z(g[809]) );
  AN2D0 C4314 ( .A1(a[810]), .A2(b[810]), .Z(g[810]) );
  AN2D0 C4313 ( .A1(a[811]), .A2(b[811]), .Z(g[811]) );
  AN2D0 C4312 ( .A1(a[812]), .A2(b[812]), .Z(g[812]) );
  AN2D0 C4311 ( .A1(a[813]), .A2(b[813]), .Z(g[813]) );
  AN2D0 C4310 ( .A1(a[814]), .A2(b[814]), .Z(g[814]) );
  AN2D0 C4309 ( .A1(a[815]), .A2(b[815]), .Z(g[815]) );
  AN2D0 C4308 ( .A1(a[816]), .A2(b[816]), .Z(g[816]) );
  AN2D0 C4307 ( .A1(a[817]), .A2(b[817]), .Z(g[817]) );
  AN2D0 C4306 ( .A1(a[818]), .A2(b[818]), .Z(g[818]) );
  AN2D0 C4305 ( .A1(a[819]), .A2(b[819]), .Z(g[819]) );
  AN2D0 C4304 ( .A1(a[820]), .A2(b[820]), .Z(g[820]) );
  AN2D0 C4303 ( .A1(a[821]), .A2(b[821]), .Z(g[821]) );
  AN2D0 C4302 ( .A1(a[822]), .A2(b[822]), .Z(g[822]) );
  AN2D0 C4301 ( .A1(a[823]), .A2(b[823]), .Z(g[823]) );
  AN2D0 C4300 ( .A1(a[824]), .A2(b[824]), .Z(g[824]) );
  AN2D0 C4299 ( .A1(a[825]), .A2(b[825]), .Z(g[825]) );
  AN2D0 C4298 ( .A1(a[826]), .A2(b[826]), .Z(g[826]) );
  AN2D0 C4297 ( .A1(a[827]), .A2(b[827]), .Z(g[827]) );
  AN2D0 C4296 ( .A1(a[828]), .A2(b[828]), .Z(g[828]) );
  AN2D0 C4295 ( .A1(a[829]), .A2(b[829]), .Z(g[829]) );
  AN2D0 C4294 ( .A1(a[830]), .A2(b[830]), .Z(g[830]) );
  AN2D0 C4293 ( .A1(a[831]), .A2(b[831]), .Z(g[831]) );
  AN2D0 C4292 ( .A1(a[832]), .A2(b[832]), .Z(g[832]) );
  AN2D0 C4291 ( .A1(a[833]), .A2(b[833]), .Z(g[833]) );
  AN2D0 C4290 ( .A1(a[834]), .A2(b[834]), .Z(g[834]) );
  AN2D0 C4289 ( .A1(a[835]), .A2(b[835]), .Z(g[835]) );
  AN2D0 C4288 ( .A1(a[836]), .A2(b[836]), .Z(g[836]) );
  AN2D0 C4287 ( .A1(a[837]), .A2(b[837]), .Z(g[837]) );
  AN2D0 C4286 ( .A1(a[838]), .A2(b[838]), .Z(g[838]) );
  AN2D0 C4285 ( .A1(a[839]), .A2(b[839]), .Z(g[839]) );
  AN2D0 C4284 ( .A1(a[840]), .A2(b[840]), .Z(g[840]) );
  AN2D0 C4283 ( .A1(a[841]), .A2(b[841]), .Z(g[841]) );
  AN2D0 C4282 ( .A1(a[842]), .A2(b[842]), .Z(g[842]) );
  AN2D0 C4281 ( .A1(a[843]), .A2(b[843]), .Z(g[843]) );
  AN2D0 C4280 ( .A1(a[844]), .A2(b[844]), .Z(g[844]) );
  AN2D0 C4279 ( .A1(a[845]), .A2(b[845]), .Z(g[845]) );
  AN2D0 C4278 ( .A1(a[846]), .A2(b[846]), .Z(g[846]) );
  AN2D0 C4277 ( .A1(a[847]), .A2(b[847]), .Z(g[847]) );
  AN2D0 C4276 ( .A1(a[848]), .A2(b[848]), .Z(g[848]) );
  AN2D0 C4275 ( .A1(a[849]), .A2(b[849]), .Z(g[849]) );
  AN2D0 C4274 ( .A1(a[850]), .A2(b[850]), .Z(g[850]) );
  AN2D0 C4273 ( .A1(a[851]), .A2(b[851]), .Z(g[851]) );
  AN2D0 C4272 ( .A1(a[852]), .A2(b[852]), .Z(g[852]) );
  AN2D0 C4271 ( .A1(a[853]), .A2(b[853]), .Z(g[853]) );
  AN2D0 C4270 ( .A1(a[854]), .A2(b[854]), .Z(g[854]) );
  AN2D0 C4269 ( .A1(a[855]), .A2(b[855]), .Z(g[855]) );
  AN2D0 C4268 ( .A1(a[856]), .A2(b[856]), .Z(g[856]) );
  AN2D0 C4267 ( .A1(a[857]), .A2(b[857]), .Z(g[857]) );
  AN2D0 C4266 ( .A1(a[858]), .A2(b[858]), .Z(g[858]) );
  AN2D0 C4265 ( .A1(a[859]), .A2(b[859]), .Z(g[859]) );
  AN2D0 C4264 ( .A1(a[860]), .A2(b[860]), .Z(g[860]) );
  AN2D0 C4263 ( .A1(a[861]), .A2(b[861]), .Z(g[861]) );
  AN2D0 C4262 ( .A1(a[862]), .A2(b[862]), .Z(g[862]) );
  AN2D0 C4261 ( .A1(a[863]), .A2(b[863]), .Z(g[863]) );
  AN2D0 C4260 ( .A1(a[864]), .A2(b[864]), .Z(g[864]) );
  AN2D0 C4259 ( .A1(a[865]), .A2(b[865]), .Z(g[865]) );
  AN2D0 C4258 ( .A1(a[866]), .A2(b[866]), .Z(g[866]) );
  AN2D0 C4257 ( .A1(a[867]), .A2(b[867]), .Z(g[867]) );
  AN2D0 C4256 ( .A1(a[868]), .A2(b[868]), .Z(g[868]) );
  AN2D0 C4255 ( .A1(a[869]), .A2(b[869]), .Z(g[869]) );
  AN2D0 C4254 ( .A1(a[870]), .A2(b[870]), .Z(g[870]) );
  AN2D0 C4253 ( .A1(a[871]), .A2(b[871]), .Z(g[871]) );
  AN2D0 C4252 ( .A1(a[872]), .A2(b[872]), .Z(g[872]) );
  AN2D0 C4251 ( .A1(a[873]), .A2(b[873]), .Z(g[873]) );
  AN2D0 C4250 ( .A1(a[874]), .A2(b[874]), .Z(g[874]) );
  AN2D0 C4249 ( .A1(a[875]), .A2(b[875]), .Z(g[875]) );
  AN2D0 C4248 ( .A1(a[876]), .A2(b[876]), .Z(g[876]) );
  AN2D0 C4247 ( .A1(a[877]), .A2(b[877]), .Z(g[877]) );
  AN2D0 C4246 ( .A1(a[878]), .A2(b[878]), .Z(g[878]) );
  AN2D0 C4245 ( .A1(a[879]), .A2(b[879]), .Z(g[879]) );
  AN2D0 C4244 ( .A1(a[880]), .A2(b[880]), .Z(g[880]) );
  AN2D0 C4243 ( .A1(a[881]), .A2(b[881]), .Z(g[881]) );
  AN2D0 C4242 ( .A1(a[882]), .A2(b[882]), .Z(g[882]) );
  AN2D0 C4241 ( .A1(a[883]), .A2(b[883]), .Z(g[883]) );
  AN2D0 C4240 ( .A1(a[884]), .A2(b[884]), .Z(g[884]) );
  AN2D0 C4239 ( .A1(a[885]), .A2(b[885]), .Z(g[885]) );
  AN2D0 C4238 ( .A1(a[886]), .A2(b[886]), .Z(g[886]) );
  AN2D0 C4237 ( .A1(a[887]), .A2(b[887]), .Z(g[887]) );
  AN2D0 C4236 ( .A1(a[888]), .A2(b[888]), .Z(g[888]) );
  AN2D0 C4235 ( .A1(a[889]), .A2(b[889]), .Z(g[889]) );
  AN2D0 C4234 ( .A1(a[890]), .A2(b[890]), .Z(g[890]) );
  AN2D0 C4233 ( .A1(a[891]), .A2(b[891]), .Z(g[891]) );
  AN2D0 C4232 ( .A1(a[892]), .A2(b[892]), .Z(g[892]) );
  AN2D0 C4231 ( .A1(a[893]), .A2(b[893]), .Z(g[893]) );
  AN2D0 C4230 ( .A1(a[894]), .A2(b[894]), .Z(g[894]) );
  AN2D0 C4229 ( .A1(a[895]), .A2(b[895]), .Z(g[895]) );
  AN2D0 C4228 ( .A1(a[896]), .A2(b[896]), .Z(g[896]) );
  AN2D0 C4227 ( .A1(a[897]), .A2(b[897]), .Z(g[897]) );
  AN2D0 C4226 ( .A1(a[898]), .A2(b[898]), .Z(g[898]) );
  AN2D0 C4225 ( .A1(a[899]), .A2(b[899]), .Z(g[899]) );
  AN2D0 C4224 ( .A1(a[900]), .A2(b[900]), .Z(g[900]) );
  AN2D0 C4223 ( .A1(a[901]), .A2(b[901]), .Z(g[901]) );
  AN2D0 C4222 ( .A1(a[902]), .A2(b[902]), .Z(g[902]) );
  AN2D0 C4221 ( .A1(a[903]), .A2(b[903]), .Z(g[903]) );
  AN2D0 C4220 ( .A1(a[904]), .A2(b[904]), .Z(g[904]) );
  AN2D0 C4219 ( .A1(a[905]), .A2(b[905]), .Z(g[905]) );
  AN2D0 C4218 ( .A1(a[906]), .A2(b[906]), .Z(g[906]) );
  AN2D0 C4217 ( .A1(a[907]), .A2(b[907]), .Z(g[907]) );
  AN2D0 C4216 ( .A1(a[908]), .A2(b[908]), .Z(g[908]) );
  AN2D0 C4215 ( .A1(a[909]), .A2(b[909]), .Z(g[909]) );
  AN2D0 C4214 ( .A1(a[910]), .A2(b[910]), .Z(g[910]) );
  AN2D0 C4213 ( .A1(a[911]), .A2(b[911]), .Z(g[911]) );
  AN2D0 C4212 ( .A1(a[912]), .A2(b[912]), .Z(g[912]) );
  AN2D0 C4211 ( .A1(a[913]), .A2(b[913]), .Z(g[913]) );
  AN2D0 C4210 ( .A1(a[914]), .A2(b[914]), .Z(g[914]) );
  AN2D0 C4209 ( .A1(a[915]), .A2(b[915]), .Z(g[915]) );
  AN2D0 C4208 ( .A1(a[916]), .A2(b[916]), .Z(g[916]) );
  AN2D0 C4207 ( .A1(a[917]), .A2(b[917]), .Z(g[917]) );
  AN2D0 C4206 ( .A1(a[918]), .A2(b[918]), .Z(g[918]) );
  AN2D0 C4205 ( .A1(a[919]), .A2(b[919]), .Z(g[919]) );
  AN2D0 C4204 ( .A1(a[920]), .A2(b[920]), .Z(g[920]) );
  AN2D0 C4203 ( .A1(a[921]), .A2(b[921]), .Z(g[921]) );
  AN2D0 C4202 ( .A1(a[922]), .A2(b[922]), .Z(g[922]) );
  AN2D0 C4201 ( .A1(a[923]), .A2(b[923]), .Z(g[923]) );
  AN2D0 C4200 ( .A1(a[924]), .A2(b[924]), .Z(g[924]) );
  AN2D0 C4199 ( .A1(a[925]), .A2(b[925]), .Z(g[925]) );
  AN2D0 C4198 ( .A1(a[926]), .A2(b[926]), .Z(g[926]) );
  AN2D0 C4197 ( .A1(a[927]), .A2(b[927]), .Z(g[927]) );
  AN2D0 C4196 ( .A1(a[928]), .A2(b[928]), .Z(g[928]) );
  AN2D0 C4195 ( .A1(a[929]), .A2(b[929]), .Z(g[929]) );
  AN2D0 C4194 ( .A1(a[930]), .A2(b[930]), .Z(g[930]) );
  AN2D0 C4193 ( .A1(a[931]), .A2(b[931]), .Z(g[931]) );
  AN2D0 C4192 ( .A1(a[932]), .A2(b[932]), .Z(g[932]) );
  AN2D0 C4191 ( .A1(a[933]), .A2(b[933]), .Z(g[933]) );
  AN2D0 C4190 ( .A1(a[934]), .A2(b[934]), .Z(g[934]) );
  AN2D0 C4189 ( .A1(a[935]), .A2(b[935]), .Z(g[935]) );
  AN2D0 C4188 ( .A1(a[936]), .A2(b[936]), .Z(g[936]) );
  AN2D0 C4187 ( .A1(a[937]), .A2(b[937]), .Z(g[937]) );
  AN2D0 C4186 ( .A1(a[938]), .A2(b[938]), .Z(g[938]) );
  AN2D0 C4185 ( .A1(a[939]), .A2(b[939]), .Z(g[939]) );
  AN2D0 C4184 ( .A1(a[940]), .A2(b[940]), .Z(g[940]) );
  AN2D0 C4183 ( .A1(a[941]), .A2(b[941]), .Z(g[941]) );
  AN2D0 C4182 ( .A1(a[942]), .A2(b[942]), .Z(g[942]) );
  AN2D0 C4181 ( .A1(a[943]), .A2(b[943]), .Z(g[943]) );
  AN2D0 C4180 ( .A1(a[944]), .A2(b[944]), .Z(g[944]) );
  AN2D0 C4179 ( .A1(a[945]), .A2(b[945]), .Z(g[945]) );
  AN2D0 C4178 ( .A1(a[946]), .A2(b[946]), .Z(g[946]) );
  AN2D0 C4177 ( .A1(a[947]), .A2(b[947]), .Z(g[947]) );
  AN2D0 C4176 ( .A1(a[948]), .A2(b[948]), .Z(g[948]) );
  AN2D0 C4175 ( .A1(a[949]), .A2(b[949]), .Z(g[949]) );
  AN2D0 C4174 ( .A1(a[950]), .A2(b[950]), .Z(g[950]) );
  AN2D0 C4173 ( .A1(a[951]), .A2(b[951]), .Z(g[951]) );
  AN2D0 C4172 ( .A1(a[952]), .A2(b[952]), .Z(g[952]) );
  AN2D0 C4171 ( .A1(a[953]), .A2(b[953]), .Z(g[953]) );
  AN2D0 C4170 ( .A1(a[954]), .A2(b[954]), .Z(g[954]) );
  AN2D0 C4169 ( .A1(a[955]), .A2(b[955]), .Z(g[955]) );
  AN2D0 C4168 ( .A1(a[956]), .A2(b[956]), .Z(g[956]) );
  AN2D0 C4167 ( .A1(a[957]), .A2(b[957]), .Z(g[957]) );
  AN2D0 C4166 ( .A1(a[958]), .A2(b[958]), .Z(g[958]) );
  AN2D0 C4165 ( .A1(a[959]), .A2(b[959]), .Z(g[959]) );
  AN2D0 C4164 ( .A1(a[960]), .A2(b[960]), .Z(g[960]) );
  AN2D0 C4163 ( .A1(a[961]), .A2(b[961]), .Z(g[961]) );
  AN2D0 C4162 ( .A1(a[962]), .A2(b[962]), .Z(g[962]) );
  AN2D0 C4161 ( .A1(a[963]), .A2(b[963]), .Z(g[963]) );
  AN2D0 C4160 ( .A1(a[964]), .A2(b[964]), .Z(g[964]) );
  AN2D0 C4159 ( .A1(a[965]), .A2(b[965]), .Z(g[965]) );
  AN2D0 C4158 ( .A1(a[966]), .A2(b[966]), .Z(g[966]) );
  AN2D0 C4157 ( .A1(a[967]), .A2(b[967]), .Z(g[967]) );
  AN2D0 C4156 ( .A1(a[968]), .A2(b[968]), .Z(g[968]) );
  AN2D0 C4155 ( .A1(a[969]), .A2(b[969]), .Z(g[969]) );
  AN2D0 C4154 ( .A1(a[970]), .A2(b[970]), .Z(g[970]) );
  AN2D0 C4153 ( .A1(a[971]), .A2(b[971]), .Z(g[971]) );
  AN2D0 C4152 ( .A1(a[972]), .A2(b[972]), .Z(g[972]) );
  AN2D0 C4151 ( .A1(a[973]), .A2(b[973]), .Z(g[973]) );
  AN2D0 C4150 ( .A1(a[974]), .A2(b[974]), .Z(g[974]) );
  AN2D0 C4149 ( .A1(a[975]), .A2(b[975]), .Z(g[975]) );
  AN2D0 C4148 ( .A1(a[976]), .A2(b[976]), .Z(g[976]) );
  AN2D0 C4147 ( .A1(a[977]), .A2(b[977]), .Z(g[977]) );
  AN2D0 C4146 ( .A1(a[978]), .A2(b[978]), .Z(g[978]) );
  AN2D0 C4145 ( .A1(a[979]), .A2(b[979]), .Z(g[979]) );
  AN2D0 C4144 ( .A1(a[980]), .A2(b[980]), .Z(g[980]) );
  AN2D0 C4143 ( .A1(a[981]), .A2(b[981]), .Z(g[981]) );
  AN2D0 C4142 ( .A1(a[982]), .A2(b[982]), .Z(g[982]) );
  AN2D0 C4141 ( .A1(a[983]), .A2(b[983]), .Z(g[983]) );
  AN2D0 C4140 ( .A1(a[984]), .A2(b[984]), .Z(g[984]) );
  AN2D0 C4139 ( .A1(a[985]), .A2(b[985]), .Z(g[985]) );
  AN2D0 C4138 ( .A1(a[986]), .A2(b[986]), .Z(g[986]) );
  AN2D0 C4137 ( .A1(a[987]), .A2(b[987]), .Z(g[987]) );
  AN2D0 C4136 ( .A1(a[988]), .A2(b[988]), .Z(g[988]) );
  AN2D0 C4135 ( .A1(a[989]), .A2(b[989]), .Z(g[989]) );
  AN2D0 C4134 ( .A1(a[990]), .A2(b[990]), .Z(g[990]) );
  AN2D0 C4133 ( .A1(a[991]), .A2(b[991]), .Z(g[991]) );
  AN2D0 C4132 ( .A1(a[992]), .A2(b[992]), .Z(g[992]) );
  AN2D0 C4131 ( .A1(a[993]), .A2(b[993]), .Z(g[993]) );
  AN2D0 C4130 ( .A1(a[994]), .A2(b[994]), .Z(g[994]) );
  AN2D0 C4129 ( .A1(a[995]), .A2(b[995]), .Z(g[995]) );
  AN2D0 C4128 ( .A1(a[996]), .A2(b[996]), .Z(g[996]) );
  AN2D0 C4127 ( .A1(a[997]), .A2(b[997]), .Z(g[997]) );
  AN2D0 C4126 ( .A1(a[998]), .A2(b[998]), .Z(g[998]) );
  AN2D0 C4125 ( .A1(a[999]), .A2(b[999]), .Z(g[999]) );
  AN2D0 C4124 ( .A1(a[1000]), .A2(b[1000]), .Z(g[1000]) );
  AN2D0 C4123 ( .A1(a[1001]), .A2(b[1001]), .Z(g[1001]) );
  AN2D0 C4122 ( .A1(a[1002]), .A2(b[1002]), .Z(g[1002]) );
  AN2D0 C4121 ( .A1(a[1003]), .A2(b[1003]), .Z(g[1003]) );
  AN2D0 C4120 ( .A1(a[1004]), .A2(b[1004]), .Z(g[1004]) );
  AN2D0 C4119 ( .A1(a[1005]), .A2(b[1005]), .Z(g[1005]) );
  AN2D0 C4118 ( .A1(a[1006]), .A2(b[1006]), .Z(g[1006]) );
  AN2D0 C4117 ( .A1(a[1007]), .A2(b[1007]), .Z(g[1007]) );
  AN2D0 C4116 ( .A1(a[1008]), .A2(b[1008]), .Z(g[1008]) );
  AN2D0 C4115 ( .A1(a[1009]), .A2(b[1009]), .Z(g[1009]) );
  AN2D0 C4114 ( .A1(a[1010]), .A2(b[1010]), .Z(g[1010]) );
  AN2D0 C4113 ( .A1(a[1011]), .A2(b[1011]), .Z(g[1011]) );
  AN2D0 C4112 ( .A1(a[1012]), .A2(b[1012]), .Z(g[1012]) );
  AN2D0 C4111 ( .A1(a[1013]), .A2(b[1013]), .Z(g[1013]) );
  AN2D0 C4110 ( .A1(a[1014]), .A2(b[1014]), .Z(g[1014]) );
  AN2D0 C4109 ( .A1(a[1015]), .A2(b[1015]), .Z(g[1015]) );
  AN2D0 C4108 ( .A1(a[1016]), .A2(b[1016]), .Z(g[1016]) );
  AN2D0 C4107 ( .A1(a[1017]), .A2(b[1017]), .Z(g[1017]) );
  AN2D0 C4106 ( .A1(a[1018]), .A2(b[1018]), .Z(g[1018]) );
  AN2D0 C4105 ( .A1(a[1019]), .A2(b[1019]), .Z(g[1019]) );
  AN2D0 C4104 ( .A1(a[1020]), .A2(b[1020]), .Z(g[1020]) );
  AN2D0 C4103 ( .A1(a[1021]), .A2(b[1021]), .Z(g[1021]) );
  AN2D0 C4102 ( .A1(a[1022]), .A2(b[1022]), .Z(g[1022]) );
endmodule

