
module gen_linear_part ( a, b, n, s );
  input [7:0] a;
  input [7:0] b;
  input [501:0] n;
  output [7:0] s;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501;

  XOR2D0 U1 ( .A1(n1), .A2(n2), .Z(s[7]) );
  XOR2D0 U2 ( .A1(a[7]), .A2(n3), .Z(n2) );
  XOR2D0 U3 ( .A1(n4), .A2(n5), .Z(n3) );
  XOR2D0 U4 ( .A1(n6), .A2(n7), .Z(n5) );
  XOR2D0 U5 ( .A1(n[492]), .A2(n8), .Z(n7) );
  XOR2D0 U6 ( .A1(n9), .A2(n10), .Z(n8) );
  XOR2D0 U7 ( .A1(n11), .A2(n12), .Z(n10) );
  XOR2D0 U8 ( .A1(n[485]), .A2(n13), .Z(n12) );
  XOR2D0 U9 ( .A1(n14), .A2(n15), .Z(n13) );
  XOR2D0 U10 ( .A1(n16), .A2(n17), .Z(n15) );
  XOR2D0 U11 ( .A1(n[478]), .A2(n18), .Z(n17) );
  XOR2D0 U12 ( .A1(n19), .A2(n20), .Z(n18) );
  XOR2D0 U13 ( .A1(n21), .A2(n22), .Z(n20) );
  XOR2D0 U14 ( .A1(n[471]), .A2(n23), .Z(n22) );
  XOR2D0 U15 ( .A1(n24), .A2(n25), .Z(n23) );
  XOR2D0 U16 ( .A1(n26), .A2(n27), .Z(n25) );
  XOR2D0 U17 ( .A1(n[464]), .A2(n28), .Z(n27) );
  XOR2D0 U18 ( .A1(n29), .A2(n30), .Z(n28) );
  XOR2D0 U19 ( .A1(n31), .A2(n32), .Z(n30) );
  XOR2D0 U20 ( .A1(n[457]), .A2(n33), .Z(n32) );
  XOR2D0 U21 ( .A1(n34), .A2(n35), .Z(n33) );
  XOR2D0 U22 ( .A1(n36), .A2(n37), .Z(n35) );
  XOR2D0 U23 ( .A1(n[450]), .A2(n38), .Z(n37) );
  XOR2D0 U24 ( .A1(n39), .A2(n40), .Z(n38) );
  XOR2D0 U25 ( .A1(n41), .A2(n42), .Z(n40) );
  XOR2D0 U26 ( .A1(n[443]), .A2(n43), .Z(n42) );
  XOR2D0 U27 ( .A1(n44), .A2(n45), .Z(n43) );
  XOR2D0 U28 ( .A1(n46), .A2(n47), .Z(n45) );
  XOR2D0 U29 ( .A1(n[436]), .A2(n48), .Z(n47) );
  XOR2D0 U30 ( .A1(n49), .A2(n50), .Z(n48) );
  XOR2D0 U31 ( .A1(n51), .A2(n52), .Z(n50) );
  XOR2D0 U32 ( .A1(n[429]), .A2(n53), .Z(n52) );
  XOR2D0 U33 ( .A1(n54), .A2(n55), .Z(n53) );
  XOR2D0 U34 ( .A1(n56), .A2(n57), .Z(n55) );
  XOR2D0 U35 ( .A1(n[422]), .A2(n58), .Z(n57) );
  XOR2D0 U36 ( .A1(n59), .A2(n60), .Z(n58) );
  XOR2D0 U37 ( .A1(n61), .A2(n62), .Z(n60) );
  XOR2D0 U38 ( .A1(n[415]), .A2(n63), .Z(n62) );
  XOR2D0 U39 ( .A1(n64), .A2(n65), .Z(n63) );
  XOR2D0 U40 ( .A1(n66), .A2(n67), .Z(n65) );
  XOR2D0 U41 ( .A1(n[408]), .A2(n68), .Z(n67) );
  XOR2D0 U42 ( .A1(n69), .A2(n70), .Z(n68) );
  XOR2D0 U43 ( .A1(n71), .A2(n72), .Z(n70) );
  XOR2D0 U44 ( .A1(n[401]), .A2(n73), .Z(n72) );
  XOR2D0 U45 ( .A1(n74), .A2(n75), .Z(n73) );
  XOR2D0 U46 ( .A1(n76), .A2(n77), .Z(n75) );
  XOR2D0 U47 ( .A1(n[394]), .A2(n78), .Z(n77) );
  XOR2D0 U48 ( .A1(n79), .A2(n80), .Z(n78) );
  XOR2D0 U49 ( .A1(n81), .A2(n82), .Z(n80) );
  XOR2D0 U50 ( .A1(n[387]), .A2(n83), .Z(n82) );
  XOR2D0 U51 ( .A1(n84), .A2(n85), .Z(n83) );
  XOR2D0 U52 ( .A1(n86), .A2(n87), .Z(n85) );
  XOR2D0 U53 ( .A1(n[380]), .A2(n88), .Z(n87) );
  XOR2D0 U54 ( .A1(n89), .A2(n90), .Z(n88) );
  XOR2D0 U55 ( .A1(n91), .A2(n92), .Z(n90) );
  XOR2D0 U56 ( .A1(n[373]), .A2(n93), .Z(n92) );
  XOR2D0 U57 ( .A1(n94), .A2(n95), .Z(n93) );
  XOR2D0 U58 ( .A1(n96), .A2(n97), .Z(n95) );
  XOR2D0 U59 ( .A1(n[366]), .A2(n98), .Z(n97) );
  XOR2D0 U60 ( .A1(n99), .A2(n100), .Z(n98) );
  XOR2D0 U61 ( .A1(n101), .A2(n102), .Z(n100) );
  XOR2D0 U62 ( .A1(n[359]), .A2(n103), .Z(n102) );
  XOR2D0 U63 ( .A1(n104), .A2(n105), .Z(n103) );
  XOR2D0 U64 ( .A1(n106), .A2(n107), .Z(n105) );
  XOR2D0 U65 ( .A1(n[352]), .A2(n108), .Z(n107) );
  XOR2D0 U66 ( .A1(n109), .A2(n110), .Z(n108) );
  XOR2D0 U67 ( .A1(n111), .A2(n112), .Z(n110) );
  XOR2D0 U68 ( .A1(n[345]), .A2(n113), .Z(n112) );
  XOR2D0 U69 ( .A1(n114), .A2(n115), .Z(n113) );
  XOR2D0 U70 ( .A1(n116), .A2(n117), .Z(n115) );
  XOR2D0 U71 ( .A1(n[338]), .A2(n118), .Z(n117) );
  XOR2D0 U72 ( .A1(n119), .A2(n120), .Z(n118) );
  XOR2D0 U73 ( .A1(n121), .A2(n122), .Z(n120) );
  XOR2D0 U74 ( .A1(n[331]), .A2(n123), .Z(n122) );
  XOR2D0 U75 ( .A1(n124), .A2(n125), .Z(n123) );
  XOR2D0 U76 ( .A1(n126), .A2(n127), .Z(n125) );
  XOR2D0 U77 ( .A1(n[324]), .A2(n128), .Z(n127) );
  XOR2D0 U78 ( .A1(n129), .A2(n130), .Z(n128) );
  XOR2D0 U79 ( .A1(n131), .A2(n132), .Z(n130) );
  XOR2D0 U80 ( .A1(n[317]), .A2(n133), .Z(n132) );
  XOR2D0 U81 ( .A1(n134), .A2(n135), .Z(n133) );
  XOR2D0 U82 ( .A1(n136), .A2(n137), .Z(n135) );
  XOR2D0 U83 ( .A1(n[310]), .A2(n138), .Z(n137) );
  XOR2D0 U84 ( .A1(n139), .A2(n140), .Z(n138) );
  XOR2D0 U85 ( .A1(n141), .A2(n142), .Z(n140) );
  XOR2D0 U86 ( .A1(n[303]), .A2(n143), .Z(n142) );
  XOR2D0 U87 ( .A1(n144), .A2(n145), .Z(n143) );
  XOR2D0 U88 ( .A1(n146), .A2(n147), .Z(n145) );
  XOR2D0 U89 ( .A1(n[296]), .A2(n148), .Z(n147) );
  XOR2D0 U90 ( .A1(n149), .A2(n150), .Z(n148) );
  XOR2D0 U91 ( .A1(n151), .A2(n152), .Z(n150) );
  XOR2D0 U92 ( .A1(n[289]), .A2(n153), .Z(n152) );
  XOR2D0 U93 ( .A1(n154), .A2(n155), .Z(n153) );
  XOR2D0 U94 ( .A1(n156), .A2(n157), .Z(n155) );
  XOR2D0 U95 ( .A1(n[282]), .A2(n158), .Z(n157) );
  XOR2D0 U96 ( .A1(n159), .A2(n160), .Z(n158) );
  XOR2D0 U97 ( .A1(n161), .A2(n162), .Z(n160) );
  XOR2D0 U98 ( .A1(n[275]), .A2(n163), .Z(n162) );
  XOR2D0 U99 ( .A1(n164), .A2(n165), .Z(n163) );
  XOR2D0 U100 ( .A1(n166), .A2(n167), .Z(n165) );
  XOR2D0 U101 ( .A1(n[268]), .A2(n168), .Z(n167) );
  XOR2D0 U102 ( .A1(n169), .A2(n170), .Z(n168) );
  XOR2D0 U103 ( .A1(n171), .A2(n172), .Z(n170) );
  XOR2D0 U104 ( .A1(n[261]), .A2(n173), .Z(n172) );
  XOR2D0 U105 ( .A1(n174), .A2(n175), .Z(n173) );
  XOR2D0 U106 ( .A1(n176), .A2(n177), .Z(n175) );
  XOR2D0 U107 ( .A1(n[254]), .A2(n178), .Z(n177) );
  XOR2D0 U108 ( .A1(n179), .A2(n180), .Z(n178) );
  XOR2D0 U109 ( .A1(n181), .A2(n182), .Z(n180) );
  XOR2D0 U110 ( .A1(n[247]), .A2(n[246]), .Z(n182) );
  XOR2D0 U111 ( .A1(n[249]), .A2(n[248]), .Z(n181) );
  XOR2D0 U112 ( .A1(n183), .A2(n184), .Z(n179) );
  XOR2D0 U113 ( .A1(n[251]), .A2(n[250]), .Z(n184) );
  XOR2D0 U114 ( .A1(n[253]), .A2(n[252]), .Z(n183) );
  XOR2D0 U115 ( .A1(n[256]), .A2(n[255]), .Z(n176) );
  XOR2D0 U116 ( .A1(n185), .A2(n186), .Z(n174) );
  XOR2D0 U117 ( .A1(n[258]), .A2(n[257]), .Z(n186) );
  XOR2D0 U118 ( .A1(n[260]), .A2(n[259]), .Z(n185) );
  XOR2D0 U119 ( .A1(n[263]), .A2(n[262]), .Z(n171) );
  XOR2D0 U120 ( .A1(n187), .A2(n188), .Z(n169) );
  XOR2D0 U121 ( .A1(n[265]), .A2(n[264]), .Z(n188) );
  XOR2D0 U122 ( .A1(n[267]), .A2(n[266]), .Z(n187) );
  XOR2D0 U123 ( .A1(n[270]), .A2(n[269]), .Z(n166) );
  XOR2D0 U124 ( .A1(n189), .A2(n190), .Z(n164) );
  XOR2D0 U125 ( .A1(n[272]), .A2(n[271]), .Z(n190) );
  XOR2D0 U126 ( .A1(n[274]), .A2(n[273]), .Z(n189) );
  XOR2D0 U127 ( .A1(n[277]), .A2(n[276]), .Z(n161) );
  XOR2D0 U128 ( .A1(n191), .A2(n192), .Z(n159) );
  XOR2D0 U129 ( .A1(n[279]), .A2(n[278]), .Z(n192) );
  XOR2D0 U130 ( .A1(n[281]), .A2(n[280]), .Z(n191) );
  XOR2D0 U131 ( .A1(n[284]), .A2(n[283]), .Z(n156) );
  XOR2D0 U132 ( .A1(n193), .A2(n194), .Z(n154) );
  XOR2D0 U133 ( .A1(n[286]), .A2(n[285]), .Z(n194) );
  XOR2D0 U134 ( .A1(n[288]), .A2(n[287]), .Z(n193) );
  XOR2D0 U135 ( .A1(n[291]), .A2(n[290]), .Z(n151) );
  XOR2D0 U136 ( .A1(n195), .A2(n196), .Z(n149) );
  XOR2D0 U137 ( .A1(n[293]), .A2(n[292]), .Z(n196) );
  XOR2D0 U138 ( .A1(n[295]), .A2(n[294]), .Z(n195) );
  XOR2D0 U139 ( .A1(n[298]), .A2(n[297]), .Z(n146) );
  XOR2D0 U140 ( .A1(n197), .A2(n198), .Z(n144) );
  XOR2D0 U141 ( .A1(n[300]), .A2(n[299]), .Z(n198) );
  XOR2D0 U142 ( .A1(n[302]), .A2(n[301]), .Z(n197) );
  XOR2D0 U143 ( .A1(n[305]), .A2(n[304]), .Z(n141) );
  XOR2D0 U144 ( .A1(n199), .A2(n200), .Z(n139) );
  XOR2D0 U145 ( .A1(n[307]), .A2(n[306]), .Z(n200) );
  XOR2D0 U146 ( .A1(n[309]), .A2(n[308]), .Z(n199) );
  XOR2D0 U147 ( .A1(n[312]), .A2(n[311]), .Z(n136) );
  XOR2D0 U148 ( .A1(n201), .A2(n202), .Z(n134) );
  XOR2D0 U149 ( .A1(n[314]), .A2(n[313]), .Z(n202) );
  XOR2D0 U150 ( .A1(n[316]), .A2(n[315]), .Z(n201) );
  XOR2D0 U151 ( .A1(n[319]), .A2(n[318]), .Z(n131) );
  XOR2D0 U152 ( .A1(n203), .A2(n204), .Z(n129) );
  XOR2D0 U153 ( .A1(n[321]), .A2(n[320]), .Z(n204) );
  XOR2D0 U154 ( .A1(n[323]), .A2(n[322]), .Z(n203) );
  XOR2D0 U155 ( .A1(n[326]), .A2(n[325]), .Z(n126) );
  XOR2D0 U156 ( .A1(n205), .A2(n206), .Z(n124) );
  XOR2D0 U157 ( .A1(n[328]), .A2(n[327]), .Z(n206) );
  XOR2D0 U158 ( .A1(n[330]), .A2(n[329]), .Z(n205) );
  XOR2D0 U159 ( .A1(n[333]), .A2(n[332]), .Z(n121) );
  XOR2D0 U160 ( .A1(n207), .A2(n208), .Z(n119) );
  XOR2D0 U161 ( .A1(n[335]), .A2(n[334]), .Z(n208) );
  XOR2D0 U162 ( .A1(n[337]), .A2(n[336]), .Z(n207) );
  XOR2D0 U163 ( .A1(n[340]), .A2(n[339]), .Z(n116) );
  XOR2D0 U164 ( .A1(n209), .A2(n210), .Z(n114) );
  XOR2D0 U165 ( .A1(n[342]), .A2(n[341]), .Z(n210) );
  XOR2D0 U166 ( .A1(n[344]), .A2(n[343]), .Z(n209) );
  XOR2D0 U167 ( .A1(n[347]), .A2(n[346]), .Z(n111) );
  XOR2D0 U168 ( .A1(n211), .A2(n212), .Z(n109) );
  XOR2D0 U169 ( .A1(n[349]), .A2(n[348]), .Z(n212) );
  XOR2D0 U170 ( .A1(n[351]), .A2(n[350]), .Z(n211) );
  XOR2D0 U171 ( .A1(n[354]), .A2(n[353]), .Z(n106) );
  XOR2D0 U172 ( .A1(n213), .A2(n214), .Z(n104) );
  XOR2D0 U173 ( .A1(n[356]), .A2(n[355]), .Z(n214) );
  XOR2D0 U174 ( .A1(n[358]), .A2(n[357]), .Z(n213) );
  XOR2D0 U175 ( .A1(n[361]), .A2(n[360]), .Z(n101) );
  XOR2D0 U176 ( .A1(n215), .A2(n216), .Z(n99) );
  XOR2D0 U177 ( .A1(n[363]), .A2(n[362]), .Z(n216) );
  XOR2D0 U178 ( .A1(n[365]), .A2(n[364]), .Z(n215) );
  XOR2D0 U179 ( .A1(n[368]), .A2(n[367]), .Z(n96) );
  XOR2D0 U180 ( .A1(n217), .A2(n218), .Z(n94) );
  XOR2D0 U181 ( .A1(n[370]), .A2(n[369]), .Z(n218) );
  XOR2D0 U182 ( .A1(n[372]), .A2(n[371]), .Z(n217) );
  XOR2D0 U183 ( .A1(n[375]), .A2(n[374]), .Z(n91) );
  XOR2D0 U184 ( .A1(n219), .A2(n220), .Z(n89) );
  XOR2D0 U185 ( .A1(n[377]), .A2(n[376]), .Z(n220) );
  XOR2D0 U186 ( .A1(n[379]), .A2(n[378]), .Z(n219) );
  XOR2D0 U187 ( .A1(n[382]), .A2(n[381]), .Z(n86) );
  XOR2D0 U188 ( .A1(n221), .A2(n222), .Z(n84) );
  XOR2D0 U189 ( .A1(n[384]), .A2(n[383]), .Z(n222) );
  XOR2D0 U190 ( .A1(n[386]), .A2(n[385]), .Z(n221) );
  XOR2D0 U191 ( .A1(n[389]), .A2(n[388]), .Z(n81) );
  XOR2D0 U192 ( .A1(n223), .A2(n224), .Z(n79) );
  XOR2D0 U193 ( .A1(n[391]), .A2(n[390]), .Z(n224) );
  XOR2D0 U194 ( .A1(n[393]), .A2(n[392]), .Z(n223) );
  XOR2D0 U195 ( .A1(n[396]), .A2(n[395]), .Z(n76) );
  XOR2D0 U196 ( .A1(n225), .A2(n226), .Z(n74) );
  XOR2D0 U197 ( .A1(n[398]), .A2(n[397]), .Z(n226) );
  XOR2D0 U198 ( .A1(n[400]), .A2(n[399]), .Z(n225) );
  XOR2D0 U199 ( .A1(n[403]), .A2(n[402]), .Z(n71) );
  XOR2D0 U200 ( .A1(n227), .A2(n228), .Z(n69) );
  XOR2D0 U201 ( .A1(n[405]), .A2(n[404]), .Z(n228) );
  XOR2D0 U202 ( .A1(n[407]), .A2(n[406]), .Z(n227) );
  XOR2D0 U203 ( .A1(n[410]), .A2(n[409]), .Z(n66) );
  XOR2D0 U204 ( .A1(n229), .A2(n230), .Z(n64) );
  XOR2D0 U205 ( .A1(n[412]), .A2(n[411]), .Z(n230) );
  XOR2D0 U206 ( .A1(n[414]), .A2(n[413]), .Z(n229) );
  XOR2D0 U207 ( .A1(n[417]), .A2(n[416]), .Z(n61) );
  XOR2D0 U208 ( .A1(n231), .A2(n232), .Z(n59) );
  XOR2D0 U209 ( .A1(n[419]), .A2(n[418]), .Z(n232) );
  XOR2D0 U210 ( .A1(n[421]), .A2(n[420]), .Z(n231) );
  XOR2D0 U211 ( .A1(n[424]), .A2(n[423]), .Z(n56) );
  XOR2D0 U212 ( .A1(n233), .A2(n234), .Z(n54) );
  XOR2D0 U213 ( .A1(n[426]), .A2(n[425]), .Z(n234) );
  XOR2D0 U214 ( .A1(n[428]), .A2(n[427]), .Z(n233) );
  XOR2D0 U215 ( .A1(n[431]), .A2(n[430]), .Z(n51) );
  XOR2D0 U216 ( .A1(n235), .A2(n236), .Z(n49) );
  XOR2D0 U217 ( .A1(n[433]), .A2(n[432]), .Z(n236) );
  XOR2D0 U218 ( .A1(n[435]), .A2(n[434]), .Z(n235) );
  XOR2D0 U219 ( .A1(n[438]), .A2(n[437]), .Z(n46) );
  XOR2D0 U220 ( .A1(n237), .A2(n238), .Z(n44) );
  XOR2D0 U221 ( .A1(n[440]), .A2(n[439]), .Z(n238) );
  XOR2D0 U222 ( .A1(n[442]), .A2(n[441]), .Z(n237) );
  XOR2D0 U223 ( .A1(n[445]), .A2(n[444]), .Z(n41) );
  XOR2D0 U224 ( .A1(n239), .A2(n240), .Z(n39) );
  XOR2D0 U225 ( .A1(n[447]), .A2(n[446]), .Z(n240) );
  XOR2D0 U226 ( .A1(n[449]), .A2(n[448]), .Z(n239) );
  XOR2D0 U227 ( .A1(n[452]), .A2(n[451]), .Z(n36) );
  XOR2D0 U228 ( .A1(n241), .A2(n242), .Z(n34) );
  XOR2D0 U229 ( .A1(n[454]), .A2(n[453]), .Z(n242) );
  XOR2D0 U230 ( .A1(n[456]), .A2(n[455]), .Z(n241) );
  XOR2D0 U231 ( .A1(n[459]), .A2(n[458]), .Z(n31) );
  XOR2D0 U232 ( .A1(n243), .A2(n244), .Z(n29) );
  XOR2D0 U233 ( .A1(n[461]), .A2(n[460]), .Z(n244) );
  XOR2D0 U234 ( .A1(n[463]), .A2(n[462]), .Z(n243) );
  XOR2D0 U235 ( .A1(n[466]), .A2(n[465]), .Z(n26) );
  XOR2D0 U236 ( .A1(n245), .A2(n246), .Z(n24) );
  XOR2D0 U237 ( .A1(n[468]), .A2(n[467]), .Z(n246) );
  XOR2D0 U238 ( .A1(n[470]), .A2(n[469]), .Z(n245) );
  XOR2D0 U239 ( .A1(n[473]), .A2(n[472]), .Z(n21) );
  XOR2D0 U240 ( .A1(n247), .A2(n248), .Z(n19) );
  XOR2D0 U241 ( .A1(n[475]), .A2(n[474]), .Z(n248) );
  XOR2D0 U242 ( .A1(n[477]), .A2(n[476]), .Z(n247) );
  XOR2D0 U243 ( .A1(n[480]), .A2(n[479]), .Z(n16) );
  XOR2D0 U244 ( .A1(n249), .A2(n250), .Z(n14) );
  XOR2D0 U245 ( .A1(n[482]), .A2(n[481]), .Z(n250) );
  XOR2D0 U246 ( .A1(n[484]), .A2(n[483]), .Z(n249) );
  XOR2D0 U247 ( .A1(n[487]), .A2(n[486]), .Z(n11) );
  XOR2D0 U248 ( .A1(n251), .A2(n252), .Z(n9) );
  XOR2D0 U249 ( .A1(n[489]), .A2(n[488]), .Z(n252) );
  XOR2D0 U250 ( .A1(n[491]), .A2(n[490]), .Z(n251) );
  XOR2D0 U251 ( .A1(n[494]), .A2(n[493]), .Z(n6) );
  XOR2D0 U252 ( .A1(n253), .A2(n254), .Z(n4) );
  XOR2D0 U253 ( .A1(n[496]), .A2(n[495]), .Z(n254) );
  XOR2D0 U254 ( .A1(n[498]), .A2(n[497]), .Z(n253) );
  XOR2D0 U255 ( .A1(b[7]), .A2(n255), .Z(n1) );
  XOR2D0 U256 ( .A1(n[500]), .A2(n[499]), .Z(n255) );
  XOR2D0 U257 ( .A1(n256), .A2(n257), .Z(s[6]) );
  XOR2D0 U258 ( .A1(b[6]), .A2(a[6]), .Z(n257) );
  XOR2D0 U259 ( .A1(n258), .A2(n259), .Z(n256) );
  XOR2D0 U260 ( .A1(n260), .A2(n261), .Z(n259) );
  XOR2D0 U261 ( .A1(n[239]), .A2(n262), .Z(n261) );
  XOR2D0 U262 ( .A1(n263), .A2(n264), .Z(n262) );
  XOR2D0 U263 ( .A1(n265), .A2(n266), .Z(n264) );
  XOR2D0 U264 ( .A1(n[232]), .A2(n267), .Z(n266) );
  XOR2D0 U265 ( .A1(n268), .A2(n269), .Z(n267) );
  XOR2D0 U266 ( .A1(n270), .A2(n271), .Z(n269) );
  XOR2D0 U267 ( .A1(n[225]), .A2(n272), .Z(n271) );
  XOR2D0 U268 ( .A1(n273), .A2(n274), .Z(n272) );
  XOR2D0 U269 ( .A1(n275), .A2(n276), .Z(n274) );
  XOR2D0 U270 ( .A1(n[218]), .A2(n277), .Z(n276) );
  XOR2D0 U271 ( .A1(n278), .A2(n279), .Z(n277) );
  XOR2D0 U272 ( .A1(n280), .A2(n281), .Z(n279) );
  XOR2D0 U273 ( .A1(n[211]), .A2(n282), .Z(n281) );
  XOR2D0 U274 ( .A1(n283), .A2(n284), .Z(n282) );
  XOR2D0 U275 ( .A1(n285), .A2(n286), .Z(n284) );
  XOR2D0 U276 ( .A1(n[204]), .A2(n287), .Z(n286) );
  XOR2D0 U277 ( .A1(n288), .A2(n289), .Z(n287) );
  XOR2D0 U278 ( .A1(n290), .A2(n291), .Z(n289) );
  XOR2D0 U279 ( .A1(n[197]), .A2(n292), .Z(n291) );
  XOR2D0 U280 ( .A1(n293), .A2(n294), .Z(n292) );
  XOR2D0 U281 ( .A1(n295), .A2(n296), .Z(n294) );
  XOR2D0 U282 ( .A1(n[190]), .A2(n297), .Z(n296) );
  XOR2D0 U283 ( .A1(n298), .A2(n299), .Z(n297) );
  XOR2D0 U284 ( .A1(n300), .A2(n301), .Z(n299) );
  XOR2D0 U285 ( .A1(n[183]), .A2(n302), .Z(n301) );
  XOR2D0 U286 ( .A1(n303), .A2(n304), .Z(n302) );
  XOR2D0 U287 ( .A1(n305), .A2(n306), .Z(n304) );
  XOR2D0 U288 ( .A1(n[176]), .A2(n307), .Z(n306) );
  XOR2D0 U289 ( .A1(n308), .A2(n309), .Z(n307) );
  XOR2D0 U290 ( .A1(n310), .A2(n311), .Z(n309) );
  XOR2D0 U291 ( .A1(n[169]), .A2(n312), .Z(n311) );
  XOR2D0 U292 ( .A1(n313), .A2(n314), .Z(n312) );
  XOR2D0 U293 ( .A1(n315), .A2(n316), .Z(n314) );
  XOR2D0 U294 ( .A1(n[162]), .A2(n317), .Z(n316) );
  XOR2D0 U295 ( .A1(n318), .A2(n319), .Z(n317) );
  XOR2D0 U296 ( .A1(n320), .A2(n321), .Z(n319) );
  XOR2D0 U297 ( .A1(n[155]), .A2(n322), .Z(n321) );
  XOR2D0 U298 ( .A1(n323), .A2(n324), .Z(n322) );
  XOR2D0 U299 ( .A1(n325), .A2(n326), .Z(n324) );
  XOR2D0 U300 ( .A1(n[148]), .A2(n327), .Z(n326) );
  XOR2D0 U301 ( .A1(n328), .A2(n329), .Z(n327) );
  XOR2D0 U302 ( .A1(n330), .A2(n331), .Z(n329) );
  XOR2D0 U303 ( .A1(n[141]), .A2(n332), .Z(n331) );
  XOR2D0 U304 ( .A1(n333), .A2(n334), .Z(n332) );
  XOR2D0 U305 ( .A1(n335), .A2(n336), .Z(n334) );
  XOR2D0 U306 ( .A1(n[134]), .A2(n337), .Z(n336) );
  XOR2D0 U307 ( .A1(n338), .A2(n339), .Z(n337) );
  XOR2D0 U308 ( .A1(n340), .A2(n341), .Z(n339) );
  XOR2D0 U309 ( .A1(n[127]), .A2(n342), .Z(n341) );
  XOR2D0 U310 ( .A1(n343), .A2(n344), .Z(n342) );
  XOR2D0 U311 ( .A1(n345), .A2(n346), .Z(n344) );
  XOR2D0 U312 ( .A1(n[120]), .A2(n[119]), .Z(n346) );
  XOR2D0 U313 ( .A1(n[122]), .A2(n[121]), .Z(n345) );
  XOR2D0 U314 ( .A1(n347), .A2(n348), .Z(n343) );
  XOR2D0 U315 ( .A1(n[124]), .A2(n[123]), .Z(n348) );
  XOR2D0 U316 ( .A1(n[126]), .A2(n[125]), .Z(n347) );
  XOR2D0 U317 ( .A1(n[129]), .A2(n[128]), .Z(n340) );
  XOR2D0 U318 ( .A1(n349), .A2(n350), .Z(n338) );
  XOR2D0 U319 ( .A1(n[131]), .A2(n[130]), .Z(n350) );
  XOR2D0 U320 ( .A1(n[133]), .A2(n[132]), .Z(n349) );
  XOR2D0 U321 ( .A1(n[136]), .A2(n[135]), .Z(n335) );
  XOR2D0 U322 ( .A1(n351), .A2(n352), .Z(n333) );
  XOR2D0 U323 ( .A1(n[138]), .A2(n[137]), .Z(n352) );
  XOR2D0 U324 ( .A1(n[140]), .A2(n[139]), .Z(n351) );
  XOR2D0 U325 ( .A1(n[143]), .A2(n[142]), .Z(n330) );
  XOR2D0 U326 ( .A1(n353), .A2(n354), .Z(n328) );
  XOR2D0 U327 ( .A1(n[145]), .A2(n[144]), .Z(n354) );
  XOR2D0 U328 ( .A1(n[147]), .A2(n[146]), .Z(n353) );
  XOR2D0 U329 ( .A1(n[150]), .A2(n[149]), .Z(n325) );
  XOR2D0 U330 ( .A1(n355), .A2(n356), .Z(n323) );
  XOR2D0 U331 ( .A1(n[152]), .A2(n[151]), .Z(n356) );
  XOR2D0 U332 ( .A1(n[154]), .A2(n[153]), .Z(n355) );
  XOR2D0 U333 ( .A1(n[157]), .A2(n[156]), .Z(n320) );
  XOR2D0 U334 ( .A1(n357), .A2(n358), .Z(n318) );
  XOR2D0 U335 ( .A1(n[159]), .A2(n[158]), .Z(n358) );
  XOR2D0 U336 ( .A1(n[161]), .A2(n[160]), .Z(n357) );
  XOR2D0 U337 ( .A1(n[164]), .A2(n[163]), .Z(n315) );
  XOR2D0 U338 ( .A1(n359), .A2(n360), .Z(n313) );
  XOR2D0 U339 ( .A1(n[166]), .A2(n[165]), .Z(n360) );
  XOR2D0 U340 ( .A1(n[168]), .A2(n[167]), .Z(n359) );
  XOR2D0 U341 ( .A1(n[171]), .A2(n[170]), .Z(n310) );
  XOR2D0 U342 ( .A1(n361), .A2(n362), .Z(n308) );
  XOR2D0 U343 ( .A1(n[173]), .A2(n[172]), .Z(n362) );
  XOR2D0 U344 ( .A1(n[175]), .A2(n[174]), .Z(n361) );
  XOR2D0 U345 ( .A1(n[178]), .A2(n[177]), .Z(n305) );
  XOR2D0 U346 ( .A1(n363), .A2(n364), .Z(n303) );
  XOR2D0 U347 ( .A1(n[180]), .A2(n[179]), .Z(n364) );
  XOR2D0 U348 ( .A1(n[182]), .A2(n[181]), .Z(n363) );
  XOR2D0 U349 ( .A1(n[185]), .A2(n[184]), .Z(n300) );
  XOR2D0 U350 ( .A1(n365), .A2(n366), .Z(n298) );
  XOR2D0 U351 ( .A1(n[187]), .A2(n[186]), .Z(n366) );
  XOR2D0 U352 ( .A1(n[189]), .A2(n[188]), .Z(n365) );
  XOR2D0 U353 ( .A1(n[192]), .A2(n[191]), .Z(n295) );
  XOR2D0 U354 ( .A1(n367), .A2(n368), .Z(n293) );
  XOR2D0 U355 ( .A1(n[194]), .A2(n[193]), .Z(n368) );
  XOR2D0 U356 ( .A1(n[196]), .A2(n[195]), .Z(n367) );
  XOR2D0 U357 ( .A1(n[199]), .A2(n[198]), .Z(n290) );
  XOR2D0 U358 ( .A1(n369), .A2(n370), .Z(n288) );
  XOR2D0 U359 ( .A1(n[201]), .A2(n[200]), .Z(n370) );
  XOR2D0 U360 ( .A1(n[203]), .A2(n[202]), .Z(n369) );
  XOR2D0 U361 ( .A1(n[206]), .A2(n[205]), .Z(n285) );
  XOR2D0 U362 ( .A1(n371), .A2(n372), .Z(n283) );
  XOR2D0 U363 ( .A1(n[208]), .A2(n[207]), .Z(n372) );
  XOR2D0 U364 ( .A1(n[210]), .A2(n[209]), .Z(n371) );
  XOR2D0 U365 ( .A1(n[213]), .A2(n[212]), .Z(n280) );
  XOR2D0 U366 ( .A1(n373), .A2(n374), .Z(n278) );
  XOR2D0 U367 ( .A1(n[215]), .A2(n[214]), .Z(n374) );
  XOR2D0 U368 ( .A1(n[217]), .A2(n[216]), .Z(n373) );
  XOR2D0 U369 ( .A1(n[220]), .A2(n[219]), .Z(n275) );
  XOR2D0 U370 ( .A1(n375), .A2(n376), .Z(n273) );
  XOR2D0 U371 ( .A1(n[222]), .A2(n[221]), .Z(n376) );
  XOR2D0 U372 ( .A1(n[224]), .A2(n[223]), .Z(n375) );
  XOR2D0 U373 ( .A1(n[227]), .A2(n[226]), .Z(n270) );
  XOR2D0 U374 ( .A1(n377), .A2(n378), .Z(n268) );
  XOR2D0 U375 ( .A1(n[229]), .A2(n[228]), .Z(n378) );
  XOR2D0 U376 ( .A1(n[231]), .A2(n[230]), .Z(n377) );
  XOR2D0 U377 ( .A1(n[234]), .A2(n[233]), .Z(n265) );
  XOR2D0 U378 ( .A1(n379), .A2(n380), .Z(n263) );
  XOR2D0 U379 ( .A1(n[236]), .A2(n[235]), .Z(n380) );
  XOR2D0 U380 ( .A1(n[238]), .A2(n[237]), .Z(n379) );
  XOR2D0 U381 ( .A1(n[241]), .A2(n[240]), .Z(n260) );
  XOR2D0 U382 ( .A1(n381), .A2(n382), .Z(n258) );
  XOR2D0 U383 ( .A1(n[243]), .A2(n[242]), .Z(n382) );
  XOR2D0 U384 ( .A1(n[245]), .A2(n[244]), .Z(n381) );
  XOR2D0 U385 ( .A1(n383), .A2(n384), .Z(s[5]) );
  XOR2D0 U386 ( .A1(n[115]), .A2(n385), .Z(n384) );
  XOR2D0 U387 ( .A1(n386), .A2(n387), .Z(n385) );
  XOR2D0 U388 ( .A1(a[5]), .A2(n388), .Z(n387) );
  XOR2D0 U389 ( .A1(n389), .A2(n390), .Z(n388) );
  XOR2D0 U390 ( .A1(n391), .A2(n392), .Z(n390) );
  XOR2D0 U391 ( .A1(n[106]), .A2(n393), .Z(n392) );
  XOR2D0 U392 ( .A1(n394), .A2(n395), .Z(n393) );
  XOR2D0 U393 ( .A1(n396), .A2(n397), .Z(n395) );
  XOR2D0 U394 ( .A1(n[100]), .A2(n398), .Z(n397) );
  XOR2D0 U395 ( .A1(n399), .A2(n400), .Z(n398) );
  XOR2D0 U396 ( .A1(n401), .A2(n402), .Z(n400) );
  XOR2D0 U397 ( .A1(n[92]), .A2(n403), .Z(n402) );
  XOR2D0 U398 ( .A1(n404), .A2(n405), .Z(n403) );
  XOR2D0 U399 ( .A1(n406), .A2(n407), .Z(n405) );
  XOR2D0 U400 ( .A1(n[85]), .A2(n408), .Z(n407) );
  XOR2D0 U401 ( .A1(n409), .A2(n410), .Z(n408) );
  XOR2D0 U402 ( .A1(n411), .A2(n412), .Z(n410) );
  XOR2D0 U403 ( .A1(n[78]), .A2(n413), .Z(n412) );
  XOR2D0 U404 ( .A1(n414), .A2(n415), .Z(n413) );
  XOR2D0 U405 ( .A1(n416), .A2(n417), .Z(n415) );
  XOR2D0 U406 ( .A1(n[71]), .A2(n418), .Z(n417) );
  XOR2D0 U407 ( .A1(n419), .A2(n420), .Z(n418) );
  XOR2D0 U408 ( .A1(n421), .A2(n422), .Z(n420) );
  XOR2D0 U409 ( .A1(n[64]), .A2(n423), .Z(n422) );
  XOR2D0 U410 ( .A1(n424), .A2(n425), .Z(n423) );
  XOR2D0 U411 ( .A1(n426), .A2(n427), .Z(n425) );
  XOR2D0 U412 ( .A1(n[57]), .A2(n[56]), .Z(n427) );
  XOR2D0 U413 ( .A1(n[59]), .A2(n[58]), .Z(n426) );
  XOR2D0 U414 ( .A1(n428), .A2(n429), .Z(n424) );
  XOR2D0 U415 ( .A1(n[61]), .A2(n[60]), .Z(n429) );
  XOR2D0 U416 ( .A1(n[63]), .A2(n[62]), .Z(n428) );
  XOR2D0 U417 ( .A1(n[66]), .A2(n[65]), .Z(n421) );
  XOR2D0 U418 ( .A1(n430), .A2(n431), .Z(n419) );
  XOR2D0 U419 ( .A1(n[68]), .A2(n[67]), .Z(n431) );
  XOR2D0 U420 ( .A1(n[70]), .A2(n[69]), .Z(n430) );
  XOR2D0 U421 ( .A1(n[73]), .A2(n[72]), .Z(n416) );
  XOR2D0 U422 ( .A1(n432), .A2(n433), .Z(n414) );
  XOR2D0 U423 ( .A1(n[75]), .A2(n[74]), .Z(n433) );
  XOR2D0 U424 ( .A1(n[77]), .A2(n[76]), .Z(n432) );
  XOR2D0 U425 ( .A1(n[80]), .A2(n[79]), .Z(n411) );
  XOR2D0 U426 ( .A1(n434), .A2(n435), .Z(n409) );
  XOR2D0 U427 ( .A1(n[82]), .A2(n[81]), .Z(n435) );
  XOR2D0 U428 ( .A1(n[84]), .A2(n[83]), .Z(n434) );
  XOR2D0 U429 ( .A1(n[87]), .A2(n[86]), .Z(n406) );
  XOR2D0 U430 ( .A1(n436), .A2(n437), .Z(n404) );
  XOR2D0 U431 ( .A1(n[89]), .A2(n[88]), .Z(n437) );
  XOR2D0 U432 ( .A1(n[91]), .A2(n[90]), .Z(n436) );
  XOR2D0 U433 ( .A1(n[94]), .A2(n[93]), .Z(n401) );
  XOR2D0 U434 ( .A1(n438), .A2(n439), .Z(n399) );
  XOR2D0 U435 ( .A1(n[96]), .A2(n[95]), .Z(n439) );
  XOR2D0 U436 ( .A1(n[98]), .A2(n[97]), .Z(n438) );
  XOR2D0 U437 ( .A1(n[102]), .A2(n[101]), .Z(n396) );
  XOR2D0 U438 ( .A1(n440), .A2(n441), .Z(n394) );
  XOR2D0 U439 ( .A1(n[104]), .A2(n[103]), .Z(n441) );
  XOR2D0 U440 ( .A1(n[99]), .A2(n[105]), .Z(n440) );
  XOR2D0 U441 ( .A1(n[108]), .A2(n[107]), .Z(n391) );
  XOR2D0 U442 ( .A1(n442), .A2(n443), .Z(n389) );
  XOR2D0 U443 ( .A1(n[110]), .A2(n[109]), .Z(n443) );
  XOR2D0 U444 ( .A1(n[112]), .A2(n[111]), .Z(n442) );
  XOR2D0 U445 ( .A1(b[5]), .A2(n444), .Z(n386) );
  XOR2D0 U446 ( .A1(n[114]), .A2(n[113]), .Z(n444) );
  XOR2D0 U447 ( .A1(n[116]), .A2(n445), .Z(n383) );
  XOR2D0 U448 ( .A1(n[118]), .A2(n[117]), .Z(n445) );
  XOR2D0 U449 ( .A1(n446), .A2(n447), .Z(s[4]) );
  XOR2D0 U450 ( .A1(a[4]), .A2(n448), .Z(n447) );
  XOR2D0 U451 ( .A1(n449), .A2(n450), .Z(n448) );
  XOR2D0 U452 ( .A1(n451), .A2(n452), .Z(n450) );
  XOR2D0 U453 ( .A1(n[47]), .A2(n453), .Z(n452) );
  XOR2D0 U454 ( .A1(n454), .A2(n455), .Z(n453) );
  XOR2D0 U455 ( .A1(n456), .A2(n457), .Z(n455) );
  XOR2D0 U456 ( .A1(n[40]), .A2(n458), .Z(n457) );
  XOR2D0 U457 ( .A1(n459), .A2(n460), .Z(n458) );
  XOR2D0 U458 ( .A1(n461), .A2(n462), .Z(n460) );
  XOR2D0 U459 ( .A1(n[33]), .A2(n463), .Z(n462) );
  XOR2D0 U460 ( .A1(n464), .A2(n465), .Z(n463) );
  XOR2D0 U461 ( .A1(n466), .A2(n467), .Z(n465) );
  XOR2D0 U462 ( .A1(n[26]), .A2(n[25]), .Z(n467) );
  XOR2D0 U463 ( .A1(n[28]), .A2(n[27]), .Z(n466) );
  XOR2D0 U464 ( .A1(n468), .A2(n469), .Z(n464) );
  XOR2D0 U465 ( .A1(n[30]), .A2(n[29]), .Z(n469) );
  XOR2D0 U466 ( .A1(n[32]), .A2(n[31]), .Z(n468) );
  XOR2D0 U467 ( .A1(n[35]), .A2(n[34]), .Z(n461) );
  XOR2D0 U468 ( .A1(n470), .A2(n471), .Z(n459) );
  XOR2D0 U469 ( .A1(n[37]), .A2(n[36]), .Z(n471) );
  XOR2D0 U470 ( .A1(n[39]), .A2(n[38]), .Z(n470) );
  XOR2D0 U471 ( .A1(n[42]), .A2(n[41]), .Z(n456) );
  XOR2D0 U472 ( .A1(n472), .A2(n473), .Z(n454) );
  XOR2D0 U473 ( .A1(n[44]), .A2(n[43]), .Z(n473) );
  XOR2D0 U474 ( .A1(n[46]), .A2(n[45]), .Z(n472) );
  XOR2D0 U475 ( .A1(n[49]), .A2(n[48]), .Z(n451) );
  XOR2D0 U476 ( .A1(n474), .A2(n475), .Z(n449) );
  XOR2D0 U477 ( .A1(n[51]), .A2(n[50]), .Z(n475) );
  XOR2D0 U478 ( .A1(n[53]), .A2(n[52]), .Z(n474) );
  XOR2D0 U479 ( .A1(b[4]), .A2(n476), .Z(n446) );
  XOR2D0 U480 ( .A1(n[55]), .A2(n[54]), .Z(n476) );
  XOR2D0 U481 ( .A1(n477), .A2(n478), .Z(s[3]) );
  XOR2D0 U482 ( .A1(b[3]), .A2(a[3]), .Z(n478) );
  XOR2D0 U483 ( .A1(n479), .A2(n480), .Z(n477) );
  XOR2D0 U484 ( .A1(n481), .A2(n482), .Z(n480) );
  XOR2D0 U485 ( .A1(n[18]), .A2(n483), .Z(n482) );
  XOR2D0 U486 ( .A1(n484), .A2(n485), .Z(n483) );
  XOR2D0 U487 ( .A1(n486), .A2(n487), .Z(n485) );
  XOR2D0 U488 ( .A1(n[11]), .A2(n[10]), .Z(n487) );
  XOR2D0 U489 ( .A1(n[13]), .A2(n[12]), .Z(n486) );
  XOR2D0 U490 ( .A1(n488), .A2(n489), .Z(n484) );
  XOR2D0 U491 ( .A1(n[15]), .A2(n[14]), .Z(n489) );
  XOR2D0 U492 ( .A1(n[17]), .A2(n[16]), .Z(n488) );
  XOR2D0 U493 ( .A1(n[20]), .A2(n[19]), .Z(n481) );
  XOR2D0 U494 ( .A1(n490), .A2(n491), .Z(n479) );
  XOR2D0 U495 ( .A1(n[22]), .A2(n[21]), .Z(n491) );
  XOR2D0 U496 ( .A1(n[24]), .A2(n[23]), .Z(n490) );
  XOR2D0 U497 ( .A1(n492), .A2(n493), .Z(s[2]) );
  XOR2D0 U498 ( .A1(n[6]), .A2(n494), .Z(n493) );
  XOR2D0 U499 ( .A1(n495), .A2(n496), .Z(n494) );
  XOR2D0 U500 ( .A1(b[2]), .A2(a[2]), .Z(n496) );
  XOR2D0 U501 ( .A1(n[3]), .A2(n497), .Z(n495) );
  XOR2D0 U502 ( .A1(n[5]), .A2(n[4]), .Z(n497) );
  XOR2D0 U503 ( .A1(n[7]), .A2(n498), .Z(n492) );
  XOR2D0 U504 ( .A1(n[9]), .A2(n[8]), .Z(n498) );
  XOR2D0 U505 ( .A1(n499), .A2(n500), .Z(s[1]) );
  XOR2D0 U506 ( .A1(b[1]), .A2(a[1]), .Z(n500) );
  XOR2D0 U507 ( .A1(n[0]), .A2(n501), .Z(n499) );
  XOR2D0 U508 ( .A1(n[2]), .A2(n[1]), .Z(n501) );
  XOR2D0 U509 ( .A1(b[0]), .A2(a[0]), .Z(s[0]) );
endmodule


module gen_nonlinear_part ( a, b, n );
  input [7:0] a;
  input [7:0] b;
  output [501:0] n;
  wire   n_498, n_495, n_494, n_491, n_488, n_487, n_486, n_483, n_480, n_479,
         n_476, n_473, n_472, n_471, n_470, n_467, n_464, n_463, n_460, n_457,
         n_456, n_455, n_452, n_449, n_448, n_445, n_442, n_441, n_440, n_439,
         n_438, n_435, n_432, n_431, n_428, n_425, n_424, n_423, n_420, n_417,
         n_416, n_413, n_410, n_409, n_408, n_407, n_404, n_401, n_400, n_397,
         n_394, n_393, n_392, n_389, n_386, n_385, n_382, n_379, n_378, n_377,
         n_376, n_375, n_374, n_371, n_368, n_367, n_364, n_361, n_360, n_359,
         n_356, n_353, n_352, n_349, n_346, n_345, n_344, n_343, n_340, n_337,
         n_336, n_333, n_330, n_329, n_328, n_325, n_322, n_321, n_318, n_315,
         n_314, n_313, n_312, n_311, n_308, n_305, n_304, n_301, n_298, n_297,
         n_296, n_293, n_290, n_289, n_286, n_283, n_282, n_281, n_280, n_277,
         n_274, n_273, n_270, n_267, n_266, n_265, n_262, n_259, n_258, n_255,
         n_243, n_240, n_239, n_236, n_233, n_232, n_231, n_228, n_225, n_224,
         n_221, n_218, n_217, n_216, n_215, n_212, n_209, n_208, n_205, n_202,
         n_201, n_200, n_197, n_194, n_193, n_190, n_187, n_186, n_185, n_184,
         n_183, n_180, n_177, n_176, n_173, n_170, n_169, n_168, n_165, n_162,
         n_161, n_158, n_155, n_154, n_153, n_152, n_149, n_146, n_145, n_142,
         n_139, n_138, n_137, n_134, n_131, n_130, n_127, n_124, n_123, n_122,
         n_121, n_120, n_119, n_116, n_113, n_112, n_109, n_106, n_105, n_104,
         n_101, n_98, n_97, n_94, n_91, n_90, n_89, n_88, n_85, n_82, n_81,
         n_78, n_75, n_74, n_73, n_70, n_67, n_66, n_63, n_60, n_59, n_58,
         n_57, n_56, n_53, n_50, n_49, n_46, n_43, n_42, n_41, n_38, n_35,
         n_34, n_31, n_28, n_27, n_26, n_25, n_22, n_19, n_18, n_15, n_12,
         n_11, n_10, n_7, n_4, n_3, n_0, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65;
  assign n[498] = n_498;
  assign n[495] = n_495;
  assign n[494] = n_494;
  assign n[491] = n_491;
  assign n[488] = n_488;
  assign n[487] = n_487;
  assign n[486] = n_486;
  assign n[483] = n_483;
  assign n[480] = n_480;
  assign n[479] = n_479;
  assign n[476] = n_476;
  assign n[473] = n_473;
  assign n[472] = n_472;
  assign n[471] = n_471;
  assign n[470] = n_470;
  assign n[467] = n_467;
  assign n[464] = n_464;
  assign n[463] = n_463;
  assign n[460] = n_460;
  assign n[457] = n_457;
  assign n[456] = n_456;
  assign n[455] = n_455;
  assign n[452] = n_452;
  assign n[449] = n_449;
  assign n[448] = n_448;
  assign n[445] = n_445;
  assign n[442] = n_442;
  assign n[441] = n_441;
  assign n[440] = n_440;
  assign n[439] = n_439;
  assign n[438] = n_438;
  assign n[435] = n_435;
  assign n[432] = n_432;
  assign n[431] = n_431;
  assign n[428] = n_428;
  assign n[425] = n_425;
  assign n[424] = n_424;
  assign n[423] = n_423;
  assign n[420] = n_420;
  assign n[417] = n_417;
  assign n[416] = n_416;
  assign n[413] = n_413;
  assign n[410] = n_410;
  assign n[409] = n_409;
  assign n[408] = n_408;
  assign n[407] = n_407;
  assign n[404] = n_404;
  assign n[401] = n_401;
  assign n[400] = n_400;
  assign n[397] = n_397;
  assign n[394] = n_394;
  assign n[393] = n_393;
  assign n[392] = n_392;
  assign n[389] = n_389;
  assign n[386] = n_386;
  assign n[385] = n_385;
  assign n[382] = n_382;
  assign n[379] = n_379;
  assign n[378] = n_378;
  assign n[377] = n_377;
  assign n[376] = n_376;
  assign n[375] = n_375;
  assign n[374] = n_374;
  assign n[371] = n_371;
  assign n[368] = n_368;
  assign n[367] = n_367;
  assign n[364] = n_364;
  assign n[361] = n_361;
  assign n[360] = n_360;
  assign n[359] = n_359;
  assign n[356] = n_356;
  assign n[353] = n_353;
  assign n[352] = n_352;
  assign n[349] = n_349;
  assign n[346] = n_346;
  assign n[345] = n_345;
  assign n[344] = n_344;
  assign n[343] = n_343;
  assign n[340] = n_340;
  assign n[337] = n_337;
  assign n[336] = n_336;
  assign n[333] = n_333;
  assign n[330] = n_330;
  assign n[329] = n_329;
  assign n[328] = n_328;
  assign n[325] = n_325;
  assign n[322] = n_322;
  assign n[321] = n_321;
  assign n[318] = n_318;
  assign n[315] = n_315;
  assign n[314] = n_314;
  assign n[313] = n_313;
  assign n[312] = n_312;
  assign n[311] = n_311;
  assign n[308] = n_308;
  assign n[305] = n_305;
  assign n[304] = n_304;
  assign n[301] = n_301;
  assign n[298] = n_298;
  assign n[297] = n_297;
  assign n[296] = n_296;
  assign n[293] = n_293;
  assign n[290] = n_290;
  assign n[289] = n_289;
  assign n[286] = n_286;
  assign n[283] = n_283;
  assign n[282] = n_282;
  assign n[281] = n_281;
  assign n[280] = n_280;
  assign n[277] = n_277;
  assign n[274] = n_274;
  assign n[273] = n_273;
  assign n[270] = n_270;
  assign n[267] = n_267;
  assign n[266] = n_266;
  assign n[265] = n_265;
  assign n[262] = n_262;
  assign n[259] = n_259;
  assign n[258] = n_258;
  assign n[255] = n_255;
  assign n[243] = n_243;
  assign n[240] = n_240;
  assign n[239] = n_239;
  assign n[236] = n_236;
  assign n[233] = n_233;
  assign n[232] = n_232;
  assign n[231] = n_231;
  assign n[228] = n_228;
  assign n[225] = n_225;
  assign n[224] = n_224;
  assign n[221] = n_221;
  assign n[218] = n_218;
  assign n[217] = n_217;
  assign n[216] = n_216;
  assign n[215] = n_215;
  assign n[212] = n_212;
  assign n[209] = n_209;
  assign n[208] = n_208;
  assign n[205] = n_205;
  assign n[202] = n_202;
  assign n[201] = n_201;
  assign n[200] = n_200;
  assign n[197] = n_197;
  assign n[194] = n_194;
  assign n[193] = n_193;
  assign n[190] = n_190;
  assign n[187] = n_187;
  assign n[186] = n_186;
  assign n[185] = n_185;
  assign n[184] = n_184;
  assign n[183] = n_183;
  assign n[180] = n_180;
  assign n[177] = n_177;
  assign n[176] = n_176;
  assign n[173] = n_173;
  assign n[170] = n_170;
  assign n[169] = n_169;
  assign n[168] = n_168;
  assign n[165] = n_165;
  assign n[162] = n_162;
  assign n[161] = n_161;
  assign n[158] = n_158;
  assign n[155] = n_155;
  assign n[154] = n_154;
  assign n[153] = n_153;
  assign n[152] = n_152;
  assign n[149] = n_149;
  assign n[146] = n_146;
  assign n[145] = n_145;
  assign n[142] = n_142;
  assign n[139] = n_139;
  assign n[138] = n_138;
  assign n[137] = n_137;
  assign n[134] = n_134;
  assign n[131] = n_131;
  assign n[130] = n_130;
  assign n[127] = n_127;
  assign n[124] = n_124;
  assign n[123] = n_123;
  assign n[122] = n_122;
  assign n[121] = n_121;
  assign n[120] = n_120;
  assign n[119] = n_119;
  assign n[116] = n_116;
  assign n[113] = n_113;
  assign n[112] = n_112;
  assign n[109] = n_109;
  assign n[106] = n_106;
  assign n[105] = n_105;
  assign n[104] = n_104;
  assign n[101] = n_101;
  assign n[98] = n_98;
  assign n[97] = n_97;
  assign n[94] = n_94;
  assign n[91] = n_91;
  assign n[90] = n_90;
  assign n[89] = n_89;
  assign n[88] = n_88;
  assign n[85] = n_85;
  assign n[82] = n_82;
  assign n[81] = n_81;
  assign n[78] = n_78;
  assign n[75] = n_75;
  assign n[74] = n_74;
  assign n[73] = n_73;
  assign n[70] = n_70;
  assign n[67] = n_67;
  assign n[66] = n_66;
  assign n[63] = n_63;
  assign n[60] = n_60;
  assign n[59] = n_59;
  assign n[58] = n_58;
  assign n[57] = n_57;
  assign n[56] = n_56;
  assign n[53] = n_53;
  assign n[50] = n_50;
  assign n[49] = n_49;
  assign n[46] = n_46;
  assign n[43] = n_43;
  assign n[42] = n_42;
  assign n[41] = n_41;
  assign n[38] = n_38;
  assign n[35] = n_35;
  assign n[34] = n_34;
  assign n[31] = n_31;
  assign n[28] = n_28;
  assign n[27] = n_27;
  assign n[26] = n_26;
  assign n[25] = n_25;
  assign n[22] = n_22;
  assign n[19] = n_19;
  assign n[18] = n_18;
  assign n[15] = n_15;
  assign n[12] = n_12;
  assign n[11] = n_11;
  assign n[10] = n_10;
  assign n[7] = n_7;
  assign n[4] = n_4;
  assign n[3] = n_3;
  assign n[0] = n_0;

  NR2D0 U2 ( .A1(n1), .A2(n2), .ZN(n_498) );
  NR2D0 U3 ( .A1(n2), .A2(n3), .ZN(n_495) );
  NR2D0 U4 ( .A1(n2), .A2(n4), .ZN(n_494) );
  NR2D0 U5 ( .A1(n2), .A2(n5), .ZN(n_491) );
  NR2D0 U6 ( .A1(n2), .A2(n6), .ZN(n_488) );
  NR2D0 U7 ( .A1(n2), .A2(n7), .ZN(n_487) );
  NR2D0 U8 ( .A1(n2), .A2(n8), .ZN(n_486) );
  NR2D0 U9 ( .A1(n2), .A2(n9), .ZN(n_483) );
  NR2D0 U10 ( .A1(n2), .A2(n10), .ZN(n_480) );
  NR2D0 U11 ( .A1(n2), .A2(n11), .ZN(n_479) );
  NR2D0 U12 ( .A1(n2), .A2(n12), .ZN(n_476) );
  NR2D0 U13 ( .A1(n2), .A2(n13), .ZN(n_473) );
  NR2D0 U14 ( .A1(n2), .A2(n14), .ZN(n_472) );
  NR2D0 U15 ( .A1(n2), .A2(n15), .ZN(n_471) );
  NR2D0 U16 ( .A1(n2), .A2(n16), .ZN(n_470) );
  NR2D0 U17 ( .A1(n2), .A2(n17), .ZN(n_467) );
  NR2D0 U18 ( .A1(n2), .A2(n18), .ZN(n_464) );
  NR2D0 U19 ( .A1(n2), .A2(n19), .ZN(n_463) );
  NR2D0 U20 ( .A1(n2), .A2(n20), .ZN(n_460) );
  NR2D0 U21 ( .A1(n2), .A2(n21), .ZN(n_457) );
  NR2D0 U22 ( .A1(n2), .A2(n22), .ZN(n_456) );
  NR2D0 U23 ( .A1(n2), .A2(n23), .ZN(n_455) );
  NR2D0 U24 ( .A1(n2), .A2(n24), .ZN(n_452) );
  NR2D0 U25 ( .A1(n2), .A2(n25), .ZN(n_449) );
  NR2D0 U26 ( .A1(n2), .A2(n26), .ZN(n_448) );
  NR2D0 U27 ( .A1(n2), .A2(n27), .ZN(n_445) );
  NR2D0 U28 ( .A1(n2), .A2(n28), .ZN(n_442) );
  NR2D0 U29 ( .A1(n2), .A2(n29), .ZN(n_441) );
  NR2D0 U30 ( .A1(n2), .A2(n30), .ZN(n_440) );
  NR2D0 U31 ( .A1(n2), .A2(n31), .ZN(n_439) );
  NR2D0 U32 ( .A1(n2), .A2(n32), .ZN(n_438) );
  NR2D0 U33 ( .A1(n2), .A2(n33), .ZN(n_435) );
  NR2D0 U34 ( .A1(n2), .A2(n34), .ZN(n_432) );
  NR2D0 U35 ( .A1(n2), .A2(n35), .ZN(n_431) );
  NR2D0 U36 ( .A1(n2), .A2(n36), .ZN(n_428) );
  NR2D0 U37 ( .A1(n2), .A2(n37), .ZN(n_425) );
  NR2D0 U38 ( .A1(n2), .A2(n38), .ZN(n_424) );
  NR2D0 U39 ( .A1(n2), .A2(n39), .ZN(n_423) );
  NR2D0 U40 ( .A1(n2), .A2(n40), .ZN(n_420) );
  NR2D0 U41 ( .A1(n2), .A2(n41), .ZN(n_417) );
  NR2D0 U42 ( .A1(n2), .A2(n42), .ZN(n_416) );
  NR2D0 U43 ( .A1(n2), .A2(n43), .ZN(n_413) );
  NR2D0 U44 ( .A1(n2), .A2(n44), .ZN(n_410) );
  NR2D0 U45 ( .A1(n2), .A2(n45), .ZN(n_409) );
  NR2D0 U46 ( .A1(n2), .A2(n46), .ZN(n_408) );
  NR2D0 U47 ( .A1(n2), .A2(n47), .ZN(n_407) );
  NR2D0 U48 ( .A1(n2), .A2(n48), .ZN(n_404) );
  NR2D0 U49 ( .A1(n2), .A2(n49), .ZN(n_401) );
  NR2D0 U50 ( .A1(n2), .A2(n50), .ZN(n_400) );
  NR2D0 U51 ( .A1(n2), .A2(n51), .ZN(n_397) );
  NR2D0 U52 ( .A1(n2), .A2(n52), .ZN(n_394) );
  NR2D0 U53 ( .A1(n2), .A2(n53), .ZN(n_393) );
  NR2D0 U54 ( .A1(n2), .A2(n54), .ZN(n_392) );
  NR2D0 U55 ( .A1(n2), .A2(n55), .ZN(n_389) );
  NR2D0 U56 ( .A1(n2), .A2(n56), .ZN(n_386) );
  NR2D0 U57 ( .A1(n2), .A2(n57), .ZN(n_385) );
  NR2D0 U58 ( .A1(n2), .A2(n58), .ZN(n_382) );
  NR2D0 U59 ( .A1(n2), .A2(n59), .ZN(n_379) );
  NR2D0 U60 ( .A1(n2), .A2(n60), .ZN(n_378) );
  NR2D0 U61 ( .A1(n2), .A2(n61), .ZN(n_377) );
  NR2D0 U62 ( .A1(n2), .A2(n62), .ZN(n_376) );
  NR2D0 U63 ( .A1(n2), .A2(n63), .ZN(n_375) );
  NR2D0 U64 ( .A1(n2), .A2(n64), .ZN(n_374) );
  NR2D0 U65 ( .A1(n1), .A2(n65), .ZN(n_371) );
  NR2D0 U66 ( .A1(n3), .A2(n65), .ZN(n_368) );
  NR2D0 U67 ( .A1(n4), .A2(n65), .ZN(n_367) );
  NR2D0 U68 ( .A1(n5), .A2(n65), .ZN(n_364) );
  NR2D0 U69 ( .A1(n6), .A2(n65), .ZN(n_361) );
  NR2D0 U70 ( .A1(n7), .A2(n65), .ZN(n_360) );
  NR2D0 U71 ( .A1(n8), .A2(n65), .ZN(n_359) );
  NR2D0 U72 ( .A1(n9), .A2(n65), .ZN(n_356) );
  NR2D0 U73 ( .A1(n10), .A2(n65), .ZN(n_353) );
  NR2D0 U74 ( .A1(n11), .A2(n65), .ZN(n_352) );
  NR2D0 U75 ( .A1(n12), .A2(n65), .ZN(n_349) );
  NR2D0 U76 ( .A1(n13), .A2(n65), .ZN(n_346) );
  NR2D0 U77 ( .A1(n14), .A2(n65), .ZN(n_345) );
  NR2D0 U78 ( .A1(n15), .A2(n65), .ZN(n_344) );
  NR2D0 U79 ( .A1(n16), .A2(n65), .ZN(n_343) );
  NR2D0 U80 ( .A1(n17), .A2(n65), .ZN(n_340) );
  NR2D0 U81 ( .A1(n18), .A2(n65), .ZN(n_337) );
  NR2D0 U82 ( .A1(n19), .A2(n65), .ZN(n_336) );
  NR2D0 U83 ( .A1(n20), .A2(n65), .ZN(n_333) );
  NR2D0 U84 ( .A1(n21), .A2(n65), .ZN(n_330) );
  NR2D0 U85 ( .A1(n22), .A2(n65), .ZN(n_329) );
  NR2D0 U86 ( .A1(n23), .A2(n65), .ZN(n_328) );
  NR2D0 U87 ( .A1(n24), .A2(n65), .ZN(n_325) );
  NR2D0 U88 ( .A1(n25), .A2(n65), .ZN(n_322) );
  NR2D0 U89 ( .A1(n26), .A2(n65), .ZN(n_321) );
  NR2D0 U90 ( .A1(n27), .A2(n65), .ZN(n_318) );
  NR2D0 U91 ( .A1(n28), .A2(n65), .ZN(n_315) );
  NR2D0 U92 ( .A1(n29), .A2(n65), .ZN(n_314) );
  NR2D0 U93 ( .A1(n30), .A2(n65), .ZN(n_313) );
  NR2D0 U94 ( .A1(n31), .A2(n65), .ZN(n_312) );
  NR2D0 U95 ( .A1(n32), .A2(n65), .ZN(n_311) );
  NR2D0 U96 ( .A1(n33), .A2(n65), .ZN(n_308) );
  NR2D0 U97 ( .A1(n34), .A2(n65), .ZN(n_305) );
  NR2D0 U98 ( .A1(n35), .A2(n65), .ZN(n_304) );
  NR2D0 U99 ( .A1(n36), .A2(n65), .ZN(n_301) );
  NR2D0 U100 ( .A1(n37), .A2(n65), .ZN(n_298) );
  NR2D0 U101 ( .A1(n38), .A2(n65), .ZN(n_297) );
  NR2D0 U102 ( .A1(n39), .A2(n65), .ZN(n_296) );
  NR2D0 U103 ( .A1(n40), .A2(n65), .ZN(n_293) );
  NR2D0 U104 ( .A1(n41), .A2(n65), .ZN(n_290) );
  NR2D0 U105 ( .A1(n42), .A2(n65), .ZN(n_289) );
  NR2D0 U106 ( .A1(n43), .A2(n65), .ZN(n_286) );
  NR2D0 U107 ( .A1(n44), .A2(n65), .ZN(n_283) );
  NR2D0 U108 ( .A1(n45), .A2(n65), .ZN(n_282) );
  NR2D0 U109 ( .A1(n46), .A2(n65), .ZN(n_281) );
  NR2D0 U110 ( .A1(n47), .A2(n65), .ZN(n_280) );
  NR2D0 U111 ( .A1(n48), .A2(n65), .ZN(n_277) );
  NR2D0 U112 ( .A1(n49), .A2(n65), .ZN(n_274) );
  NR2D0 U113 ( .A1(n50), .A2(n65), .ZN(n_273) );
  NR2D0 U114 ( .A1(n51), .A2(n65), .ZN(n_270) );
  NR2D0 U115 ( .A1(n52), .A2(n65), .ZN(n_267) );
  NR2D0 U116 ( .A1(n53), .A2(n65), .ZN(n_266) );
  NR2D0 U117 ( .A1(n54), .A2(n65), .ZN(n_265) );
  NR2D0 U118 ( .A1(n55), .A2(n65), .ZN(n_262) );
  NR2D0 U119 ( .A1(n56), .A2(n65), .ZN(n_259) );
  NR2D0 U120 ( .A1(n57), .A2(n65), .ZN(n_258) );
  NR2D0 U121 ( .A1(n58), .A2(n65), .ZN(n_255) );
  INVD0 U122 ( .I(n1), .ZN(n_243) );
  ND2D0 U123 ( .A1(b[5]), .A2(n_116), .ZN(n1) );
  INVD0 U124 ( .I(n3), .ZN(n_240) );
  ND2D0 U125 ( .A1(n_113), .A2(b[5]), .ZN(n3) );
  INVD0 U126 ( .I(n4), .ZN(n_239) );
  ND2D0 U127 ( .A1(n_112), .A2(b[5]), .ZN(n4) );
  INVD0 U128 ( .I(n5), .ZN(n_236) );
  ND2D0 U129 ( .A1(n_109), .A2(b[5]), .ZN(n5) );
  INVD0 U130 ( .I(n6), .ZN(n_233) );
  ND2D0 U131 ( .A1(n_106), .A2(b[5]), .ZN(n6) );
  INVD0 U132 ( .I(n7), .ZN(n_232) );
  ND2D0 U133 ( .A1(n_105), .A2(b[5]), .ZN(n7) );
  INVD0 U134 ( .I(n8), .ZN(n_231) );
  ND2D0 U135 ( .A1(n_104), .A2(b[5]), .ZN(n8) );
  INVD0 U136 ( .I(n9), .ZN(n_228) );
  ND2D0 U137 ( .A1(n_101), .A2(b[5]), .ZN(n9) );
  INVD0 U138 ( .I(n10), .ZN(n_225) );
  ND2D0 U139 ( .A1(n_98), .A2(b[5]), .ZN(n10) );
  INVD0 U140 ( .I(n11), .ZN(n_224) );
  ND2D0 U141 ( .A1(n_97), .A2(b[5]), .ZN(n11) );
  INVD0 U142 ( .I(n12), .ZN(n_221) );
  ND2D0 U143 ( .A1(n_94), .A2(b[5]), .ZN(n12) );
  INVD0 U144 ( .I(n13), .ZN(n_218) );
  ND2D0 U145 ( .A1(n_91), .A2(b[5]), .ZN(n13) );
  INVD0 U146 ( .I(n14), .ZN(n_217) );
  ND2D0 U147 ( .A1(n_90), .A2(b[5]), .ZN(n14) );
  INVD0 U148 ( .I(n15), .ZN(n_216) );
  ND2D0 U149 ( .A1(n_89), .A2(b[5]), .ZN(n15) );
  INVD0 U150 ( .I(n16), .ZN(n_215) );
  ND2D0 U151 ( .A1(n_88), .A2(b[5]), .ZN(n16) );
  INVD0 U152 ( .I(n17), .ZN(n_212) );
  ND2D0 U153 ( .A1(n_85), .A2(b[5]), .ZN(n17) );
  INVD0 U154 ( .I(n18), .ZN(n_209) );
  ND2D0 U155 ( .A1(n_82), .A2(b[5]), .ZN(n18) );
  INVD0 U156 ( .I(n19), .ZN(n_208) );
  ND2D0 U157 ( .A1(n_81), .A2(b[5]), .ZN(n19) );
  INVD0 U158 ( .I(n20), .ZN(n_205) );
  ND2D0 U159 ( .A1(n_78), .A2(b[5]), .ZN(n20) );
  INVD0 U160 ( .I(n21), .ZN(n_202) );
  ND2D0 U161 ( .A1(n_75), .A2(b[5]), .ZN(n21) );
  INVD0 U162 ( .I(n22), .ZN(n_201) );
  ND2D0 U163 ( .A1(n_74), .A2(b[5]), .ZN(n22) );
  INVD0 U164 ( .I(n23), .ZN(n_200) );
  ND2D0 U165 ( .A1(n_73), .A2(b[5]), .ZN(n23) );
  INVD0 U166 ( .I(n24), .ZN(n_197) );
  ND2D0 U167 ( .A1(n_70), .A2(b[5]), .ZN(n24) );
  INVD0 U168 ( .I(n25), .ZN(n_194) );
  ND2D0 U169 ( .A1(n_67), .A2(b[5]), .ZN(n25) );
  INVD0 U170 ( .I(n26), .ZN(n_193) );
  ND2D0 U171 ( .A1(n_66), .A2(b[5]), .ZN(n26) );
  INVD0 U172 ( .I(n27), .ZN(n_190) );
  ND2D0 U173 ( .A1(n_63), .A2(b[5]), .ZN(n27) );
  INVD0 U174 ( .I(n28), .ZN(n_187) );
  ND2D0 U175 ( .A1(n_60), .A2(b[5]), .ZN(n28) );
  INVD0 U176 ( .I(n29), .ZN(n_186) );
  ND2D0 U177 ( .A1(n_59), .A2(b[5]), .ZN(n29) );
  INVD0 U178 ( .I(n30), .ZN(n_185) );
  ND2D0 U179 ( .A1(n_58), .A2(b[5]), .ZN(n30) );
  INVD0 U180 ( .I(n31), .ZN(n_184) );
  ND2D0 U181 ( .A1(n_57), .A2(b[5]), .ZN(n31) );
  INVD0 U182 ( .I(n32), .ZN(n_183) );
  ND2D0 U183 ( .A1(n_56), .A2(b[5]), .ZN(n32) );
  INVD0 U184 ( .I(n33), .ZN(n_180) );
  ND2D0 U185 ( .A1(a[5]), .A2(n_116), .ZN(n33) );
  INVD0 U186 ( .I(n34), .ZN(n_177) );
  ND2D0 U187 ( .A1(a[5]), .A2(n_113), .ZN(n34) );
  INVD0 U188 ( .I(n35), .ZN(n_176) );
  ND2D0 U189 ( .A1(a[5]), .A2(n_112), .ZN(n35) );
  INVD0 U190 ( .I(n36), .ZN(n_173) );
  ND2D0 U191 ( .A1(a[5]), .A2(n_109), .ZN(n36) );
  INVD0 U192 ( .I(n37), .ZN(n_170) );
  ND2D0 U193 ( .A1(a[5]), .A2(n_106), .ZN(n37) );
  INVD0 U194 ( .I(n38), .ZN(n_169) );
  ND2D0 U195 ( .A1(a[5]), .A2(n_105), .ZN(n38) );
  INVD0 U196 ( .I(n39), .ZN(n_168) );
  ND2D0 U197 ( .A1(a[5]), .A2(n_104), .ZN(n39) );
  INVD0 U198 ( .I(n40), .ZN(n_165) );
  ND2D0 U199 ( .A1(a[5]), .A2(n_101), .ZN(n40) );
  INVD0 U200 ( .I(n41), .ZN(n_162) );
  ND2D0 U201 ( .A1(a[5]), .A2(n_98), .ZN(n41) );
  AN2D0 U202 ( .A1(b[4]), .A2(n_35), .Z(n_98) );
  INVD0 U203 ( .I(n42), .ZN(n_161) );
  ND2D0 U204 ( .A1(a[5]), .A2(n_97), .ZN(n42) );
  AN2D0 U205 ( .A1(n_34), .A2(b[4]), .Z(n_97) );
  INVD0 U206 ( .I(n43), .ZN(n_158) );
  ND2D0 U207 ( .A1(a[5]), .A2(n_94), .ZN(n43) );
  AN2D0 U208 ( .A1(n_31), .A2(b[4]), .Z(n_94) );
  INVD0 U209 ( .I(n44), .ZN(n_155) );
  ND2D0 U210 ( .A1(a[5]), .A2(n_91), .ZN(n44) );
  AN2D0 U211 ( .A1(n_28), .A2(b[4]), .Z(n_91) );
  INVD0 U212 ( .I(n45), .ZN(n_154) );
  ND2D0 U213 ( .A1(a[5]), .A2(n_90), .ZN(n45) );
  AN2D0 U214 ( .A1(n_27), .A2(b[4]), .Z(n_90) );
  INVD0 U215 ( .I(n46), .ZN(n_153) );
  ND2D0 U216 ( .A1(a[5]), .A2(n_89), .ZN(n46) );
  AN2D0 U217 ( .A1(n_26), .A2(b[4]), .Z(n_89) );
  INVD0 U218 ( .I(n47), .ZN(n_152) );
  ND2D0 U219 ( .A1(a[5]), .A2(n_88), .ZN(n47) );
  AN2D0 U220 ( .A1(n_25), .A2(b[4]), .Z(n_88) );
  INVD0 U221 ( .I(n48), .ZN(n_149) );
  ND2D0 U222 ( .A1(a[5]), .A2(n_85), .ZN(n48) );
  AN2D0 U223 ( .A1(a[4]), .A2(n_53), .Z(n_85) );
  INVD0 U224 ( .I(n49), .ZN(n_146) );
  ND2D0 U225 ( .A1(a[5]), .A2(n_82), .ZN(n49) );
  AN2D0 U226 ( .A1(n_50), .A2(a[4]), .Z(n_82) );
  INVD0 U227 ( .I(n50), .ZN(n_145) );
  ND2D0 U228 ( .A1(a[5]), .A2(n_81), .ZN(n50) );
  AN2D0 U229 ( .A1(n_49), .A2(a[4]), .Z(n_81) );
  INVD0 U230 ( .I(n51), .ZN(n_142) );
  ND2D0 U231 ( .A1(a[5]), .A2(n_78), .ZN(n51) );
  AN2D0 U232 ( .A1(n_46), .A2(a[4]), .Z(n_78) );
  INVD0 U233 ( .I(n52), .ZN(n_139) );
  ND2D0 U234 ( .A1(a[5]), .A2(n_75), .ZN(n52) );
  AN2D0 U235 ( .A1(n_43), .A2(a[4]), .Z(n_75) );
  INVD0 U236 ( .I(n53), .ZN(n_138) );
  ND2D0 U237 ( .A1(a[5]), .A2(n_74), .ZN(n53) );
  AN2D0 U238 ( .A1(n_42), .A2(a[4]), .Z(n_74) );
  INVD0 U239 ( .I(n54), .ZN(n_137) );
  ND2D0 U240 ( .A1(a[5]), .A2(n_73), .ZN(n54) );
  AN2D0 U241 ( .A1(n_41), .A2(a[4]), .Z(n_73) );
  INVD0 U242 ( .I(n55), .ZN(n_134) );
  ND2D0 U243 ( .A1(a[5]), .A2(n_70), .ZN(n55) );
  AN2D0 U244 ( .A1(n_38), .A2(a[4]), .Z(n_70) );
  INVD0 U245 ( .I(n56), .ZN(n_131) );
  ND2D0 U246 ( .A1(a[5]), .A2(n_67), .ZN(n56) );
  AN2D0 U247 ( .A1(a[4]), .A2(n_35), .Z(n_67) );
  AN2D0 U248 ( .A1(a[3]), .A2(n_19), .Z(n_35) );
  INVD0 U249 ( .I(n57), .ZN(n_130) );
  ND2D0 U250 ( .A1(a[5]), .A2(n_66), .ZN(n57) );
  AN2D0 U251 ( .A1(a[4]), .A2(n_34), .Z(n_66) );
  AN2D0 U252 ( .A1(n_18), .A2(a[3]), .Z(n_34) );
  INVD0 U253 ( .I(n58), .ZN(n_127) );
  ND2D0 U254 ( .A1(a[5]), .A2(n_63), .ZN(n58) );
  AN2D0 U255 ( .A1(a[4]), .A2(n_31), .Z(n_63) );
  AN2D0 U256 ( .A1(n_15), .A2(a[3]), .Z(n_31) );
  INVD0 U257 ( .I(n59), .ZN(n_124) );
  INVD0 U258 ( .I(n60), .ZN(n_123) );
  INVD0 U259 ( .I(n61), .ZN(n_122) );
  INVD0 U260 ( .I(n62), .ZN(n_121) );
  INVD0 U261 ( .I(n63), .ZN(n_120) );
  INVD0 U262 ( .I(n64), .ZN(n_119) );
  AN2D0 U263 ( .A1(n_53), .A2(b[4]), .Z(n_116) );
  AN2D0 U264 ( .A1(n_22), .A2(b[3]), .Z(n_53) );
  AN2D0 U265 ( .A1(n_50), .A2(b[4]), .Z(n_113) );
  AN2D0 U266 ( .A1(b[3]), .A2(n_19), .Z(n_50) );
  AN2D0 U267 ( .A1(b[2]), .A2(n_4), .Z(n_19) );
  AN2D0 U268 ( .A1(n_49), .A2(b[4]), .Z(n_112) );
  AN2D0 U269 ( .A1(b[3]), .A2(n_18), .Z(n_49) );
  AN2D0 U270 ( .A1(n_3), .A2(b[2]), .Z(n_18) );
  AN2D0 U271 ( .A1(n_46), .A2(b[4]), .Z(n_109) );
  AN2D0 U272 ( .A1(b[3]), .A2(n_15), .Z(n_46) );
  AN2D0 U273 ( .A1(a[2]), .A2(n_7), .Z(n_15) );
  AN2D0 U274 ( .A1(n_43), .A2(b[4]), .Z(n_106) );
  AN2D0 U275 ( .A1(b[3]), .A2(n_12), .Z(n_43) );
  AN2D0 U276 ( .A1(n_42), .A2(b[4]), .Z(n_105) );
  AN2D0 U277 ( .A1(b[3]), .A2(n_11), .Z(n_42) );
  AN2D0 U278 ( .A1(n_41), .A2(b[4]), .Z(n_104) );
  AN2D0 U279 ( .A1(b[3]), .A2(n_10), .Z(n_41) );
  AN2D0 U280 ( .A1(n_38), .A2(b[4]), .Z(n_101) );
  AN2D0 U281 ( .A1(n_22), .A2(a[3]), .Z(n_38) );
  AN2D0 U282 ( .A1(n_7), .A2(b[2]), .Z(n_22) );
  AN2D0 U283 ( .A1(b[1]), .A2(n_0), .Z(n_7) );
  NR2D0 U284 ( .A1(n59), .A2(n65), .ZN(n[252]) );
  ND2D0 U285 ( .A1(a[5]), .A2(n_60), .ZN(n59) );
  AN2D0 U286 ( .A1(a[4]), .A2(n_28), .Z(n_60) );
  AN2D0 U287 ( .A1(n_12), .A2(a[3]), .Z(n_28) );
  AN2D0 U288 ( .A1(a[2]), .A2(n_4), .Z(n_12) );
  AN2D0 U289 ( .A1(a[1]), .A2(n_0), .Z(n_4) );
  AN2D0 U290 ( .A1(b[0]), .A2(a[0]), .Z(n_0) );
  NR2D0 U291 ( .A1(n60), .A2(n65), .ZN(n[251]) );
  ND2D0 U292 ( .A1(a[5]), .A2(n_59), .ZN(n60) );
  AN2D0 U293 ( .A1(a[4]), .A2(n_27), .Z(n_59) );
  AN2D0 U294 ( .A1(n_11), .A2(a[3]), .Z(n_27) );
  AN2D0 U295 ( .A1(a[2]), .A2(n_3), .Z(n_11) );
  AN2D0 U296 ( .A1(b[1]), .A2(a[1]), .Z(n_3) );
  NR2D0 U297 ( .A1(n61), .A2(n65), .ZN(n[250]) );
  ND2D0 U298 ( .A1(a[5]), .A2(n_58), .ZN(n61) );
  AN2D0 U299 ( .A1(a[4]), .A2(n_26), .Z(n_58) );
  AN2D0 U300 ( .A1(n_10), .A2(a[3]), .Z(n_26) );
  AN2D0 U301 ( .A1(a[2]), .A2(b[2]), .Z(n_10) );
  NR2D0 U302 ( .A1(n62), .A2(n65), .ZN(n[249]) );
  ND2D0 U303 ( .A1(a[5]), .A2(n_57), .ZN(n62) );
  AN2D0 U304 ( .A1(a[4]), .A2(n_25), .Z(n_57) );
  AN2D0 U305 ( .A1(b[3]), .A2(a[3]), .Z(n_25) );
  NR2D0 U306 ( .A1(n63), .A2(n65), .ZN(n[248]) );
  ND2D0 U307 ( .A1(a[5]), .A2(n_56), .ZN(n63) );
  AN2D0 U308 ( .A1(a[4]), .A2(b[4]), .Z(n_56) );
  NR2D0 U309 ( .A1(n64), .A2(n65), .ZN(n[247]) );
  ND2D0 U310 ( .A1(a[5]), .A2(b[5]), .ZN(n64) );
  NR2D0 U311 ( .A1(n2), .A2(n65), .ZN(n[246]) );
  INVD1 U312 ( .I(1'b1), .ZN(n[1]) );
  INVD1 U314 ( .I(1'b1), .ZN(n[2]) );
  INVD1 U316 ( .I(1'b1), .ZN(n[5]) );
  INVD1 U318 ( .I(1'b1), .ZN(n[6]) );
  INVD1 U320 ( .I(1'b1), .ZN(n[8]) );
  INVD1 U322 ( .I(1'b1), .ZN(n[9]) );
  INVD1 U324 ( .I(1'b1), .ZN(n[13]) );
  INVD1 U326 ( .I(1'b1), .ZN(n[14]) );
  INVD1 U328 ( .I(1'b1), .ZN(n[16]) );
  INVD1 U330 ( .I(1'b1), .ZN(n[17]) );
  INVD1 U332 ( .I(1'b1), .ZN(n[20]) );
  INVD1 U334 ( .I(1'b1), .ZN(n[21]) );
  INVD1 U336 ( .I(1'b1), .ZN(n[23]) );
  INVD1 U338 ( .I(1'b1), .ZN(n[24]) );
  INVD1 U340 ( .I(1'b1), .ZN(n[29]) );
  INVD1 U342 ( .I(1'b1), .ZN(n[30]) );
  INVD1 U344 ( .I(1'b1), .ZN(n[32]) );
  INVD1 U346 ( .I(1'b1), .ZN(n[33]) );
  INVD1 U348 ( .I(1'b1), .ZN(n[36]) );
  INVD1 U350 ( .I(1'b1), .ZN(n[37]) );
  INVD1 U352 ( .I(1'b1), .ZN(n[39]) );
  INVD1 U354 ( .I(1'b1), .ZN(n[40]) );
  INVD1 U356 ( .I(1'b1), .ZN(n[44]) );
  INVD1 U358 ( .I(1'b1), .ZN(n[45]) );
  INVD1 U360 ( .I(1'b1), .ZN(n[47]) );
  INVD1 U362 ( .I(1'b1), .ZN(n[48]) );
  INVD1 U364 ( .I(1'b1), .ZN(n[51]) );
  INVD1 U366 ( .I(1'b1), .ZN(n[52]) );
  INVD1 U368 ( .I(1'b1), .ZN(n[54]) );
  INVD1 U370 ( .I(1'b1), .ZN(n[55]) );
  INVD1 U372 ( .I(1'b1), .ZN(n[61]) );
  INVD1 U374 ( .I(1'b1), .ZN(n[62]) );
  INVD1 U376 ( .I(1'b1), .ZN(n[64]) );
  INVD1 U378 ( .I(1'b1), .ZN(n[65]) );
  INVD1 U380 ( .I(1'b1), .ZN(n[68]) );
  INVD1 U382 ( .I(1'b1), .ZN(n[69]) );
  INVD1 U384 ( .I(1'b1), .ZN(n[71]) );
  INVD1 U386 ( .I(1'b1), .ZN(n[72]) );
  INVD1 U388 ( .I(1'b1), .ZN(n[76]) );
  INVD1 U390 ( .I(1'b1), .ZN(n[77]) );
  INVD1 U392 ( .I(1'b1), .ZN(n[79]) );
  INVD1 U394 ( .I(1'b1), .ZN(n[80]) );
  INVD1 U396 ( .I(1'b1), .ZN(n[83]) );
  INVD1 U398 ( .I(1'b1), .ZN(n[84]) );
  INVD1 U400 ( .I(1'b1), .ZN(n[86]) );
  INVD1 U402 ( .I(1'b1), .ZN(n[87]) );
  INVD1 U404 ( .I(1'b1), .ZN(n[92]) );
  INVD1 U406 ( .I(1'b1), .ZN(n[93]) );
  INVD1 U408 ( .I(1'b1), .ZN(n[95]) );
  INVD1 U410 ( .I(1'b1), .ZN(n[96]) );
  INVD1 U412 ( .I(1'b1), .ZN(n[99]) );
  INVD1 U414 ( .I(1'b1), .ZN(n[100]) );
  INVD1 U416 ( .I(1'b1), .ZN(n[102]) );
  INVD1 U418 ( .I(1'b1), .ZN(n[103]) );
  INVD1 U420 ( .I(1'b1), .ZN(n[107]) );
  INVD1 U422 ( .I(1'b1), .ZN(n[108]) );
  INVD1 U424 ( .I(1'b1), .ZN(n[110]) );
  INVD1 U426 ( .I(1'b1), .ZN(n[111]) );
  INVD1 U428 ( .I(1'b1), .ZN(n[114]) );
  INVD1 U430 ( .I(1'b1), .ZN(n[115]) );
  INVD1 U432 ( .I(1'b1), .ZN(n[117]) );
  INVD1 U434 ( .I(1'b1), .ZN(n[118]) );
  INVD1 U436 ( .I(1'b1), .ZN(n[125]) );
  INVD1 U438 ( .I(1'b1), .ZN(n[126]) );
  INVD1 U440 ( .I(1'b1), .ZN(n[128]) );
  INVD1 U442 ( .I(1'b1), .ZN(n[129]) );
  INVD1 U444 ( .I(1'b1), .ZN(n[132]) );
  INVD1 U446 ( .I(1'b1), .ZN(n[133]) );
  INVD1 U448 ( .I(1'b1), .ZN(n[135]) );
  INVD1 U450 ( .I(1'b1), .ZN(n[136]) );
  INVD1 U452 ( .I(1'b1), .ZN(n[140]) );
  INVD1 U454 ( .I(1'b1), .ZN(n[141]) );
  INVD1 U456 ( .I(1'b1), .ZN(n[143]) );
  INVD1 U458 ( .I(1'b1), .ZN(n[144]) );
  INVD1 U460 ( .I(1'b1), .ZN(n[147]) );
  INVD1 U462 ( .I(1'b1), .ZN(n[148]) );
  INVD1 U464 ( .I(1'b1), .ZN(n[150]) );
  INVD1 U466 ( .I(1'b1), .ZN(n[151]) );
  INVD1 U468 ( .I(1'b1), .ZN(n[156]) );
  INVD1 U470 ( .I(1'b1), .ZN(n[157]) );
  INVD1 U472 ( .I(1'b1), .ZN(n[159]) );
  INVD1 U474 ( .I(1'b1), .ZN(n[160]) );
  INVD1 U476 ( .I(1'b1), .ZN(n[163]) );
  INVD1 U478 ( .I(1'b1), .ZN(n[164]) );
  INVD1 U480 ( .I(1'b1), .ZN(n[166]) );
  INVD1 U482 ( .I(1'b1), .ZN(n[167]) );
  INVD1 U484 ( .I(1'b1), .ZN(n[171]) );
  INVD1 U486 ( .I(1'b1), .ZN(n[172]) );
  INVD1 U488 ( .I(1'b1), .ZN(n[174]) );
  INVD1 U490 ( .I(1'b1), .ZN(n[175]) );
  INVD1 U492 ( .I(1'b1), .ZN(n[178]) );
  INVD1 U494 ( .I(1'b1), .ZN(n[179]) );
  INVD1 U496 ( .I(1'b1), .ZN(n[181]) );
  INVD1 U498 ( .I(1'b1), .ZN(n[182]) );
  INVD1 U500 ( .I(1'b1), .ZN(n[188]) );
  INVD1 U502 ( .I(1'b1), .ZN(n[189]) );
  INVD1 U504 ( .I(1'b1), .ZN(n[191]) );
  INVD1 U506 ( .I(1'b1), .ZN(n[192]) );
  INVD1 U508 ( .I(1'b1), .ZN(n[195]) );
  INVD1 U510 ( .I(1'b1), .ZN(n[196]) );
  INVD1 U512 ( .I(1'b1), .ZN(n[198]) );
  INVD1 U514 ( .I(1'b1), .ZN(n[199]) );
  INVD1 U516 ( .I(1'b1), .ZN(n[203]) );
  INVD1 U518 ( .I(1'b1), .ZN(n[204]) );
  INVD1 U520 ( .I(1'b1), .ZN(n[206]) );
  INVD1 U522 ( .I(1'b1), .ZN(n[207]) );
  INVD1 U524 ( .I(1'b1), .ZN(n[210]) );
  INVD1 U526 ( .I(1'b1), .ZN(n[211]) );
  INVD1 U528 ( .I(1'b1), .ZN(n[213]) );
  INVD1 U530 ( .I(1'b1), .ZN(n[214]) );
  INVD1 U532 ( .I(1'b1), .ZN(n[219]) );
  INVD1 U534 ( .I(1'b1), .ZN(n[220]) );
  INVD1 U536 ( .I(1'b1), .ZN(n[222]) );
  INVD1 U538 ( .I(1'b1), .ZN(n[223]) );
  INVD1 U540 ( .I(1'b1), .ZN(n[226]) );
  INVD1 U542 ( .I(1'b1), .ZN(n[227]) );
  INVD1 U544 ( .I(1'b1), .ZN(n[229]) );
  INVD1 U546 ( .I(1'b1), .ZN(n[230]) );
  INVD1 U548 ( .I(1'b1), .ZN(n[234]) );
  INVD1 U550 ( .I(1'b1), .ZN(n[235]) );
  INVD1 U552 ( .I(1'b1), .ZN(n[237]) );
  INVD1 U554 ( .I(1'b1), .ZN(n[238]) );
  INVD1 U556 ( .I(1'b1), .ZN(n[241]) );
  INVD1 U558 ( .I(1'b1), .ZN(n[242]) );
  INVD1 U560 ( .I(1'b1), .ZN(n[244]) );
  INVD1 U562 ( .I(1'b1), .ZN(n[245]) );
  INVD1 U564 ( .I(1'b1), .ZN(n[253]) );
  INVD1 U566 ( .I(1'b1), .ZN(n[254]) );
  INVD1 U568 ( .I(1'b1), .ZN(n[256]) );
  INVD1 U570 ( .I(1'b1), .ZN(n[257]) );
  INVD1 U572 ( .I(1'b1), .ZN(n[260]) );
  INVD1 U574 ( .I(1'b1), .ZN(n[261]) );
  INVD1 U576 ( .I(1'b1), .ZN(n[263]) );
  INVD1 U578 ( .I(1'b1), .ZN(n[264]) );
  INVD1 U580 ( .I(1'b1), .ZN(n[268]) );
  INVD1 U582 ( .I(1'b1), .ZN(n[269]) );
  INVD1 U584 ( .I(1'b1), .ZN(n[271]) );
  INVD1 U586 ( .I(1'b1), .ZN(n[272]) );
  INVD1 U588 ( .I(1'b1), .ZN(n[275]) );
  INVD1 U590 ( .I(1'b1), .ZN(n[276]) );
  INVD1 U592 ( .I(1'b1), .ZN(n[278]) );
  INVD1 U594 ( .I(1'b1), .ZN(n[279]) );
  INVD1 U596 ( .I(1'b1), .ZN(n[284]) );
  INVD1 U598 ( .I(1'b1), .ZN(n[285]) );
  INVD1 U600 ( .I(1'b1), .ZN(n[287]) );
  INVD1 U602 ( .I(1'b1), .ZN(n[288]) );
  INVD1 U604 ( .I(1'b1), .ZN(n[291]) );
  INVD1 U606 ( .I(1'b1), .ZN(n[292]) );
  INVD1 U608 ( .I(1'b1), .ZN(n[294]) );
  INVD1 U610 ( .I(1'b1), .ZN(n[295]) );
  INVD1 U612 ( .I(1'b1), .ZN(n[299]) );
  INVD1 U614 ( .I(1'b1), .ZN(n[300]) );
  INVD1 U616 ( .I(1'b1), .ZN(n[302]) );
  INVD1 U618 ( .I(1'b1), .ZN(n[303]) );
  INVD1 U620 ( .I(1'b1), .ZN(n[306]) );
  INVD1 U622 ( .I(1'b1), .ZN(n[307]) );
  INVD1 U624 ( .I(1'b1), .ZN(n[309]) );
  INVD1 U626 ( .I(1'b1), .ZN(n[310]) );
  INVD1 U628 ( .I(1'b1), .ZN(n[316]) );
  INVD1 U630 ( .I(1'b1), .ZN(n[317]) );
  INVD1 U632 ( .I(1'b1), .ZN(n[319]) );
  INVD1 U634 ( .I(1'b1), .ZN(n[320]) );
  INVD1 U636 ( .I(1'b1), .ZN(n[323]) );
  INVD1 U638 ( .I(1'b1), .ZN(n[324]) );
  INVD1 U640 ( .I(1'b1), .ZN(n[326]) );
  INVD1 U642 ( .I(1'b1), .ZN(n[327]) );
  INVD1 U644 ( .I(1'b1), .ZN(n[331]) );
  INVD1 U646 ( .I(1'b1), .ZN(n[332]) );
  INVD1 U648 ( .I(1'b1), .ZN(n[334]) );
  INVD1 U650 ( .I(1'b1), .ZN(n[335]) );
  INVD1 U652 ( .I(1'b1), .ZN(n[338]) );
  INVD1 U654 ( .I(1'b1), .ZN(n[339]) );
  INVD1 U656 ( .I(1'b1), .ZN(n[341]) );
  INVD1 U658 ( .I(1'b1), .ZN(n[342]) );
  INVD1 U660 ( .I(1'b1), .ZN(n[347]) );
  INVD1 U662 ( .I(1'b1), .ZN(n[348]) );
  INVD1 U664 ( .I(1'b1), .ZN(n[350]) );
  INVD1 U666 ( .I(1'b1), .ZN(n[351]) );
  INVD1 U668 ( .I(1'b1), .ZN(n[354]) );
  INVD1 U670 ( .I(1'b1), .ZN(n[355]) );
  INVD1 U672 ( .I(1'b1), .ZN(n[357]) );
  INVD1 U674 ( .I(1'b1), .ZN(n[358]) );
  INVD1 U676 ( .I(1'b1), .ZN(n[362]) );
  INVD1 U678 ( .I(1'b1), .ZN(n[363]) );
  INVD1 U680 ( .I(1'b1), .ZN(n[365]) );
  INVD1 U682 ( .I(1'b1), .ZN(n[366]) );
  INVD1 U684 ( .I(1'b1), .ZN(n[369]) );
  INVD1 U686 ( .I(1'b1), .ZN(n[370]) );
  INVD1 U688 ( .I(1'b1), .ZN(n[372]) );
  INVD1 U690 ( .I(1'b1), .ZN(n[373]) );
  INVD1 U692 ( .I(1'b1), .ZN(n[380]) );
  INVD1 U694 ( .I(1'b1), .ZN(n[381]) );
  INVD1 U696 ( .I(1'b1), .ZN(n[383]) );
  INVD1 U698 ( .I(1'b1), .ZN(n[384]) );
  INVD1 U700 ( .I(1'b1), .ZN(n[387]) );
  INVD1 U702 ( .I(1'b1), .ZN(n[388]) );
  INVD1 U704 ( .I(1'b1), .ZN(n[390]) );
  INVD1 U706 ( .I(1'b1), .ZN(n[391]) );
  INVD1 U708 ( .I(1'b1), .ZN(n[395]) );
  INVD1 U710 ( .I(1'b1), .ZN(n[396]) );
  INVD1 U712 ( .I(1'b1), .ZN(n[398]) );
  INVD1 U714 ( .I(1'b1), .ZN(n[399]) );
  INVD1 U716 ( .I(1'b1), .ZN(n[402]) );
  INVD1 U718 ( .I(1'b1), .ZN(n[403]) );
  INVD1 U720 ( .I(1'b1), .ZN(n[405]) );
  INVD1 U722 ( .I(1'b1), .ZN(n[406]) );
  INVD1 U724 ( .I(1'b1), .ZN(n[411]) );
  INVD1 U726 ( .I(1'b1), .ZN(n[412]) );
  INVD1 U728 ( .I(1'b1), .ZN(n[414]) );
  INVD1 U730 ( .I(1'b1), .ZN(n[415]) );
  INVD1 U732 ( .I(1'b1), .ZN(n[418]) );
  INVD1 U734 ( .I(1'b1), .ZN(n[419]) );
  INVD1 U736 ( .I(1'b1), .ZN(n[421]) );
  INVD1 U738 ( .I(1'b1), .ZN(n[422]) );
  INVD1 U740 ( .I(1'b1), .ZN(n[426]) );
  INVD1 U742 ( .I(1'b1), .ZN(n[427]) );
  INVD1 U744 ( .I(1'b1), .ZN(n[429]) );
  INVD1 U746 ( .I(1'b1), .ZN(n[430]) );
  INVD1 U748 ( .I(1'b1), .ZN(n[433]) );
  INVD1 U750 ( .I(1'b1), .ZN(n[434]) );
  INVD1 U752 ( .I(1'b1), .ZN(n[436]) );
  INVD1 U754 ( .I(1'b1), .ZN(n[437]) );
  INVD1 U756 ( .I(1'b1), .ZN(n[443]) );
  INVD1 U758 ( .I(1'b1), .ZN(n[444]) );
  INVD1 U760 ( .I(1'b1), .ZN(n[446]) );
  INVD1 U762 ( .I(1'b1), .ZN(n[447]) );
  INVD1 U764 ( .I(1'b1), .ZN(n[450]) );
  INVD1 U766 ( .I(1'b1), .ZN(n[451]) );
  INVD1 U768 ( .I(1'b1), .ZN(n[453]) );
  INVD1 U770 ( .I(1'b1), .ZN(n[454]) );
  INVD1 U772 ( .I(1'b1), .ZN(n[458]) );
  INVD1 U774 ( .I(1'b1), .ZN(n[459]) );
  INVD1 U776 ( .I(1'b1), .ZN(n[461]) );
  INVD1 U778 ( .I(1'b1), .ZN(n[462]) );
  INVD1 U780 ( .I(1'b1), .ZN(n[465]) );
  INVD1 U782 ( .I(1'b1), .ZN(n[466]) );
  INVD1 U784 ( .I(1'b1), .ZN(n[468]) );
  INVD1 U786 ( .I(1'b1), .ZN(n[469]) );
  INVD1 U788 ( .I(1'b1), .ZN(n[474]) );
  INVD1 U790 ( .I(1'b1), .ZN(n[475]) );
  INVD1 U792 ( .I(1'b1), .ZN(n[477]) );
  INVD1 U794 ( .I(1'b1), .ZN(n[478]) );
  INVD1 U796 ( .I(1'b1), .ZN(n[481]) );
  INVD1 U798 ( .I(1'b1), .ZN(n[482]) );
  INVD1 U800 ( .I(1'b1), .ZN(n[484]) );
  INVD1 U802 ( .I(1'b1), .ZN(n[485]) );
  INVD1 U804 ( .I(1'b1), .ZN(n[489]) );
  INVD1 U806 ( .I(1'b1), .ZN(n[490]) );
  INVD1 U808 ( .I(1'b1), .ZN(n[492]) );
  INVD1 U810 ( .I(1'b1), .ZN(n[493]) );
  INVD1 U812 ( .I(1'b1), .ZN(n[496]) );
  INVD1 U814 ( .I(1'b1), .ZN(n[497]) );
  INVD1 U816 ( .I(1'b1), .ZN(n[499]) );
  INVD1 U818 ( .I(1'b1), .ZN(n[500]) );
  INVD1 U820 ( .I(1'b1), .ZN(n[501]) );
  INVD1 U822 ( .I(a[6]), .ZN(n65) );
  INVD1 U823 ( .I(b[6]), .ZN(n2) );
endmodule


module gen_cla_decomposed ( a, b, s );
  input [7:0] a;
  input [7:0] b;
  output [7:0] s;

  wire   [501:0] n;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, 
        SYNOPSYS_UNCONNECTED__172, SYNOPSYS_UNCONNECTED__173, 
        SYNOPSYS_UNCONNECTED__174, SYNOPSYS_UNCONNECTED__175, 
        SYNOPSYS_UNCONNECTED__176, SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178, SYNOPSYS_UNCONNECTED__179, 
        SYNOPSYS_UNCONNECTED__180, SYNOPSYS_UNCONNECTED__181, 
        SYNOPSYS_UNCONNECTED__182, SYNOPSYS_UNCONNECTED__183, 
        SYNOPSYS_UNCONNECTED__184, SYNOPSYS_UNCONNECTED__185, 
        SYNOPSYS_UNCONNECTED__186, SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191, 
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        SYNOPSYS_UNCONNECTED__200, SYNOPSYS_UNCONNECTED__201, 
        SYNOPSYS_UNCONNECTED__202, SYNOPSYS_UNCONNECTED__203, 
        SYNOPSYS_UNCONNECTED__204, SYNOPSYS_UNCONNECTED__205, 
        SYNOPSYS_UNCONNECTED__206, SYNOPSYS_UNCONNECTED__207, 
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, 
        SYNOPSYS_UNCONNECTED__212, SYNOPSYS_UNCONNECTED__213, 
        SYNOPSYS_UNCONNECTED__214, SYNOPSYS_UNCONNECTED__215, 
        SYNOPSYS_UNCONNECTED__216, SYNOPSYS_UNCONNECTED__217, 
        SYNOPSYS_UNCONNECTED__218, SYNOPSYS_UNCONNECTED__219, 
        SYNOPSYS_UNCONNECTED__220, SYNOPSYS_UNCONNECTED__221, 
        SYNOPSYS_UNCONNECTED__222, SYNOPSYS_UNCONNECTED__223, 
        SYNOPSYS_UNCONNECTED__224, SYNOPSYS_UNCONNECTED__225, 
        SYNOPSYS_UNCONNECTED__226, SYNOPSYS_UNCONNECTED__227, 
        SYNOPSYS_UNCONNECTED__228, SYNOPSYS_UNCONNECTED__229, 
        SYNOPSYS_UNCONNECTED__230, SYNOPSYS_UNCONNECTED__231, 
        SYNOPSYS_UNCONNECTED__232, SYNOPSYS_UNCONNECTED__233, 
        SYNOPSYS_UNCONNECTED__234, SYNOPSYS_UNCONNECTED__235, 
        SYNOPSYS_UNCONNECTED__236, SYNOPSYS_UNCONNECTED__237, 
        SYNOPSYS_UNCONNECTED__238, SYNOPSYS_UNCONNECTED__239, 
        SYNOPSYS_UNCONNECTED__240, SYNOPSYS_UNCONNECTED__241, 
        SYNOPSYS_UNCONNECTED__242, SYNOPSYS_UNCONNECTED__243, 
        SYNOPSYS_UNCONNECTED__244, SYNOPSYS_UNCONNECTED__245, 
        SYNOPSYS_UNCONNECTED__246, SYNOPSYS_UNCONNECTED__247, 
        SYNOPSYS_UNCONNECTED__248, SYNOPSYS_UNCONNECTED__249, 
        SYNOPSYS_UNCONNECTED__250, SYNOPSYS_UNCONNECTED__251, 
        SYNOPSYS_UNCONNECTED__252, SYNOPSYS_UNCONNECTED__253, 
        SYNOPSYS_UNCONNECTED__254;

  gen_nonlinear_part NLIN ( .a(a), .b(b), .n({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, n[498], 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, n[495:494], 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, n[491], 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, n[488:486], 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, n[483], 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, n[480:479], 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, n[476], 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, n[473:470], 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, n[467], 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, n[464:463], 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, n[460], 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, n[457:455], 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, n[452], 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, n[449:448], 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, n[445], 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, n[442:438], 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, n[435], 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, n[432:431], 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, n[428], 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, n[425:423], 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, n[420], 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, n[417:416], 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, n[413], 
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, n[410:407], 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, n[404], 
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, n[401:400], 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, n[397], 
        SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, n[394:392], 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58, n[389], 
        SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, n[386:385], 
        SYNOPSYS_UNCONNECTED__61, SYNOPSYS_UNCONNECTED__62, n[382], 
        SYNOPSYS_UNCONNECTED__63, SYNOPSYS_UNCONNECTED__64, n[379:374], 
        SYNOPSYS_UNCONNECTED__65, SYNOPSYS_UNCONNECTED__66, n[371], 
        SYNOPSYS_UNCONNECTED__67, SYNOPSYS_UNCONNECTED__68, n[368:367], 
        SYNOPSYS_UNCONNECTED__69, SYNOPSYS_UNCONNECTED__70, n[364], 
        SYNOPSYS_UNCONNECTED__71, SYNOPSYS_UNCONNECTED__72, n[361:359], 
        SYNOPSYS_UNCONNECTED__73, SYNOPSYS_UNCONNECTED__74, n[356], 
        SYNOPSYS_UNCONNECTED__75, SYNOPSYS_UNCONNECTED__76, n[353:352], 
        SYNOPSYS_UNCONNECTED__77, SYNOPSYS_UNCONNECTED__78, n[349], 
        SYNOPSYS_UNCONNECTED__79, SYNOPSYS_UNCONNECTED__80, n[346:343], 
        SYNOPSYS_UNCONNECTED__81, SYNOPSYS_UNCONNECTED__82, n[340], 
        SYNOPSYS_UNCONNECTED__83, SYNOPSYS_UNCONNECTED__84, n[337:336], 
        SYNOPSYS_UNCONNECTED__85, SYNOPSYS_UNCONNECTED__86, n[333], 
        SYNOPSYS_UNCONNECTED__87, SYNOPSYS_UNCONNECTED__88, n[330:328], 
        SYNOPSYS_UNCONNECTED__89, SYNOPSYS_UNCONNECTED__90, n[325], 
        SYNOPSYS_UNCONNECTED__91, SYNOPSYS_UNCONNECTED__92, n[322:321], 
        SYNOPSYS_UNCONNECTED__93, SYNOPSYS_UNCONNECTED__94, n[318], 
        SYNOPSYS_UNCONNECTED__95, SYNOPSYS_UNCONNECTED__96, n[315:311], 
        SYNOPSYS_UNCONNECTED__97, SYNOPSYS_UNCONNECTED__98, n[308], 
        SYNOPSYS_UNCONNECTED__99, SYNOPSYS_UNCONNECTED__100, n[305:304], 
        SYNOPSYS_UNCONNECTED__101, SYNOPSYS_UNCONNECTED__102, n[301], 
        SYNOPSYS_UNCONNECTED__103, SYNOPSYS_UNCONNECTED__104, n[298:296], 
        SYNOPSYS_UNCONNECTED__105, SYNOPSYS_UNCONNECTED__106, n[293], 
        SYNOPSYS_UNCONNECTED__107, SYNOPSYS_UNCONNECTED__108, n[290:289], 
        SYNOPSYS_UNCONNECTED__109, SYNOPSYS_UNCONNECTED__110, n[286], 
        SYNOPSYS_UNCONNECTED__111, SYNOPSYS_UNCONNECTED__112, n[283:280], 
        SYNOPSYS_UNCONNECTED__113, SYNOPSYS_UNCONNECTED__114, n[277], 
        SYNOPSYS_UNCONNECTED__115, SYNOPSYS_UNCONNECTED__116, n[274:273], 
        SYNOPSYS_UNCONNECTED__117, SYNOPSYS_UNCONNECTED__118, n[270], 
        SYNOPSYS_UNCONNECTED__119, SYNOPSYS_UNCONNECTED__120, n[267:265], 
        SYNOPSYS_UNCONNECTED__121, SYNOPSYS_UNCONNECTED__122, n[262], 
        SYNOPSYS_UNCONNECTED__123, SYNOPSYS_UNCONNECTED__124, n[259:258], 
        SYNOPSYS_UNCONNECTED__125, SYNOPSYS_UNCONNECTED__126, n[255], 
        SYNOPSYS_UNCONNECTED__127, SYNOPSYS_UNCONNECTED__128, n[252:246], 
        SYNOPSYS_UNCONNECTED__129, SYNOPSYS_UNCONNECTED__130, n[243], 
        SYNOPSYS_UNCONNECTED__131, SYNOPSYS_UNCONNECTED__132, n[240:239], 
        SYNOPSYS_UNCONNECTED__133, SYNOPSYS_UNCONNECTED__134, n[236], 
        SYNOPSYS_UNCONNECTED__135, SYNOPSYS_UNCONNECTED__136, n[233:231], 
        SYNOPSYS_UNCONNECTED__137, SYNOPSYS_UNCONNECTED__138, n[228], 
        SYNOPSYS_UNCONNECTED__139, SYNOPSYS_UNCONNECTED__140, n[225:224], 
        SYNOPSYS_UNCONNECTED__141, SYNOPSYS_UNCONNECTED__142, n[221], 
        SYNOPSYS_UNCONNECTED__143, SYNOPSYS_UNCONNECTED__144, n[218:215], 
        SYNOPSYS_UNCONNECTED__145, SYNOPSYS_UNCONNECTED__146, n[212], 
        SYNOPSYS_UNCONNECTED__147, SYNOPSYS_UNCONNECTED__148, n[209:208], 
        SYNOPSYS_UNCONNECTED__149, SYNOPSYS_UNCONNECTED__150, n[205], 
        SYNOPSYS_UNCONNECTED__151, SYNOPSYS_UNCONNECTED__152, n[202:200], 
        SYNOPSYS_UNCONNECTED__153, SYNOPSYS_UNCONNECTED__154, n[197], 
        SYNOPSYS_UNCONNECTED__155, SYNOPSYS_UNCONNECTED__156, n[194:193], 
        SYNOPSYS_UNCONNECTED__157, SYNOPSYS_UNCONNECTED__158, n[190], 
        SYNOPSYS_UNCONNECTED__159, SYNOPSYS_UNCONNECTED__160, n[187:183], 
        SYNOPSYS_UNCONNECTED__161, SYNOPSYS_UNCONNECTED__162, n[180], 
        SYNOPSYS_UNCONNECTED__163, SYNOPSYS_UNCONNECTED__164, n[177:176], 
        SYNOPSYS_UNCONNECTED__165, SYNOPSYS_UNCONNECTED__166, n[173], 
        SYNOPSYS_UNCONNECTED__167, SYNOPSYS_UNCONNECTED__168, n[170:168], 
        SYNOPSYS_UNCONNECTED__169, SYNOPSYS_UNCONNECTED__170, n[165], 
        SYNOPSYS_UNCONNECTED__171, SYNOPSYS_UNCONNECTED__172, n[162:161], 
        SYNOPSYS_UNCONNECTED__173, SYNOPSYS_UNCONNECTED__174, n[158], 
        SYNOPSYS_UNCONNECTED__175, SYNOPSYS_UNCONNECTED__176, n[155:152], 
        SYNOPSYS_UNCONNECTED__177, SYNOPSYS_UNCONNECTED__178, n[149], 
        SYNOPSYS_UNCONNECTED__179, SYNOPSYS_UNCONNECTED__180, n[146:145], 
        SYNOPSYS_UNCONNECTED__181, SYNOPSYS_UNCONNECTED__182, n[142], 
        SYNOPSYS_UNCONNECTED__183, SYNOPSYS_UNCONNECTED__184, n[139:137], 
        SYNOPSYS_UNCONNECTED__185, SYNOPSYS_UNCONNECTED__186, n[134], 
        SYNOPSYS_UNCONNECTED__187, SYNOPSYS_UNCONNECTED__188, n[131:130], 
        SYNOPSYS_UNCONNECTED__189, SYNOPSYS_UNCONNECTED__190, n[127], 
        SYNOPSYS_UNCONNECTED__191, SYNOPSYS_UNCONNECTED__192, n[124:119], 
        SYNOPSYS_UNCONNECTED__193, SYNOPSYS_UNCONNECTED__194, n[116], 
        SYNOPSYS_UNCONNECTED__195, SYNOPSYS_UNCONNECTED__196, n[113:112], 
        SYNOPSYS_UNCONNECTED__197, SYNOPSYS_UNCONNECTED__198, n[109], 
        SYNOPSYS_UNCONNECTED__199, SYNOPSYS_UNCONNECTED__200, n[106:104], 
        SYNOPSYS_UNCONNECTED__201, SYNOPSYS_UNCONNECTED__202, n[101], 
        SYNOPSYS_UNCONNECTED__203, SYNOPSYS_UNCONNECTED__204, n[98:97], 
        SYNOPSYS_UNCONNECTED__205, SYNOPSYS_UNCONNECTED__206, n[94], 
        SYNOPSYS_UNCONNECTED__207, SYNOPSYS_UNCONNECTED__208, n[91:88], 
        SYNOPSYS_UNCONNECTED__209, SYNOPSYS_UNCONNECTED__210, n[85], 
        SYNOPSYS_UNCONNECTED__211, SYNOPSYS_UNCONNECTED__212, n[82:81], 
        SYNOPSYS_UNCONNECTED__213, SYNOPSYS_UNCONNECTED__214, n[78], 
        SYNOPSYS_UNCONNECTED__215, SYNOPSYS_UNCONNECTED__216, n[75:73], 
        SYNOPSYS_UNCONNECTED__217, SYNOPSYS_UNCONNECTED__218, n[70], 
        SYNOPSYS_UNCONNECTED__219, SYNOPSYS_UNCONNECTED__220, n[67:66], 
        SYNOPSYS_UNCONNECTED__221, SYNOPSYS_UNCONNECTED__222, n[63], 
        SYNOPSYS_UNCONNECTED__223, SYNOPSYS_UNCONNECTED__224, n[60:56], 
        SYNOPSYS_UNCONNECTED__225, SYNOPSYS_UNCONNECTED__226, n[53], 
        SYNOPSYS_UNCONNECTED__227, SYNOPSYS_UNCONNECTED__228, n[50:49], 
        SYNOPSYS_UNCONNECTED__229, SYNOPSYS_UNCONNECTED__230, n[46], 
        SYNOPSYS_UNCONNECTED__231, SYNOPSYS_UNCONNECTED__232, n[43:41], 
        SYNOPSYS_UNCONNECTED__233, SYNOPSYS_UNCONNECTED__234, n[38], 
        SYNOPSYS_UNCONNECTED__235, SYNOPSYS_UNCONNECTED__236, n[35:34], 
        SYNOPSYS_UNCONNECTED__237, SYNOPSYS_UNCONNECTED__238, n[31], 
        SYNOPSYS_UNCONNECTED__239, SYNOPSYS_UNCONNECTED__240, n[28:25], 
        SYNOPSYS_UNCONNECTED__241, SYNOPSYS_UNCONNECTED__242, n[22], 
        SYNOPSYS_UNCONNECTED__243, SYNOPSYS_UNCONNECTED__244, n[19:18], 
        SYNOPSYS_UNCONNECTED__245, SYNOPSYS_UNCONNECTED__246, n[15], 
        SYNOPSYS_UNCONNECTED__247, SYNOPSYS_UNCONNECTED__248, n[12:10], 
        SYNOPSYS_UNCONNECTED__249, SYNOPSYS_UNCONNECTED__250, n[7], 
        SYNOPSYS_UNCONNECTED__251, SYNOPSYS_UNCONNECTED__252, n[4:3], 
        SYNOPSYS_UNCONNECTED__253, SYNOPSYS_UNCONNECTED__254, n[0]}) );
  gen_linear_part LIN ( .a(a), .b(b), .n({1'b0, 1'b0, 1'b0, n[498], 1'b0, 1'b0, 
        n[495:494], 1'b0, 1'b0, n[491], 1'b0, 1'b0, n[488:486], 1'b0, 1'b0, 
        n[483], 1'b0, 1'b0, n[480:479], 1'b0, 1'b0, n[476], 1'b0, 1'b0, 
        n[473:470], 1'b0, 1'b0, n[467], 1'b0, 1'b0, n[464:463], 1'b0, 1'b0, 
        n[460], 1'b0, 1'b0, n[457:455], 1'b0, 1'b0, n[452], 1'b0, 1'b0, 
        n[449:448], 1'b0, 1'b0, n[445], 1'b0, 1'b0, n[442:438], 1'b0, 1'b0, 
        n[435], 1'b0, 1'b0, n[432:431], 1'b0, 1'b0, n[428], 1'b0, 1'b0, 
        n[425:423], 1'b0, 1'b0, n[420], 1'b0, 1'b0, n[417:416], 1'b0, 1'b0, 
        n[413], 1'b0, 1'b0, n[410:407], 1'b0, 1'b0, n[404], 1'b0, 1'b0, 
        n[401:400], 1'b0, 1'b0, n[397], 1'b0, 1'b0, n[394:392], 1'b0, 1'b0, 
        n[389], 1'b0, 1'b0, n[386:385], 1'b0, 1'b0, n[382], 1'b0, 1'b0, 
        n[379:374], 1'b0, 1'b0, n[371], 1'b0, 1'b0, n[368:367], 1'b0, 1'b0, 
        n[364], 1'b0, 1'b0, n[361:359], 1'b0, 1'b0, n[356], 1'b0, 1'b0, 
        n[353:352], 1'b0, 1'b0, n[349], 1'b0, 1'b0, n[346:343], 1'b0, 1'b0, 
        n[340], 1'b0, 1'b0, n[337:336], 1'b0, 1'b0, n[333], 1'b0, 1'b0, 
        n[330:328], 1'b0, 1'b0, n[325], 1'b0, 1'b0, n[322:321], 1'b0, 1'b0, 
        n[318], 1'b0, 1'b0, n[315:311], 1'b0, 1'b0, n[308], 1'b0, 1'b0, 
        n[305:304], 1'b0, 1'b0, n[301], 1'b0, 1'b0, n[298:296], 1'b0, 1'b0, 
        n[293], 1'b0, 1'b0, n[290:289], 1'b0, 1'b0, n[286], 1'b0, 1'b0, 
        n[283:280], 1'b0, 1'b0, n[277], 1'b0, 1'b0, n[274:273], 1'b0, 1'b0, 
        n[270], 1'b0, 1'b0, n[267:265], 1'b0, 1'b0, n[262], 1'b0, 1'b0, 
        n[259:258], 1'b0, 1'b0, n[255], 1'b0, 1'b0, n[252:246], 1'b0, 1'b0, 
        n[243], 1'b0, 1'b0, n[240:239], 1'b0, 1'b0, n[236], 1'b0, 1'b0, 
        n[233:231], 1'b0, 1'b0, n[228], 1'b0, 1'b0, n[225:224], 1'b0, 1'b0, 
        n[221], 1'b0, 1'b0, n[218:215], 1'b0, 1'b0, n[212], 1'b0, 1'b0, 
        n[209:208], 1'b0, 1'b0, n[205], 1'b0, 1'b0, n[202:200], 1'b0, 1'b0, 
        n[197], 1'b0, 1'b0, n[194:193], 1'b0, 1'b0, n[190], 1'b0, 1'b0, 
        n[187:183], 1'b0, 1'b0, n[180], 1'b0, 1'b0, n[177:176], 1'b0, 1'b0, 
        n[173], 1'b0, 1'b0, n[170:168], 1'b0, 1'b0, n[165], 1'b0, 1'b0, 
        n[162:161], 1'b0, 1'b0, n[158], 1'b0, 1'b0, n[155:152], 1'b0, 1'b0, 
        n[149], 1'b0, 1'b0, n[146:145], 1'b0, 1'b0, n[142], 1'b0, 1'b0, 
        n[139:137], 1'b0, 1'b0, n[134], 1'b0, 1'b0, n[131:130], 1'b0, 1'b0, 
        n[127], 1'b0, 1'b0, n[124:119], 1'b0, 1'b0, n[116], 1'b0, 1'b0, 
        n[113:112], 1'b0, 1'b0, n[109], 1'b0, 1'b0, n[106:104], 1'b0, 1'b0, 
        n[101], 1'b0, 1'b0, n[98:97], 1'b0, 1'b0, n[94], 1'b0, 1'b0, n[91:88], 
        1'b0, 1'b0, n[85], 1'b0, 1'b0, n[82:81], 1'b0, 1'b0, n[78], 1'b0, 1'b0, 
        n[75:73], 1'b0, 1'b0, n[70], 1'b0, 1'b0, n[67:66], 1'b0, 1'b0, n[63], 
        1'b0, 1'b0, n[60:56], 1'b0, 1'b0, n[53], 1'b0, 1'b0, n[50:49], 1'b0, 
        1'b0, n[46], 1'b0, 1'b0, n[43:41], 1'b0, 1'b0, n[38], 1'b0, 1'b0, 
        n[35:34], 1'b0, 1'b0, n[31], 1'b0, 1'b0, n[28:25], 1'b0, 1'b0, n[22], 
        1'b0, 1'b0, n[19:18], 1'b0, 1'b0, n[15], 1'b0, 1'b0, n[12:10], 1'b0, 
        1'b0, n[7], 1'b0, 1'b0, n[4:3], 1'b0, 1'b0, n[0]}), .s(s) );
endmodule

