module normal_adder (a,b,s);
parameter NBIT = 8;
input [NBIT-1:0] a,b;
output reg [NBIT:0] s;
//assign s = a + b;
always @(*)
begin
    casex({a,b})
	{8'd0,8'd0} : s = 0;
	{8'd0,8'd1} : s = 1;
	{8'd0,8'd2} : s = 2;
	{8'd0,8'd3} : s = 3;
	{8'd0,8'd4} : s = 4;
	{8'd0,8'd5} : s = 5;
	{8'd0,8'd6} : s = 6;
	{8'd0,8'd7} : s = 7;
	{8'd0,8'd8} : s = 8;
	{8'd0,8'd9} : s = 9;
	{8'd0,8'd10} : s = 10;
	{8'd0,8'd11} : s = 11;
	{8'd0,8'd12} : s = 12;
	{8'd0,8'd13} : s = 13;
	{8'd0,8'd14} : s = 14;
	{8'd0,8'd15} : s = 15;
	{8'd0,8'd16} : s = 16;
	{8'd0,8'd17} : s = 17;
	{8'd0,8'd18} : s = 18;
	{8'd0,8'd19} : s = 19;
	{8'd0,8'd20} : s = 20;
	{8'd0,8'd21} : s = 21;
	{8'd0,8'd22} : s = 22;
	{8'd0,8'd23} : s = 23;
	{8'd0,8'd24} : s = 24;
	{8'd0,8'd25} : s = 25;
	{8'd0,8'd26} : s = 26;
	{8'd0,8'd27} : s = 27;
	{8'd0,8'd28} : s = 28;
	{8'd0,8'd29} : s = 29;
	{8'd0,8'd30} : s = 30;
	{8'd0,8'd31} : s = 31;
	{8'd0,8'd32} : s = 32;
	{8'd0,8'd33} : s = 33;
	{8'd0,8'd34} : s = 34;
	{8'd0,8'd35} : s = 35;
	{8'd0,8'd36} : s = 36;
	{8'd0,8'd37} : s = 37;
	{8'd0,8'd38} : s = 38;
	{8'd0,8'd39} : s = 39;
	{8'd0,8'd40} : s = 40;
	{8'd0,8'd41} : s = 41;
	{8'd0,8'd42} : s = 42;
	{8'd0,8'd43} : s = 43;
	{8'd0,8'd44} : s = 44;
	{8'd0,8'd45} : s = 45;
	{8'd0,8'd46} : s = 46;
	{8'd0,8'd47} : s = 47;
	{8'd0,8'd48} : s = 48;
	{8'd0,8'd49} : s = 49;
	{8'd0,8'd50} : s = 50;
	{8'd0,8'd51} : s = 51;
	{8'd0,8'd52} : s = 52;
	{8'd0,8'd53} : s = 53;
	{8'd0,8'd54} : s = 54;
	{8'd0,8'd55} : s = 55;
	{8'd0,8'd56} : s = 56;
	{8'd0,8'd57} : s = 57;
	{8'd0,8'd58} : s = 58;
	{8'd0,8'd59} : s = 59;
	{8'd0,8'd60} : s = 60;
	{8'd0,8'd61} : s = 61;
	{8'd0,8'd62} : s = 62;
	{8'd0,8'd63} : s = 63;
	{8'd0,8'd64} : s = 64;
	{8'd0,8'd65} : s = 65;
	{8'd0,8'd66} : s = 66;
	{8'd0,8'd67} : s = 67;
	{8'd0,8'd68} : s = 68;
	{8'd0,8'd69} : s = 69;
	{8'd0,8'd70} : s = 70;
	{8'd0,8'd71} : s = 71;
	{8'd0,8'd72} : s = 72;
	{8'd0,8'd73} : s = 73;
	{8'd0,8'd74} : s = 74;
	{8'd0,8'd75} : s = 75;
	{8'd0,8'd76} : s = 76;
	{8'd0,8'd77} : s = 77;
	{8'd0,8'd78} : s = 78;
	{8'd0,8'd79} : s = 79;
	{8'd0,8'd80} : s = 80;
	{8'd0,8'd81} : s = 81;
	{8'd0,8'd82} : s = 82;
	{8'd0,8'd83} : s = 83;
	{8'd0,8'd84} : s = 84;
	{8'd0,8'd85} : s = 85;
	{8'd0,8'd86} : s = 86;
	{8'd0,8'd87} : s = 87;
	{8'd0,8'd88} : s = 88;
	{8'd0,8'd89} : s = 89;
	{8'd0,8'd90} : s = 90;
	{8'd0,8'd91} : s = 91;
	{8'd0,8'd92} : s = 92;
	{8'd0,8'd93} : s = 93;
	{8'd0,8'd94} : s = 94;
	{8'd0,8'd95} : s = 95;
	{8'd0,8'd96} : s = 96;
	{8'd0,8'd97} : s = 97;
	{8'd0,8'd98} : s = 98;
	{8'd0,8'd99} : s = 99;
	{8'd0,8'd100} : s = 100;
	{8'd0,8'd101} : s = 101;
	{8'd0,8'd102} : s = 102;
	{8'd0,8'd103} : s = 103;
	{8'd0,8'd104} : s = 104;
	{8'd0,8'd105} : s = 105;
	{8'd0,8'd106} : s = 106;
	{8'd0,8'd107} : s = 107;
	{8'd0,8'd108} : s = 108;
	{8'd0,8'd109} : s = 109;
	{8'd0,8'd110} : s = 110;
	{8'd0,8'd111} : s = 111;
	{8'd0,8'd112} : s = 112;
	{8'd0,8'd113} : s = 113;
	{8'd0,8'd114} : s = 114;
	{8'd0,8'd115} : s = 115;
	{8'd0,8'd116} : s = 116;
	{8'd0,8'd117} : s = 117;
	{8'd0,8'd118} : s = 118;
	{8'd0,8'd119} : s = 119;
	{8'd0,8'd120} : s = 120;
	{8'd0,8'd121} : s = 121;
	{8'd0,8'd122} : s = 122;
	{8'd0,8'd123} : s = 123;
	{8'd0,8'd124} : s = 124;
	{8'd0,8'd125} : s = 125;
	{8'd0,8'd126} : s = 126;
	{8'd0,8'd127} : s = 127;
	{8'd0,8'd128} : s = 128;
	{8'd0,8'd129} : s = 129;
	{8'd0,8'd130} : s = 130;
	{8'd0,8'd131} : s = 131;
	{8'd0,8'd132} : s = 132;
	{8'd0,8'd133} : s = 133;
	{8'd0,8'd134} : s = 134;
	{8'd0,8'd135} : s = 135;
	{8'd0,8'd136} : s = 136;
	{8'd0,8'd137} : s = 137;
	{8'd0,8'd138} : s = 138;
	{8'd0,8'd139} : s = 139;
	{8'd0,8'd140} : s = 140;
	{8'd0,8'd141} : s = 141;
	{8'd0,8'd142} : s = 142;
	{8'd0,8'd143} : s = 143;
	{8'd0,8'd144} : s = 144;
	{8'd0,8'd145} : s = 145;
	{8'd0,8'd146} : s = 146;
	{8'd0,8'd147} : s = 147;
	{8'd0,8'd148} : s = 148;
	{8'd0,8'd149} : s = 149;
	{8'd0,8'd150} : s = 150;
	{8'd0,8'd151} : s = 151;
	{8'd0,8'd152} : s = 152;
	{8'd0,8'd153} : s = 153;
	{8'd0,8'd154} : s = 154;
	{8'd0,8'd155} : s = 155;
	{8'd0,8'd156} : s = 156;
	{8'd0,8'd157} : s = 157;
	{8'd0,8'd158} : s = 158;
	{8'd0,8'd159} : s = 159;
	{8'd0,8'd160} : s = 160;
	{8'd0,8'd161} : s = 161;
	{8'd0,8'd162} : s = 162;
	{8'd0,8'd163} : s = 163;
	{8'd0,8'd164} : s = 164;
	{8'd0,8'd165} : s = 165;
	{8'd0,8'd166} : s = 166;
	{8'd0,8'd167} : s = 167;
	{8'd0,8'd168} : s = 168;
	{8'd0,8'd169} : s = 169;
	{8'd0,8'd170} : s = 170;
	{8'd0,8'd171} : s = 171;
	{8'd0,8'd172} : s = 172;
	{8'd0,8'd173} : s = 173;
	{8'd0,8'd174} : s = 174;
	{8'd0,8'd175} : s = 175;
	{8'd0,8'd176} : s = 176;
	{8'd0,8'd177} : s = 177;
	{8'd0,8'd178} : s = 178;
	{8'd0,8'd179} : s = 179;
	{8'd0,8'd180} : s = 180;
	{8'd0,8'd181} : s = 181;
	{8'd0,8'd182} : s = 182;
	{8'd0,8'd183} : s = 183;
	{8'd0,8'd184} : s = 184;
	{8'd0,8'd185} : s = 185;
	{8'd0,8'd186} : s = 186;
	{8'd0,8'd187} : s = 187;
	{8'd0,8'd188} : s = 188;
	{8'd0,8'd189} : s = 189;
	{8'd0,8'd190} : s = 190;
	{8'd0,8'd191} : s = 191;
	{8'd0,8'd192} : s = 192;
	{8'd0,8'd193} : s = 193;
	{8'd0,8'd194} : s = 194;
	{8'd0,8'd195} : s = 195;
	{8'd0,8'd196} : s = 196;
	{8'd0,8'd197} : s = 197;
	{8'd0,8'd198} : s = 198;
	{8'd0,8'd199} : s = 199;
	{8'd0,8'd200} : s = 200;
	{8'd0,8'd201} : s = 201;
	{8'd0,8'd202} : s = 202;
	{8'd0,8'd203} : s = 203;
	{8'd0,8'd204} : s = 204;
	{8'd0,8'd205} : s = 205;
	{8'd0,8'd206} : s = 206;
	{8'd0,8'd207} : s = 207;
	{8'd0,8'd208} : s = 208;
	{8'd0,8'd209} : s = 209;
	{8'd0,8'd210} : s = 210;
	{8'd0,8'd211} : s = 211;
	{8'd0,8'd212} : s = 212;
	{8'd0,8'd213} : s = 213;
	{8'd0,8'd214} : s = 214;
	{8'd0,8'd215} : s = 215;
	{8'd0,8'd216} : s = 216;
	{8'd0,8'd217} : s = 217;
	{8'd0,8'd218} : s = 218;
	{8'd0,8'd219} : s = 219;
	{8'd0,8'd220} : s = 220;
	{8'd0,8'd221} : s = 221;
	{8'd0,8'd222} : s = 222;
	{8'd0,8'd223} : s = 223;
	{8'd0,8'd224} : s = 224;
	{8'd0,8'd225} : s = 225;
	{8'd0,8'd226} : s = 226;
	{8'd0,8'd227} : s = 227;
	{8'd0,8'd228} : s = 228;
	{8'd0,8'd229} : s = 229;
	{8'd0,8'd230} : s = 230;
	{8'd0,8'd231} : s = 231;
	{8'd0,8'd232} : s = 232;
	{8'd0,8'd233} : s = 233;
	{8'd0,8'd234} : s = 234;
	{8'd0,8'd235} : s = 235;
	{8'd0,8'd236} : s = 236;
	{8'd0,8'd237} : s = 237;
	{8'd0,8'd238} : s = 238;
	{8'd0,8'd239} : s = 239;
	{8'd0,8'd240} : s = 240;
	{8'd0,8'd241} : s = 241;
	{8'd0,8'd242} : s = 242;
	{8'd0,8'd243} : s = 243;
	{8'd0,8'd244} : s = 244;
	{8'd0,8'd245} : s = 245;
	{8'd0,8'd246} : s = 246;
	{8'd0,8'd247} : s = 247;
	{8'd0,8'd248} : s = 248;
	{8'd0,8'd249} : s = 249;
	{8'd0,8'd250} : s = 250;
	{8'd0,8'd251} : s = 251;
	{8'd0,8'd252} : s = 252;
	{8'd0,8'd253} : s = 253;
	{8'd0,8'd254} : s = 254;
	{8'd0,8'd255} : s = 255;
	{8'd1,8'd0} : s = 1;
	{8'd1,8'd1} : s = 2;
	{8'd1,8'd2} : s = 3;
	{8'd1,8'd3} : s = 4;
	{8'd1,8'd4} : s = 5;
	{8'd1,8'd5} : s = 6;
	{8'd1,8'd6} : s = 7;
	{8'd1,8'd7} : s = 8;
	{8'd1,8'd8} : s = 9;
	{8'd1,8'd9} : s = 10;
	{8'd1,8'd10} : s = 11;
	{8'd1,8'd11} : s = 12;
	{8'd1,8'd12} : s = 13;
	{8'd1,8'd13} : s = 14;
	{8'd1,8'd14} : s = 15;
	{8'd1,8'd15} : s = 16;
	{8'd1,8'd16} : s = 17;
	{8'd1,8'd17} : s = 18;
	{8'd1,8'd18} : s = 19;
	{8'd1,8'd19} : s = 20;
	{8'd1,8'd20} : s = 21;
	{8'd1,8'd21} : s = 22;
	{8'd1,8'd22} : s = 23;
	{8'd1,8'd23} : s = 24;
	{8'd1,8'd24} : s = 25;
	{8'd1,8'd25} : s = 26;
	{8'd1,8'd26} : s = 27;
	{8'd1,8'd27} : s = 28;
	{8'd1,8'd28} : s = 29;
	{8'd1,8'd29} : s = 30;
	{8'd1,8'd30} : s = 31;
	{8'd1,8'd31} : s = 32;
	{8'd1,8'd32} : s = 33;
	{8'd1,8'd33} : s = 34;
	{8'd1,8'd34} : s = 35;
	{8'd1,8'd35} : s = 36;
	{8'd1,8'd36} : s = 37;
	{8'd1,8'd37} : s = 38;
	{8'd1,8'd38} : s = 39;
	{8'd1,8'd39} : s = 40;
	{8'd1,8'd40} : s = 41;
	{8'd1,8'd41} : s = 42;
	{8'd1,8'd42} : s = 43;
	{8'd1,8'd43} : s = 44;
	{8'd1,8'd44} : s = 45;
	{8'd1,8'd45} : s = 46;
	{8'd1,8'd46} : s = 47;
	{8'd1,8'd47} : s = 48;
	{8'd1,8'd48} : s = 49;
	{8'd1,8'd49} : s = 50;
	{8'd1,8'd50} : s = 51;
	{8'd1,8'd51} : s = 52;
	{8'd1,8'd52} : s = 53;
	{8'd1,8'd53} : s = 54;
	{8'd1,8'd54} : s = 55;
	{8'd1,8'd55} : s = 56;
	{8'd1,8'd56} : s = 57;
	{8'd1,8'd57} : s = 58;
	{8'd1,8'd58} : s = 59;
	{8'd1,8'd59} : s = 60;
	{8'd1,8'd60} : s = 61;
	{8'd1,8'd61} : s = 62;
	{8'd1,8'd62} : s = 63;
	{8'd1,8'd63} : s = 64;
	{8'd1,8'd64} : s = 65;
	{8'd1,8'd65} : s = 66;
	{8'd1,8'd66} : s = 67;
	{8'd1,8'd67} : s = 68;
	{8'd1,8'd68} : s = 69;
	{8'd1,8'd69} : s = 70;
	{8'd1,8'd70} : s = 71;
	{8'd1,8'd71} : s = 72;
	{8'd1,8'd72} : s = 73;
	{8'd1,8'd73} : s = 74;
	{8'd1,8'd74} : s = 75;
	{8'd1,8'd75} : s = 76;
	{8'd1,8'd76} : s = 77;
	{8'd1,8'd77} : s = 78;
	{8'd1,8'd78} : s = 79;
	{8'd1,8'd79} : s = 80;
	{8'd1,8'd80} : s = 81;
	{8'd1,8'd81} : s = 82;
	{8'd1,8'd82} : s = 83;
	{8'd1,8'd83} : s = 84;
	{8'd1,8'd84} : s = 85;
	{8'd1,8'd85} : s = 86;
	{8'd1,8'd86} : s = 87;
	{8'd1,8'd87} : s = 88;
	{8'd1,8'd88} : s = 89;
	{8'd1,8'd89} : s = 90;
	{8'd1,8'd90} : s = 91;
	{8'd1,8'd91} : s = 92;
	{8'd1,8'd92} : s = 93;
	{8'd1,8'd93} : s = 94;
	{8'd1,8'd94} : s = 95;
	{8'd1,8'd95} : s = 96;
	{8'd1,8'd96} : s = 97;
	{8'd1,8'd97} : s = 98;
	{8'd1,8'd98} : s = 99;
	{8'd1,8'd99} : s = 100;
	{8'd1,8'd100} : s = 101;
	{8'd1,8'd101} : s = 102;
	{8'd1,8'd102} : s = 103;
	{8'd1,8'd103} : s = 104;
	{8'd1,8'd104} : s = 105;
	{8'd1,8'd105} : s = 106;
	{8'd1,8'd106} : s = 107;
	{8'd1,8'd107} : s = 108;
	{8'd1,8'd108} : s = 109;
	{8'd1,8'd109} : s = 110;
	{8'd1,8'd110} : s = 111;
	{8'd1,8'd111} : s = 112;
	{8'd1,8'd112} : s = 113;
	{8'd1,8'd113} : s = 114;
	{8'd1,8'd114} : s = 115;
	{8'd1,8'd115} : s = 116;
	{8'd1,8'd116} : s = 117;
	{8'd1,8'd117} : s = 118;
	{8'd1,8'd118} : s = 119;
	{8'd1,8'd119} : s = 120;
	{8'd1,8'd120} : s = 121;
	{8'd1,8'd121} : s = 122;
	{8'd1,8'd122} : s = 123;
	{8'd1,8'd123} : s = 124;
	{8'd1,8'd124} : s = 125;
	{8'd1,8'd125} : s = 126;
	{8'd1,8'd126} : s = 127;
	{8'd1,8'd127} : s = 128;
	{8'd1,8'd128} : s = 129;
	{8'd1,8'd129} : s = 130;
	{8'd1,8'd130} : s = 131;
	{8'd1,8'd131} : s = 132;
	{8'd1,8'd132} : s = 133;
	{8'd1,8'd133} : s = 134;
	{8'd1,8'd134} : s = 135;
	{8'd1,8'd135} : s = 136;
	{8'd1,8'd136} : s = 137;
	{8'd1,8'd137} : s = 138;
	{8'd1,8'd138} : s = 139;
	{8'd1,8'd139} : s = 140;
	{8'd1,8'd140} : s = 141;
	{8'd1,8'd141} : s = 142;
	{8'd1,8'd142} : s = 143;
	{8'd1,8'd143} : s = 144;
	{8'd1,8'd144} : s = 145;
	{8'd1,8'd145} : s = 146;
	{8'd1,8'd146} : s = 147;
	{8'd1,8'd147} : s = 148;
	{8'd1,8'd148} : s = 149;
	{8'd1,8'd149} : s = 150;
	{8'd1,8'd150} : s = 151;
	{8'd1,8'd151} : s = 152;
	{8'd1,8'd152} : s = 153;
	{8'd1,8'd153} : s = 154;
	{8'd1,8'd154} : s = 155;
	{8'd1,8'd155} : s = 156;
	{8'd1,8'd156} : s = 157;
	{8'd1,8'd157} : s = 158;
	{8'd1,8'd158} : s = 159;
	{8'd1,8'd159} : s = 160;
	{8'd1,8'd160} : s = 161;
	{8'd1,8'd161} : s = 162;
	{8'd1,8'd162} : s = 163;
	{8'd1,8'd163} : s = 164;
	{8'd1,8'd164} : s = 165;
	{8'd1,8'd165} : s = 166;
	{8'd1,8'd166} : s = 167;
	{8'd1,8'd167} : s = 168;
	{8'd1,8'd168} : s = 169;
	{8'd1,8'd169} : s = 170;
	{8'd1,8'd170} : s = 171;
	{8'd1,8'd171} : s = 172;
	{8'd1,8'd172} : s = 173;
	{8'd1,8'd173} : s = 174;
	{8'd1,8'd174} : s = 175;
	{8'd1,8'd175} : s = 176;
	{8'd1,8'd176} : s = 177;
	{8'd1,8'd177} : s = 178;
	{8'd1,8'd178} : s = 179;
	{8'd1,8'd179} : s = 180;
	{8'd1,8'd180} : s = 181;
	{8'd1,8'd181} : s = 182;
	{8'd1,8'd182} : s = 183;
	{8'd1,8'd183} : s = 184;
	{8'd1,8'd184} : s = 185;
	{8'd1,8'd185} : s = 186;
	{8'd1,8'd186} : s = 187;
	{8'd1,8'd187} : s = 188;
	{8'd1,8'd188} : s = 189;
	{8'd1,8'd189} : s = 190;
	{8'd1,8'd190} : s = 191;
	{8'd1,8'd191} : s = 192;
	{8'd1,8'd192} : s = 193;
	{8'd1,8'd193} : s = 194;
	{8'd1,8'd194} : s = 195;
	{8'd1,8'd195} : s = 196;
	{8'd1,8'd196} : s = 197;
	{8'd1,8'd197} : s = 198;
	{8'd1,8'd198} : s = 199;
	{8'd1,8'd199} : s = 200;
	{8'd1,8'd200} : s = 201;
	{8'd1,8'd201} : s = 202;
	{8'd1,8'd202} : s = 203;
	{8'd1,8'd203} : s = 204;
	{8'd1,8'd204} : s = 205;
	{8'd1,8'd205} : s = 206;
	{8'd1,8'd206} : s = 207;
	{8'd1,8'd207} : s = 208;
	{8'd1,8'd208} : s = 209;
	{8'd1,8'd209} : s = 210;
	{8'd1,8'd210} : s = 211;
	{8'd1,8'd211} : s = 212;
	{8'd1,8'd212} : s = 213;
	{8'd1,8'd213} : s = 214;
	{8'd1,8'd214} : s = 215;
	{8'd1,8'd215} : s = 216;
	{8'd1,8'd216} : s = 217;
	{8'd1,8'd217} : s = 218;
	{8'd1,8'd218} : s = 219;
	{8'd1,8'd219} : s = 220;
	{8'd1,8'd220} : s = 221;
	{8'd1,8'd221} : s = 222;
	{8'd1,8'd222} : s = 223;
	{8'd1,8'd223} : s = 224;
	{8'd1,8'd224} : s = 225;
	{8'd1,8'd225} : s = 226;
	{8'd1,8'd226} : s = 227;
	{8'd1,8'd227} : s = 228;
	{8'd1,8'd228} : s = 229;
	{8'd1,8'd229} : s = 230;
	{8'd1,8'd230} : s = 231;
	{8'd1,8'd231} : s = 232;
	{8'd1,8'd232} : s = 233;
	{8'd1,8'd233} : s = 234;
	{8'd1,8'd234} : s = 235;
	{8'd1,8'd235} : s = 236;
	{8'd1,8'd236} : s = 237;
	{8'd1,8'd237} : s = 238;
	{8'd1,8'd238} : s = 239;
	{8'd1,8'd239} : s = 240;
	{8'd1,8'd240} : s = 241;
	{8'd1,8'd241} : s = 242;
	{8'd1,8'd242} : s = 243;
	{8'd1,8'd243} : s = 244;
	{8'd1,8'd244} : s = 245;
	{8'd1,8'd245} : s = 246;
	{8'd1,8'd246} : s = 247;
	{8'd1,8'd247} : s = 248;
	{8'd1,8'd248} : s = 249;
	{8'd1,8'd249} : s = 250;
	{8'd1,8'd250} : s = 251;
	{8'd1,8'd251} : s = 252;
	{8'd1,8'd252} : s = 253;
	{8'd1,8'd253} : s = 254;
	{8'd1,8'd254} : s = 255;
	{8'd1,8'd255} : s = 256;
	{8'd2,8'd0} : s = 2;
	{8'd2,8'd1} : s = 3;
	{8'd2,8'd2} : s = 4;
	{8'd2,8'd3} : s = 5;
	{8'd2,8'd4} : s = 6;
	{8'd2,8'd5} : s = 7;
	{8'd2,8'd6} : s = 8;
	{8'd2,8'd7} : s = 9;
	{8'd2,8'd8} : s = 10;
	{8'd2,8'd9} : s = 11;
	{8'd2,8'd10} : s = 12;
	{8'd2,8'd11} : s = 13;
	{8'd2,8'd12} : s = 14;
	{8'd2,8'd13} : s = 15;
	{8'd2,8'd14} : s = 16;
	{8'd2,8'd15} : s = 17;
	{8'd2,8'd16} : s = 18;
	{8'd2,8'd17} : s = 19;
	{8'd2,8'd18} : s = 20;
	{8'd2,8'd19} : s = 21;
	{8'd2,8'd20} : s = 22;
	{8'd2,8'd21} : s = 23;
	{8'd2,8'd22} : s = 24;
	{8'd2,8'd23} : s = 25;
	{8'd2,8'd24} : s = 26;
	{8'd2,8'd25} : s = 27;
	{8'd2,8'd26} : s = 28;
	{8'd2,8'd27} : s = 29;
	{8'd2,8'd28} : s = 30;
	{8'd2,8'd29} : s = 31;
	{8'd2,8'd30} : s = 32;
	{8'd2,8'd31} : s = 33;
	{8'd2,8'd32} : s = 34;
	{8'd2,8'd33} : s = 35;
	{8'd2,8'd34} : s = 36;
	{8'd2,8'd35} : s = 37;
	{8'd2,8'd36} : s = 38;
	{8'd2,8'd37} : s = 39;
	{8'd2,8'd38} : s = 40;
	{8'd2,8'd39} : s = 41;
	{8'd2,8'd40} : s = 42;
	{8'd2,8'd41} : s = 43;
	{8'd2,8'd42} : s = 44;
	{8'd2,8'd43} : s = 45;
	{8'd2,8'd44} : s = 46;
	{8'd2,8'd45} : s = 47;
	{8'd2,8'd46} : s = 48;
	{8'd2,8'd47} : s = 49;
	{8'd2,8'd48} : s = 50;
	{8'd2,8'd49} : s = 51;
	{8'd2,8'd50} : s = 52;
	{8'd2,8'd51} : s = 53;
	{8'd2,8'd52} : s = 54;
	{8'd2,8'd53} : s = 55;
	{8'd2,8'd54} : s = 56;
	{8'd2,8'd55} : s = 57;
	{8'd2,8'd56} : s = 58;
	{8'd2,8'd57} : s = 59;
	{8'd2,8'd58} : s = 60;
	{8'd2,8'd59} : s = 61;
	{8'd2,8'd60} : s = 62;
	{8'd2,8'd61} : s = 63;
	{8'd2,8'd62} : s = 64;
	{8'd2,8'd63} : s = 65;
	{8'd2,8'd64} : s = 66;
	{8'd2,8'd65} : s = 67;
	{8'd2,8'd66} : s = 68;
	{8'd2,8'd67} : s = 69;
	{8'd2,8'd68} : s = 70;
	{8'd2,8'd69} : s = 71;
	{8'd2,8'd70} : s = 72;
	{8'd2,8'd71} : s = 73;
	{8'd2,8'd72} : s = 74;
	{8'd2,8'd73} : s = 75;
	{8'd2,8'd74} : s = 76;
	{8'd2,8'd75} : s = 77;
	{8'd2,8'd76} : s = 78;
	{8'd2,8'd77} : s = 79;
	{8'd2,8'd78} : s = 80;
	{8'd2,8'd79} : s = 81;
	{8'd2,8'd80} : s = 82;
	{8'd2,8'd81} : s = 83;
	{8'd2,8'd82} : s = 84;
	{8'd2,8'd83} : s = 85;
	{8'd2,8'd84} : s = 86;
	{8'd2,8'd85} : s = 87;
	{8'd2,8'd86} : s = 88;
	{8'd2,8'd87} : s = 89;
	{8'd2,8'd88} : s = 90;
	{8'd2,8'd89} : s = 91;
	{8'd2,8'd90} : s = 92;
	{8'd2,8'd91} : s = 93;
	{8'd2,8'd92} : s = 94;
	{8'd2,8'd93} : s = 95;
	{8'd2,8'd94} : s = 96;
	{8'd2,8'd95} : s = 97;
	{8'd2,8'd96} : s = 98;
	{8'd2,8'd97} : s = 99;
	{8'd2,8'd98} : s = 100;
	{8'd2,8'd99} : s = 101;
	{8'd2,8'd100} : s = 102;
	{8'd2,8'd101} : s = 103;
	{8'd2,8'd102} : s = 104;
	{8'd2,8'd103} : s = 105;
	{8'd2,8'd104} : s = 106;
	{8'd2,8'd105} : s = 107;
	{8'd2,8'd106} : s = 108;
	{8'd2,8'd107} : s = 109;
	{8'd2,8'd108} : s = 110;
	{8'd2,8'd109} : s = 111;
	{8'd2,8'd110} : s = 112;
	{8'd2,8'd111} : s = 113;
	{8'd2,8'd112} : s = 114;
	{8'd2,8'd113} : s = 115;
	{8'd2,8'd114} : s = 116;
	{8'd2,8'd115} : s = 117;
	{8'd2,8'd116} : s = 118;
	{8'd2,8'd117} : s = 119;
	{8'd2,8'd118} : s = 120;
	{8'd2,8'd119} : s = 121;
	{8'd2,8'd120} : s = 122;
	{8'd2,8'd121} : s = 123;
	{8'd2,8'd122} : s = 124;
	{8'd2,8'd123} : s = 125;
	{8'd2,8'd124} : s = 126;
	{8'd2,8'd125} : s = 127;
	{8'd2,8'd126} : s = 128;
	{8'd2,8'd127} : s = 129;
	{8'd2,8'd128} : s = 130;
	{8'd2,8'd129} : s = 131;
	{8'd2,8'd130} : s = 132;
	{8'd2,8'd131} : s = 133;
	{8'd2,8'd132} : s = 134;
	{8'd2,8'd133} : s = 135;
	{8'd2,8'd134} : s = 136;
	{8'd2,8'd135} : s = 137;
	{8'd2,8'd136} : s = 138;
	{8'd2,8'd137} : s = 139;
	{8'd2,8'd138} : s = 140;
	{8'd2,8'd139} : s = 141;
	{8'd2,8'd140} : s = 142;
	{8'd2,8'd141} : s = 143;
	{8'd2,8'd142} : s = 144;
	{8'd2,8'd143} : s = 145;
	{8'd2,8'd144} : s = 146;
	{8'd2,8'd145} : s = 147;
	{8'd2,8'd146} : s = 148;
	{8'd2,8'd147} : s = 149;
	{8'd2,8'd148} : s = 150;
	{8'd2,8'd149} : s = 151;
	{8'd2,8'd150} : s = 152;
	{8'd2,8'd151} : s = 153;
	{8'd2,8'd152} : s = 154;
	{8'd2,8'd153} : s = 155;
	{8'd2,8'd154} : s = 156;
	{8'd2,8'd155} : s = 157;
	{8'd2,8'd156} : s = 158;
	{8'd2,8'd157} : s = 159;
	{8'd2,8'd158} : s = 160;
	{8'd2,8'd159} : s = 161;
	{8'd2,8'd160} : s = 162;
	{8'd2,8'd161} : s = 163;
	{8'd2,8'd162} : s = 164;
	{8'd2,8'd163} : s = 165;
	{8'd2,8'd164} : s = 166;
	{8'd2,8'd165} : s = 167;
	{8'd2,8'd166} : s = 168;
	{8'd2,8'd167} : s = 169;
	{8'd2,8'd168} : s = 170;
	{8'd2,8'd169} : s = 171;
	{8'd2,8'd170} : s = 172;
	{8'd2,8'd171} : s = 173;
	{8'd2,8'd172} : s = 174;
	{8'd2,8'd173} : s = 175;
	{8'd2,8'd174} : s = 176;
	{8'd2,8'd175} : s = 177;
	{8'd2,8'd176} : s = 178;
	{8'd2,8'd177} : s = 179;
	{8'd2,8'd178} : s = 180;
	{8'd2,8'd179} : s = 181;
	{8'd2,8'd180} : s = 182;
	{8'd2,8'd181} : s = 183;
	{8'd2,8'd182} : s = 184;
	{8'd2,8'd183} : s = 185;
	{8'd2,8'd184} : s = 186;
	{8'd2,8'd185} : s = 187;
	{8'd2,8'd186} : s = 188;
	{8'd2,8'd187} : s = 189;
	{8'd2,8'd188} : s = 190;
	{8'd2,8'd189} : s = 191;
	{8'd2,8'd190} : s = 192;
	{8'd2,8'd191} : s = 193;
	{8'd2,8'd192} : s = 194;
	{8'd2,8'd193} : s = 195;
	{8'd2,8'd194} : s = 196;
	{8'd2,8'd195} : s = 197;
	{8'd2,8'd196} : s = 198;
	{8'd2,8'd197} : s = 199;
	{8'd2,8'd198} : s = 200;
	{8'd2,8'd199} : s = 201;
	{8'd2,8'd200} : s = 202;
	{8'd2,8'd201} : s = 203;
	{8'd2,8'd202} : s = 204;
	{8'd2,8'd203} : s = 205;
	{8'd2,8'd204} : s = 206;
	{8'd2,8'd205} : s = 207;
	{8'd2,8'd206} : s = 208;
	{8'd2,8'd207} : s = 209;
	{8'd2,8'd208} : s = 210;
	{8'd2,8'd209} : s = 211;
	{8'd2,8'd210} : s = 212;
	{8'd2,8'd211} : s = 213;
	{8'd2,8'd212} : s = 214;
	{8'd2,8'd213} : s = 215;
	{8'd2,8'd214} : s = 216;
	{8'd2,8'd215} : s = 217;
	{8'd2,8'd216} : s = 218;
	{8'd2,8'd217} : s = 219;
	{8'd2,8'd218} : s = 220;
	{8'd2,8'd219} : s = 221;
	{8'd2,8'd220} : s = 222;
	{8'd2,8'd221} : s = 223;
	{8'd2,8'd222} : s = 224;
	{8'd2,8'd223} : s = 225;
	{8'd2,8'd224} : s = 226;
	{8'd2,8'd225} : s = 227;
	{8'd2,8'd226} : s = 228;
	{8'd2,8'd227} : s = 229;
	{8'd2,8'd228} : s = 230;
	{8'd2,8'd229} : s = 231;
	{8'd2,8'd230} : s = 232;
	{8'd2,8'd231} : s = 233;
	{8'd2,8'd232} : s = 234;
	{8'd2,8'd233} : s = 235;
	{8'd2,8'd234} : s = 236;
	{8'd2,8'd235} : s = 237;
	{8'd2,8'd236} : s = 238;
	{8'd2,8'd237} : s = 239;
	{8'd2,8'd238} : s = 240;
	{8'd2,8'd239} : s = 241;
	{8'd2,8'd240} : s = 242;
	{8'd2,8'd241} : s = 243;
	{8'd2,8'd242} : s = 244;
	{8'd2,8'd243} : s = 245;
	{8'd2,8'd244} : s = 246;
	{8'd2,8'd245} : s = 247;
	{8'd2,8'd246} : s = 248;
	{8'd2,8'd247} : s = 249;
	{8'd2,8'd248} : s = 250;
	{8'd2,8'd249} : s = 251;
	{8'd2,8'd250} : s = 252;
	{8'd2,8'd251} : s = 253;
	{8'd2,8'd252} : s = 254;
	{8'd2,8'd253} : s = 255;
	{8'd2,8'd254} : s = 256;
	{8'd2,8'd255} : s = 257;
	{8'd3,8'd0} : s = 3;
	{8'd3,8'd1} : s = 4;
	{8'd3,8'd2} : s = 5;
	{8'd3,8'd3} : s = 6;
	{8'd3,8'd4} : s = 7;
	{8'd3,8'd5} : s = 8;
	{8'd3,8'd6} : s = 9;
	{8'd3,8'd7} : s = 10;
	{8'd3,8'd8} : s = 11;
	{8'd3,8'd9} : s = 12;
	{8'd3,8'd10} : s = 13;
	{8'd3,8'd11} : s = 14;
	{8'd3,8'd12} : s = 15;
	{8'd3,8'd13} : s = 16;
	{8'd3,8'd14} : s = 17;
	{8'd3,8'd15} : s = 18;
	{8'd3,8'd16} : s = 19;
	{8'd3,8'd17} : s = 20;
	{8'd3,8'd18} : s = 21;
	{8'd3,8'd19} : s = 22;
	{8'd3,8'd20} : s = 23;
	{8'd3,8'd21} : s = 24;
	{8'd3,8'd22} : s = 25;
	{8'd3,8'd23} : s = 26;
	{8'd3,8'd24} : s = 27;
	{8'd3,8'd25} : s = 28;
	{8'd3,8'd26} : s = 29;
	{8'd3,8'd27} : s = 30;
	{8'd3,8'd28} : s = 31;
	{8'd3,8'd29} : s = 32;
	{8'd3,8'd30} : s = 33;
	{8'd3,8'd31} : s = 34;
	{8'd3,8'd32} : s = 35;
	{8'd3,8'd33} : s = 36;
	{8'd3,8'd34} : s = 37;
	{8'd3,8'd35} : s = 38;
	{8'd3,8'd36} : s = 39;
	{8'd3,8'd37} : s = 40;
	{8'd3,8'd38} : s = 41;
	{8'd3,8'd39} : s = 42;
	{8'd3,8'd40} : s = 43;
	{8'd3,8'd41} : s = 44;
	{8'd3,8'd42} : s = 45;
	{8'd3,8'd43} : s = 46;
	{8'd3,8'd44} : s = 47;
	{8'd3,8'd45} : s = 48;
	{8'd3,8'd46} : s = 49;
	{8'd3,8'd47} : s = 50;
	{8'd3,8'd48} : s = 51;
	{8'd3,8'd49} : s = 52;
	{8'd3,8'd50} : s = 53;
	{8'd3,8'd51} : s = 54;
	{8'd3,8'd52} : s = 55;
	{8'd3,8'd53} : s = 56;
	{8'd3,8'd54} : s = 57;
	{8'd3,8'd55} : s = 58;
	{8'd3,8'd56} : s = 59;
	{8'd3,8'd57} : s = 60;
	{8'd3,8'd58} : s = 61;
	{8'd3,8'd59} : s = 62;
	{8'd3,8'd60} : s = 63;
	{8'd3,8'd61} : s = 64;
	{8'd3,8'd62} : s = 65;
	{8'd3,8'd63} : s = 66;
	{8'd3,8'd64} : s = 67;
	{8'd3,8'd65} : s = 68;
	{8'd3,8'd66} : s = 69;
	{8'd3,8'd67} : s = 70;
	{8'd3,8'd68} : s = 71;
	{8'd3,8'd69} : s = 72;
	{8'd3,8'd70} : s = 73;
	{8'd3,8'd71} : s = 74;
	{8'd3,8'd72} : s = 75;
	{8'd3,8'd73} : s = 76;
	{8'd3,8'd74} : s = 77;
	{8'd3,8'd75} : s = 78;
	{8'd3,8'd76} : s = 79;
	{8'd3,8'd77} : s = 80;
	{8'd3,8'd78} : s = 81;
	{8'd3,8'd79} : s = 82;
	{8'd3,8'd80} : s = 83;
	{8'd3,8'd81} : s = 84;
	{8'd3,8'd82} : s = 85;
	{8'd3,8'd83} : s = 86;
	{8'd3,8'd84} : s = 87;
	{8'd3,8'd85} : s = 88;
	{8'd3,8'd86} : s = 89;
	{8'd3,8'd87} : s = 90;
	{8'd3,8'd88} : s = 91;
	{8'd3,8'd89} : s = 92;
	{8'd3,8'd90} : s = 93;
	{8'd3,8'd91} : s = 94;
	{8'd3,8'd92} : s = 95;
	{8'd3,8'd93} : s = 96;
	{8'd3,8'd94} : s = 97;
	{8'd3,8'd95} : s = 98;
	{8'd3,8'd96} : s = 99;
	{8'd3,8'd97} : s = 100;
	{8'd3,8'd98} : s = 101;
	{8'd3,8'd99} : s = 102;
	{8'd3,8'd100} : s = 103;
	{8'd3,8'd101} : s = 104;
	{8'd3,8'd102} : s = 105;
	{8'd3,8'd103} : s = 106;
	{8'd3,8'd104} : s = 107;
	{8'd3,8'd105} : s = 108;
	{8'd3,8'd106} : s = 109;
	{8'd3,8'd107} : s = 110;
	{8'd3,8'd108} : s = 111;
	{8'd3,8'd109} : s = 112;
	{8'd3,8'd110} : s = 113;
	{8'd3,8'd111} : s = 114;
	{8'd3,8'd112} : s = 115;
	{8'd3,8'd113} : s = 116;
	{8'd3,8'd114} : s = 117;
	{8'd3,8'd115} : s = 118;
	{8'd3,8'd116} : s = 119;
	{8'd3,8'd117} : s = 120;
	{8'd3,8'd118} : s = 121;
	{8'd3,8'd119} : s = 122;
	{8'd3,8'd120} : s = 123;
	{8'd3,8'd121} : s = 124;
	{8'd3,8'd122} : s = 125;
	{8'd3,8'd123} : s = 126;
	{8'd3,8'd124} : s = 127;
	{8'd3,8'd125} : s = 128;
	{8'd3,8'd126} : s = 129;
	{8'd3,8'd127} : s = 130;
	{8'd3,8'd128} : s = 131;
	{8'd3,8'd129} : s = 132;
	{8'd3,8'd130} : s = 133;
	{8'd3,8'd131} : s = 134;
	{8'd3,8'd132} : s = 135;
	{8'd3,8'd133} : s = 136;
	{8'd3,8'd134} : s = 137;
	{8'd3,8'd135} : s = 138;
	{8'd3,8'd136} : s = 139;
	{8'd3,8'd137} : s = 140;
	{8'd3,8'd138} : s = 141;
	{8'd3,8'd139} : s = 142;
	{8'd3,8'd140} : s = 143;
	{8'd3,8'd141} : s = 144;
	{8'd3,8'd142} : s = 145;
	{8'd3,8'd143} : s = 146;
	{8'd3,8'd144} : s = 147;
	{8'd3,8'd145} : s = 148;
	{8'd3,8'd146} : s = 149;
	{8'd3,8'd147} : s = 150;
	{8'd3,8'd148} : s = 151;
	{8'd3,8'd149} : s = 152;
	{8'd3,8'd150} : s = 153;
	{8'd3,8'd151} : s = 154;
	{8'd3,8'd152} : s = 155;
	{8'd3,8'd153} : s = 156;
	{8'd3,8'd154} : s = 157;
	{8'd3,8'd155} : s = 158;
	{8'd3,8'd156} : s = 159;
	{8'd3,8'd157} : s = 160;
	{8'd3,8'd158} : s = 161;
	{8'd3,8'd159} : s = 162;
	{8'd3,8'd160} : s = 163;
	{8'd3,8'd161} : s = 164;
	{8'd3,8'd162} : s = 165;
	{8'd3,8'd163} : s = 166;
	{8'd3,8'd164} : s = 167;
	{8'd3,8'd165} : s = 168;
	{8'd3,8'd166} : s = 169;
	{8'd3,8'd167} : s = 170;
	{8'd3,8'd168} : s = 171;
	{8'd3,8'd169} : s = 172;
	{8'd3,8'd170} : s = 173;
	{8'd3,8'd171} : s = 174;
	{8'd3,8'd172} : s = 175;
	{8'd3,8'd173} : s = 176;
	{8'd3,8'd174} : s = 177;
	{8'd3,8'd175} : s = 178;
	{8'd3,8'd176} : s = 179;
	{8'd3,8'd177} : s = 180;
	{8'd3,8'd178} : s = 181;
	{8'd3,8'd179} : s = 182;
	{8'd3,8'd180} : s = 183;
	{8'd3,8'd181} : s = 184;
	{8'd3,8'd182} : s = 185;
	{8'd3,8'd183} : s = 186;
	{8'd3,8'd184} : s = 187;
	{8'd3,8'd185} : s = 188;
	{8'd3,8'd186} : s = 189;
	{8'd3,8'd187} : s = 190;
	{8'd3,8'd188} : s = 191;
	{8'd3,8'd189} : s = 192;
	{8'd3,8'd190} : s = 193;
	{8'd3,8'd191} : s = 194;
	{8'd3,8'd192} : s = 195;
	{8'd3,8'd193} : s = 196;
	{8'd3,8'd194} : s = 197;
	{8'd3,8'd195} : s = 198;
	{8'd3,8'd196} : s = 199;
	{8'd3,8'd197} : s = 200;
	{8'd3,8'd198} : s = 201;
	{8'd3,8'd199} : s = 202;
	{8'd3,8'd200} : s = 203;
	{8'd3,8'd201} : s = 204;
	{8'd3,8'd202} : s = 205;
	{8'd3,8'd203} : s = 206;
	{8'd3,8'd204} : s = 207;
	{8'd3,8'd205} : s = 208;
	{8'd3,8'd206} : s = 209;
	{8'd3,8'd207} : s = 210;
	{8'd3,8'd208} : s = 211;
	{8'd3,8'd209} : s = 212;
	{8'd3,8'd210} : s = 213;
	{8'd3,8'd211} : s = 214;
	{8'd3,8'd212} : s = 215;
	{8'd3,8'd213} : s = 216;
	{8'd3,8'd214} : s = 217;
	{8'd3,8'd215} : s = 218;
	{8'd3,8'd216} : s = 219;
	{8'd3,8'd217} : s = 220;
	{8'd3,8'd218} : s = 221;
	{8'd3,8'd219} : s = 222;
	{8'd3,8'd220} : s = 223;
	{8'd3,8'd221} : s = 224;
	{8'd3,8'd222} : s = 225;
	{8'd3,8'd223} : s = 226;
	{8'd3,8'd224} : s = 227;
	{8'd3,8'd225} : s = 228;
	{8'd3,8'd226} : s = 229;
	{8'd3,8'd227} : s = 230;
	{8'd3,8'd228} : s = 231;
	{8'd3,8'd229} : s = 232;
	{8'd3,8'd230} : s = 233;
	{8'd3,8'd231} : s = 234;
	{8'd3,8'd232} : s = 235;
	{8'd3,8'd233} : s = 236;
	{8'd3,8'd234} : s = 237;
	{8'd3,8'd235} : s = 238;
	{8'd3,8'd236} : s = 239;
	{8'd3,8'd237} : s = 240;
	{8'd3,8'd238} : s = 241;
	{8'd3,8'd239} : s = 242;
	{8'd3,8'd240} : s = 243;
	{8'd3,8'd241} : s = 244;
	{8'd3,8'd242} : s = 245;
	{8'd3,8'd243} : s = 246;
	{8'd3,8'd244} : s = 247;
	{8'd3,8'd245} : s = 248;
	{8'd3,8'd246} : s = 249;
	{8'd3,8'd247} : s = 250;
	{8'd3,8'd248} : s = 251;
	{8'd3,8'd249} : s = 252;
	{8'd3,8'd250} : s = 253;
	{8'd3,8'd251} : s = 254;
	{8'd3,8'd252} : s = 255;
	{8'd3,8'd253} : s = 256;
	{8'd3,8'd254} : s = 257;
	{8'd3,8'd255} : s = 258;
	{8'd4,8'd0} : s = 4;
	{8'd4,8'd1} : s = 5;
	{8'd4,8'd2} : s = 6;
	{8'd4,8'd3} : s = 7;
	{8'd4,8'd4} : s = 8;
	{8'd4,8'd5} : s = 9;
	{8'd4,8'd6} : s = 10;
	{8'd4,8'd7} : s = 11;
	{8'd4,8'd8} : s = 12;
	{8'd4,8'd9} : s = 13;
	{8'd4,8'd10} : s = 14;
	{8'd4,8'd11} : s = 15;
	{8'd4,8'd12} : s = 16;
	{8'd4,8'd13} : s = 17;
	{8'd4,8'd14} : s = 18;
	{8'd4,8'd15} : s = 19;
	{8'd4,8'd16} : s = 20;
	{8'd4,8'd17} : s = 21;
	{8'd4,8'd18} : s = 22;
	{8'd4,8'd19} : s = 23;
	{8'd4,8'd20} : s = 24;
	{8'd4,8'd21} : s = 25;
	{8'd4,8'd22} : s = 26;
	{8'd4,8'd23} : s = 27;
	{8'd4,8'd24} : s = 28;
	{8'd4,8'd25} : s = 29;
	{8'd4,8'd26} : s = 30;
	{8'd4,8'd27} : s = 31;
	{8'd4,8'd28} : s = 32;
	{8'd4,8'd29} : s = 33;
	{8'd4,8'd30} : s = 34;
	{8'd4,8'd31} : s = 35;
	{8'd4,8'd32} : s = 36;
	{8'd4,8'd33} : s = 37;
	{8'd4,8'd34} : s = 38;
	{8'd4,8'd35} : s = 39;
	{8'd4,8'd36} : s = 40;
	{8'd4,8'd37} : s = 41;
	{8'd4,8'd38} : s = 42;
	{8'd4,8'd39} : s = 43;
	{8'd4,8'd40} : s = 44;
	{8'd4,8'd41} : s = 45;
	{8'd4,8'd42} : s = 46;
	{8'd4,8'd43} : s = 47;
	{8'd4,8'd44} : s = 48;
	{8'd4,8'd45} : s = 49;
	{8'd4,8'd46} : s = 50;
	{8'd4,8'd47} : s = 51;
	{8'd4,8'd48} : s = 52;
	{8'd4,8'd49} : s = 53;
	{8'd4,8'd50} : s = 54;
	{8'd4,8'd51} : s = 55;
	{8'd4,8'd52} : s = 56;
	{8'd4,8'd53} : s = 57;
	{8'd4,8'd54} : s = 58;
	{8'd4,8'd55} : s = 59;
	{8'd4,8'd56} : s = 60;
	{8'd4,8'd57} : s = 61;
	{8'd4,8'd58} : s = 62;
	{8'd4,8'd59} : s = 63;
	{8'd4,8'd60} : s = 64;
	{8'd4,8'd61} : s = 65;
	{8'd4,8'd62} : s = 66;
	{8'd4,8'd63} : s = 67;
	{8'd4,8'd64} : s = 68;
	{8'd4,8'd65} : s = 69;
	{8'd4,8'd66} : s = 70;
	{8'd4,8'd67} : s = 71;
	{8'd4,8'd68} : s = 72;
	{8'd4,8'd69} : s = 73;
	{8'd4,8'd70} : s = 74;
	{8'd4,8'd71} : s = 75;
	{8'd4,8'd72} : s = 76;
	{8'd4,8'd73} : s = 77;
	{8'd4,8'd74} : s = 78;
	{8'd4,8'd75} : s = 79;
	{8'd4,8'd76} : s = 80;
	{8'd4,8'd77} : s = 81;
	{8'd4,8'd78} : s = 82;
	{8'd4,8'd79} : s = 83;
	{8'd4,8'd80} : s = 84;
	{8'd4,8'd81} : s = 85;
	{8'd4,8'd82} : s = 86;
	{8'd4,8'd83} : s = 87;
	{8'd4,8'd84} : s = 88;
	{8'd4,8'd85} : s = 89;
	{8'd4,8'd86} : s = 90;
	{8'd4,8'd87} : s = 91;
	{8'd4,8'd88} : s = 92;
	{8'd4,8'd89} : s = 93;
	{8'd4,8'd90} : s = 94;
	{8'd4,8'd91} : s = 95;
	{8'd4,8'd92} : s = 96;
	{8'd4,8'd93} : s = 97;
	{8'd4,8'd94} : s = 98;
	{8'd4,8'd95} : s = 99;
	{8'd4,8'd96} : s = 100;
	{8'd4,8'd97} : s = 101;
	{8'd4,8'd98} : s = 102;
	{8'd4,8'd99} : s = 103;
	{8'd4,8'd100} : s = 104;
	{8'd4,8'd101} : s = 105;
	{8'd4,8'd102} : s = 106;
	{8'd4,8'd103} : s = 107;
	{8'd4,8'd104} : s = 108;
	{8'd4,8'd105} : s = 109;
	{8'd4,8'd106} : s = 110;
	{8'd4,8'd107} : s = 111;
	{8'd4,8'd108} : s = 112;
	{8'd4,8'd109} : s = 113;
	{8'd4,8'd110} : s = 114;
	{8'd4,8'd111} : s = 115;
	{8'd4,8'd112} : s = 116;
	{8'd4,8'd113} : s = 117;
	{8'd4,8'd114} : s = 118;
	{8'd4,8'd115} : s = 119;
	{8'd4,8'd116} : s = 120;
	{8'd4,8'd117} : s = 121;
	{8'd4,8'd118} : s = 122;
	{8'd4,8'd119} : s = 123;
	{8'd4,8'd120} : s = 124;
	{8'd4,8'd121} : s = 125;
	{8'd4,8'd122} : s = 126;
	{8'd4,8'd123} : s = 127;
	{8'd4,8'd124} : s = 128;
	{8'd4,8'd125} : s = 129;
	{8'd4,8'd126} : s = 130;
	{8'd4,8'd127} : s = 131;
	{8'd4,8'd128} : s = 132;
	{8'd4,8'd129} : s = 133;
	{8'd4,8'd130} : s = 134;
	{8'd4,8'd131} : s = 135;
	{8'd4,8'd132} : s = 136;
	{8'd4,8'd133} : s = 137;
	{8'd4,8'd134} : s = 138;
	{8'd4,8'd135} : s = 139;
	{8'd4,8'd136} : s = 140;
	{8'd4,8'd137} : s = 141;
	{8'd4,8'd138} : s = 142;
	{8'd4,8'd139} : s = 143;
	{8'd4,8'd140} : s = 144;
	{8'd4,8'd141} : s = 145;
	{8'd4,8'd142} : s = 146;
	{8'd4,8'd143} : s = 147;
	{8'd4,8'd144} : s = 148;
	{8'd4,8'd145} : s = 149;
	{8'd4,8'd146} : s = 150;
	{8'd4,8'd147} : s = 151;
	{8'd4,8'd148} : s = 152;
	{8'd4,8'd149} : s = 153;
	{8'd4,8'd150} : s = 154;
	{8'd4,8'd151} : s = 155;
	{8'd4,8'd152} : s = 156;
	{8'd4,8'd153} : s = 157;
	{8'd4,8'd154} : s = 158;
	{8'd4,8'd155} : s = 159;
	{8'd4,8'd156} : s = 160;
	{8'd4,8'd157} : s = 161;
	{8'd4,8'd158} : s = 162;
	{8'd4,8'd159} : s = 163;
	{8'd4,8'd160} : s = 164;
	{8'd4,8'd161} : s = 165;
	{8'd4,8'd162} : s = 166;
	{8'd4,8'd163} : s = 167;
	{8'd4,8'd164} : s = 168;
	{8'd4,8'd165} : s = 169;
	{8'd4,8'd166} : s = 170;
	{8'd4,8'd167} : s = 171;
	{8'd4,8'd168} : s = 172;
	{8'd4,8'd169} : s = 173;
	{8'd4,8'd170} : s = 174;
	{8'd4,8'd171} : s = 175;
	{8'd4,8'd172} : s = 176;
	{8'd4,8'd173} : s = 177;
	{8'd4,8'd174} : s = 178;
	{8'd4,8'd175} : s = 179;
	{8'd4,8'd176} : s = 180;
	{8'd4,8'd177} : s = 181;
	{8'd4,8'd178} : s = 182;
	{8'd4,8'd179} : s = 183;
	{8'd4,8'd180} : s = 184;
	{8'd4,8'd181} : s = 185;
	{8'd4,8'd182} : s = 186;
	{8'd4,8'd183} : s = 187;
	{8'd4,8'd184} : s = 188;
	{8'd4,8'd185} : s = 189;
	{8'd4,8'd186} : s = 190;
	{8'd4,8'd187} : s = 191;
	{8'd4,8'd188} : s = 192;
	{8'd4,8'd189} : s = 193;
	{8'd4,8'd190} : s = 194;
	{8'd4,8'd191} : s = 195;
	{8'd4,8'd192} : s = 196;
	{8'd4,8'd193} : s = 197;
	{8'd4,8'd194} : s = 198;
	{8'd4,8'd195} : s = 199;
	{8'd4,8'd196} : s = 200;
	{8'd4,8'd197} : s = 201;
	{8'd4,8'd198} : s = 202;
	{8'd4,8'd199} : s = 203;
	{8'd4,8'd200} : s = 204;
	{8'd4,8'd201} : s = 205;
	{8'd4,8'd202} : s = 206;
	{8'd4,8'd203} : s = 207;
	{8'd4,8'd204} : s = 208;
	{8'd4,8'd205} : s = 209;
	{8'd4,8'd206} : s = 210;
	{8'd4,8'd207} : s = 211;
	{8'd4,8'd208} : s = 212;
	{8'd4,8'd209} : s = 213;
	{8'd4,8'd210} : s = 214;
	{8'd4,8'd211} : s = 215;
	{8'd4,8'd212} : s = 216;
	{8'd4,8'd213} : s = 217;
	{8'd4,8'd214} : s = 218;
	{8'd4,8'd215} : s = 219;
	{8'd4,8'd216} : s = 220;
	{8'd4,8'd217} : s = 221;
	{8'd4,8'd218} : s = 222;
	{8'd4,8'd219} : s = 223;
	{8'd4,8'd220} : s = 224;
	{8'd4,8'd221} : s = 225;
	{8'd4,8'd222} : s = 226;
	{8'd4,8'd223} : s = 227;
	{8'd4,8'd224} : s = 228;
	{8'd4,8'd225} : s = 229;
	{8'd4,8'd226} : s = 230;
	{8'd4,8'd227} : s = 231;
	{8'd4,8'd228} : s = 232;
	{8'd4,8'd229} : s = 233;
	{8'd4,8'd230} : s = 234;
	{8'd4,8'd231} : s = 235;
	{8'd4,8'd232} : s = 236;
	{8'd4,8'd233} : s = 237;
	{8'd4,8'd234} : s = 238;
	{8'd4,8'd235} : s = 239;
	{8'd4,8'd236} : s = 240;
	{8'd4,8'd237} : s = 241;
	{8'd4,8'd238} : s = 242;
	{8'd4,8'd239} : s = 243;
	{8'd4,8'd240} : s = 244;
	{8'd4,8'd241} : s = 245;
	{8'd4,8'd242} : s = 246;
	{8'd4,8'd243} : s = 247;
	{8'd4,8'd244} : s = 248;
	{8'd4,8'd245} : s = 249;
	{8'd4,8'd246} : s = 250;
	{8'd4,8'd247} : s = 251;
	{8'd4,8'd248} : s = 252;
	{8'd4,8'd249} : s = 253;
	{8'd4,8'd250} : s = 254;
	{8'd4,8'd251} : s = 255;
	{8'd4,8'd252} : s = 256;
	{8'd4,8'd253} : s = 257;
	{8'd4,8'd254} : s = 258;
	{8'd4,8'd255} : s = 259;
	{8'd5,8'd0} : s = 5;
	{8'd5,8'd1} : s = 6;
	{8'd5,8'd2} : s = 7;
	{8'd5,8'd3} : s = 8;
	{8'd5,8'd4} : s = 9;
	{8'd5,8'd5} : s = 10;
	{8'd5,8'd6} : s = 11;
	{8'd5,8'd7} : s = 12;
	{8'd5,8'd8} : s = 13;
	{8'd5,8'd9} : s = 14;
	{8'd5,8'd10} : s = 15;
	{8'd5,8'd11} : s = 16;
	{8'd5,8'd12} : s = 17;
	{8'd5,8'd13} : s = 18;
	{8'd5,8'd14} : s = 19;
	{8'd5,8'd15} : s = 20;
	{8'd5,8'd16} : s = 21;
	{8'd5,8'd17} : s = 22;
	{8'd5,8'd18} : s = 23;
	{8'd5,8'd19} : s = 24;
	{8'd5,8'd20} : s = 25;
	{8'd5,8'd21} : s = 26;
	{8'd5,8'd22} : s = 27;
	{8'd5,8'd23} : s = 28;
	{8'd5,8'd24} : s = 29;
	{8'd5,8'd25} : s = 30;
	{8'd5,8'd26} : s = 31;
	{8'd5,8'd27} : s = 32;
	{8'd5,8'd28} : s = 33;
	{8'd5,8'd29} : s = 34;
	{8'd5,8'd30} : s = 35;
	{8'd5,8'd31} : s = 36;
	{8'd5,8'd32} : s = 37;
	{8'd5,8'd33} : s = 38;
	{8'd5,8'd34} : s = 39;
	{8'd5,8'd35} : s = 40;
	{8'd5,8'd36} : s = 41;
	{8'd5,8'd37} : s = 42;
	{8'd5,8'd38} : s = 43;
	{8'd5,8'd39} : s = 44;
	{8'd5,8'd40} : s = 45;
	{8'd5,8'd41} : s = 46;
	{8'd5,8'd42} : s = 47;
	{8'd5,8'd43} : s = 48;
	{8'd5,8'd44} : s = 49;
	{8'd5,8'd45} : s = 50;
	{8'd5,8'd46} : s = 51;
	{8'd5,8'd47} : s = 52;
	{8'd5,8'd48} : s = 53;
	{8'd5,8'd49} : s = 54;
	{8'd5,8'd50} : s = 55;
	{8'd5,8'd51} : s = 56;
	{8'd5,8'd52} : s = 57;
	{8'd5,8'd53} : s = 58;
	{8'd5,8'd54} : s = 59;
	{8'd5,8'd55} : s = 60;
	{8'd5,8'd56} : s = 61;
	{8'd5,8'd57} : s = 62;
	{8'd5,8'd58} : s = 63;
	{8'd5,8'd59} : s = 64;
	{8'd5,8'd60} : s = 65;
	{8'd5,8'd61} : s = 66;
	{8'd5,8'd62} : s = 67;
	{8'd5,8'd63} : s = 68;
	{8'd5,8'd64} : s = 69;
	{8'd5,8'd65} : s = 70;
	{8'd5,8'd66} : s = 71;
	{8'd5,8'd67} : s = 72;
	{8'd5,8'd68} : s = 73;
	{8'd5,8'd69} : s = 74;
	{8'd5,8'd70} : s = 75;
	{8'd5,8'd71} : s = 76;
	{8'd5,8'd72} : s = 77;
	{8'd5,8'd73} : s = 78;
	{8'd5,8'd74} : s = 79;
	{8'd5,8'd75} : s = 80;
	{8'd5,8'd76} : s = 81;
	{8'd5,8'd77} : s = 82;
	{8'd5,8'd78} : s = 83;
	{8'd5,8'd79} : s = 84;
	{8'd5,8'd80} : s = 85;
	{8'd5,8'd81} : s = 86;
	{8'd5,8'd82} : s = 87;
	{8'd5,8'd83} : s = 88;
	{8'd5,8'd84} : s = 89;
	{8'd5,8'd85} : s = 90;
	{8'd5,8'd86} : s = 91;
	{8'd5,8'd87} : s = 92;
	{8'd5,8'd88} : s = 93;
	{8'd5,8'd89} : s = 94;
	{8'd5,8'd90} : s = 95;
	{8'd5,8'd91} : s = 96;
	{8'd5,8'd92} : s = 97;
	{8'd5,8'd93} : s = 98;
	{8'd5,8'd94} : s = 99;
	{8'd5,8'd95} : s = 100;
	{8'd5,8'd96} : s = 101;
	{8'd5,8'd97} : s = 102;
	{8'd5,8'd98} : s = 103;
	{8'd5,8'd99} : s = 104;
	{8'd5,8'd100} : s = 105;
	{8'd5,8'd101} : s = 106;
	{8'd5,8'd102} : s = 107;
	{8'd5,8'd103} : s = 108;
	{8'd5,8'd104} : s = 109;
	{8'd5,8'd105} : s = 110;
	{8'd5,8'd106} : s = 111;
	{8'd5,8'd107} : s = 112;
	{8'd5,8'd108} : s = 113;
	{8'd5,8'd109} : s = 114;
	{8'd5,8'd110} : s = 115;
	{8'd5,8'd111} : s = 116;
	{8'd5,8'd112} : s = 117;
	{8'd5,8'd113} : s = 118;
	{8'd5,8'd114} : s = 119;
	{8'd5,8'd115} : s = 120;
	{8'd5,8'd116} : s = 121;
	{8'd5,8'd117} : s = 122;
	{8'd5,8'd118} : s = 123;
	{8'd5,8'd119} : s = 124;
	{8'd5,8'd120} : s = 125;
	{8'd5,8'd121} : s = 126;
	{8'd5,8'd122} : s = 127;
	{8'd5,8'd123} : s = 128;
	{8'd5,8'd124} : s = 129;
	{8'd5,8'd125} : s = 130;
	{8'd5,8'd126} : s = 131;
	{8'd5,8'd127} : s = 132;
	{8'd5,8'd128} : s = 133;
	{8'd5,8'd129} : s = 134;
	{8'd5,8'd130} : s = 135;
	{8'd5,8'd131} : s = 136;
	{8'd5,8'd132} : s = 137;
	{8'd5,8'd133} : s = 138;
	{8'd5,8'd134} : s = 139;
	{8'd5,8'd135} : s = 140;
	{8'd5,8'd136} : s = 141;
	{8'd5,8'd137} : s = 142;
	{8'd5,8'd138} : s = 143;
	{8'd5,8'd139} : s = 144;
	{8'd5,8'd140} : s = 145;
	{8'd5,8'd141} : s = 146;
	{8'd5,8'd142} : s = 147;
	{8'd5,8'd143} : s = 148;
	{8'd5,8'd144} : s = 149;
	{8'd5,8'd145} : s = 150;
	{8'd5,8'd146} : s = 151;
	{8'd5,8'd147} : s = 152;
	{8'd5,8'd148} : s = 153;
	{8'd5,8'd149} : s = 154;
	{8'd5,8'd150} : s = 155;
	{8'd5,8'd151} : s = 156;
	{8'd5,8'd152} : s = 157;
	{8'd5,8'd153} : s = 158;
	{8'd5,8'd154} : s = 159;
	{8'd5,8'd155} : s = 160;
	{8'd5,8'd156} : s = 161;
	{8'd5,8'd157} : s = 162;
	{8'd5,8'd158} : s = 163;
	{8'd5,8'd159} : s = 164;
	{8'd5,8'd160} : s = 165;
	{8'd5,8'd161} : s = 166;
	{8'd5,8'd162} : s = 167;
	{8'd5,8'd163} : s = 168;
	{8'd5,8'd164} : s = 169;
	{8'd5,8'd165} : s = 170;
	{8'd5,8'd166} : s = 171;
	{8'd5,8'd167} : s = 172;
	{8'd5,8'd168} : s = 173;
	{8'd5,8'd169} : s = 174;
	{8'd5,8'd170} : s = 175;
	{8'd5,8'd171} : s = 176;
	{8'd5,8'd172} : s = 177;
	{8'd5,8'd173} : s = 178;
	{8'd5,8'd174} : s = 179;
	{8'd5,8'd175} : s = 180;
	{8'd5,8'd176} : s = 181;
	{8'd5,8'd177} : s = 182;
	{8'd5,8'd178} : s = 183;
	{8'd5,8'd179} : s = 184;
	{8'd5,8'd180} : s = 185;
	{8'd5,8'd181} : s = 186;
	{8'd5,8'd182} : s = 187;
	{8'd5,8'd183} : s = 188;
	{8'd5,8'd184} : s = 189;
	{8'd5,8'd185} : s = 190;
	{8'd5,8'd186} : s = 191;
	{8'd5,8'd187} : s = 192;
	{8'd5,8'd188} : s = 193;
	{8'd5,8'd189} : s = 194;
	{8'd5,8'd190} : s = 195;
	{8'd5,8'd191} : s = 196;
	{8'd5,8'd192} : s = 197;
	{8'd5,8'd193} : s = 198;
	{8'd5,8'd194} : s = 199;
	{8'd5,8'd195} : s = 200;
	{8'd5,8'd196} : s = 201;
	{8'd5,8'd197} : s = 202;
	{8'd5,8'd198} : s = 203;
	{8'd5,8'd199} : s = 204;
	{8'd5,8'd200} : s = 205;
	{8'd5,8'd201} : s = 206;
	{8'd5,8'd202} : s = 207;
	{8'd5,8'd203} : s = 208;
	{8'd5,8'd204} : s = 209;
	{8'd5,8'd205} : s = 210;
	{8'd5,8'd206} : s = 211;
	{8'd5,8'd207} : s = 212;
	{8'd5,8'd208} : s = 213;
	{8'd5,8'd209} : s = 214;
	{8'd5,8'd210} : s = 215;
	{8'd5,8'd211} : s = 216;
	{8'd5,8'd212} : s = 217;
	{8'd5,8'd213} : s = 218;
	{8'd5,8'd214} : s = 219;
	{8'd5,8'd215} : s = 220;
	{8'd5,8'd216} : s = 221;
	{8'd5,8'd217} : s = 222;
	{8'd5,8'd218} : s = 223;
	{8'd5,8'd219} : s = 224;
	{8'd5,8'd220} : s = 225;
	{8'd5,8'd221} : s = 226;
	{8'd5,8'd222} : s = 227;
	{8'd5,8'd223} : s = 228;
	{8'd5,8'd224} : s = 229;
	{8'd5,8'd225} : s = 230;
	{8'd5,8'd226} : s = 231;
	{8'd5,8'd227} : s = 232;
	{8'd5,8'd228} : s = 233;
	{8'd5,8'd229} : s = 234;
	{8'd5,8'd230} : s = 235;
	{8'd5,8'd231} : s = 236;
	{8'd5,8'd232} : s = 237;
	{8'd5,8'd233} : s = 238;
	{8'd5,8'd234} : s = 239;
	{8'd5,8'd235} : s = 240;
	{8'd5,8'd236} : s = 241;
	{8'd5,8'd237} : s = 242;
	{8'd5,8'd238} : s = 243;
	{8'd5,8'd239} : s = 244;
	{8'd5,8'd240} : s = 245;
	{8'd5,8'd241} : s = 246;
	{8'd5,8'd242} : s = 247;
	{8'd5,8'd243} : s = 248;
	{8'd5,8'd244} : s = 249;
	{8'd5,8'd245} : s = 250;
	{8'd5,8'd246} : s = 251;
	{8'd5,8'd247} : s = 252;
	{8'd5,8'd248} : s = 253;
	{8'd5,8'd249} : s = 254;
	{8'd5,8'd250} : s = 255;
	{8'd5,8'd251} : s = 256;
	{8'd5,8'd252} : s = 257;
	{8'd5,8'd253} : s = 258;
	{8'd5,8'd254} : s = 259;
	{8'd5,8'd255} : s = 260;
	{8'd6,8'd0} : s = 6;
	{8'd6,8'd1} : s = 7;
	{8'd6,8'd2} : s = 8;
	{8'd6,8'd3} : s = 9;
	{8'd6,8'd4} : s = 10;
	{8'd6,8'd5} : s = 11;
	{8'd6,8'd6} : s = 12;
	{8'd6,8'd7} : s = 13;
	{8'd6,8'd8} : s = 14;
	{8'd6,8'd9} : s = 15;
	{8'd6,8'd10} : s = 16;
	{8'd6,8'd11} : s = 17;
	{8'd6,8'd12} : s = 18;
	{8'd6,8'd13} : s = 19;
	{8'd6,8'd14} : s = 20;
	{8'd6,8'd15} : s = 21;
	{8'd6,8'd16} : s = 22;
	{8'd6,8'd17} : s = 23;
	{8'd6,8'd18} : s = 24;
	{8'd6,8'd19} : s = 25;
	{8'd6,8'd20} : s = 26;
	{8'd6,8'd21} : s = 27;
	{8'd6,8'd22} : s = 28;
	{8'd6,8'd23} : s = 29;
	{8'd6,8'd24} : s = 30;
	{8'd6,8'd25} : s = 31;
	{8'd6,8'd26} : s = 32;
	{8'd6,8'd27} : s = 33;
	{8'd6,8'd28} : s = 34;
	{8'd6,8'd29} : s = 35;
	{8'd6,8'd30} : s = 36;
	{8'd6,8'd31} : s = 37;
	{8'd6,8'd32} : s = 38;
	{8'd6,8'd33} : s = 39;
	{8'd6,8'd34} : s = 40;
	{8'd6,8'd35} : s = 41;
	{8'd6,8'd36} : s = 42;
	{8'd6,8'd37} : s = 43;
	{8'd6,8'd38} : s = 44;
	{8'd6,8'd39} : s = 45;
	{8'd6,8'd40} : s = 46;
	{8'd6,8'd41} : s = 47;
	{8'd6,8'd42} : s = 48;
	{8'd6,8'd43} : s = 49;
	{8'd6,8'd44} : s = 50;
	{8'd6,8'd45} : s = 51;
	{8'd6,8'd46} : s = 52;
	{8'd6,8'd47} : s = 53;
	{8'd6,8'd48} : s = 54;
	{8'd6,8'd49} : s = 55;
	{8'd6,8'd50} : s = 56;
	{8'd6,8'd51} : s = 57;
	{8'd6,8'd52} : s = 58;
	{8'd6,8'd53} : s = 59;
	{8'd6,8'd54} : s = 60;
	{8'd6,8'd55} : s = 61;
	{8'd6,8'd56} : s = 62;
	{8'd6,8'd57} : s = 63;
	{8'd6,8'd58} : s = 64;
	{8'd6,8'd59} : s = 65;
	{8'd6,8'd60} : s = 66;
	{8'd6,8'd61} : s = 67;
	{8'd6,8'd62} : s = 68;
	{8'd6,8'd63} : s = 69;
	{8'd6,8'd64} : s = 70;
	{8'd6,8'd65} : s = 71;
	{8'd6,8'd66} : s = 72;
	{8'd6,8'd67} : s = 73;
	{8'd6,8'd68} : s = 74;
	{8'd6,8'd69} : s = 75;
	{8'd6,8'd70} : s = 76;
	{8'd6,8'd71} : s = 77;
	{8'd6,8'd72} : s = 78;
	{8'd6,8'd73} : s = 79;
	{8'd6,8'd74} : s = 80;
	{8'd6,8'd75} : s = 81;
	{8'd6,8'd76} : s = 82;
	{8'd6,8'd77} : s = 83;
	{8'd6,8'd78} : s = 84;
	{8'd6,8'd79} : s = 85;
	{8'd6,8'd80} : s = 86;
	{8'd6,8'd81} : s = 87;
	{8'd6,8'd82} : s = 88;
	{8'd6,8'd83} : s = 89;
	{8'd6,8'd84} : s = 90;
	{8'd6,8'd85} : s = 91;
	{8'd6,8'd86} : s = 92;
	{8'd6,8'd87} : s = 93;
	{8'd6,8'd88} : s = 94;
	{8'd6,8'd89} : s = 95;
	{8'd6,8'd90} : s = 96;
	{8'd6,8'd91} : s = 97;
	{8'd6,8'd92} : s = 98;
	{8'd6,8'd93} : s = 99;
	{8'd6,8'd94} : s = 100;
	{8'd6,8'd95} : s = 101;
	{8'd6,8'd96} : s = 102;
	{8'd6,8'd97} : s = 103;
	{8'd6,8'd98} : s = 104;
	{8'd6,8'd99} : s = 105;
	{8'd6,8'd100} : s = 106;
	{8'd6,8'd101} : s = 107;
	{8'd6,8'd102} : s = 108;
	{8'd6,8'd103} : s = 109;
	{8'd6,8'd104} : s = 110;
	{8'd6,8'd105} : s = 111;
	{8'd6,8'd106} : s = 112;
	{8'd6,8'd107} : s = 113;
	{8'd6,8'd108} : s = 114;
	{8'd6,8'd109} : s = 115;
	{8'd6,8'd110} : s = 116;
	{8'd6,8'd111} : s = 117;
	{8'd6,8'd112} : s = 118;
	{8'd6,8'd113} : s = 119;
	{8'd6,8'd114} : s = 120;
	{8'd6,8'd115} : s = 121;
	{8'd6,8'd116} : s = 122;
	{8'd6,8'd117} : s = 123;
	{8'd6,8'd118} : s = 124;
	{8'd6,8'd119} : s = 125;
	{8'd6,8'd120} : s = 126;
	{8'd6,8'd121} : s = 127;
	{8'd6,8'd122} : s = 128;
	{8'd6,8'd123} : s = 129;
	{8'd6,8'd124} : s = 130;
	{8'd6,8'd125} : s = 131;
	{8'd6,8'd126} : s = 132;
	{8'd6,8'd127} : s = 133;
	{8'd6,8'd128} : s = 134;
	{8'd6,8'd129} : s = 135;
	{8'd6,8'd130} : s = 136;
	{8'd6,8'd131} : s = 137;
	{8'd6,8'd132} : s = 138;
	{8'd6,8'd133} : s = 139;
	{8'd6,8'd134} : s = 140;
	{8'd6,8'd135} : s = 141;
	{8'd6,8'd136} : s = 142;
	{8'd6,8'd137} : s = 143;
	{8'd6,8'd138} : s = 144;
	{8'd6,8'd139} : s = 145;
	{8'd6,8'd140} : s = 146;
	{8'd6,8'd141} : s = 147;
	{8'd6,8'd142} : s = 148;
	{8'd6,8'd143} : s = 149;
	{8'd6,8'd144} : s = 150;
	{8'd6,8'd145} : s = 151;
	{8'd6,8'd146} : s = 152;
	{8'd6,8'd147} : s = 153;
	{8'd6,8'd148} : s = 154;
	{8'd6,8'd149} : s = 155;
	{8'd6,8'd150} : s = 156;
	{8'd6,8'd151} : s = 157;
	{8'd6,8'd152} : s = 158;
	{8'd6,8'd153} : s = 159;
	{8'd6,8'd154} : s = 160;
	{8'd6,8'd155} : s = 161;
	{8'd6,8'd156} : s = 162;
	{8'd6,8'd157} : s = 163;
	{8'd6,8'd158} : s = 164;
	{8'd6,8'd159} : s = 165;
	{8'd6,8'd160} : s = 166;
	{8'd6,8'd161} : s = 167;
	{8'd6,8'd162} : s = 168;
	{8'd6,8'd163} : s = 169;
	{8'd6,8'd164} : s = 170;
	{8'd6,8'd165} : s = 171;
	{8'd6,8'd166} : s = 172;
	{8'd6,8'd167} : s = 173;
	{8'd6,8'd168} : s = 174;
	{8'd6,8'd169} : s = 175;
	{8'd6,8'd170} : s = 176;
	{8'd6,8'd171} : s = 177;
	{8'd6,8'd172} : s = 178;
	{8'd6,8'd173} : s = 179;
	{8'd6,8'd174} : s = 180;
	{8'd6,8'd175} : s = 181;
	{8'd6,8'd176} : s = 182;
	{8'd6,8'd177} : s = 183;
	{8'd6,8'd178} : s = 184;
	{8'd6,8'd179} : s = 185;
	{8'd6,8'd180} : s = 186;
	{8'd6,8'd181} : s = 187;
	{8'd6,8'd182} : s = 188;
	{8'd6,8'd183} : s = 189;
	{8'd6,8'd184} : s = 190;
	{8'd6,8'd185} : s = 191;
	{8'd6,8'd186} : s = 192;
	{8'd6,8'd187} : s = 193;
	{8'd6,8'd188} : s = 194;
	{8'd6,8'd189} : s = 195;
	{8'd6,8'd190} : s = 196;
	{8'd6,8'd191} : s = 197;
	{8'd6,8'd192} : s = 198;
	{8'd6,8'd193} : s = 199;
	{8'd6,8'd194} : s = 200;
	{8'd6,8'd195} : s = 201;
	{8'd6,8'd196} : s = 202;
	{8'd6,8'd197} : s = 203;
	{8'd6,8'd198} : s = 204;
	{8'd6,8'd199} : s = 205;
	{8'd6,8'd200} : s = 206;
	{8'd6,8'd201} : s = 207;
	{8'd6,8'd202} : s = 208;
	{8'd6,8'd203} : s = 209;
	{8'd6,8'd204} : s = 210;
	{8'd6,8'd205} : s = 211;
	{8'd6,8'd206} : s = 212;
	{8'd6,8'd207} : s = 213;
	{8'd6,8'd208} : s = 214;
	{8'd6,8'd209} : s = 215;
	{8'd6,8'd210} : s = 216;
	{8'd6,8'd211} : s = 217;
	{8'd6,8'd212} : s = 218;
	{8'd6,8'd213} : s = 219;
	{8'd6,8'd214} : s = 220;
	{8'd6,8'd215} : s = 221;
	{8'd6,8'd216} : s = 222;
	{8'd6,8'd217} : s = 223;
	{8'd6,8'd218} : s = 224;
	{8'd6,8'd219} : s = 225;
	{8'd6,8'd220} : s = 226;
	{8'd6,8'd221} : s = 227;
	{8'd6,8'd222} : s = 228;
	{8'd6,8'd223} : s = 229;
	{8'd6,8'd224} : s = 230;
	{8'd6,8'd225} : s = 231;
	{8'd6,8'd226} : s = 232;
	{8'd6,8'd227} : s = 233;
	{8'd6,8'd228} : s = 234;
	{8'd6,8'd229} : s = 235;
	{8'd6,8'd230} : s = 236;
	{8'd6,8'd231} : s = 237;
	{8'd6,8'd232} : s = 238;
	{8'd6,8'd233} : s = 239;
	{8'd6,8'd234} : s = 240;
	{8'd6,8'd235} : s = 241;
	{8'd6,8'd236} : s = 242;
	{8'd6,8'd237} : s = 243;
	{8'd6,8'd238} : s = 244;
	{8'd6,8'd239} : s = 245;
	{8'd6,8'd240} : s = 246;
	{8'd6,8'd241} : s = 247;
	{8'd6,8'd242} : s = 248;
	{8'd6,8'd243} : s = 249;
	{8'd6,8'd244} : s = 250;
	{8'd6,8'd245} : s = 251;
	{8'd6,8'd246} : s = 252;
	{8'd6,8'd247} : s = 253;
	{8'd6,8'd248} : s = 254;
	{8'd6,8'd249} : s = 255;
	{8'd6,8'd250} : s = 256;
	{8'd6,8'd251} : s = 257;
	{8'd6,8'd252} : s = 258;
	{8'd6,8'd253} : s = 259;
	{8'd6,8'd254} : s = 260;
	{8'd6,8'd255} : s = 261;
	{8'd7,8'd0} : s = 7;
	{8'd7,8'd1} : s = 8;
	{8'd7,8'd2} : s = 9;
	{8'd7,8'd3} : s = 10;
	{8'd7,8'd4} : s = 11;
	{8'd7,8'd5} : s = 12;
	{8'd7,8'd6} : s = 13;
	{8'd7,8'd7} : s = 14;
	{8'd7,8'd8} : s = 15;
	{8'd7,8'd9} : s = 16;
	{8'd7,8'd10} : s = 17;
	{8'd7,8'd11} : s = 18;
	{8'd7,8'd12} : s = 19;
	{8'd7,8'd13} : s = 20;
	{8'd7,8'd14} : s = 21;
	{8'd7,8'd15} : s = 22;
	{8'd7,8'd16} : s = 23;
	{8'd7,8'd17} : s = 24;
	{8'd7,8'd18} : s = 25;
	{8'd7,8'd19} : s = 26;
	{8'd7,8'd20} : s = 27;
	{8'd7,8'd21} : s = 28;
	{8'd7,8'd22} : s = 29;
	{8'd7,8'd23} : s = 30;
	{8'd7,8'd24} : s = 31;
	{8'd7,8'd25} : s = 32;
	{8'd7,8'd26} : s = 33;
	{8'd7,8'd27} : s = 34;
	{8'd7,8'd28} : s = 35;
	{8'd7,8'd29} : s = 36;
	{8'd7,8'd30} : s = 37;
	{8'd7,8'd31} : s = 38;
	{8'd7,8'd32} : s = 39;
	{8'd7,8'd33} : s = 40;
	{8'd7,8'd34} : s = 41;
	{8'd7,8'd35} : s = 42;
	{8'd7,8'd36} : s = 43;
	{8'd7,8'd37} : s = 44;
	{8'd7,8'd38} : s = 45;
	{8'd7,8'd39} : s = 46;
	{8'd7,8'd40} : s = 47;
	{8'd7,8'd41} : s = 48;
	{8'd7,8'd42} : s = 49;
	{8'd7,8'd43} : s = 50;
	{8'd7,8'd44} : s = 51;
	{8'd7,8'd45} : s = 52;
	{8'd7,8'd46} : s = 53;
	{8'd7,8'd47} : s = 54;
	{8'd7,8'd48} : s = 55;
	{8'd7,8'd49} : s = 56;
	{8'd7,8'd50} : s = 57;
	{8'd7,8'd51} : s = 58;
	{8'd7,8'd52} : s = 59;
	{8'd7,8'd53} : s = 60;
	{8'd7,8'd54} : s = 61;
	{8'd7,8'd55} : s = 62;
	{8'd7,8'd56} : s = 63;
	{8'd7,8'd57} : s = 64;
	{8'd7,8'd58} : s = 65;
	{8'd7,8'd59} : s = 66;
	{8'd7,8'd60} : s = 67;
	{8'd7,8'd61} : s = 68;
	{8'd7,8'd62} : s = 69;
	{8'd7,8'd63} : s = 70;
	{8'd7,8'd64} : s = 71;
	{8'd7,8'd65} : s = 72;
	{8'd7,8'd66} : s = 73;
	{8'd7,8'd67} : s = 74;
	{8'd7,8'd68} : s = 75;
	{8'd7,8'd69} : s = 76;
	{8'd7,8'd70} : s = 77;
	{8'd7,8'd71} : s = 78;
	{8'd7,8'd72} : s = 79;
	{8'd7,8'd73} : s = 80;
	{8'd7,8'd74} : s = 81;
	{8'd7,8'd75} : s = 82;
	{8'd7,8'd76} : s = 83;
	{8'd7,8'd77} : s = 84;
	{8'd7,8'd78} : s = 85;
	{8'd7,8'd79} : s = 86;
	{8'd7,8'd80} : s = 87;
	{8'd7,8'd81} : s = 88;
	{8'd7,8'd82} : s = 89;
	{8'd7,8'd83} : s = 90;
	{8'd7,8'd84} : s = 91;
	{8'd7,8'd85} : s = 92;
	{8'd7,8'd86} : s = 93;
	{8'd7,8'd87} : s = 94;
	{8'd7,8'd88} : s = 95;
	{8'd7,8'd89} : s = 96;
	{8'd7,8'd90} : s = 97;
	{8'd7,8'd91} : s = 98;
	{8'd7,8'd92} : s = 99;
	{8'd7,8'd93} : s = 100;
	{8'd7,8'd94} : s = 101;
	{8'd7,8'd95} : s = 102;
	{8'd7,8'd96} : s = 103;
	{8'd7,8'd97} : s = 104;
	{8'd7,8'd98} : s = 105;
	{8'd7,8'd99} : s = 106;
	{8'd7,8'd100} : s = 107;
	{8'd7,8'd101} : s = 108;
	{8'd7,8'd102} : s = 109;
	{8'd7,8'd103} : s = 110;
	{8'd7,8'd104} : s = 111;
	{8'd7,8'd105} : s = 112;
	{8'd7,8'd106} : s = 113;
	{8'd7,8'd107} : s = 114;
	{8'd7,8'd108} : s = 115;
	{8'd7,8'd109} : s = 116;
	{8'd7,8'd110} : s = 117;
	{8'd7,8'd111} : s = 118;
	{8'd7,8'd112} : s = 119;
	{8'd7,8'd113} : s = 120;
	{8'd7,8'd114} : s = 121;
	{8'd7,8'd115} : s = 122;
	{8'd7,8'd116} : s = 123;
	{8'd7,8'd117} : s = 124;
	{8'd7,8'd118} : s = 125;
	{8'd7,8'd119} : s = 126;
	{8'd7,8'd120} : s = 127;
	{8'd7,8'd121} : s = 128;
	{8'd7,8'd122} : s = 129;
	{8'd7,8'd123} : s = 130;
	{8'd7,8'd124} : s = 131;
	{8'd7,8'd125} : s = 132;
	{8'd7,8'd126} : s = 133;
	{8'd7,8'd127} : s = 134;
	{8'd7,8'd128} : s = 135;
	{8'd7,8'd129} : s = 136;
	{8'd7,8'd130} : s = 137;
	{8'd7,8'd131} : s = 138;
	{8'd7,8'd132} : s = 139;
	{8'd7,8'd133} : s = 140;
	{8'd7,8'd134} : s = 141;
	{8'd7,8'd135} : s = 142;
	{8'd7,8'd136} : s = 143;
	{8'd7,8'd137} : s = 144;
	{8'd7,8'd138} : s = 145;
	{8'd7,8'd139} : s = 146;
	{8'd7,8'd140} : s = 147;
	{8'd7,8'd141} : s = 148;
	{8'd7,8'd142} : s = 149;
	{8'd7,8'd143} : s = 150;
	{8'd7,8'd144} : s = 151;
	{8'd7,8'd145} : s = 152;
	{8'd7,8'd146} : s = 153;
	{8'd7,8'd147} : s = 154;
	{8'd7,8'd148} : s = 155;
	{8'd7,8'd149} : s = 156;
	{8'd7,8'd150} : s = 157;
	{8'd7,8'd151} : s = 158;
	{8'd7,8'd152} : s = 159;
	{8'd7,8'd153} : s = 160;
	{8'd7,8'd154} : s = 161;
	{8'd7,8'd155} : s = 162;
	{8'd7,8'd156} : s = 163;
	{8'd7,8'd157} : s = 164;
	{8'd7,8'd158} : s = 165;
	{8'd7,8'd159} : s = 166;
	{8'd7,8'd160} : s = 167;
	{8'd7,8'd161} : s = 168;
	{8'd7,8'd162} : s = 169;
	{8'd7,8'd163} : s = 170;
	{8'd7,8'd164} : s = 171;
	{8'd7,8'd165} : s = 172;
	{8'd7,8'd166} : s = 173;
	{8'd7,8'd167} : s = 174;
	{8'd7,8'd168} : s = 175;
	{8'd7,8'd169} : s = 176;
	{8'd7,8'd170} : s = 177;
	{8'd7,8'd171} : s = 178;
	{8'd7,8'd172} : s = 179;
	{8'd7,8'd173} : s = 180;
	{8'd7,8'd174} : s = 181;
	{8'd7,8'd175} : s = 182;
	{8'd7,8'd176} : s = 183;
	{8'd7,8'd177} : s = 184;
	{8'd7,8'd178} : s = 185;
	{8'd7,8'd179} : s = 186;
	{8'd7,8'd180} : s = 187;
	{8'd7,8'd181} : s = 188;
	{8'd7,8'd182} : s = 189;
	{8'd7,8'd183} : s = 190;
	{8'd7,8'd184} : s = 191;
	{8'd7,8'd185} : s = 192;
	{8'd7,8'd186} : s = 193;
	{8'd7,8'd187} : s = 194;
	{8'd7,8'd188} : s = 195;
	{8'd7,8'd189} : s = 196;
	{8'd7,8'd190} : s = 197;
	{8'd7,8'd191} : s = 198;
	{8'd7,8'd192} : s = 199;
	{8'd7,8'd193} : s = 200;
	{8'd7,8'd194} : s = 201;
	{8'd7,8'd195} : s = 202;
	{8'd7,8'd196} : s = 203;
	{8'd7,8'd197} : s = 204;
	{8'd7,8'd198} : s = 205;
	{8'd7,8'd199} : s = 206;
	{8'd7,8'd200} : s = 207;
	{8'd7,8'd201} : s = 208;
	{8'd7,8'd202} : s = 209;
	{8'd7,8'd203} : s = 210;
	{8'd7,8'd204} : s = 211;
	{8'd7,8'd205} : s = 212;
	{8'd7,8'd206} : s = 213;
	{8'd7,8'd207} : s = 214;
	{8'd7,8'd208} : s = 215;
	{8'd7,8'd209} : s = 216;
	{8'd7,8'd210} : s = 217;
	{8'd7,8'd211} : s = 218;
	{8'd7,8'd212} : s = 219;
	{8'd7,8'd213} : s = 220;
	{8'd7,8'd214} : s = 221;
	{8'd7,8'd215} : s = 222;
	{8'd7,8'd216} : s = 223;
	{8'd7,8'd217} : s = 224;
	{8'd7,8'd218} : s = 225;
	{8'd7,8'd219} : s = 226;
	{8'd7,8'd220} : s = 227;
	{8'd7,8'd221} : s = 228;
	{8'd7,8'd222} : s = 229;
	{8'd7,8'd223} : s = 230;
	{8'd7,8'd224} : s = 231;
	{8'd7,8'd225} : s = 232;
	{8'd7,8'd226} : s = 233;
	{8'd7,8'd227} : s = 234;
	{8'd7,8'd228} : s = 235;
	{8'd7,8'd229} : s = 236;
	{8'd7,8'd230} : s = 237;
	{8'd7,8'd231} : s = 238;
	{8'd7,8'd232} : s = 239;
	{8'd7,8'd233} : s = 240;
	{8'd7,8'd234} : s = 241;
	{8'd7,8'd235} : s = 242;
	{8'd7,8'd236} : s = 243;
	{8'd7,8'd237} : s = 244;
	{8'd7,8'd238} : s = 245;
	{8'd7,8'd239} : s = 246;
	{8'd7,8'd240} : s = 247;
	{8'd7,8'd241} : s = 248;
	{8'd7,8'd242} : s = 249;
	{8'd7,8'd243} : s = 250;
	{8'd7,8'd244} : s = 251;
	{8'd7,8'd245} : s = 252;
	{8'd7,8'd246} : s = 253;
	{8'd7,8'd247} : s = 254;
	{8'd7,8'd248} : s = 255;
	{8'd7,8'd249} : s = 256;
	{8'd7,8'd250} : s = 257;
	{8'd7,8'd251} : s = 258;
	{8'd7,8'd252} : s = 259;
	{8'd7,8'd253} : s = 260;
	{8'd7,8'd254} : s = 261;
	{8'd7,8'd255} : s = 262;
	{8'd8,8'd0} : s = 8;
	{8'd8,8'd1} : s = 9;
	{8'd8,8'd2} : s = 10;
	{8'd8,8'd3} : s = 11;
	{8'd8,8'd4} : s = 12;
	{8'd8,8'd5} : s = 13;
	{8'd8,8'd6} : s = 14;
	{8'd8,8'd7} : s = 15;
	{8'd8,8'd8} : s = 16;
	{8'd8,8'd9} : s = 17;
	{8'd8,8'd10} : s = 18;
	{8'd8,8'd11} : s = 19;
	{8'd8,8'd12} : s = 20;
	{8'd8,8'd13} : s = 21;
	{8'd8,8'd14} : s = 22;
	{8'd8,8'd15} : s = 23;
	{8'd8,8'd16} : s = 24;
	{8'd8,8'd17} : s = 25;
	{8'd8,8'd18} : s = 26;
	{8'd8,8'd19} : s = 27;
	{8'd8,8'd20} : s = 28;
	{8'd8,8'd21} : s = 29;
	{8'd8,8'd22} : s = 30;
	{8'd8,8'd23} : s = 31;
	{8'd8,8'd24} : s = 32;
	{8'd8,8'd25} : s = 33;
	{8'd8,8'd26} : s = 34;
	{8'd8,8'd27} : s = 35;
	{8'd8,8'd28} : s = 36;
	{8'd8,8'd29} : s = 37;
	{8'd8,8'd30} : s = 38;
	{8'd8,8'd31} : s = 39;
	{8'd8,8'd32} : s = 40;
	{8'd8,8'd33} : s = 41;
	{8'd8,8'd34} : s = 42;
	{8'd8,8'd35} : s = 43;
	{8'd8,8'd36} : s = 44;
	{8'd8,8'd37} : s = 45;
	{8'd8,8'd38} : s = 46;
	{8'd8,8'd39} : s = 47;
	{8'd8,8'd40} : s = 48;
	{8'd8,8'd41} : s = 49;
	{8'd8,8'd42} : s = 50;
	{8'd8,8'd43} : s = 51;
	{8'd8,8'd44} : s = 52;
	{8'd8,8'd45} : s = 53;
	{8'd8,8'd46} : s = 54;
	{8'd8,8'd47} : s = 55;
	{8'd8,8'd48} : s = 56;
	{8'd8,8'd49} : s = 57;
	{8'd8,8'd50} : s = 58;
	{8'd8,8'd51} : s = 59;
	{8'd8,8'd52} : s = 60;
	{8'd8,8'd53} : s = 61;
	{8'd8,8'd54} : s = 62;
	{8'd8,8'd55} : s = 63;
	{8'd8,8'd56} : s = 64;
	{8'd8,8'd57} : s = 65;
	{8'd8,8'd58} : s = 66;
	{8'd8,8'd59} : s = 67;
	{8'd8,8'd60} : s = 68;
	{8'd8,8'd61} : s = 69;
	{8'd8,8'd62} : s = 70;
	{8'd8,8'd63} : s = 71;
	{8'd8,8'd64} : s = 72;
	{8'd8,8'd65} : s = 73;
	{8'd8,8'd66} : s = 74;
	{8'd8,8'd67} : s = 75;
	{8'd8,8'd68} : s = 76;
	{8'd8,8'd69} : s = 77;
	{8'd8,8'd70} : s = 78;
	{8'd8,8'd71} : s = 79;
	{8'd8,8'd72} : s = 80;
	{8'd8,8'd73} : s = 81;
	{8'd8,8'd74} : s = 82;
	{8'd8,8'd75} : s = 83;
	{8'd8,8'd76} : s = 84;
	{8'd8,8'd77} : s = 85;
	{8'd8,8'd78} : s = 86;
	{8'd8,8'd79} : s = 87;
	{8'd8,8'd80} : s = 88;
	{8'd8,8'd81} : s = 89;
	{8'd8,8'd82} : s = 90;
	{8'd8,8'd83} : s = 91;
	{8'd8,8'd84} : s = 92;
	{8'd8,8'd85} : s = 93;
	{8'd8,8'd86} : s = 94;
	{8'd8,8'd87} : s = 95;
	{8'd8,8'd88} : s = 96;
	{8'd8,8'd89} : s = 97;
	{8'd8,8'd90} : s = 98;
	{8'd8,8'd91} : s = 99;
	{8'd8,8'd92} : s = 100;
	{8'd8,8'd93} : s = 101;
	{8'd8,8'd94} : s = 102;
	{8'd8,8'd95} : s = 103;
	{8'd8,8'd96} : s = 104;
	{8'd8,8'd97} : s = 105;
	{8'd8,8'd98} : s = 106;
	{8'd8,8'd99} : s = 107;
	{8'd8,8'd100} : s = 108;
	{8'd8,8'd101} : s = 109;
	{8'd8,8'd102} : s = 110;
	{8'd8,8'd103} : s = 111;
	{8'd8,8'd104} : s = 112;
	{8'd8,8'd105} : s = 113;
	{8'd8,8'd106} : s = 114;
	{8'd8,8'd107} : s = 115;
	{8'd8,8'd108} : s = 116;
	{8'd8,8'd109} : s = 117;
	{8'd8,8'd110} : s = 118;
	{8'd8,8'd111} : s = 119;
	{8'd8,8'd112} : s = 120;
	{8'd8,8'd113} : s = 121;
	{8'd8,8'd114} : s = 122;
	{8'd8,8'd115} : s = 123;
	{8'd8,8'd116} : s = 124;
	{8'd8,8'd117} : s = 125;
	{8'd8,8'd118} : s = 126;
	{8'd8,8'd119} : s = 127;
	{8'd8,8'd120} : s = 128;
	{8'd8,8'd121} : s = 129;
	{8'd8,8'd122} : s = 130;
	{8'd8,8'd123} : s = 131;
	{8'd8,8'd124} : s = 132;
	{8'd8,8'd125} : s = 133;
	{8'd8,8'd126} : s = 134;
	{8'd8,8'd127} : s = 135;
	{8'd8,8'd128} : s = 136;
	{8'd8,8'd129} : s = 137;
	{8'd8,8'd130} : s = 138;
	{8'd8,8'd131} : s = 139;
	{8'd8,8'd132} : s = 140;
	{8'd8,8'd133} : s = 141;
	{8'd8,8'd134} : s = 142;
	{8'd8,8'd135} : s = 143;
	{8'd8,8'd136} : s = 144;
	{8'd8,8'd137} : s = 145;
	{8'd8,8'd138} : s = 146;
	{8'd8,8'd139} : s = 147;
	{8'd8,8'd140} : s = 148;
	{8'd8,8'd141} : s = 149;
	{8'd8,8'd142} : s = 150;
	{8'd8,8'd143} : s = 151;
	{8'd8,8'd144} : s = 152;
	{8'd8,8'd145} : s = 153;
	{8'd8,8'd146} : s = 154;
	{8'd8,8'd147} : s = 155;
	{8'd8,8'd148} : s = 156;
	{8'd8,8'd149} : s = 157;
	{8'd8,8'd150} : s = 158;
	{8'd8,8'd151} : s = 159;
	{8'd8,8'd152} : s = 160;
	{8'd8,8'd153} : s = 161;
	{8'd8,8'd154} : s = 162;
	{8'd8,8'd155} : s = 163;
	{8'd8,8'd156} : s = 164;
	{8'd8,8'd157} : s = 165;
	{8'd8,8'd158} : s = 166;
	{8'd8,8'd159} : s = 167;
	{8'd8,8'd160} : s = 168;
	{8'd8,8'd161} : s = 169;
	{8'd8,8'd162} : s = 170;
	{8'd8,8'd163} : s = 171;
	{8'd8,8'd164} : s = 172;
	{8'd8,8'd165} : s = 173;
	{8'd8,8'd166} : s = 174;
	{8'd8,8'd167} : s = 175;
	{8'd8,8'd168} : s = 176;
	{8'd8,8'd169} : s = 177;
	{8'd8,8'd170} : s = 178;
	{8'd8,8'd171} : s = 179;
	{8'd8,8'd172} : s = 180;
	{8'd8,8'd173} : s = 181;
	{8'd8,8'd174} : s = 182;
	{8'd8,8'd175} : s = 183;
	{8'd8,8'd176} : s = 184;
	{8'd8,8'd177} : s = 185;
	{8'd8,8'd178} : s = 186;
	{8'd8,8'd179} : s = 187;
	{8'd8,8'd180} : s = 188;
	{8'd8,8'd181} : s = 189;
	{8'd8,8'd182} : s = 190;
	{8'd8,8'd183} : s = 191;
	{8'd8,8'd184} : s = 192;
	{8'd8,8'd185} : s = 193;
	{8'd8,8'd186} : s = 194;
	{8'd8,8'd187} : s = 195;
	{8'd8,8'd188} : s = 196;
	{8'd8,8'd189} : s = 197;
	{8'd8,8'd190} : s = 198;
	{8'd8,8'd191} : s = 199;
	{8'd8,8'd192} : s = 200;
	{8'd8,8'd193} : s = 201;
	{8'd8,8'd194} : s = 202;
	{8'd8,8'd195} : s = 203;
	{8'd8,8'd196} : s = 204;
	{8'd8,8'd197} : s = 205;
	{8'd8,8'd198} : s = 206;
	{8'd8,8'd199} : s = 207;
	{8'd8,8'd200} : s = 208;
	{8'd8,8'd201} : s = 209;
	{8'd8,8'd202} : s = 210;
	{8'd8,8'd203} : s = 211;
	{8'd8,8'd204} : s = 212;
	{8'd8,8'd205} : s = 213;
	{8'd8,8'd206} : s = 214;
	{8'd8,8'd207} : s = 215;
	{8'd8,8'd208} : s = 216;
	{8'd8,8'd209} : s = 217;
	{8'd8,8'd210} : s = 218;
	{8'd8,8'd211} : s = 219;
	{8'd8,8'd212} : s = 220;
	{8'd8,8'd213} : s = 221;
	{8'd8,8'd214} : s = 222;
	{8'd8,8'd215} : s = 223;
	{8'd8,8'd216} : s = 224;
	{8'd8,8'd217} : s = 225;
	{8'd8,8'd218} : s = 226;
	{8'd8,8'd219} : s = 227;
	{8'd8,8'd220} : s = 228;
	{8'd8,8'd221} : s = 229;
	{8'd8,8'd222} : s = 230;
	{8'd8,8'd223} : s = 231;
	{8'd8,8'd224} : s = 232;
	{8'd8,8'd225} : s = 233;
	{8'd8,8'd226} : s = 234;
	{8'd8,8'd227} : s = 235;
	{8'd8,8'd228} : s = 236;
	{8'd8,8'd229} : s = 237;
	{8'd8,8'd230} : s = 238;
	{8'd8,8'd231} : s = 239;
	{8'd8,8'd232} : s = 240;
	{8'd8,8'd233} : s = 241;
	{8'd8,8'd234} : s = 242;
	{8'd8,8'd235} : s = 243;
	{8'd8,8'd236} : s = 244;
	{8'd8,8'd237} : s = 245;
	{8'd8,8'd238} : s = 246;
	{8'd8,8'd239} : s = 247;
	{8'd8,8'd240} : s = 248;
	{8'd8,8'd241} : s = 249;
	{8'd8,8'd242} : s = 250;
	{8'd8,8'd243} : s = 251;
	{8'd8,8'd244} : s = 252;
	{8'd8,8'd245} : s = 253;
	{8'd8,8'd246} : s = 254;
	{8'd8,8'd247} : s = 255;
	{8'd8,8'd248} : s = 256;
	{8'd8,8'd249} : s = 257;
	{8'd8,8'd250} : s = 258;
	{8'd8,8'd251} : s = 259;
	{8'd8,8'd252} : s = 260;
	{8'd8,8'd253} : s = 261;
	{8'd8,8'd254} : s = 262;
	{8'd8,8'd255} : s = 263;
	{8'd9,8'd0} : s = 9;
	{8'd9,8'd1} : s = 10;
	{8'd9,8'd2} : s = 11;
	{8'd9,8'd3} : s = 12;
	{8'd9,8'd4} : s = 13;
	{8'd9,8'd5} : s = 14;
	{8'd9,8'd6} : s = 15;
	{8'd9,8'd7} : s = 16;
	{8'd9,8'd8} : s = 17;
	{8'd9,8'd9} : s = 18;
	{8'd9,8'd10} : s = 19;
	{8'd9,8'd11} : s = 20;
	{8'd9,8'd12} : s = 21;
	{8'd9,8'd13} : s = 22;
	{8'd9,8'd14} : s = 23;
	{8'd9,8'd15} : s = 24;
	{8'd9,8'd16} : s = 25;
	{8'd9,8'd17} : s = 26;
	{8'd9,8'd18} : s = 27;
	{8'd9,8'd19} : s = 28;
	{8'd9,8'd20} : s = 29;
	{8'd9,8'd21} : s = 30;
	{8'd9,8'd22} : s = 31;
	{8'd9,8'd23} : s = 32;
	{8'd9,8'd24} : s = 33;
	{8'd9,8'd25} : s = 34;
	{8'd9,8'd26} : s = 35;
	{8'd9,8'd27} : s = 36;
	{8'd9,8'd28} : s = 37;
	{8'd9,8'd29} : s = 38;
	{8'd9,8'd30} : s = 39;
	{8'd9,8'd31} : s = 40;
	{8'd9,8'd32} : s = 41;
	{8'd9,8'd33} : s = 42;
	{8'd9,8'd34} : s = 43;
	{8'd9,8'd35} : s = 44;
	{8'd9,8'd36} : s = 45;
	{8'd9,8'd37} : s = 46;
	{8'd9,8'd38} : s = 47;
	{8'd9,8'd39} : s = 48;
	{8'd9,8'd40} : s = 49;
	{8'd9,8'd41} : s = 50;
	{8'd9,8'd42} : s = 51;
	{8'd9,8'd43} : s = 52;
	{8'd9,8'd44} : s = 53;
	{8'd9,8'd45} : s = 54;
	{8'd9,8'd46} : s = 55;
	{8'd9,8'd47} : s = 56;
	{8'd9,8'd48} : s = 57;
	{8'd9,8'd49} : s = 58;
	{8'd9,8'd50} : s = 59;
	{8'd9,8'd51} : s = 60;
	{8'd9,8'd52} : s = 61;
	{8'd9,8'd53} : s = 62;
	{8'd9,8'd54} : s = 63;
	{8'd9,8'd55} : s = 64;
	{8'd9,8'd56} : s = 65;
	{8'd9,8'd57} : s = 66;
	{8'd9,8'd58} : s = 67;
	{8'd9,8'd59} : s = 68;
	{8'd9,8'd60} : s = 69;
	{8'd9,8'd61} : s = 70;
	{8'd9,8'd62} : s = 71;
	{8'd9,8'd63} : s = 72;
	{8'd9,8'd64} : s = 73;
	{8'd9,8'd65} : s = 74;
	{8'd9,8'd66} : s = 75;
	{8'd9,8'd67} : s = 76;
	{8'd9,8'd68} : s = 77;
	{8'd9,8'd69} : s = 78;
	{8'd9,8'd70} : s = 79;
	{8'd9,8'd71} : s = 80;
	{8'd9,8'd72} : s = 81;
	{8'd9,8'd73} : s = 82;
	{8'd9,8'd74} : s = 83;
	{8'd9,8'd75} : s = 84;
	{8'd9,8'd76} : s = 85;
	{8'd9,8'd77} : s = 86;
	{8'd9,8'd78} : s = 87;
	{8'd9,8'd79} : s = 88;
	{8'd9,8'd80} : s = 89;
	{8'd9,8'd81} : s = 90;
	{8'd9,8'd82} : s = 91;
	{8'd9,8'd83} : s = 92;
	{8'd9,8'd84} : s = 93;
	{8'd9,8'd85} : s = 94;
	{8'd9,8'd86} : s = 95;
	{8'd9,8'd87} : s = 96;
	{8'd9,8'd88} : s = 97;
	{8'd9,8'd89} : s = 98;
	{8'd9,8'd90} : s = 99;
	{8'd9,8'd91} : s = 100;
	{8'd9,8'd92} : s = 101;
	{8'd9,8'd93} : s = 102;
	{8'd9,8'd94} : s = 103;
	{8'd9,8'd95} : s = 104;
	{8'd9,8'd96} : s = 105;
	{8'd9,8'd97} : s = 106;
	{8'd9,8'd98} : s = 107;
	{8'd9,8'd99} : s = 108;
	{8'd9,8'd100} : s = 109;
	{8'd9,8'd101} : s = 110;
	{8'd9,8'd102} : s = 111;
	{8'd9,8'd103} : s = 112;
	{8'd9,8'd104} : s = 113;
	{8'd9,8'd105} : s = 114;
	{8'd9,8'd106} : s = 115;
	{8'd9,8'd107} : s = 116;
	{8'd9,8'd108} : s = 117;
	{8'd9,8'd109} : s = 118;
	{8'd9,8'd110} : s = 119;
	{8'd9,8'd111} : s = 120;
	{8'd9,8'd112} : s = 121;
	{8'd9,8'd113} : s = 122;
	{8'd9,8'd114} : s = 123;
	{8'd9,8'd115} : s = 124;
	{8'd9,8'd116} : s = 125;
	{8'd9,8'd117} : s = 126;
	{8'd9,8'd118} : s = 127;
	{8'd9,8'd119} : s = 128;
	{8'd9,8'd120} : s = 129;
	{8'd9,8'd121} : s = 130;
	{8'd9,8'd122} : s = 131;
	{8'd9,8'd123} : s = 132;
	{8'd9,8'd124} : s = 133;
	{8'd9,8'd125} : s = 134;
	{8'd9,8'd126} : s = 135;
	{8'd9,8'd127} : s = 136;
	{8'd9,8'd128} : s = 137;
	{8'd9,8'd129} : s = 138;
	{8'd9,8'd130} : s = 139;
	{8'd9,8'd131} : s = 140;
	{8'd9,8'd132} : s = 141;
	{8'd9,8'd133} : s = 142;
	{8'd9,8'd134} : s = 143;
	{8'd9,8'd135} : s = 144;
	{8'd9,8'd136} : s = 145;
	{8'd9,8'd137} : s = 146;
	{8'd9,8'd138} : s = 147;
	{8'd9,8'd139} : s = 148;
	{8'd9,8'd140} : s = 149;
	{8'd9,8'd141} : s = 150;
	{8'd9,8'd142} : s = 151;
	{8'd9,8'd143} : s = 152;
	{8'd9,8'd144} : s = 153;
	{8'd9,8'd145} : s = 154;
	{8'd9,8'd146} : s = 155;
	{8'd9,8'd147} : s = 156;
	{8'd9,8'd148} : s = 157;
	{8'd9,8'd149} : s = 158;
	{8'd9,8'd150} : s = 159;
	{8'd9,8'd151} : s = 160;
	{8'd9,8'd152} : s = 161;
	{8'd9,8'd153} : s = 162;
	{8'd9,8'd154} : s = 163;
	{8'd9,8'd155} : s = 164;
	{8'd9,8'd156} : s = 165;
	{8'd9,8'd157} : s = 166;
	{8'd9,8'd158} : s = 167;
	{8'd9,8'd159} : s = 168;
	{8'd9,8'd160} : s = 169;
	{8'd9,8'd161} : s = 170;
	{8'd9,8'd162} : s = 171;
	{8'd9,8'd163} : s = 172;
	{8'd9,8'd164} : s = 173;
	{8'd9,8'd165} : s = 174;
	{8'd9,8'd166} : s = 175;
	{8'd9,8'd167} : s = 176;
	{8'd9,8'd168} : s = 177;
	{8'd9,8'd169} : s = 178;
	{8'd9,8'd170} : s = 179;
	{8'd9,8'd171} : s = 180;
	{8'd9,8'd172} : s = 181;
	{8'd9,8'd173} : s = 182;
	{8'd9,8'd174} : s = 183;
	{8'd9,8'd175} : s = 184;
	{8'd9,8'd176} : s = 185;
	{8'd9,8'd177} : s = 186;
	{8'd9,8'd178} : s = 187;
	{8'd9,8'd179} : s = 188;
	{8'd9,8'd180} : s = 189;
	{8'd9,8'd181} : s = 190;
	{8'd9,8'd182} : s = 191;
	{8'd9,8'd183} : s = 192;
	{8'd9,8'd184} : s = 193;
	{8'd9,8'd185} : s = 194;
	{8'd9,8'd186} : s = 195;
	{8'd9,8'd187} : s = 196;
	{8'd9,8'd188} : s = 197;
	{8'd9,8'd189} : s = 198;
	{8'd9,8'd190} : s = 199;
	{8'd9,8'd191} : s = 200;
	{8'd9,8'd192} : s = 201;
	{8'd9,8'd193} : s = 202;
	{8'd9,8'd194} : s = 203;
	{8'd9,8'd195} : s = 204;
	{8'd9,8'd196} : s = 205;
	{8'd9,8'd197} : s = 206;
	{8'd9,8'd198} : s = 207;
	{8'd9,8'd199} : s = 208;
	{8'd9,8'd200} : s = 209;
	{8'd9,8'd201} : s = 210;
	{8'd9,8'd202} : s = 211;
	{8'd9,8'd203} : s = 212;
	{8'd9,8'd204} : s = 213;
	{8'd9,8'd205} : s = 214;
	{8'd9,8'd206} : s = 215;
	{8'd9,8'd207} : s = 216;
	{8'd9,8'd208} : s = 217;
	{8'd9,8'd209} : s = 218;
	{8'd9,8'd210} : s = 219;
	{8'd9,8'd211} : s = 220;
	{8'd9,8'd212} : s = 221;
	{8'd9,8'd213} : s = 222;
	{8'd9,8'd214} : s = 223;
	{8'd9,8'd215} : s = 224;
	{8'd9,8'd216} : s = 225;
	{8'd9,8'd217} : s = 226;
	{8'd9,8'd218} : s = 227;
	{8'd9,8'd219} : s = 228;
	{8'd9,8'd220} : s = 229;
	{8'd9,8'd221} : s = 230;
	{8'd9,8'd222} : s = 231;
	{8'd9,8'd223} : s = 232;
	{8'd9,8'd224} : s = 233;
	{8'd9,8'd225} : s = 234;
	{8'd9,8'd226} : s = 235;
	{8'd9,8'd227} : s = 236;
	{8'd9,8'd228} : s = 237;
	{8'd9,8'd229} : s = 238;
	{8'd9,8'd230} : s = 239;
	{8'd9,8'd231} : s = 240;
	{8'd9,8'd232} : s = 241;
	{8'd9,8'd233} : s = 242;
	{8'd9,8'd234} : s = 243;
	{8'd9,8'd235} : s = 244;
	{8'd9,8'd236} : s = 245;
	{8'd9,8'd237} : s = 246;
	{8'd9,8'd238} : s = 247;
	{8'd9,8'd239} : s = 248;
	{8'd9,8'd240} : s = 249;
	{8'd9,8'd241} : s = 250;
	{8'd9,8'd242} : s = 251;
	{8'd9,8'd243} : s = 252;
	{8'd9,8'd244} : s = 253;
	{8'd9,8'd245} : s = 254;
	{8'd9,8'd246} : s = 255;
	{8'd9,8'd247} : s = 256;
	{8'd9,8'd248} : s = 257;
	{8'd9,8'd249} : s = 258;
	{8'd9,8'd250} : s = 259;
	{8'd9,8'd251} : s = 260;
	{8'd9,8'd252} : s = 261;
	{8'd9,8'd253} : s = 262;
	{8'd9,8'd254} : s = 263;
	{8'd9,8'd255} : s = 264;
	{8'd10,8'd0} : s = 10;
	{8'd10,8'd1} : s = 11;
	{8'd10,8'd2} : s = 12;
	{8'd10,8'd3} : s = 13;
	{8'd10,8'd4} : s = 14;
	{8'd10,8'd5} : s = 15;
	{8'd10,8'd6} : s = 16;
	{8'd10,8'd7} : s = 17;
	{8'd10,8'd8} : s = 18;
	{8'd10,8'd9} : s = 19;
	{8'd10,8'd10} : s = 20;
	{8'd10,8'd11} : s = 21;
	{8'd10,8'd12} : s = 22;
	{8'd10,8'd13} : s = 23;
	{8'd10,8'd14} : s = 24;
	{8'd10,8'd15} : s = 25;
	{8'd10,8'd16} : s = 26;
	{8'd10,8'd17} : s = 27;
	{8'd10,8'd18} : s = 28;
	{8'd10,8'd19} : s = 29;
	{8'd10,8'd20} : s = 30;
	{8'd10,8'd21} : s = 31;
	{8'd10,8'd22} : s = 32;
	{8'd10,8'd23} : s = 33;
	{8'd10,8'd24} : s = 34;
	{8'd10,8'd25} : s = 35;
	{8'd10,8'd26} : s = 36;
	{8'd10,8'd27} : s = 37;
	{8'd10,8'd28} : s = 38;
	{8'd10,8'd29} : s = 39;
	{8'd10,8'd30} : s = 40;
	{8'd10,8'd31} : s = 41;
	{8'd10,8'd32} : s = 42;
	{8'd10,8'd33} : s = 43;
	{8'd10,8'd34} : s = 44;
	{8'd10,8'd35} : s = 45;
	{8'd10,8'd36} : s = 46;
	{8'd10,8'd37} : s = 47;
	{8'd10,8'd38} : s = 48;
	{8'd10,8'd39} : s = 49;
	{8'd10,8'd40} : s = 50;
	{8'd10,8'd41} : s = 51;
	{8'd10,8'd42} : s = 52;
	{8'd10,8'd43} : s = 53;
	{8'd10,8'd44} : s = 54;
	{8'd10,8'd45} : s = 55;
	{8'd10,8'd46} : s = 56;
	{8'd10,8'd47} : s = 57;
	{8'd10,8'd48} : s = 58;
	{8'd10,8'd49} : s = 59;
	{8'd10,8'd50} : s = 60;
	{8'd10,8'd51} : s = 61;
	{8'd10,8'd52} : s = 62;
	{8'd10,8'd53} : s = 63;
	{8'd10,8'd54} : s = 64;
	{8'd10,8'd55} : s = 65;
	{8'd10,8'd56} : s = 66;
	{8'd10,8'd57} : s = 67;
	{8'd10,8'd58} : s = 68;
	{8'd10,8'd59} : s = 69;
	{8'd10,8'd60} : s = 70;
	{8'd10,8'd61} : s = 71;
	{8'd10,8'd62} : s = 72;
	{8'd10,8'd63} : s = 73;
	{8'd10,8'd64} : s = 74;
	{8'd10,8'd65} : s = 75;
	{8'd10,8'd66} : s = 76;
	{8'd10,8'd67} : s = 77;
	{8'd10,8'd68} : s = 78;
	{8'd10,8'd69} : s = 79;
	{8'd10,8'd70} : s = 80;
	{8'd10,8'd71} : s = 81;
	{8'd10,8'd72} : s = 82;
	{8'd10,8'd73} : s = 83;
	{8'd10,8'd74} : s = 84;
	{8'd10,8'd75} : s = 85;
	{8'd10,8'd76} : s = 86;
	{8'd10,8'd77} : s = 87;
	{8'd10,8'd78} : s = 88;
	{8'd10,8'd79} : s = 89;
	{8'd10,8'd80} : s = 90;
	{8'd10,8'd81} : s = 91;
	{8'd10,8'd82} : s = 92;
	{8'd10,8'd83} : s = 93;
	{8'd10,8'd84} : s = 94;
	{8'd10,8'd85} : s = 95;
	{8'd10,8'd86} : s = 96;
	{8'd10,8'd87} : s = 97;
	{8'd10,8'd88} : s = 98;
	{8'd10,8'd89} : s = 99;
	{8'd10,8'd90} : s = 100;
	{8'd10,8'd91} : s = 101;
	{8'd10,8'd92} : s = 102;
	{8'd10,8'd93} : s = 103;
	{8'd10,8'd94} : s = 104;
	{8'd10,8'd95} : s = 105;
	{8'd10,8'd96} : s = 106;
	{8'd10,8'd97} : s = 107;
	{8'd10,8'd98} : s = 108;
	{8'd10,8'd99} : s = 109;
	{8'd10,8'd100} : s = 110;
	{8'd10,8'd101} : s = 111;
	{8'd10,8'd102} : s = 112;
	{8'd10,8'd103} : s = 113;
	{8'd10,8'd104} : s = 114;
	{8'd10,8'd105} : s = 115;
	{8'd10,8'd106} : s = 116;
	{8'd10,8'd107} : s = 117;
	{8'd10,8'd108} : s = 118;
	{8'd10,8'd109} : s = 119;
	{8'd10,8'd110} : s = 120;
	{8'd10,8'd111} : s = 121;
	{8'd10,8'd112} : s = 122;
	{8'd10,8'd113} : s = 123;
	{8'd10,8'd114} : s = 124;
	{8'd10,8'd115} : s = 125;
	{8'd10,8'd116} : s = 126;
	{8'd10,8'd117} : s = 127;
	{8'd10,8'd118} : s = 128;
	{8'd10,8'd119} : s = 129;
	{8'd10,8'd120} : s = 130;
	{8'd10,8'd121} : s = 131;
	{8'd10,8'd122} : s = 132;
	{8'd10,8'd123} : s = 133;
	{8'd10,8'd124} : s = 134;
	{8'd10,8'd125} : s = 135;
	{8'd10,8'd126} : s = 136;
	{8'd10,8'd127} : s = 137;
	{8'd10,8'd128} : s = 138;
	{8'd10,8'd129} : s = 139;
	{8'd10,8'd130} : s = 140;
	{8'd10,8'd131} : s = 141;
	{8'd10,8'd132} : s = 142;
	{8'd10,8'd133} : s = 143;
	{8'd10,8'd134} : s = 144;
	{8'd10,8'd135} : s = 145;
	{8'd10,8'd136} : s = 146;
	{8'd10,8'd137} : s = 147;
	{8'd10,8'd138} : s = 148;
	{8'd10,8'd139} : s = 149;
	{8'd10,8'd140} : s = 150;
	{8'd10,8'd141} : s = 151;
	{8'd10,8'd142} : s = 152;
	{8'd10,8'd143} : s = 153;
	{8'd10,8'd144} : s = 154;
	{8'd10,8'd145} : s = 155;
	{8'd10,8'd146} : s = 156;
	{8'd10,8'd147} : s = 157;
	{8'd10,8'd148} : s = 158;
	{8'd10,8'd149} : s = 159;
	{8'd10,8'd150} : s = 160;
	{8'd10,8'd151} : s = 161;
	{8'd10,8'd152} : s = 162;
	{8'd10,8'd153} : s = 163;
	{8'd10,8'd154} : s = 164;
	{8'd10,8'd155} : s = 165;
	{8'd10,8'd156} : s = 166;
	{8'd10,8'd157} : s = 167;
	{8'd10,8'd158} : s = 168;
	{8'd10,8'd159} : s = 169;
	{8'd10,8'd160} : s = 170;
	{8'd10,8'd161} : s = 171;
	{8'd10,8'd162} : s = 172;
	{8'd10,8'd163} : s = 173;
	{8'd10,8'd164} : s = 174;
	{8'd10,8'd165} : s = 175;
	{8'd10,8'd166} : s = 176;
	{8'd10,8'd167} : s = 177;
	{8'd10,8'd168} : s = 178;
	{8'd10,8'd169} : s = 179;
	{8'd10,8'd170} : s = 180;
	{8'd10,8'd171} : s = 181;
	{8'd10,8'd172} : s = 182;
	{8'd10,8'd173} : s = 183;
	{8'd10,8'd174} : s = 184;
	{8'd10,8'd175} : s = 185;
	{8'd10,8'd176} : s = 186;
	{8'd10,8'd177} : s = 187;
	{8'd10,8'd178} : s = 188;
	{8'd10,8'd179} : s = 189;
	{8'd10,8'd180} : s = 190;
	{8'd10,8'd181} : s = 191;
	{8'd10,8'd182} : s = 192;
	{8'd10,8'd183} : s = 193;
	{8'd10,8'd184} : s = 194;
	{8'd10,8'd185} : s = 195;
	{8'd10,8'd186} : s = 196;
	{8'd10,8'd187} : s = 197;
	{8'd10,8'd188} : s = 198;
	{8'd10,8'd189} : s = 199;
	{8'd10,8'd190} : s = 200;
	{8'd10,8'd191} : s = 201;
	{8'd10,8'd192} : s = 202;
	{8'd10,8'd193} : s = 203;
	{8'd10,8'd194} : s = 204;
	{8'd10,8'd195} : s = 205;
	{8'd10,8'd196} : s = 206;
	{8'd10,8'd197} : s = 207;
	{8'd10,8'd198} : s = 208;
	{8'd10,8'd199} : s = 209;
	{8'd10,8'd200} : s = 210;
	{8'd10,8'd201} : s = 211;
	{8'd10,8'd202} : s = 212;
	{8'd10,8'd203} : s = 213;
	{8'd10,8'd204} : s = 214;
	{8'd10,8'd205} : s = 215;
	{8'd10,8'd206} : s = 216;
	{8'd10,8'd207} : s = 217;
	{8'd10,8'd208} : s = 218;
	{8'd10,8'd209} : s = 219;
	{8'd10,8'd210} : s = 220;
	{8'd10,8'd211} : s = 221;
	{8'd10,8'd212} : s = 222;
	{8'd10,8'd213} : s = 223;
	{8'd10,8'd214} : s = 224;
	{8'd10,8'd215} : s = 225;
	{8'd10,8'd216} : s = 226;
	{8'd10,8'd217} : s = 227;
	{8'd10,8'd218} : s = 228;
	{8'd10,8'd219} : s = 229;
	{8'd10,8'd220} : s = 230;
	{8'd10,8'd221} : s = 231;
	{8'd10,8'd222} : s = 232;
	{8'd10,8'd223} : s = 233;
	{8'd10,8'd224} : s = 234;
	{8'd10,8'd225} : s = 235;
	{8'd10,8'd226} : s = 236;
	{8'd10,8'd227} : s = 237;
	{8'd10,8'd228} : s = 238;
	{8'd10,8'd229} : s = 239;
	{8'd10,8'd230} : s = 240;
	{8'd10,8'd231} : s = 241;
	{8'd10,8'd232} : s = 242;
	{8'd10,8'd233} : s = 243;
	{8'd10,8'd234} : s = 244;
	{8'd10,8'd235} : s = 245;
	{8'd10,8'd236} : s = 246;
	{8'd10,8'd237} : s = 247;
	{8'd10,8'd238} : s = 248;
	{8'd10,8'd239} : s = 249;
	{8'd10,8'd240} : s = 250;
	{8'd10,8'd241} : s = 251;
	{8'd10,8'd242} : s = 252;
	{8'd10,8'd243} : s = 253;
	{8'd10,8'd244} : s = 254;
	{8'd10,8'd245} : s = 255;
	{8'd10,8'd246} : s = 256;
	{8'd10,8'd247} : s = 257;
	{8'd10,8'd248} : s = 258;
	{8'd10,8'd249} : s = 259;
	{8'd10,8'd250} : s = 260;
	{8'd10,8'd251} : s = 261;
	{8'd10,8'd252} : s = 262;
	{8'd10,8'd253} : s = 263;
	{8'd10,8'd254} : s = 264;
	{8'd10,8'd255} : s = 265;
	{8'd11,8'd0} : s = 11;
	{8'd11,8'd1} : s = 12;
	{8'd11,8'd2} : s = 13;
	{8'd11,8'd3} : s = 14;
	{8'd11,8'd4} : s = 15;
	{8'd11,8'd5} : s = 16;
	{8'd11,8'd6} : s = 17;
	{8'd11,8'd7} : s = 18;
	{8'd11,8'd8} : s = 19;
	{8'd11,8'd9} : s = 20;
	{8'd11,8'd10} : s = 21;
	{8'd11,8'd11} : s = 22;
	{8'd11,8'd12} : s = 23;
	{8'd11,8'd13} : s = 24;
	{8'd11,8'd14} : s = 25;
	{8'd11,8'd15} : s = 26;
	{8'd11,8'd16} : s = 27;
	{8'd11,8'd17} : s = 28;
	{8'd11,8'd18} : s = 29;
	{8'd11,8'd19} : s = 30;
	{8'd11,8'd20} : s = 31;
	{8'd11,8'd21} : s = 32;
	{8'd11,8'd22} : s = 33;
	{8'd11,8'd23} : s = 34;
	{8'd11,8'd24} : s = 35;
	{8'd11,8'd25} : s = 36;
	{8'd11,8'd26} : s = 37;
	{8'd11,8'd27} : s = 38;
	{8'd11,8'd28} : s = 39;
	{8'd11,8'd29} : s = 40;
	{8'd11,8'd30} : s = 41;
	{8'd11,8'd31} : s = 42;
	{8'd11,8'd32} : s = 43;
	{8'd11,8'd33} : s = 44;
	{8'd11,8'd34} : s = 45;
	{8'd11,8'd35} : s = 46;
	{8'd11,8'd36} : s = 47;
	{8'd11,8'd37} : s = 48;
	{8'd11,8'd38} : s = 49;
	{8'd11,8'd39} : s = 50;
	{8'd11,8'd40} : s = 51;
	{8'd11,8'd41} : s = 52;
	{8'd11,8'd42} : s = 53;
	{8'd11,8'd43} : s = 54;
	{8'd11,8'd44} : s = 55;
	{8'd11,8'd45} : s = 56;
	{8'd11,8'd46} : s = 57;
	{8'd11,8'd47} : s = 58;
	{8'd11,8'd48} : s = 59;
	{8'd11,8'd49} : s = 60;
	{8'd11,8'd50} : s = 61;
	{8'd11,8'd51} : s = 62;
	{8'd11,8'd52} : s = 63;
	{8'd11,8'd53} : s = 64;
	{8'd11,8'd54} : s = 65;
	{8'd11,8'd55} : s = 66;
	{8'd11,8'd56} : s = 67;
	{8'd11,8'd57} : s = 68;
	{8'd11,8'd58} : s = 69;
	{8'd11,8'd59} : s = 70;
	{8'd11,8'd60} : s = 71;
	{8'd11,8'd61} : s = 72;
	{8'd11,8'd62} : s = 73;
	{8'd11,8'd63} : s = 74;
	{8'd11,8'd64} : s = 75;
	{8'd11,8'd65} : s = 76;
	{8'd11,8'd66} : s = 77;
	{8'd11,8'd67} : s = 78;
	{8'd11,8'd68} : s = 79;
	{8'd11,8'd69} : s = 80;
	{8'd11,8'd70} : s = 81;
	{8'd11,8'd71} : s = 82;
	{8'd11,8'd72} : s = 83;
	{8'd11,8'd73} : s = 84;
	{8'd11,8'd74} : s = 85;
	{8'd11,8'd75} : s = 86;
	{8'd11,8'd76} : s = 87;
	{8'd11,8'd77} : s = 88;
	{8'd11,8'd78} : s = 89;
	{8'd11,8'd79} : s = 90;
	{8'd11,8'd80} : s = 91;
	{8'd11,8'd81} : s = 92;
	{8'd11,8'd82} : s = 93;
	{8'd11,8'd83} : s = 94;
	{8'd11,8'd84} : s = 95;
	{8'd11,8'd85} : s = 96;
	{8'd11,8'd86} : s = 97;
	{8'd11,8'd87} : s = 98;
	{8'd11,8'd88} : s = 99;
	{8'd11,8'd89} : s = 100;
	{8'd11,8'd90} : s = 101;
	{8'd11,8'd91} : s = 102;
	{8'd11,8'd92} : s = 103;
	{8'd11,8'd93} : s = 104;
	{8'd11,8'd94} : s = 105;
	{8'd11,8'd95} : s = 106;
	{8'd11,8'd96} : s = 107;
	{8'd11,8'd97} : s = 108;
	{8'd11,8'd98} : s = 109;
	{8'd11,8'd99} : s = 110;
	{8'd11,8'd100} : s = 111;
	{8'd11,8'd101} : s = 112;
	{8'd11,8'd102} : s = 113;
	{8'd11,8'd103} : s = 114;
	{8'd11,8'd104} : s = 115;
	{8'd11,8'd105} : s = 116;
	{8'd11,8'd106} : s = 117;
	{8'd11,8'd107} : s = 118;
	{8'd11,8'd108} : s = 119;
	{8'd11,8'd109} : s = 120;
	{8'd11,8'd110} : s = 121;
	{8'd11,8'd111} : s = 122;
	{8'd11,8'd112} : s = 123;
	{8'd11,8'd113} : s = 124;
	{8'd11,8'd114} : s = 125;
	{8'd11,8'd115} : s = 126;
	{8'd11,8'd116} : s = 127;
	{8'd11,8'd117} : s = 128;
	{8'd11,8'd118} : s = 129;
	{8'd11,8'd119} : s = 130;
	{8'd11,8'd120} : s = 131;
	{8'd11,8'd121} : s = 132;
	{8'd11,8'd122} : s = 133;
	{8'd11,8'd123} : s = 134;
	{8'd11,8'd124} : s = 135;
	{8'd11,8'd125} : s = 136;
	{8'd11,8'd126} : s = 137;
	{8'd11,8'd127} : s = 138;
	{8'd11,8'd128} : s = 139;
	{8'd11,8'd129} : s = 140;
	{8'd11,8'd130} : s = 141;
	{8'd11,8'd131} : s = 142;
	{8'd11,8'd132} : s = 143;
	{8'd11,8'd133} : s = 144;
	{8'd11,8'd134} : s = 145;
	{8'd11,8'd135} : s = 146;
	{8'd11,8'd136} : s = 147;
	{8'd11,8'd137} : s = 148;
	{8'd11,8'd138} : s = 149;
	{8'd11,8'd139} : s = 150;
	{8'd11,8'd140} : s = 151;
	{8'd11,8'd141} : s = 152;
	{8'd11,8'd142} : s = 153;
	{8'd11,8'd143} : s = 154;
	{8'd11,8'd144} : s = 155;
	{8'd11,8'd145} : s = 156;
	{8'd11,8'd146} : s = 157;
	{8'd11,8'd147} : s = 158;
	{8'd11,8'd148} : s = 159;
	{8'd11,8'd149} : s = 160;
	{8'd11,8'd150} : s = 161;
	{8'd11,8'd151} : s = 162;
	{8'd11,8'd152} : s = 163;
	{8'd11,8'd153} : s = 164;
	{8'd11,8'd154} : s = 165;
	{8'd11,8'd155} : s = 166;
	{8'd11,8'd156} : s = 167;
	{8'd11,8'd157} : s = 168;
	{8'd11,8'd158} : s = 169;
	{8'd11,8'd159} : s = 170;
	{8'd11,8'd160} : s = 171;
	{8'd11,8'd161} : s = 172;
	{8'd11,8'd162} : s = 173;
	{8'd11,8'd163} : s = 174;
	{8'd11,8'd164} : s = 175;
	{8'd11,8'd165} : s = 176;
	{8'd11,8'd166} : s = 177;
	{8'd11,8'd167} : s = 178;
	{8'd11,8'd168} : s = 179;
	{8'd11,8'd169} : s = 180;
	{8'd11,8'd170} : s = 181;
	{8'd11,8'd171} : s = 182;
	{8'd11,8'd172} : s = 183;
	{8'd11,8'd173} : s = 184;
	{8'd11,8'd174} : s = 185;
	{8'd11,8'd175} : s = 186;
	{8'd11,8'd176} : s = 187;
	{8'd11,8'd177} : s = 188;
	{8'd11,8'd178} : s = 189;
	{8'd11,8'd179} : s = 190;
	{8'd11,8'd180} : s = 191;
	{8'd11,8'd181} : s = 192;
	{8'd11,8'd182} : s = 193;
	{8'd11,8'd183} : s = 194;
	{8'd11,8'd184} : s = 195;
	{8'd11,8'd185} : s = 196;
	{8'd11,8'd186} : s = 197;
	{8'd11,8'd187} : s = 198;
	{8'd11,8'd188} : s = 199;
	{8'd11,8'd189} : s = 200;
	{8'd11,8'd190} : s = 201;
	{8'd11,8'd191} : s = 202;
	{8'd11,8'd192} : s = 203;
	{8'd11,8'd193} : s = 204;
	{8'd11,8'd194} : s = 205;
	{8'd11,8'd195} : s = 206;
	{8'd11,8'd196} : s = 207;
	{8'd11,8'd197} : s = 208;
	{8'd11,8'd198} : s = 209;
	{8'd11,8'd199} : s = 210;
	{8'd11,8'd200} : s = 211;
	{8'd11,8'd201} : s = 212;
	{8'd11,8'd202} : s = 213;
	{8'd11,8'd203} : s = 214;
	{8'd11,8'd204} : s = 215;
	{8'd11,8'd205} : s = 216;
	{8'd11,8'd206} : s = 217;
	{8'd11,8'd207} : s = 218;
	{8'd11,8'd208} : s = 219;
	{8'd11,8'd209} : s = 220;
	{8'd11,8'd210} : s = 221;
	{8'd11,8'd211} : s = 222;
	{8'd11,8'd212} : s = 223;
	{8'd11,8'd213} : s = 224;
	{8'd11,8'd214} : s = 225;
	{8'd11,8'd215} : s = 226;
	{8'd11,8'd216} : s = 227;
	{8'd11,8'd217} : s = 228;
	{8'd11,8'd218} : s = 229;
	{8'd11,8'd219} : s = 230;
	{8'd11,8'd220} : s = 231;
	{8'd11,8'd221} : s = 232;
	{8'd11,8'd222} : s = 233;
	{8'd11,8'd223} : s = 234;
	{8'd11,8'd224} : s = 235;
	{8'd11,8'd225} : s = 236;
	{8'd11,8'd226} : s = 237;
	{8'd11,8'd227} : s = 238;
	{8'd11,8'd228} : s = 239;
	{8'd11,8'd229} : s = 240;
	{8'd11,8'd230} : s = 241;
	{8'd11,8'd231} : s = 242;
	{8'd11,8'd232} : s = 243;
	{8'd11,8'd233} : s = 244;
	{8'd11,8'd234} : s = 245;
	{8'd11,8'd235} : s = 246;
	{8'd11,8'd236} : s = 247;
	{8'd11,8'd237} : s = 248;
	{8'd11,8'd238} : s = 249;
	{8'd11,8'd239} : s = 250;
	{8'd11,8'd240} : s = 251;
	{8'd11,8'd241} : s = 252;
	{8'd11,8'd242} : s = 253;
	{8'd11,8'd243} : s = 254;
	{8'd11,8'd244} : s = 255;
	{8'd11,8'd245} : s = 256;
	{8'd11,8'd246} : s = 257;
	{8'd11,8'd247} : s = 258;
	{8'd11,8'd248} : s = 259;
	{8'd11,8'd249} : s = 260;
	{8'd11,8'd250} : s = 261;
	{8'd11,8'd251} : s = 262;
	{8'd11,8'd252} : s = 263;
	{8'd11,8'd253} : s = 264;
	{8'd11,8'd254} : s = 265;
	{8'd11,8'd255} : s = 266;
	{8'd12,8'd0} : s = 12;
	{8'd12,8'd1} : s = 13;
	{8'd12,8'd2} : s = 14;
	{8'd12,8'd3} : s = 15;
	{8'd12,8'd4} : s = 16;
	{8'd12,8'd5} : s = 17;
	{8'd12,8'd6} : s = 18;
	{8'd12,8'd7} : s = 19;
	{8'd12,8'd8} : s = 20;
	{8'd12,8'd9} : s = 21;
	{8'd12,8'd10} : s = 22;
	{8'd12,8'd11} : s = 23;
	{8'd12,8'd12} : s = 24;
	{8'd12,8'd13} : s = 25;
	{8'd12,8'd14} : s = 26;
	{8'd12,8'd15} : s = 27;
	{8'd12,8'd16} : s = 28;
	{8'd12,8'd17} : s = 29;
	{8'd12,8'd18} : s = 30;
	{8'd12,8'd19} : s = 31;
	{8'd12,8'd20} : s = 32;
	{8'd12,8'd21} : s = 33;
	{8'd12,8'd22} : s = 34;
	{8'd12,8'd23} : s = 35;
	{8'd12,8'd24} : s = 36;
	{8'd12,8'd25} : s = 37;
	{8'd12,8'd26} : s = 38;
	{8'd12,8'd27} : s = 39;
	{8'd12,8'd28} : s = 40;
	{8'd12,8'd29} : s = 41;
	{8'd12,8'd30} : s = 42;
	{8'd12,8'd31} : s = 43;
	{8'd12,8'd32} : s = 44;
	{8'd12,8'd33} : s = 45;
	{8'd12,8'd34} : s = 46;
	{8'd12,8'd35} : s = 47;
	{8'd12,8'd36} : s = 48;
	{8'd12,8'd37} : s = 49;
	{8'd12,8'd38} : s = 50;
	{8'd12,8'd39} : s = 51;
	{8'd12,8'd40} : s = 52;
	{8'd12,8'd41} : s = 53;
	{8'd12,8'd42} : s = 54;
	{8'd12,8'd43} : s = 55;
	{8'd12,8'd44} : s = 56;
	{8'd12,8'd45} : s = 57;
	{8'd12,8'd46} : s = 58;
	{8'd12,8'd47} : s = 59;
	{8'd12,8'd48} : s = 60;
	{8'd12,8'd49} : s = 61;
	{8'd12,8'd50} : s = 62;
	{8'd12,8'd51} : s = 63;
	{8'd12,8'd52} : s = 64;
	{8'd12,8'd53} : s = 65;
	{8'd12,8'd54} : s = 66;
	{8'd12,8'd55} : s = 67;
	{8'd12,8'd56} : s = 68;
	{8'd12,8'd57} : s = 69;
	{8'd12,8'd58} : s = 70;
	{8'd12,8'd59} : s = 71;
	{8'd12,8'd60} : s = 72;
	{8'd12,8'd61} : s = 73;
	{8'd12,8'd62} : s = 74;
	{8'd12,8'd63} : s = 75;
	{8'd12,8'd64} : s = 76;
	{8'd12,8'd65} : s = 77;
	{8'd12,8'd66} : s = 78;
	{8'd12,8'd67} : s = 79;
	{8'd12,8'd68} : s = 80;
	{8'd12,8'd69} : s = 81;
	{8'd12,8'd70} : s = 82;
	{8'd12,8'd71} : s = 83;
	{8'd12,8'd72} : s = 84;
	{8'd12,8'd73} : s = 85;
	{8'd12,8'd74} : s = 86;
	{8'd12,8'd75} : s = 87;
	{8'd12,8'd76} : s = 88;
	{8'd12,8'd77} : s = 89;
	{8'd12,8'd78} : s = 90;
	{8'd12,8'd79} : s = 91;
	{8'd12,8'd80} : s = 92;
	{8'd12,8'd81} : s = 93;
	{8'd12,8'd82} : s = 94;
	{8'd12,8'd83} : s = 95;
	{8'd12,8'd84} : s = 96;
	{8'd12,8'd85} : s = 97;
	{8'd12,8'd86} : s = 98;
	{8'd12,8'd87} : s = 99;
	{8'd12,8'd88} : s = 100;
	{8'd12,8'd89} : s = 101;
	{8'd12,8'd90} : s = 102;
	{8'd12,8'd91} : s = 103;
	{8'd12,8'd92} : s = 104;
	{8'd12,8'd93} : s = 105;
	{8'd12,8'd94} : s = 106;
	{8'd12,8'd95} : s = 107;
	{8'd12,8'd96} : s = 108;
	{8'd12,8'd97} : s = 109;
	{8'd12,8'd98} : s = 110;
	{8'd12,8'd99} : s = 111;
	{8'd12,8'd100} : s = 112;
	{8'd12,8'd101} : s = 113;
	{8'd12,8'd102} : s = 114;
	{8'd12,8'd103} : s = 115;
	{8'd12,8'd104} : s = 116;
	{8'd12,8'd105} : s = 117;
	{8'd12,8'd106} : s = 118;
	{8'd12,8'd107} : s = 119;
	{8'd12,8'd108} : s = 120;
	{8'd12,8'd109} : s = 121;
	{8'd12,8'd110} : s = 122;
	{8'd12,8'd111} : s = 123;
	{8'd12,8'd112} : s = 124;
	{8'd12,8'd113} : s = 125;
	{8'd12,8'd114} : s = 126;
	{8'd12,8'd115} : s = 127;
	{8'd12,8'd116} : s = 128;
	{8'd12,8'd117} : s = 129;
	{8'd12,8'd118} : s = 130;
	{8'd12,8'd119} : s = 131;
	{8'd12,8'd120} : s = 132;
	{8'd12,8'd121} : s = 133;
	{8'd12,8'd122} : s = 134;
	{8'd12,8'd123} : s = 135;
	{8'd12,8'd124} : s = 136;
	{8'd12,8'd125} : s = 137;
	{8'd12,8'd126} : s = 138;
	{8'd12,8'd127} : s = 139;
	{8'd12,8'd128} : s = 140;
	{8'd12,8'd129} : s = 141;
	{8'd12,8'd130} : s = 142;
	{8'd12,8'd131} : s = 143;
	{8'd12,8'd132} : s = 144;
	{8'd12,8'd133} : s = 145;
	{8'd12,8'd134} : s = 146;
	{8'd12,8'd135} : s = 147;
	{8'd12,8'd136} : s = 148;
	{8'd12,8'd137} : s = 149;
	{8'd12,8'd138} : s = 150;
	{8'd12,8'd139} : s = 151;
	{8'd12,8'd140} : s = 152;
	{8'd12,8'd141} : s = 153;
	{8'd12,8'd142} : s = 154;
	{8'd12,8'd143} : s = 155;
	{8'd12,8'd144} : s = 156;
	{8'd12,8'd145} : s = 157;
	{8'd12,8'd146} : s = 158;
	{8'd12,8'd147} : s = 159;
	{8'd12,8'd148} : s = 160;
	{8'd12,8'd149} : s = 161;
	{8'd12,8'd150} : s = 162;
	{8'd12,8'd151} : s = 163;
	{8'd12,8'd152} : s = 164;
	{8'd12,8'd153} : s = 165;
	{8'd12,8'd154} : s = 166;
	{8'd12,8'd155} : s = 167;
	{8'd12,8'd156} : s = 168;
	{8'd12,8'd157} : s = 169;
	{8'd12,8'd158} : s = 170;
	{8'd12,8'd159} : s = 171;
	{8'd12,8'd160} : s = 172;
	{8'd12,8'd161} : s = 173;
	{8'd12,8'd162} : s = 174;
	{8'd12,8'd163} : s = 175;
	{8'd12,8'd164} : s = 176;
	{8'd12,8'd165} : s = 177;
	{8'd12,8'd166} : s = 178;
	{8'd12,8'd167} : s = 179;
	{8'd12,8'd168} : s = 180;
	{8'd12,8'd169} : s = 181;
	{8'd12,8'd170} : s = 182;
	{8'd12,8'd171} : s = 183;
	{8'd12,8'd172} : s = 184;
	{8'd12,8'd173} : s = 185;
	{8'd12,8'd174} : s = 186;
	{8'd12,8'd175} : s = 187;
	{8'd12,8'd176} : s = 188;
	{8'd12,8'd177} : s = 189;
	{8'd12,8'd178} : s = 190;
	{8'd12,8'd179} : s = 191;
	{8'd12,8'd180} : s = 192;
	{8'd12,8'd181} : s = 193;
	{8'd12,8'd182} : s = 194;
	{8'd12,8'd183} : s = 195;
	{8'd12,8'd184} : s = 196;
	{8'd12,8'd185} : s = 197;
	{8'd12,8'd186} : s = 198;
	{8'd12,8'd187} : s = 199;
	{8'd12,8'd188} : s = 200;
	{8'd12,8'd189} : s = 201;
	{8'd12,8'd190} : s = 202;
	{8'd12,8'd191} : s = 203;
	{8'd12,8'd192} : s = 204;
	{8'd12,8'd193} : s = 205;
	{8'd12,8'd194} : s = 206;
	{8'd12,8'd195} : s = 207;
	{8'd12,8'd196} : s = 208;
	{8'd12,8'd197} : s = 209;
	{8'd12,8'd198} : s = 210;
	{8'd12,8'd199} : s = 211;
	{8'd12,8'd200} : s = 212;
	{8'd12,8'd201} : s = 213;
	{8'd12,8'd202} : s = 214;
	{8'd12,8'd203} : s = 215;
	{8'd12,8'd204} : s = 216;
	{8'd12,8'd205} : s = 217;
	{8'd12,8'd206} : s = 218;
	{8'd12,8'd207} : s = 219;
	{8'd12,8'd208} : s = 220;
	{8'd12,8'd209} : s = 221;
	{8'd12,8'd210} : s = 222;
	{8'd12,8'd211} : s = 223;
	{8'd12,8'd212} : s = 224;
	{8'd12,8'd213} : s = 225;
	{8'd12,8'd214} : s = 226;
	{8'd12,8'd215} : s = 227;
	{8'd12,8'd216} : s = 228;
	{8'd12,8'd217} : s = 229;
	{8'd12,8'd218} : s = 230;
	{8'd12,8'd219} : s = 231;
	{8'd12,8'd220} : s = 232;
	{8'd12,8'd221} : s = 233;
	{8'd12,8'd222} : s = 234;
	{8'd12,8'd223} : s = 235;
	{8'd12,8'd224} : s = 236;
	{8'd12,8'd225} : s = 237;
	{8'd12,8'd226} : s = 238;
	{8'd12,8'd227} : s = 239;
	{8'd12,8'd228} : s = 240;
	{8'd12,8'd229} : s = 241;
	{8'd12,8'd230} : s = 242;
	{8'd12,8'd231} : s = 243;
	{8'd12,8'd232} : s = 244;
	{8'd12,8'd233} : s = 245;
	{8'd12,8'd234} : s = 246;
	{8'd12,8'd235} : s = 247;
	{8'd12,8'd236} : s = 248;
	{8'd12,8'd237} : s = 249;
	{8'd12,8'd238} : s = 250;
	{8'd12,8'd239} : s = 251;
	{8'd12,8'd240} : s = 252;
	{8'd12,8'd241} : s = 253;
	{8'd12,8'd242} : s = 254;
	{8'd12,8'd243} : s = 255;
	{8'd12,8'd244} : s = 256;
	{8'd12,8'd245} : s = 257;
	{8'd12,8'd246} : s = 258;
	{8'd12,8'd247} : s = 259;
	{8'd12,8'd248} : s = 260;
	{8'd12,8'd249} : s = 261;
	{8'd12,8'd250} : s = 262;
	{8'd12,8'd251} : s = 263;
	{8'd12,8'd252} : s = 264;
	{8'd12,8'd253} : s = 265;
	{8'd12,8'd254} : s = 266;
	{8'd12,8'd255} : s = 267;
	{8'd13,8'd0} : s = 13;
	{8'd13,8'd1} : s = 14;
	{8'd13,8'd2} : s = 15;
	{8'd13,8'd3} : s = 16;
	{8'd13,8'd4} : s = 17;
	{8'd13,8'd5} : s = 18;
	{8'd13,8'd6} : s = 19;
	{8'd13,8'd7} : s = 20;
	{8'd13,8'd8} : s = 21;
	{8'd13,8'd9} : s = 22;
	{8'd13,8'd10} : s = 23;
	{8'd13,8'd11} : s = 24;
	{8'd13,8'd12} : s = 25;
	{8'd13,8'd13} : s = 26;
	{8'd13,8'd14} : s = 27;
	{8'd13,8'd15} : s = 28;
	{8'd13,8'd16} : s = 29;
	{8'd13,8'd17} : s = 30;
	{8'd13,8'd18} : s = 31;
	{8'd13,8'd19} : s = 32;
	{8'd13,8'd20} : s = 33;
	{8'd13,8'd21} : s = 34;
	{8'd13,8'd22} : s = 35;
	{8'd13,8'd23} : s = 36;
	{8'd13,8'd24} : s = 37;
	{8'd13,8'd25} : s = 38;
	{8'd13,8'd26} : s = 39;
	{8'd13,8'd27} : s = 40;
	{8'd13,8'd28} : s = 41;
	{8'd13,8'd29} : s = 42;
	{8'd13,8'd30} : s = 43;
	{8'd13,8'd31} : s = 44;
	{8'd13,8'd32} : s = 45;
	{8'd13,8'd33} : s = 46;
	{8'd13,8'd34} : s = 47;
	{8'd13,8'd35} : s = 48;
	{8'd13,8'd36} : s = 49;
	{8'd13,8'd37} : s = 50;
	{8'd13,8'd38} : s = 51;
	{8'd13,8'd39} : s = 52;
	{8'd13,8'd40} : s = 53;
	{8'd13,8'd41} : s = 54;
	{8'd13,8'd42} : s = 55;
	{8'd13,8'd43} : s = 56;
	{8'd13,8'd44} : s = 57;
	{8'd13,8'd45} : s = 58;
	{8'd13,8'd46} : s = 59;
	{8'd13,8'd47} : s = 60;
	{8'd13,8'd48} : s = 61;
	{8'd13,8'd49} : s = 62;
	{8'd13,8'd50} : s = 63;
	{8'd13,8'd51} : s = 64;
	{8'd13,8'd52} : s = 65;
	{8'd13,8'd53} : s = 66;
	{8'd13,8'd54} : s = 67;
	{8'd13,8'd55} : s = 68;
	{8'd13,8'd56} : s = 69;
	{8'd13,8'd57} : s = 70;
	{8'd13,8'd58} : s = 71;
	{8'd13,8'd59} : s = 72;
	{8'd13,8'd60} : s = 73;
	{8'd13,8'd61} : s = 74;
	{8'd13,8'd62} : s = 75;
	{8'd13,8'd63} : s = 76;
	{8'd13,8'd64} : s = 77;
	{8'd13,8'd65} : s = 78;
	{8'd13,8'd66} : s = 79;
	{8'd13,8'd67} : s = 80;
	{8'd13,8'd68} : s = 81;
	{8'd13,8'd69} : s = 82;
	{8'd13,8'd70} : s = 83;
	{8'd13,8'd71} : s = 84;
	{8'd13,8'd72} : s = 85;
	{8'd13,8'd73} : s = 86;
	{8'd13,8'd74} : s = 87;
	{8'd13,8'd75} : s = 88;
	{8'd13,8'd76} : s = 89;
	{8'd13,8'd77} : s = 90;
	{8'd13,8'd78} : s = 91;
	{8'd13,8'd79} : s = 92;
	{8'd13,8'd80} : s = 93;
	{8'd13,8'd81} : s = 94;
	{8'd13,8'd82} : s = 95;
	{8'd13,8'd83} : s = 96;
	{8'd13,8'd84} : s = 97;
	{8'd13,8'd85} : s = 98;
	{8'd13,8'd86} : s = 99;
	{8'd13,8'd87} : s = 100;
	{8'd13,8'd88} : s = 101;
	{8'd13,8'd89} : s = 102;
	{8'd13,8'd90} : s = 103;
	{8'd13,8'd91} : s = 104;
	{8'd13,8'd92} : s = 105;
	{8'd13,8'd93} : s = 106;
	{8'd13,8'd94} : s = 107;
	{8'd13,8'd95} : s = 108;
	{8'd13,8'd96} : s = 109;
	{8'd13,8'd97} : s = 110;
	{8'd13,8'd98} : s = 111;
	{8'd13,8'd99} : s = 112;
	{8'd13,8'd100} : s = 113;
	{8'd13,8'd101} : s = 114;
	{8'd13,8'd102} : s = 115;
	{8'd13,8'd103} : s = 116;
	{8'd13,8'd104} : s = 117;
	{8'd13,8'd105} : s = 118;
	{8'd13,8'd106} : s = 119;
	{8'd13,8'd107} : s = 120;
	{8'd13,8'd108} : s = 121;
	{8'd13,8'd109} : s = 122;
	{8'd13,8'd110} : s = 123;
	{8'd13,8'd111} : s = 124;
	{8'd13,8'd112} : s = 125;
	{8'd13,8'd113} : s = 126;
	{8'd13,8'd114} : s = 127;
	{8'd13,8'd115} : s = 128;
	{8'd13,8'd116} : s = 129;
	{8'd13,8'd117} : s = 130;
	{8'd13,8'd118} : s = 131;
	{8'd13,8'd119} : s = 132;
	{8'd13,8'd120} : s = 133;
	{8'd13,8'd121} : s = 134;
	{8'd13,8'd122} : s = 135;
	{8'd13,8'd123} : s = 136;
	{8'd13,8'd124} : s = 137;
	{8'd13,8'd125} : s = 138;
	{8'd13,8'd126} : s = 139;
	{8'd13,8'd127} : s = 140;
	{8'd13,8'd128} : s = 141;
	{8'd13,8'd129} : s = 142;
	{8'd13,8'd130} : s = 143;
	{8'd13,8'd131} : s = 144;
	{8'd13,8'd132} : s = 145;
	{8'd13,8'd133} : s = 146;
	{8'd13,8'd134} : s = 147;
	{8'd13,8'd135} : s = 148;
	{8'd13,8'd136} : s = 149;
	{8'd13,8'd137} : s = 150;
	{8'd13,8'd138} : s = 151;
	{8'd13,8'd139} : s = 152;
	{8'd13,8'd140} : s = 153;
	{8'd13,8'd141} : s = 154;
	{8'd13,8'd142} : s = 155;
	{8'd13,8'd143} : s = 156;
	{8'd13,8'd144} : s = 157;
	{8'd13,8'd145} : s = 158;
	{8'd13,8'd146} : s = 159;
	{8'd13,8'd147} : s = 160;
	{8'd13,8'd148} : s = 161;
	{8'd13,8'd149} : s = 162;
	{8'd13,8'd150} : s = 163;
	{8'd13,8'd151} : s = 164;
	{8'd13,8'd152} : s = 165;
	{8'd13,8'd153} : s = 166;
	{8'd13,8'd154} : s = 167;
	{8'd13,8'd155} : s = 168;
	{8'd13,8'd156} : s = 169;
	{8'd13,8'd157} : s = 170;
	{8'd13,8'd158} : s = 171;
	{8'd13,8'd159} : s = 172;
	{8'd13,8'd160} : s = 173;
	{8'd13,8'd161} : s = 174;
	{8'd13,8'd162} : s = 175;
	{8'd13,8'd163} : s = 176;
	{8'd13,8'd164} : s = 177;
	{8'd13,8'd165} : s = 178;
	{8'd13,8'd166} : s = 179;
	{8'd13,8'd167} : s = 180;
	{8'd13,8'd168} : s = 181;
	{8'd13,8'd169} : s = 182;
	{8'd13,8'd170} : s = 183;
	{8'd13,8'd171} : s = 184;
	{8'd13,8'd172} : s = 185;
	{8'd13,8'd173} : s = 186;
	{8'd13,8'd174} : s = 187;
	{8'd13,8'd175} : s = 188;
	{8'd13,8'd176} : s = 189;
	{8'd13,8'd177} : s = 190;
	{8'd13,8'd178} : s = 191;
	{8'd13,8'd179} : s = 192;
	{8'd13,8'd180} : s = 193;
	{8'd13,8'd181} : s = 194;
	{8'd13,8'd182} : s = 195;
	{8'd13,8'd183} : s = 196;
	{8'd13,8'd184} : s = 197;
	{8'd13,8'd185} : s = 198;
	{8'd13,8'd186} : s = 199;
	{8'd13,8'd187} : s = 200;
	{8'd13,8'd188} : s = 201;
	{8'd13,8'd189} : s = 202;
	{8'd13,8'd190} : s = 203;
	{8'd13,8'd191} : s = 204;
	{8'd13,8'd192} : s = 205;
	{8'd13,8'd193} : s = 206;
	{8'd13,8'd194} : s = 207;
	{8'd13,8'd195} : s = 208;
	{8'd13,8'd196} : s = 209;
	{8'd13,8'd197} : s = 210;
	{8'd13,8'd198} : s = 211;
	{8'd13,8'd199} : s = 212;
	{8'd13,8'd200} : s = 213;
	{8'd13,8'd201} : s = 214;
	{8'd13,8'd202} : s = 215;
	{8'd13,8'd203} : s = 216;
	{8'd13,8'd204} : s = 217;
	{8'd13,8'd205} : s = 218;
	{8'd13,8'd206} : s = 219;
	{8'd13,8'd207} : s = 220;
	{8'd13,8'd208} : s = 221;
	{8'd13,8'd209} : s = 222;
	{8'd13,8'd210} : s = 223;
	{8'd13,8'd211} : s = 224;
	{8'd13,8'd212} : s = 225;
	{8'd13,8'd213} : s = 226;
	{8'd13,8'd214} : s = 227;
	{8'd13,8'd215} : s = 228;
	{8'd13,8'd216} : s = 229;
	{8'd13,8'd217} : s = 230;
	{8'd13,8'd218} : s = 231;
	{8'd13,8'd219} : s = 232;
	{8'd13,8'd220} : s = 233;
	{8'd13,8'd221} : s = 234;
	{8'd13,8'd222} : s = 235;
	{8'd13,8'd223} : s = 236;
	{8'd13,8'd224} : s = 237;
	{8'd13,8'd225} : s = 238;
	{8'd13,8'd226} : s = 239;
	{8'd13,8'd227} : s = 240;
	{8'd13,8'd228} : s = 241;
	{8'd13,8'd229} : s = 242;
	{8'd13,8'd230} : s = 243;
	{8'd13,8'd231} : s = 244;
	{8'd13,8'd232} : s = 245;
	{8'd13,8'd233} : s = 246;
	{8'd13,8'd234} : s = 247;
	{8'd13,8'd235} : s = 248;
	{8'd13,8'd236} : s = 249;
	{8'd13,8'd237} : s = 250;
	{8'd13,8'd238} : s = 251;
	{8'd13,8'd239} : s = 252;
	{8'd13,8'd240} : s = 253;
	{8'd13,8'd241} : s = 254;
	{8'd13,8'd242} : s = 255;
	{8'd13,8'd243} : s = 256;
	{8'd13,8'd244} : s = 257;
	{8'd13,8'd245} : s = 258;
	{8'd13,8'd246} : s = 259;
	{8'd13,8'd247} : s = 260;
	{8'd13,8'd248} : s = 261;
	{8'd13,8'd249} : s = 262;
	{8'd13,8'd250} : s = 263;
	{8'd13,8'd251} : s = 264;
	{8'd13,8'd252} : s = 265;
	{8'd13,8'd253} : s = 266;
	{8'd13,8'd254} : s = 267;
	{8'd13,8'd255} : s = 268;
	{8'd14,8'd0} : s = 14;
	{8'd14,8'd1} : s = 15;
	{8'd14,8'd2} : s = 16;
	{8'd14,8'd3} : s = 17;
	{8'd14,8'd4} : s = 18;
	{8'd14,8'd5} : s = 19;
	{8'd14,8'd6} : s = 20;
	{8'd14,8'd7} : s = 21;
	{8'd14,8'd8} : s = 22;
	{8'd14,8'd9} : s = 23;
	{8'd14,8'd10} : s = 24;
	{8'd14,8'd11} : s = 25;
	{8'd14,8'd12} : s = 26;
	{8'd14,8'd13} : s = 27;
	{8'd14,8'd14} : s = 28;
	{8'd14,8'd15} : s = 29;
	{8'd14,8'd16} : s = 30;
	{8'd14,8'd17} : s = 31;
	{8'd14,8'd18} : s = 32;
	{8'd14,8'd19} : s = 33;
	{8'd14,8'd20} : s = 34;
	{8'd14,8'd21} : s = 35;
	{8'd14,8'd22} : s = 36;
	{8'd14,8'd23} : s = 37;
	{8'd14,8'd24} : s = 38;
	{8'd14,8'd25} : s = 39;
	{8'd14,8'd26} : s = 40;
	{8'd14,8'd27} : s = 41;
	{8'd14,8'd28} : s = 42;
	{8'd14,8'd29} : s = 43;
	{8'd14,8'd30} : s = 44;
	{8'd14,8'd31} : s = 45;
	{8'd14,8'd32} : s = 46;
	{8'd14,8'd33} : s = 47;
	{8'd14,8'd34} : s = 48;
	{8'd14,8'd35} : s = 49;
	{8'd14,8'd36} : s = 50;
	{8'd14,8'd37} : s = 51;
	{8'd14,8'd38} : s = 52;
	{8'd14,8'd39} : s = 53;
	{8'd14,8'd40} : s = 54;
	{8'd14,8'd41} : s = 55;
	{8'd14,8'd42} : s = 56;
	{8'd14,8'd43} : s = 57;
	{8'd14,8'd44} : s = 58;
	{8'd14,8'd45} : s = 59;
	{8'd14,8'd46} : s = 60;
	{8'd14,8'd47} : s = 61;
	{8'd14,8'd48} : s = 62;
	{8'd14,8'd49} : s = 63;
	{8'd14,8'd50} : s = 64;
	{8'd14,8'd51} : s = 65;
	{8'd14,8'd52} : s = 66;
	{8'd14,8'd53} : s = 67;
	{8'd14,8'd54} : s = 68;
	{8'd14,8'd55} : s = 69;
	{8'd14,8'd56} : s = 70;
	{8'd14,8'd57} : s = 71;
	{8'd14,8'd58} : s = 72;
	{8'd14,8'd59} : s = 73;
	{8'd14,8'd60} : s = 74;
	{8'd14,8'd61} : s = 75;
	{8'd14,8'd62} : s = 76;
	{8'd14,8'd63} : s = 77;
	{8'd14,8'd64} : s = 78;
	{8'd14,8'd65} : s = 79;
	{8'd14,8'd66} : s = 80;
	{8'd14,8'd67} : s = 81;
	{8'd14,8'd68} : s = 82;
	{8'd14,8'd69} : s = 83;
	{8'd14,8'd70} : s = 84;
	{8'd14,8'd71} : s = 85;
	{8'd14,8'd72} : s = 86;
	{8'd14,8'd73} : s = 87;
	{8'd14,8'd74} : s = 88;
	{8'd14,8'd75} : s = 89;
	{8'd14,8'd76} : s = 90;
	{8'd14,8'd77} : s = 91;
	{8'd14,8'd78} : s = 92;
	{8'd14,8'd79} : s = 93;
	{8'd14,8'd80} : s = 94;
	{8'd14,8'd81} : s = 95;
	{8'd14,8'd82} : s = 96;
	{8'd14,8'd83} : s = 97;
	{8'd14,8'd84} : s = 98;
	{8'd14,8'd85} : s = 99;
	{8'd14,8'd86} : s = 100;
	{8'd14,8'd87} : s = 101;
	{8'd14,8'd88} : s = 102;
	{8'd14,8'd89} : s = 103;
	{8'd14,8'd90} : s = 104;
	{8'd14,8'd91} : s = 105;
	{8'd14,8'd92} : s = 106;
	{8'd14,8'd93} : s = 107;
	{8'd14,8'd94} : s = 108;
	{8'd14,8'd95} : s = 109;
	{8'd14,8'd96} : s = 110;
	{8'd14,8'd97} : s = 111;
	{8'd14,8'd98} : s = 112;
	{8'd14,8'd99} : s = 113;
	{8'd14,8'd100} : s = 114;
	{8'd14,8'd101} : s = 115;
	{8'd14,8'd102} : s = 116;
	{8'd14,8'd103} : s = 117;
	{8'd14,8'd104} : s = 118;
	{8'd14,8'd105} : s = 119;
	{8'd14,8'd106} : s = 120;
	{8'd14,8'd107} : s = 121;
	{8'd14,8'd108} : s = 122;
	{8'd14,8'd109} : s = 123;
	{8'd14,8'd110} : s = 124;
	{8'd14,8'd111} : s = 125;
	{8'd14,8'd112} : s = 126;
	{8'd14,8'd113} : s = 127;
	{8'd14,8'd114} : s = 128;
	{8'd14,8'd115} : s = 129;
	{8'd14,8'd116} : s = 130;
	{8'd14,8'd117} : s = 131;
	{8'd14,8'd118} : s = 132;
	{8'd14,8'd119} : s = 133;
	{8'd14,8'd120} : s = 134;
	{8'd14,8'd121} : s = 135;
	{8'd14,8'd122} : s = 136;
	{8'd14,8'd123} : s = 137;
	{8'd14,8'd124} : s = 138;
	{8'd14,8'd125} : s = 139;
	{8'd14,8'd126} : s = 140;
	{8'd14,8'd127} : s = 141;
	{8'd14,8'd128} : s = 142;
	{8'd14,8'd129} : s = 143;
	{8'd14,8'd130} : s = 144;
	{8'd14,8'd131} : s = 145;
	{8'd14,8'd132} : s = 146;
	{8'd14,8'd133} : s = 147;
	{8'd14,8'd134} : s = 148;
	{8'd14,8'd135} : s = 149;
	{8'd14,8'd136} : s = 150;
	{8'd14,8'd137} : s = 151;
	{8'd14,8'd138} : s = 152;
	{8'd14,8'd139} : s = 153;
	{8'd14,8'd140} : s = 154;
	{8'd14,8'd141} : s = 155;
	{8'd14,8'd142} : s = 156;
	{8'd14,8'd143} : s = 157;
	{8'd14,8'd144} : s = 158;
	{8'd14,8'd145} : s = 159;
	{8'd14,8'd146} : s = 160;
	{8'd14,8'd147} : s = 161;
	{8'd14,8'd148} : s = 162;
	{8'd14,8'd149} : s = 163;
	{8'd14,8'd150} : s = 164;
	{8'd14,8'd151} : s = 165;
	{8'd14,8'd152} : s = 166;
	{8'd14,8'd153} : s = 167;
	{8'd14,8'd154} : s = 168;
	{8'd14,8'd155} : s = 169;
	{8'd14,8'd156} : s = 170;
	{8'd14,8'd157} : s = 171;
	{8'd14,8'd158} : s = 172;
	{8'd14,8'd159} : s = 173;
	{8'd14,8'd160} : s = 174;
	{8'd14,8'd161} : s = 175;
	{8'd14,8'd162} : s = 176;
	{8'd14,8'd163} : s = 177;
	{8'd14,8'd164} : s = 178;
	{8'd14,8'd165} : s = 179;
	{8'd14,8'd166} : s = 180;
	{8'd14,8'd167} : s = 181;
	{8'd14,8'd168} : s = 182;
	{8'd14,8'd169} : s = 183;
	{8'd14,8'd170} : s = 184;
	{8'd14,8'd171} : s = 185;
	{8'd14,8'd172} : s = 186;
	{8'd14,8'd173} : s = 187;
	{8'd14,8'd174} : s = 188;
	{8'd14,8'd175} : s = 189;
	{8'd14,8'd176} : s = 190;
	{8'd14,8'd177} : s = 191;
	{8'd14,8'd178} : s = 192;
	{8'd14,8'd179} : s = 193;
	{8'd14,8'd180} : s = 194;
	{8'd14,8'd181} : s = 195;
	{8'd14,8'd182} : s = 196;
	{8'd14,8'd183} : s = 197;
	{8'd14,8'd184} : s = 198;
	{8'd14,8'd185} : s = 199;
	{8'd14,8'd186} : s = 200;
	{8'd14,8'd187} : s = 201;
	{8'd14,8'd188} : s = 202;
	{8'd14,8'd189} : s = 203;
	{8'd14,8'd190} : s = 204;
	{8'd14,8'd191} : s = 205;
	{8'd14,8'd192} : s = 206;
	{8'd14,8'd193} : s = 207;
	{8'd14,8'd194} : s = 208;
	{8'd14,8'd195} : s = 209;
	{8'd14,8'd196} : s = 210;
	{8'd14,8'd197} : s = 211;
	{8'd14,8'd198} : s = 212;
	{8'd14,8'd199} : s = 213;
	{8'd14,8'd200} : s = 214;
	{8'd14,8'd201} : s = 215;
	{8'd14,8'd202} : s = 216;
	{8'd14,8'd203} : s = 217;
	{8'd14,8'd204} : s = 218;
	{8'd14,8'd205} : s = 219;
	{8'd14,8'd206} : s = 220;
	{8'd14,8'd207} : s = 221;
	{8'd14,8'd208} : s = 222;
	{8'd14,8'd209} : s = 223;
	{8'd14,8'd210} : s = 224;
	{8'd14,8'd211} : s = 225;
	{8'd14,8'd212} : s = 226;
	{8'd14,8'd213} : s = 227;
	{8'd14,8'd214} : s = 228;
	{8'd14,8'd215} : s = 229;
	{8'd14,8'd216} : s = 230;
	{8'd14,8'd217} : s = 231;
	{8'd14,8'd218} : s = 232;
	{8'd14,8'd219} : s = 233;
	{8'd14,8'd220} : s = 234;
	{8'd14,8'd221} : s = 235;
	{8'd14,8'd222} : s = 236;
	{8'd14,8'd223} : s = 237;
	{8'd14,8'd224} : s = 238;
	{8'd14,8'd225} : s = 239;
	{8'd14,8'd226} : s = 240;
	{8'd14,8'd227} : s = 241;
	{8'd14,8'd228} : s = 242;
	{8'd14,8'd229} : s = 243;
	{8'd14,8'd230} : s = 244;
	{8'd14,8'd231} : s = 245;
	{8'd14,8'd232} : s = 246;
	{8'd14,8'd233} : s = 247;
	{8'd14,8'd234} : s = 248;
	{8'd14,8'd235} : s = 249;
	{8'd14,8'd236} : s = 250;
	{8'd14,8'd237} : s = 251;
	{8'd14,8'd238} : s = 252;
	{8'd14,8'd239} : s = 253;
	{8'd14,8'd240} : s = 254;
	{8'd14,8'd241} : s = 255;
	{8'd14,8'd242} : s = 256;
	{8'd14,8'd243} : s = 257;
	{8'd14,8'd244} : s = 258;
	{8'd14,8'd245} : s = 259;
	{8'd14,8'd246} : s = 260;
	{8'd14,8'd247} : s = 261;
	{8'd14,8'd248} : s = 262;
	{8'd14,8'd249} : s = 263;
	{8'd14,8'd250} : s = 264;
	{8'd14,8'd251} : s = 265;
	{8'd14,8'd252} : s = 266;
	{8'd14,8'd253} : s = 267;
	{8'd14,8'd254} : s = 268;
	{8'd14,8'd255} : s = 269;
	{8'd15,8'd0} : s = 15;
	{8'd15,8'd1} : s = 16;
	{8'd15,8'd2} : s = 17;
	{8'd15,8'd3} : s = 18;
	{8'd15,8'd4} : s = 19;
	{8'd15,8'd5} : s = 20;
	{8'd15,8'd6} : s = 21;
	{8'd15,8'd7} : s = 22;
	{8'd15,8'd8} : s = 23;
	{8'd15,8'd9} : s = 24;
	{8'd15,8'd10} : s = 25;
	{8'd15,8'd11} : s = 26;
	{8'd15,8'd12} : s = 27;
	{8'd15,8'd13} : s = 28;
	{8'd15,8'd14} : s = 29;
	{8'd15,8'd15} : s = 30;
	{8'd15,8'd16} : s = 31;
	{8'd15,8'd17} : s = 32;
	{8'd15,8'd18} : s = 33;
	{8'd15,8'd19} : s = 34;
	{8'd15,8'd20} : s = 35;
	{8'd15,8'd21} : s = 36;
	{8'd15,8'd22} : s = 37;
	{8'd15,8'd23} : s = 38;
	{8'd15,8'd24} : s = 39;
	{8'd15,8'd25} : s = 40;
	{8'd15,8'd26} : s = 41;
	{8'd15,8'd27} : s = 42;
	{8'd15,8'd28} : s = 43;
	{8'd15,8'd29} : s = 44;
	{8'd15,8'd30} : s = 45;
	{8'd15,8'd31} : s = 46;
	{8'd15,8'd32} : s = 47;
	{8'd15,8'd33} : s = 48;
	{8'd15,8'd34} : s = 49;
	{8'd15,8'd35} : s = 50;
	{8'd15,8'd36} : s = 51;
	{8'd15,8'd37} : s = 52;
	{8'd15,8'd38} : s = 53;
	{8'd15,8'd39} : s = 54;
	{8'd15,8'd40} : s = 55;
	{8'd15,8'd41} : s = 56;
	{8'd15,8'd42} : s = 57;
	{8'd15,8'd43} : s = 58;
	{8'd15,8'd44} : s = 59;
	{8'd15,8'd45} : s = 60;
	{8'd15,8'd46} : s = 61;
	{8'd15,8'd47} : s = 62;
	{8'd15,8'd48} : s = 63;
	{8'd15,8'd49} : s = 64;
	{8'd15,8'd50} : s = 65;
	{8'd15,8'd51} : s = 66;
	{8'd15,8'd52} : s = 67;
	{8'd15,8'd53} : s = 68;
	{8'd15,8'd54} : s = 69;
	{8'd15,8'd55} : s = 70;
	{8'd15,8'd56} : s = 71;
	{8'd15,8'd57} : s = 72;
	{8'd15,8'd58} : s = 73;
	{8'd15,8'd59} : s = 74;
	{8'd15,8'd60} : s = 75;
	{8'd15,8'd61} : s = 76;
	{8'd15,8'd62} : s = 77;
	{8'd15,8'd63} : s = 78;
	{8'd15,8'd64} : s = 79;
	{8'd15,8'd65} : s = 80;
	{8'd15,8'd66} : s = 81;
	{8'd15,8'd67} : s = 82;
	{8'd15,8'd68} : s = 83;
	{8'd15,8'd69} : s = 84;
	{8'd15,8'd70} : s = 85;
	{8'd15,8'd71} : s = 86;
	{8'd15,8'd72} : s = 87;
	{8'd15,8'd73} : s = 88;
	{8'd15,8'd74} : s = 89;
	{8'd15,8'd75} : s = 90;
	{8'd15,8'd76} : s = 91;
	{8'd15,8'd77} : s = 92;
	{8'd15,8'd78} : s = 93;
	{8'd15,8'd79} : s = 94;
	{8'd15,8'd80} : s = 95;
	{8'd15,8'd81} : s = 96;
	{8'd15,8'd82} : s = 97;
	{8'd15,8'd83} : s = 98;
	{8'd15,8'd84} : s = 99;
	{8'd15,8'd85} : s = 100;
	{8'd15,8'd86} : s = 101;
	{8'd15,8'd87} : s = 102;
	{8'd15,8'd88} : s = 103;
	{8'd15,8'd89} : s = 104;
	{8'd15,8'd90} : s = 105;
	{8'd15,8'd91} : s = 106;
	{8'd15,8'd92} : s = 107;
	{8'd15,8'd93} : s = 108;
	{8'd15,8'd94} : s = 109;
	{8'd15,8'd95} : s = 110;
	{8'd15,8'd96} : s = 111;
	{8'd15,8'd97} : s = 112;
	{8'd15,8'd98} : s = 113;
	{8'd15,8'd99} : s = 114;
	{8'd15,8'd100} : s = 115;
	{8'd15,8'd101} : s = 116;
	{8'd15,8'd102} : s = 117;
	{8'd15,8'd103} : s = 118;
	{8'd15,8'd104} : s = 119;
	{8'd15,8'd105} : s = 120;
	{8'd15,8'd106} : s = 121;
	{8'd15,8'd107} : s = 122;
	{8'd15,8'd108} : s = 123;
	{8'd15,8'd109} : s = 124;
	{8'd15,8'd110} : s = 125;
	{8'd15,8'd111} : s = 126;
	{8'd15,8'd112} : s = 127;
	{8'd15,8'd113} : s = 128;
	{8'd15,8'd114} : s = 129;
	{8'd15,8'd115} : s = 130;
	{8'd15,8'd116} : s = 131;
	{8'd15,8'd117} : s = 132;
	{8'd15,8'd118} : s = 133;
	{8'd15,8'd119} : s = 134;
	{8'd15,8'd120} : s = 135;
	{8'd15,8'd121} : s = 136;
	{8'd15,8'd122} : s = 137;
	{8'd15,8'd123} : s = 138;
	{8'd15,8'd124} : s = 139;
	{8'd15,8'd125} : s = 140;
	{8'd15,8'd126} : s = 141;
	{8'd15,8'd127} : s = 142;
	{8'd15,8'd128} : s = 143;
	{8'd15,8'd129} : s = 144;
	{8'd15,8'd130} : s = 145;
	{8'd15,8'd131} : s = 146;
	{8'd15,8'd132} : s = 147;
	{8'd15,8'd133} : s = 148;
	{8'd15,8'd134} : s = 149;
	{8'd15,8'd135} : s = 150;
	{8'd15,8'd136} : s = 151;
	{8'd15,8'd137} : s = 152;
	{8'd15,8'd138} : s = 153;
	{8'd15,8'd139} : s = 154;
	{8'd15,8'd140} : s = 155;
	{8'd15,8'd141} : s = 156;
	{8'd15,8'd142} : s = 157;
	{8'd15,8'd143} : s = 158;
	{8'd15,8'd144} : s = 159;
	{8'd15,8'd145} : s = 160;
	{8'd15,8'd146} : s = 161;
	{8'd15,8'd147} : s = 162;
	{8'd15,8'd148} : s = 163;
	{8'd15,8'd149} : s = 164;
	{8'd15,8'd150} : s = 165;
	{8'd15,8'd151} : s = 166;
	{8'd15,8'd152} : s = 167;
	{8'd15,8'd153} : s = 168;
	{8'd15,8'd154} : s = 169;
	{8'd15,8'd155} : s = 170;
	{8'd15,8'd156} : s = 171;
	{8'd15,8'd157} : s = 172;
	{8'd15,8'd158} : s = 173;
	{8'd15,8'd159} : s = 174;
	{8'd15,8'd160} : s = 175;
	{8'd15,8'd161} : s = 176;
	{8'd15,8'd162} : s = 177;
	{8'd15,8'd163} : s = 178;
	{8'd15,8'd164} : s = 179;
	{8'd15,8'd165} : s = 180;
	{8'd15,8'd166} : s = 181;
	{8'd15,8'd167} : s = 182;
	{8'd15,8'd168} : s = 183;
	{8'd15,8'd169} : s = 184;
	{8'd15,8'd170} : s = 185;
	{8'd15,8'd171} : s = 186;
	{8'd15,8'd172} : s = 187;
	{8'd15,8'd173} : s = 188;
	{8'd15,8'd174} : s = 189;
	{8'd15,8'd175} : s = 190;
	{8'd15,8'd176} : s = 191;
	{8'd15,8'd177} : s = 192;
	{8'd15,8'd178} : s = 193;
	{8'd15,8'd179} : s = 194;
	{8'd15,8'd180} : s = 195;
	{8'd15,8'd181} : s = 196;
	{8'd15,8'd182} : s = 197;
	{8'd15,8'd183} : s = 198;
	{8'd15,8'd184} : s = 199;
	{8'd15,8'd185} : s = 200;
	{8'd15,8'd186} : s = 201;
	{8'd15,8'd187} : s = 202;
	{8'd15,8'd188} : s = 203;
	{8'd15,8'd189} : s = 204;
	{8'd15,8'd190} : s = 205;
	{8'd15,8'd191} : s = 206;
	{8'd15,8'd192} : s = 207;
	{8'd15,8'd193} : s = 208;
	{8'd15,8'd194} : s = 209;
	{8'd15,8'd195} : s = 210;
	{8'd15,8'd196} : s = 211;
	{8'd15,8'd197} : s = 212;
	{8'd15,8'd198} : s = 213;
	{8'd15,8'd199} : s = 214;
	{8'd15,8'd200} : s = 215;
	{8'd15,8'd201} : s = 216;
	{8'd15,8'd202} : s = 217;
	{8'd15,8'd203} : s = 218;
	{8'd15,8'd204} : s = 219;
	{8'd15,8'd205} : s = 220;
	{8'd15,8'd206} : s = 221;
	{8'd15,8'd207} : s = 222;
	{8'd15,8'd208} : s = 223;
	{8'd15,8'd209} : s = 224;
	{8'd15,8'd210} : s = 225;
	{8'd15,8'd211} : s = 226;
	{8'd15,8'd212} : s = 227;
	{8'd15,8'd213} : s = 228;
	{8'd15,8'd214} : s = 229;
	{8'd15,8'd215} : s = 230;
	{8'd15,8'd216} : s = 231;
	{8'd15,8'd217} : s = 232;
	{8'd15,8'd218} : s = 233;
	{8'd15,8'd219} : s = 234;
	{8'd15,8'd220} : s = 235;
	{8'd15,8'd221} : s = 236;
	{8'd15,8'd222} : s = 237;
	{8'd15,8'd223} : s = 238;
	{8'd15,8'd224} : s = 239;
	{8'd15,8'd225} : s = 240;
	{8'd15,8'd226} : s = 241;
	{8'd15,8'd227} : s = 242;
	{8'd15,8'd228} : s = 243;
	{8'd15,8'd229} : s = 244;
	{8'd15,8'd230} : s = 245;
	{8'd15,8'd231} : s = 246;
	{8'd15,8'd232} : s = 247;
	{8'd15,8'd233} : s = 248;
	{8'd15,8'd234} : s = 249;
	{8'd15,8'd235} : s = 250;
	{8'd15,8'd236} : s = 251;
	{8'd15,8'd237} : s = 252;
	{8'd15,8'd238} : s = 253;
	{8'd15,8'd239} : s = 254;
	{8'd15,8'd240} : s = 255;
	{8'd15,8'd241} : s = 256;
	{8'd15,8'd242} : s = 257;
	{8'd15,8'd243} : s = 258;
	{8'd15,8'd244} : s = 259;
	{8'd15,8'd245} : s = 260;
	{8'd15,8'd246} : s = 261;
	{8'd15,8'd247} : s = 262;
	{8'd15,8'd248} : s = 263;
	{8'd15,8'd249} : s = 264;
	{8'd15,8'd250} : s = 265;
	{8'd15,8'd251} : s = 266;
	{8'd15,8'd252} : s = 267;
	{8'd15,8'd253} : s = 268;
	{8'd15,8'd254} : s = 269;
	{8'd15,8'd255} : s = 270;
	{8'd16,8'd0} : s = 16;
	{8'd16,8'd1} : s = 17;
	{8'd16,8'd2} : s = 18;
	{8'd16,8'd3} : s = 19;
	{8'd16,8'd4} : s = 20;
	{8'd16,8'd5} : s = 21;
	{8'd16,8'd6} : s = 22;
	{8'd16,8'd7} : s = 23;
	{8'd16,8'd8} : s = 24;
	{8'd16,8'd9} : s = 25;
	{8'd16,8'd10} : s = 26;
	{8'd16,8'd11} : s = 27;
	{8'd16,8'd12} : s = 28;
	{8'd16,8'd13} : s = 29;
	{8'd16,8'd14} : s = 30;
	{8'd16,8'd15} : s = 31;
	{8'd16,8'd16} : s = 32;
	{8'd16,8'd17} : s = 33;
	{8'd16,8'd18} : s = 34;
	{8'd16,8'd19} : s = 35;
	{8'd16,8'd20} : s = 36;
	{8'd16,8'd21} : s = 37;
	{8'd16,8'd22} : s = 38;
	{8'd16,8'd23} : s = 39;
	{8'd16,8'd24} : s = 40;
	{8'd16,8'd25} : s = 41;
	{8'd16,8'd26} : s = 42;
	{8'd16,8'd27} : s = 43;
	{8'd16,8'd28} : s = 44;
	{8'd16,8'd29} : s = 45;
	{8'd16,8'd30} : s = 46;
	{8'd16,8'd31} : s = 47;
	{8'd16,8'd32} : s = 48;
	{8'd16,8'd33} : s = 49;
	{8'd16,8'd34} : s = 50;
	{8'd16,8'd35} : s = 51;
	{8'd16,8'd36} : s = 52;
	{8'd16,8'd37} : s = 53;
	{8'd16,8'd38} : s = 54;
	{8'd16,8'd39} : s = 55;
	{8'd16,8'd40} : s = 56;
	{8'd16,8'd41} : s = 57;
	{8'd16,8'd42} : s = 58;
	{8'd16,8'd43} : s = 59;
	{8'd16,8'd44} : s = 60;
	{8'd16,8'd45} : s = 61;
	{8'd16,8'd46} : s = 62;
	{8'd16,8'd47} : s = 63;
	{8'd16,8'd48} : s = 64;
	{8'd16,8'd49} : s = 65;
	{8'd16,8'd50} : s = 66;
	{8'd16,8'd51} : s = 67;
	{8'd16,8'd52} : s = 68;
	{8'd16,8'd53} : s = 69;
	{8'd16,8'd54} : s = 70;
	{8'd16,8'd55} : s = 71;
	{8'd16,8'd56} : s = 72;
	{8'd16,8'd57} : s = 73;
	{8'd16,8'd58} : s = 74;
	{8'd16,8'd59} : s = 75;
	{8'd16,8'd60} : s = 76;
	{8'd16,8'd61} : s = 77;
	{8'd16,8'd62} : s = 78;
	{8'd16,8'd63} : s = 79;
	{8'd16,8'd64} : s = 80;
	{8'd16,8'd65} : s = 81;
	{8'd16,8'd66} : s = 82;
	{8'd16,8'd67} : s = 83;
	{8'd16,8'd68} : s = 84;
	{8'd16,8'd69} : s = 85;
	{8'd16,8'd70} : s = 86;
	{8'd16,8'd71} : s = 87;
	{8'd16,8'd72} : s = 88;
	{8'd16,8'd73} : s = 89;
	{8'd16,8'd74} : s = 90;
	{8'd16,8'd75} : s = 91;
	{8'd16,8'd76} : s = 92;
	{8'd16,8'd77} : s = 93;
	{8'd16,8'd78} : s = 94;
	{8'd16,8'd79} : s = 95;
	{8'd16,8'd80} : s = 96;
	{8'd16,8'd81} : s = 97;
	{8'd16,8'd82} : s = 98;
	{8'd16,8'd83} : s = 99;
	{8'd16,8'd84} : s = 100;
	{8'd16,8'd85} : s = 101;
	{8'd16,8'd86} : s = 102;
	{8'd16,8'd87} : s = 103;
	{8'd16,8'd88} : s = 104;
	{8'd16,8'd89} : s = 105;
	{8'd16,8'd90} : s = 106;
	{8'd16,8'd91} : s = 107;
	{8'd16,8'd92} : s = 108;
	{8'd16,8'd93} : s = 109;
	{8'd16,8'd94} : s = 110;
	{8'd16,8'd95} : s = 111;
	{8'd16,8'd96} : s = 112;
	{8'd16,8'd97} : s = 113;
	{8'd16,8'd98} : s = 114;
	{8'd16,8'd99} : s = 115;
	{8'd16,8'd100} : s = 116;
	{8'd16,8'd101} : s = 117;
	{8'd16,8'd102} : s = 118;
	{8'd16,8'd103} : s = 119;
	{8'd16,8'd104} : s = 120;
	{8'd16,8'd105} : s = 121;
	{8'd16,8'd106} : s = 122;
	{8'd16,8'd107} : s = 123;
	{8'd16,8'd108} : s = 124;
	{8'd16,8'd109} : s = 125;
	{8'd16,8'd110} : s = 126;
	{8'd16,8'd111} : s = 127;
	{8'd16,8'd112} : s = 128;
	{8'd16,8'd113} : s = 129;
	{8'd16,8'd114} : s = 130;
	{8'd16,8'd115} : s = 131;
	{8'd16,8'd116} : s = 132;
	{8'd16,8'd117} : s = 133;
	{8'd16,8'd118} : s = 134;
	{8'd16,8'd119} : s = 135;
	{8'd16,8'd120} : s = 136;
	{8'd16,8'd121} : s = 137;
	{8'd16,8'd122} : s = 138;
	{8'd16,8'd123} : s = 139;
	{8'd16,8'd124} : s = 140;
	{8'd16,8'd125} : s = 141;
	{8'd16,8'd126} : s = 142;
	{8'd16,8'd127} : s = 143;
	{8'd16,8'd128} : s = 144;
	{8'd16,8'd129} : s = 145;
	{8'd16,8'd130} : s = 146;
	{8'd16,8'd131} : s = 147;
	{8'd16,8'd132} : s = 148;
	{8'd16,8'd133} : s = 149;
	{8'd16,8'd134} : s = 150;
	{8'd16,8'd135} : s = 151;
	{8'd16,8'd136} : s = 152;
	{8'd16,8'd137} : s = 153;
	{8'd16,8'd138} : s = 154;
	{8'd16,8'd139} : s = 155;
	{8'd16,8'd140} : s = 156;
	{8'd16,8'd141} : s = 157;
	{8'd16,8'd142} : s = 158;
	{8'd16,8'd143} : s = 159;
	{8'd16,8'd144} : s = 160;
	{8'd16,8'd145} : s = 161;
	{8'd16,8'd146} : s = 162;
	{8'd16,8'd147} : s = 163;
	{8'd16,8'd148} : s = 164;
	{8'd16,8'd149} : s = 165;
	{8'd16,8'd150} : s = 166;
	{8'd16,8'd151} : s = 167;
	{8'd16,8'd152} : s = 168;
	{8'd16,8'd153} : s = 169;
	{8'd16,8'd154} : s = 170;
	{8'd16,8'd155} : s = 171;
	{8'd16,8'd156} : s = 172;
	{8'd16,8'd157} : s = 173;
	{8'd16,8'd158} : s = 174;
	{8'd16,8'd159} : s = 175;
	{8'd16,8'd160} : s = 176;
	{8'd16,8'd161} : s = 177;
	{8'd16,8'd162} : s = 178;
	{8'd16,8'd163} : s = 179;
	{8'd16,8'd164} : s = 180;
	{8'd16,8'd165} : s = 181;
	{8'd16,8'd166} : s = 182;
	{8'd16,8'd167} : s = 183;
	{8'd16,8'd168} : s = 184;
	{8'd16,8'd169} : s = 185;
	{8'd16,8'd170} : s = 186;
	{8'd16,8'd171} : s = 187;
	{8'd16,8'd172} : s = 188;
	{8'd16,8'd173} : s = 189;
	{8'd16,8'd174} : s = 190;
	{8'd16,8'd175} : s = 191;
	{8'd16,8'd176} : s = 192;
	{8'd16,8'd177} : s = 193;
	{8'd16,8'd178} : s = 194;
	{8'd16,8'd179} : s = 195;
	{8'd16,8'd180} : s = 196;
	{8'd16,8'd181} : s = 197;
	{8'd16,8'd182} : s = 198;
	{8'd16,8'd183} : s = 199;
	{8'd16,8'd184} : s = 200;
	{8'd16,8'd185} : s = 201;
	{8'd16,8'd186} : s = 202;
	{8'd16,8'd187} : s = 203;
	{8'd16,8'd188} : s = 204;
	{8'd16,8'd189} : s = 205;
	{8'd16,8'd190} : s = 206;
	{8'd16,8'd191} : s = 207;
	{8'd16,8'd192} : s = 208;
	{8'd16,8'd193} : s = 209;
	{8'd16,8'd194} : s = 210;
	{8'd16,8'd195} : s = 211;
	{8'd16,8'd196} : s = 212;
	{8'd16,8'd197} : s = 213;
	{8'd16,8'd198} : s = 214;
	{8'd16,8'd199} : s = 215;
	{8'd16,8'd200} : s = 216;
	{8'd16,8'd201} : s = 217;
	{8'd16,8'd202} : s = 218;
	{8'd16,8'd203} : s = 219;
	{8'd16,8'd204} : s = 220;
	{8'd16,8'd205} : s = 221;
	{8'd16,8'd206} : s = 222;
	{8'd16,8'd207} : s = 223;
	{8'd16,8'd208} : s = 224;
	{8'd16,8'd209} : s = 225;
	{8'd16,8'd210} : s = 226;
	{8'd16,8'd211} : s = 227;
	{8'd16,8'd212} : s = 228;
	{8'd16,8'd213} : s = 229;
	{8'd16,8'd214} : s = 230;
	{8'd16,8'd215} : s = 231;
	{8'd16,8'd216} : s = 232;
	{8'd16,8'd217} : s = 233;
	{8'd16,8'd218} : s = 234;
	{8'd16,8'd219} : s = 235;
	{8'd16,8'd220} : s = 236;
	{8'd16,8'd221} : s = 237;
	{8'd16,8'd222} : s = 238;
	{8'd16,8'd223} : s = 239;
	{8'd16,8'd224} : s = 240;
	{8'd16,8'd225} : s = 241;
	{8'd16,8'd226} : s = 242;
	{8'd16,8'd227} : s = 243;
	{8'd16,8'd228} : s = 244;
	{8'd16,8'd229} : s = 245;
	{8'd16,8'd230} : s = 246;
	{8'd16,8'd231} : s = 247;
	{8'd16,8'd232} : s = 248;
	{8'd16,8'd233} : s = 249;
	{8'd16,8'd234} : s = 250;
	{8'd16,8'd235} : s = 251;
	{8'd16,8'd236} : s = 252;
	{8'd16,8'd237} : s = 253;
	{8'd16,8'd238} : s = 254;
	{8'd16,8'd239} : s = 255;
	{8'd16,8'd240} : s = 256;
	{8'd16,8'd241} : s = 257;
	{8'd16,8'd242} : s = 258;
	{8'd16,8'd243} : s = 259;
	{8'd16,8'd244} : s = 260;
	{8'd16,8'd245} : s = 261;
	{8'd16,8'd246} : s = 262;
	{8'd16,8'd247} : s = 263;
	{8'd16,8'd248} : s = 264;
	{8'd16,8'd249} : s = 265;
	{8'd16,8'd250} : s = 266;
	{8'd16,8'd251} : s = 267;
	{8'd16,8'd252} : s = 268;
	{8'd16,8'd253} : s = 269;
	{8'd16,8'd254} : s = 270;
	{8'd16,8'd255} : s = 271;
	{8'd17,8'd0} : s = 17;
	{8'd17,8'd1} : s = 18;
	{8'd17,8'd2} : s = 19;
	{8'd17,8'd3} : s = 20;
	{8'd17,8'd4} : s = 21;
	{8'd17,8'd5} : s = 22;
	{8'd17,8'd6} : s = 23;
	{8'd17,8'd7} : s = 24;
	{8'd17,8'd8} : s = 25;
	{8'd17,8'd9} : s = 26;
	{8'd17,8'd10} : s = 27;
	{8'd17,8'd11} : s = 28;
	{8'd17,8'd12} : s = 29;
	{8'd17,8'd13} : s = 30;
	{8'd17,8'd14} : s = 31;
	{8'd17,8'd15} : s = 32;
	{8'd17,8'd16} : s = 33;
	{8'd17,8'd17} : s = 34;
	{8'd17,8'd18} : s = 35;
	{8'd17,8'd19} : s = 36;
	{8'd17,8'd20} : s = 37;
	{8'd17,8'd21} : s = 38;
	{8'd17,8'd22} : s = 39;
	{8'd17,8'd23} : s = 40;
	{8'd17,8'd24} : s = 41;
	{8'd17,8'd25} : s = 42;
	{8'd17,8'd26} : s = 43;
	{8'd17,8'd27} : s = 44;
	{8'd17,8'd28} : s = 45;
	{8'd17,8'd29} : s = 46;
	{8'd17,8'd30} : s = 47;
	{8'd17,8'd31} : s = 48;
	{8'd17,8'd32} : s = 49;
	{8'd17,8'd33} : s = 50;
	{8'd17,8'd34} : s = 51;
	{8'd17,8'd35} : s = 52;
	{8'd17,8'd36} : s = 53;
	{8'd17,8'd37} : s = 54;
	{8'd17,8'd38} : s = 55;
	{8'd17,8'd39} : s = 56;
	{8'd17,8'd40} : s = 57;
	{8'd17,8'd41} : s = 58;
	{8'd17,8'd42} : s = 59;
	{8'd17,8'd43} : s = 60;
	{8'd17,8'd44} : s = 61;
	{8'd17,8'd45} : s = 62;
	{8'd17,8'd46} : s = 63;
	{8'd17,8'd47} : s = 64;
	{8'd17,8'd48} : s = 65;
	{8'd17,8'd49} : s = 66;
	{8'd17,8'd50} : s = 67;
	{8'd17,8'd51} : s = 68;
	{8'd17,8'd52} : s = 69;
	{8'd17,8'd53} : s = 70;
	{8'd17,8'd54} : s = 71;
	{8'd17,8'd55} : s = 72;
	{8'd17,8'd56} : s = 73;
	{8'd17,8'd57} : s = 74;
	{8'd17,8'd58} : s = 75;
	{8'd17,8'd59} : s = 76;
	{8'd17,8'd60} : s = 77;
	{8'd17,8'd61} : s = 78;
	{8'd17,8'd62} : s = 79;
	{8'd17,8'd63} : s = 80;
	{8'd17,8'd64} : s = 81;
	{8'd17,8'd65} : s = 82;
	{8'd17,8'd66} : s = 83;
	{8'd17,8'd67} : s = 84;
	{8'd17,8'd68} : s = 85;
	{8'd17,8'd69} : s = 86;
	{8'd17,8'd70} : s = 87;
	{8'd17,8'd71} : s = 88;
	{8'd17,8'd72} : s = 89;
	{8'd17,8'd73} : s = 90;
	{8'd17,8'd74} : s = 91;
	{8'd17,8'd75} : s = 92;
	{8'd17,8'd76} : s = 93;
	{8'd17,8'd77} : s = 94;
	{8'd17,8'd78} : s = 95;
	{8'd17,8'd79} : s = 96;
	{8'd17,8'd80} : s = 97;
	{8'd17,8'd81} : s = 98;
	{8'd17,8'd82} : s = 99;
	{8'd17,8'd83} : s = 100;
	{8'd17,8'd84} : s = 101;
	{8'd17,8'd85} : s = 102;
	{8'd17,8'd86} : s = 103;
	{8'd17,8'd87} : s = 104;
	{8'd17,8'd88} : s = 105;
	{8'd17,8'd89} : s = 106;
	{8'd17,8'd90} : s = 107;
	{8'd17,8'd91} : s = 108;
	{8'd17,8'd92} : s = 109;
	{8'd17,8'd93} : s = 110;
	{8'd17,8'd94} : s = 111;
	{8'd17,8'd95} : s = 112;
	{8'd17,8'd96} : s = 113;
	{8'd17,8'd97} : s = 114;
	{8'd17,8'd98} : s = 115;
	{8'd17,8'd99} : s = 116;
	{8'd17,8'd100} : s = 117;
	{8'd17,8'd101} : s = 118;
	{8'd17,8'd102} : s = 119;
	{8'd17,8'd103} : s = 120;
	{8'd17,8'd104} : s = 121;
	{8'd17,8'd105} : s = 122;
	{8'd17,8'd106} : s = 123;
	{8'd17,8'd107} : s = 124;
	{8'd17,8'd108} : s = 125;
	{8'd17,8'd109} : s = 126;
	{8'd17,8'd110} : s = 127;
	{8'd17,8'd111} : s = 128;
	{8'd17,8'd112} : s = 129;
	{8'd17,8'd113} : s = 130;
	{8'd17,8'd114} : s = 131;
	{8'd17,8'd115} : s = 132;
	{8'd17,8'd116} : s = 133;
	{8'd17,8'd117} : s = 134;
	{8'd17,8'd118} : s = 135;
	{8'd17,8'd119} : s = 136;
	{8'd17,8'd120} : s = 137;
	{8'd17,8'd121} : s = 138;
	{8'd17,8'd122} : s = 139;
	{8'd17,8'd123} : s = 140;
	{8'd17,8'd124} : s = 141;
	{8'd17,8'd125} : s = 142;
	{8'd17,8'd126} : s = 143;
	{8'd17,8'd127} : s = 144;
	{8'd17,8'd128} : s = 145;
	{8'd17,8'd129} : s = 146;
	{8'd17,8'd130} : s = 147;
	{8'd17,8'd131} : s = 148;
	{8'd17,8'd132} : s = 149;
	{8'd17,8'd133} : s = 150;
	{8'd17,8'd134} : s = 151;
	{8'd17,8'd135} : s = 152;
	{8'd17,8'd136} : s = 153;
	{8'd17,8'd137} : s = 154;
	{8'd17,8'd138} : s = 155;
	{8'd17,8'd139} : s = 156;
	{8'd17,8'd140} : s = 157;
	{8'd17,8'd141} : s = 158;
	{8'd17,8'd142} : s = 159;
	{8'd17,8'd143} : s = 160;
	{8'd17,8'd144} : s = 161;
	{8'd17,8'd145} : s = 162;
	{8'd17,8'd146} : s = 163;
	{8'd17,8'd147} : s = 164;
	{8'd17,8'd148} : s = 165;
	{8'd17,8'd149} : s = 166;
	{8'd17,8'd150} : s = 167;
	{8'd17,8'd151} : s = 168;
	{8'd17,8'd152} : s = 169;
	{8'd17,8'd153} : s = 170;
	{8'd17,8'd154} : s = 171;
	{8'd17,8'd155} : s = 172;
	{8'd17,8'd156} : s = 173;
	{8'd17,8'd157} : s = 174;
	{8'd17,8'd158} : s = 175;
	{8'd17,8'd159} : s = 176;
	{8'd17,8'd160} : s = 177;
	{8'd17,8'd161} : s = 178;
	{8'd17,8'd162} : s = 179;
	{8'd17,8'd163} : s = 180;
	{8'd17,8'd164} : s = 181;
	{8'd17,8'd165} : s = 182;
	{8'd17,8'd166} : s = 183;
	{8'd17,8'd167} : s = 184;
	{8'd17,8'd168} : s = 185;
	{8'd17,8'd169} : s = 186;
	{8'd17,8'd170} : s = 187;
	{8'd17,8'd171} : s = 188;
	{8'd17,8'd172} : s = 189;
	{8'd17,8'd173} : s = 190;
	{8'd17,8'd174} : s = 191;
	{8'd17,8'd175} : s = 192;
	{8'd17,8'd176} : s = 193;
	{8'd17,8'd177} : s = 194;
	{8'd17,8'd178} : s = 195;
	{8'd17,8'd179} : s = 196;
	{8'd17,8'd180} : s = 197;
	{8'd17,8'd181} : s = 198;
	{8'd17,8'd182} : s = 199;
	{8'd17,8'd183} : s = 200;
	{8'd17,8'd184} : s = 201;
	{8'd17,8'd185} : s = 202;
	{8'd17,8'd186} : s = 203;
	{8'd17,8'd187} : s = 204;
	{8'd17,8'd188} : s = 205;
	{8'd17,8'd189} : s = 206;
	{8'd17,8'd190} : s = 207;
	{8'd17,8'd191} : s = 208;
	{8'd17,8'd192} : s = 209;
	{8'd17,8'd193} : s = 210;
	{8'd17,8'd194} : s = 211;
	{8'd17,8'd195} : s = 212;
	{8'd17,8'd196} : s = 213;
	{8'd17,8'd197} : s = 214;
	{8'd17,8'd198} : s = 215;
	{8'd17,8'd199} : s = 216;
	{8'd17,8'd200} : s = 217;
	{8'd17,8'd201} : s = 218;
	{8'd17,8'd202} : s = 219;
	{8'd17,8'd203} : s = 220;
	{8'd17,8'd204} : s = 221;
	{8'd17,8'd205} : s = 222;
	{8'd17,8'd206} : s = 223;
	{8'd17,8'd207} : s = 224;
	{8'd17,8'd208} : s = 225;
	{8'd17,8'd209} : s = 226;
	{8'd17,8'd210} : s = 227;
	{8'd17,8'd211} : s = 228;
	{8'd17,8'd212} : s = 229;
	{8'd17,8'd213} : s = 230;
	{8'd17,8'd214} : s = 231;
	{8'd17,8'd215} : s = 232;
	{8'd17,8'd216} : s = 233;
	{8'd17,8'd217} : s = 234;
	{8'd17,8'd218} : s = 235;
	{8'd17,8'd219} : s = 236;
	{8'd17,8'd220} : s = 237;
	{8'd17,8'd221} : s = 238;
	{8'd17,8'd222} : s = 239;
	{8'd17,8'd223} : s = 240;
	{8'd17,8'd224} : s = 241;
	{8'd17,8'd225} : s = 242;
	{8'd17,8'd226} : s = 243;
	{8'd17,8'd227} : s = 244;
	{8'd17,8'd228} : s = 245;
	{8'd17,8'd229} : s = 246;
	{8'd17,8'd230} : s = 247;
	{8'd17,8'd231} : s = 248;
	{8'd17,8'd232} : s = 249;
	{8'd17,8'd233} : s = 250;
	{8'd17,8'd234} : s = 251;
	{8'd17,8'd235} : s = 252;
	{8'd17,8'd236} : s = 253;
	{8'd17,8'd237} : s = 254;
	{8'd17,8'd238} : s = 255;
	{8'd17,8'd239} : s = 256;
	{8'd17,8'd240} : s = 257;
	{8'd17,8'd241} : s = 258;
	{8'd17,8'd242} : s = 259;
	{8'd17,8'd243} : s = 260;
	{8'd17,8'd244} : s = 261;
	{8'd17,8'd245} : s = 262;
	{8'd17,8'd246} : s = 263;
	{8'd17,8'd247} : s = 264;
	{8'd17,8'd248} : s = 265;
	{8'd17,8'd249} : s = 266;
	{8'd17,8'd250} : s = 267;
	{8'd17,8'd251} : s = 268;
	{8'd17,8'd252} : s = 269;
	{8'd17,8'd253} : s = 270;
	{8'd17,8'd254} : s = 271;
	{8'd17,8'd255} : s = 272;
	{8'd18,8'd0} : s = 18;
	{8'd18,8'd1} : s = 19;
	{8'd18,8'd2} : s = 20;
	{8'd18,8'd3} : s = 21;
	{8'd18,8'd4} : s = 22;
	{8'd18,8'd5} : s = 23;
	{8'd18,8'd6} : s = 24;
	{8'd18,8'd7} : s = 25;
	{8'd18,8'd8} : s = 26;
	{8'd18,8'd9} : s = 27;
	{8'd18,8'd10} : s = 28;
	{8'd18,8'd11} : s = 29;
	{8'd18,8'd12} : s = 30;
	{8'd18,8'd13} : s = 31;
	{8'd18,8'd14} : s = 32;
	{8'd18,8'd15} : s = 33;
	{8'd18,8'd16} : s = 34;
	{8'd18,8'd17} : s = 35;
	{8'd18,8'd18} : s = 36;
	{8'd18,8'd19} : s = 37;
	{8'd18,8'd20} : s = 38;
	{8'd18,8'd21} : s = 39;
	{8'd18,8'd22} : s = 40;
	{8'd18,8'd23} : s = 41;
	{8'd18,8'd24} : s = 42;
	{8'd18,8'd25} : s = 43;
	{8'd18,8'd26} : s = 44;
	{8'd18,8'd27} : s = 45;
	{8'd18,8'd28} : s = 46;
	{8'd18,8'd29} : s = 47;
	{8'd18,8'd30} : s = 48;
	{8'd18,8'd31} : s = 49;
	{8'd18,8'd32} : s = 50;
	{8'd18,8'd33} : s = 51;
	{8'd18,8'd34} : s = 52;
	{8'd18,8'd35} : s = 53;
	{8'd18,8'd36} : s = 54;
	{8'd18,8'd37} : s = 55;
	{8'd18,8'd38} : s = 56;
	{8'd18,8'd39} : s = 57;
	{8'd18,8'd40} : s = 58;
	{8'd18,8'd41} : s = 59;
	{8'd18,8'd42} : s = 60;
	{8'd18,8'd43} : s = 61;
	{8'd18,8'd44} : s = 62;
	{8'd18,8'd45} : s = 63;
	{8'd18,8'd46} : s = 64;
	{8'd18,8'd47} : s = 65;
	{8'd18,8'd48} : s = 66;
	{8'd18,8'd49} : s = 67;
	{8'd18,8'd50} : s = 68;
	{8'd18,8'd51} : s = 69;
	{8'd18,8'd52} : s = 70;
	{8'd18,8'd53} : s = 71;
	{8'd18,8'd54} : s = 72;
	{8'd18,8'd55} : s = 73;
	{8'd18,8'd56} : s = 74;
	{8'd18,8'd57} : s = 75;
	{8'd18,8'd58} : s = 76;
	{8'd18,8'd59} : s = 77;
	{8'd18,8'd60} : s = 78;
	{8'd18,8'd61} : s = 79;
	{8'd18,8'd62} : s = 80;
	{8'd18,8'd63} : s = 81;
	{8'd18,8'd64} : s = 82;
	{8'd18,8'd65} : s = 83;
	{8'd18,8'd66} : s = 84;
	{8'd18,8'd67} : s = 85;
	{8'd18,8'd68} : s = 86;
	{8'd18,8'd69} : s = 87;
	{8'd18,8'd70} : s = 88;
	{8'd18,8'd71} : s = 89;
	{8'd18,8'd72} : s = 90;
	{8'd18,8'd73} : s = 91;
	{8'd18,8'd74} : s = 92;
	{8'd18,8'd75} : s = 93;
	{8'd18,8'd76} : s = 94;
	{8'd18,8'd77} : s = 95;
	{8'd18,8'd78} : s = 96;
	{8'd18,8'd79} : s = 97;
	{8'd18,8'd80} : s = 98;
	{8'd18,8'd81} : s = 99;
	{8'd18,8'd82} : s = 100;
	{8'd18,8'd83} : s = 101;
	{8'd18,8'd84} : s = 102;
	{8'd18,8'd85} : s = 103;
	{8'd18,8'd86} : s = 104;
	{8'd18,8'd87} : s = 105;
	{8'd18,8'd88} : s = 106;
	{8'd18,8'd89} : s = 107;
	{8'd18,8'd90} : s = 108;
	{8'd18,8'd91} : s = 109;
	{8'd18,8'd92} : s = 110;
	{8'd18,8'd93} : s = 111;
	{8'd18,8'd94} : s = 112;
	{8'd18,8'd95} : s = 113;
	{8'd18,8'd96} : s = 114;
	{8'd18,8'd97} : s = 115;
	{8'd18,8'd98} : s = 116;
	{8'd18,8'd99} : s = 117;
	{8'd18,8'd100} : s = 118;
	{8'd18,8'd101} : s = 119;
	{8'd18,8'd102} : s = 120;
	{8'd18,8'd103} : s = 121;
	{8'd18,8'd104} : s = 122;
	{8'd18,8'd105} : s = 123;
	{8'd18,8'd106} : s = 124;
	{8'd18,8'd107} : s = 125;
	{8'd18,8'd108} : s = 126;
	{8'd18,8'd109} : s = 127;
	{8'd18,8'd110} : s = 128;
	{8'd18,8'd111} : s = 129;
	{8'd18,8'd112} : s = 130;
	{8'd18,8'd113} : s = 131;
	{8'd18,8'd114} : s = 132;
	{8'd18,8'd115} : s = 133;
	{8'd18,8'd116} : s = 134;
	{8'd18,8'd117} : s = 135;
	{8'd18,8'd118} : s = 136;
	{8'd18,8'd119} : s = 137;
	{8'd18,8'd120} : s = 138;
	{8'd18,8'd121} : s = 139;
	{8'd18,8'd122} : s = 140;
	{8'd18,8'd123} : s = 141;
	{8'd18,8'd124} : s = 142;
	{8'd18,8'd125} : s = 143;
	{8'd18,8'd126} : s = 144;
	{8'd18,8'd127} : s = 145;
	{8'd18,8'd128} : s = 146;
	{8'd18,8'd129} : s = 147;
	{8'd18,8'd130} : s = 148;
	{8'd18,8'd131} : s = 149;
	{8'd18,8'd132} : s = 150;
	{8'd18,8'd133} : s = 151;
	{8'd18,8'd134} : s = 152;
	{8'd18,8'd135} : s = 153;
	{8'd18,8'd136} : s = 154;
	{8'd18,8'd137} : s = 155;
	{8'd18,8'd138} : s = 156;
	{8'd18,8'd139} : s = 157;
	{8'd18,8'd140} : s = 158;
	{8'd18,8'd141} : s = 159;
	{8'd18,8'd142} : s = 160;
	{8'd18,8'd143} : s = 161;
	{8'd18,8'd144} : s = 162;
	{8'd18,8'd145} : s = 163;
	{8'd18,8'd146} : s = 164;
	{8'd18,8'd147} : s = 165;
	{8'd18,8'd148} : s = 166;
	{8'd18,8'd149} : s = 167;
	{8'd18,8'd150} : s = 168;
	{8'd18,8'd151} : s = 169;
	{8'd18,8'd152} : s = 170;
	{8'd18,8'd153} : s = 171;
	{8'd18,8'd154} : s = 172;
	{8'd18,8'd155} : s = 173;
	{8'd18,8'd156} : s = 174;
	{8'd18,8'd157} : s = 175;
	{8'd18,8'd158} : s = 176;
	{8'd18,8'd159} : s = 177;
	{8'd18,8'd160} : s = 178;
	{8'd18,8'd161} : s = 179;
	{8'd18,8'd162} : s = 180;
	{8'd18,8'd163} : s = 181;
	{8'd18,8'd164} : s = 182;
	{8'd18,8'd165} : s = 183;
	{8'd18,8'd166} : s = 184;
	{8'd18,8'd167} : s = 185;
	{8'd18,8'd168} : s = 186;
	{8'd18,8'd169} : s = 187;
	{8'd18,8'd170} : s = 188;
	{8'd18,8'd171} : s = 189;
	{8'd18,8'd172} : s = 190;
	{8'd18,8'd173} : s = 191;
	{8'd18,8'd174} : s = 192;
	{8'd18,8'd175} : s = 193;
	{8'd18,8'd176} : s = 194;
	{8'd18,8'd177} : s = 195;
	{8'd18,8'd178} : s = 196;
	{8'd18,8'd179} : s = 197;
	{8'd18,8'd180} : s = 198;
	{8'd18,8'd181} : s = 199;
	{8'd18,8'd182} : s = 200;
	{8'd18,8'd183} : s = 201;
	{8'd18,8'd184} : s = 202;
	{8'd18,8'd185} : s = 203;
	{8'd18,8'd186} : s = 204;
	{8'd18,8'd187} : s = 205;
	{8'd18,8'd188} : s = 206;
	{8'd18,8'd189} : s = 207;
	{8'd18,8'd190} : s = 208;
	{8'd18,8'd191} : s = 209;
	{8'd18,8'd192} : s = 210;
	{8'd18,8'd193} : s = 211;
	{8'd18,8'd194} : s = 212;
	{8'd18,8'd195} : s = 213;
	{8'd18,8'd196} : s = 214;
	{8'd18,8'd197} : s = 215;
	{8'd18,8'd198} : s = 216;
	{8'd18,8'd199} : s = 217;
	{8'd18,8'd200} : s = 218;
	{8'd18,8'd201} : s = 219;
	{8'd18,8'd202} : s = 220;
	{8'd18,8'd203} : s = 221;
	{8'd18,8'd204} : s = 222;
	{8'd18,8'd205} : s = 223;
	{8'd18,8'd206} : s = 224;
	{8'd18,8'd207} : s = 225;
	{8'd18,8'd208} : s = 226;
	{8'd18,8'd209} : s = 227;
	{8'd18,8'd210} : s = 228;
	{8'd18,8'd211} : s = 229;
	{8'd18,8'd212} : s = 230;
	{8'd18,8'd213} : s = 231;
	{8'd18,8'd214} : s = 232;
	{8'd18,8'd215} : s = 233;
	{8'd18,8'd216} : s = 234;
	{8'd18,8'd217} : s = 235;
	{8'd18,8'd218} : s = 236;
	{8'd18,8'd219} : s = 237;
	{8'd18,8'd220} : s = 238;
	{8'd18,8'd221} : s = 239;
	{8'd18,8'd222} : s = 240;
	{8'd18,8'd223} : s = 241;
	{8'd18,8'd224} : s = 242;
	{8'd18,8'd225} : s = 243;
	{8'd18,8'd226} : s = 244;
	{8'd18,8'd227} : s = 245;
	{8'd18,8'd228} : s = 246;
	{8'd18,8'd229} : s = 247;
	{8'd18,8'd230} : s = 248;
	{8'd18,8'd231} : s = 249;
	{8'd18,8'd232} : s = 250;
	{8'd18,8'd233} : s = 251;
	{8'd18,8'd234} : s = 252;
	{8'd18,8'd235} : s = 253;
	{8'd18,8'd236} : s = 254;
	{8'd18,8'd237} : s = 255;
	{8'd18,8'd238} : s = 256;
	{8'd18,8'd239} : s = 257;
	{8'd18,8'd240} : s = 258;
	{8'd18,8'd241} : s = 259;
	{8'd18,8'd242} : s = 260;
	{8'd18,8'd243} : s = 261;
	{8'd18,8'd244} : s = 262;
	{8'd18,8'd245} : s = 263;
	{8'd18,8'd246} : s = 264;
	{8'd18,8'd247} : s = 265;
	{8'd18,8'd248} : s = 266;
	{8'd18,8'd249} : s = 267;
	{8'd18,8'd250} : s = 268;
	{8'd18,8'd251} : s = 269;
	{8'd18,8'd252} : s = 270;
	{8'd18,8'd253} : s = 271;
	{8'd18,8'd254} : s = 272;
	{8'd18,8'd255} : s = 273;
	{8'd19,8'd0} : s = 19;
	{8'd19,8'd1} : s = 20;
	{8'd19,8'd2} : s = 21;
	{8'd19,8'd3} : s = 22;
	{8'd19,8'd4} : s = 23;
	{8'd19,8'd5} : s = 24;
	{8'd19,8'd6} : s = 25;
	{8'd19,8'd7} : s = 26;
	{8'd19,8'd8} : s = 27;
	{8'd19,8'd9} : s = 28;
	{8'd19,8'd10} : s = 29;
	{8'd19,8'd11} : s = 30;
	{8'd19,8'd12} : s = 31;
	{8'd19,8'd13} : s = 32;
	{8'd19,8'd14} : s = 33;
	{8'd19,8'd15} : s = 34;
	{8'd19,8'd16} : s = 35;
	{8'd19,8'd17} : s = 36;
	{8'd19,8'd18} : s = 37;
	{8'd19,8'd19} : s = 38;
	{8'd19,8'd20} : s = 39;
	{8'd19,8'd21} : s = 40;
	{8'd19,8'd22} : s = 41;
	{8'd19,8'd23} : s = 42;
	{8'd19,8'd24} : s = 43;
	{8'd19,8'd25} : s = 44;
	{8'd19,8'd26} : s = 45;
	{8'd19,8'd27} : s = 46;
	{8'd19,8'd28} : s = 47;
	{8'd19,8'd29} : s = 48;
	{8'd19,8'd30} : s = 49;
	{8'd19,8'd31} : s = 50;
	{8'd19,8'd32} : s = 51;
	{8'd19,8'd33} : s = 52;
	{8'd19,8'd34} : s = 53;
	{8'd19,8'd35} : s = 54;
	{8'd19,8'd36} : s = 55;
	{8'd19,8'd37} : s = 56;
	{8'd19,8'd38} : s = 57;
	{8'd19,8'd39} : s = 58;
	{8'd19,8'd40} : s = 59;
	{8'd19,8'd41} : s = 60;
	{8'd19,8'd42} : s = 61;
	{8'd19,8'd43} : s = 62;
	{8'd19,8'd44} : s = 63;
	{8'd19,8'd45} : s = 64;
	{8'd19,8'd46} : s = 65;
	{8'd19,8'd47} : s = 66;
	{8'd19,8'd48} : s = 67;
	{8'd19,8'd49} : s = 68;
	{8'd19,8'd50} : s = 69;
	{8'd19,8'd51} : s = 70;
	{8'd19,8'd52} : s = 71;
	{8'd19,8'd53} : s = 72;
	{8'd19,8'd54} : s = 73;
	{8'd19,8'd55} : s = 74;
	{8'd19,8'd56} : s = 75;
	{8'd19,8'd57} : s = 76;
	{8'd19,8'd58} : s = 77;
	{8'd19,8'd59} : s = 78;
	{8'd19,8'd60} : s = 79;
	{8'd19,8'd61} : s = 80;
	{8'd19,8'd62} : s = 81;
	{8'd19,8'd63} : s = 82;
	{8'd19,8'd64} : s = 83;
	{8'd19,8'd65} : s = 84;
	{8'd19,8'd66} : s = 85;
	{8'd19,8'd67} : s = 86;
	{8'd19,8'd68} : s = 87;
	{8'd19,8'd69} : s = 88;
	{8'd19,8'd70} : s = 89;
	{8'd19,8'd71} : s = 90;
	{8'd19,8'd72} : s = 91;
	{8'd19,8'd73} : s = 92;
	{8'd19,8'd74} : s = 93;
	{8'd19,8'd75} : s = 94;
	{8'd19,8'd76} : s = 95;
	{8'd19,8'd77} : s = 96;
	{8'd19,8'd78} : s = 97;
	{8'd19,8'd79} : s = 98;
	{8'd19,8'd80} : s = 99;
	{8'd19,8'd81} : s = 100;
	{8'd19,8'd82} : s = 101;
	{8'd19,8'd83} : s = 102;
	{8'd19,8'd84} : s = 103;
	{8'd19,8'd85} : s = 104;
	{8'd19,8'd86} : s = 105;
	{8'd19,8'd87} : s = 106;
	{8'd19,8'd88} : s = 107;
	{8'd19,8'd89} : s = 108;
	{8'd19,8'd90} : s = 109;
	{8'd19,8'd91} : s = 110;
	{8'd19,8'd92} : s = 111;
	{8'd19,8'd93} : s = 112;
	{8'd19,8'd94} : s = 113;
	{8'd19,8'd95} : s = 114;
	{8'd19,8'd96} : s = 115;
	{8'd19,8'd97} : s = 116;
	{8'd19,8'd98} : s = 117;
	{8'd19,8'd99} : s = 118;
	{8'd19,8'd100} : s = 119;
	{8'd19,8'd101} : s = 120;
	{8'd19,8'd102} : s = 121;
	{8'd19,8'd103} : s = 122;
	{8'd19,8'd104} : s = 123;
	{8'd19,8'd105} : s = 124;
	{8'd19,8'd106} : s = 125;
	{8'd19,8'd107} : s = 126;
	{8'd19,8'd108} : s = 127;
	{8'd19,8'd109} : s = 128;
	{8'd19,8'd110} : s = 129;
	{8'd19,8'd111} : s = 130;
	{8'd19,8'd112} : s = 131;
	{8'd19,8'd113} : s = 132;
	{8'd19,8'd114} : s = 133;
	{8'd19,8'd115} : s = 134;
	{8'd19,8'd116} : s = 135;
	{8'd19,8'd117} : s = 136;
	{8'd19,8'd118} : s = 137;
	{8'd19,8'd119} : s = 138;
	{8'd19,8'd120} : s = 139;
	{8'd19,8'd121} : s = 140;
	{8'd19,8'd122} : s = 141;
	{8'd19,8'd123} : s = 142;
	{8'd19,8'd124} : s = 143;
	{8'd19,8'd125} : s = 144;
	{8'd19,8'd126} : s = 145;
	{8'd19,8'd127} : s = 146;
	{8'd19,8'd128} : s = 147;
	{8'd19,8'd129} : s = 148;
	{8'd19,8'd130} : s = 149;
	{8'd19,8'd131} : s = 150;
	{8'd19,8'd132} : s = 151;
	{8'd19,8'd133} : s = 152;
	{8'd19,8'd134} : s = 153;
	{8'd19,8'd135} : s = 154;
	{8'd19,8'd136} : s = 155;
	{8'd19,8'd137} : s = 156;
	{8'd19,8'd138} : s = 157;
	{8'd19,8'd139} : s = 158;
	{8'd19,8'd140} : s = 159;
	{8'd19,8'd141} : s = 160;
	{8'd19,8'd142} : s = 161;
	{8'd19,8'd143} : s = 162;
	{8'd19,8'd144} : s = 163;
	{8'd19,8'd145} : s = 164;
	{8'd19,8'd146} : s = 165;
	{8'd19,8'd147} : s = 166;
	{8'd19,8'd148} : s = 167;
	{8'd19,8'd149} : s = 168;
	{8'd19,8'd150} : s = 169;
	{8'd19,8'd151} : s = 170;
	{8'd19,8'd152} : s = 171;
	{8'd19,8'd153} : s = 172;
	{8'd19,8'd154} : s = 173;
	{8'd19,8'd155} : s = 174;
	{8'd19,8'd156} : s = 175;
	{8'd19,8'd157} : s = 176;
	{8'd19,8'd158} : s = 177;
	{8'd19,8'd159} : s = 178;
	{8'd19,8'd160} : s = 179;
	{8'd19,8'd161} : s = 180;
	{8'd19,8'd162} : s = 181;
	{8'd19,8'd163} : s = 182;
	{8'd19,8'd164} : s = 183;
	{8'd19,8'd165} : s = 184;
	{8'd19,8'd166} : s = 185;
	{8'd19,8'd167} : s = 186;
	{8'd19,8'd168} : s = 187;
	{8'd19,8'd169} : s = 188;
	{8'd19,8'd170} : s = 189;
	{8'd19,8'd171} : s = 190;
	{8'd19,8'd172} : s = 191;
	{8'd19,8'd173} : s = 192;
	{8'd19,8'd174} : s = 193;
	{8'd19,8'd175} : s = 194;
	{8'd19,8'd176} : s = 195;
	{8'd19,8'd177} : s = 196;
	{8'd19,8'd178} : s = 197;
	{8'd19,8'd179} : s = 198;
	{8'd19,8'd180} : s = 199;
	{8'd19,8'd181} : s = 200;
	{8'd19,8'd182} : s = 201;
	{8'd19,8'd183} : s = 202;
	{8'd19,8'd184} : s = 203;
	{8'd19,8'd185} : s = 204;
	{8'd19,8'd186} : s = 205;
	{8'd19,8'd187} : s = 206;
	{8'd19,8'd188} : s = 207;
	{8'd19,8'd189} : s = 208;
	{8'd19,8'd190} : s = 209;
	{8'd19,8'd191} : s = 210;
	{8'd19,8'd192} : s = 211;
	{8'd19,8'd193} : s = 212;
	{8'd19,8'd194} : s = 213;
	{8'd19,8'd195} : s = 214;
	{8'd19,8'd196} : s = 215;
	{8'd19,8'd197} : s = 216;
	{8'd19,8'd198} : s = 217;
	{8'd19,8'd199} : s = 218;
	{8'd19,8'd200} : s = 219;
	{8'd19,8'd201} : s = 220;
	{8'd19,8'd202} : s = 221;
	{8'd19,8'd203} : s = 222;
	{8'd19,8'd204} : s = 223;
	{8'd19,8'd205} : s = 224;
	{8'd19,8'd206} : s = 225;
	{8'd19,8'd207} : s = 226;
	{8'd19,8'd208} : s = 227;
	{8'd19,8'd209} : s = 228;
	{8'd19,8'd210} : s = 229;
	{8'd19,8'd211} : s = 230;
	{8'd19,8'd212} : s = 231;
	{8'd19,8'd213} : s = 232;
	{8'd19,8'd214} : s = 233;
	{8'd19,8'd215} : s = 234;
	{8'd19,8'd216} : s = 235;
	{8'd19,8'd217} : s = 236;
	{8'd19,8'd218} : s = 237;
	{8'd19,8'd219} : s = 238;
	{8'd19,8'd220} : s = 239;
	{8'd19,8'd221} : s = 240;
	{8'd19,8'd222} : s = 241;
	{8'd19,8'd223} : s = 242;
	{8'd19,8'd224} : s = 243;
	{8'd19,8'd225} : s = 244;
	{8'd19,8'd226} : s = 245;
	{8'd19,8'd227} : s = 246;
	{8'd19,8'd228} : s = 247;
	{8'd19,8'd229} : s = 248;
	{8'd19,8'd230} : s = 249;
	{8'd19,8'd231} : s = 250;
	{8'd19,8'd232} : s = 251;
	{8'd19,8'd233} : s = 252;
	{8'd19,8'd234} : s = 253;
	{8'd19,8'd235} : s = 254;
	{8'd19,8'd236} : s = 255;
	{8'd19,8'd237} : s = 256;
	{8'd19,8'd238} : s = 257;
	{8'd19,8'd239} : s = 258;
	{8'd19,8'd240} : s = 259;
	{8'd19,8'd241} : s = 260;
	{8'd19,8'd242} : s = 261;
	{8'd19,8'd243} : s = 262;
	{8'd19,8'd244} : s = 263;
	{8'd19,8'd245} : s = 264;
	{8'd19,8'd246} : s = 265;
	{8'd19,8'd247} : s = 266;
	{8'd19,8'd248} : s = 267;
	{8'd19,8'd249} : s = 268;
	{8'd19,8'd250} : s = 269;
	{8'd19,8'd251} : s = 270;
	{8'd19,8'd252} : s = 271;
	{8'd19,8'd253} : s = 272;
	{8'd19,8'd254} : s = 273;
	{8'd19,8'd255} : s = 274;
	{8'd20,8'd0} : s = 20;
	{8'd20,8'd1} : s = 21;
	{8'd20,8'd2} : s = 22;
	{8'd20,8'd3} : s = 23;
	{8'd20,8'd4} : s = 24;
	{8'd20,8'd5} : s = 25;
	{8'd20,8'd6} : s = 26;
	{8'd20,8'd7} : s = 27;
	{8'd20,8'd8} : s = 28;
	{8'd20,8'd9} : s = 29;
	{8'd20,8'd10} : s = 30;
	{8'd20,8'd11} : s = 31;
	{8'd20,8'd12} : s = 32;
	{8'd20,8'd13} : s = 33;
	{8'd20,8'd14} : s = 34;
	{8'd20,8'd15} : s = 35;
	{8'd20,8'd16} : s = 36;
	{8'd20,8'd17} : s = 37;
	{8'd20,8'd18} : s = 38;
	{8'd20,8'd19} : s = 39;
	{8'd20,8'd20} : s = 40;
	{8'd20,8'd21} : s = 41;
	{8'd20,8'd22} : s = 42;
	{8'd20,8'd23} : s = 43;
	{8'd20,8'd24} : s = 44;
	{8'd20,8'd25} : s = 45;
	{8'd20,8'd26} : s = 46;
	{8'd20,8'd27} : s = 47;
	{8'd20,8'd28} : s = 48;
	{8'd20,8'd29} : s = 49;
	{8'd20,8'd30} : s = 50;
	{8'd20,8'd31} : s = 51;
	{8'd20,8'd32} : s = 52;
	{8'd20,8'd33} : s = 53;
	{8'd20,8'd34} : s = 54;
	{8'd20,8'd35} : s = 55;
	{8'd20,8'd36} : s = 56;
	{8'd20,8'd37} : s = 57;
	{8'd20,8'd38} : s = 58;
	{8'd20,8'd39} : s = 59;
	{8'd20,8'd40} : s = 60;
	{8'd20,8'd41} : s = 61;
	{8'd20,8'd42} : s = 62;
	{8'd20,8'd43} : s = 63;
	{8'd20,8'd44} : s = 64;
	{8'd20,8'd45} : s = 65;
	{8'd20,8'd46} : s = 66;
	{8'd20,8'd47} : s = 67;
	{8'd20,8'd48} : s = 68;
	{8'd20,8'd49} : s = 69;
	{8'd20,8'd50} : s = 70;
	{8'd20,8'd51} : s = 71;
	{8'd20,8'd52} : s = 72;
	{8'd20,8'd53} : s = 73;
	{8'd20,8'd54} : s = 74;
	{8'd20,8'd55} : s = 75;
	{8'd20,8'd56} : s = 76;
	{8'd20,8'd57} : s = 77;
	{8'd20,8'd58} : s = 78;
	{8'd20,8'd59} : s = 79;
	{8'd20,8'd60} : s = 80;
	{8'd20,8'd61} : s = 81;
	{8'd20,8'd62} : s = 82;
	{8'd20,8'd63} : s = 83;
	{8'd20,8'd64} : s = 84;
	{8'd20,8'd65} : s = 85;
	{8'd20,8'd66} : s = 86;
	{8'd20,8'd67} : s = 87;
	{8'd20,8'd68} : s = 88;
	{8'd20,8'd69} : s = 89;
	{8'd20,8'd70} : s = 90;
	{8'd20,8'd71} : s = 91;
	{8'd20,8'd72} : s = 92;
	{8'd20,8'd73} : s = 93;
	{8'd20,8'd74} : s = 94;
	{8'd20,8'd75} : s = 95;
	{8'd20,8'd76} : s = 96;
	{8'd20,8'd77} : s = 97;
	{8'd20,8'd78} : s = 98;
	{8'd20,8'd79} : s = 99;
	{8'd20,8'd80} : s = 100;
	{8'd20,8'd81} : s = 101;
	{8'd20,8'd82} : s = 102;
	{8'd20,8'd83} : s = 103;
	{8'd20,8'd84} : s = 104;
	{8'd20,8'd85} : s = 105;
	{8'd20,8'd86} : s = 106;
	{8'd20,8'd87} : s = 107;
	{8'd20,8'd88} : s = 108;
	{8'd20,8'd89} : s = 109;
	{8'd20,8'd90} : s = 110;
	{8'd20,8'd91} : s = 111;
	{8'd20,8'd92} : s = 112;
	{8'd20,8'd93} : s = 113;
	{8'd20,8'd94} : s = 114;
	{8'd20,8'd95} : s = 115;
	{8'd20,8'd96} : s = 116;
	{8'd20,8'd97} : s = 117;
	{8'd20,8'd98} : s = 118;
	{8'd20,8'd99} : s = 119;
	{8'd20,8'd100} : s = 120;
	{8'd20,8'd101} : s = 121;
	{8'd20,8'd102} : s = 122;
	{8'd20,8'd103} : s = 123;
	{8'd20,8'd104} : s = 124;
	{8'd20,8'd105} : s = 125;
	{8'd20,8'd106} : s = 126;
	{8'd20,8'd107} : s = 127;
	{8'd20,8'd108} : s = 128;
	{8'd20,8'd109} : s = 129;
	{8'd20,8'd110} : s = 130;
	{8'd20,8'd111} : s = 131;
	{8'd20,8'd112} : s = 132;
	{8'd20,8'd113} : s = 133;
	{8'd20,8'd114} : s = 134;
	{8'd20,8'd115} : s = 135;
	{8'd20,8'd116} : s = 136;
	{8'd20,8'd117} : s = 137;
	{8'd20,8'd118} : s = 138;
	{8'd20,8'd119} : s = 139;
	{8'd20,8'd120} : s = 140;
	{8'd20,8'd121} : s = 141;
	{8'd20,8'd122} : s = 142;
	{8'd20,8'd123} : s = 143;
	{8'd20,8'd124} : s = 144;
	{8'd20,8'd125} : s = 145;
	{8'd20,8'd126} : s = 146;
	{8'd20,8'd127} : s = 147;
	{8'd20,8'd128} : s = 148;
	{8'd20,8'd129} : s = 149;
	{8'd20,8'd130} : s = 150;
	{8'd20,8'd131} : s = 151;
	{8'd20,8'd132} : s = 152;
	{8'd20,8'd133} : s = 153;
	{8'd20,8'd134} : s = 154;
	{8'd20,8'd135} : s = 155;
	{8'd20,8'd136} : s = 156;
	{8'd20,8'd137} : s = 157;
	{8'd20,8'd138} : s = 158;
	{8'd20,8'd139} : s = 159;
	{8'd20,8'd140} : s = 160;
	{8'd20,8'd141} : s = 161;
	{8'd20,8'd142} : s = 162;
	{8'd20,8'd143} : s = 163;
	{8'd20,8'd144} : s = 164;
	{8'd20,8'd145} : s = 165;
	{8'd20,8'd146} : s = 166;
	{8'd20,8'd147} : s = 167;
	{8'd20,8'd148} : s = 168;
	{8'd20,8'd149} : s = 169;
	{8'd20,8'd150} : s = 170;
	{8'd20,8'd151} : s = 171;
	{8'd20,8'd152} : s = 172;
	{8'd20,8'd153} : s = 173;
	{8'd20,8'd154} : s = 174;
	{8'd20,8'd155} : s = 175;
	{8'd20,8'd156} : s = 176;
	{8'd20,8'd157} : s = 177;
	{8'd20,8'd158} : s = 178;
	{8'd20,8'd159} : s = 179;
	{8'd20,8'd160} : s = 180;
	{8'd20,8'd161} : s = 181;
	{8'd20,8'd162} : s = 182;
	{8'd20,8'd163} : s = 183;
	{8'd20,8'd164} : s = 184;
	{8'd20,8'd165} : s = 185;
	{8'd20,8'd166} : s = 186;
	{8'd20,8'd167} : s = 187;
	{8'd20,8'd168} : s = 188;
	{8'd20,8'd169} : s = 189;
	{8'd20,8'd170} : s = 190;
	{8'd20,8'd171} : s = 191;
	{8'd20,8'd172} : s = 192;
	{8'd20,8'd173} : s = 193;
	{8'd20,8'd174} : s = 194;
	{8'd20,8'd175} : s = 195;
	{8'd20,8'd176} : s = 196;
	{8'd20,8'd177} : s = 197;
	{8'd20,8'd178} : s = 198;
	{8'd20,8'd179} : s = 199;
	{8'd20,8'd180} : s = 200;
	{8'd20,8'd181} : s = 201;
	{8'd20,8'd182} : s = 202;
	{8'd20,8'd183} : s = 203;
	{8'd20,8'd184} : s = 204;
	{8'd20,8'd185} : s = 205;
	{8'd20,8'd186} : s = 206;
	{8'd20,8'd187} : s = 207;
	{8'd20,8'd188} : s = 208;
	{8'd20,8'd189} : s = 209;
	{8'd20,8'd190} : s = 210;
	{8'd20,8'd191} : s = 211;
	{8'd20,8'd192} : s = 212;
	{8'd20,8'd193} : s = 213;
	{8'd20,8'd194} : s = 214;
	{8'd20,8'd195} : s = 215;
	{8'd20,8'd196} : s = 216;
	{8'd20,8'd197} : s = 217;
	{8'd20,8'd198} : s = 218;
	{8'd20,8'd199} : s = 219;
	{8'd20,8'd200} : s = 220;
	{8'd20,8'd201} : s = 221;
	{8'd20,8'd202} : s = 222;
	{8'd20,8'd203} : s = 223;
	{8'd20,8'd204} : s = 224;
	{8'd20,8'd205} : s = 225;
	{8'd20,8'd206} : s = 226;
	{8'd20,8'd207} : s = 227;
	{8'd20,8'd208} : s = 228;
	{8'd20,8'd209} : s = 229;
	{8'd20,8'd210} : s = 230;
	{8'd20,8'd211} : s = 231;
	{8'd20,8'd212} : s = 232;
	{8'd20,8'd213} : s = 233;
	{8'd20,8'd214} : s = 234;
	{8'd20,8'd215} : s = 235;
	{8'd20,8'd216} : s = 236;
	{8'd20,8'd217} : s = 237;
	{8'd20,8'd218} : s = 238;
	{8'd20,8'd219} : s = 239;
	{8'd20,8'd220} : s = 240;
	{8'd20,8'd221} : s = 241;
	{8'd20,8'd222} : s = 242;
	{8'd20,8'd223} : s = 243;
	{8'd20,8'd224} : s = 244;
	{8'd20,8'd225} : s = 245;
	{8'd20,8'd226} : s = 246;
	{8'd20,8'd227} : s = 247;
	{8'd20,8'd228} : s = 248;
	{8'd20,8'd229} : s = 249;
	{8'd20,8'd230} : s = 250;
	{8'd20,8'd231} : s = 251;
	{8'd20,8'd232} : s = 252;
	{8'd20,8'd233} : s = 253;
	{8'd20,8'd234} : s = 254;
	{8'd20,8'd235} : s = 255;
	{8'd20,8'd236} : s = 256;
	{8'd20,8'd237} : s = 257;
	{8'd20,8'd238} : s = 258;
	{8'd20,8'd239} : s = 259;
	{8'd20,8'd240} : s = 260;
	{8'd20,8'd241} : s = 261;
	{8'd20,8'd242} : s = 262;
	{8'd20,8'd243} : s = 263;
	{8'd20,8'd244} : s = 264;
	{8'd20,8'd245} : s = 265;
	{8'd20,8'd246} : s = 266;
	{8'd20,8'd247} : s = 267;
	{8'd20,8'd248} : s = 268;
	{8'd20,8'd249} : s = 269;
	{8'd20,8'd250} : s = 270;
	{8'd20,8'd251} : s = 271;
	{8'd20,8'd252} : s = 272;
	{8'd20,8'd253} : s = 273;
	{8'd20,8'd254} : s = 274;
	{8'd20,8'd255} : s = 275;
	{8'd21,8'd0} : s = 21;
	{8'd21,8'd1} : s = 22;
	{8'd21,8'd2} : s = 23;
	{8'd21,8'd3} : s = 24;
	{8'd21,8'd4} : s = 25;
	{8'd21,8'd5} : s = 26;
	{8'd21,8'd6} : s = 27;
	{8'd21,8'd7} : s = 28;
	{8'd21,8'd8} : s = 29;
	{8'd21,8'd9} : s = 30;
	{8'd21,8'd10} : s = 31;
	{8'd21,8'd11} : s = 32;
	{8'd21,8'd12} : s = 33;
	{8'd21,8'd13} : s = 34;
	{8'd21,8'd14} : s = 35;
	{8'd21,8'd15} : s = 36;
	{8'd21,8'd16} : s = 37;
	{8'd21,8'd17} : s = 38;
	{8'd21,8'd18} : s = 39;
	{8'd21,8'd19} : s = 40;
	{8'd21,8'd20} : s = 41;
	{8'd21,8'd21} : s = 42;
	{8'd21,8'd22} : s = 43;
	{8'd21,8'd23} : s = 44;
	{8'd21,8'd24} : s = 45;
	{8'd21,8'd25} : s = 46;
	{8'd21,8'd26} : s = 47;
	{8'd21,8'd27} : s = 48;
	{8'd21,8'd28} : s = 49;
	{8'd21,8'd29} : s = 50;
	{8'd21,8'd30} : s = 51;
	{8'd21,8'd31} : s = 52;
	{8'd21,8'd32} : s = 53;
	{8'd21,8'd33} : s = 54;
	{8'd21,8'd34} : s = 55;
	{8'd21,8'd35} : s = 56;
	{8'd21,8'd36} : s = 57;
	{8'd21,8'd37} : s = 58;
	{8'd21,8'd38} : s = 59;
	{8'd21,8'd39} : s = 60;
	{8'd21,8'd40} : s = 61;
	{8'd21,8'd41} : s = 62;
	{8'd21,8'd42} : s = 63;
	{8'd21,8'd43} : s = 64;
	{8'd21,8'd44} : s = 65;
	{8'd21,8'd45} : s = 66;
	{8'd21,8'd46} : s = 67;
	{8'd21,8'd47} : s = 68;
	{8'd21,8'd48} : s = 69;
	{8'd21,8'd49} : s = 70;
	{8'd21,8'd50} : s = 71;
	{8'd21,8'd51} : s = 72;
	{8'd21,8'd52} : s = 73;
	{8'd21,8'd53} : s = 74;
	{8'd21,8'd54} : s = 75;
	{8'd21,8'd55} : s = 76;
	{8'd21,8'd56} : s = 77;
	{8'd21,8'd57} : s = 78;
	{8'd21,8'd58} : s = 79;
	{8'd21,8'd59} : s = 80;
	{8'd21,8'd60} : s = 81;
	{8'd21,8'd61} : s = 82;
	{8'd21,8'd62} : s = 83;
	{8'd21,8'd63} : s = 84;
	{8'd21,8'd64} : s = 85;
	{8'd21,8'd65} : s = 86;
	{8'd21,8'd66} : s = 87;
	{8'd21,8'd67} : s = 88;
	{8'd21,8'd68} : s = 89;
	{8'd21,8'd69} : s = 90;
	{8'd21,8'd70} : s = 91;
	{8'd21,8'd71} : s = 92;
	{8'd21,8'd72} : s = 93;
	{8'd21,8'd73} : s = 94;
	{8'd21,8'd74} : s = 95;
	{8'd21,8'd75} : s = 96;
	{8'd21,8'd76} : s = 97;
	{8'd21,8'd77} : s = 98;
	{8'd21,8'd78} : s = 99;
	{8'd21,8'd79} : s = 100;
	{8'd21,8'd80} : s = 101;
	{8'd21,8'd81} : s = 102;
	{8'd21,8'd82} : s = 103;
	{8'd21,8'd83} : s = 104;
	{8'd21,8'd84} : s = 105;
	{8'd21,8'd85} : s = 106;
	{8'd21,8'd86} : s = 107;
	{8'd21,8'd87} : s = 108;
	{8'd21,8'd88} : s = 109;
	{8'd21,8'd89} : s = 110;
	{8'd21,8'd90} : s = 111;
	{8'd21,8'd91} : s = 112;
	{8'd21,8'd92} : s = 113;
	{8'd21,8'd93} : s = 114;
	{8'd21,8'd94} : s = 115;
	{8'd21,8'd95} : s = 116;
	{8'd21,8'd96} : s = 117;
	{8'd21,8'd97} : s = 118;
	{8'd21,8'd98} : s = 119;
	{8'd21,8'd99} : s = 120;
	{8'd21,8'd100} : s = 121;
	{8'd21,8'd101} : s = 122;
	{8'd21,8'd102} : s = 123;
	{8'd21,8'd103} : s = 124;
	{8'd21,8'd104} : s = 125;
	{8'd21,8'd105} : s = 126;
	{8'd21,8'd106} : s = 127;
	{8'd21,8'd107} : s = 128;
	{8'd21,8'd108} : s = 129;
	{8'd21,8'd109} : s = 130;
	{8'd21,8'd110} : s = 131;
	{8'd21,8'd111} : s = 132;
	{8'd21,8'd112} : s = 133;
	{8'd21,8'd113} : s = 134;
	{8'd21,8'd114} : s = 135;
	{8'd21,8'd115} : s = 136;
	{8'd21,8'd116} : s = 137;
	{8'd21,8'd117} : s = 138;
	{8'd21,8'd118} : s = 139;
	{8'd21,8'd119} : s = 140;
	{8'd21,8'd120} : s = 141;
	{8'd21,8'd121} : s = 142;
	{8'd21,8'd122} : s = 143;
	{8'd21,8'd123} : s = 144;
	{8'd21,8'd124} : s = 145;
	{8'd21,8'd125} : s = 146;
	{8'd21,8'd126} : s = 147;
	{8'd21,8'd127} : s = 148;
	{8'd21,8'd128} : s = 149;
	{8'd21,8'd129} : s = 150;
	{8'd21,8'd130} : s = 151;
	{8'd21,8'd131} : s = 152;
	{8'd21,8'd132} : s = 153;
	{8'd21,8'd133} : s = 154;
	{8'd21,8'd134} : s = 155;
	{8'd21,8'd135} : s = 156;
	{8'd21,8'd136} : s = 157;
	{8'd21,8'd137} : s = 158;
	{8'd21,8'd138} : s = 159;
	{8'd21,8'd139} : s = 160;
	{8'd21,8'd140} : s = 161;
	{8'd21,8'd141} : s = 162;
	{8'd21,8'd142} : s = 163;
	{8'd21,8'd143} : s = 164;
	{8'd21,8'd144} : s = 165;
	{8'd21,8'd145} : s = 166;
	{8'd21,8'd146} : s = 167;
	{8'd21,8'd147} : s = 168;
	{8'd21,8'd148} : s = 169;
	{8'd21,8'd149} : s = 170;
	{8'd21,8'd150} : s = 171;
	{8'd21,8'd151} : s = 172;
	{8'd21,8'd152} : s = 173;
	{8'd21,8'd153} : s = 174;
	{8'd21,8'd154} : s = 175;
	{8'd21,8'd155} : s = 176;
	{8'd21,8'd156} : s = 177;
	{8'd21,8'd157} : s = 178;
	{8'd21,8'd158} : s = 179;
	{8'd21,8'd159} : s = 180;
	{8'd21,8'd160} : s = 181;
	{8'd21,8'd161} : s = 182;
	{8'd21,8'd162} : s = 183;
	{8'd21,8'd163} : s = 184;
	{8'd21,8'd164} : s = 185;
	{8'd21,8'd165} : s = 186;
	{8'd21,8'd166} : s = 187;
	{8'd21,8'd167} : s = 188;
	{8'd21,8'd168} : s = 189;
	{8'd21,8'd169} : s = 190;
	{8'd21,8'd170} : s = 191;
	{8'd21,8'd171} : s = 192;
	{8'd21,8'd172} : s = 193;
	{8'd21,8'd173} : s = 194;
	{8'd21,8'd174} : s = 195;
	{8'd21,8'd175} : s = 196;
	{8'd21,8'd176} : s = 197;
	{8'd21,8'd177} : s = 198;
	{8'd21,8'd178} : s = 199;
	{8'd21,8'd179} : s = 200;
	{8'd21,8'd180} : s = 201;
	{8'd21,8'd181} : s = 202;
	{8'd21,8'd182} : s = 203;
	{8'd21,8'd183} : s = 204;
	{8'd21,8'd184} : s = 205;
	{8'd21,8'd185} : s = 206;
	{8'd21,8'd186} : s = 207;
	{8'd21,8'd187} : s = 208;
	{8'd21,8'd188} : s = 209;
	{8'd21,8'd189} : s = 210;
	{8'd21,8'd190} : s = 211;
	{8'd21,8'd191} : s = 212;
	{8'd21,8'd192} : s = 213;
	{8'd21,8'd193} : s = 214;
	{8'd21,8'd194} : s = 215;
	{8'd21,8'd195} : s = 216;
	{8'd21,8'd196} : s = 217;
	{8'd21,8'd197} : s = 218;
	{8'd21,8'd198} : s = 219;
	{8'd21,8'd199} : s = 220;
	{8'd21,8'd200} : s = 221;
	{8'd21,8'd201} : s = 222;
	{8'd21,8'd202} : s = 223;
	{8'd21,8'd203} : s = 224;
	{8'd21,8'd204} : s = 225;
	{8'd21,8'd205} : s = 226;
	{8'd21,8'd206} : s = 227;
	{8'd21,8'd207} : s = 228;
	{8'd21,8'd208} : s = 229;
	{8'd21,8'd209} : s = 230;
	{8'd21,8'd210} : s = 231;
	{8'd21,8'd211} : s = 232;
	{8'd21,8'd212} : s = 233;
	{8'd21,8'd213} : s = 234;
	{8'd21,8'd214} : s = 235;
	{8'd21,8'd215} : s = 236;
	{8'd21,8'd216} : s = 237;
	{8'd21,8'd217} : s = 238;
	{8'd21,8'd218} : s = 239;
	{8'd21,8'd219} : s = 240;
	{8'd21,8'd220} : s = 241;
	{8'd21,8'd221} : s = 242;
	{8'd21,8'd222} : s = 243;
	{8'd21,8'd223} : s = 244;
	{8'd21,8'd224} : s = 245;
	{8'd21,8'd225} : s = 246;
	{8'd21,8'd226} : s = 247;
	{8'd21,8'd227} : s = 248;
	{8'd21,8'd228} : s = 249;
	{8'd21,8'd229} : s = 250;
	{8'd21,8'd230} : s = 251;
	{8'd21,8'd231} : s = 252;
	{8'd21,8'd232} : s = 253;
	{8'd21,8'd233} : s = 254;
	{8'd21,8'd234} : s = 255;
	{8'd21,8'd235} : s = 256;
	{8'd21,8'd236} : s = 257;
	{8'd21,8'd237} : s = 258;
	{8'd21,8'd238} : s = 259;
	{8'd21,8'd239} : s = 260;
	{8'd21,8'd240} : s = 261;
	{8'd21,8'd241} : s = 262;
	{8'd21,8'd242} : s = 263;
	{8'd21,8'd243} : s = 264;
	{8'd21,8'd244} : s = 265;
	{8'd21,8'd245} : s = 266;
	{8'd21,8'd246} : s = 267;
	{8'd21,8'd247} : s = 268;
	{8'd21,8'd248} : s = 269;
	{8'd21,8'd249} : s = 270;
	{8'd21,8'd250} : s = 271;
	{8'd21,8'd251} : s = 272;
	{8'd21,8'd252} : s = 273;
	{8'd21,8'd253} : s = 274;
	{8'd21,8'd254} : s = 275;
	{8'd21,8'd255} : s = 276;
	{8'd22,8'd0} : s = 22;
	{8'd22,8'd1} : s = 23;
	{8'd22,8'd2} : s = 24;
	{8'd22,8'd3} : s = 25;
	{8'd22,8'd4} : s = 26;
	{8'd22,8'd5} : s = 27;
	{8'd22,8'd6} : s = 28;
	{8'd22,8'd7} : s = 29;
	{8'd22,8'd8} : s = 30;
	{8'd22,8'd9} : s = 31;
	{8'd22,8'd10} : s = 32;
	{8'd22,8'd11} : s = 33;
	{8'd22,8'd12} : s = 34;
	{8'd22,8'd13} : s = 35;
	{8'd22,8'd14} : s = 36;
	{8'd22,8'd15} : s = 37;
	{8'd22,8'd16} : s = 38;
	{8'd22,8'd17} : s = 39;
	{8'd22,8'd18} : s = 40;
	{8'd22,8'd19} : s = 41;
	{8'd22,8'd20} : s = 42;
	{8'd22,8'd21} : s = 43;
	{8'd22,8'd22} : s = 44;
	{8'd22,8'd23} : s = 45;
	{8'd22,8'd24} : s = 46;
	{8'd22,8'd25} : s = 47;
	{8'd22,8'd26} : s = 48;
	{8'd22,8'd27} : s = 49;
	{8'd22,8'd28} : s = 50;
	{8'd22,8'd29} : s = 51;
	{8'd22,8'd30} : s = 52;
	{8'd22,8'd31} : s = 53;
	{8'd22,8'd32} : s = 54;
	{8'd22,8'd33} : s = 55;
	{8'd22,8'd34} : s = 56;
	{8'd22,8'd35} : s = 57;
	{8'd22,8'd36} : s = 58;
	{8'd22,8'd37} : s = 59;
	{8'd22,8'd38} : s = 60;
	{8'd22,8'd39} : s = 61;
	{8'd22,8'd40} : s = 62;
	{8'd22,8'd41} : s = 63;
	{8'd22,8'd42} : s = 64;
	{8'd22,8'd43} : s = 65;
	{8'd22,8'd44} : s = 66;
	{8'd22,8'd45} : s = 67;
	{8'd22,8'd46} : s = 68;
	{8'd22,8'd47} : s = 69;
	{8'd22,8'd48} : s = 70;
	{8'd22,8'd49} : s = 71;
	{8'd22,8'd50} : s = 72;
	{8'd22,8'd51} : s = 73;
	{8'd22,8'd52} : s = 74;
	{8'd22,8'd53} : s = 75;
	{8'd22,8'd54} : s = 76;
	{8'd22,8'd55} : s = 77;
	{8'd22,8'd56} : s = 78;
	{8'd22,8'd57} : s = 79;
	{8'd22,8'd58} : s = 80;
	{8'd22,8'd59} : s = 81;
	{8'd22,8'd60} : s = 82;
	{8'd22,8'd61} : s = 83;
	{8'd22,8'd62} : s = 84;
	{8'd22,8'd63} : s = 85;
	{8'd22,8'd64} : s = 86;
	{8'd22,8'd65} : s = 87;
	{8'd22,8'd66} : s = 88;
	{8'd22,8'd67} : s = 89;
	{8'd22,8'd68} : s = 90;
	{8'd22,8'd69} : s = 91;
	{8'd22,8'd70} : s = 92;
	{8'd22,8'd71} : s = 93;
	{8'd22,8'd72} : s = 94;
	{8'd22,8'd73} : s = 95;
	{8'd22,8'd74} : s = 96;
	{8'd22,8'd75} : s = 97;
	{8'd22,8'd76} : s = 98;
	{8'd22,8'd77} : s = 99;
	{8'd22,8'd78} : s = 100;
	{8'd22,8'd79} : s = 101;
	{8'd22,8'd80} : s = 102;
	{8'd22,8'd81} : s = 103;
	{8'd22,8'd82} : s = 104;
	{8'd22,8'd83} : s = 105;
	{8'd22,8'd84} : s = 106;
	{8'd22,8'd85} : s = 107;
	{8'd22,8'd86} : s = 108;
	{8'd22,8'd87} : s = 109;
	{8'd22,8'd88} : s = 110;
	{8'd22,8'd89} : s = 111;
	{8'd22,8'd90} : s = 112;
	{8'd22,8'd91} : s = 113;
	{8'd22,8'd92} : s = 114;
	{8'd22,8'd93} : s = 115;
	{8'd22,8'd94} : s = 116;
	{8'd22,8'd95} : s = 117;
	{8'd22,8'd96} : s = 118;
	{8'd22,8'd97} : s = 119;
	{8'd22,8'd98} : s = 120;
	{8'd22,8'd99} : s = 121;
	{8'd22,8'd100} : s = 122;
	{8'd22,8'd101} : s = 123;
	{8'd22,8'd102} : s = 124;
	{8'd22,8'd103} : s = 125;
	{8'd22,8'd104} : s = 126;
	{8'd22,8'd105} : s = 127;
	{8'd22,8'd106} : s = 128;
	{8'd22,8'd107} : s = 129;
	{8'd22,8'd108} : s = 130;
	{8'd22,8'd109} : s = 131;
	{8'd22,8'd110} : s = 132;
	{8'd22,8'd111} : s = 133;
	{8'd22,8'd112} : s = 134;
	{8'd22,8'd113} : s = 135;
	{8'd22,8'd114} : s = 136;
	{8'd22,8'd115} : s = 137;
	{8'd22,8'd116} : s = 138;
	{8'd22,8'd117} : s = 139;
	{8'd22,8'd118} : s = 140;
	{8'd22,8'd119} : s = 141;
	{8'd22,8'd120} : s = 142;
	{8'd22,8'd121} : s = 143;
	{8'd22,8'd122} : s = 144;
	{8'd22,8'd123} : s = 145;
	{8'd22,8'd124} : s = 146;
	{8'd22,8'd125} : s = 147;
	{8'd22,8'd126} : s = 148;
	{8'd22,8'd127} : s = 149;
	{8'd22,8'd128} : s = 150;
	{8'd22,8'd129} : s = 151;
	{8'd22,8'd130} : s = 152;
	{8'd22,8'd131} : s = 153;
	{8'd22,8'd132} : s = 154;
	{8'd22,8'd133} : s = 155;
	{8'd22,8'd134} : s = 156;
	{8'd22,8'd135} : s = 157;
	{8'd22,8'd136} : s = 158;
	{8'd22,8'd137} : s = 159;
	{8'd22,8'd138} : s = 160;
	{8'd22,8'd139} : s = 161;
	{8'd22,8'd140} : s = 162;
	{8'd22,8'd141} : s = 163;
	{8'd22,8'd142} : s = 164;
	{8'd22,8'd143} : s = 165;
	{8'd22,8'd144} : s = 166;
	{8'd22,8'd145} : s = 167;
	{8'd22,8'd146} : s = 168;
	{8'd22,8'd147} : s = 169;
	{8'd22,8'd148} : s = 170;
	{8'd22,8'd149} : s = 171;
	{8'd22,8'd150} : s = 172;
	{8'd22,8'd151} : s = 173;
	{8'd22,8'd152} : s = 174;
	{8'd22,8'd153} : s = 175;
	{8'd22,8'd154} : s = 176;
	{8'd22,8'd155} : s = 177;
	{8'd22,8'd156} : s = 178;
	{8'd22,8'd157} : s = 179;
	{8'd22,8'd158} : s = 180;
	{8'd22,8'd159} : s = 181;
	{8'd22,8'd160} : s = 182;
	{8'd22,8'd161} : s = 183;
	{8'd22,8'd162} : s = 184;
	{8'd22,8'd163} : s = 185;
	{8'd22,8'd164} : s = 186;
	{8'd22,8'd165} : s = 187;
	{8'd22,8'd166} : s = 188;
	{8'd22,8'd167} : s = 189;
	{8'd22,8'd168} : s = 190;
	{8'd22,8'd169} : s = 191;
	{8'd22,8'd170} : s = 192;
	{8'd22,8'd171} : s = 193;
	{8'd22,8'd172} : s = 194;
	{8'd22,8'd173} : s = 195;
	{8'd22,8'd174} : s = 196;
	{8'd22,8'd175} : s = 197;
	{8'd22,8'd176} : s = 198;
	{8'd22,8'd177} : s = 199;
	{8'd22,8'd178} : s = 200;
	{8'd22,8'd179} : s = 201;
	{8'd22,8'd180} : s = 202;
	{8'd22,8'd181} : s = 203;
	{8'd22,8'd182} : s = 204;
	{8'd22,8'd183} : s = 205;
	{8'd22,8'd184} : s = 206;
	{8'd22,8'd185} : s = 207;
	{8'd22,8'd186} : s = 208;
	{8'd22,8'd187} : s = 209;
	{8'd22,8'd188} : s = 210;
	{8'd22,8'd189} : s = 211;
	{8'd22,8'd190} : s = 212;
	{8'd22,8'd191} : s = 213;
	{8'd22,8'd192} : s = 214;
	{8'd22,8'd193} : s = 215;
	{8'd22,8'd194} : s = 216;
	{8'd22,8'd195} : s = 217;
	{8'd22,8'd196} : s = 218;
	{8'd22,8'd197} : s = 219;
	{8'd22,8'd198} : s = 220;
	{8'd22,8'd199} : s = 221;
	{8'd22,8'd200} : s = 222;
	{8'd22,8'd201} : s = 223;
	{8'd22,8'd202} : s = 224;
	{8'd22,8'd203} : s = 225;
	{8'd22,8'd204} : s = 226;
	{8'd22,8'd205} : s = 227;
	{8'd22,8'd206} : s = 228;
	{8'd22,8'd207} : s = 229;
	{8'd22,8'd208} : s = 230;
	{8'd22,8'd209} : s = 231;
	{8'd22,8'd210} : s = 232;
	{8'd22,8'd211} : s = 233;
	{8'd22,8'd212} : s = 234;
	{8'd22,8'd213} : s = 235;
	{8'd22,8'd214} : s = 236;
	{8'd22,8'd215} : s = 237;
	{8'd22,8'd216} : s = 238;
	{8'd22,8'd217} : s = 239;
	{8'd22,8'd218} : s = 240;
	{8'd22,8'd219} : s = 241;
	{8'd22,8'd220} : s = 242;
	{8'd22,8'd221} : s = 243;
	{8'd22,8'd222} : s = 244;
	{8'd22,8'd223} : s = 245;
	{8'd22,8'd224} : s = 246;
	{8'd22,8'd225} : s = 247;
	{8'd22,8'd226} : s = 248;
	{8'd22,8'd227} : s = 249;
	{8'd22,8'd228} : s = 250;
	{8'd22,8'd229} : s = 251;
	{8'd22,8'd230} : s = 252;
	{8'd22,8'd231} : s = 253;
	{8'd22,8'd232} : s = 254;
	{8'd22,8'd233} : s = 255;
	{8'd22,8'd234} : s = 256;
	{8'd22,8'd235} : s = 257;
	{8'd22,8'd236} : s = 258;
	{8'd22,8'd237} : s = 259;
	{8'd22,8'd238} : s = 260;
	{8'd22,8'd239} : s = 261;
	{8'd22,8'd240} : s = 262;
	{8'd22,8'd241} : s = 263;
	{8'd22,8'd242} : s = 264;
	{8'd22,8'd243} : s = 265;
	{8'd22,8'd244} : s = 266;
	{8'd22,8'd245} : s = 267;
	{8'd22,8'd246} : s = 268;
	{8'd22,8'd247} : s = 269;
	{8'd22,8'd248} : s = 270;
	{8'd22,8'd249} : s = 271;
	{8'd22,8'd250} : s = 272;
	{8'd22,8'd251} : s = 273;
	{8'd22,8'd252} : s = 274;
	{8'd22,8'd253} : s = 275;
	{8'd22,8'd254} : s = 276;
	{8'd22,8'd255} : s = 277;
	{8'd23,8'd0} : s = 23;
	{8'd23,8'd1} : s = 24;
	{8'd23,8'd2} : s = 25;
	{8'd23,8'd3} : s = 26;
	{8'd23,8'd4} : s = 27;
	{8'd23,8'd5} : s = 28;
	{8'd23,8'd6} : s = 29;
	{8'd23,8'd7} : s = 30;
	{8'd23,8'd8} : s = 31;
	{8'd23,8'd9} : s = 32;
	{8'd23,8'd10} : s = 33;
	{8'd23,8'd11} : s = 34;
	{8'd23,8'd12} : s = 35;
	{8'd23,8'd13} : s = 36;
	{8'd23,8'd14} : s = 37;
	{8'd23,8'd15} : s = 38;
	{8'd23,8'd16} : s = 39;
	{8'd23,8'd17} : s = 40;
	{8'd23,8'd18} : s = 41;
	{8'd23,8'd19} : s = 42;
	{8'd23,8'd20} : s = 43;
	{8'd23,8'd21} : s = 44;
	{8'd23,8'd22} : s = 45;
	{8'd23,8'd23} : s = 46;
	{8'd23,8'd24} : s = 47;
	{8'd23,8'd25} : s = 48;
	{8'd23,8'd26} : s = 49;
	{8'd23,8'd27} : s = 50;
	{8'd23,8'd28} : s = 51;
	{8'd23,8'd29} : s = 52;
	{8'd23,8'd30} : s = 53;
	{8'd23,8'd31} : s = 54;
	{8'd23,8'd32} : s = 55;
	{8'd23,8'd33} : s = 56;
	{8'd23,8'd34} : s = 57;
	{8'd23,8'd35} : s = 58;
	{8'd23,8'd36} : s = 59;
	{8'd23,8'd37} : s = 60;
	{8'd23,8'd38} : s = 61;
	{8'd23,8'd39} : s = 62;
	{8'd23,8'd40} : s = 63;
	{8'd23,8'd41} : s = 64;
	{8'd23,8'd42} : s = 65;
	{8'd23,8'd43} : s = 66;
	{8'd23,8'd44} : s = 67;
	{8'd23,8'd45} : s = 68;
	{8'd23,8'd46} : s = 69;
	{8'd23,8'd47} : s = 70;
	{8'd23,8'd48} : s = 71;
	{8'd23,8'd49} : s = 72;
	{8'd23,8'd50} : s = 73;
	{8'd23,8'd51} : s = 74;
	{8'd23,8'd52} : s = 75;
	{8'd23,8'd53} : s = 76;
	{8'd23,8'd54} : s = 77;
	{8'd23,8'd55} : s = 78;
	{8'd23,8'd56} : s = 79;
	{8'd23,8'd57} : s = 80;
	{8'd23,8'd58} : s = 81;
	{8'd23,8'd59} : s = 82;
	{8'd23,8'd60} : s = 83;
	{8'd23,8'd61} : s = 84;
	{8'd23,8'd62} : s = 85;
	{8'd23,8'd63} : s = 86;
	{8'd23,8'd64} : s = 87;
	{8'd23,8'd65} : s = 88;
	{8'd23,8'd66} : s = 89;
	{8'd23,8'd67} : s = 90;
	{8'd23,8'd68} : s = 91;
	{8'd23,8'd69} : s = 92;
	{8'd23,8'd70} : s = 93;
	{8'd23,8'd71} : s = 94;
	{8'd23,8'd72} : s = 95;
	{8'd23,8'd73} : s = 96;
	{8'd23,8'd74} : s = 97;
	{8'd23,8'd75} : s = 98;
	{8'd23,8'd76} : s = 99;
	{8'd23,8'd77} : s = 100;
	{8'd23,8'd78} : s = 101;
	{8'd23,8'd79} : s = 102;
	{8'd23,8'd80} : s = 103;
	{8'd23,8'd81} : s = 104;
	{8'd23,8'd82} : s = 105;
	{8'd23,8'd83} : s = 106;
	{8'd23,8'd84} : s = 107;
	{8'd23,8'd85} : s = 108;
	{8'd23,8'd86} : s = 109;
	{8'd23,8'd87} : s = 110;
	{8'd23,8'd88} : s = 111;
	{8'd23,8'd89} : s = 112;
	{8'd23,8'd90} : s = 113;
	{8'd23,8'd91} : s = 114;
	{8'd23,8'd92} : s = 115;
	{8'd23,8'd93} : s = 116;
	{8'd23,8'd94} : s = 117;
	{8'd23,8'd95} : s = 118;
	{8'd23,8'd96} : s = 119;
	{8'd23,8'd97} : s = 120;
	{8'd23,8'd98} : s = 121;
	{8'd23,8'd99} : s = 122;
	{8'd23,8'd100} : s = 123;
	{8'd23,8'd101} : s = 124;
	{8'd23,8'd102} : s = 125;
	{8'd23,8'd103} : s = 126;
	{8'd23,8'd104} : s = 127;
	{8'd23,8'd105} : s = 128;
	{8'd23,8'd106} : s = 129;
	{8'd23,8'd107} : s = 130;
	{8'd23,8'd108} : s = 131;
	{8'd23,8'd109} : s = 132;
	{8'd23,8'd110} : s = 133;
	{8'd23,8'd111} : s = 134;
	{8'd23,8'd112} : s = 135;
	{8'd23,8'd113} : s = 136;
	{8'd23,8'd114} : s = 137;
	{8'd23,8'd115} : s = 138;
	{8'd23,8'd116} : s = 139;
	{8'd23,8'd117} : s = 140;
	{8'd23,8'd118} : s = 141;
	{8'd23,8'd119} : s = 142;
	{8'd23,8'd120} : s = 143;
	{8'd23,8'd121} : s = 144;
	{8'd23,8'd122} : s = 145;
	{8'd23,8'd123} : s = 146;
	{8'd23,8'd124} : s = 147;
	{8'd23,8'd125} : s = 148;
	{8'd23,8'd126} : s = 149;
	{8'd23,8'd127} : s = 150;
	{8'd23,8'd128} : s = 151;
	{8'd23,8'd129} : s = 152;
	{8'd23,8'd130} : s = 153;
	{8'd23,8'd131} : s = 154;
	{8'd23,8'd132} : s = 155;
	{8'd23,8'd133} : s = 156;
	{8'd23,8'd134} : s = 157;
	{8'd23,8'd135} : s = 158;
	{8'd23,8'd136} : s = 159;
	{8'd23,8'd137} : s = 160;
	{8'd23,8'd138} : s = 161;
	{8'd23,8'd139} : s = 162;
	{8'd23,8'd140} : s = 163;
	{8'd23,8'd141} : s = 164;
	{8'd23,8'd142} : s = 165;
	{8'd23,8'd143} : s = 166;
	{8'd23,8'd144} : s = 167;
	{8'd23,8'd145} : s = 168;
	{8'd23,8'd146} : s = 169;
	{8'd23,8'd147} : s = 170;
	{8'd23,8'd148} : s = 171;
	{8'd23,8'd149} : s = 172;
	{8'd23,8'd150} : s = 173;
	{8'd23,8'd151} : s = 174;
	{8'd23,8'd152} : s = 175;
	{8'd23,8'd153} : s = 176;
	{8'd23,8'd154} : s = 177;
	{8'd23,8'd155} : s = 178;
	{8'd23,8'd156} : s = 179;
	{8'd23,8'd157} : s = 180;
	{8'd23,8'd158} : s = 181;
	{8'd23,8'd159} : s = 182;
	{8'd23,8'd160} : s = 183;
	{8'd23,8'd161} : s = 184;
	{8'd23,8'd162} : s = 185;
	{8'd23,8'd163} : s = 186;
	{8'd23,8'd164} : s = 187;
	{8'd23,8'd165} : s = 188;
	{8'd23,8'd166} : s = 189;
	{8'd23,8'd167} : s = 190;
	{8'd23,8'd168} : s = 191;
	{8'd23,8'd169} : s = 192;
	{8'd23,8'd170} : s = 193;
	{8'd23,8'd171} : s = 194;
	{8'd23,8'd172} : s = 195;
	{8'd23,8'd173} : s = 196;
	{8'd23,8'd174} : s = 197;
	{8'd23,8'd175} : s = 198;
	{8'd23,8'd176} : s = 199;
	{8'd23,8'd177} : s = 200;
	{8'd23,8'd178} : s = 201;
	{8'd23,8'd179} : s = 202;
	{8'd23,8'd180} : s = 203;
	{8'd23,8'd181} : s = 204;
	{8'd23,8'd182} : s = 205;
	{8'd23,8'd183} : s = 206;
	{8'd23,8'd184} : s = 207;
	{8'd23,8'd185} : s = 208;
	{8'd23,8'd186} : s = 209;
	{8'd23,8'd187} : s = 210;
	{8'd23,8'd188} : s = 211;
	{8'd23,8'd189} : s = 212;
	{8'd23,8'd190} : s = 213;
	{8'd23,8'd191} : s = 214;
	{8'd23,8'd192} : s = 215;
	{8'd23,8'd193} : s = 216;
	{8'd23,8'd194} : s = 217;
	{8'd23,8'd195} : s = 218;
	{8'd23,8'd196} : s = 219;
	{8'd23,8'd197} : s = 220;
	{8'd23,8'd198} : s = 221;
	{8'd23,8'd199} : s = 222;
	{8'd23,8'd200} : s = 223;
	{8'd23,8'd201} : s = 224;
	{8'd23,8'd202} : s = 225;
	{8'd23,8'd203} : s = 226;
	{8'd23,8'd204} : s = 227;
	{8'd23,8'd205} : s = 228;
	{8'd23,8'd206} : s = 229;
	{8'd23,8'd207} : s = 230;
	{8'd23,8'd208} : s = 231;
	{8'd23,8'd209} : s = 232;
	{8'd23,8'd210} : s = 233;
	{8'd23,8'd211} : s = 234;
	{8'd23,8'd212} : s = 235;
	{8'd23,8'd213} : s = 236;
	{8'd23,8'd214} : s = 237;
	{8'd23,8'd215} : s = 238;
	{8'd23,8'd216} : s = 239;
	{8'd23,8'd217} : s = 240;
	{8'd23,8'd218} : s = 241;
	{8'd23,8'd219} : s = 242;
	{8'd23,8'd220} : s = 243;
	{8'd23,8'd221} : s = 244;
	{8'd23,8'd222} : s = 245;
	{8'd23,8'd223} : s = 246;
	{8'd23,8'd224} : s = 247;
	{8'd23,8'd225} : s = 248;
	{8'd23,8'd226} : s = 249;
	{8'd23,8'd227} : s = 250;
	{8'd23,8'd228} : s = 251;
	{8'd23,8'd229} : s = 252;
	{8'd23,8'd230} : s = 253;
	{8'd23,8'd231} : s = 254;
	{8'd23,8'd232} : s = 255;
	{8'd23,8'd233} : s = 256;
	{8'd23,8'd234} : s = 257;
	{8'd23,8'd235} : s = 258;
	{8'd23,8'd236} : s = 259;
	{8'd23,8'd237} : s = 260;
	{8'd23,8'd238} : s = 261;
	{8'd23,8'd239} : s = 262;
	{8'd23,8'd240} : s = 263;
	{8'd23,8'd241} : s = 264;
	{8'd23,8'd242} : s = 265;
	{8'd23,8'd243} : s = 266;
	{8'd23,8'd244} : s = 267;
	{8'd23,8'd245} : s = 268;
	{8'd23,8'd246} : s = 269;
	{8'd23,8'd247} : s = 270;
	{8'd23,8'd248} : s = 271;
	{8'd23,8'd249} : s = 272;
	{8'd23,8'd250} : s = 273;
	{8'd23,8'd251} : s = 274;
	{8'd23,8'd252} : s = 275;
	{8'd23,8'd253} : s = 276;
	{8'd23,8'd254} : s = 277;
	{8'd23,8'd255} : s = 278;
	{8'd24,8'd0} : s = 24;
	{8'd24,8'd1} : s = 25;
	{8'd24,8'd2} : s = 26;
	{8'd24,8'd3} : s = 27;
	{8'd24,8'd4} : s = 28;
	{8'd24,8'd5} : s = 29;
	{8'd24,8'd6} : s = 30;
	{8'd24,8'd7} : s = 31;
	{8'd24,8'd8} : s = 32;
	{8'd24,8'd9} : s = 33;
	{8'd24,8'd10} : s = 34;
	{8'd24,8'd11} : s = 35;
	{8'd24,8'd12} : s = 36;
	{8'd24,8'd13} : s = 37;
	{8'd24,8'd14} : s = 38;
	{8'd24,8'd15} : s = 39;
	{8'd24,8'd16} : s = 40;
	{8'd24,8'd17} : s = 41;
	{8'd24,8'd18} : s = 42;
	{8'd24,8'd19} : s = 43;
	{8'd24,8'd20} : s = 44;
	{8'd24,8'd21} : s = 45;
	{8'd24,8'd22} : s = 46;
	{8'd24,8'd23} : s = 47;
	{8'd24,8'd24} : s = 48;
	{8'd24,8'd25} : s = 49;
	{8'd24,8'd26} : s = 50;
	{8'd24,8'd27} : s = 51;
	{8'd24,8'd28} : s = 52;
	{8'd24,8'd29} : s = 53;
	{8'd24,8'd30} : s = 54;
	{8'd24,8'd31} : s = 55;
	{8'd24,8'd32} : s = 56;
	{8'd24,8'd33} : s = 57;
	{8'd24,8'd34} : s = 58;
	{8'd24,8'd35} : s = 59;
	{8'd24,8'd36} : s = 60;
	{8'd24,8'd37} : s = 61;
	{8'd24,8'd38} : s = 62;
	{8'd24,8'd39} : s = 63;
	{8'd24,8'd40} : s = 64;
	{8'd24,8'd41} : s = 65;
	{8'd24,8'd42} : s = 66;
	{8'd24,8'd43} : s = 67;
	{8'd24,8'd44} : s = 68;
	{8'd24,8'd45} : s = 69;
	{8'd24,8'd46} : s = 70;
	{8'd24,8'd47} : s = 71;
	{8'd24,8'd48} : s = 72;
	{8'd24,8'd49} : s = 73;
	{8'd24,8'd50} : s = 74;
	{8'd24,8'd51} : s = 75;
	{8'd24,8'd52} : s = 76;
	{8'd24,8'd53} : s = 77;
	{8'd24,8'd54} : s = 78;
	{8'd24,8'd55} : s = 79;
	{8'd24,8'd56} : s = 80;
	{8'd24,8'd57} : s = 81;
	{8'd24,8'd58} : s = 82;
	{8'd24,8'd59} : s = 83;
	{8'd24,8'd60} : s = 84;
	{8'd24,8'd61} : s = 85;
	{8'd24,8'd62} : s = 86;
	{8'd24,8'd63} : s = 87;
	{8'd24,8'd64} : s = 88;
	{8'd24,8'd65} : s = 89;
	{8'd24,8'd66} : s = 90;
	{8'd24,8'd67} : s = 91;
	{8'd24,8'd68} : s = 92;
	{8'd24,8'd69} : s = 93;
	{8'd24,8'd70} : s = 94;
	{8'd24,8'd71} : s = 95;
	{8'd24,8'd72} : s = 96;
	{8'd24,8'd73} : s = 97;
	{8'd24,8'd74} : s = 98;
	{8'd24,8'd75} : s = 99;
	{8'd24,8'd76} : s = 100;
	{8'd24,8'd77} : s = 101;
	{8'd24,8'd78} : s = 102;
	{8'd24,8'd79} : s = 103;
	{8'd24,8'd80} : s = 104;
	{8'd24,8'd81} : s = 105;
	{8'd24,8'd82} : s = 106;
	{8'd24,8'd83} : s = 107;
	{8'd24,8'd84} : s = 108;
	{8'd24,8'd85} : s = 109;
	{8'd24,8'd86} : s = 110;
	{8'd24,8'd87} : s = 111;
	{8'd24,8'd88} : s = 112;
	{8'd24,8'd89} : s = 113;
	{8'd24,8'd90} : s = 114;
	{8'd24,8'd91} : s = 115;
	{8'd24,8'd92} : s = 116;
	{8'd24,8'd93} : s = 117;
	{8'd24,8'd94} : s = 118;
	{8'd24,8'd95} : s = 119;
	{8'd24,8'd96} : s = 120;
	{8'd24,8'd97} : s = 121;
	{8'd24,8'd98} : s = 122;
	{8'd24,8'd99} : s = 123;
	{8'd24,8'd100} : s = 124;
	{8'd24,8'd101} : s = 125;
	{8'd24,8'd102} : s = 126;
	{8'd24,8'd103} : s = 127;
	{8'd24,8'd104} : s = 128;
	{8'd24,8'd105} : s = 129;
	{8'd24,8'd106} : s = 130;
	{8'd24,8'd107} : s = 131;
	{8'd24,8'd108} : s = 132;
	{8'd24,8'd109} : s = 133;
	{8'd24,8'd110} : s = 134;
	{8'd24,8'd111} : s = 135;
	{8'd24,8'd112} : s = 136;
	{8'd24,8'd113} : s = 137;
	{8'd24,8'd114} : s = 138;
	{8'd24,8'd115} : s = 139;
	{8'd24,8'd116} : s = 140;
	{8'd24,8'd117} : s = 141;
	{8'd24,8'd118} : s = 142;
	{8'd24,8'd119} : s = 143;
	{8'd24,8'd120} : s = 144;
	{8'd24,8'd121} : s = 145;
	{8'd24,8'd122} : s = 146;
	{8'd24,8'd123} : s = 147;
	{8'd24,8'd124} : s = 148;
	{8'd24,8'd125} : s = 149;
	{8'd24,8'd126} : s = 150;
	{8'd24,8'd127} : s = 151;
	{8'd24,8'd128} : s = 152;
	{8'd24,8'd129} : s = 153;
	{8'd24,8'd130} : s = 154;
	{8'd24,8'd131} : s = 155;
	{8'd24,8'd132} : s = 156;
	{8'd24,8'd133} : s = 157;
	{8'd24,8'd134} : s = 158;
	{8'd24,8'd135} : s = 159;
	{8'd24,8'd136} : s = 160;
	{8'd24,8'd137} : s = 161;
	{8'd24,8'd138} : s = 162;
	{8'd24,8'd139} : s = 163;
	{8'd24,8'd140} : s = 164;
	{8'd24,8'd141} : s = 165;
	{8'd24,8'd142} : s = 166;
	{8'd24,8'd143} : s = 167;
	{8'd24,8'd144} : s = 168;
	{8'd24,8'd145} : s = 169;
	{8'd24,8'd146} : s = 170;
	{8'd24,8'd147} : s = 171;
	{8'd24,8'd148} : s = 172;
	{8'd24,8'd149} : s = 173;
	{8'd24,8'd150} : s = 174;
	{8'd24,8'd151} : s = 175;
	{8'd24,8'd152} : s = 176;
	{8'd24,8'd153} : s = 177;
	{8'd24,8'd154} : s = 178;
	{8'd24,8'd155} : s = 179;
	{8'd24,8'd156} : s = 180;
	{8'd24,8'd157} : s = 181;
	{8'd24,8'd158} : s = 182;
	{8'd24,8'd159} : s = 183;
	{8'd24,8'd160} : s = 184;
	{8'd24,8'd161} : s = 185;
	{8'd24,8'd162} : s = 186;
	{8'd24,8'd163} : s = 187;
	{8'd24,8'd164} : s = 188;
	{8'd24,8'd165} : s = 189;
	{8'd24,8'd166} : s = 190;
	{8'd24,8'd167} : s = 191;
	{8'd24,8'd168} : s = 192;
	{8'd24,8'd169} : s = 193;
	{8'd24,8'd170} : s = 194;
	{8'd24,8'd171} : s = 195;
	{8'd24,8'd172} : s = 196;
	{8'd24,8'd173} : s = 197;
	{8'd24,8'd174} : s = 198;
	{8'd24,8'd175} : s = 199;
	{8'd24,8'd176} : s = 200;
	{8'd24,8'd177} : s = 201;
	{8'd24,8'd178} : s = 202;
	{8'd24,8'd179} : s = 203;
	{8'd24,8'd180} : s = 204;
	{8'd24,8'd181} : s = 205;
	{8'd24,8'd182} : s = 206;
	{8'd24,8'd183} : s = 207;
	{8'd24,8'd184} : s = 208;
	{8'd24,8'd185} : s = 209;
	{8'd24,8'd186} : s = 210;
	{8'd24,8'd187} : s = 211;
	{8'd24,8'd188} : s = 212;
	{8'd24,8'd189} : s = 213;
	{8'd24,8'd190} : s = 214;
	{8'd24,8'd191} : s = 215;
	{8'd24,8'd192} : s = 216;
	{8'd24,8'd193} : s = 217;
	{8'd24,8'd194} : s = 218;
	{8'd24,8'd195} : s = 219;
	{8'd24,8'd196} : s = 220;
	{8'd24,8'd197} : s = 221;
	{8'd24,8'd198} : s = 222;
	{8'd24,8'd199} : s = 223;
	{8'd24,8'd200} : s = 224;
	{8'd24,8'd201} : s = 225;
	{8'd24,8'd202} : s = 226;
	{8'd24,8'd203} : s = 227;
	{8'd24,8'd204} : s = 228;
	{8'd24,8'd205} : s = 229;
	{8'd24,8'd206} : s = 230;
	{8'd24,8'd207} : s = 231;
	{8'd24,8'd208} : s = 232;
	{8'd24,8'd209} : s = 233;
	{8'd24,8'd210} : s = 234;
	{8'd24,8'd211} : s = 235;
	{8'd24,8'd212} : s = 236;
	{8'd24,8'd213} : s = 237;
	{8'd24,8'd214} : s = 238;
	{8'd24,8'd215} : s = 239;
	{8'd24,8'd216} : s = 240;
	{8'd24,8'd217} : s = 241;
	{8'd24,8'd218} : s = 242;
	{8'd24,8'd219} : s = 243;
	{8'd24,8'd220} : s = 244;
	{8'd24,8'd221} : s = 245;
	{8'd24,8'd222} : s = 246;
	{8'd24,8'd223} : s = 247;
	{8'd24,8'd224} : s = 248;
	{8'd24,8'd225} : s = 249;
	{8'd24,8'd226} : s = 250;
	{8'd24,8'd227} : s = 251;
	{8'd24,8'd228} : s = 252;
	{8'd24,8'd229} : s = 253;
	{8'd24,8'd230} : s = 254;
	{8'd24,8'd231} : s = 255;
	{8'd24,8'd232} : s = 256;
	{8'd24,8'd233} : s = 257;
	{8'd24,8'd234} : s = 258;
	{8'd24,8'd235} : s = 259;
	{8'd24,8'd236} : s = 260;
	{8'd24,8'd237} : s = 261;
	{8'd24,8'd238} : s = 262;
	{8'd24,8'd239} : s = 263;
	{8'd24,8'd240} : s = 264;
	{8'd24,8'd241} : s = 265;
	{8'd24,8'd242} : s = 266;
	{8'd24,8'd243} : s = 267;
	{8'd24,8'd244} : s = 268;
	{8'd24,8'd245} : s = 269;
	{8'd24,8'd246} : s = 270;
	{8'd24,8'd247} : s = 271;
	{8'd24,8'd248} : s = 272;
	{8'd24,8'd249} : s = 273;
	{8'd24,8'd250} : s = 274;
	{8'd24,8'd251} : s = 275;
	{8'd24,8'd252} : s = 276;
	{8'd24,8'd253} : s = 277;
	{8'd24,8'd254} : s = 278;
	{8'd24,8'd255} : s = 279;
	{8'd25,8'd0} : s = 25;
	{8'd25,8'd1} : s = 26;
	{8'd25,8'd2} : s = 27;
	{8'd25,8'd3} : s = 28;
	{8'd25,8'd4} : s = 29;
	{8'd25,8'd5} : s = 30;
	{8'd25,8'd6} : s = 31;
	{8'd25,8'd7} : s = 32;
	{8'd25,8'd8} : s = 33;
	{8'd25,8'd9} : s = 34;
	{8'd25,8'd10} : s = 35;
	{8'd25,8'd11} : s = 36;
	{8'd25,8'd12} : s = 37;
	{8'd25,8'd13} : s = 38;
	{8'd25,8'd14} : s = 39;
	{8'd25,8'd15} : s = 40;
	{8'd25,8'd16} : s = 41;
	{8'd25,8'd17} : s = 42;
	{8'd25,8'd18} : s = 43;
	{8'd25,8'd19} : s = 44;
	{8'd25,8'd20} : s = 45;
	{8'd25,8'd21} : s = 46;
	{8'd25,8'd22} : s = 47;
	{8'd25,8'd23} : s = 48;
	{8'd25,8'd24} : s = 49;
	{8'd25,8'd25} : s = 50;
	{8'd25,8'd26} : s = 51;
	{8'd25,8'd27} : s = 52;
	{8'd25,8'd28} : s = 53;
	{8'd25,8'd29} : s = 54;
	{8'd25,8'd30} : s = 55;
	{8'd25,8'd31} : s = 56;
	{8'd25,8'd32} : s = 57;
	{8'd25,8'd33} : s = 58;
	{8'd25,8'd34} : s = 59;
	{8'd25,8'd35} : s = 60;
	{8'd25,8'd36} : s = 61;
	{8'd25,8'd37} : s = 62;
	{8'd25,8'd38} : s = 63;
	{8'd25,8'd39} : s = 64;
	{8'd25,8'd40} : s = 65;
	{8'd25,8'd41} : s = 66;
	{8'd25,8'd42} : s = 67;
	{8'd25,8'd43} : s = 68;
	{8'd25,8'd44} : s = 69;
	{8'd25,8'd45} : s = 70;
	{8'd25,8'd46} : s = 71;
	{8'd25,8'd47} : s = 72;
	{8'd25,8'd48} : s = 73;
	{8'd25,8'd49} : s = 74;
	{8'd25,8'd50} : s = 75;
	{8'd25,8'd51} : s = 76;
	{8'd25,8'd52} : s = 77;
	{8'd25,8'd53} : s = 78;
	{8'd25,8'd54} : s = 79;
	{8'd25,8'd55} : s = 80;
	{8'd25,8'd56} : s = 81;
	{8'd25,8'd57} : s = 82;
	{8'd25,8'd58} : s = 83;
	{8'd25,8'd59} : s = 84;
	{8'd25,8'd60} : s = 85;
	{8'd25,8'd61} : s = 86;
	{8'd25,8'd62} : s = 87;
	{8'd25,8'd63} : s = 88;
	{8'd25,8'd64} : s = 89;
	{8'd25,8'd65} : s = 90;
	{8'd25,8'd66} : s = 91;
	{8'd25,8'd67} : s = 92;
	{8'd25,8'd68} : s = 93;
	{8'd25,8'd69} : s = 94;
	{8'd25,8'd70} : s = 95;
	{8'd25,8'd71} : s = 96;
	{8'd25,8'd72} : s = 97;
	{8'd25,8'd73} : s = 98;
	{8'd25,8'd74} : s = 99;
	{8'd25,8'd75} : s = 100;
	{8'd25,8'd76} : s = 101;
	{8'd25,8'd77} : s = 102;
	{8'd25,8'd78} : s = 103;
	{8'd25,8'd79} : s = 104;
	{8'd25,8'd80} : s = 105;
	{8'd25,8'd81} : s = 106;
	{8'd25,8'd82} : s = 107;
	{8'd25,8'd83} : s = 108;
	{8'd25,8'd84} : s = 109;
	{8'd25,8'd85} : s = 110;
	{8'd25,8'd86} : s = 111;
	{8'd25,8'd87} : s = 112;
	{8'd25,8'd88} : s = 113;
	{8'd25,8'd89} : s = 114;
	{8'd25,8'd90} : s = 115;
	{8'd25,8'd91} : s = 116;
	{8'd25,8'd92} : s = 117;
	{8'd25,8'd93} : s = 118;
	{8'd25,8'd94} : s = 119;
	{8'd25,8'd95} : s = 120;
	{8'd25,8'd96} : s = 121;
	{8'd25,8'd97} : s = 122;
	{8'd25,8'd98} : s = 123;
	{8'd25,8'd99} : s = 124;
	{8'd25,8'd100} : s = 125;
	{8'd25,8'd101} : s = 126;
	{8'd25,8'd102} : s = 127;
	{8'd25,8'd103} : s = 128;
	{8'd25,8'd104} : s = 129;
	{8'd25,8'd105} : s = 130;
	{8'd25,8'd106} : s = 131;
	{8'd25,8'd107} : s = 132;
	{8'd25,8'd108} : s = 133;
	{8'd25,8'd109} : s = 134;
	{8'd25,8'd110} : s = 135;
	{8'd25,8'd111} : s = 136;
	{8'd25,8'd112} : s = 137;
	{8'd25,8'd113} : s = 138;
	{8'd25,8'd114} : s = 139;
	{8'd25,8'd115} : s = 140;
	{8'd25,8'd116} : s = 141;
	{8'd25,8'd117} : s = 142;
	{8'd25,8'd118} : s = 143;
	{8'd25,8'd119} : s = 144;
	{8'd25,8'd120} : s = 145;
	{8'd25,8'd121} : s = 146;
	{8'd25,8'd122} : s = 147;
	{8'd25,8'd123} : s = 148;
	{8'd25,8'd124} : s = 149;
	{8'd25,8'd125} : s = 150;
	{8'd25,8'd126} : s = 151;
	{8'd25,8'd127} : s = 152;
	{8'd25,8'd128} : s = 153;
	{8'd25,8'd129} : s = 154;
	{8'd25,8'd130} : s = 155;
	{8'd25,8'd131} : s = 156;
	{8'd25,8'd132} : s = 157;
	{8'd25,8'd133} : s = 158;
	{8'd25,8'd134} : s = 159;
	{8'd25,8'd135} : s = 160;
	{8'd25,8'd136} : s = 161;
	{8'd25,8'd137} : s = 162;
	{8'd25,8'd138} : s = 163;
	{8'd25,8'd139} : s = 164;
	{8'd25,8'd140} : s = 165;
	{8'd25,8'd141} : s = 166;
	{8'd25,8'd142} : s = 167;
	{8'd25,8'd143} : s = 168;
	{8'd25,8'd144} : s = 169;
	{8'd25,8'd145} : s = 170;
	{8'd25,8'd146} : s = 171;
	{8'd25,8'd147} : s = 172;
	{8'd25,8'd148} : s = 173;
	{8'd25,8'd149} : s = 174;
	{8'd25,8'd150} : s = 175;
	{8'd25,8'd151} : s = 176;
	{8'd25,8'd152} : s = 177;
	{8'd25,8'd153} : s = 178;
	{8'd25,8'd154} : s = 179;
	{8'd25,8'd155} : s = 180;
	{8'd25,8'd156} : s = 181;
	{8'd25,8'd157} : s = 182;
	{8'd25,8'd158} : s = 183;
	{8'd25,8'd159} : s = 184;
	{8'd25,8'd160} : s = 185;
	{8'd25,8'd161} : s = 186;
	{8'd25,8'd162} : s = 187;
	{8'd25,8'd163} : s = 188;
	{8'd25,8'd164} : s = 189;
	{8'd25,8'd165} : s = 190;
	{8'd25,8'd166} : s = 191;
	{8'd25,8'd167} : s = 192;
	{8'd25,8'd168} : s = 193;
	{8'd25,8'd169} : s = 194;
	{8'd25,8'd170} : s = 195;
	{8'd25,8'd171} : s = 196;
	{8'd25,8'd172} : s = 197;
	{8'd25,8'd173} : s = 198;
	{8'd25,8'd174} : s = 199;
	{8'd25,8'd175} : s = 200;
	{8'd25,8'd176} : s = 201;
	{8'd25,8'd177} : s = 202;
	{8'd25,8'd178} : s = 203;
	{8'd25,8'd179} : s = 204;
	{8'd25,8'd180} : s = 205;
	{8'd25,8'd181} : s = 206;
	{8'd25,8'd182} : s = 207;
	{8'd25,8'd183} : s = 208;
	{8'd25,8'd184} : s = 209;
	{8'd25,8'd185} : s = 210;
	{8'd25,8'd186} : s = 211;
	{8'd25,8'd187} : s = 212;
	{8'd25,8'd188} : s = 213;
	{8'd25,8'd189} : s = 214;
	{8'd25,8'd190} : s = 215;
	{8'd25,8'd191} : s = 216;
	{8'd25,8'd192} : s = 217;
	{8'd25,8'd193} : s = 218;
	{8'd25,8'd194} : s = 219;
	{8'd25,8'd195} : s = 220;
	{8'd25,8'd196} : s = 221;
	{8'd25,8'd197} : s = 222;
	{8'd25,8'd198} : s = 223;
	{8'd25,8'd199} : s = 224;
	{8'd25,8'd200} : s = 225;
	{8'd25,8'd201} : s = 226;
	{8'd25,8'd202} : s = 227;
	{8'd25,8'd203} : s = 228;
	{8'd25,8'd204} : s = 229;
	{8'd25,8'd205} : s = 230;
	{8'd25,8'd206} : s = 231;
	{8'd25,8'd207} : s = 232;
	{8'd25,8'd208} : s = 233;
	{8'd25,8'd209} : s = 234;
	{8'd25,8'd210} : s = 235;
	{8'd25,8'd211} : s = 236;
	{8'd25,8'd212} : s = 237;
	{8'd25,8'd213} : s = 238;
	{8'd25,8'd214} : s = 239;
	{8'd25,8'd215} : s = 240;
	{8'd25,8'd216} : s = 241;
	{8'd25,8'd217} : s = 242;
	{8'd25,8'd218} : s = 243;
	{8'd25,8'd219} : s = 244;
	{8'd25,8'd220} : s = 245;
	{8'd25,8'd221} : s = 246;
	{8'd25,8'd222} : s = 247;
	{8'd25,8'd223} : s = 248;
	{8'd25,8'd224} : s = 249;
	{8'd25,8'd225} : s = 250;
	{8'd25,8'd226} : s = 251;
	{8'd25,8'd227} : s = 252;
	{8'd25,8'd228} : s = 253;
	{8'd25,8'd229} : s = 254;
	{8'd25,8'd230} : s = 255;
	{8'd25,8'd231} : s = 256;
	{8'd25,8'd232} : s = 257;
	{8'd25,8'd233} : s = 258;
	{8'd25,8'd234} : s = 259;
	{8'd25,8'd235} : s = 260;
	{8'd25,8'd236} : s = 261;
	{8'd25,8'd237} : s = 262;
	{8'd25,8'd238} : s = 263;
	{8'd25,8'd239} : s = 264;
	{8'd25,8'd240} : s = 265;
	{8'd25,8'd241} : s = 266;
	{8'd25,8'd242} : s = 267;
	{8'd25,8'd243} : s = 268;
	{8'd25,8'd244} : s = 269;
	{8'd25,8'd245} : s = 270;
	{8'd25,8'd246} : s = 271;
	{8'd25,8'd247} : s = 272;
	{8'd25,8'd248} : s = 273;
	{8'd25,8'd249} : s = 274;
	{8'd25,8'd250} : s = 275;
	{8'd25,8'd251} : s = 276;
	{8'd25,8'd252} : s = 277;
	{8'd25,8'd253} : s = 278;
	{8'd25,8'd254} : s = 279;
	{8'd25,8'd255} : s = 280;
	{8'd26,8'd0} : s = 26;
	{8'd26,8'd1} : s = 27;
	{8'd26,8'd2} : s = 28;
	{8'd26,8'd3} : s = 29;
	{8'd26,8'd4} : s = 30;
	{8'd26,8'd5} : s = 31;
	{8'd26,8'd6} : s = 32;
	{8'd26,8'd7} : s = 33;
	{8'd26,8'd8} : s = 34;
	{8'd26,8'd9} : s = 35;
	{8'd26,8'd10} : s = 36;
	{8'd26,8'd11} : s = 37;
	{8'd26,8'd12} : s = 38;
	{8'd26,8'd13} : s = 39;
	{8'd26,8'd14} : s = 40;
	{8'd26,8'd15} : s = 41;
	{8'd26,8'd16} : s = 42;
	{8'd26,8'd17} : s = 43;
	{8'd26,8'd18} : s = 44;
	{8'd26,8'd19} : s = 45;
	{8'd26,8'd20} : s = 46;
	{8'd26,8'd21} : s = 47;
	{8'd26,8'd22} : s = 48;
	{8'd26,8'd23} : s = 49;
	{8'd26,8'd24} : s = 50;
	{8'd26,8'd25} : s = 51;
	{8'd26,8'd26} : s = 52;
	{8'd26,8'd27} : s = 53;
	{8'd26,8'd28} : s = 54;
	{8'd26,8'd29} : s = 55;
	{8'd26,8'd30} : s = 56;
	{8'd26,8'd31} : s = 57;
	{8'd26,8'd32} : s = 58;
	{8'd26,8'd33} : s = 59;
	{8'd26,8'd34} : s = 60;
	{8'd26,8'd35} : s = 61;
	{8'd26,8'd36} : s = 62;
	{8'd26,8'd37} : s = 63;
	{8'd26,8'd38} : s = 64;
	{8'd26,8'd39} : s = 65;
	{8'd26,8'd40} : s = 66;
	{8'd26,8'd41} : s = 67;
	{8'd26,8'd42} : s = 68;
	{8'd26,8'd43} : s = 69;
	{8'd26,8'd44} : s = 70;
	{8'd26,8'd45} : s = 71;
	{8'd26,8'd46} : s = 72;
	{8'd26,8'd47} : s = 73;
	{8'd26,8'd48} : s = 74;
	{8'd26,8'd49} : s = 75;
	{8'd26,8'd50} : s = 76;
	{8'd26,8'd51} : s = 77;
	{8'd26,8'd52} : s = 78;
	{8'd26,8'd53} : s = 79;
	{8'd26,8'd54} : s = 80;
	{8'd26,8'd55} : s = 81;
	{8'd26,8'd56} : s = 82;
	{8'd26,8'd57} : s = 83;
	{8'd26,8'd58} : s = 84;
	{8'd26,8'd59} : s = 85;
	{8'd26,8'd60} : s = 86;
	{8'd26,8'd61} : s = 87;
	{8'd26,8'd62} : s = 88;
	{8'd26,8'd63} : s = 89;
	{8'd26,8'd64} : s = 90;
	{8'd26,8'd65} : s = 91;
	{8'd26,8'd66} : s = 92;
	{8'd26,8'd67} : s = 93;
	{8'd26,8'd68} : s = 94;
	{8'd26,8'd69} : s = 95;
	{8'd26,8'd70} : s = 96;
	{8'd26,8'd71} : s = 97;
	{8'd26,8'd72} : s = 98;
	{8'd26,8'd73} : s = 99;
	{8'd26,8'd74} : s = 100;
	{8'd26,8'd75} : s = 101;
	{8'd26,8'd76} : s = 102;
	{8'd26,8'd77} : s = 103;
	{8'd26,8'd78} : s = 104;
	{8'd26,8'd79} : s = 105;
	{8'd26,8'd80} : s = 106;
	{8'd26,8'd81} : s = 107;
	{8'd26,8'd82} : s = 108;
	{8'd26,8'd83} : s = 109;
	{8'd26,8'd84} : s = 110;
	{8'd26,8'd85} : s = 111;
	{8'd26,8'd86} : s = 112;
	{8'd26,8'd87} : s = 113;
	{8'd26,8'd88} : s = 114;
	{8'd26,8'd89} : s = 115;
	{8'd26,8'd90} : s = 116;
	{8'd26,8'd91} : s = 117;
	{8'd26,8'd92} : s = 118;
	{8'd26,8'd93} : s = 119;
	{8'd26,8'd94} : s = 120;
	{8'd26,8'd95} : s = 121;
	{8'd26,8'd96} : s = 122;
	{8'd26,8'd97} : s = 123;
	{8'd26,8'd98} : s = 124;
	{8'd26,8'd99} : s = 125;
	{8'd26,8'd100} : s = 126;
	{8'd26,8'd101} : s = 127;
	{8'd26,8'd102} : s = 128;
	{8'd26,8'd103} : s = 129;
	{8'd26,8'd104} : s = 130;
	{8'd26,8'd105} : s = 131;
	{8'd26,8'd106} : s = 132;
	{8'd26,8'd107} : s = 133;
	{8'd26,8'd108} : s = 134;
	{8'd26,8'd109} : s = 135;
	{8'd26,8'd110} : s = 136;
	{8'd26,8'd111} : s = 137;
	{8'd26,8'd112} : s = 138;
	{8'd26,8'd113} : s = 139;
	{8'd26,8'd114} : s = 140;
	{8'd26,8'd115} : s = 141;
	{8'd26,8'd116} : s = 142;
	{8'd26,8'd117} : s = 143;
	{8'd26,8'd118} : s = 144;
	{8'd26,8'd119} : s = 145;
	{8'd26,8'd120} : s = 146;
	{8'd26,8'd121} : s = 147;
	{8'd26,8'd122} : s = 148;
	{8'd26,8'd123} : s = 149;
	{8'd26,8'd124} : s = 150;
	{8'd26,8'd125} : s = 151;
	{8'd26,8'd126} : s = 152;
	{8'd26,8'd127} : s = 153;
	{8'd26,8'd128} : s = 154;
	{8'd26,8'd129} : s = 155;
	{8'd26,8'd130} : s = 156;
	{8'd26,8'd131} : s = 157;
	{8'd26,8'd132} : s = 158;
	{8'd26,8'd133} : s = 159;
	{8'd26,8'd134} : s = 160;
	{8'd26,8'd135} : s = 161;
	{8'd26,8'd136} : s = 162;
	{8'd26,8'd137} : s = 163;
	{8'd26,8'd138} : s = 164;
	{8'd26,8'd139} : s = 165;
	{8'd26,8'd140} : s = 166;
	{8'd26,8'd141} : s = 167;
	{8'd26,8'd142} : s = 168;
	{8'd26,8'd143} : s = 169;
	{8'd26,8'd144} : s = 170;
	{8'd26,8'd145} : s = 171;
	{8'd26,8'd146} : s = 172;
	{8'd26,8'd147} : s = 173;
	{8'd26,8'd148} : s = 174;
	{8'd26,8'd149} : s = 175;
	{8'd26,8'd150} : s = 176;
	{8'd26,8'd151} : s = 177;
	{8'd26,8'd152} : s = 178;
	{8'd26,8'd153} : s = 179;
	{8'd26,8'd154} : s = 180;
	{8'd26,8'd155} : s = 181;
	{8'd26,8'd156} : s = 182;
	{8'd26,8'd157} : s = 183;
	{8'd26,8'd158} : s = 184;
	{8'd26,8'd159} : s = 185;
	{8'd26,8'd160} : s = 186;
	{8'd26,8'd161} : s = 187;
	{8'd26,8'd162} : s = 188;
	{8'd26,8'd163} : s = 189;
	{8'd26,8'd164} : s = 190;
	{8'd26,8'd165} : s = 191;
	{8'd26,8'd166} : s = 192;
	{8'd26,8'd167} : s = 193;
	{8'd26,8'd168} : s = 194;
	{8'd26,8'd169} : s = 195;
	{8'd26,8'd170} : s = 196;
	{8'd26,8'd171} : s = 197;
	{8'd26,8'd172} : s = 198;
	{8'd26,8'd173} : s = 199;
	{8'd26,8'd174} : s = 200;
	{8'd26,8'd175} : s = 201;
	{8'd26,8'd176} : s = 202;
	{8'd26,8'd177} : s = 203;
	{8'd26,8'd178} : s = 204;
	{8'd26,8'd179} : s = 205;
	{8'd26,8'd180} : s = 206;
	{8'd26,8'd181} : s = 207;
	{8'd26,8'd182} : s = 208;
	{8'd26,8'd183} : s = 209;
	{8'd26,8'd184} : s = 210;
	{8'd26,8'd185} : s = 211;
	{8'd26,8'd186} : s = 212;
	{8'd26,8'd187} : s = 213;
	{8'd26,8'd188} : s = 214;
	{8'd26,8'd189} : s = 215;
	{8'd26,8'd190} : s = 216;
	{8'd26,8'd191} : s = 217;
	{8'd26,8'd192} : s = 218;
	{8'd26,8'd193} : s = 219;
	{8'd26,8'd194} : s = 220;
	{8'd26,8'd195} : s = 221;
	{8'd26,8'd196} : s = 222;
	{8'd26,8'd197} : s = 223;
	{8'd26,8'd198} : s = 224;
	{8'd26,8'd199} : s = 225;
	{8'd26,8'd200} : s = 226;
	{8'd26,8'd201} : s = 227;
	{8'd26,8'd202} : s = 228;
	{8'd26,8'd203} : s = 229;
	{8'd26,8'd204} : s = 230;
	{8'd26,8'd205} : s = 231;
	{8'd26,8'd206} : s = 232;
	{8'd26,8'd207} : s = 233;
	{8'd26,8'd208} : s = 234;
	{8'd26,8'd209} : s = 235;
	{8'd26,8'd210} : s = 236;
	{8'd26,8'd211} : s = 237;
	{8'd26,8'd212} : s = 238;
	{8'd26,8'd213} : s = 239;
	{8'd26,8'd214} : s = 240;
	{8'd26,8'd215} : s = 241;
	{8'd26,8'd216} : s = 242;
	{8'd26,8'd217} : s = 243;
	{8'd26,8'd218} : s = 244;
	{8'd26,8'd219} : s = 245;
	{8'd26,8'd220} : s = 246;
	{8'd26,8'd221} : s = 247;
	{8'd26,8'd222} : s = 248;
	{8'd26,8'd223} : s = 249;
	{8'd26,8'd224} : s = 250;
	{8'd26,8'd225} : s = 251;
	{8'd26,8'd226} : s = 252;
	{8'd26,8'd227} : s = 253;
	{8'd26,8'd228} : s = 254;
	{8'd26,8'd229} : s = 255;
	{8'd26,8'd230} : s = 256;
	{8'd26,8'd231} : s = 257;
	{8'd26,8'd232} : s = 258;
	{8'd26,8'd233} : s = 259;
	{8'd26,8'd234} : s = 260;
	{8'd26,8'd235} : s = 261;
	{8'd26,8'd236} : s = 262;
	{8'd26,8'd237} : s = 263;
	{8'd26,8'd238} : s = 264;
	{8'd26,8'd239} : s = 265;
	{8'd26,8'd240} : s = 266;
	{8'd26,8'd241} : s = 267;
	{8'd26,8'd242} : s = 268;
	{8'd26,8'd243} : s = 269;
	{8'd26,8'd244} : s = 270;
	{8'd26,8'd245} : s = 271;
	{8'd26,8'd246} : s = 272;
	{8'd26,8'd247} : s = 273;
	{8'd26,8'd248} : s = 274;
	{8'd26,8'd249} : s = 275;
	{8'd26,8'd250} : s = 276;
	{8'd26,8'd251} : s = 277;
	{8'd26,8'd252} : s = 278;
	{8'd26,8'd253} : s = 279;
	{8'd26,8'd254} : s = 280;
	{8'd26,8'd255} : s = 281;
	{8'd27,8'd0} : s = 27;
	{8'd27,8'd1} : s = 28;
	{8'd27,8'd2} : s = 29;
	{8'd27,8'd3} : s = 30;
	{8'd27,8'd4} : s = 31;
	{8'd27,8'd5} : s = 32;
	{8'd27,8'd6} : s = 33;
	{8'd27,8'd7} : s = 34;
	{8'd27,8'd8} : s = 35;
	{8'd27,8'd9} : s = 36;
	{8'd27,8'd10} : s = 37;
	{8'd27,8'd11} : s = 38;
	{8'd27,8'd12} : s = 39;
	{8'd27,8'd13} : s = 40;
	{8'd27,8'd14} : s = 41;
	{8'd27,8'd15} : s = 42;
	{8'd27,8'd16} : s = 43;
	{8'd27,8'd17} : s = 44;
	{8'd27,8'd18} : s = 45;
	{8'd27,8'd19} : s = 46;
	{8'd27,8'd20} : s = 47;
	{8'd27,8'd21} : s = 48;
	{8'd27,8'd22} : s = 49;
	{8'd27,8'd23} : s = 50;
	{8'd27,8'd24} : s = 51;
	{8'd27,8'd25} : s = 52;
	{8'd27,8'd26} : s = 53;
	{8'd27,8'd27} : s = 54;
	{8'd27,8'd28} : s = 55;
	{8'd27,8'd29} : s = 56;
	{8'd27,8'd30} : s = 57;
	{8'd27,8'd31} : s = 58;
	{8'd27,8'd32} : s = 59;
	{8'd27,8'd33} : s = 60;
	{8'd27,8'd34} : s = 61;
	{8'd27,8'd35} : s = 62;
	{8'd27,8'd36} : s = 63;
	{8'd27,8'd37} : s = 64;
	{8'd27,8'd38} : s = 65;
	{8'd27,8'd39} : s = 66;
	{8'd27,8'd40} : s = 67;
	{8'd27,8'd41} : s = 68;
	{8'd27,8'd42} : s = 69;
	{8'd27,8'd43} : s = 70;
	{8'd27,8'd44} : s = 71;
	{8'd27,8'd45} : s = 72;
	{8'd27,8'd46} : s = 73;
	{8'd27,8'd47} : s = 74;
	{8'd27,8'd48} : s = 75;
	{8'd27,8'd49} : s = 76;
	{8'd27,8'd50} : s = 77;
	{8'd27,8'd51} : s = 78;
	{8'd27,8'd52} : s = 79;
	{8'd27,8'd53} : s = 80;
	{8'd27,8'd54} : s = 81;
	{8'd27,8'd55} : s = 82;
	{8'd27,8'd56} : s = 83;
	{8'd27,8'd57} : s = 84;
	{8'd27,8'd58} : s = 85;
	{8'd27,8'd59} : s = 86;
	{8'd27,8'd60} : s = 87;
	{8'd27,8'd61} : s = 88;
	{8'd27,8'd62} : s = 89;
	{8'd27,8'd63} : s = 90;
	{8'd27,8'd64} : s = 91;
	{8'd27,8'd65} : s = 92;
	{8'd27,8'd66} : s = 93;
	{8'd27,8'd67} : s = 94;
	{8'd27,8'd68} : s = 95;
	{8'd27,8'd69} : s = 96;
	{8'd27,8'd70} : s = 97;
	{8'd27,8'd71} : s = 98;
	{8'd27,8'd72} : s = 99;
	{8'd27,8'd73} : s = 100;
	{8'd27,8'd74} : s = 101;
	{8'd27,8'd75} : s = 102;
	{8'd27,8'd76} : s = 103;
	{8'd27,8'd77} : s = 104;
	{8'd27,8'd78} : s = 105;
	{8'd27,8'd79} : s = 106;
	{8'd27,8'd80} : s = 107;
	{8'd27,8'd81} : s = 108;
	{8'd27,8'd82} : s = 109;
	{8'd27,8'd83} : s = 110;
	{8'd27,8'd84} : s = 111;
	{8'd27,8'd85} : s = 112;
	{8'd27,8'd86} : s = 113;
	{8'd27,8'd87} : s = 114;
	{8'd27,8'd88} : s = 115;
	{8'd27,8'd89} : s = 116;
	{8'd27,8'd90} : s = 117;
	{8'd27,8'd91} : s = 118;
	{8'd27,8'd92} : s = 119;
	{8'd27,8'd93} : s = 120;
	{8'd27,8'd94} : s = 121;
	{8'd27,8'd95} : s = 122;
	{8'd27,8'd96} : s = 123;
	{8'd27,8'd97} : s = 124;
	{8'd27,8'd98} : s = 125;
	{8'd27,8'd99} : s = 126;
	{8'd27,8'd100} : s = 127;
	{8'd27,8'd101} : s = 128;
	{8'd27,8'd102} : s = 129;
	{8'd27,8'd103} : s = 130;
	{8'd27,8'd104} : s = 131;
	{8'd27,8'd105} : s = 132;
	{8'd27,8'd106} : s = 133;
	{8'd27,8'd107} : s = 134;
	{8'd27,8'd108} : s = 135;
	{8'd27,8'd109} : s = 136;
	{8'd27,8'd110} : s = 137;
	{8'd27,8'd111} : s = 138;
	{8'd27,8'd112} : s = 139;
	{8'd27,8'd113} : s = 140;
	{8'd27,8'd114} : s = 141;
	{8'd27,8'd115} : s = 142;
	{8'd27,8'd116} : s = 143;
	{8'd27,8'd117} : s = 144;
	{8'd27,8'd118} : s = 145;
	{8'd27,8'd119} : s = 146;
	{8'd27,8'd120} : s = 147;
	{8'd27,8'd121} : s = 148;
	{8'd27,8'd122} : s = 149;
	{8'd27,8'd123} : s = 150;
	{8'd27,8'd124} : s = 151;
	{8'd27,8'd125} : s = 152;
	{8'd27,8'd126} : s = 153;
	{8'd27,8'd127} : s = 154;
	{8'd27,8'd128} : s = 155;
	{8'd27,8'd129} : s = 156;
	{8'd27,8'd130} : s = 157;
	{8'd27,8'd131} : s = 158;
	{8'd27,8'd132} : s = 159;
	{8'd27,8'd133} : s = 160;
	{8'd27,8'd134} : s = 161;
	{8'd27,8'd135} : s = 162;
	{8'd27,8'd136} : s = 163;
	{8'd27,8'd137} : s = 164;
	{8'd27,8'd138} : s = 165;
	{8'd27,8'd139} : s = 166;
	{8'd27,8'd140} : s = 167;
	{8'd27,8'd141} : s = 168;
	{8'd27,8'd142} : s = 169;
	{8'd27,8'd143} : s = 170;
	{8'd27,8'd144} : s = 171;
	{8'd27,8'd145} : s = 172;
	{8'd27,8'd146} : s = 173;
	{8'd27,8'd147} : s = 174;
	{8'd27,8'd148} : s = 175;
	{8'd27,8'd149} : s = 176;
	{8'd27,8'd150} : s = 177;
	{8'd27,8'd151} : s = 178;
	{8'd27,8'd152} : s = 179;
	{8'd27,8'd153} : s = 180;
	{8'd27,8'd154} : s = 181;
	{8'd27,8'd155} : s = 182;
	{8'd27,8'd156} : s = 183;
	{8'd27,8'd157} : s = 184;
	{8'd27,8'd158} : s = 185;
	{8'd27,8'd159} : s = 186;
	{8'd27,8'd160} : s = 187;
	{8'd27,8'd161} : s = 188;
	{8'd27,8'd162} : s = 189;
	{8'd27,8'd163} : s = 190;
	{8'd27,8'd164} : s = 191;
	{8'd27,8'd165} : s = 192;
	{8'd27,8'd166} : s = 193;
	{8'd27,8'd167} : s = 194;
	{8'd27,8'd168} : s = 195;
	{8'd27,8'd169} : s = 196;
	{8'd27,8'd170} : s = 197;
	{8'd27,8'd171} : s = 198;
	{8'd27,8'd172} : s = 199;
	{8'd27,8'd173} : s = 200;
	{8'd27,8'd174} : s = 201;
	{8'd27,8'd175} : s = 202;
	{8'd27,8'd176} : s = 203;
	{8'd27,8'd177} : s = 204;
	{8'd27,8'd178} : s = 205;
	{8'd27,8'd179} : s = 206;
	{8'd27,8'd180} : s = 207;
	{8'd27,8'd181} : s = 208;
	{8'd27,8'd182} : s = 209;
	{8'd27,8'd183} : s = 210;
	{8'd27,8'd184} : s = 211;
	{8'd27,8'd185} : s = 212;
	{8'd27,8'd186} : s = 213;
	{8'd27,8'd187} : s = 214;
	{8'd27,8'd188} : s = 215;
	{8'd27,8'd189} : s = 216;
	{8'd27,8'd190} : s = 217;
	{8'd27,8'd191} : s = 218;
	{8'd27,8'd192} : s = 219;
	{8'd27,8'd193} : s = 220;
	{8'd27,8'd194} : s = 221;
	{8'd27,8'd195} : s = 222;
	{8'd27,8'd196} : s = 223;
	{8'd27,8'd197} : s = 224;
	{8'd27,8'd198} : s = 225;
	{8'd27,8'd199} : s = 226;
	{8'd27,8'd200} : s = 227;
	{8'd27,8'd201} : s = 228;
	{8'd27,8'd202} : s = 229;
	{8'd27,8'd203} : s = 230;
	{8'd27,8'd204} : s = 231;
	{8'd27,8'd205} : s = 232;
	{8'd27,8'd206} : s = 233;
	{8'd27,8'd207} : s = 234;
	{8'd27,8'd208} : s = 235;
	{8'd27,8'd209} : s = 236;
	{8'd27,8'd210} : s = 237;
	{8'd27,8'd211} : s = 238;
	{8'd27,8'd212} : s = 239;
	{8'd27,8'd213} : s = 240;
	{8'd27,8'd214} : s = 241;
	{8'd27,8'd215} : s = 242;
	{8'd27,8'd216} : s = 243;
	{8'd27,8'd217} : s = 244;
	{8'd27,8'd218} : s = 245;
	{8'd27,8'd219} : s = 246;
	{8'd27,8'd220} : s = 247;
	{8'd27,8'd221} : s = 248;
	{8'd27,8'd222} : s = 249;
	{8'd27,8'd223} : s = 250;
	{8'd27,8'd224} : s = 251;
	{8'd27,8'd225} : s = 252;
	{8'd27,8'd226} : s = 253;
	{8'd27,8'd227} : s = 254;
	{8'd27,8'd228} : s = 255;
	{8'd27,8'd229} : s = 256;
	{8'd27,8'd230} : s = 257;
	{8'd27,8'd231} : s = 258;
	{8'd27,8'd232} : s = 259;
	{8'd27,8'd233} : s = 260;
	{8'd27,8'd234} : s = 261;
	{8'd27,8'd235} : s = 262;
	{8'd27,8'd236} : s = 263;
	{8'd27,8'd237} : s = 264;
	{8'd27,8'd238} : s = 265;
	{8'd27,8'd239} : s = 266;
	{8'd27,8'd240} : s = 267;
	{8'd27,8'd241} : s = 268;
	{8'd27,8'd242} : s = 269;
	{8'd27,8'd243} : s = 270;
	{8'd27,8'd244} : s = 271;
	{8'd27,8'd245} : s = 272;
	{8'd27,8'd246} : s = 273;
	{8'd27,8'd247} : s = 274;
	{8'd27,8'd248} : s = 275;
	{8'd27,8'd249} : s = 276;
	{8'd27,8'd250} : s = 277;
	{8'd27,8'd251} : s = 278;
	{8'd27,8'd252} : s = 279;
	{8'd27,8'd253} : s = 280;
	{8'd27,8'd254} : s = 281;
	{8'd27,8'd255} : s = 282;
	{8'd28,8'd0} : s = 28;
	{8'd28,8'd1} : s = 29;
	{8'd28,8'd2} : s = 30;
	{8'd28,8'd3} : s = 31;
	{8'd28,8'd4} : s = 32;
	{8'd28,8'd5} : s = 33;
	{8'd28,8'd6} : s = 34;
	{8'd28,8'd7} : s = 35;
	{8'd28,8'd8} : s = 36;
	{8'd28,8'd9} : s = 37;
	{8'd28,8'd10} : s = 38;
	{8'd28,8'd11} : s = 39;
	{8'd28,8'd12} : s = 40;
	{8'd28,8'd13} : s = 41;
	{8'd28,8'd14} : s = 42;
	{8'd28,8'd15} : s = 43;
	{8'd28,8'd16} : s = 44;
	{8'd28,8'd17} : s = 45;
	{8'd28,8'd18} : s = 46;
	{8'd28,8'd19} : s = 47;
	{8'd28,8'd20} : s = 48;
	{8'd28,8'd21} : s = 49;
	{8'd28,8'd22} : s = 50;
	{8'd28,8'd23} : s = 51;
	{8'd28,8'd24} : s = 52;
	{8'd28,8'd25} : s = 53;
	{8'd28,8'd26} : s = 54;
	{8'd28,8'd27} : s = 55;
	{8'd28,8'd28} : s = 56;
	{8'd28,8'd29} : s = 57;
	{8'd28,8'd30} : s = 58;
	{8'd28,8'd31} : s = 59;
	{8'd28,8'd32} : s = 60;
	{8'd28,8'd33} : s = 61;
	{8'd28,8'd34} : s = 62;
	{8'd28,8'd35} : s = 63;
	{8'd28,8'd36} : s = 64;
	{8'd28,8'd37} : s = 65;
	{8'd28,8'd38} : s = 66;
	{8'd28,8'd39} : s = 67;
	{8'd28,8'd40} : s = 68;
	{8'd28,8'd41} : s = 69;
	{8'd28,8'd42} : s = 70;
	{8'd28,8'd43} : s = 71;
	{8'd28,8'd44} : s = 72;
	{8'd28,8'd45} : s = 73;
	{8'd28,8'd46} : s = 74;
	{8'd28,8'd47} : s = 75;
	{8'd28,8'd48} : s = 76;
	{8'd28,8'd49} : s = 77;
	{8'd28,8'd50} : s = 78;
	{8'd28,8'd51} : s = 79;
	{8'd28,8'd52} : s = 80;
	{8'd28,8'd53} : s = 81;
	{8'd28,8'd54} : s = 82;
	{8'd28,8'd55} : s = 83;
	{8'd28,8'd56} : s = 84;
	{8'd28,8'd57} : s = 85;
	{8'd28,8'd58} : s = 86;
	{8'd28,8'd59} : s = 87;
	{8'd28,8'd60} : s = 88;
	{8'd28,8'd61} : s = 89;
	{8'd28,8'd62} : s = 90;
	{8'd28,8'd63} : s = 91;
	{8'd28,8'd64} : s = 92;
	{8'd28,8'd65} : s = 93;
	{8'd28,8'd66} : s = 94;
	{8'd28,8'd67} : s = 95;
	{8'd28,8'd68} : s = 96;
	{8'd28,8'd69} : s = 97;
	{8'd28,8'd70} : s = 98;
	{8'd28,8'd71} : s = 99;
	{8'd28,8'd72} : s = 100;
	{8'd28,8'd73} : s = 101;
	{8'd28,8'd74} : s = 102;
	{8'd28,8'd75} : s = 103;
	{8'd28,8'd76} : s = 104;
	{8'd28,8'd77} : s = 105;
	{8'd28,8'd78} : s = 106;
	{8'd28,8'd79} : s = 107;
	{8'd28,8'd80} : s = 108;
	{8'd28,8'd81} : s = 109;
	{8'd28,8'd82} : s = 110;
	{8'd28,8'd83} : s = 111;
	{8'd28,8'd84} : s = 112;
	{8'd28,8'd85} : s = 113;
	{8'd28,8'd86} : s = 114;
	{8'd28,8'd87} : s = 115;
	{8'd28,8'd88} : s = 116;
	{8'd28,8'd89} : s = 117;
	{8'd28,8'd90} : s = 118;
	{8'd28,8'd91} : s = 119;
	{8'd28,8'd92} : s = 120;
	{8'd28,8'd93} : s = 121;
	{8'd28,8'd94} : s = 122;
	{8'd28,8'd95} : s = 123;
	{8'd28,8'd96} : s = 124;
	{8'd28,8'd97} : s = 125;
	{8'd28,8'd98} : s = 126;
	{8'd28,8'd99} : s = 127;
	{8'd28,8'd100} : s = 128;
	{8'd28,8'd101} : s = 129;
	{8'd28,8'd102} : s = 130;
	{8'd28,8'd103} : s = 131;
	{8'd28,8'd104} : s = 132;
	{8'd28,8'd105} : s = 133;
	{8'd28,8'd106} : s = 134;
	{8'd28,8'd107} : s = 135;
	{8'd28,8'd108} : s = 136;
	{8'd28,8'd109} : s = 137;
	{8'd28,8'd110} : s = 138;
	{8'd28,8'd111} : s = 139;
	{8'd28,8'd112} : s = 140;
	{8'd28,8'd113} : s = 141;
	{8'd28,8'd114} : s = 142;
	{8'd28,8'd115} : s = 143;
	{8'd28,8'd116} : s = 144;
	{8'd28,8'd117} : s = 145;
	{8'd28,8'd118} : s = 146;
	{8'd28,8'd119} : s = 147;
	{8'd28,8'd120} : s = 148;
	{8'd28,8'd121} : s = 149;
	{8'd28,8'd122} : s = 150;
	{8'd28,8'd123} : s = 151;
	{8'd28,8'd124} : s = 152;
	{8'd28,8'd125} : s = 153;
	{8'd28,8'd126} : s = 154;
	{8'd28,8'd127} : s = 155;
	{8'd28,8'd128} : s = 156;
	{8'd28,8'd129} : s = 157;
	{8'd28,8'd130} : s = 158;
	{8'd28,8'd131} : s = 159;
	{8'd28,8'd132} : s = 160;
	{8'd28,8'd133} : s = 161;
	{8'd28,8'd134} : s = 162;
	{8'd28,8'd135} : s = 163;
	{8'd28,8'd136} : s = 164;
	{8'd28,8'd137} : s = 165;
	{8'd28,8'd138} : s = 166;
	{8'd28,8'd139} : s = 167;
	{8'd28,8'd140} : s = 168;
	{8'd28,8'd141} : s = 169;
	{8'd28,8'd142} : s = 170;
	{8'd28,8'd143} : s = 171;
	{8'd28,8'd144} : s = 172;
	{8'd28,8'd145} : s = 173;
	{8'd28,8'd146} : s = 174;
	{8'd28,8'd147} : s = 175;
	{8'd28,8'd148} : s = 176;
	{8'd28,8'd149} : s = 177;
	{8'd28,8'd150} : s = 178;
	{8'd28,8'd151} : s = 179;
	{8'd28,8'd152} : s = 180;
	{8'd28,8'd153} : s = 181;
	{8'd28,8'd154} : s = 182;
	{8'd28,8'd155} : s = 183;
	{8'd28,8'd156} : s = 184;
	{8'd28,8'd157} : s = 185;
	{8'd28,8'd158} : s = 186;
	{8'd28,8'd159} : s = 187;
	{8'd28,8'd160} : s = 188;
	{8'd28,8'd161} : s = 189;
	{8'd28,8'd162} : s = 190;
	{8'd28,8'd163} : s = 191;
	{8'd28,8'd164} : s = 192;
	{8'd28,8'd165} : s = 193;
	{8'd28,8'd166} : s = 194;
	{8'd28,8'd167} : s = 195;
	{8'd28,8'd168} : s = 196;
	{8'd28,8'd169} : s = 197;
	{8'd28,8'd170} : s = 198;
	{8'd28,8'd171} : s = 199;
	{8'd28,8'd172} : s = 200;
	{8'd28,8'd173} : s = 201;
	{8'd28,8'd174} : s = 202;
	{8'd28,8'd175} : s = 203;
	{8'd28,8'd176} : s = 204;
	{8'd28,8'd177} : s = 205;
	{8'd28,8'd178} : s = 206;
	{8'd28,8'd179} : s = 207;
	{8'd28,8'd180} : s = 208;
	{8'd28,8'd181} : s = 209;
	{8'd28,8'd182} : s = 210;
	{8'd28,8'd183} : s = 211;
	{8'd28,8'd184} : s = 212;
	{8'd28,8'd185} : s = 213;
	{8'd28,8'd186} : s = 214;
	{8'd28,8'd187} : s = 215;
	{8'd28,8'd188} : s = 216;
	{8'd28,8'd189} : s = 217;
	{8'd28,8'd190} : s = 218;
	{8'd28,8'd191} : s = 219;
	{8'd28,8'd192} : s = 220;
	{8'd28,8'd193} : s = 221;
	{8'd28,8'd194} : s = 222;
	{8'd28,8'd195} : s = 223;
	{8'd28,8'd196} : s = 224;
	{8'd28,8'd197} : s = 225;
	{8'd28,8'd198} : s = 226;
	{8'd28,8'd199} : s = 227;
	{8'd28,8'd200} : s = 228;
	{8'd28,8'd201} : s = 229;
	{8'd28,8'd202} : s = 230;
	{8'd28,8'd203} : s = 231;
	{8'd28,8'd204} : s = 232;
	{8'd28,8'd205} : s = 233;
	{8'd28,8'd206} : s = 234;
	{8'd28,8'd207} : s = 235;
	{8'd28,8'd208} : s = 236;
	{8'd28,8'd209} : s = 237;
	{8'd28,8'd210} : s = 238;
	{8'd28,8'd211} : s = 239;
	{8'd28,8'd212} : s = 240;
	{8'd28,8'd213} : s = 241;
	{8'd28,8'd214} : s = 242;
	{8'd28,8'd215} : s = 243;
	{8'd28,8'd216} : s = 244;
	{8'd28,8'd217} : s = 245;
	{8'd28,8'd218} : s = 246;
	{8'd28,8'd219} : s = 247;
	{8'd28,8'd220} : s = 248;
	{8'd28,8'd221} : s = 249;
	{8'd28,8'd222} : s = 250;
	{8'd28,8'd223} : s = 251;
	{8'd28,8'd224} : s = 252;
	{8'd28,8'd225} : s = 253;
	{8'd28,8'd226} : s = 254;
	{8'd28,8'd227} : s = 255;
	{8'd28,8'd228} : s = 256;
	{8'd28,8'd229} : s = 257;
	{8'd28,8'd230} : s = 258;
	{8'd28,8'd231} : s = 259;
	{8'd28,8'd232} : s = 260;
	{8'd28,8'd233} : s = 261;
	{8'd28,8'd234} : s = 262;
	{8'd28,8'd235} : s = 263;
	{8'd28,8'd236} : s = 264;
	{8'd28,8'd237} : s = 265;
	{8'd28,8'd238} : s = 266;
	{8'd28,8'd239} : s = 267;
	{8'd28,8'd240} : s = 268;
	{8'd28,8'd241} : s = 269;
	{8'd28,8'd242} : s = 270;
	{8'd28,8'd243} : s = 271;
	{8'd28,8'd244} : s = 272;
	{8'd28,8'd245} : s = 273;
	{8'd28,8'd246} : s = 274;
	{8'd28,8'd247} : s = 275;
	{8'd28,8'd248} : s = 276;
	{8'd28,8'd249} : s = 277;
	{8'd28,8'd250} : s = 278;
	{8'd28,8'd251} : s = 279;
	{8'd28,8'd252} : s = 280;
	{8'd28,8'd253} : s = 281;
	{8'd28,8'd254} : s = 282;
	{8'd28,8'd255} : s = 283;
	{8'd29,8'd0} : s = 29;
	{8'd29,8'd1} : s = 30;
	{8'd29,8'd2} : s = 31;
	{8'd29,8'd3} : s = 32;
	{8'd29,8'd4} : s = 33;
	{8'd29,8'd5} : s = 34;
	{8'd29,8'd6} : s = 35;
	{8'd29,8'd7} : s = 36;
	{8'd29,8'd8} : s = 37;
	{8'd29,8'd9} : s = 38;
	{8'd29,8'd10} : s = 39;
	{8'd29,8'd11} : s = 40;
	{8'd29,8'd12} : s = 41;
	{8'd29,8'd13} : s = 42;
	{8'd29,8'd14} : s = 43;
	{8'd29,8'd15} : s = 44;
	{8'd29,8'd16} : s = 45;
	{8'd29,8'd17} : s = 46;
	{8'd29,8'd18} : s = 47;
	{8'd29,8'd19} : s = 48;
	{8'd29,8'd20} : s = 49;
	{8'd29,8'd21} : s = 50;
	{8'd29,8'd22} : s = 51;
	{8'd29,8'd23} : s = 52;
	{8'd29,8'd24} : s = 53;
	{8'd29,8'd25} : s = 54;
	{8'd29,8'd26} : s = 55;
	{8'd29,8'd27} : s = 56;
	{8'd29,8'd28} : s = 57;
	{8'd29,8'd29} : s = 58;
	{8'd29,8'd30} : s = 59;
	{8'd29,8'd31} : s = 60;
	{8'd29,8'd32} : s = 61;
	{8'd29,8'd33} : s = 62;
	{8'd29,8'd34} : s = 63;
	{8'd29,8'd35} : s = 64;
	{8'd29,8'd36} : s = 65;
	{8'd29,8'd37} : s = 66;
	{8'd29,8'd38} : s = 67;
	{8'd29,8'd39} : s = 68;
	{8'd29,8'd40} : s = 69;
	{8'd29,8'd41} : s = 70;
	{8'd29,8'd42} : s = 71;
	{8'd29,8'd43} : s = 72;
	{8'd29,8'd44} : s = 73;
	{8'd29,8'd45} : s = 74;
	{8'd29,8'd46} : s = 75;
	{8'd29,8'd47} : s = 76;
	{8'd29,8'd48} : s = 77;
	{8'd29,8'd49} : s = 78;
	{8'd29,8'd50} : s = 79;
	{8'd29,8'd51} : s = 80;
	{8'd29,8'd52} : s = 81;
	{8'd29,8'd53} : s = 82;
	{8'd29,8'd54} : s = 83;
	{8'd29,8'd55} : s = 84;
	{8'd29,8'd56} : s = 85;
	{8'd29,8'd57} : s = 86;
	{8'd29,8'd58} : s = 87;
	{8'd29,8'd59} : s = 88;
	{8'd29,8'd60} : s = 89;
	{8'd29,8'd61} : s = 90;
	{8'd29,8'd62} : s = 91;
	{8'd29,8'd63} : s = 92;
	{8'd29,8'd64} : s = 93;
	{8'd29,8'd65} : s = 94;
	{8'd29,8'd66} : s = 95;
	{8'd29,8'd67} : s = 96;
	{8'd29,8'd68} : s = 97;
	{8'd29,8'd69} : s = 98;
	{8'd29,8'd70} : s = 99;
	{8'd29,8'd71} : s = 100;
	{8'd29,8'd72} : s = 101;
	{8'd29,8'd73} : s = 102;
	{8'd29,8'd74} : s = 103;
	{8'd29,8'd75} : s = 104;
	{8'd29,8'd76} : s = 105;
	{8'd29,8'd77} : s = 106;
	{8'd29,8'd78} : s = 107;
	{8'd29,8'd79} : s = 108;
	{8'd29,8'd80} : s = 109;
	{8'd29,8'd81} : s = 110;
	{8'd29,8'd82} : s = 111;
	{8'd29,8'd83} : s = 112;
	{8'd29,8'd84} : s = 113;
	{8'd29,8'd85} : s = 114;
	{8'd29,8'd86} : s = 115;
	{8'd29,8'd87} : s = 116;
	{8'd29,8'd88} : s = 117;
	{8'd29,8'd89} : s = 118;
	{8'd29,8'd90} : s = 119;
	{8'd29,8'd91} : s = 120;
	{8'd29,8'd92} : s = 121;
	{8'd29,8'd93} : s = 122;
	{8'd29,8'd94} : s = 123;
	{8'd29,8'd95} : s = 124;
	{8'd29,8'd96} : s = 125;
	{8'd29,8'd97} : s = 126;
	{8'd29,8'd98} : s = 127;
	{8'd29,8'd99} : s = 128;
	{8'd29,8'd100} : s = 129;
	{8'd29,8'd101} : s = 130;
	{8'd29,8'd102} : s = 131;
	{8'd29,8'd103} : s = 132;
	{8'd29,8'd104} : s = 133;
	{8'd29,8'd105} : s = 134;
	{8'd29,8'd106} : s = 135;
	{8'd29,8'd107} : s = 136;
	{8'd29,8'd108} : s = 137;
	{8'd29,8'd109} : s = 138;
	{8'd29,8'd110} : s = 139;
	{8'd29,8'd111} : s = 140;
	{8'd29,8'd112} : s = 141;
	{8'd29,8'd113} : s = 142;
	{8'd29,8'd114} : s = 143;
	{8'd29,8'd115} : s = 144;
	{8'd29,8'd116} : s = 145;
	{8'd29,8'd117} : s = 146;
	{8'd29,8'd118} : s = 147;
	{8'd29,8'd119} : s = 148;
	{8'd29,8'd120} : s = 149;
	{8'd29,8'd121} : s = 150;
	{8'd29,8'd122} : s = 151;
	{8'd29,8'd123} : s = 152;
	{8'd29,8'd124} : s = 153;
	{8'd29,8'd125} : s = 154;
	{8'd29,8'd126} : s = 155;
	{8'd29,8'd127} : s = 156;
	{8'd29,8'd128} : s = 157;
	{8'd29,8'd129} : s = 158;
	{8'd29,8'd130} : s = 159;
	{8'd29,8'd131} : s = 160;
	{8'd29,8'd132} : s = 161;
	{8'd29,8'd133} : s = 162;
	{8'd29,8'd134} : s = 163;
	{8'd29,8'd135} : s = 164;
	{8'd29,8'd136} : s = 165;
	{8'd29,8'd137} : s = 166;
	{8'd29,8'd138} : s = 167;
	{8'd29,8'd139} : s = 168;
	{8'd29,8'd140} : s = 169;
	{8'd29,8'd141} : s = 170;
	{8'd29,8'd142} : s = 171;
	{8'd29,8'd143} : s = 172;
	{8'd29,8'd144} : s = 173;
	{8'd29,8'd145} : s = 174;
	{8'd29,8'd146} : s = 175;
	{8'd29,8'd147} : s = 176;
	{8'd29,8'd148} : s = 177;
	{8'd29,8'd149} : s = 178;
	{8'd29,8'd150} : s = 179;
	{8'd29,8'd151} : s = 180;
	{8'd29,8'd152} : s = 181;
	{8'd29,8'd153} : s = 182;
	{8'd29,8'd154} : s = 183;
	{8'd29,8'd155} : s = 184;
	{8'd29,8'd156} : s = 185;
	{8'd29,8'd157} : s = 186;
	{8'd29,8'd158} : s = 187;
	{8'd29,8'd159} : s = 188;
	{8'd29,8'd160} : s = 189;
	{8'd29,8'd161} : s = 190;
	{8'd29,8'd162} : s = 191;
	{8'd29,8'd163} : s = 192;
	{8'd29,8'd164} : s = 193;
	{8'd29,8'd165} : s = 194;
	{8'd29,8'd166} : s = 195;
	{8'd29,8'd167} : s = 196;
	{8'd29,8'd168} : s = 197;
	{8'd29,8'd169} : s = 198;
	{8'd29,8'd170} : s = 199;
	{8'd29,8'd171} : s = 200;
	{8'd29,8'd172} : s = 201;
	{8'd29,8'd173} : s = 202;
	{8'd29,8'd174} : s = 203;
	{8'd29,8'd175} : s = 204;
	{8'd29,8'd176} : s = 205;
	{8'd29,8'd177} : s = 206;
	{8'd29,8'd178} : s = 207;
	{8'd29,8'd179} : s = 208;
	{8'd29,8'd180} : s = 209;
	{8'd29,8'd181} : s = 210;
	{8'd29,8'd182} : s = 211;
	{8'd29,8'd183} : s = 212;
	{8'd29,8'd184} : s = 213;
	{8'd29,8'd185} : s = 214;
	{8'd29,8'd186} : s = 215;
	{8'd29,8'd187} : s = 216;
	{8'd29,8'd188} : s = 217;
	{8'd29,8'd189} : s = 218;
	{8'd29,8'd190} : s = 219;
	{8'd29,8'd191} : s = 220;
	{8'd29,8'd192} : s = 221;
	{8'd29,8'd193} : s = 222;
	{8'd29,8'd194} : s = 223;
	{8'd29,8'd195} : s = 224;
	{8'd29,8'd196} : s = 225;
	{8'd29,8'd197} : s = 226;
	{8'd29,8'd198} : s = 227;
	{8'd29,8'd199} : s = 228;
	{8'd29,8'd200} : s = 229;
	{8'd29,8'd201} : s = 230;
	{8'd29,8'd202} : s = 231;
	{8'd29,8'd203} : s = 232;
	{8'd29,8'd204} : s = 233;
	{8'd29,8'd205} : s = 234;
	{8'd29,8'd206} : s = 235;
	{8'd29,8'd207} : s = 236;
	{8'd29,8'd208} : s = 237;
	{8'd29,8'd209} : s = 238;
	{8'd29,8'd210} : s = 239;
	{8'd29,8'd211} : s = 240;
	{8'd29,8'd212} : s = 241;
	{8'd29,8'd213} : s = 242;
	{8'd29,8'd214} : s = 243;
	{8'd29,8'd215} : s = 244;
	{8'd29,8'd216} : s = 245;
	{8'd29,8'd217} : s = 246;
	{8'd29,8'd218} : s = 247;
	{8'd29,8'd219} : s = 248;
	{8'd29,8'd220} : s = 249;
	{8'd29,8'd221} : s = 250;
	{8'd29,8'd222} : s = 251;
	{8'd29,8'd223} : s = 252;
	{8'd29,8'd224} : s = 253;
	{8'd29,8'd225} : s = 254;
	{8'd29,8'd226} : s = 255;
	{8'd29,8'd227} : s = 256;
	{8'd29,8'd228} : s = 257;
	{8'd29,8'd229} : s = 258;
	{8'd29,8'd230} : s = 259;
	{8'd29,8'd231} : s = 260;
	{8'd29,8'd232} : s = 261;
	{8'd29,8'd233} : s = 262;
	{8'd29,8'd234} : s = 263;
	{8'd29,8'd235} : s = 264;
	{8'd29,8'd236} : s = 265;
	{8'd29,8'd237} : s = 266;
	{8'd29,8'd238} : s = 267;
	{8'd29,8'd239} : s = 268;
	{8'd29,8'd240} : s = 269;
	{8'd29,8'd241} : s = 270;
	{8'd29,8'd242} : s = 271;
	{8'd29,8'd243} : s = 272;
	{8'd29,8'd244} : s = 273;
	{8'd29,8'd245} : s = 274;
	{8'd29,8'd246} : s = 275;
	{8'd29,8'd247} : s = 276;
	{8'd29,8'd248} : s = 277;
	{8'd29,8'd249} : s = 278;
	{8'd29,8'd250} : s = 279;
	{8'd29,8'd251} : s = 280;
	{8'd29,8'd252} : s = 281;
	{8'd29,8'd253} : s = 282;
	{8'd29,8'd254} : s = 283;
	{8'd29,8'd255} : s = 284;
	{8'd30,8'd0} : s = 30;
	{8'd30,8'd1} : s = 31;
	{8'd30,8'd2} : s = 32;
	{8'd30,8'd3} : s = 33;
	{8'd30,8'd4} : s = 34;
	{8'd30,8'd5} : s = 35;
	{8'd30,8'd6} : s = 36;
	{8'd30,8'd7} : s = 37;
	{8'd30,8'd8} : s = 38;
	{8'd30,8'd9} : s = 39;
	{8'd30,8'd10} : s = 40;
	{8'd30,8'd11} : s = 41;
	{8'd30,8'd12} : s = 42;
	{8'd30,8'd13} : s = 43;
	{8'd30,8'd14} : s = 44;
	{8'd30,8'd15} : s = 45;
	{8'd30,8'd16} : s = 46;
	{8'd30,8'd17} : s = 47;
	{8'd30,8'd18} : s = 48;
	{8'd30,8'd19} : s = 49;
	{8'd30,8'd20} : s = 50;
	{8'd30,8'd21} : s = 51;
	{8'd30,8'd22} : s = 52;
	{8'd30,8'd23} : s = 53;
	{8'd30,8'd24} : s = 54;
	{8'd30,8'd25} : s = 55;
	{8'd30,8'd26} : s = 56;
	{8'd30,8'd27} : s = 57;
	{8'd30,8'd28} : s = 58;
	{8'd30,8'd29} : s = 59;
	{8'd30,8'd30} : s = 60;
	{8'd30,8'd31} : s = 61;
	{8'd30,8'd32} : s = 62;
	{8'd30,8'd33} : s = 63;
	{8'd30,8'd34} : s = 64;
	{8'd30,8'd35} : s = 65;
	{8'd30,8'd36} : s = 66;
	{8'd30,8'd37} : s = 67;
	{8'd30,8'd38} : s = 68;
	{8'd30,8'd39} : s = 69;
	{8'd30,8'd40} : s = 70;
	{8'd30,8'd41} : s = 71;
	{8'd30,8'd42} : s = 72;
	{8'd30,8'd43} : s = 73;
	{8'd30,8'd44} : s = 74;
	{8'd30,8'd45} : s = 75;
	{8'd30,8'd46} : s = 76;
	{8'd30,8'd47} : s = 77;
	{8'd30,8'd48} : s = 78;
	{8'd30,8'd49} : s = 79;
	{8'd30,8'd50} : s = 80;
	{8'd30,8'd51} : s = 81;
	{8'd30,8'd52} : s = 82;
	{8'd30,8'd53} : s = 83;
	{8'd30,8'd54} : s = 84;
	{8'd30,8'd55} : s = 85;
	{8'd30,8'd56} : s = 86;
	{8'd30,8'd57} : s = 87;
	{8'd30,8'd58} : s = 88;
	{8'd30,8'd59} : s = 89;
	{8'd30,8'd60} : s = 90;
	{8'd30,8'd61} : s = 91;
	{8'd30,8'd62} : s = 92;
	{8'd30,8'd63} : s = 93;
	{8'd30,8'd64} : s = 94;
	{8'd30,8'd65} : s = 95;
	{8'd30,8'd66} : s = 96;
	{8'd30,8'd67} : s = 97;
	{8'd30,8'd68} : s = 98;
	{8'd30,8'd69} : s = 99;
	{8'd30,8'd70} : s = 100;
	{8'd30,8'd71} : s = 101;
	{8'd30,8'd72} : s = 102;
	{8'd30,8'd73} : s = 103;
	{8'd30,8'd74} : s = 104;
	{8'd30,8'd75} : s = 105;
	{8'd30,8'd76} : s = 106;
	{8'd30,8'd77} : s = 107;
	{8'd30,8'd78} : s = 108;
	{8'd30,8'd79} : s = 109;
	{8'd30,8'd80} : s = 110;
	{8'd30,8'd81} : s = 111;
	{8'd30,8'd82} : s = 112;
	{8'd30,8'd83} : s = 113;
	{8'd30,8'd84} : s = 114;
	{8'd30,8'd85} : s = 115;
	{8'd30,8'd86} : s = 116;
	{8'd30,8'd87} : s = 117;
	{8'd30,8'd88} : s = 118;
	{8'd30,8'd89} : s = 119;
	{8'd30,8'd90} : s = 120;
	{8'd30,8'd91} : s = 121;
	{8'd30,8'd92} : s = 122;
	{8'd30,8'd93} : s = 123;
	{8'd30,8'd94} : s = 124;
	{8'd30,8'd95} : s = 125;
	{8'd30,8'd96} : s = 126;
	{8'd30,8'd97} : s = 127;
	{8'd30,8'd98} : s = 128;
	{8'd30,8'd99} : s = 129;
	{8'd30,8'd100} : s = 130;
	{8'd30,8'd101} : s = 131;
	{8'd30,8'd102} : s = 132;
	{8'd30,8'd103} : s = 133;
	{8'd30,8'd104} : s = 134;
	{8'd30,8'd105} : s = 135;
	{8'd30,8'd106} : s = 136;
	{8'd30,8'd107} : s = 137;
	{8'd30,8'd108} : s = 138;
	{8'd30,8'd109} : s = 139;
	{8'd30,8'd110} : s = 140;
	{8'd30,8'd111} : s = 141;
	{8'd30,8'd112} : s = 142;
	{8'd30,8'd113} : s = 143;
	{8'd30,8'd114} : s = 144;
	{8'd30,8'd115} : s = 145;
	{8'd30,8'd116} : s = 146;
	{8'd30,8'd117} : s = 147;
	{8'd30,8'd118} : s = 148;
	{8'd30,8'd119} : s = 149;
	{8'd30,8'd120} : s = 150;
	{8'd30,8'd121} : s = 151;
	{8'd30,8'd122} : s = 152;
	{8'd30,8'd123} : s = 153;
	{8'd30,8'd124} : s = 154;
	{8'd30,8'd125} : s = 155;
	{8'd30,8'd126} : s = 156;
	{8'd30,8'd127} : s = 157;
	{8'd30,8'd128} : s = 158;
	{8'd30,8'd129} : s = 159;
	{8'd30,8'd130} : s = 160;
	{8'd30,8'd131} : s = 161;
	{8'd30,8'd132} : s = 162;
	{8'd30,8'd133} : s = 163;
	{8'd30,8'd134} : s = 164;
	{8'd30,8'd135} : s = 165;
	{8'd30,8'd136} : s = 166;
	{8'd30,8'd137} : s = 167;
	{8'd30,8'd138} : s = 168;
	{8'd30,8'd139} : s = 169;
	{8'd30,8'd140} : s = 170;
	{8'd30,8'd141} : s = 171;
	{8'd30,8'd142} : s = 172;
	{8'd30,8'd143} : s = 173;
	{8'd30,8'd144} : s = 174;
	{8'd30,8'd145} : s = 175;
	{8'd30,8'd146} : s = 176;
	{8'd30,8'd147} : s = 177;
	{8'd30,8'd148} : s = 178;
	{8'd30,8'd149} : s = 179;
	{8'd30,8'd150} : s = 180;
	{8'd30,8'd151} : s = 181;
	{8'd30,8'd152} : s = 182;
	{8'd30,8'd153} : s = 183;
	{8'd30,8'd154} : s = 184;
	{8'd30,8'd155} : s = 185;
	{8'd30,8'd156} : s = 186;
	{8'd30,8'd157} : s = 187;
	{8'd30,8'd158} : s = 188;
	{8'd30,8'd159} : s = 189;
	{8'd30,8'd160} : s = 190;
	{8'd30,8'd161} : s = 191;
	{8'd30,8'd162} : s = 192;
	{8'd30,8'd163} : s = 193;
	{8'd30,8'd164} : s = 194;
	{8'd30,8'd165} : s = 195;
	{8'd30,8'd166} : s = 196;
	{8'd30,8'd167} : s = 197;
	{8'd30,8'd168} : s = 198;
	{8'd30,8'd169} : s = 199;
	{8'd30,8'd170} : s = 200;
	{8'd30,8'd171} : s = 201;
	{8'd30,8'd172} : s = 202;
	{8'd30,8'd173} : s = 203;
	{8'd30,8'd174} : s = 204;
	{8'd30,8'd175} : s = 205;
	{8'd30,8'd176} : s = 206;
	{8'd30,8'd177} : s = 207;
	{8'd30,8'd178} : s = 208;
	{8'd30,8'd179} : s = 209;
	{8'd30,8'd180} : s = 210;
	{8'd30,8'd181} : s = 211;
	{8'd30,8'd182} : s = 212;
	{8'd30,8'd183} : s = 213;
	{8'd30,8'd184} : s = 214;
	{8'd30,8'd185} : s = 215;
	{8'd30,8'd186} : s = 216;
	{8'd30,8'd187} : s = 217;
	{8'd30,8'd188} : s = 218;
	{8'd30,8'd189} : s = 219;
	{8'd30,8'd190} : s = 220;
	{8'd30,8'd191} : s = 221;
	{8'd30,8'd192} : s = 222;
	{8'd30,8'd193} : s = 223;
	{8'd30,8'd194} : s = 224;
	{8'd30,8'd195} : s = 225;
	{8'd30,8'd196} : s = 226;
	{8'd30,8'd197} : s = 227;
	{8'd30,8'd198} : s = 228;
	{8'd30,8'd199} : s = 229;
	{8'd30,8'd200} : s = 230;
	{8'd30,8'd201} : s = 231;
	{8'd30,8'd202} : s = 232;
	{8'd30,8'd203} : s = 233;
	{8'd30,8'd204} : s = 234;
	{8'd30,8'd205} : s = 235;
	{8'd30,8'd206} : s = 236;
	{8'd30,8'd207} : s = 237;
	{8'd30,8'd208} : s = 238;
	{8'd30,8'd209} : s = 239;
	{8'd30,8'd210} : s = 240;
	{8'd30,8'd211} : s = 241;
	{8'd30,8'd212} : s = 242;
	{8'd30,8'd213} : s = 243;
	{8'd30,8'd214} : s = 244;
	{8'd30,8'd215} : s = 245;
	{8'd30,8'd216} : s = 246;
	{8'd30,8'd217} : s = 247;
	{8'd30,8'd218} : s = 248;
	{8'd30,8'd219} : s = 249;
	{8'd30,8'd220} : s = 250;
	{8'd30,8'd221} : s = 251;
	{8'd30,8'd222} : s = 252;
	{8'd30,8'd223} : s = 253;
	{8'd30,8'd224} : s = 254;
	{8'd30,8'd225} : s = 255;
	{8'd30,8'd226} : s = 256;
	{8'd30,8'd227} : s = 257;
	{8'd30,8'd228} : s = 258;
	{8'd30,8'd229} : s = 259;
	{8'd30,8'd230} : s = 260;
	{8'd30,8'd231} : s = 261;
	{8'd30,8'd232} : s = 262;
	{8'd30,8'd233} : s = 263;
	{8'd30,8'd234} : s = 264;
	{8'd30,8'd235} : s = 265;
	{8'd30,8'd236} : s = 266;
	{8'd30,8'd237} : s = 267;
	{8'd30,8'd238} : s = 268;
	{8'd30,8'd239} : s = 269;
	{8'd30,8'd240} : s = 270;
	{8'd30,8'd241} : s = 271;
	{8'd30,8'd242} : s = 272;
	{8'd30,8'd243} : s = 273;
	{8'd30,8'd244} : s = 274;
	{8'd30,8'd245} : s = 275;
	{8'd30,8'd246} : s = 276;
	{8'd30,8'd247} : s = 277;
	{8'd30,8'd248} : s = 278;
	{8'd30,8'd249} : s = 279;
	{8'd30,8'd250} : s = 280;
	{8'd30,8'd251} : s = 281;
	{8'd30,8'd252} : s = 282;
	{8'd30,8'd253} : s = 283;
	{8'd30,8'd254} : s = 284;
	{8'd30,8'd255} : s = 285;
	{8'd31,8'd0} : s = 31;
	{8'd31,8'd1} : s = 32;
	{8'd31,8'd2} : s = 33;
	{8'd31,8'd3} : s = 34;
	{8'd31,8'd4} : s = 35;
	{8'd31,8'd5} : s = 36;
	{8'd31,8'd6} : s = 37;
	{8'd31,8'd7} : s = 38;
	{8'd31,8'd8} : s = 39;
	{8'd31,8'd9} : s = 40;
	{8'd31,8'd10} : s = 41;
	{8'd31,8'd11} : s = 42;
	{8'd31,8'd12} : s = 43;
	{8'd31,8'd13} : s = 44;
	{8'd31,8'd14} : s = 45;
	{8'd31,8'd15} : s = 46;
	{8'd31,8'd16} : s = 47;
	{8'd31,8'd17} : s = 48;
	{8'd31,8'd18} : s = 49;
	{8'd31,8'd19} : s = 50;
	{8'd31,8'd20} : s = 51;
	{8'd31,8'd21} : s = 52;
	{8'd31,8'd22} : s = 53;
	{8'd31,8'd23} : s = 54;
	{8'd31,8'd24} : s = 55;
	{8'd31,8'd25} : s = 56;
	{8'd31,8'd26} : s = 57;
	{8'd31,8'd27} : s = 58;
	{8'd31,8'd28} : s = 59;
	{8'd31,8'd29} : s = 60;
	{8'd31,8'd30} : s = 61;
	{8'd31,8'd31} : s = 62;
	{8'd31,8'd32} : s = 63;
	{8'd31,8'd33} : s = 64;
	{8'd31,8'd34} : s = 65;
	{8'd31,8'd35} : s = 66;
	{8'd31,8'd36} : s = 67;
	{8'd31,8'd37} : s = 68;
	{8'd31,8'd38} : s = 69;
	{8'd31,8'd39} : s = 70;
	{8'd31,8'd40} : s = 71;
	{8'd31,8'd41} : s = 72;
	{8'd31,8'd42} : s = 73;
	{8'd31,8'd43} : s = 74;
	{8'd31,8'd44} : s = 75;
	{8'd31,8'd45} : s = 76;
	{8'd31,8'd46} : s = 77;
	{8'd31,8'd47} : s = 78;
	{8'd31,8'd48} : s = 79;
	{8'd31,8'd49} : s = 80;
	{8'd31,8'd50} : s = 81;
	{8'd31,8'd51} : s = 82;
	{8'd31,8'd52} : s = 83;
	{8'd31,8'd53} : s = 84;
	{8'd31,8'd54} : s = 85;
	{8'd31,8'd55} : s = 86;
	{8'd31,8'd56} : s = 87;
	{8'd31,8'd57} : s = 88;
	{8'd31,8'd58} : s = 89;
	{8'd31,8'd59} : s = 90;
	{8'd31,8'd60} : s = 91;
	{8'd31,8'd61} : s = 92;
	{8'd31,8'd62} : s = 93;
	{8'd31,8'd63} : s = 94;
	{8'd31,8'd64} : s = 95;
	{8'd31,8'd65} : s = 96;
	{8'd31,8'd66} : s = 97;
	{8'd31,8'd67} : s = 98;
	{8'd31,8'd68} : s = 99;
	{8'd31,8'd69} : s = 100;
	{8'd31,8'd70} : s = 101;
	{8'd31,8'd71} : s = 102;
	{8'd31,8'd72} : s = 103;
	{8'd31,8'd73} : s = 104;
	{8'd31,8'd74} : s = 105;
	{8'd31,8'd75} : s = 106;
	{8'd31,8'd76} : s = 107;
	{8'd31,8'd77} : s = 108;
	{8'd31,8'd78} : s = 109;
	{8'd31,8'd79} : s = 110;
	{8'd31,8'd80} : s = 111;
	{8'd31,8'd81} : s = 112;
	{8'd31,8'd82} : s = 113;
	{8'd31,8'd83} : s = 114;
	{8'd31,8'd84} : s = 115;
	{8'd31,8'd85} : s = 116;
	{8'd31,8'd86} : s = 117;
	{8'd31,8'd87} : s = 118;
	{8'd31,8'd88} : s = 119;
	{8'd31,8'd89} : s = 120;
	{8'd31,8'd90} : s = 121;
	{8'd31,8'd91} : s = 122;
	{8'd31,8'd92} : s = 123;
	{8'd31,8'd93} : s = 124;
	{8'd31,8'd94} : s = 125;
	{8'd31,8'd95} : s = 126;
	{8'd31,8'd96} : s = 127;
	{8'd31,8'd97} : s = 128;
	{8'd31,8'd98} : s = 129;
	{8'd31,8'd99} : s = 130;
	{8'd31,8'd100} : s = 131;
	{8'd31,8'd101} : s = 132;
	{8'd31,8'd102} : s = 133;
	{8'd31,8'd103} : s = 134;
	{8'd31,8'd104} : s = 135;
	{8'd31,8'd105} : s = 136;
	{8'd31,8'd106} : s = 137;
	{8'd31,8'd107} : s = 138;
	{8'd31,8'd108} : s = 139;
	{8'd31,8'd109} : s = 140;
	{8'd31,8'd110} : s = 141;
	{8'd31,8'd111} : s = 142;
	{8'd31,8'd112} : s = 143;
	{8'd31,8'd113} : s = 144;
	{8'd31,8'd114} : s = 145;
	{8'd31,8'd115} : s = 146;
	{8'd31,8'd116} : s = 147;
	{8'd31,8'd117} : s = 148;
	{8'd31,8'd118} : s = 149;
	{8'd31,8'd119} : s = 150;
	{8'd31,8'd120} : s = 151;
	{8'd31,8'd121} : s = 152;
	{8'd31,8'd122} : s = 153;
	{8'd31,8'd123} : s = 154;
	{8'd31,8'd124} : s = 155;
	{8'd31,8'd125} : s = 156;
	{8'd31,8'd126} : s = 157;
	{8'd31,8'd127} : s = 158;
	{8'd31,8'd128} : s = 159;
	{8'd31,8'd129} : s = 160;
	{8'd31,8'd130} : s = 161;
	{8'd31,8'd131} : s = 162;
	{8'd31,8'd132} : s = 163;
	{8'd31,8'd133} : s = 164;
	{8'd31,8'd134} : s = 165;
	{8'd31,8'd135} : s = 166;
	{8'd31,8'd136} : s = 167;
	{8'd31,8'd137} : s = 168;
	{8'd31,8'd138} : s = 169;
	{8'd31,8'd139} : s = 170;
	{8'd31,8'd140} : s = 171;
	{8'd31,8'd141} : s = 172;
	{8'd31,8'd142} : s = 173;
	{8'd31,8'd143} : s = 174;
	{8'd31,8'd144} : s = 175;
	{8'd31,8'd145} : s = 176;
	{8'd31,8'd146} : s = 177;
	{8'd31,8'd147} : s = 178;
	{8'd31,8'd148} : s = 179;
	{8'd31,8'd149} : s = 180;
	{8'd31,8'd150} : s = 181;
	{8'd31,8'd151} : s = 182;
	{8'd31,8'd152} : s = 183;
	{8'd31,8'd153} : s = 184;
	{8'd31,8'd154} : s = 185;
	{8'd31,8'd155} : s = 186;
	{8'd31,8'd156} : s = 187;
	{8'd31,8'd157} : s = 188;
	{8'd31,8'd158} : s = 189;
	{8'd31,8'd159} : s = 190;
	{8'd31,8'd160} : s = 191;
	{8'd31,8'd161} : s = 192;
	{8'd31,8'd162} : s = 193;
	{8'd31,8'd163} : s = 194;
	{8'd31,8'd164} : s = 195;
	{8'd31,8'd165} : s = 196;
	{8'd31,8'd166} : s = 197;
	{8'd31,8'd167} : s = 198;
	{8'd31,8'd168} : s = 199;
	{8'd31,8'd169} : s = 200;
	{8'd31,8'd170} : s = 201;
	{8'd31,8'd171} : s = 202;
	{8'd31,8'd172} : s = 203;
	{8'd31,8'd173} : s = 204;
	{8'd31,8'd174} : s = 205;
	{8'd31,8'd175} : s = 206;
	{8'd31,8'd176} : s = 207;
	{8'd31,8'd177} : s = 208;
	{8'd31,8'd178} : s = 209;
	{8'd31,8'd179} : s = 210;
	{8'd31,8'd180} : s = 211;
	{8'd31,8'd181} : s = 212;
	{8'd31,8'd182} : s = 213;
	{8'd31,8'd183} : s = 214;
	{8'd31,8'd184} : s = 215;
	{8'd31,8'd185} : s = 216;
	{8'd31,8'd186} : s = 217;
	{8'd31,8'd187} : s = 218;
	{8'd31,8'd188} : s = 219;
	{8'd31,8'd189} : s = 220;
	{8'd31,8'd190} : s = 221;
	{8'd31,8'd191} : s = 222;
	{8'd31,8'd192} : s = 223;
	{8'd31,8'd193} : s = 224;
	{8'd31,8'd194} : s = 225;
	{8'd31,8'd195} : s = 226;
	{8'd31,8'd196} : s = 227;
	{8'd31,8'd197} : s = 228;
	{8'd31,8'd198} : s = 229;
	{8'd31,8'd199} : s = 230;
	{8'd31,8'd200} : s = 231;
	{8'd31,8'd201} : s = 232;
	{8'd31,8'd202} : s = 233;
	{8'd31,8'd203} : s = 234;
	{8'd31,8'd204} : s = 235;
	{8'd31,8'd205} : s = 236;
	{8'd31,8'd206} : s = 237;
	{8'd31,8'd207} : s = 238;
	{8'd31,8'd208} : s = 239;
	{8'd31,8'd209} : s = 240;
	{8'd31,8'd210} : s = 241;
	{8'd31,8'd211} : s = 242;
	{8'd31,8'd212} : s = 243;
	{8'd31,8'd213} : s = 244;
	{8'd31,8'd214} : s = 245;
	{8'd31,8'd215} : s = 246;
	{8'd31,8'd216} : s = 247;
	{8'd31,8'd217} : s = 248;
	{8'd31,8'd218} : s = 249;
	{8'd31,8'd219} : s = 250;
	{8'd31,8'd220} : s = 251;
	{8'd31,8'd221} : s = 252;
	{8'd31,8'd222} : s = 253;
	{8'd31,8'd223} : s = 254;
	{8'd31,8'd224} : s = 255;
	{8'd31,8'd225} : s = 256;
	{8'd31,8'd226} : s = 257;
	{8'd31,8'd227} : s = 258;
	{8'd31,8'd228} : s = 259;
	{8'd31,8'd229} : s = 260;
	{8'd31,8'd230} : s = 261;
	{8'd31,8'd231} : s = 262;
	{8'd31,8'd232} : s = 263;
	{8'd31,8'd233} : s = 264;
	{8'd31,8'd234} : s = 265;
	{8'd31,8'd235} : s = 266;
	{8'd31,8'd236} : s = 267;
	{8'd31,8'd237} : s = 268;
	{8'd31,8'd238} : s = 269;
	{8'd31,8'd239} : s = 270;
	{8'd31,8'd240} : s = 271;
	{8'd31,8'd241} : s = 272;
	{8'd31,8'd242} : s = 273;
	{8'd31,8'd243} : s = 274;
	{8'd31,8'd244} : s = 275;
	{8'd31,8'd245} : s = 276;
	{8'd31,8'd246} : s = 277;
	{8'd31,8'd247} : s = 278;
	{8'd31,8'd248} : s = 279;
	{8'd31,8'd249} : s = 280;
	{8'd31,8'd250} : s = 281;
	{8'd31,8'd251} : s = 282;
	{8'd31,8'd252} : s = 283;
	{8'd31,8'd253} : s = 284;
	{8'd31,8'd254} : s = 285;
	{8'd31,8'd255} : s = 286;
	{8'd32,8'd0} : s = 32;
	{8'd32,8'd1} : s = 33;
	{8'd32,8'd2} : s = 34;
	{8'd32,8'd3} : s = 35;
	{8'd32,8'd4} : s = 36;
	{8'd32,8'd5} : s = 37;
	{8'd32,8'd6} : s = 38;
	{8'd32,8'd7} : s = 39;
	{8'd32,8'd8} : s = 40;
	{8'd32,8'd9} : s = 41;
	{8'd32,8'd10} : s = 42;
	{8'd32,8'd11} : s = 43;
	{8'd32,8'd12} : s = 44;
	{8'd32,8'd13} : s = 45;
	{8'd32,8'd14} : s = 46;
	{8'd32,8'd15} : s = 47;
	{8'd32,8'd16} : s = 48;
	{8'd32,8'd17} : s = 49;
	{8'd32,8'd18} : s = 50;
	{8'd32,8'd19} : s = 51;
	{8'd32,8'd20} : s = 52;
	{8'd32,8'd21} : s = 53;
	{8'd32,8'd22} : s = 54;
	{8'd32,8'd23} : s = 55;
	{8'd32,8'd24} : s = 56;
	{8'd32,8'd25} : s = 57;
	{8'd32,8'd26} : s = 58;
	{8'd32,8'd27} : s = 59;
	{8'd32,8'd28} : s = 60;
	{8'd32,8'd29} : s = 61;
	{8'd32,8'd30} : s = 62;
	{8'd32,8'd31} : s = 63;
	{8'd32,8'd32} : s = 64;
	{8'd32,8'd33} : s = 65;
	{8'd32,8'd34} : s = 66;
	{8'd32,8'd35} : s = 67;
	{8'd32,8'd36} : s = 68;
	{8'd32,8'd37} : s = 69;
	{8'd32,8'd38} : s = 70;
	{8'd32,8'd39} : s = 71;
	{8'd32,8'd40} : s = 72;
	{8'd32,8'd41} : s = 73;
	{8'd32,8'd42} : s = 74;
	{8'd32,8'd43} : s = 75;
	{8'd32,8'd44} : s = 76;
	{8'd32,8'd45} : s = 77;
	{8'd32,8'd46} : s = 78;
	{8'd32,8'd47} : s = 79;
	{8'd32,8'd48} : s = 80;
	{8'd32,8'd49} : s = 81;
	{8'd32,8'd50} : s = 82;
	{8'd32,8'd51} : s = 83;
	{8'd32,8'd52} : s = 84;
	{8'd32,8'd53} : s = 85;
	{8'd32,8'd54} : s = 86;
	{8'd32,8'd55} : s = 87;
	{8'd32,8'd56} : s = 88;
	{8'd32,8'd57} : s = 89;
	{8'd32,8'd58} : s = 90;
	{8'd32,8'd59} : s = 91;
	{8'd32,8'd60} : s = 92;
	{8'd32,8'd61} : s = 93;
	{8'd32,8'd62} : s = 94;
	{8'd32,8'd63} : s = 95;
	{8'd32,8'd64} : s = 96;
	{8'd32,8'd65} : s = 97;
	{8'd32,8'd66} : s = 98;
	{8'd32,8'd67} : s = 99;
	{8'd32,8'd68} : s = 100;
	{8'd32,8'd69} : s = 101;
	{8'd32,8'd70} : s = 102;
	{8'd32,8'd71} : s = 103;
	{8'd32,8'd72} : s = 104;
	{8'd32,8'd73} : s = 105;
	{8'd32,8'd74} : s = 106;
	{8'd32,8'd75} : s = 107;
	{8'd32,8'd76} : s = 108;
	{8'd32,8'd77} : s = 109;
	{8'd32,8'd78} : s = 110;
	{8'd32,8'd79} : s = 111;
	{8'd32,8'd80} : s = 112;
	{8'd32,8'd81} : s = 113;
	{8'd32,8'd82} : s = 114;
	{8'd32,8'd83} : s = 115;
	{8'd32,8'd84} : s = 116;
	{8'd32,8'd85} : s = 117;
	{8'd32,8'd86} : s = 118;
	{8'd32,8'd87} : s = 119;
	{8'd32,8'd88} : s = 120;
	{8'd32,8'd89} : s = 121;
	{8'd32,8'd90} : s = 122;
	{8'd32,8'd91} : s = 123;
	{8'd32,8'd92} : s = 124;
	{8'd32,8'd93} : s = 125;
	{8'd32,8'd94} : s = 126;
	{8'd32,8'd95} : s = 127;
	{8'd32,8'd96} : s = 128;
	{8'd32,8'd97} : s = 129;
	{8'd32,8'd98} : s = 130;
	{8'd32,8'd99} : s = 131;
	{8'd32,8'd100} : s = 132;
	{8'd32,8'd101} : s = 133;
	{8'd32,8'd102} : s = 134;
	{8'd32,8'd103} : s = 135;
	{8'd32,8'd104} : s = 136;
	{8'd32,8'd105} : s = 137;
	{8'd32,8'd106} : s = 138;
	{8'd32,8'd107} : s = 139;
	{8'd32,8'd108} : s = 140;
	{8'd32,8'd109} : s = 141;
	{8'd32,8'd110} : s = 142;
	{8'd32,8'd111} : s = 143;
	{8'd32,8'd112} : s = 144;
	{8'd32,8'd113} : s = 145;
	{8'd32,8'd114} : s = 146;
	{8'd32,8'd115} : s = 147;
	{8'd32,8'd116} : s = 148;
	{8'd32,8'd117} : s = 149;
	{8'd32,8'd118} : s = 150;
	{8'd32,8'd119} : s = 151;
	{8'd32,8'd120} : s = 152;
	{8'd32,8'd121} : s = 153;
	{8'd32,8'd122} : s = 154;
	{8'd32,8'd123} : s = 155;
	{8'd32,8'd124} : s = 156;
	{8'd32,8'd125} : s = 157;
	{8'd32,8'd126} : s = 158;
	{8'd32,8'd127} : s = 159;
	{8'd32,8'd128} : s = 160;
	{8'd32,8'd129} : s = 161;
	{8'd32,8'd130} : s = 162;
	{8'd32,8'd131} : s = 163;
	{8'd32,8'd132} : s = 164;
	{8'd32,8'd133} : s = 165;
	{8'd32,8'd134} : s = 166;
	{8'd32,8'd135} : s = 167;
	{8'd32,8'd136} : s = 168;
	{8'd32,8'd137} : s = 169;
	{8'd32,8'd138} : s = 170;
	{8'd32,8'd139} : s = 171;
	{8'd32,8'd140} : s = 172;
	{8'd32,8'd141} : s = 173;
	{8'd32,8'd142} : s = 174;
	{8'd32,8'd143} : s = 175;
	{8'd32,8'd144} : s = 176;
	{8'd32,8'd145} : s = 177;
	{8'd32,8'd146} : s = 178;
	{8'd32,8'd147} : s = 179;
	{8'd32,8'd148} : s = 180;
	{8'd32,8'd149} : s = 181;
	{8'd32,8'd150} : s = 182;
	{8'd32,8'd151} : s = 183;
	{8'd32,8'd152} : s = 184;
	{8'd32,8'd153} : s = 185;
	{8'd32,8'd154} : s = 186;
	{8'd32,8'd155} : s = 187;
	{8'd32,8'd156} : s = 188;
	{8'd32,8'd157} : s = 189;
	{8'd32,8'd158} : s = 190;
	{8'd32,8'd159} : s = 191;
	{8'd32,8'd160} : s = 192;
	{8'd32,8'd161} : s = 193;
	{8'd32,8'd162} : s = 194;
	{8'd32,8'd163} : s = 195;
	{8'd32,8'd164} : s = 196;
	{8'd32,8'd165} : s = 197;
	{8'd32,8'd166} : s = 198;
	{8'd32,8'd167} : s = 199;
	{8'd32,8'd168} : s = 200;
	{8'd32,8'd169} : s = 201;
	{8'd32,8'd170} : s = 202;
	{8'd32,8'd171} : s = 203;
	{8'd32,8'd172} : s = 204;
	{8'd32,8'd173} : s = 205;
	{8'd32,8'd174} : s = 206;
	{8'd32,8'd175} : s = 207;
	{8'd32,8'd176} : s = 208;
	{8'd32,8'd177} : s = 209;
	{8'd32,8'd178} : s = 210;
	{8'd32,8'd179} : s = 211;
	{8'd32,8'd180} : s = 212;
	{8'd32,8'd181} : s = 213;
	{8'd32,8'd182} : s = 214;
	{8'd32,8'd183} : s = 215;
	{8'd32,8'd184} : s = 216;
	{8'd32,8'd185} : s = 217;
	{8'd32,8'd186} : s = 218;
	{8'd32,8'd187} : s = 219;
	{8'd32,8'd188} : s = 220;
	{8'd32,8'd189} : s = 221;
	{8'd32,8'd190} : s = 222;
	{8'd32,8'd191} : s = 223;
	{8'd32,8'd192} : s = 224;
	{8'd32,8'd193} : s = 225;
	{8'd32,8'd194} : s = 226;
	{8'd32,8'd195} : s = 227;
	{8'd32,8'd196} : s = 228;
	{8'd32,8'd197} : s = 229;
	{8'd32,8'd198} : s = 230;
	{8'd32,8'd199} : s = 231;
	{8'd32,8'd200} : s = 232;
	{8'd32,8'd201} : s = 233;
	{8'd32,8'd202} : s = 234;
	{8'd32,8'd203} : s = 235;
	{8'd32,8'd204} : s = 236;
	{8'd32,8'd205} : s = 237;
	{8'd32,8'd206} : s = 238;
	{8'd32,8'd207} : s = 239;
	{8'd32,8'd208} : s = 240;
	{8'd32,8'd209} : s = 241;
	{8'd32,8'd210} : s = 242;
	{8'd32,8'd211} : s = 243;
	{8'd32,8'd212} : s = 244;
	{8'd32,8'd213} : s = 245;
	{8'd32,8'd214} : s = 246;
	{8'd32,8'd215} : s = 247;
	{8'd32,8'd216} : s = 248;
	{8'd32,8'd217} : s = 249;
	{8'd32,8'd218} : s = 250;
	{8'd32,8'd219} : s = 251;
	{8'd32,8'd220} : s = 252;
	{8'd32,8'd221} : s = 253;
	{8'd32,8'd222} : s = 254;
	{8'd32,8'd223} : s = 255;
	{8'd32,8'd224} : s = 256;
	{8'd32,8'd225} : s = 257;
	{8'd32,8'd226} : s = 258;
	{8'd32,8'd227} : s = 259;
	{8'd32,8'd228} : s = 260;
	{8'd32,8'd229} : s = 261;
	{8'd32,8'd230} : s = 262;
	{8'd32,8'd231} : s = 263;
	{8'd32,8'd232} : s = 264;
	{8'd32,8'd233} : s = 265;
	{8'd32,8'd234} : s = 266;
	{8'd32,8'd235} : s = 267;
	{8'd32,8'd236} : s = 268;
	{8'd32,8'd237} : s = 269;
	{8'd32,8'd238} : s = 270;
	{8'd32,8'd239} : s = 271;
	{8'd32,8'd240} : s = 272;
	{8'd32,8'd241} : s = 273;
	{8'd32,8'd242} : s = 274;
	{8'd32,8'd243} : s = 275;
	{8'd32,8'd244} : s = 276;
	{8'd32,8'd245} : s = 277;
	{8'd32,8'd246} : s = 278;
	{8'd32,8'd247} : s = 279;
	{8'd32,8'd248} : s = 280;
	{8'd32,8'd249} : s = 281;
	{8'd32,8'd250} : s = 282;
	{8'd32,8'd251} : s = 283;
	{8'd32,8'd252} : s = 284;
	{8'd32,8'd253} : s = 285;
	{8'd32,8'd254} : s = 286;
	{8'd32,8'd255} : s = 287;
	{8'd33,8'd0} : s = 33;
	{8'd33,8'd1} : s = 34;
	{8'd33,8'd2} : s = 35;
	{8'd33,8'd3} : s = 36;
	{8'd33,8'd4} : s = 37;
	{8'd33,8'd5} : s = 38;
	{8'd33,8'd6} : s = 39;
	{8'd33,8'd7} : s = 40;
	{8'd33,8'd8} : s = 41;
	{8'd33,8'd9} : s = 42;
	{8'd33,8'd10} : s = 43;
	{8'd33,8'd11} : s = 44;
	{8'd33,8'd12} : s = 45;
	{8'd33,8'd13} : s = 46;
	{8'd33,8'd14} : s = 47;
	{8'd33,8'd15} : s = 48;
	{8'd33,8'd16} : s = 49;
	{8'd33,8'd17} : s = 50;
	{8'd33,8'd18} : s = 51;
	{8'd33,8'd19} : s = 52;
	{8'd33,8'd20} : s = 53;
	{8'd33,8'd21} : s = 54;
	{8'd33,8'd22} : s = 55;
	{8'd33,8'd23} : s = 56;
	{8'd33,8'd24} : s = 57;
	{8'd33,8'd25} : s = 58;
	{8'd33,8'd26} : s = 59;
	{8'd33,8'd27} : s = 60;
	{8'd33,8'd28} : s = 61;
	{8'd33,8'd29} : s = 62;
	{8'd33,8'd30} : s = 63;
	{8'd33,8'd31} : s = 64;
	{8'd33,8'd32} : s = 65;
	{8'd33,8'd33} : s = 66;
	{8'd33,8'd34} : s = 67;
	{8'd33,8'd35} : s = 68;
	{8'd33,8'd36} : s = 69;
	{8'd33,8'd37} : s = 70;
	{8'd33,8'd38} : s = 71;
	{8'd33,8'd39} : s = 72;
	{8'd33,8'd40} : s = 73;
	{8'd33,8'd41} : s = 74;
	{8'd33,8'd42} : s = 75;
	{8'd33,8'd43} : s = 76;
	{8'd33,8'd44} : s = 77;
	{8'd33,8'd45} : s = 78;
	{8'd33,8'd46} : s = 79;
	{8'd33,8'd47} : s = 80;
	{8'd33,8'd48} : s = 81;
	{8'd33,8'd49} : s = 82;
	{8'd33,8'd50} : s = 83;
	{8'd33,8'd51} : s = 84;
	{8'd33,8'd52} : s = 85;
	{8'd33,8'd53} : s = 86;
	{8'd33,8'd54} : s = 87;
	{8'd33,8'd55} : s = 88;
	{8'd33,8'd56} : s = 89;
	{8'd33,8'd57} : s = 90;
	{8'd33,8'd58} : s = 91;
	{8'd33,8'd59} : s = 92;
	{8'd33,8'd60} : s = 93;
	{8'd33,8'd61} : s = 94;
	{8'd33,8'd62} : s = 95;
	{8'd33,8'd63} : s = 96;
	{8'd33,8'd64} : s = 97;
	{8'd33,8'd65} : s = 98;
	{8'd33,8'd66} : s = 99;
	{8'd33,8'd67} : s = 100;
	{8'd33,8'd68} : s = 101;
	{8'd33,8'd69} : s = 102;
	{8'd33,8'd70} : s = 103;
	{8'd33,8'd71} : s = 104;
	{8'd33,8'd72} : s = 105;
	{8'd33,8'd73} : s = 106;
	{8'd33,8'd74} : s = 107;
	{8'd33,8'd75} : s = 108;
	{8'd33,8'd76} : s = 109;
	{8'd33,8'd77} : s = 110;
	{8'd33,8'd78} : s = 111;
	{8'd33,8'd79} : s = 112;
	{8'd33,8'd80} : s = 113;
	{8'd33,8'd81} : s = 114;
	{8'd33,8'd82} : s = 115;
	{8'd33,8'd83} : s = 116;
	{8'd33,8'd84} : s = 117;
	{8'd33,8'd85} : s = 118;
	{8'd33,8'd86} : s = 119;
	{8'd33,8'd87} : s = 120;
	{8'd33,8'd88} : s = 121;
	{8'd33,8'd89} : s = 122;
	{8'd33,8'd90} : s = 123;
	{8'd33,8'd91} : s = 124;
	{8'd33,8'd92} : s = 125;
	{8'd33,8'd93} : s = 126;
	{8'd33,8'd94} : s = 127;
	{8'd33,8'd95} : s = 128;
	{8'd33,8'd96} : s = 129;
	{8'd33,8'd97} : s = 130;
	{8'd33,8'd98} : s = 131;
	{8'd33,8'd99} : s = 132;
	{8'd33,8'd100} : s = 133;
	{8'd33,8'd101} : s = 134;
	{8'd33,8'd102} : s = 135;
	{8'd33,8'd103} : s = 136;
	{8'd33,8'd104} : s = 137;
	{8'd33,8'd105} : s = 138;
	{8'd33,8'd106} : s = 139;
	{8'd33,8'd107} : s = 140;
	{8'd33,8'd108} : s = 141;
	{8'd33,8'd109} : s = 142;
	{8'd33,8'd110} : s = 143;
	{8'd33,8'd111} : s = 144;
	{8'd33,8'd112} : s = 145;
	{8'd33,8'd113} : s = 146;
	{8'd33,8'd114} : s = 147;
	{8'd33,8'd115} : s = 148;
	{8'd33,8'd116} : s = 149;
	{8'd33,8'd117} : s = 150;
	{8'd33,8'd118} : s = 151;
	{8'd33,8'd119} : s = 152;
	{8'd33,8'd120} : s = 153;
	{8'd33,8'd121} : s = 154;
	{8'd33,8'd122} : s = 155;
	{8'd33,8'd123} : s = 156;
	{8'd33,8'd124} : s = 157;
	{8'd33,8'd125} : s = 158;
	{8'd33,8'd126} : s = 159;
	{8'd33,8'd127} : s = 160;
	{8'd33,8'd128} : s = 161;
	{8'd33,8'd129} : s = 162;
	{8'd33,8'd130} : s = 163;
	{8'd33,8'd131} : s = 164;
	{8'd33,8'd132} : s = 165;
	{8'd33,8'd133} : s = 166;
	{8'd33,8'd134} : s = 167;
	{8'd33,8'd135} : s = 168;
	{8'd33,8'd136} : s = 169;
	{8'd33,8'd137} : s = 170;
	{8'd33,8'd138} : s = 171;
	{8'd33,8'd139} : s = 172;
	{8'd33,8'd140} : s = 173;
	{8'd33,8'd141} : s = 174;
	{8'd33,8'd142} : s = 175;
	{8'd33,8'd143} : s = 176;
	{8'd33,8'd144} : s = 177;
	{8'd33,8'd145} : s = 178;
	{8'd33,8'd146} : s = 179;
	{8'd33,8'd147} : s = 180;
	{8'd33,8'd148} : s = 181;
	{8'd33,8'd149} : s = 182;
	{8'd33,8'd150} : s = 183;
	{8'd33,8'd151} : s = 184;
	{8'd33,8'd152} : s = 185;
	{8'd33,8'd153} : s = 186;
	{8'd33,8'd154} : s = 187;
	{8'd33,8'd155} : s = 188;
	{8'd33,8'd156} : s = 189;
	{8'd33,8'd157} : s = 190;
	{8'd33,8'd158} : s = 191;
	{8'd33,8'd159} : s = 192;
	{8'd33,8'd160} : s = 193;
	{8'd33,8'd161} : s = 194;
	{8'd33,8'd162} : s = 195;
	{8'd33,8'd163} : s = 196;
	{8'd33,8'd164} : s = 197;
	{8'd33,8'd165} : s = 198;
	{8'd33,8'd166} : s = 199;
	{8'd33,8'd167} : s = 200;
	{8'd33,8'd168} : s = 201;
	{8'd33,8'd169} : s = 202;
	{8'd33,8'd170} : s = 203;
	{8'd33,8'd171} : s = 204;
	{8'd33,8'd172} : s = 205;
	{8'd33,8'd173} : s = 206;
	{8'd33,8'd174} : s = 207;
	{8'd33,8'd175} : s = 208;
	{8'd33,8'd176} : s = 209;
	{8'd33,8'd177} : s = 210;
	{8'd33,8'd178} : s = 211;
	{8'd33,8'd179} : s = 212;
	{8'd33,8'd180} : s = 213;
	{8'd33,8'd181} : s = 214;
	{8'd33,8'd182} : s = 215;
	{8'd33,8'd183} : s = 216;
	{8'd33,8'd184} : s = 217;
	{8'd33,8'd185} : s = 218;
	{8'd33,8'd186} : s = 219;
	{8'd33,8'd187} : s = 220;
	{8'd33,8'd188} : s = 221;
	{8'd33,8'd189} : s = 222;
	{8'd33,8'd190} : s = 223;
	{8'd33,8'd191} : s = 224;
	{8'd33,8'd192} : s = 225;
	{8'd33,8'd193} : s = 226;
	{8'd33,8'd194} : s = 227;
	{8'd33,8'd195} : s = 228;
	{8'd33,8'd196} : s = 229;
	{8'd33,8'd197} : s = 230;
	{8'd33,8'd198} : s = 231;
	{8'd33,8'd199} : s = 232;
	{8'd33,8'd200} : s = 233;
	{8'd33,8'd201} : s = 234;
	{8'd33,8'd202} : s = 235;
	{8'd33,8'd203} : s = 236;
	{8'd33,8'd204} : s = 237;
	{8'd33,8'd205} : s = 238;
	{8'd33,8'd206} : s = 239;
	{8'd33,8'd207} : s = 240;
	{8'd33,8'd208} : s = 241;
	{8'd33,8'd209} : s = 242;
	{8'd33,8'd210} : s = 243;
	{8'd33,8'd211} : s = 244;
	{8'd33,8'd212} : s = 245;
	{8'd33,8'd213} : s = 246;
	{8'd33,8'd214} : s = 247;
	{8'd33,8'd215} : s = 248;
	{8'd33,8'd216} : s = 249;
	{8'd33,8'd217} : s = 250;
	{8'd33,8'd218} : s = 251;
	{8'd33,8'd219} : s = 252;
	{8'd33,8'd220} : s = 253;
	{8'd33,8'd221} : s = 254;
	{8'd33,8'd222} : s = 255;
	{8'd33,8'd223} : s = 256;
	{8'd33,8'd224} : s = 257;
	{8'd33,8'd225} : s = 258;
	{8'd33,8'd226} : s = 259;
	{8'd33,8'd227} : s = 260;
	{8'd33,8'd228} : s = 261;
	{8'd33,8'd229} : s = 262;
	{8'd33,8'd230} : s = 263;
	{8'd33,8'd231} : s = 264;
	{8'd33,8'd232} : s = 265;
	{8'd33,8'd233} : s = 266;
	{8'd33,8'd234} : s = 267;
	{8'd33,8'd235} : s = 268;
	{8'd33,8'd236} : s = 269;
	{8'd33,8'd237} : s = 270;
	{8'd33,8'd238} : s = 271;
	{8'd33,8'd239} : s = 272;
	{8'd33,8'd240} : s = 273;
	{8'd33,8'd241} : s = 274;
	{8'd33,8'd242} : s = 275;
	{8'd33,8'd243} : s = 276;
	{8'd33,8'd244} : s = 277;
	{8'd33,8'd245} : s = 278;
	{8'd33,8'd246} : s = 279;
	{8'd33,8'd247} : s = 280;
	{8'd33,8'd248} : s = 281;
	{8'd33,8'd249} : s = 282;
	{8'd33,8'd250} : s = 283;
	{8'd33,8'd251} : s = 284;
	{8'd33,8'd252} : s = 285;
	{8'd33,8'd253} : s = 286;
	{8'd33,8'd254} : s = 287;
	{8'd33,8'd255} : s = 288;
	{8'd34,8'd0} : s = 34;
	{8'd34,8'd1} : s = 35;
	{8'd34,8'd2} : s = 36;
	{8'd34,8'd3} : s = 37;
	{8'd34,8'd4} : s = 38;
	{8'd34,8'd5} : s = 39;
	{8'd34,8'd6} : s = 40;
	{8'd34,8'd7} : s = 41;
	{8'd34,8'd8} : s = 42;
	{8'd34,8'd9} : s = 43;
	{8'd34,8'd10} : s = 44;
	{8'd34,8'd11} : s = 45;
	{8'd34,8'd12} : s = 46;
	{8'd34,8'd13} : s = 47;
	{8'd34,8'd14} : s = 48;
	{8'd34,8'd15} : s = 49;
	{8'd34,8'd16} : s = 50;
	{8'd34,8'd17} : s = 51;
	{8'd34,8'd18} : s = 52;
	{8'd34,8'd19} : s = 53;
	{8'd34,8'd20} : s = 54;
	{8'd34,8'd21} : s = 55;
	{8'd34,8'd22} : s = 56;
	{8'd34,8'd23} : s = 57;
	{8'd34,8'd24} : s = 58;
	{8'd34,8'd25} : s = 59;
	{8'd34,8'd26} : s = 60;
	{8'd34,8'd27} : s = 61;
	{8'd34,8'd28} : s = 62;
	{8'd34,8'd29} : s = 63;
	{8'd34,8'd30} : s = 64;
	{8'd34,8'd31} : s = 65;
	{8'd34,8'd32} : s = 66;
	{8'd34,8'd33} : s = 67;
	{8'd34,8'd34} : s = 68;
	{8'd34,8'd35} : s = 69;
	{8'd34,8'd36} : s = 70;
	{8'd34,8'd37} : s = 71;
	{8'd34,8'd38} : s = 72;
	{8'd34,8'd39} : s = 73;
	{8'd34,8'd40} : s = 74;
	{8'd34,8'd41} : s = 75;
	{8'd34,8'd42} : s = 76;
	{8'd34,8'd43} : s = 77;
	{8'd34,8'd44} : s = 78;
	{8'd34,8'd45} : s = 79;
	{8'd34,8'd46} : s = 80;
	{8'd34,8'd47} : s = 81;
	{8'd34,8'd48} : s = 82;
	{8'd34,8'd49} : s = 83;
	{8'd34,8'd50} : s = 84;
	{8'd34,8'd51} : s = 85;
	{8'd34,8'd52} : s = 86;
	{8'd34,8'd53} : s = 87;
	{8'd34,8'd54} : s = 88;
	{8'd34,8'd55} : s = 89;
	{8'd34,8'd56} : s = 90;
	{8'd34,8'd57} : s = 91;
	{8'd34,8'd58} : s = 92;
	{8'd34,8'd59} : s = 93;
	{8'd34,8'd60} : s = 94;
	{8'd34,8'd61} : s = 95;
	{8'd34,8'd62} : s = 96;
	{8'd34,8'd63} : s = 97;
	{8'd34,8'd64} : s = 98;
	{8'd34,8'd65} : s = 99;
	{8'd34,8'd66} : s = 100;
	{8'd34,8'd67} : s = 101;
	{8'd34,8'd68} : s = 102;
	{8'd34,8'd69} : s = 103;
	{8'd34,8'd70} : s = 104;
	{8'd34,8'd71} : s = 105;
	{8'd34,8'd72} : s = 106;
	{8'd34,8'd73} : s = 107;
	{8'd34,8'd74} : s = 108;
	{8'd34,8'd75} : s = 109;
	{8'd34,8'd76} : s = 110;
	{8'd34,8'd77} : s = 111;
	{8'd34,8'd78} : s = 112;
	{8'd34,8'd79} : s = 113;
	{8'd34,8'd80} : s = 114;
	{8'd34,8'd81} : s = 115;
	{8'd34,8'd82} : s = 116;
	{8'd34,8'd83} : s = 117;
	{8'd34,8'd84} : s = 118;
	{8'd34,8'd85} : s = 119;
	{8'd34,8'd86} : s = 120;
	{8'd34,8'd87} : s = 121;
	{8'd34,8'd88} : s = 122;
	{8'd34,8'd89} : s = 123;
	{8'd34,8'd90} : s = 124;
	{8'd34,8'd91} : s = 125;
	{8'd34,8'd92} : s = 126;
	{8'd34,8'd93} : s = 127;
	{8'd34,8'd94} : s = 128;
	{8'd34,8'd95} : s = 129;
	{8'd34,8'd96} : s = 130;
	{8'd34,8'd97} : s = 131;
	{8'd34,8'd98} : s = 132;
	{8'd34,8'd99} : s = 133;
	{8'd34,8'd100} : s = 134;
	{8'd34,8'd101} : s = 135;
	{8'd34,8'd102} : s = 136;
	{8'd34,8'd103} : s = 137;
	{8'd34,8'd104} : s = 138;
	{8'd34,8'd105} : s = 139;
	{8'd34,8'd106} : s = 140;
	{8'd34,8'd107} : s = 141;
	{8'd34,8'd108} : s = 142;
	{8'd34,8'd109} : s = 143;
	{8'd34,8'd110} : s = 144;
	{8'd34,8'd111} : s = 145;
	{8'd34,8'd112} : s = 146;
	{8'd34,8'd113} : s = 147;
	{8'd34,8'd114} : s = 148;
	{8'd34,8'd115} : s = 149;
	{8'd34,8'd116} : s = 150;
	{8'd34,8'd117} : s = 151;
	{8'd34,8'd118} : s = 152;
	{8'd34,8'd119} : s = 153;
	{8'd34,8'd120} : s = 154;
	{8'd34,8'd121} : s = 155;
	{8'd34,8'd122} : s = 156;
	{8'd34,8'd123} : s = 157;
	{8'd34,8'd124} : s = 158;
	{8'd34,8'd125} : s = 159;
	{8'd34,8'd126} : s = 160;
	{8'd34,8'd127} : s = 161;
	{8'd34,8'd128} : s = 162;
	{8'd34,8'd129} : s = 163;
	{8'd34,8'd130} : s = 164;
	{8'd34,8'd131} : s = 165;
	{8'd34,8'd132} : s = 166;
	{8'd34,8'd133} : s = 167;
	{8'd34,8'd134} : s = 168;
	{8'd34,8'd135} : s = 169;
	{8'd34,8'd136} : s = 170;
	{8'd34,8'd137} : s = 171;
	{8'd34,8'd138} : s = 172;
	{8'd34,8'd139} : s = 173;
	{8'd34,8'd140} : s = 174;
	{8'd34,8'd141} : s = 175;
	{8'd34,8'd142} : s = 176;
	{8'd34,8'd143} : s = 177;
	{8'd34,8'd144} : s = 178;
	{8'd34,8'd145} : s = 179;
	{8'd34,8'd146} : s = 180;
	{8'd34,8'd147} : s = 181;
	{8'd34,8'd148} : s = 182;
	{8'd34,8'd149} : s = 183;
	{8'd34,8'd150} : s = 184;
	{8'd34,8'd151} : s = 185;
	{8'd34,8'd152} : s = 186;
	{8'd34,8'd153} : s = 187;
	{8'd34,8'd154} : s = 188;
	{8'd34,8'd155} : s = 189;
	{8'd34,8'd156} : s = 190;
	{8'd34,8'd157} : s = 191;
	{8'd34,8'd158} : s = 192;
	{8'd34,8'd159} : s = 193;
	{8'd34,8'd160} : s = 194;
	{8'd34,8'd161} : s = 195;
	{8'd34,8'd162} : s = 196;
	{8'd34,8'd163} : s = 197;
	{8'd34,8'd164} : s = 198;
	{8'd34,8'd165} : s = 199;
	{8'd34,8'd166} : s = 200;
	{8'd34,8'd167} : s = 201;
	{8'd34,8'd168} : s = 202;
	{8'd34,8'd169} : s = 203;
	{8'd34,8'd170} : s = 204;
	{8'd34,8'd171} : s = 205;
	{8'd34,8'd172} : s = 206;
	{8'd34,8'd173} : s = 207;
	{8'd34,8'd174} : s = 208;
	{8'd34,8'd175} : s = 209;
	{8'd34,8'd176} : s = 210;
	{8'd34,8'd177} : s = 211;
	{8'd34,8'd178} : s = 212;
	{8'd34,8'd179} : s = 213;
	{8'd34,8'd180} : s = 214;
	{8'd34,8'd181} : s = 215;
	{8'd34,8'd182} : s = 216;
	{8'd34,8'd183} : s = 217;
	{8'd34,8'd184} : s = 218;
	{8'd34,8'd185} : s = 219;
	{8'd34,8'd186} : s = 220;
	{8'd34,8'd187} : s = 221;
	{8'd34,8'd188} : s = 222;
	{8'd34,8'd189} : s = 223;
	{8'd34,8'd190} : s = 224;
	{8'd34,8'd191} : s = 225;
	{8'd34,8'd192} : s = 226;
	{8'd34,8'd193} : s = 227;
	{8'd34,8'd194} : s = 228;
	{8'd34,8'd195} : s = 229;
	{8'd34,8'd196} : s = 230;
	{8'd34,8'd197} : s = 231;
	{8'd34,8'd198} : s = 232;
	{8'd34,8'd199} : s = 233;
	{8'd34,8'd200} : s = 234;
	{8'd34,8'd201} : s = 235;
	{8'd34,8'd202} : s = 236;
	{8'd34,8'd203} : s = 237;
	{8'd34,8'd204} : s = 238;
	{8'd34,8'd205} : s = 239;
	{8'd34,8'd206} : s = 240;
	{8'd34,8'd207} : s = 241;
	{8'd34,8'd208} : s = 242;
	{8'd34,8'd209} : s = 243;
	{8'd34,8'd210} : s = 244;
	{8'd34,8'd211} : s = 245;
	{8'd34,8'd212} : s = 246;
	{8'd34,8'd213} : s = 247;
	{8'd34,8'd214} : s = 248;
	{8'd34,8'd215} : s = 249;
	{8'd34,8'd216} : s = 250;
	{8'd34,8'd217} : s = 251;
	{8'd34,8'd218} : s = 252;
	{8'd34,8'd219} : s = 253;
	{8'd34,8'd220} : s = 254;
	{8'd34,8'd221} : s = 255;
	{8'd34,8'd222} : s = 256;
	{8'd34,8'd223} : s = 257;
	{8'd34,8'd224} : s = 258;
	{8'd34,8'd225} : s = 259;
	{8'd34,8'd226} : s = 260;
	{8'd34,8'd227} : s = 261;
	{8'd34,8'd228} : s = 262;
	{8'd34,8'd229} : s = 263;
	{8'd34,8'd230} : s = 264;
	{8'd34,8'd231} : s = 265;
	{8'd34,8'd232} : s = 266;
	{8'd34,8'd233} : s = 267;
	{8'd34,8'd234} : s = 268;
	{8'd34,8'd235} : s = 269;
	{8'd34,8'd236} : s = 270;
	{8'd34,8'd237} : s = 271;
	{8'd34,8'd238} : s = 272;
	{8'd34,8'd239} : s = 273;
	{8'd34,8'd240} : s = 274;
	{8'd34,8'd241} : s = 275;
	{8'd34,8'd242} : s = 276;
	{8'd34,8'd243} : s = 277;
	{8'd34,8'd244} : s = 278;
	{8'd34,8'd245} : s = 279;
	{8'd34,8'd246} : s = 280;
	{8'd34,8'd247} : s = 281;
	{8'd34,8'd248} : s = 282;
	{8'd34,8'd249} : s = 283;
	{8'd34,8'd250} : s = 284;
	{8'd34,8'd251} : s = 285;
	{8'd34,8'd252} : s = 286;
	{8'd34,8'd253} : s = 287;
	{8'd34,8'd254} : s = 288;
	{8'd34,8'd255} : s = 289;
	{8'd35,8'd0} : s = 35;
	{8'd35,8'd1} : s = 36;
	{8'd35,8'd2} : s = 37;
	{8'd35,8'd3} : s = 38;
	{8'd35,8'd4} : s = 39;
	{8'd35,8'd5} : s = 40;
	{8'd35,8'd6} : s = 41;
	{8'd35,8'd7} : s = 42;
	{8'd35,8'd8} : s = 43;
	{8'd35,8'd9} : s = 44;
	{8'd35,8'd10} : s = 45;
	{8'd35,8'd11} : s = 46;
	{8'd35,8'd12} : s = 47;
	{8'd35,8'd13} : s = 48;
	{8'd35,8'd14} : s = 49;
	{8'd35,8'd15} : s = 50;
	{8'd35,8'd16} : s = 51;
	{8'd35,8'd17} : s = 52;
	{8'd35,8'd18} : s = 53;
	{8'd35,8'd19} : s = 54;
	{8'd35,8'd20} : s = 55;
	{8'd35,8'd21} : s = 56;
	{8'd35,8'd22} : s = 57;
	{8'd35,8'd23} : s = 58;
	{8'd35,8'd24} : s = 59;
	{8'd35,8'd25} : s = 60;
	{8'd35,8'd26} : s = 61;
	{8'd35,8'd27} : s = 62;
	{8'd35,8'd28} : s = 63;
	{8'd35,8'd29} : s = 64;
	{8'd35,8'd30} : s = 65;
	{8'd35,8'd31} : s = 66;
	{8'd35,8'd32} : s = 67;
	{8'd35,8'd33} : s = 68;
	{8'd35,8'd34} : s = 69;
	{8'd35,8'd35} : s = 70;
	{8'd35,8'd36} : s = 71;
	{8'd35,8'd37} : s = 72;
	{8'd35,8'd38} : s = 73;
	{8'd35,8'd39} : s = 74;
	{8'd35,8'd40} : s = 75;
	{8'd35,8'd41} : s = 76;
	{8'd35,8'd42} : s = 77;
	{8'd35,8'd43} : s = 78;
	{8'd35,8'd44} : s = 79;
	{8'd35,8'd45} : s = 80;
	{8'd35,8'd46} : s = 81;
	{8'd35,8'd47} : s = 82;
	{8'd35,8'd48} : s = 83;
	{8'd35,8'd49} : s = 84;
	{8'd35,8'd50} : s = 85;
	{8'd35,8'd51} : s = 86;
	{8'd35,8'd52} : s = 87;
	{8'd35,8'd53} : s = 88;
	{8'd35,8'd54} : s = 89;
	{8'd35,8'd55} : s = 90;
	{8'd35,8'd56} : s = 91;
	{8'd35,8'd57} : s = 92;
	{8'd35,8'd58} : s = 93;
	{8'd35,8'd59} : s = 94;
	{8'd35,8'd60} : s = 95;
	{8'd35,8'd61} : s = 96;
	{8'd35,8'd62} : s = 97;
	{8'd35,8'd63} : s = 98;
	{8'd35,8'd64} : s = 99;
	{8'd35,8'd65} : s = 100;
	{8'd35,8'd66} : s = 101;
	{8'd35,8'd67} : s = 102;
	{8'd35,8'd68} : s = 103;
	{8'd35,8'd69} : s = 104;
	{8'd35,8'd70} : s = 105;
	{8'd35,8'd71} : s = 106;
	{8'd35,8'd72} : s = 107;
	{8'd35,8'd73} : s = 108;
	{8'd35,8'd74} : s = 109;
	{8'd35,8'd75} : s = 110;
	{8'd35,8'd76} : s = 111;
	{8'd35,8'd77} : s = 112;
	{8'd35,8'd78} : s = 113;
	{8'd35,8'd79} : s = 114;
	{8'd35,8'd80} : s = 115;
	{8'd35,8'd81} : s = 116;
	{8'd35,8'd82} : s = 117;
	{8'd35,8'd83} : s = 118;
	{8'd35,8'd84} : s = 119;
	{8'd35,8'd85} : s = 120;
	{8'd35,8'd86} : s = 121;
	{8'd35,8'd87} : s = 122;
	{8'd35,8'd88} : s = 123;
	{8'd35,8'd89} : s = 124;
	{8'd35,8'd90} : s = 125;
	{8'd35,8'd91} : s = 126;
	{8'd35,8'd92} : s = 127;
	{8'd35,8'd93} : s = 128;
	{8'd35,8'd94} : s = 129;
	{8'd35,8'd95} : s = 130;
	{8'd35,8'd96} : s = 131;
	{8'd35,8'd97} : s = 132;
	{8'd35,8'd98} : s = 133;
	{8'd35,8'd99} : s = 134;
	{8'd35,8'd100} : s = 135;
	{8'd35,8'd101} : s = 136;
	{8'd35,8'd102} : s = 137;
	{8'd35,8'd103} : s = 138;
	{8'd35,8'd104} : s = 139;
	{8'd35,8'd105} : s = 140;
	{8'd35,8'd106} : s = 141;
	{8'd35,8'd107} : s = 142;
	{8'd35,8'd108} : s = 143;
	{8'd35,8'd109} : s = 144;
	{8'd35,8'd110} : s = 145;
	{8'd35,8'd111} : s = 146;
	{8'd35,8'd112} : s = 147;
	{8'd35,8'd113} : s = 148;
	{8'd35,8'd114} : s = 149;
	{8'd35,8'd115} : s = 150;
	{8'd35,8'd116} : s = 151;
	{8'd35,8'd117} : s = 152;
	{8'd35,8'd118} : s = 153;
	{8'd35,8'd119} : s = 154;
	{8'd35,8'd120} : s = 155;
	{8'd35,8'd121} : s = 156;
	{8'd35,8'd122} : s = 157;
	{8'd35,8'd123} : s = 158;
	{8'd35,8'd124} : s = 159;
	{8'd35,8'd125} : s = 160;
	{8'd35,8'd126} : s = 161;
	{8'd35,8'd127} : s = 162;
	{8'd35,8'd128} : s = 163;
	{8'd35,8'd129} : s = 164;
	{8'd35,8'd130} : s = 165;
	{8'd35,8'd131} : s = 166;
	{8'd35,8'd132} : s = 167;
	{8'd35,8'd133} : s = 168;
	{8'd35,8'd134} : s = 169;
	{8'd35,8'd135} : s = 170;
	{8'd35,8'd136} : s = 171;
	{8'd35,8'd137} : s = 172;
	{8'd35,8'd138} : s = 173;
	{8'd35,8'd139} : s = 174;
	{8'd35,8'd140} : s = 175;
	{8'd35,8'd141} : s = 176;
	{8'd35,8'd142} : s = 177;
	{8'd35,8'd143} : s = 178;
	{8'd35,8'd144} : s = 179;
	{8'd35,8'd145} : s = 180;
	{8'd35,8'd146} : s = 181;
	{8'd35,8'd147} : s = 182;
	{8'd35,8'd148} : s = 183;
	{8'd35,8'd149} : s = 184;
	{8'd35,8'd150} : s = 185;
	{8'd35,8'd151} : s = 186;
	{8'd35,8'd152} : s = 187;
	{8'd35,8'd153} : s = 188;
	{8'd35,8'd154} : s = 189;
	{8'd35,8'd155} : s = 190;
	{8'd35,8'd156} : s = 191;
	{8'd35,8'd157} : s = 192;
	{8'd35,8'd158} : s = 193;
	{8'd35,8'd159} : s = 194;
	{8'd35,8'd160} : s = 195;
	{8'd35,8'd161} : s = 196;
	{8'd35,8'd162} : s = 197;
	{8'd35,8'd163} : s = 198;
	{8'd35,8'd164} : s = 199;
	{8'd35,8'd165} : s = 200;
	{8'd35,8'd166} : s = 201;
	{8'd35,8'd167} : s = 202;
	{8'd35,8'd168} : s = 203;
	{8'd35,8'd169} : s = 204;
	{8'd35,8'd170} : s = 205;
	{8'd35,8'd171} : s = 206;
	{8'd35,8'd172} : s = 207;
	{8'd35,8'd173} : s = 208;
	{8'd35,8'd174} : s = 209;
	{8'd35,8'd175} : s = 210;
	{8'd35,8'd176} : s = 211;
	{8'd35,8'd177} : s = 212;
	{8'd35,8'd178} : s = 213;
	{8'd35,8'd179} : s = 214;
	{8'd35,8'd180} : s = 215;
	{8'd35,8'd181} : s = 216;
	{8'd35,8'd182} : s = 217;
	{8'd35,8'd183} : s = 218;
	{8'd35,8'd184} : s = 219;
	{8'd35,8'd185} : s = 220;
	{8'd35,8'd186} : s = 221;
	{8'd35,8'd187} : s = 222;
	{8'd35,8'd188} : s = 223;
	{8'd35,8'd189} : s = 224;
	{8'd35,8'd190} : s = 225;
	{8'd35,8'd191} : s = 226;
	{8'd35,8'd192} : s = 227;
	{8'd35,8'd193} : s = 228;
	{8'd35,8'd194} : s = 229;
	{8'd35,8'd195} : s = 230;
	{8'd35,8'd196} : s = 231;
	{8'd35,8'd197} : s = 232;
	{8'd35,8'd198} : s = 233;
	{8'd35,8'd199} : s = 234;
	{8'd35,8'd200} : s = 235;
	{8'd35,8'd201} : s = 236;
	{8'd35,8'd202} : s = 237;
	{8'd35,8'd203} : s = 238;
	{8'd35,8'd204} : s = 239;
	{8'd35,8'd205} : s = 240;
	{8'd35,8'd206} : s = 241;
	{8'd35,8'd207} : s = 242;
	{8'd35,8'd208} : s = 243;
	{8'd35,8'd209} : s = 244;
	{8'd35,8'd210} : s = 245;
	{8'd35,8'd211} : s = 246;
	{8'd35,8'd212} : s = 247;
	{8'd35,8'd213} : s = 248;
	{8'd35,8'd214} : s = 249;
	{8'd35,8'd215} : s = 250;
	{8'd35,8'd216} : s = 251;
	{8'd35,8'd217} : s = 252;
	{8'd35,8'd218} : s = 253;
	{8'd35,8'd219} : s = 254;
	{8'd35,8'd220} : s = 255;
	{8'd35,8'd221} : s = 256;
	{8'd35,8'd222} : s = 257;
	{8'd35,8'd223} : s = 258;
	{8'd35,8'd224} : s = 259;
	{8'd35,8'd225} : s = 260;
	{8'd35,8'd226} : s = 261;
	{8'd35,8'd227} : s = 262;
	{8'd35,8'd228} : s = 263;
	{8'd35,8'd229} : s = 264;
	{8'd35,8'd230} : s = 265;
	{8'd35,8'd231} : s = 266;
	{8'd35,8'd232} : s = 267;
	{8'd35,8'd233} : s = 268;
	{8'd35,8'd234} : s = 269;
	{8'd35,8'd235} : s = 270;
	{8'd35,8'd236} : s = 271;
	{8'd35,8'd237} : s = 272;
	{8'd35,8'd238} : s = 273;
	{8'd35,8'd239} : s = 274;
	{8'd35,8'd240} : s = 275;
	{8'd35,8'd241} : s = 276;
	{8'd35,8'd242} : s = 277;
	{8'd35,8'd243} : s = 278;
	{8'd35,8'd244} : s = 279;
	{8'd35,8'd245} : s = 280;
	{8'd35,8'd246} : s = 281;
	{8'd35,8'd247} : s = 282;
	{8'd35,8'd248} : s = 283;
	{8'd35,8'd249} : s = 284;
	{8'd35,8'd250} : s = 285;
	{8'd35,8'd251} : s = 286;
	{8'd35,8'd252} : s = 287;
	{8'd35,8'd253} : s = 288;
	{8'd35,8'd254} : s = 289;
	{8'd35,8'd255} : s = 290;
	{8'd36,8'd0} : s = 36;
	{8'd36,8'd1} : s = 37;
	{8'd36,8'd2} : s = 38;
	{8'd36,8'd3} : s = 39;
	{8'd36,8'd4} : s = 40;
	{8'd36,8'd5} : s = 41;
	{8'd36,8'd6} : s = 42;
	{8'd36,8'd7} : s = 43;
	{8'd36,8'd8} : s = 44;
	{8'd36,8'd9} : s = 45;
	{8'd36,8'd10} : s = 46;
	{8'd36,8'd11} : s = 47;
	{8'd36,8'd12} : s = 48;
	{8'd36,8'd13} : s = 49;
	{8'd36,8'd14} : s = 50;
	{8'd36,8'd15} : s = 51;
	{8'd36,8'd16} : s = 52;
	{8'd36,8'd17} : s = 53;
	{8'd36,8'd18} : s = 54;
	{8'd36,8'd19} : s = 55;
	{8'd36,8'd20} : s = 56;
	{8'd36,8'd21} : s = 57;
	{8'd36,8'd22} : s = 58;
	{8'd36,8'd23} : s = 59;
	{8'd36,8'd24} : s = 60;
	{8'd36,8'd25} : s = 61;
	{8'd36,8'd26} : s = 62;
	{8'd36,8'd27} : s = 63;
	{8'd36,8'd28} : s = 64;
	{8'd36,8'd29} : s = 65;
	{8'd36,8'd30} : s = 66;
	{8'd36,8'd31} : s = 67;
	{8'd36,8'd32} : s = 68;
	{8'd36,8'd33} : s = 69;
	{8'd36,8'd34} : s = 70;
	{8'd36,8'd35} : s = 71;
	{8'd36,8'd36} : s = 72;
	{8'd36,8'd37} : s = 73;
	{8'd36,8'd38} : s = 74;
	{8'd36,8'd39} : s = 75;
	{8'd36,8'd40} : s = 76;
	{8'd36,8'd41} : s = 77;
	{8'd36,8'd42} : s = 78;
	{8'd36,8'd43} : s = 79;
	{8'd36,8'd44} : s = 80;
	{8'd36,8'd45} : s = 81;
	{8'd36,8'd46} : s = 82;
	{8'd36,8'd47} : s = 83;
	{8'd36,8'd48} : s = 84;
	{8'd36,8'd49} : s = 85;
	{8'd36,8'd50} : s = 86;
	{8'd36,8'd51} : s = 87;
	{8'd36,8'd52} : s = 88;
	{8'd36,8'd53} : s = 89;
	{8'd36,8'd54} : s = 90;
	{8'd36,8'd55} : s = 91;
	{8'd36,8'd56} : s = 92;
	{8'd36,8'd57} : s = 93;
	{8'd36,8'd58} : s = 94;
	{8'd36,8'd59} : s = 95;
	{8'd36,8'd60} : s = 96;
	{8'd36,8'd61} : s = 97;
	{8'd36,8'd62} : s = 98;
	{8'd36,8'd63} : s = 99;
	{8'd36,8'd64} : s = 100;
	{8'd36,8'd65} : s = 101;
	{8'd36,8'd66} : s = 102;
	{8'd36,8'd67} : s = 103;
	{8'd36,8'd68} : s = 104;
	{8'd36,8'd69} : s = 105;
	{8'd36,8'd70} : s = 106;
	{8'd36,8'd71} : s = 107;
	{8'd36,8'd72} : s = 108;
	{8'd36,8'd73} : s = 109;
	{8'd36,8'd74} : s = 110;
	{8'd36,8'd75} : s = 111;
	{8'd36,8'd76} : s = 112;
	{8'd36,8'd77} : s = 113;
	{8'd36,8'd78} : s = 114;
	{8'd36,8'd79} : s = 115;
	{8'd36,8'd80} : s = 116;
	{8'd36,8'd81} : s = 117;
	{8'd36,8'd82} : s = 118;
	{8'd36,8'd83} : s = 119;
	{8'd36,8'd84} : s = 120;
	{8'd36,8'd85} : s = 121;
	{8'd36,8'd86} : s = 122;
	{8'd36,8'd87} : s = 123;
	{8'd36,8'd88} : s = 124;
	{8'd36,8'd89} : s = 125;
	{8'd36,8'd90} : s = 126;
	{8'd36,8'd91} : s = 127;
	{8'd36,8'd92} : s = 128;
	{8'd36,8'd93} : s = 129;
	{8'd36,8'd94} : s = 130;
	{8'd36,8'd95} : s = 131;
	{8'd36,8'd96} : s = 132;
	{8'd36,8'd97} : s = 133;
	{8'd36,8'd98} : s = 134;
	{8'd36,8'd99} : s = 135;
	{8'd36,8'd100} : s = 136;
	{8'd36,8'd101} : s = 137;
	{8'd36,8'd102} : s = 138;
	{8'd36,8'd103} : s = 139;
	{8'd36,8'd104} : s = 140;
	{8'd36,8'd105} : s = 141;
	{8'd36,8'd106} : s = 142;
	{8'd36,8'd107} : s = 143;
	{8'd36,8'd108} : s = 144;
	{8'd36,8'd109} : s = 145;
	{8'd36,8'd110} : s = 146;
	{8'd36,8'd111} : s = 147;
	{8'd36,8'd112} : s = 148;
	{8'd36,8'd113} : s = 149;
	{8'd36,8'd114} : s = 150;
	{8'd36,8'd115} : s = 151;
	{8'd36,8'd116} : s = 152;
	{8'd36,8'd117} : s = 153;
	{8'd36,8'd118} : s = 154;
	{8'd36,8'd119} : s = 155;
	{8'd36,8'd120} : s = 156;
	{8'd36,8'd121} : s = 157;
	{8'd36,8'd122} : s = 158;
	{8'd36,8'd123} : s = 159;
	{8'd36,8'd124} : s = 160;
	{8'd36,8'd125} : s = 161;
	{8'd36,8'd126} : s = 162;
	{8'd36,8'd127} : s = 163;
	{8'd36,8'd128} : s = 164;
	{8'd36,8'd129} : s = 165;
	{8'd36,8'd130} : s = 166;
	{8'd36,8'd131} : s = 167;
	{8'd36,8'd132} : s = 168;
	{8'd36,8'd133} : s = 169;
	{8'd36,8'd134} : s = 170;
	{8'd36,8'd135} : s = 171;
	{8'd36,8'd136} : s = 172;
	{8'd36,8'd137} : s = 173;
	{8'd36,8'd138} : s = 174;
	{8'd36,8'd139} : s = 175;
	{8'd36,8'd140} : s = 176;
	{8'd36,8'd141} : s = 177;
	{8'd36,8'd142} : s = 178;
	{8'd36,8'd143} : s = 179;
	{8'd36,8'd144} : s = 180;
	{8'd36,8'd145} : s = 181;
	{8'd36,8'd146} : s = 182;
	{8'd36,8'd147} : s = 183;
	{8'd36,8'd148} : s = 184;
	{8'd36,8'd149} : s = 185;
	{8'd36,8'd150} : s = 186;
	{8'd36,8'd151} : s = 187;
	{8'd36,8'd152} : s = 188;
	{8'd36,8'd153} : s = 189;
	{8'd36,8'd154} : s = 190;
	{8'd36,8'd155} : s = 191;
	{8'd36,8'd156} : s = 192;
	{8'd36,8'd157} : s = 193;
	{8'd36,8'd158} : s = 194;
	{8'd36,8'd159} : s = 195;
	{8'd36,8'd160} : s = 196;
	{8'd36,8'd161} : s = 197;
	{8'd36,8'd162} : s = 198;
	{8'd36,8'd163} : s = 199;
	{8'd36,8'd164} : s = 200;
	{8'd36,8'd165} : s = 201;
	{8'd36,8'd166} : s = 202;
	{8'd36,8'd167} : s = 203;
	{8'd36,8'd168} : s = 204;
	{8'd36,8'd169} : s = 205;
	{8'd36,8'd170} : s = 206;
	{8'd36,8'd171} : s = 207;
	{8'd36,8'd172} : s = 208;
	{8'd36,8'd173} : s = 209;
	{8'd36,8'd174} : s = 210;
	{8'd36,8'd175} : s = 211;
	{8'd36,8'd176} : s = 212;
	{8'd36,8'd177} : s = 213;
	{8'd36,8'd178} : s = 214;
	{8'd36,8'd179} : s = 215;
	{8'd36,8'd180} : s = 216;
	{8'd36,8'd181} : s = 217;
	{8'd36,8'd182} : s = 218;
	{8'd36,8'd183} : s = 219;
	{8'd36,8'd184} : s = 220;
	{8'd36,8'd185} : s = 221;
	{8'd36,8'd186} : s = 222;
	{8'd36,8'd187} : s = 223;
	{8'd36,8'd188} : s = 224;
	{8'd36,8'd189} : s = 225;
	{8'd36,8'd190} : s = 226;
	{8'd36,8'd191} : s = 227;
	{8'd36,8'd192} : s = 228;
	{8'd36,8'd193} : s = 229;
	{8'd36,8'd194} : s = 230;
	{8'd36,8'd195} : s = 231;
	{8'd36,8'd196} : s = 232;
	{8'd36,8'd197} : s = 233;
	{8'd36,8'd198} : s = 234;
	{8'd36,8'd199} : s = 235;
	{8'd36,8'd200} : s = 236;
	{8'd36,8'd201} : s = 237;
	{8'd36,8'd202} : s = 238;
	{8'd36,8'd203} : s = 239;
	{8'd36,8'd204} : s = 240;
	{8'd36,8'd205} : s = 241;
	{8'd36,8'd206} : s = 242;
	{8'd36,8'd207} : s = 243;
	{8'd36,8'd208} : s = 244;
	{8'd36,8'd209} : s = 245;
	{8'd36,8'd210} : s = 246;
	{8'd36,8'd211} : s = 247;
	{8'd36,8'd212} : s = 248;
	{8'd36,8'd213} : s = 249;
	{8'd36,8'd214} : s = 250;
	{8'd36,8'd215} : s = 251;
	{8'd36,8'd216} : s = 252;
	{8'd36,8'd217} : s = 253;
	{8'd36,8'd218} : s = 254;
	{8'd36,8'd219} : s = 255;
	{8'd36,8'd220} : s = 256;
	{8'd36,8'd221} : s = 257;
	{8'd36,8'd222} : s = 258;
	{8'd36,8'd223} : s = 259;
	{8'd36,8'd224} : s = 260;
	{8'd36,8'd225} : s = 261;
	{8'd36,8'd226} : s = 262;
	{8'd36,8'd227} : s = 263;
	{8'd36,8'd228} : s = 264;
	{8'd36,8'd229} : s = 265;
	{8'd36,8'd230} : s = 266;
	{8'd36,8'd231} : s = 267;
	{8'd36,8'd232} : s = 268;
	{8'd36,8'd233} : s = 269;
	{8'd36,8'd234} : s = 270;
	{8'd36,8'd235} : s = 271;
	{8'd36,8'd236} : s = 272;
	{8'd36,8'd237} : s = 273;
	{8'd36,8'd238} : s = 274;
	{8'd36,8'd239} : s = 275;
	{8'd36,8'd240} : s = 276;
	{8'd36,8'd241} : s = 277;
	{8'd36,8'd242} : s = 278;
	{8'd36,8'd243} : s = 279;
	{8'd36,8'd244} : s = 280;
	{8'd36,8'd245} : s = 281;
	{8'd36,8'd246} : s = 282;
	{8'd36,8'd247} : s = 283;
	{8'd36,8'd248} : s = 284;
	{8'd36,8'd249} : s = 285;
	{8'd36,8'd250} : s = 286;
	{8'd36,8'd251} : s = 287;
	{8'd36,8'd252} : s = 288;
	{8'd36,8'd253} : s = 289;
	{8'd36,8'd254} : s = 290;
	{8'd36,8'd255} : s = 291;
	{8'd37,8'd0} : s = 37;
	{8'd37,8'd1} : s = 38;
	{8'd37,8'd2} : s = 39;
	{8'd37,8'd3} : s = 40;
	{8'd37,8'd4} : s = 41;
	{8'd37,8'd5} : s = 42;
	{8'd37,8'd6} : s = 43;
	{8'd37,8'd7} : s = 44;
	{8'd37,8'd8} : s = 45;
	{8'd37,8'd9} : s = 46;
	{8'd37,8'd10} : s = 47;
	{8'd37,8'd11} : s = 48;
	{8'd37,8'd12} : s = 49;
	{8'd37,8'd13} : s = 50;
	{8'd37,8'd14} : s = 51;
	{8'd37,8'd15} : s = 52;
	{8'd37,8'd16} : s = 53;
	{8'd37,8'd17} : s = 54;
	{8'd37,8'd18} : s = 55;
	{8'd37,8'd19} : s = 56;
	{8'd37,8'd20} : s = 57;
	{8'd37,8'd21} : s = 58;
	{8'd37,8'd22} : s = 59;
	{8'd37,8'd23} : s = 60;
	{8'd37,8'd24} : s = 61;
	{8'd37,8'd25} : s = 62;
	{8'd37,8'd26} : s = 63;
	{8'd37,8'd27} : s = 64;
	{8'd37,8'd28} : s = 65;
	{8'd37,8'd29} : s = 66;
	{8'd37,8'd30} : s = 67;
	{8'd37,8'd31} : s = 68;
	{8'd37,8'd32} : s = 69;
	{8'd37,8'd33} : s = 70;
	{8'd37,8'd34} : s = 71;
	{8'd37,8'd35} : s = 72;
	{8'd37,8'd36} : s = 73;
	{8'd37,8'd37} : s = 74;
	{8'd37,8'd38} : s = 75;
	{8'd37,8'd39} : s = 76;
	{8'd37,8'd40} : s = 77;
	{8'd37,8'd41} : s = 78;
	{8'd37,8'd42} : s = 79;
	{8'd37,8'd43} : s = 80;
	{8'd37,8'd44} : s = 81;
	{8'd37,8'd45} : s = 82;
	{8'd37,8'd46} : s = 83;
	{8'd37,8'd47} : s = 84;
	{8'd37,8'd48} : s = 85;
	{8'd37,8'd49} : s = 86;
	{8'd37,8'd50} : s = 87;
	{8'd37,8'd51} : s = 88;
	{8'd37,8'd52} : s = 89;
	{8'd37,8'd53} : s = 90;
	{8'd37,8'd54} : s = 91;
	{8'd37,8'd55} : s = 92;
	{8'd37,8'd56} : s = 93;
	{8'd37,8'd57} : s = 94;
	{8'd37,8'd58} : s = 95;
	{8'd37,8'd59} : s = 96;
	{8'd37,8'd60} : s = 97;
	{8'd37,8'd61} : s = 98;
	{8'd37,8'd62} : s = 99;
	{8'd37,8'd63} : s = 100;
	{8'd37,8'd64} : s = 101;
	{8'd37,8'd65} : s = 102;
	{8'd37,8'd66} : s = 103;
	{8'd37,8'd67} : s = 104;
	{8'd37,8'd68} : s = 105;
	{8'd37,8'd69} : s = 106;
	{8'd37,8'd70} : s = 107;
	{8'd37,8'd71} : s = 108;
	{8'd37,8'd72} : s = 109;
	{8'd37,8'd73} : s = 110;
	{8'd37,8'd74} : s = 111;
	{8'd37,8'd75} : s = 112;
	{8'd37,8'd76} : s = 113;
	{8'd37,8'd77} : s = 114;
	{8'd37,8'd78} : s = 115;
	{8'd37,8'd79} : s = 116;
	{8'd37,8'd80} : s = 117;
	{8'd37,8'd81} : s = 118;
	{8'd37,8'd82} : s = 119;
	{8'd37,8'd83} : s = 120;
	{8'd37,8'd84} : s = 121;
	{8'd37,8'd85} : s = 122;
	{8'd37,8'd86} : s = 123;
	{8'd37,8'd87} : s = 124;
	{8'd37,8'd88} : s = 125;
	{8'd37,8'd89} : s = 126;
	{8'd37,8'd90} : s = 127;
	{8'd37,8'd91} : s = 128;
	{8'd37,8'd92} : s = 129;
	{8'd37,8'd93} : s = 130;
	{8'd37,8'd94} : s = 131;
	{8'd37,8'd95} : s = 132;
	{8'd37,8'd96} : s = 133;
	{8'd37,8'd97} : s = 134;
	{8'd37,8'd98} : s = 135;
	{8'd37,8'd99} : s = 136;
	{8'd37,8'd100} : s = 137;
	{8'd37,8'd101} : s = 138;
	{8'd37,8'd102} : s = 139;
	{8'd37,8'd103} : s = 140;
	{8'd37,8'd104} : s = 141;
	{8'd37,8'd105} : s = 142;
	{8'd37,8'd106} : s = 143;
	{8'd37,8'd107} : s = 144;
	{8'd37,8'd108} : s = 145;
	{8'd37,8'd109} : s = 146;
	{8'd37,8'd110} : s = 147;
	{8'd37,8'd111} : s = 148;
	{8'd37,8'd112} : s = 149;
	{8'd37,8'd113} : s = 150;
	{8'd37,8'd114} : s = 151;
	{8'd37,8'd115} : s = 152;
	{8'd37,8'd116} : s = 153;
	{8'd37,8'd117} : s = 154;
	{8'd37,8'd118} : s = 155;
	{8'd37,8'd119} : s = 156;
	{8'd37,8'd120} : s = 157;
	{8'd37,8'd121} : s = 158;
	{8'd37,8'd122} : s = 159;
	{8'd37,8'd123} : s = 160;
	{8'd37,8'd124} : s = 161;
	{8'd37,8'd125} : s = 162;
	{8'd37,8'd126} : s = 163;
	{8'd37,8'd127} : s = 164;
	{8'd37,8'd128} : s = 165;
	{8'd37,8'd129} : s = 166;
	{8'd37,8'd130} : s = 167;
	{8'd37,8'd131} : s = 168;
	{8'd37,8'd132} : s = 169;
	{8'd37,8'd133} : s = 170;
	{8'd37,8'd134} : s = 171;
	{8'd37,8'd135} : s = 172;
	{8'd37,8'd136} : s = 173;
	{8'd37,8'd137} : s = 174;
	{8'd37,8'd138} : s = 175;
	{8'd37,8'd139} : s = 176;
	{8'd37,8'd140} : s = 177;
	{8'd37,8'd141} : s = 178;
	{8'd37,8'd142} : s = 179;
	{8'd37,8'd143} : s = 180;
	{8'd37,8'd144} : s = 181;
	{8'd37,8'd145} : s = 182;
	{8'd37,8'd146} : s = 183;
	{8'd37,8'd147} : s = 184;
	{8'd37,8'd148} : s = 185;
	{8'd37,8'd149} : s = 186;
	{8'd37,8'd150} : s = 187;
	{8'd37,8'd151} : s = 188;
	{8'd37,8'd152} : s = 189;
	{8'd37,8'd153} : s = 190;
	{8'd37,8'd154} : s = 191;
	{8'd37,8'd155} : s = 192;
	{8'd37,8'd156} : s = 193;
	{8'd37,8'd157} : s = 194;
	{8'd37,8'd158} : s = 195;
	{8'd37,8'd159} : s = 196;
	{8'd37,8'd160} : s = 197;
	{8'd37,8'd161} : s = 198;
	{8'd37,8'd162} : s = 199;
	{8'd37,8'd163} : s = 200;
	{8'd37,8'd164} : s = 201;
	{8'd37,8'd165} : s = 202;
	{8'd37,8'd166} : s = 203;
	{8'd37,8'd167} : s = 204;
	{8'd37,8'd168} : s = 205;
	{8'd37,8'd169} : s = 206;
	{8'd37,8'd170} : s = 207;
	{8'd37,8'd171} : s = 208;
	{8'd37,8'd172} : s = 209;
	{8'd37,8'd173} : s = 210;
	{8'd37,8'd174} : s = 211;
	{8'd37,8'd175} : s = 212;
	{8'd37,8'd176} : s = 213;
	{8'd37,8'd177} : s = 214;
	{8'd37,8'd178} : s = 215;
	{8'd37,8'd179} : s = 216;
	{8'd37,8'd180} : s = 217;
	{8'd37,8'd181} : s = 218;
	{8'd37,8'd182} : s = 219;
	{8'd37,8'd183} : s = 220;
	{8'd37,8'd184} : s = 221;
	{8'd37,8'd185} : s = 222;
	{8'd37,8'd186} : s = 223;
	{8'd37,8'd187} : s = 224;
	{8'd37,8'd188} : s = 225;
	{8'd37,8'd189} : s = 226;
	{8'd37,8'd190} : s = 227;
	{8'd37,8'd191} : s = 228;
	{8'd37,8'd192} : s = 229;
	{8'd37,8'd193} : s = 230;
	{8'd37,8'd194} : s = 231;
	{8'd37,8'd195} : s = 232;
	{8'd37,8'd196} : s = 233;
	{8'd37,8'd197} : s = 234;
	{8'd37,8'd198} : s = 235;
	{8'd37,8'd199} : s = 236;
	{8'd37,8'd200} : s = 237;
	{8'd37,8'd201} : s = 238;
	{8'd37,8'd202} : s = 239;
	{8'd37,8'd203} : s = 240;
	{8'd37,8'd204} : s = 241;
	{8'd37,8'd205} : s = 242;
	{8'd37,8'd206} : s = 243;
	{8'd37,8'd207} : s = 244;
	{8'd37,8'd208} : s = 245;
	{8'd37,8'd209} : s = 246;
	{8'd37,8'd210} : s = 247;
	{8'd37,8'd211} : s = 248;
	{8'd37,8'd212} : s = 249;
	{8'd37,8'd213} : s = 250;
	{8'd37,8'd214} : s = 251;
	{8'd37,8'd215} : s = 252;
	{8'd37,8'd216} : s = 253;
	{8'd37,8'd217} : s = 254;
	{8'd37,8'd218} : s = 255;
	{8'd37,8'd219} : s = 256;
	{8'd37,8'd220} : s = 257;
	{8'd37,8'd221} : s = 258;
	{8'd37,8'd222} : s = 259;
	{8'd37,8'd223} : s = 260;
	{8'd37,8'd224} : s = 261;
	{8'd37,8'd225} : s = 262;
	{8'd37,8'd226} : s = 263;
	{8'd37,8'd227} : s = 264;
	{8'd37,8'd228} : s = 265;
	{8'd37,8'd229} : s = 266;
	{8'd37,8'd230} : s = 267;
	{8'd37,8'd231} : s = 268;
	{8'd37,8'd232} : s = 269;
	{8'd37,8'd233} : s = 270;
	{8'd37,8'd234} : s = 271;
	{8'd37,8'd235} : s = 272;
	{8'd37,8'd236} : s = 273;
	{8'd37,8'd237} : s = 274;
	{8'd37,8'd238} : s = 275;
	{8'd37,8'd239} : s = 276;
	{8'd37,8'd240} : s = 277;
	{8'd37,8'd241} : s = 278;
	{8'd37,8'd242} : s = 279;
	{8'd37,8'd243} : s = 280;
	{8'd37,8'd244} : s = 281;
	{8'd37,8'd245} : s = 282;
	{8'd37,8'd246} : s = 283;
	{8'd37,8'd247} : s = 284;
	{8'd37,8'd248} : s = 285;
	{8'd37,8'd249} : s = 286;
	{8'd37,8'd250} : s = 287;
	{8'd37,8'd251} : s = 288;
	{8'd37,8'd252} : s = 289;
	{8'd37,8'd253} : s = 290;
	{8'd37,8'd254} : s = 291;
	{8'd37,8'd255} : s = 292;
	{8'd38,8'd0} : s = 38;
	{8'd38,8'd1} : s = 39;
	{8'd38,8'd2} : s = 40;
	{8'd38,8'd3} : s = 41;
	{8'd38,8'd4} : s = 42;
	{8'd38,8'd5} : s = 43;
	{8'd38,8'd6} : s = 44;
	{8'd38,8'd7} : s = 45;
	{8'd38,8'd8} : s = 46;
	{8'd38,8'd9} : s = 47;
	{8'd38,8'd10} : s = 48;
	{8'd38,8'd11} : s = 49;
	{8'd38,8'd12} : s = 50;
	{8'd38,8'd13} : s = 51;
	{8'd38,8'd14} : s = 52;
	{8'd38,8'd15} : s = 53;
	{8'd38,8'd16} : s = 54;
	{8'd38,8'd17} : s = 55;
	{8'd38,8'd18} : s = 56;
	{8'd38,8'd19} : s = 57;
	{8'd38,8'd20} : s = 58;
	{8'd38,8'd21} : s = 59;
	{8'd38,8'd22} : s = 60;
	{8'd38,8'd23} : s = 61;
	{8'd38,8'd24} : s = 62;
	{8'd38,8'd25} : s = 63;
	{8'd38,8'd26} : s = 64;
	{8'd38,8'd27} : s = 65;
	{8'd38,8'd28} : s = 66;
	{8'd38,8'd29} : s = 67;
	{8'd38,8'd30} : s = 68;
	{8'd38,8'd31} : s = 69;
	{8'd38,8'd32} : s = 70;
	{8'd38,8'd33} : s = 71;
	{8'd38,8'd34} : s = 72;
	{8'd38,8'd35} : s = 73;
	{8'd38,8'd36} : s = 74;
	{8'd38,8'd37} : s = 75;
	{8'd38,8'd38} : s = 76;
	{8'd38,8'd39} : s = 77;
	{8'd38,8'd40} : s = 78;
	{8'd38,8'd41} : s = 79;
	{8'd38,8'd42} : s = 80;
	{8'd38,8'd43} : s = 81;
	{8'd38,8'd44} : s = 82;
	{8'd38,8'd45} : s = 83;
	{8'd38,8'd46} : s = 84;
	{8'd38,8'd47} : s = 85;
	{8'd38,8'd48} : s = 86;
	{8'd38,8'd49} : s = 87;
	{8'd38,8'd50} : s = 88;
	{8'd38,8'd51} : s = 89;
	{8'd38,8'd52} : s = 90;
	{8'd38,8'd53} : s = 91;
	{8'd38,8'd54} : s = 92;
	{8'd38,8'd55} : s = 93;
	{8'd38,8'd56} : s = 94;
	{8'd38,8'd57} : s = 95;
	{8'd38,8'd58} : s = 96;
	{8'd38,8'd59} : s = 97;
	{8'd38,8'd60} : s = 98;
	{8'd38,8'd61} : s = 99;
	{8'd38,8'd62} : s = 100;
	{8'd38,8'd63} : s = 101;
	{8'd38,8'd64} : s = 102;
	{8'd38,8'd65} : s = 103;
	{8'd38,8'd66} : s = 104;
	{8'd38,8'd67} : s = 105;
	{8'd38,8'd68} : s = 106;
	{8'd38,8'd69} : s = 107;
	{8'd38,8'd70} : s = 108;
	{8'd38,8'd71} : s = 109;
	{8'd38,8'd72} : s = 110;
	{8'd38,8'd73} : s = 111;
	{8'd38,8'd74} : s = 112;
	{8'd38,8'd75} : s = 113;
	{8'd38,8'd76} : s = 114;
	{8'd38,8'd77} : s = 115;
	{8'd38,8'd78} : s = 116;
	{8'd38,8'd79} : s = 117;
	{8'd38,8'd80} : s = 118;
	{8'd38,8'd81} : s = 119;
	{8'd38,8'd82} : s = 120;
	{8'd38,8'd83} : s = 121;
	{8'd38,8'd84} : s = 122;
	{8'd38,8'd85} : s = 123;
	{8'd38,8'd86} : s = 124;
	{8'd38,8'd87} : s = 125;
	{8'd38,8'd88} : s = 126;
	{8'd38,8'd89} : s = 127;
	{8'd38,8'd90} : s = 128;
	{8'd38,8'd91} : s = 129;
	{8'd38,8'd92} : s = 130;
	{8'd38,8'd93} : s = 131;
	{8'd38,8'd94} : s = 132;
	{8'd38,8'd95} : s = 133;
	{8'd38,8'd96} : s = 134;
	{8'd38,8'd97} : s = 135;
	{8'd38,8'd98} : s = 136;
	{8'd38,8'd99} : s = 137;
	{8'd38,8'd100} : s = 138;
	{8'd38,8'd101} : s = 139;
	{8'd38,8'd102} : s = 140;
	{8'd38,8'd103} : s = 141;
	{8'd38,8'd104} : s = 142;
	{8'd38,8'd105} : s = 143;
	{8'd38,8'd106} : s = 144;
	{8'd38,8'd107} : s = 145;
	{8'd38,8'd108} : s = 146;
	{8'd38,8'd109} : s = 147;
	{8'd38,8'd110} : s = 148;
	{8'd38,8'd111} : s = 149;
	{8'd38,8'd112} : s = 150;
	{8'd38,8'd113} : s = 151;
	{8'd38,8'd114} : s = 152;
	{8'd38,8'd115} : s = 153;
	{8'd38,8'd116} : s = 154;
	{8'd38,8'd117} : s = 155;
	{8'd38,8'd118} : s = 156;
	{8'd38,8'd119} : s = 157;
	{8'd38,8'd120} : s = 158;
	{8'd38,8'd121} : s = 159;
	{8'd38,8'd122} : s = 160;
	{8'd38,8'd123} : s = 161;
	{8'd38,8'd124} : s = 162;
	{8'd38,8'd125} : s = 163;
	{8'd38,8'd126} : s = 164;
	{8'd38,8'd127} : s = 165;
	{8'd38,8'd128} : s = 166;
	{8'd38,8'd129} : s = 167;
	{8'd38,8'd130} : s = 168;
	{8'd38,8'd131} : s = 169;
	{8'd38,8'd132} : s = 170;
	{8'd38,8'd133} : s = 171;
	{8'd38,8'd134} : s = 172;
	{8'd38,8'd135} : s = 173;
	{8'd38,8'd136} : s = 174;
	{8'd38,8'd137} : s = 175;
	{8'd38,8'd138} : s = 176;
	{8'd38,8'd139} : s = 177;
	{8'd38,8'd140} : s = 178;
	{8'd38,8'd141} : s = 179;
	{8'd38,8'd142} : s = 180;
	{8'd38,8'd143} : s = 181;
	{8'd38,8'd144} : s = 182;
	{8'd38,8'd145} : s = 183;
	{8'd38,8'd146} : s = 184;
	{8'd38,8'd147} : s = 185;
	{8'd38,8'd148} : s = 186;
	{8'd38,8'd149} : s = 187;
	{8'd38,8'd150} : s = 188;
	{8'd38,8'd151} : s = 189;
	{8'd38,8'd152} : s = 190;
	{8'd38,8'd153} : s = 191;
	{8'd38,8'd154} : s = 192;
	{8'd38,8'd155} : s = 193;
	{8'd38,8'd156} : s = 194;
	{8'd38,8'd157} : s = 195;
	{8'd38,8'd158} : s = 196;
	{8'd38,8'd159} : s = 197;
	{8'd38,8'd160} : s = 198;
	{8'd38,8'd161} : s = 199;
	{8'd38,8'd162} : s = 200;
	{8'd38,8'd163} : s = 201;
	{8'd38,8'd164} : s = 202;
	{8'd38,8'd165} : s = 203;
	{8'd38,8'd166} : s = 204;
	{8'd38,8'd167} : s = 205;
	{8'd38,8'd168} : s = 206;
	{8'd38,8'd169} : s = 207;
	{8'd38,8'd170} : s = 208;
	{8'd38,8'd171} : s = 209;
	{8'd38,8'd172} : s = 210;
	{8'd38,8'd173} : s = 211;
	{8'd38,8'd174} : s = 212;
	{8'd38,8'd175} : s = 213;
	{8'd38,8'd176} : s = 214;
	{8'd38,8'd177} : s = 215;
	{8'd38,8'd178} : s = 216;
	{8'd38,8'd179} : s = 217;
	{8'd38,8'd180} : s = 218;
	{8'd38,8'd181} : s = 219;
	{8'd38,8'd182} : s = 220;
	{8'd38,8'd183} : s = 221;
	{8'd38,8'd184} : s = 222;
	{8'd38,8'd185} : s = 223;
	{8'd38,8'd186} : s = 224;
	{8'd38,8'd187} : s = 225;
	{8'd38,8'd188} : s = 226;
	{8'd38,8'd189} : s = 227;
	{8'd38,8'd190} : s = 228;
	{8'd38,8'd191} : s = 229;
	{8'd38,8'd192} : s = 230;
	{8'd38,8'd193} : s = 231;
	{8'd38,8'd194} : s = 232;
	{8'd38,8'd195} : s = 233;
	{8'd38,8'd196} : s = 234;
	{8'd38,8'd197} : s = 235;
	{8'd38,8'd198} : s = 236;
	{8'd38,8'd199} : s = 237;
	{8'd38,8'd200} : s = 238;
	{8'd38,8'd201} : s = 239;
	{8'd38,8'd202} : s = 240;
	{8'd38,8'd203} : s = 241;
	{8'd38,8'd204} : s = 242;
	{8'd38,8'd205} : s = 243;
	{8'd38,8'd206} : s = 244;
	{8'd38,8'd207} : s = 245;
	{8'd38,8'd208} : s = 246;
	{8'd38,8'd209} : s = 247;
	{8'd38,8'd210} : s = 248;
	{8'd38,8'd211} : s = 249;
	{8'd38,8'd212} : s = 250;
	{8'd38,8'd213} : s = 251;
	{8'd38,8'd214} : s = 252;
	{8'd38,8'd215} : s = 253;
	{8'd38,8'd216} : s = 254;
	{8'd38,8'd217} : s = 255;
	{8'd38,8'd218} : s = 256;
	{8'd38,8'd219} : s = 257;
	{8'd38,8'd220} : s = 258;
	{8'd38,8'd221} : s = 259;
	{8'd38,8'd222} : s = 260;
	{8'd38,8'd223} : s = 261;
	{8'd38,8'd224} : s = 262;
	{8'd38,8'd225} : s = 263;
	{8'd38,8'd226} : s = 264;
	{8'd38,8'd227} : s = 265;
	{8'd38,8'd228} : s = 266;
	{8'd38,8'd229} : s = 267;
	{8'd38,8'd230} : s = 268;
	{8'd38,8'd231} : s = 269;
	{8'd38,8'd232} : s = 270;
	{8'd38,8'd233} : s = 271;
	{8'd38,8'd234} : s = 272;
	{8'd38,8'd235} : s = 273;
	{8'd38,8'd236} : s = 274;
	{8'd38,8'd237} : s = 275;
	{8'd38,8'd238} : s = 276;
	{8'd38,8'd239} : s = 277;
	{8'd38,8'd240} : s = 278;
	{8'd38,8'd241} : s = 279;
	{8'd38,8'd242} : s = 280;
	{8'd38,8'd243} : s = 281;
	{8'd38,8'd244} : s = 282;
	{8'd38,8'd245} : s = 283;
	{8'd38,8'd246} : s = 284;
	{8'd38,8'd247} : s = 285;
	{8'd38,8'd248} : s = 286;
	{8'd38,8'd249} : s = 287;
	{8'd38,8'd250} : s = 288;
	{8'd38,8'd251} : s = 289;
	{8'd38,8'd252} : s = 290;
	{8'd38,8'd253} : s = 291;
	{8'd38,8'd254} : s = 292;
	{8'd38,8'd255} : s = 293;
	{8'd39,8'd0} : s = 39;
	{8'd39,8'd1} : s = 40;
	{8'd39,8'd2} : s = 41;
	{8'd39,8'd3} : s = 42;
	{8'd39,8'd4} : s = 43;
	{8'd39,8'd5} : s = 44;
	{8'd39,8'd6} : s = 45;
	{8'd39,8'd7} : s = 46;
	{8'd39,8'd8} : s = 47;
	{8'd39,8'd9} : s = 48;
	{8'd39,8'd10} : s = 49;
	{8'd39,8'd11} : s = 50;
	{8'd39,8'd12} : s = 51;
	{8'd39,8'd13} : s = 52;
	{8'd39,8'd14} : s = 53;
	{8'd39,8'd15} : s = 54;
	{8'd39,8'd16} : s = 55;
	{8'd39,8'd17} : s = 56;
	{8'd39,8'd18} : s = 57;
	{8'd39,8'd19} : s = 58;
	{8'd39,8'd20} : s = 59;
	{8'd39,8'd21} : s = 60;
	{8'd39,8'd22} : s = 61;
	{8'd39,8'd23} : s = 62;
	{8'd39,8'd24} : s = 63;
	{8'd39,8'd25} : s = 64;
	{8'd39,8'd26} : s = 65;
	{8'd39,8'd27} : s = 66;
	{8'd39,8'd28} : s = 67;
	{8'd39,8'd29} : s = 68;
	{8'd39,8'd30} : s = 69;
	{8'd39,8'd31} : s = 70;
	{8'd39,8'd32} : s = 71;
	{8'd39,8'd33} : s = 72;
	{8'd39,8'd34} : s = 73;
	{8'd39,8'd35} : s = 74;
	{8'd39,8'd36} : s = 75;
	{8'd39,8'd37} : s = 76;
	{8'd39,8'd38} : s = 77;
	{8'd39,8'd39} : s = 78;
	{8'd39,8'd40} : s = 79;
	{8'd39,8'd41} : s = 80;
	{8'd39,8'd42} : s = 81;
	{8'd39,8'd43} : s = 82;
	{8'd39,8'd44} : s = 83;
	{8'd39,8'd45} : s = 84;
	{8'd39,8'd46} : s = 85;
	{8'd39,8'd47} : s = 86;
	{8'd39,8'd48} : s = 87;
	{8'd39,8'd49} : s = 88;
	{8'd39,8'd50} : s = 89;
	{8'd39,8'd51} : s = 90;
	{8'd39,8'd52} : s = 91;
	{8'd39,8'd53} : s = 92;
	{8'd39,8'd54} : s = 93;
	{8'd39,8'd55} : s = 94;
	{8'd39,8'd56} : s = 95;
	{8'd39,8'd57} : s = 96;
	{8'd39,8'd58} : s = 97;
	{8'd39,8'd59} : s = 98;
	{8'd39,8'd60} : s = 99;
	{8'd39,8'd61} : s = 100;
	{8'd39,8'd62} : s = 101;
	{8'd39,8'd63} : s = 102;
	{8'd39,8'd64} : s = 103;
	{8'd39,8'd65} : s = 104;
	{8'd39,8'd66} : s = 105;
	{8'd39,8'd67} : s = 106;
	{8'd39,8'd68} : s = 107;
	{8'd39,8'd69} : s = 108;
	{8'd39,8'd70} : s = 109;
	{8'd39,8'd71} : s = 110;
	{8'd39,8'd72} : s = 111;
	{8'd39,8'd73} : s = 112;
	{8'd39,8'd74} : s = 113;
	{8'd39,8'd75} : s = 114;
	{8'd39,8'd76} : s = 115;
	{8'd39,8'd77} : s = 116;
	{8'd39,8'd78} : s = 117;
	{8'd39,8'd79} : s = 118;
	{8'd39,8'd80} : s = 119;
	{8'd39,8'd81} : s = 120;
	{8'd39,8'd82} : s = 121;
	{8'd39,8'd83} : s = 122;
	{8'd39,8'd84} : s = 123;
	{8'd39,8'd85} : s = 124;
	{8'd39,8'd86} : s = 125;
	{8'd39,8'd87} : s = 126;
	{8'd39,8'd88} : s = 127;
	{8'd39,8'd89} : s = 128;
	{8'd39,8'd90} : s = 129;
	{8'd39,8'd91} : s = 130;
	{8'd39,8'd92} : s = 131;
	{8'd39,8'd93} : s = 132;
	{8'd39,8'd94} : s = 133;
	{8'd39,8'd95} : s = 134;
	{8'd39,8'd96} : s = 135;
	{8'd39,8'd97} : s = 136;
	{8'd39,8'd98} : s = 137;
	{8'd39,8'd99} : s = 138;
	{8'd39,8'd100} : s = 139;
	{8'd39,8'd101} : s = 140;
	{8'd39,8'd102} : s = 141;
	{8'd39,8'd103} : s = 142;
	{8'd39,8'd104} : s = 143;
	{8'd39,8'd105} : s = 144;
	{8'd39,8'd106} : s = 145;
	{8'd39,8'd107} : s = 146;
	{8'd39,8'd108} : s = 147;
	{8'd39,8'd109} : s = 148;
	{8'd39,8'd110} : s = 149;
	{8'd39,8'd111} : s = 150;
	{8'd39,8'd112} : s = 151;
	{8'd39,8'd113} : s = 152;
	{8'd39,8'd114} : s = 153;
	{8'd39,8'd115} : s = 154;
	{8'd39,8'd116} : s = 155;
	{8'd39,8'd117} : s = 156;
	{8'd39,8'd118} : s = 157;
	{8'd39,8'd119} : s = 158;
	{8'd39,8'd120} : s = 159;
	{8'd39,8'd121} : s = 160;
	{8'd39,8'd122} : s = 161;
	{8'd39,8'd123} : s = 162;
	{8'd39,8'd124} : s = 163;
	{8'd39,8'd125} : s = 164;
	{8'd39,8'd126} : s = 165;
	{8'd39,8'd127} : s = 166;
	{8'd39,8'd128} : s = 167;
	{8'd39,8'd129} : s = 168;
	{8'd39,8'd130} : s = 169;
	{8'd39,8'd131} : s = 170;
	{8'd39,8'd132} : s = 171;
	{8'd39,8'd133} : s = 172;
	{8'd39,8'd134} : s = 173;
	{8'd39,8'd135} : s = 174;
	{8'd39,8'd136} : s = 175;
	{8'd39,8'd137} : s = 176;
	{8'd39,8'd138} : s = 177;
	{8'd39,8'd139} : s = 178;
	{8'd39,8'd140} : s = 179;
	{8'd39,8'd141} : s = 180;
	{8'd39,8'd142} : s = 181;
	{8'd39,8'd143} : s = 182;
	{8'd39,8'd144} : s = 183;
	{8'd39,8'd145} : s = 184;
	{8'd39,8'd146} : s = 185;
	{8'd39,8'd147} : s = 186;
	{8'd39,8'd148} : s = 187;
	{8'd39,8'd149} : s = 188;
	{8'd39,8'd150} : s = 189;
	{8'd39,8'd151} : s = 190;
	{8'd39,8'd152} : s = 191;
	{8'd39,8'd153} : s = 192;
	{8'd39,8'd154} : s = 193;
	{8'd39,8'd155} : s = 194;
	{8'd39,8'd156} : s = 195;
	{8'd39,8'd157} : s = 196;
	{8'd39,8'd158} : s = 197;
	{8'd39,8'd159} : s = 198;
	{8'd39,8'd160} : s = 199;
	{8'd39,8'd161} : s = 200;
	{8'd39,8'd162} : s = 201;
	{8'd39,8'd163} : s = 202;
	{8'd39,8'd164} : s = 203;
	{8'd39,8'd165} : s = 204;
	{8'd39,8'd166} : s = 205;
	{8'd39,8'd167} : s = 206;
	{8'd39,8'd168} : s = 207;
	{8'd39,8'd169} : s = 208;
	{8'd39,8'd170} : s = 209;
	{8'd39,8'd171} : s = 210;
	{8'd39,8'd172} : s = 211;
	{8'd39,8'd173} : s = 212;
	{8'd39,8'd174} : s = 213;
	{8'd39,8'd175} : s = 214;
	{8'd39,8'd176} : s = 215;
	{8'd39,8'd177} : s = 216;
	{8'd39,8'd178} : s = 217;
	{8'd39,8'd179} : s = 218;
	{8'd39,8'd180} : s = 219;
	{8'd39,8'd181} : s = 220;
	{8'd39,8'd182} : s = 221;
	{8'd39,8'd183} : s = 222;
	{8'd39,8'd184} : s = 223;
	{8'd39,8'd185} : s = 224;
	{8'd39,8'd186} : s = 225;
	{8'd39,8'd187} : s = 226;
	{8'd39,8'd188} : s = 227;
	{8'd39,8'd189} : s = 228;
	{8'd39,8'd190} : s = 229;
	{8'd39,8'd191} : s = 230;
	{8'd39,8'd192} : s = 231;
	{8'd39,8'd193} : s = 232;
	{8'd39,8'd194} : s = 233;
	{8'd39,8'd195} : s = 234;
	{8'd39,8'd196} : s = 235;
	{8'd39,8'd197} : s = 236;
	{8'd39,8'd198} : s = 237;
	{8'd39,8'd199} : s = 238;
	{8'd39,8'd200} : s = 239;
	{8'd39,8'd201} : s = 240;
	{8'd39,8'd202} : s = 241;
	{8'd39,8'd203} : s = 242;
	{8'd39,8'd204} : s = 243;
	{8'd39,8'd205} : s = 244;
	{8'd39,8'd206} : s = 245;
	{8'd39,8'd207} : s = 246;
	{8'd39,8'd208} : s = 247;
	{8'd39,8'd209} : s = 248;
	{8'd39,8'd210} : s = 249;
	{8'd39,8'd211} : s = 250;
	{8'd39,8'd212} : s = 251;
	{8'd39,8'd213} : s = 252;
	{8'd39,8'd214} : s = 253;
	{8'd39,8'd215} : s = 254;
	{8'd39,8'd216} : s = 255;
	{8'd39,8'd217} : s = 256;
	{8'd39,8'd218} : s = 257;
	{8'd39,8'd219} : s = 258;
	{8'd39,8'd220} : s = 259;
	{8'd39,8'd221} : s = 260;
	{8'd39,8'd222} : s = 261;
	{8'd39,8'd223} : s = 262;
	{8'd39,8'd224} : s = 263;
	{8'd39,8'd225} : s = 264;
	{8'd39,8'd226} : s = 265;
	{8'd39,8'd227} : s = 266;
	{8'd39,8'd228} : s = 267;
	{8'd39,8'd229} : s = 268;
	{8'd39,8'd230} : s = 269;
	{8'd39,8'd231} : s = 270;
	{8'd39,8'd232} : s = 271;
	{8'd39,8'd233} : s = 272;
	{8'd39,8'd234} : s = 273;
	{8'd39,8'd235} : s = 274;
	{8'd39,8'd236} : s = 275;
	{8'd39,8'd237} : s = 276;
	{8'd39,8'd238} : s = 277;
	{8'd39,8'd239} : s = 278;
	{8'd39,8'd240} : s = 279;
	{8'd39,8'd241} : s = 280;
	{8'd39,8'd242} : s = 281;
	{8'd39,8'd243} : s = 282;
	{8'd39,8'd244} : s = 283;
	{8'd39,8'd245} : s = 284;
	{8'd39,8'd246} : s = 285;
	{8'd39,8'd247} : s = 286;
	{8'd39,8'd248} : s = 287;
	{8'd39,8'd249} : s = 288;
	{8'd39,8'd250} : s = 289;
	{8'd39,8'd251} : s = 290;
	{8'd39,8'd252} : s = 291;
	{8'd39,8'd253} : s = 292;
	{8'd39,8'd254} : s = 293;
	{8'd39,8'd255} : s = 294;
	{8'd40,8'd0} : s = 40;
	{8'd40,8'd1} : s = 41;
	{8'd40,8'd2} : s = 42;
	{8'd40,8'd3} : s = 43;
	{8'd40,8'd4} : s = 44;
	{8'd40,8'd5} : s = 45;
	{8'd40,8'd6} : s = 46;
	{8'd40,8'd7} : s = 47;
	{8'd40,8'd8} : s = 48;
	{8'd40,8'd9} : s = 49;
	{8'd40,8'd10} : s = 50;
	{8'd40,8'd11} : s = 51;
	{8'd40,8'd12} : s = 52;
	{8'd40,8'd13} : s = 53;
	{8'd40,8'd14} : s = 54;
	{8'd40,8'd15} : s = 55;
	{8'd40,8'd16} : s = 56;
	{8'd40,8'd17} : s = 57;
	{8'd40,8'd18} : s = 58;
	{8'd40,8'd19} : s = 59;
	{8'd40,8'd20} : s = 60;
	{8'd40,8'd21} : s = 61;
	{8'd40,8'd22} : s = 62;
	{8'd40,8'd23} : s = 63;
	{8'd40,8'd24} : s = 64;
	{8'd40,8'd25} : s = 65;
	{8'd40,8'd26} : s = 66;
	{8'd40,8'd27} : s = 67;
	{8'd40,8'd28} : s = 68;
	{8'd40,8'd29} : s = 69;
	{8'd40,8'd30} : s = 70;
	{8'd40,8'd31} : s = 71;
	{8'd40,8'd32} : s = 72;
	{8'd40,8'd33} : s = 73;
	{8'd40,8'd34} : s = 74;
	{8'd40,8'd35} : s = 75;
	{8'd40,8'd36} : s = 76;
	{8'd40,8'd37} : s = 77;
	{8'd40,8'd38} : s = 78;
	{8'd40,8'd39} : s = 79;
	{8'd40,8'd40} : s = 80;
	{8'd40,8'd41} : s = 81;
	{8'd40,8'd42} : s = 82;
	{8'd40,8'd43} : s = 83;
	{8'd40,8'd44} : s = 84;
	{8'd40,8'd45} : s = 85;
	{8'd40,8'd46} : s = 86;
	{8'd40,8'd47} : s = 87;
	{8'd40,8'd48} : s = 88;
	{8'd40,8'd49} : s = 89;
	{8'd40,8'd50} : s = 90;
	{8'd40,8'd51} : s = 91;
	{8'd40,8'd52} : s = 92;
	{8'd40,8'd53} : s = 93;
	{8'd40,8'd54} : s = 94;
	{8'd40,8'd55} : s = 95;
	{8'd40,8'd56} : s = 96;
	{8'd40,8'd57} : s = 97;
	{8'd40,8'd58} : s = 98;
	{8'd40,8'd59} : s = 99;
	{8'd40,8'd60} : s = 100;
	{8'd40,8'd61} : s = 101;
	{8'd40,8'd62} : s = 102;
	{8'd40,8'd63} : s = 103;
	{8'd40,8'd64} : s = 104;
	{8'd40,8'd65} : s = 105;
	{8'd40,8'd66} : s = 106;
	{8'd40,8'd67} : s = 107;
	{8'd40,8'd68} : s = 108;
	{8'd40,8'd69} : s = 109;
	{8'd40,8'd70} : s = 110;
	{8'd40,8'd71} : s = 111;
	{8'd40,8'd72} : s = 112;
	{8'd40,8'd73} : s = 113;
	{8'd40,8'd74} : s = 114;
	{8'd40,8'd75} : s = 115;
	{8'd40,8'd76} : s = 116;
	{8'd40,8'd77} : s = 117;
	{8'd40,8'd78} : s = 118;
	{8'd40,8'd79} : s = 119;
	{8'd40,8'd80} : s = 120;
	{8'd40,8'd81} : s = 121;
	{8'd40,8'd82} : s = 122;
	{8'd40,8'd83} : s = 123;
	{8'd40,8'd84} : s = 124;
	{8'd40,8'd85} : s = 125;
	{8'd40,8'd86} : s = 126;
	{8'd40,8'd87} : s = 127;
	{8'd40,8'd88} : s = 128;
	{8'd40,8'd89} : s = 129;
	{8'd40,8'd90} : s = 130;
	{8'd40,8'd91} : s = 131;
	{8'd40,8'd92} : s = 132;
	{8'd40,8'd93} : s = 133;
	{8'd40,8'd94} : s = 134;
	{8'd40,8'd95} : s = 135;
	{8'd40,8'd96} : s = 136;
	{8'd40,8'd97} : s = 137;
	{8'd40,8'd98} : s = 138;
	{8'd40,8'd99} : s = 139;
	{8'd40,8'd100} : s = 140;
	{8'd40,8'd101} : s = 141;
	{8'd40,8'd102} : s = 142;
	{8'd40,8'd103} : s = 143;
	{8'd40,8'd104} : s = 144;
	{8'd40,8'd105} : s = 145;
	{8'd40,8'd106} : s = 146;
	{8'd40,8'd107} : s = 147;
	{8'd40,8'd108} : s = 148;
	{8'd40,8'd109} : s = 149;
	{8'd40,8'd110} : s = 150;
	{8'd40,8'd111} : s = 151;
	{8'd40,8'd112} : s = 152;
	{8'd40,8'd113} : s = 153;
	{8'd40,8'd114} : s = 154;
	{8'd40,8'd115} : s = 155;
	{8'd40,8'd116} : s = 156;
	{8'd40,8'd117} : s = 157;
	{8'd40,8'd118} : s = 158;
	{8'd40,8'd119} : s = 159;
	{8'd40,8'd120} : s = 160;
	{8'd40,8'd121} : s = 161;
	{8'd40,8'd122} : s = 162;
	{8'd40,8'd123} : s = 163;
	{8'd40,8'd124} : s = 164;
	{8'd40,8'd125} : s = 165;
	{8'd40,8'd126} : s = 166;
	{8'd40,8'd127} : s = 167;
	{8'd40,8'd128} : s = 168;
	{8'd40,8'd129} : s = 169;
	{8'd40,8'd130} : s = 170;
	{8'd40,8'd131} : s = 171;
	{8'd40,8'd132} : s = 172;
	{8'd40,8'd133} : s = 173;
	{8'd40,8'd134} : s = 174;
	{8'd40,8'd135} : s = 175;
	{8'd40,8'd136} : s = 176;
	{8'd40,8'd137} : s = 177;
	{8'd40,8'd138} : s = 178;
	{8'd40,8'd139} : s = 179;
	{8'd40,8'd140} : s = 180;
	{8'd40,8'd141} : s = 181;
	{8'd40,8'd142} : s = 182;
	{8'd40,8'd143} : s = 183;
	{8'd40,8'd144} : s = 184;
	{8'd40,8'd145} : s = 185;
	{8'd40,8'd146} : s = 186;
	{8'd40,8'd147} : s = 187;
	{8'd40,8'd148} : s = 188;
	{8'd40,8'd149} : s = 189;
	{8'd40,8'd150} : s = 190;
	{8'd40,8'd151} : s = 191;
	{8'd40,8'd152} : s = 192;
	{8'd40,8'd153} : s = 193;
	{8'd40,8'd154} : s = 194;
	{8'd40,8'd155} : s = 195;
	{8'd40,8'd156} : s = 196;
	{8'd40,8'd157} : s = 197;
	{8'd40,8'd158} : s = 198;
	{8'd40,8'd159} : s = 199;
	{8'd40,8'd160} : s = 200;
	{8'd40,8'd161} : s = 201;
	{8'd40,8'd162} : s = 202;
	{8'd40,8'd163} : s = 203;
	{8'd40,8'd164} : s = 204;
	{8'd40,8'd165} : s = 205;
	{8'd40,8'd166} : s = 206;
	{8'd40,8'd167} : s = 207;
	{8'd40,8'd168} : s = 208;
	{8'd40,8'd169} : s = 209;
	{8'd40,8'd170} : s = 210;
	{8'd40,8'd171} : s = 211;
	{8'd40,8'd172} : s = 212;
	{8'd40,8'd173} : s = 213;
	{8'd40,8'd174} : s = 214;
	{8'd40,8'd175} : s = 215;
	{8'd40,8'd176} : s = 216;
	{8'd40,8'd177} : s = 217;
	{8'd40,8'd178} : s = 218;
	{8'd40,8'd179} : s = 219;
	{8'd40,8'd180} : s = 220;
	{8'd40,8'd181} : s = 221;
	{8'd40,8'd182} : s = 222;
	{8'd40,8'd183} : s = 223;
	{8'd40,8'd184} : s = 224;
	{8'd40,8'd185} : s = 225;
	{8'd40,8'd186} : s = 226;
	{8'd40,8'd187} : s = 227;
	{8'd40,8'd188} : s = 228;
	{8'd40,8'd189} : s = 229;
	{8'd40,8'd190} : s = 230;
	{8'd40,8'd191} : s = 231;
	{8'd40,8'd192} : s = 232;
	{8'd40,8'd193} : s = 233;
	{8'd40,8'd194} : s = 234;
	{8'd40,8'd195} : s = 235;
	{8'd40,8'd196} : s = 236;
	{8'd40,8'd197} : s = 237;
	{8'd40,8'd198} : s = 238;
	{8'd40,8'd199} : s = 239;
	{8'd40,8'd200} : s = 240;
	{8'd40,8'd201} : s = 241;
	{8'd40,8'd202} : s = 242;
	{8'd40,8'd203} : s = 243;
	{8'd40,8'd204} : s = 244;
	{8'd40,8'd205} : s = 245;
	{8'd40,8'd206} : s = 246;
	{8'd40,8'd207} : s = 247;
	{8'd40,8'd208} : s = 248;
	{8'd40,8'd209} : s = 249;
	{8'd40,8'd210} : s = 250;
	{8'd40,8'd211} : s = 251;
	{8'd40,8'd212} : s = 252;
	{8'd40,8'd213} : s = 253;
	{8'd40,8'd214} : s = 254;
	{8'd40,8'd215} : s = 255;
	{8'd40,8'd216} : s = 256;
	{8'd40,8'd217} : s = 257;
	{8'd40,8'd218} : s = 258;
	{8'd40,8'd219} : s = 259;
	{8'd40,8'd220} : s = 260;
	{8'd40,8'd221} : s = 261;
	{8'd40,8'd222} : s = 262;
	{8'd40,8'd223} : s = 263;
	{8'd40,8'd224} : s = 264;
	{8'd40,8'd225} : s = 265;
	{8'd40,8'd226} : s = 266;
	{8'd40,8'd227} : s = 267;
	{8'd40,8'd228} : s = 268;
	{8'd40,8'd229} : s = 269;
	{8'd40,8'd230} : s = 270;
	{8'd40,8'd231} : s = 271;
	{8'd40,8'd232} : s = 272;
	{8'd40,8'd233} : s = 273;
	{8'd40,8'd234} : s = 274;
	{8'd40,8'd235} : s = 275;
	{8'd40,8'd236} : s = 276;
	{8'd40,8'd237} : s = 277;
	{8'd40,8'd238} : s = 278;
	{8'd40,8'd239} : s = 279;
	{8'd40,8'd240} : s = 280;
	{8'd40,8'd241} : s = 281;
	{8'd40,8'd242} : s = 282;
	{8'd40,8'd243} : s = 283;
	{8'd40,8'd244} : s = 284;
	{8'd40,8'd245} : s = 285;
	{8'd40,8'd246} : s = 286;
	{8'd40,8'd247} : s = 287;
	{8'd40,8'd248} : s = 288;
	{8'd40,8'd249} : s = 289;
	{8'd40,8'd250} : s = 290;
	{8'd40,8'd251} : s = 291;
	{8'd40,8'd252} : s = 292;
	{8'd40,8'd253} : s = 293;
	{8'd40,8'd254} : s = 294;
	{8'd40,8'd255} : s = 295;
	{8'd41,8'd0} : s = 41;
	{8'd41,8'd1} : s = 42;
	{8'd41,8'd2} : s = 43;
	{8'd41,8'd3} : s = 44;
	{8'd41,8'd4} : s = 45;
	{8'd41,8'd5} : s = 46;
	{8'd41,8'd6} : s = 47;
	{8'd41,8'd7} : s = 48;
	{8'd41,8'd8} : s = 49;
	{8'd41,8'd9} : s = 50;
	{8'd41,8'd10} : s = 51;
	{8'd41,8'd11} : s = 52;
	{8'd41,8'd12} : s = 53;
	{8'd41,8'd13} : s = 54;
	{8'd41,8'd14} : s = 55;
	{8'd41,8'd15} : s = 56;
	{8'd41,8'd16} : s = 57;
	{8'd41,8'd17} : s = 58;
	{8'd41,8'd18} : s = 59;
	{8'd41,8'd19} : s = 60;
	{8'd41,8'd20} : s = 61;
	{8'd41,8'd21} : s = 62;
	{8'd41,8'd22} : s = 63;
	{8'd41,8'd23} : s = 64;
	{8'd41,8'd24} : s = 65;
	{8'd41,8'd25} : s = 66;
	{8'd41,8'd26} : s = 67;
	{8'd41,8'd27} : s = 68;
	{8'd41,8'd28} : s = 69;
	{8'd41,8'd29} : s = 70;
	{8'd41,8'd30} : s = 71;
	{8'd41,8'd31} : s = 72;
	{8'd41,8'd32} : s = 73;
	{8'd41,8'd33} : s = 74;
	{8'd41,8'd34} : s = 75;
	{8'd41,8'd35} : s = 76;
	{8'd41,8'd36} : s = 77;
	{8'd41,8'd37} : s = 78;
	{8'd41,8'd38} : s = 79;
	{8'd41,8'd39} : s = 80;
	{8'd41,8'd40} : s = 81;
	{8'd41,8'd41} : s = 82;
	{8'd41,8'd42} : s = 83;
	{8'd41,8'd43} : s = 84;
	{8'd41,8'd44} : s = 85;
	{8'd41,8'd45} : s = 86;
	{8'd41,8'd46} : s = 87;
	{8'd41,8'd47} : s = 88;
	{8'd41,8'd48} : s = 89;
	{8'd41,8'd49} : s = 90;
	{8'd41,8'd50} : s = 91;
	{8'd41,8'd51} : s = 92;
	{8'd41,8'd52} : s = 93;
	{8'd41,8'd53} : s = 94;
	{8'd41,8'd54} : s = 95;
	{8'd41,8'd55} : s = 96;
	{8'd41,8'd56} : s = 97;
	{8'd41,8'd57} : s = 98;
	{8'd41,8'd58} : s = 99;
	{8'd41,8'd59} : s = 100;
	{8'd41,8'd60} : s = 101;
	{8'd41,8'd61} : s = 102;
	{8'd41,8'd62} : s = 103;
	{8'd41,8'd63} : s = 104;
	{8'd41,8'd64} : s = 105;
	{8'd41,8'd65} : s = 106;
	{8'd41,8'd66} : s = 107;
	{8'd41,8'd67} : s = 108;
	{8'd41,8'd68} : s = 109;
	{8'd41,8'd69} : s = 110;
	{8'd41,8'd70} : s = 111;
	{8'd41,8'd71} : s = 112;
	{8'd41,8'd72} : s = 113;
	{8'd41,8'd73} : s = 114;
	{8'd41,8'd74} : s = 115;
	{8'd41,8'd75} : s = 116;
	{8'd41,8'd76} : s = 117;
	{8'd41,8'd77} : s = 118;
	{8'd41,8'd78} : s = 119;
	{8'd41,8'd79} : s = 120;
	{8'd41,8'd80} : s = 121;
	{8'd41,8'd81} : s = 122;
	{8'd41,8'd82} : s = 123;
	{8'd41,8'd83} : s = 124;
	{8'd41,8'd84} : s = 125;
	{8'd41,8'd85} : s = 126;
	{8'd41,8'd86} : s = 127;
	{8'd41,8'd87} : s = 128;
	{8'd41,8'd88} : s = 129;
	{8'd41,8'd89} : s = 130;
	{8'd41,8'd90} : s = 131;
	{8'd41,8'd91} : s = 132;
	{8'd41,8'd92} : s = 133;
	{8'd41,8'd93} : s = 134;
	{8'd41,8'd94} : s = 135;
	{8'd41,8'd95} : s = 136;
	{8'd41,8'd96} : s = 137;
	{8'd41,8'd97} : s = 138;
	{8'd41,8'd98} : s = 139;
	{8'd41,8'd99} : s = 140;
	{8'd41,8'd100} : s = 141;
	{8'd41,8'd101} : s = 142;
	{8'd41,8'd102} : s = 143;
	{8'd41,8'd103} : s = 144;
	{8'd41,8'd104} : s = 145;
	{8'd41,8'd105} : s = 146;
	{8'd41,8'd106} : s = 147;
	{8'd41,8'd107} : s = 148;
	{8'd41,8'd108} : s = 149;
	{8'd41,8'd109} : s = 150;
	{8'd41,8'd110} : s = 151;
	{8'd41,8'd111} : s = 152;
	{8'd41,8'd112} : s = 153;
	{8'd41,8'd113} : s = 154;
	{8'd41,8'd114} : s = 155;
	{8'd41,8'd115} : s = 156;
	{8'd41,8'd116} : s = 157;
	{8'd41,8'd117} : s = 158;
	{8'd41,8'd118} : s = 159;
	{8'd41,8'd119} : s = 160;
	{8'd41,8'd120} : s = 161;
	{8'd41,8'd121} : s = 162;
	{8'd41,8'd122} : s = 163;
	{8'd41,8'd123} : s = 164;
	{8'd41,8'd124} : s = 165;
	{8'd41,8'd125} : s = 166;
	{8'd41,8'd126} : s = 167;
	{8'd41,8'd127} : s = 168;
	{8'd41,8'd128} : s = 169;
	{8'd41,8'd129} : s = 170;
	{8'd41,8'd130} : s = 171;
	{8'd41,8'd131} : s = 172;
	{8'd41,8'd132} : s = 173;
	{8'd41,8'd133} : s = 174;
	{8'd41,8'd134} : s = 175;
	{8'd41,8'd135} : s = 176;
	{8'd41,8'd136} : s = 177;
	{8'd41,8'd137} : s = 178;
	{8'd41,8'd138} : s = 179;
	{8'd41,8'd139} : s = 180;
	{8'd41,8'd140} : s = 181;
	{8'd41,8'd141} : s = 182;
	{8'd41,8'd142} : s = 183;
	{8'd41,8'd143} : s = 184;
	{8'd41,8'd144} : s = 185;
	{8'd41,8'd145} : s = 186;
	{8'd41,8'd146} : s = 187;
	{8'd41,8'd147} : s = 188;
	{8'd41,8'd148} : s = 189;
	{8'd41,8'd149} : s = 190;
	{8'd41,8'd150} : s = 191;
	{8'd41,8'd151} : s = 192;
	{8'd41,8'd152} : s = 193;
	{8'd41,8'd153} : s = 194;
	{8'd41,8'd154} : s = 195;
	{8'd41,8'd155} : s = 196;
	{8'd41,8'd156} : s = 197;
	{8'd41,8'd157} : s = 198;
	{8'd41,8'd158} : s = 199;
	{8'd41,8'd159} : s = 200;
	{8'd41,8'd160} : s = 201;
	{8'd41,8'd161} : s = 202;
	{8'd41,8'd162} : s = 203;
	{8'd41,8'd163} : s = 204;
	{8'd41,8'd164} : s = 205;
	{8'd41,8'd165} : s = 206;
	{8'd41,8'd166} : s = 207;
	{8'd41,8'd167} : s = 208;
	{8'd41,8'd168} : s = 209;
	{8'd41,8'd169} : s = 210;
	{8'd41,8'd170} : s = 211;
	{8'd41,8'd171} : s = 212;
	{8'd41,8'd172} : s = 213;
	{8'd41,8'd173} : s = 214;
	{8'd41,8'd174} : s = 215;
	{8'd41,8'd175} : s = 216;
	{8'd41,8'd176} : s = 217;
	{8'd41,8'd177} : s = 218;
	{8'd41,8'd178} : s = 219;
	{8'd41,8'd179} : s = 220;
	{8'd41,8'd180} : s = 221;
	{8'd41,8'd181} : s = 222;
	{8'd41,8'd182} : s = 223;
	{8'd41,8'd183} : s = 224;
	{8'd41,8'd184} : s = 225;
	{8'd41,8'd185} : s = 226;
	{8'd41,8'd186} : s = 227;
	{8'd41,8'd187} : s = 228;
	{8'd41,8'd188} : s = 229;
	{8'd41,8'd189} : s = 230;
	{8'd41,8'd190} : s = 231;
	{8'd41,8'd191} : s = 232;
	{8'd41,8'd192} : s = 233;
	{8'd41,8'd193} : s = 234;
	{8'd41,8'd194} : s = 235;
	{8'd41,8'd195} : s = 236;
	{8'd41,8'd196} : s = 237;
	{8'd41,8'd197} : s = 238;
	{8'd41,8'd198} : s = 239;
	{8'd41,8'd199} : s = 240;
	{8'd41,8'd200} : s = 241;
	{8'd41,8'd201} : s = 242;
	{8'd41,8'd202} : s = 243;
	{8'd41,8'd203} : s = 244;
	{8'd41,8'd204} : s = 245;
	{8'd41,8'd205} : s = 246;
	{8'd41,8'd206} : s = 247;
	{8'd41,8'd207} : s = 248;
	{8'd41,8'd208} : s = 249;
	{8'd41,8'd209} : s = 250;
	{8'd41,8'd210} : s = 251;
	{8'd41,8'd211} : s = 252;
	{8'd41,8'd212} : s = 253;
	{8'd41,8'd213} : s = 254;
	{8'd41,8'd214} : s = 255;
	{8'd41,8'd215} : s = 256;
	{8'd41,8'd216} : s = 257;
	{8'd41,8'd217} : s = 258;
	{8'd41,8'd218} : s = 259;
	{8'd41,8'd219} : s = 260;
	{8'd41,8'd220} : s = 261;
	{8'd41,8'd221} : s = 262;
	{8'd41,8'd222} : s = 263;
	{8'd41,8'd223} : s = 264;
	{8'd41,8'd224} : s = 265;
	{8'd41,8'd225} : s = 266;
	{8'd41,8'd226} : s = 267;
	{8'd41,8'd227} : s = 268;
	{8'd41,8'd228} : s = 269;
	{8'd41,8'd229} : s = 270;
	{8'd41,8'd230} : s = 271;
	{8'd41,8'd231} : s = 272;
	{8'd41,8'd232} : s = 273;
	{8'd41,8'd233} : s = 274;
	{8'd41,8'd234} : s = 275;
	{8'd41,8'd235} : s = 276;
	{8'd41,8'd236} : s = 277;
	{8'd41,8'd237} : s = 278;
	{8'd41,8'd238} : s = 279;
	{8'd41,8'd239} : s = 280;
	{8'd41,8'd240} : s = 281;
	{8'd41,8'd241} : s = 282;
	{8'd41,8'd242} : s = 283;
	{8'd41,8'd243} : s = 284;
	{8'd41,8'd244} : s = 285;
	{8'd41,8'd245} : s = 286;
	{8'd41,8'd246} : s = 287;
	{8'd41,8'd247} : s = 288;
	{8'd41,8'd248} : s = 289;
	{8'd41,8'd249} : s = 290;
	{8'd41,8'd250} : s = 291;
	{8'd41,8'd251} : s = 292;
	{8'd41,8'd252} : s = 293;
	{8'd41,8'd253} : s = 294;
	{8'd41,8'd254} : s = 295;
	{8'd41,8'd255} : s = 296;
	{8'd42,8'd0} : s = 42;
	{8'd42,8'd1} : s = 43;
	{8'd42,8'd2} : s = 44;
	{8'd42,8'd3} : s = 45;
	{8'd42,8'd4} : s = 46;
	{8'd42,8'd5} : s = 47;
	{8'd42,8'd6} : s = 48;
	{8'd42,8'd7} : s = 49;
	{8'd42,8'd8} : s = 50;
	{8'd42,8'd9} : s = 51;
	{8'd42,8'd10} : s = 52;
	{8'd42,8'd11} : s = 53;
	{8'd42,8'd12} : s = 54;
	{8'd42,8'd13} : s = 55;
	{8'd42,8'd14} : s = 56;
	{8'd42,8'd15} : s = 57;
	{8'd42,8'd16} : s = 58;
	{8'd42,8'd17} : s = 59;
	{8'd42,8'd18} : s = 60;
	{8'd42,8'd19} : s = 61;
	{8'd42,8'd20} : s = 62;
	{8'd42,8'd21} : s = 63;
	{8'd42,8'd22} : s = 64;
	{8'd42,8'd23} : s = 65;
	{8'd42,8'd24} : s = 66;
	{8'd42,8'd25} : s = 67;
	{8'd42,8'd26} : s = 68;
	{8'd42,8'd27} : s = 69;
	{8'd42,8'd28} : s = 70;
	{8'd42,8'd29} : s = 71;
	{8'd42,8'd30} : s = 72;
	{8'd42,8'd31} : s = 73;
	{8'd42,8'd32} : s = 74;
	{8'd42,8'd33} : s = 75;
	{8'd42,8'd34} : s = 76;
	{8'd42,8'd35} : s = 77;
	{8'd42,8'd36} : s = 78;
	{8'd42,8'd37} : s = 79;
	{8'd42,8'd38} : s = 80;
	{8'd42,8'd39} : s = 81;
	{8'd42,8'd40} : s = 82;
	{8'd42,8'd41} : s = 83;
	{8'd42,8'd42} : s = 84;
	{8'd42,8'd43} : s = 85;
	{8'd42,8'd44} : s = 86;
	{8'd42,8'd45} : s = 87;
	{8'd42,8'd46} : s = 88;
	{8'd42,8'd47} : s = 89;
	{8'd42,8'd48} : s = 90;
	{8'd42,8'd49} : s = 91;
	{8'd42,8'd50} : s = 92;
	{8'd42,8'd51} : s = 93;
	{8'd42,8'd52} : s = 94;
	{8'd42,8'd53} : s = 95;
	{8'd42,8'd54} : s = 96;
	{8'd42,8'd55} : s = 97;
	{8'd42,8'd56} : s = 98;
	{8'd42,8'd57} : s = 99;
	{8'd42,8'd58} : s = 100;
	{8'd42,8'd59} : s = 101;
	{8'd42,8'd60} : s = 102;
	{8'd42,8'd61} : s = 103;
	{8'd42,8'd62} : s = 104;
	{8'd42,8'd63} : s = 105;
	{8'd42,8'd64} : s = 106;
	{8'd42,8'd65} : s = 107;
	{8'd42,8'd66} : s = 108;
	{8'd42,8'd67} : s = 109;
	{8'd42,8'd68} : s = 110;
	{8'd42,8'd69} : s = 111;
	{8'd42,8'd70} : s = 112;
	{8'd42,8'd71} : s = 113;
	{8'd42,8'd72} : s = 114;
	{8'd42,8'd73} : s = 115;
	{8'd42,8'd74} : s = 116;
	{8'd42,8'd75} : s = 117;
	{8'd42,8'd76} : s = 118;
	{8'd42,8'd77} : s = 119;
	{8'd42,8'd78} : s = 120;
	{8'd42,8'd79} : s = 121;
	{8'd42,8'd80} : s = 122;
	{8'd42,8'd81} : s = 123;
	{8'd42,8'd82} : s = 124;
	{8'd42,8'd83} : s = 125;
	{8'd42,8'd84} : s = 126;
	{8'd42,8'd85} : s = 127;
	{8'd42,8'd86} : s = 128;
	{8'd42,8'd87} : s = 129;
	{8'd42,8'd88} : s = 130;
	{8'd42,8'd89} : s = 131;
	{8'd42,8'd90} : s = 132;
	{8'd42,8'd91} : s = 133;
	{8'd42,8'd92} : s = 134;
	{8'd42,8'd93} : s = 135;
	{8'd42,8'd94} : s = 136;
	{8'd42,8'd95} : s = 137;
	{8'd42,8'd96} : s = 138;
	{8'd42,8'd97} : s = 139;
	{8'd42,8'd98} : s = 140;
	{8'd42,8'd99} : s = 141;
	{8'd42,8'd100} : s = 142;
	{8'd42,8'd101} : s = 143;
	{8'd42,8'd102} : s = 144;
	{8'd42,8'd103} : s = 145;
	{8'd42,8'd104} : s = 146;
	{8'd42,8'd105} : s = 147;
	{8'd42,8'd106} : s = 148;
	{8'd42,8'd107} : s = 149;
	{8'd42,8'd108} : s = 150;
	{8'd42,8'd109} : s = 151;
	{8'd42,8'd110} : s = 152;
	{8'd42,8'd111} : s = 153;
	{8'd42,8'd112} : s = 154;
	{8'd42,8'd113} : s = 155;
	{8'd42,8'd114} : s = 156;
	{8'd42,8'd115} : s = 157;
	{8'd42,8'd116} : s = 158;
	{8'd42,8'd117} : s = 159;
	{8'd42,8'd118} : s = 160;
	{8'd42,8'd119} : s = 161;
	{8'd42,8'd120} : s = 162;
	{8'd42,8'd121} : s = 163;
	{8'd42,8'd122} : s = 164;
	{8'd42,8'd123} : s = 165;
	{8'd42,8'd124} : s = 166;
	{8'd42,8'd125} : s = 167;
	{8'd42,8'd126} : s = 168;
	{8'd42,8'd127} : s = 169;
	{8'd42,8'd128} : s = 170;
	{8'd42,8'd129} : s = 171;
	{8'd42,8'd130} : s = 172;
	{8'd42,8'd131} : s = 173;
	{8'd42,8'd132} : s = 174;
	{8'd42,8'd133} : s = 175;
	{8'd42,8'd134} : s = 176;
	{8'd42,8'd135} : s = 177;
	{8'd42,8'd136} : s = 178;
	{8'd42,8'd137} : s = 179;
	{8'd42,8'd138} : s = 180;
	{8'd42,8'd139} : s = 181;
	{8'd42,8'd140} : s = 182;
	{8'd42,8'd141} : s = 183;
	{8'd42,8'd142} : s = 184;
	{8'd42,8'd143} : s = 185;
	{8'd42,8'd144} : s = 186;
	{8'd42,8'd145} : s = 187;
	{8'd42,8'd146} : s = 188;
	{8'd42,8'd147} : s = 189;
	{8'd42,8'd148} : s = 190;
	{8'd42,8'd149} : s = 191;
	{8'd42,8'd150} : s = 192;
	{8'd42,8'd151} : s = 193;
	{8'd42,8'd152} : s = 194;
	{8'd42,8'd153} : s = 195;
	{8'd42,8'd154} : s = 196;
	{8'd42,8'd155} : s = 197;
	{8'd42,8'd156} : s = 198;
	{8'd42,8'd157} : s = 199;
	{8'd42,8'd158} : s = 200;
	{8'd42,8'd159} : s = 201;
	{8'd42,8'd160} : s = 202;
	{8'd42,8'd161} : s = 203;
	{8'd42,8'd162} : s = 204;
	{8'd42,8'd163} : s = 205;
	{8'd42,8'd164} : s = 206;
	{8'd42,8'd165} : s = 207;
	{8'd42,8'd166} : s = 208;
	{8'd42,8'd167} : s = 209;
	{8'd42,8'd168} : s = 210;
	{8'd42,8'd169} : s = 211;
	{8'd42,8'd170} : s = 212;
	{8'd42,8'd171} : s = 213;
	{8'd42,8'd172} : s = 214;
	{8'd42,8'd173} : s = 215;
	{8'd42,8'd174} : s = 216;
	{8'd42,8'd175} : s = 217;
	{8'd42,8'd176} : s = 218;
	{8'd42,8'd177} : s = 219;
	{8'd42,8'd178} : s = 220;
	{8'd42,8'd179} : s = 221;
	{8'd42,8'd180} : s = 222;
	{8'd42,8'd181} : s = 223;
	{8'd42,8'd182} : s = 224;
	{8'd42,8'd183} : s = 225;
	{8'd42,8'd184} : s = 226;
	{8'd42,8'd185} : s = 227;
	{8'd42,8'd186} : s = 228;
	{8'd42,8'd187} : s = 229;
	{8'd42,8'd188} : s = 230;
	{8'd42,8'd189} : s = 231;
	{8'd42,8'd190} : s = 232;
	{8'd42,8'd191} : s = 233;
	{8'd42,8'd192} : s = 234;
	{8'd42,8'd193} : s = 235;
	{8'd42,8'd194} : s = 236;
	{8'd42,8'd195} : s = 237;
	{8'd42,8'd196} : s = 238;
	{8'd42,8'd197} : s = 239;
	{8'd42,8'd198} : s = 240;
	{8'd42,8'd199} : s = 241;
	{8'd42,8'd200} : s = 242;
	{8'd42,8'd201} : s = 243;
	{8'd42,8'd202} : s = 244;
	{8'd42,8'd203} : s = 245;
	{8'd42,8'd204} : s = 246;
	{8'd42,8'd205} : s = 247;
	{8'd42,8'd206} : s = 248;
	{8'd42,8'd207} : s = 249;
	{8'd42,8'd208} : s = 250;
	{8'd42,8'd209} : s = 251;
	{8'd42,8'd210} : s = 252;
	{8'd42,8'd211} : s = 253;
	{8'd42,8'd212} : s = 254;
	{8'd42,8'd213} : s = 255;
	{8'd42,8'd214} : s = 256;
	{8'd42,8'd215} : s = 257;
	{8'd42,8'd216} : s = 258;
	{8'd42,8'd217} : s = 259;
	{8'd42,8'd218} : s = 260;
	{8'd42,8'd219} : s = 261;
	{8'd42,8'd220} : s = 262;
	{8'd42,8'd221} : s = 263;
	{8'd42,8'd222} : s = 264;
	{8'd42,8'd223} : s = 265;
	{8'd42,8'd224} : s = 266;
	{8'd42,8'd225} : s = 267;
	{8'd42,8'd226} : s = 268;
	{8'd42,8'd227} : s = 269;
	{8'd42,8'd228} : s = 270;
	{8'd42,8'd229} : s = 271;
	{8'd42,8'd230} : s = 272;
	{8'd42,8'd231} : s = 273;
	{8'd42,8'd232} : s = 274;
	{8'd42,8'd233} : s = 275;
	{8'd42,8'd234} : s = 276;
	{8'd42,8'd235} : s = 277;
	{8'd42,8'd236} : s = 278;
	{8'd42,8'd237} : s = 279;
	{8'd42,8'd238} : s = 280;
	{8'd42,8'd239} : s = 281;
	{8'd42,8'd240} : s = 282;
	{8'd42,8'd241} : s = 283;
	{8'd42,8'd242} : s = 284;
	{8'd42,8'd243} : s = 285;
	{8'd42,8'd244} : s = 286;
	{8'd42,8'd245} : s = 287;
	{8'd42,8'd246} : s = 288;
	{8'd42,8'd247} : s = 289;
	{8'd42,8'd248} : s = 290;
	{8'd42,8'd249} : s = 291;
	{8'd42,8'd250} : s = 292;
	{8'd42,8'd251} : s = 293;
	{8'd42,8'd252} : s = 294;
	{8'd42,8'd253} : s = 295;
	{8'd42,8'd254} : s = 296;
	{8'd42,8'd255} : s = 297;
	{8'd43,8'd0} : s = 43;
	{8'd43,8'd1} : s = 44;
	{8'd43,8'd2} : s = 45;
	{8'd43,8'd3} : s = 46;
	{8'd43,8'd4} : s = 47;
	{8'd43,8'd5} : s = 48;
	{8'd43,8'd6} : s = 49;
	{8'd43,8'd7} : s = 50;
	{8'd43,8'd8} : s = 51;
	{8'd43,8'd9} : s = 52;
	{8'd43,8'd10} : s = 53;
	{8'd43,8'd11} : s = 54;
	{8'd43,8'd12} : s = 55;
	{8'd43,8'd13} : s = 56;
	{8'd43,8'd14} : s = 57;
	{8'd43,8'd15} : s = 58;
	{8'd43,8'd16} : s = 59;
	{8'd43,8'd17} : s = 60;
	{8'd43,8'd18} : s = 61;
	{8'd43,8'd19} : s = 62;
	{8'd43,8'd20} : s = 63;
	{8'd43,8'd21} : s = 64;
	{8'd43,8'd22} : s = 65;
	{8'd43,8'd23} : s = 66;
	{8'd43,8'd24} : s = 67;
	{8'd43,8'd25} : s = 68;
	{8'd43,8'd26} : s = 69;
	{8'd43,8'd27} : s = 70;
	{8'd43,8'd28} : s = 71;
	{8'd43,8'd29} : s = 72;
	{8'd43,8'd30} : s = 73;
	{8'd43,8'd31} : s = 74;
	{8'd43,8'd32} : s = 75;
	{8'd43,8'd33} : s = 76;
	{8'd43,8'd34} : s = 77;
	{8'd43,8'd35} : s = 78;
	{8'd43,8'd36} : s = 79;
	{8'd43,8'd37} : s = 80;
	{8'd43,8'd38} : s = 81;
	{8'd43,8'd39} : s = 82;
	{8'd43,8'd40} : s = 83;
	{8'd43,8'd41} : s = 84;
	{8'd43,8'd42} : s = 85;
	{8'd43,8'd43} : s = 86;
	{8'd43,8'd44} : s = 87;
	{8'd43,8'd45} : s = 88;
	{8'd43,8'd46} : s = 89;
	{8'd43,8'd47} : s = 90;
	{8'd43,8'd48} : s = 91;
	{8'd43,8'd49} : s = 92;
	{8'd43,8'd50} : s = 93;
	{8'd43,8'd51} : s = 94;
	{8'd43,8'd52} : s = 95;
	{8'd43,8'd53} : s = 96;
	{8'd43,8'd54} : s = 97;
	{8'd43,8'd55} : s = 98;
	{8'd43,8'd56} : s = 99;
	{8'd43,8'd57} : s = 100;
	{8'd43,8'd58} : s = 101;
	{8'd43,8'd59} : s = 102;
	{8'd43,8'd60} : s = 103;
	{8'd43,8'd61} : s = 104;
	{8'd43,8'd62} : s = 105;
	{8'd43,8'd63} : s = 106;
	{8'd43,8'd64} : s = 107;
	{8'd43,8'd65} : s = 108;
	{8'd43,8'd66} : s = 109;
	{8'd43,8'd67} : s = 110;
	{8'd43,8'd68} : s = 111;
	{8'd43,8'd69} : s = 112;
	{8'd43,8'd70} : s = 113;
	{8'd43,8'd71} : s = 114;
	{8'd43,8'd72} : s = 115;
	{8'd43,8'd73} : s = 116;
	{8'd43,8'd74} : s = 117;
	{8'd43,8'd75} : s = 118;
	{8'd43,8'd76} : s = 119;
	{8'd43,8'd77} : s = 120;
	{8'd43,8'd78} : s = 121;
	{8'd43,8'd79} : s = 122;
	{8'd43,8'd80} : s = 123;
	{8'd43,8'd81} : s = 124;
	{8'd43,8'd82} : s = 125;
	{8'd43,8'd83} : s = 126;
	{8'd43,8'd84} : s = 127;
	{8'd43,8'd85} : s = 128;
	{8'd43,8'd86} : s = 129;
	{8'd43,8'd87} : s = 130;
	{8'd43,8'd88} : s = 131;
	{8'd43,8'd89} : s = 132;
	{8'd43,8'd90} : s = 133;
	{8'd43,8'd91} : s = 134;
	{8'd43,8'd92} : s = 135;
	{8'd43,8'd93} : s = 136;
	{8'd43,8'd94} : s = 137;
	{8'd43,8'd95} : s = 138;
	{8'd43,8'd96} : s = 139;
	{8'd43,8'd97} : s = 140;
	{8'd43,8'd98} : s = 141;
	{8'd43,8'd99} : s = 142;
	{8'd43,8'd100} : s = 143;
	{8'd43,8'd101} : s = 144;
	{8'd43,8'd102} : s = 145;
	{8'd43,8'd103} : s = 146;
	{8'd43,8'd104} : s = 147;
	{8'd43,8'd105} : s = 148;
	{8'd43,8'd106} : s = 149;
	{8'd43,8'd107} : s = 150;
	{8'd43,8'd108} : s = 151;
	{8'd43,8'd109} : s = 152;
	{8'd43,8'd110} : s = 153;
	{8'd43,8'd111} : s = 154;
	{8'd43,8'd112} : s = 155;
	{8'd43,8'd113} : s = 156;
	{8'd43,8'd114} : s = 157;
	{8'd43,8'd115} : s = 158;
	{8'd43,8'd116} : s = 159;
	{8'd43,8'd117} : s = 160;
	{8'd43,8'd118} : s = 161;
	{8'd43,8'd119} : s = 162;
	{8'd43,8'd120} : s = 163;
	{8'd43,8'd121} : s = 164;
	{8'd43,8'd122} : s = 165;
	{8'd43,8'd123} : s = 166;
	{8'd43,8'd124} : s = 167;
	{8'd43,8'd125} : s = 168;
	{8'd43,8'd126} : s = 169;
	{8'd43,8'd127} : s = 170;
	{8'd43,8'd128} : s = 171;
	{8'd43,8'd129} : s = 172;
	{8'd43,8'd130} : s = 173;
	{8'd43,8'd131} : s = 174;
	{8'd43,8'd132} : s = 175;
	{8'd43,8'd133} : s = 176;
	{8'd43,8'd134} : s = 177;
	{8'd43,8'd135} : s = 178;
	{8'd43,8'd136} : s = 179;
	{8'd43,8'd137} : s = 180;
	{8'd43,8'd138} : s = 181;
	{8'd43,8'd139} : s = 182;
	{8'd43,8'd140} : s = 183;
	{8'd43,8'd141} : s = 184;
	{8'd43,8'd142} : s = 185;
	{8'd43,8'd143} : s = 186;
	{8'd43,8'd144} : s = 187;
	{8'd43,8'd145} : s = 188;
	{8'd43,8'd146} : s = 189;
	{8'd43,8'd147} : s = 190;
	{8'd43,8'd148} : s = 191;
	{8'd43,8'd149} : s = 192;
	{8'd43,8'd150} : s = 193;
	{8'd43,8'd151} : s = 194;
	{8'd43,8'd152} : s = 195;
	{8'd43,8'd153} : s = 196;
	{8'd43,8'd154} : s = 197;
	{8'd43,8'd155} : s = 198;
	{8'd43,8'd156} : s = 199;
	{8'd43,8'd157} : s = 200;
	{8'd43,8'd158} : s = 201;
	{8'd43,8'd159} : s = 202;
	{8'd43,8'd160} : s = 203;
	{8'd43,8'd161} : s = 204;
	{8'd43,8'd162} : s = 205;
	{8'd43,8'd163} : s = 206;
	{8'd43,8'd164} : s = 207;
	{8'd43,8'd165} : s = 208;
	{8'd43,8'd166} : s = 209;
	{8'd43,8'd167} : s = 210;
	{8'd43,8'd168} : s = 211;
	{8'd43,8'd169} : s = 212;
	{8'd43,8'd170} : s = 213;
	{8'd43,8'd171} : s = 214;
	{8'd43,8'd172} : s = 215;
	{8'd43,8'd173} : s = 216;
	{8'd43,8'd174} : s = 217;
	{8'd43,8'd175} : s = 218;
	{8'd43,8'd176} : s = 219;
	{8'd43,8'd177} : s = 220;
	{8'd43,8'd178} : s = 221;
	{8'd43,8'd179} : s = 222;
	{8'd43,8'd180} : s = 223;
	{8'd43,8'd181} : s = 224;
	{8'd43,8'd182} : s = 225;
	{8'd43,8'd183} : s = 226;
	{8'd43,8'd184} : s = 227;
	{8'd43,8'd185} : s = 228;
	{8'd43,8'd186} : s = 229;
	{8'd43,8'd187} : s = 230;
	{8'd43,8'd188} : s = 231;
	{8'd43,8'd189} : s = 232;
	{8'd43,8'd190} : s = 233;
	{8'd43,8'd191} : s = 234;
	{8'd43,8'd192} : s = 235;
	{8'd43,8'd193} : s = 236;
	{8'd43,8'd194} : s = 237;
	{8'd43,8'd195} : s = 238;
	{8'd43,8'd196} : s = 239;
	{8'd43,8'd197} : s = 240;
	{8'd43,8'd198} : s = 241;
	{8'd43,8'd199} : s = 242;
	{8'd43,8'd200} : s = 243;
	{8'd43,8'd201} : s = 244;
	{8'd43,8'd202} : s = 245;
	{8'd43,8'd203} : s = 246;
	{8'd43,8'd204} : s = 247;
	{8'd43,8'd205} : s = 248;
	{8'd43,8'd206} : s = 249;
	{8'd43,8'd207} : s = 250;
	{8'd43,8'd208} : s = 251;
	{8'd43,8'd209} : s = 252;
	{8'd43,8'd210} : s = 253;
	{8'd43,8'd211} : s = 254;
	{8'd43,8'd212} : s = 255;
	{8'd43,8'd213} : s = 256;
	{8'd43,8'd214} : s = 257;
	{8'd43,8'd215} : s = 258;
	{8'd43,8'd216} : s = 259;
	{8'd43,8'd217} : s = 260;
	{8'd43,8'd218} : s = 261;
	{8'd43,8'd219} : s = 262;
	{8'd43,8'd220} : s = 263;
	{8'd43,8'd221} : s = 264;
	{8'd43,8'd222} : s = 265;
	{8'd43,8'd223} : s = 266;
	{8'd43,8'd224} : s = 267;
	{8'd43,8'd225} : s = 268;
	{8'd43,8'd226} : s = 269;
	{8'd43,8'd227} : s = 270;
	{8'd43,8'd228} : s = 271;
	{8'd43,8'd229} : s = 272;
	{8'd43,8'd230} : s = 273;
	{8'd43,8'd231} : s = 274;
	{8'd43,8'd232} : s = 275;
	{8'd43,8'd233} : s = 276;
	{8'd43,8'd234} : s = 277;
	{8'd43,8'd235} : s = 278;
	{8'd43,8'd236} : s = 279;
	{8'd43,8'd237} : s = 280;
	{8'd43,8'd238} : s = 281;
	{8'd43,8'd239} : s = 282;
	{8'd43,8'd240} : s = 283;
	{8'd43,8'd241} : s = 284;
	{8'd43,8'd242} : s = 285;
	{8'd43,8'd243} : s = 286;
	{8'd43,8'd244} : s = 287;
	{8'd43,8'd245} : s = 288;
	{8'd43,8'd246} : s = 289;
	{8'd43,8'd247} : s = 290;
	{8'd43,8'd248} : s = 291;
	{8'd43,8'd249} : s = 292;
	{8'd43,8'd250} : s = 293;
	{8'd43,8'd251} : s = 294;
	{8'd43,8'd252} : s = 295;
	{8'd43,8'd253} : s = 296;
	{8'd43,8'd254} : s = 297;
	{8'd43,8'd255} : s = 298;
	{8'd44,8'd0} : s = 44;
	{8'd44,8'd1} : s = 45;
	{8'd44,8'd2} : s = 46;
	{8'd44,8'd3} : s = 47;
	{8'd44,8'd4} : s = 48;
	{8'd44,8'd5} : s = 49;
	{8'd44,8'd6} : s = 50;
	{8'd44,8'd7} : s = 51;
	{8'd44,8'd8} : s = 52;
	{8'd44,8'd9} : s = 53;
	{8'd44,8'd10} : s = 54;
	{8'd44,8'd11} : s = 55;
	{8'd44,8'd12} : s = 56;
	{8'd44,8'd13} : s = 57;
	{8'd44,8'd14} : s = 58;
	{8'd44,8'd15} : s = 59;
	{8'd44,8'd16} : s = 60;
	{8'd44,8'd17} : s = 61;
	{8'd44,8'd18} : s = 62;
	{8'd44,8'd19} : s = 63;
	{8'd44,8'd20} : s = 64;
	{8'd44,8'd21} : s = 65;
	{8'd44,8'd22} : s = 66;
	{8'd44,8'd23} : s = 67;
	{8'd44,8'd24} : s = 68;
	{8'd44,8'd25} : s = 69;
	{8'd44,8'd26} : s = 70;
	{8'd44,8'd27} : s = 71;
	{8'd44,8'd28} : s = 72;
	{8'd44,8'd29} : s = 73;
	{8'd44,8'd30} : s = 74;
	{8'd44,8'd31} : s = 75;
	{8'd44,8'd32} : s = 76;
	{8'd44,8'd33} : s = 77;
	{8'd44,8'd34} : s = 78;
	{8'd44,8'd35} : s = 79;
	{8'd44,8'd36} : s = 80;
	{8'd44,8'd37} : s = 81;
	{8'd44,8'd38} : s = 82;
	{8'd44,8'd39} : s = 83;
	{8'd44,8'd40} : s = 84;
	{8'd44,8'd41} : s = 85;
	{8'd44,8'd42} : s = 86;
	{8'd44,8'd43} : s = 87;
	{8'd44,8'd44} : s = 88;
	{8'd44,8'd45} : s = 89;
	{8'd44,8'd46} : s = 90;
	{8'd44,8'd47} : s = 91;
	{8'd44,8'd48} : s = 92;
	{8'd44,8'd49} : s = 93;
	{8'd44,8'd50} : s = 94;
	{8'd44,8'd51} : s = 95;
	{8'd44,8'd52} : s = 96;
	{8'd44,8'd53} : s = 97;
	{8'd44,8'd54} : s = 98;
	{8'd44,8'd55} : s = 99;
	{8'd44,8'd56} : s = 100;
	{8'd44,8'd57} : s = 101;
	{8'd44,8'd58} : s = 102;
	{8'd44,8'd59} : s = 103;
	{8'd44,8'd60} : s = 104;
	{8'd44,8'd61} : s = 105;
	{8'd44,8'd62} : s = 106;
	{8'd44,8'd63} : s = 107;
	{8'd44,8'd64} : s = 108;
	{8'd44,8'd65} : s = 109;
	{8'd44,8'd66} : s = 110;
	{8'd44,8'd67} : s = 111;
	{8'd44,8'd68} : s = 112;
	{8'd44,8'd69} : s = 113;
	{8'd44,8'd70} : s = 114;
	{8'd44,8'd71} : s = 115;
	{8'd44,8'd72} : s = 116;
	{8'd44,8'd73} : s = 117;
	{8'd44,8'd74} : s = 118;
	{8'd44,8'd75} : s = 119;
	{8'd44,8'd76} : s = 120;
	{8'd44,8'd77} : s = 121;
	{8'd44,8'd78} : s = 122;
	{8'd44,8'd79} : s = 123;
	{8'd44,8'd80} : s = 124;
	{8'd44,8'd81} : s = 125;
	{8'd44,8'd82} : s = 126;
	{8'd44,8'd83} : s = 127;
	{8'd44,8'd84} : s = 128;
	{8'd44,8'd85} : s = 129;
	{8'd44,8'd86} : s = 130;
	{8'd44,8'd87} : s = 131;
	{8'd44,8'd88} : s = 132;
	{8'd44,8'd89} : s = 133;
	{8'd44,8'd90} : s = 134;
	{8'd44,8'd91} : s = 135;
	{8'd44,8'd92} : s = 136;
	{8'd44,8'd93} : s = 137;
	{8'd44,8'd94} : s = 138;
	{8'd44,8'd95} : s = 139;
	{8'd44,8'd96} : s = 140;
	{8'd44,8'd97} : s = 141;
	{8'd44,8'd98} : s = 142;
	{8'd44,8'd99} : s = 143;
	{8'd44,8'd100} : s = 144;
	{8'd44,8'd101} : s = 145;
	{8'd44,8'd102} : s = 146;
	{8'd44,8'd103} : s = 147;
	{8'd44,8'd104} : s = 148;
	{8'd44,8'd105} : s = 149;
	{8'd44,8'd106} : s = 150;
	{8'd44,8'd107} : s = 151;
	{8'd44,8'd108} : s = 152;
	{8'd44,8'd109} : s = 153;
	{8'd44,8'd110} : s = 154;
	{8'd44,8'd111} : s = 155;
	{8'd44,8'd112} : s = 156;
	{8'd44,8'd113} : s = 157;
	{8'd44,8'd114} : s = 158;
	{8'd44,8'd115} : s = 159;
	{8'd44,8'd116} : s = 160;
	{8'd44,8'd117} : s = 161;
	{8'd44,8'd118} : s = 162;
	{8'd44,8'd119} : s = 163;
	{8'd44,8'd120} : s = 164;
	{8'd44,8'd121} : s = 165;
	{8'd44,8'd122} : s = 166;
	{8'd44,8'd123} : s = 167;
	{8'd44,8'd124} : s = 168;
	{8'd44,8'd125} : s = 169;
	{8'd44,8'd126} : s = 170;
	{8'd44,8'd127} : s = 171;
	{8'd44,8'd128} : s = 172;
	{8'd44,8'd129} : s = 173;
	{8'd44,8'd130} : s = 174;
	{8'd44,8'd131} : s = 175;
	{8'd44,8'd132} : s = 176;
	{8'd44,8'd133} : s = 177;
	{8'd44,8'd134} : s = 178;
	{8'd44,8'd135} : s = 179;
	{8'd44,8'd136} : s = 180;
	{8'd44,8'd137} : s = 181;
	{8'd44,8'd138} : s = 182;
	{8'd44,8'd139} : s = 183;
	{8'd44,8'd140} : s = 184;
	{8'd44,8'd141} : s = 185;
	{8'd44,8'd142} : s = 186;
	{8'd44,8'd143} : s = 187;
	{8'd44,8'd144} : s = 188;
	{8'd44,8'd145} : s = 189;
	{8'd44,8'd146} : s = 190;
	{8'd44,8'd147} : s = 191;
	{8'd44,8'd148} : s = 192;
	{8'd44,8'd149} : s = 193;
	{8'd44,8'd150} : s = 194;
	{8'd44,8'd151} : s = 195;
	{8'd44,8'd152} : s = 196;
	{8'd44,8'd153} : s = 197;
	{8'd44,8'd154} : s = 198;
	{8'd44,8'd155} : s = 199;
	{8'd44,8'd156} : s = 200;
	{8'd44,8'd157} : s = 201;
	{8'd44,8'd158} : s = 202;
	{8'd44,8'd159} : s = 203;
	{8'd44,8'd160} : s = 204;
	{8'd44,8'd161} : s = 205;
	{8'd44,8'd162} : s = 206;
	{8'd44,8'd163} : s = 207;
	{8'd44,8'd164} : s = 208;
	{8'd44,8'd165} : s = 209;
	{8'd44,8'd166} : s = 210;
	{8'd44,8'd167} : s = 211;
	{8'd44,8'd168} : s = 212;
	{8'd44,8'd169} : s = 213;
	{8'd44,8'd170} : s = 214;
	{8'd44,8'd171} : s = 215;
	{8'd44,8'd172} : s = 216;
	{8'd44,8'd173} : s = 217;
	{8'd44,8'd174} : s = 218;
	{8'd44,8'd175} : s = 219;
	{8'd44,8'd176} : s = 220;
	{8'd44,8'd177} : s = 221;
	{8'd44,8'd178} : s = 222;
	{8'd44,8'd179} : s = 223;
	{8'd44,8'd180} : s = 224;
	{8'd44,8'd181} : s = 225;
	{8'd44,8'd182} : s = 226;
	{8'd44,8'd183} : s = 227;
	{8'd44,8'd184} : s = 228;
	{8'd44,8'd185} : s = 229;
	{8'd44,8'd186} : s = 230;
	{8'd44,8'd187} : s = 231;
	{8'd44,8'd188} : s = 232;
	{8'd44,8'd189} : s = 233;
	{8'd44,8'd190} : s = 234;
	{8'd44,8'd191} : s = 235;
	{8'd44,8'd192} : s = 236;
	{8'd44,8'd193} : s = 237;
	{8'd44,8'd194} : s = 238;
	{8'd44,8'd195} : s = 239;
	{8'd44,8'd196} : s = 240;
	{8'd44,8'd197} : s = 241;
	{8'd44,8'd198} : s = 242;
	{8'd44,8'd199} : s = 243;
	{8'd44,8'd200} : s = 244;
	{8'd44,8'd201} : s = 245;
	{8'd44,8'd202} : s = 246;
	{8'd44,8'd203} : s = 247;
	{8'd44,8'd204} : s = 248;
	{8'd44,8'd205} : s = 249;
	{8'd44,8'd206} : s = 250;
	{8'd44,8'd207} : s = 251;
	{8'd44,8'd208} : s = 252;
	{8'd44,8'd209} : s = 253;
	{8'd44,8'd210} : s = 254;
	{8'd44,8'd211} : s = 255;
	{8'd44,8'd212} : s = 256;
	{8'd44,8'd213} : s = 257;
	{8'd44,8'd214} : s = 258;
	{8'd44,8'd215} : s = 259;
	{8'd44,8'd216} : s = 260;
	{8'd44,8'd217} : s = 261;
	{8'd44,8'd218} : s = 262;
	{8'd44,8'd219} : s = 263;
	{8'd44,8'd220} : s = 264;
	{8'd44,8'd221} : s = 265;
	{8'd44,8'd222} : s = 266;
	{8'd44,8'd223} : s = 267;
	{8'd44,8'd224} : s = 268;
	{8'd44,8'd225} : s = 269;
	{8'd44,8'd226} : s = 270;
	{8'd44,8'd227} : s = 271;
	{8'd44,8'd228} : s = 272;
	{8'd44,8'd229} : s = 273;
	{8'd44,8'd230} : s = 274;
	{8'd44,8'd231} : s = 275;
	{8'd44,8'd232} : s = 276;
	{8'd44,8'd233} : s = 277;
	{8'd44,8'd234} : s = 278;
	{8'd44,8'd235} : s = 279;
	{8'd44,8'd236} : s = 280;
	{8'd44,8'd237} : s = 281;
	{8'd44,8'd238} : s = 282;
	{8'd44,8'd239} : s = 283;
	{8'd44,8'd240} : s = 284;
	{8'd44,8'd241} : s = 285;
	{8'd44,8'd242} : s = 286;
	{8'd44,8'd243} : s = 287;
	{8'd44,8'd244} : s = 288;
	{8'd44,8'd245} : s = 289;
	{8'd44,8'd246} : s = 290;
	{8'd44,8'd247} : s = 291;
	{8'd44,8'd248} : s = 292;
	{8'd44,8'd249} : s = 293;
	{8'd44,8'd250} : s = 294;
	{8'd44,8'd251} : s = 295;
	{8'd44,8'd252} : s = 296;
	{8'd44,8'd253} : s = 297;
	{8'd44,8'd254} : s = 298;
	{8'd44,8'd255} : s = 299;
	{8'd45,8'd0} : s = 45;
	{8'd45,8'd1} : s = 46;
	{8'd45,8'd2} : s = 47;
	{8'd45,8'd3} : s = 48;
	{8'd45,8'd4} : s = 49;
	{8'd45,8'd5} : s = 50;
	{8'd45,8'd6} : s = 51;
	{8'd45,8'd7} : s = 52;
	{8'd45,8'd8} : s = 53;
	{8'd45,8'd9} : s = 54;
	{8'd45,8'd10} : s = 55;
	{8'd45,8'd11} : s = 56;
	{8'd45,8'd12} : s = 57;
	{8'd45,8'd13} : s = 58;
	{8'd45,8'd14} : s = 59;
	{8'd45,8'd15} : s = 60;
	{8'd45,8'd16} : s = 61;
	{8'd45,8'd17} : s = 62;
	{8'd45,8'd18} : s = 63;
	{8'd45,8'd19} : s = 64;
	{8'd45,8'd20} : s = 65;
	{8'd45,8'd21} : s = 66;
	{8'd45,8'd22} : s = 67;
	{8'd45,8'd23} : s = 68;
	{8'd45,8'd24} : s = 69;
	{8'd45,8'd25} : s = 70;
	{8'd45,8'd26} : s = 71;
	{8'd45,8'd27} : s = 72;
	{8'd45,8'd28} : s = 73;
	{8'd45,8'd29} : s = 74;
	{8'd45,8'd30} : s = 75;
	{8'd45,8'd31} : s = 76;
	{8'd45,8'd32} : s = 77;
	{8'd45,8'd33} : s = 78;
	{8'd45,8'd34} : s = 79;
	{8'd45,8'd35} : s = 80;
	{8'd45,8'd36} : s = 81;
	{8'd45,8'd37} : s = 82;
	{8'd45,8'd38} : s = 83;
	{8'd45,8'd39} : s = 84;
	{8'd45,8'd40} : s = 85;
	{8'd45,8'd41} : s = 86;
	{8'd45,8'd42} : s = 87;
	{8'd45,8'd43} : s = 88;
	{8'd45,8'd44} : s = 89;
	{8'd45,8'd45} : s = 90;
	{8'd45,8'd46} : s = 91;
	{8'd45,8'd47} : s = 92;
	{8'd45,8'd48} : s = 93;
	{8'd45,8'd49} : s = 94;
	{8'd45,8'd50} : s = 95;
	{8'd45,8'd51} : s = 96;
	{8'd45,8'd52} : s = 97;
	{8'd45,8'd53} : s = 98;
	{8'd45,8'd54} : s = 99;
	{8'd45,8'd55} : s = 100;
	{8'd45,8'd56} : s = 101;
	{8'd45,8'd57} : s = 102;
	{8'd45,8'd58} : s = 103;
	{8'd45,8'd59} : s = 104;
	{8'd45,8'd60} : s = 105;
	{8'd45,8'd61} : s = 106;
	{8'd45,8'd62} : s = 107;
	{8'd45,8'd63} : s = 108;
	{8'd45,8'd64} : s = 109;
	{8'd45,8'd65} : s = 110;
	{8'd45,8'd66} : s = 111;
	{8'd45,8'd67} : s = 112;
	{8'd45,8'd68} : s = 113;
	{8'd45,8'd69} : s = 114;
	{8'd45,8'd70} : s = 115;
	{8'd45,8'd71} : s = 116;
	{8'd45,8'd72} : s = 117;
	{8'd45,8'd73} : s = 118;
	{8'd45,8'd74} : s = 119;
	{8'd45,8'd75} : s = 120;
	{8'd45,8'd76} : s = 121;
	{8'd45,8'd77} : s = 122;
	{8'd45,8'd78} : s = 123;
	{8'd45,8'd79} : s = 124;
	{8'd45,8'd80} : s = 125;
	{8'd45,8'd81} : s = 126;
	{8'd45,8'd82} : s = 127;
	{8'd45,8'd83} : s = 128;
	{8'd45,8'd84} : s = 129;
	{8'd45,8'd85} : s = 130;
	{8'd45,8'd86} : s = 131;
	{8'd45,8'd87} : s = 132;
	{8'd45,8'd88} : s = 133;
	{8'd45,8'd89} : s = 134;
	{8'd45,8'd90} : s = 135;
	{8'd45,8'd91} : s = 136;
	{8'd45,8'd92} : s = 137;
	{8'd45,8'd93} : s = 138;
	{8'd45,8'd94} : s = 139;
	{8'd45,8'd95} : s = 140;
	{8'd45,8'd96} : s = 141;
	{8'd45,8'd97} : s = 142;
	{8'd45,8'd98} : s = 143;
	{8'd45,8'd99} : s = 144;
	{8'd45,8'd100} : s = 145;
	{8'd45,8'd101} : s = 146;
	{8'd45,8'd102} : s = 147;
	{8'd45,8'd103} : s = 148;
	{8'd45,8'd104} : s = 149;
	{8'd45,8'd105} : s = 150;
	{8'd45,8'd106} : s = 151;
	{8'd45,8'd107} : s = 152;
	{8'd45,8'd108} : s = 153;
	{8'd45,8'd109} : s = 154;
	{8'd45,8'd110} : s = 155;
	{8'd45,8'd111} : s = 156;
	{8'd45,8'd112} : s = 157;
	{8'd45,8'd113} : s = 158;
	{8'd45,8'd114} : s = 159;
	{8'd45,8'd115} : s = 160;
	{8'd45,8'd116} : s = 161;
	{8'd45,8'd117} : s = 162;
	{8'd45,8'd118} : s = 163;
	{8'd45,8'd119} : s = 164;
	{8'd45,8'd120} : s = 165;
	{8'd45,8'd121} : s = 166;
	{8'd45,8'd122} : s = 167;
	{8'd45,8'd123} : s = 168;
	{8'd45,8'd124} : s = 169;
	{8'd45,8'd125} : s = 170;
	{8'd45,8'd126} : s = 171;
	{8'd45,8'd127} : s = 172;
	{8'd45,8'd128} : s = 173;
	{8'd45,8'd129} : s = 174;
	{8'd45,8'd130} : s = 175;
	{8'd45,8'd131} : s = 176;
	{8'd45,8'd132} : s = 177;
	{8'd45,8'd133} : s = 178;
	{8'd45,8'd134} : s = 179;
	{8'd45,8'd135} : s = 180;
	{8'd45,8'd136} : s = 181;
	{8'd45,8'd137} : s = 182;
	{8'd45,8'd138} : s = 183;
	{8'd45,8'd139} : s = 184;
	{8'd45,8'd140} : s = 185;
	{8'd45,8'd141} : s = 186;
	{8'd45,8'd142} : s = 187;
	{8'd45,8'd143} : s = 188;
	{8'd45,8'd144} : s = 189;
	{8'd45,8'd145} : s = 190;
	{8'd45,8'd146} : s = 191;
	{8'd45,8'd147} : s = 192;
	{8'd45,8'd148} : s = 193;
	{8'd45,8'd149} : s = 194;
	{8'd45,8'd150} : s = 195;
	{8'd45,8'd151} : s = 196;
	{8'd45,8'd152} : s = 197;
	{8'd45,8'd153} : s = 198;
	{8'd45,8'd154} : s = 199;
	{8'd45,8'd155} : s = 200;
	{8'd45,8'd156} : s = 201;
	{8'd45,8'd157} : s = 202;
	{8'd45,8'd158} : s = 203;
	{8'd45,8'd159} : s = 204;
	{8'd45,8'd160} : s = 205;
	{8'd45,8'd161} : s = 206;
	{8'd45,8'd162} : s = 207;
	{8'd45,8'd163} : s = 208;
	{8'd45,8'd164} : s = 209;
	{8'd45,8'd165} : s = 210;
	{8'd45,8'd166} : s = 211;
	{8'd45,8'd167} : s = 212;
	{8'd45,8'd168} : s = 213;
	{8'd45,8'd169} : s = 214;
	{8'd45,8'd170} : s = 215;
	{8'd45,8'd171} : s = 216;
	{8'd45,8'd172} : s = 217;
	{8'd45,8'd173} : s = 218;
	{8'd45,8'd174} : s = 219;
	{8'd45,8'd175} : s = 220;
	{8'd45,8'd176} : s = 221;
	{8'd45,8'd177} : s = 222;
	{8'd45,8'd178} : s = 223;
	{8'd45,8'd179} : s = 224;
	{8'd45,8'd180} : s = 225;
	{8'd45,8'd181} : s = 226;
	{8'd45,8'd182} : s = 227;
	{8'd45,8'd183} : s = 228;
	{8'd45,8'd184} : s = 229;
	{8'd45,8'd185} : s = 230;
	{8'd45,8'd186} : s = 231;
	{8'd45,8'd187} : s = 232;
	{8'd45,8'd188} : s = 233;
	{8'd45,8'd189} : s = 234;
	{8'd45,8'd190} : s = 235;
	{8'd45,8'd191} : s = 236;
	{8'd45,8'd192} : s = 237;
	{8'd45,8'd193} : s = 238;
	{8'd45,8'd194} : s = 239;
	{8'd45,8'd195} : s = 240;
	{8'd45,8'd196} : s = 241;
	{8'd45,8'd197} : s = 242;
	{8'd45,8'd198} : s = 243;
	{8'd45,8'd199} : s = 244;
	{8'd45,8'd200} : s = 245;
	{8'd45,8'd201} : s = 246;
	{8'd45,8'd202} : s = 247;
	{8'd45,8'd203} : s = 248;
	{8'd45,8'd204} : s = 249;
	{8'd45,8'd205} : s = 250;
	{8'd45,8'd206} : s = 251;
	{8'd45,8'd207} : s = 252;
	{8'd45,8'd208} : s = 253;
	{8'd45,8'd209} : s = 254;
	{8'd45,8'd210} : s = 255;
	{8'd45,8'd211} : s = 256;
	{8'd45,8'd212} : s = 257;
	{8'd45,8'd213} : s = 258;
	{8'd45,8'd214} : s = 259;
	{8'd45,8'd215} : s = 260;
	{8'd45,8'd216} : s = 261;
	{8'd45,8'd217} : s = 262;
	{8'd45,8'd218} : s = 263;
	{8'd45,8'd219} : s = 264;
	{8'd45,8'd220} : s = 265;
	{8'd45,8'd221} : s = 266;
	{8'd45,8'd222} : s = 267;
	{8'd45,8'd223} : s = 268;
	{8'd45,8'd224} : s = 269;
	{8'd45,8'd225} : s = 270;
	{8'd45,8'd226} : s = 271;
	{8'd45,8'd227} : s = 272;
	{8'd45,8'd228} : s = 273;
	{8'd45,8'd229} : s = 274;
	{8'd45,8'd230} : s = 275;
	{8'd45,8'd231} : s = 276;
	{8'd45,8'd232} : s = 277;
	{8'd45,8'd233} : s = 278;
	{8'd45,8'd234} : s = 279;
	{8'd45,8'd235} : s = 280;
	{8'd45,8'd236} : s = 281;
	{8'd45,8'd237} : s = 282;
	{8'd45,8'd238} : s = 283;
	{8'd45,8'd239} : s = 284;
	{8'd45,8'd240} : s = 285;
	{8'd45,8'd241} : s = 286;
	{8'd45,8'd242} : s = 287;
	{8'd45,8'd243} : s = 288;
	{8'd45,8'd244} : s = 289;
	{8'd45,8'd245} : s = 290;
	{8'd45,8'd246} : s = 291;
	{8'd45,8'd247} : s = 292;
	{8'd45,8'd248} : s = 293;
	{8'd45,8'd249} : s = 294;
	{8'd45,8'd250} : s = 295;
	{8'd45,8'd251} : s = 296;
	{8'd45,8'd252} : s = 297;
	{8'd45,8'd253} : s = 298;
	{8'd45,8'd254} : s = 299;
	{8'd45,8'd255} : s = 300;
	{8'd46,8'd0} : s = 46;
	{8'd46,8'd1} : s = 47;
	{8'd46,8'd2} : s = 48;
	{8'd46,8'd3} : s = 49;
	{8'd46,8'd4} : s = 50;
	{8'd46,8'd5} : s = 51;
	{8'd46,8'd6} : s = 52;
	{8'd46,8'd7} : s = 53;
	{8'd46,8'd8} : s = 54;
	{8'd46,8'd9} : s = 55;
	{8'd46,8'd10} : s = 56;
	{8'd46,8'd11} : s = 57;
	{8'd46,8'd12} : s = 58;
	{8'd46,8'd13} : s = 59;
	{8'd46,8'd14} : s = 60;
	{8'd46,8'd15} : s = 61;
	{8'd46,8'd16} : s = 62;
	{8'd46,8'd17} : s = 63;
	{8'd46,8'd18} : s = 64;
	{8'd46,8'd19} : s = 65;
	{8'd46,8'd20} : s = 66;
	{8'd46,8'd21} : s = 67;
	{8'd46,8'd22} : s = 68;
	{8'd46,8'd23} : s = 69;
	{8'd46,8'd24} : s = 70;
	{8'd46,8'd25} : s = 71;
	{8'd46,8'd26} : s = 72;
	{8'd46,8'd27} : s = 73;
	{8'd46,8'd28} : s = 74;
	{8'd46,8'd29} : s = 75;
	{8'd46,8'd30} : s = 76;
	{8'd46,8'd31} : s = 77;
	{8'd46,8'd32} : s = 78;
	{8'd46,8'd33} : s = 79;
	{8'd46,8'd34} : s = 80;
	{8'd46,8'd35} : s = 81;
	{8'd46,8'd36} : s = 82;
	{8'd46,8'd37} : s = 83;
	{8'd46,8'd38} : s = 84;
	{8'd46,8'd39} : s = 85;
	{8'd46,8'd40} : s = 86;
	{8'd46,8'd41} : s = 87;
	{8'd46,8'd42} : s = 88;
	{8'd46,8'd43} : s = 89;
	{8'd46,8'd44} : s = 90;
	{8'd46,8'd45} : s = 91;
	{8'd46,8'd46} : s = 92;
	{8'd46,8'd47} : s = 93;
	{8'd46,8'd48} : s = 94;
	{8'd46,8'd49} : s = 95;
	{8'd46,8'd50} : s = 96;
	{8'd46,8'd51} : s = 97;
	{8'd46,8'd52} : s = 98;
	{8'd46,8'd53} : s = 99;
	{8'd46,8'd54} : s = 100;
	{8'd46,8'd55} : s = 101;
	{8'd46,8'd56} : s = 102;
	{8'd46,8'd57} : s = 103;
	{8'd46,8'd58} : s = 104;
	{8'd46,8'd59} : s = 105;
	{8'd46,8'd60} : s = 106;
	{8'd46,8'd61} : s = 107;
	{8'd46,8'd62} : s = 108;
	{8'd46,8'd63} : s = 109;
	{8'd46,8'd64} : s = 110;
	{8'd46,8'd65} : s = 111;
	{8'd46,8'd66} : s = 112;
	{8'd46,8'd67} : s = 113;
	{8'd46,8'd68} : s = 114;
	{8'd46,8'd69} : s = 115;
	{8'd46,8'd70} : s = 116;
	{8'd46,8'd71} : s = 117;
	{8'd46,8'd72} : s = 118;
	{8'd46,8'd73} : s = 119;
	{8'd46,8'd74} : s = 120;
	{8'd46,8'd75} : s = 121;
	{8'd46,8'd76} : s = 122;
	{8'd46,8'd77} : s = 123;
	{8'd46,8'd78} : s = 124;
	{8'd46,8'd79} : s = 125;
	{8'd46,8'd80} : s = 126;
	{8'd46,8'd81} : s = 127;
	{8'd46,8'd82} : s = 128;
	{8'd46,8'd83} : s = 129;
	{8'd46,8'd84} : s = 130;
	{8'd46,8'd85} : s = 131;
	{8'd46,8'd86} : s = 132;
	{8'd46,8'd87} : s = 133;
	{8'd46,8'd88} : s = 134;
	{8'd46,8'd89} : s = 135;
	{8'd46,8'd90} : s = 136;
	{8'd46,8'd91} : s = 137;
	{8'd46,8'd92} : s = 138;
	{8'd46,8'd93} : s = 139;
	{8'd46,8'd94} : s = 140;
	{8'd46,8'd95} : s = 141;
	{8'd46,8'd96} : s = 142;
	{8'd46,8'd97} : s = 143;
	{8'd46,8'd98} : s = 144;
	{8'd46,8'd99} : s = 145;
	{8'd46,8'd100} : s = 146;
	{8'd46,8'd101} : s = 147;
	{8'd46,8'd102} : s = 148;
	{8'd46,8'd103} : s = 149;
	{8'd46,8'd104} : s = 150;
	{8'd46,8'd105} : s = 151;
	{8'd46,8'd106} : s = 152;
	{8'd46,8'd107} : s = 153;
	{8'd46,8'd108} : s = 154;
	{8'd46,8'd109} : s = 155;
	{8'd46,8'd110} : s = 156;
	{8'd46,8'd111} : s = 157;
	{8'd46,8'd112} : s = 158;
	{8'd46,8'd113} : s = 159;
	{8'd46,8'd114} : s = 160;
	{8'd46,8'd115} : s = 161;
	{8'd46,8'd116} : s = 162;
	{8'd46,8'd117} : s = 163;
	{8'd46,8'd118} : s = 164;
	{8'd46,8'd119} : s = 165;
	{8'd46,8'd120} : s = 166;
	{8'd46,8'd121} : s = 167;
	{8'd46,8'd122} : s = 168;
	{8'd46,8'd123} : s = 169;
	{8'd46,8'd124} : s = 170;
	{8'd46,8'd125} : s = 171;
	{8'd46,8'd126} : s = 172;
	{8'd46,8'd127} : s = 173;
	{8'd46,8'd128} : s = 174;
	{8'd46,8'd129} : s = 175;
	{8'd46,8'd130} : s = 176;
	{8'd46,8'd131} : s = 177;
	{8'd46,8'd132} : s = 178;
	{8'd46,8'd133} : s = 179;
	{8'd46,8'd134} : s = 180;
	{8'd46,8'd135} : s = 181;
	{8'd46,8'd136} : s = 182;
	{8'd46,8'd137} : s = 183;
	{8'd46,8'd138} : s = 184;
	{8'd46,8'd139} : s = 185;
	{8'd46,8'd140} : s = 186;
	{8'd46,8'd141} : s = 187;
	{8'd46,8'd142} : s = 188;
	{8'd46,8'd143} : s = 189;
	{8'd46,8'd144} : s = 190;
	{8'd46,8'd145} : s = 191;
	{8'd46,8'd146} : s = 192;
	{8'd46,8'd147} : s = 193;
	{8'd46,8'd148} : s = 194;
	{8'd46,8'd149} : s = 195;
	{8'd46,8'd150} : s = 196;
	{8'd46,8'd151} : s = 197;
	{8'd46,8'd152} : s = 198;
	{8'd46,8'd153} : s = 199;
	{8'd46,8'd154} : s = 200;
	{8'd46,8'd155} : s = 201;
	{8'd46,8'd156} : s = 202;
	{8'd46,8'd157} : s = 203;
	{8'd46,8'd158} : s = 204;
	{8'd46,8'd159} : s = 205;
	{8'd46,8'd160} : s = 206;
	{8'd46,8'd161} : s = 207;
	{8'd46,8'd162} : s = 208;
	{8'd46,8'd163} : s = 209;
	{8'd46,8'd164} : s = 210;
	{8'd46,8'd165} : s = 211;
	{8'd46,8'd166} : s = 212;
	{8'd46,8'd167} : s = 213;
	{8'd46,8'd168} : s = 214;
	{8'd46,8'd169} : s = 215;
	{8'd46,8'd170} : s = 216;
	{8'd46,8'd171} : s = 217;
	{8'd46,8'd172} : s = 218;
	{8'd46,8'd173} : s = 219;
	{8'd46,8'd174} : s = 220;
	{8'd46,8'd175} : s = 221;
	{8'd46,8'd176} : s = 222;
	{8'd46,8'd177} : s = 223;
	{8'd46,8'd178} : s = 224;
	{8'd46,8'd179} : s = 225;
	{8'd46,8'd180} : s = 226;
	{8'd46,8'd181} : s = 227;
	{8'd46,8'd182} : s = 228;
	{8'd46,8'd183} : s = 229;
	{8'd46,8'd184} : s = 230;
	{8'd46,8'd185} : s = 231;
	{8'd46,8'd186} : s = 232;
	{8'd46,8'd187} : s = 233;
	{8'd46,8'd188} : s = 234;
	{8'd46,8'd189} : s = 235;
	{8'd46,8'd190} : s = 236;
	{8'd46,8'd191} : s = 237;
	{8'd46,8'd192} : s = 238;
	{8'd46,8'd193} : s = 239;
	{8'd46,8'd194} : s = 240;
	{8'd46,8'd195} : s = 241;
	{8'd46,8'd196} : s = 242;
	{8'd46,8'd197} : s = 243;
	{8'd46,8'd198} : s = 244;
	{8'd46,8'd199} : s = 245;
	{8'd46,8'd200} : s = 246;
	{8'd46,8'd201} : s = 247;
	{8'd46,8'd202} : s = 248;
	{8'd46,8'd203} : s = 249;
	{8'd46,8'd204} : s = 250;
	{8'd46,8'd205} : s = 251;
	{8'd46,8'd206} : s = 252;
	{8'd46,8'd207} : s = 253;
	{8'd46,8'd208} : s = 254;
	{8'd46,8'd209} : s = 255;
	{8'd46,8'd210} : s = 256;
	{8'd46,8'd211} : s = 257;
	{8'd46,8'd212} : s = 258;
	{8'd46,8'd213} : s = 259;
	{8'd46,8'd214} : s = 260;
	{8'd46,8'd215} : s = 261;
	{8'd46,8'd216} : s = 262;
	{8'd46,8'd217} : s = 263;
	{8'd46,8'd218} : s = 264;
	{8'd46,8'd219} : s = 265;
	{8'd46,8'd220} : s = 266;
	{8'd46,8'd221} : s = 267;
	{8'd46,8'd222} : s = 268;
	{8'd46,8'd223} : s = 269;
	{8'd46,8'd224} : s = 270;
	{8'd46,8'd225} : s = 271;
	{8'd46,8'd226} : s = 272;
	{8'd46,8'd227} : s = 273;
	{8'd46,8'd228} : s = 274;
	{8'd46,8'd229} : s = 275;
	{8'd46,8'd230} : s = 276;
	{8'd46,8'd231} : s = 277;
	{8'd46,8'd232} : s = 278;
	{8'd46,8'd233} : s = 279;
	{8'd46,8'd234} : s = 280;
	{8'd46,8'd235} : s = 281;
	{8'd46,8'd236} : s = 282;
	{8'd46,8'd237} : s = 283;
	{8'd46,8'd238} : s = 284;
	{8'd46,8'd239} : s = 285;
	{8'd46,8'd240} : s = 286;
	{8'd46,8'd241} : s = 287;
	{8'd46,8'd242} : s = 288;
	{8'd46,8'd243} : s = 289;
	{8'd46,8'd244} : s = 290;
	{8'd46,8'd245} : s = 291;
	{8'd46,8'd246} : s = 292;
	{8'd46,8'd247} : s = 293;
	{8'd46,8'd248} : s = 294;
	{8'd46,8'd249} : s = 295;
	{8'd46,8'd250} : s = 296;
	{8'd46,8'd251} : s = 297;
	{8'd46,8'd252} : s = 298;
	{8'd46,8'd253} : s = 299;
	{8'd46,8'd254} : s = 300;
	{8'd46,8'd255} : s = 301;
	{8'd47,8'd0} : s = 47;
	{8'd47,8'd1} : s = 48;
	{8'd47,8'd2} : s = 49;
	{8'd47,8'd3} : s = 50;
	{8'd47,8'd4} : s = 51;
	{8'd47,8'd5} : s = 52;
	{8'd47,8'd6} : s = 53;
	{8'd47,8'd7} : s = 54;
	{8'd47,8'd8} : s = 55;
	{8'd47,8'd9} : s = 56;
	{8'd47,8'd10} : s = 57;
	{8'd47,8'd11} : s = 58;
	{8'd47,8'd12} : s = 59;
	{8'd47,8'd13} : s = 60;
	{8'd47,8'd14} : s = 61;
	{8'd47,8'd15} : s = 62;
	{8'd47,8'd16} : s = 63;
	{8'd47,8'd17} : s = 64;
	{8'd47,8'd18} : s = 65;
	{8'd47,8'd19} : s = 66;
	{8'd47,8'd20} : s = 67;
	{8'd47,8'd21} : s = 68;
	{8'd47,8'd22} : s = 69;
	{8'd47,8'd23} : s = 70;
	{8'd47,8'd24} : s = 71;
	{8'd47,8'd25} : s = 72;
	{8'd47,8'd26} : s = 73;
	{8'd47,8'd27} : s = 74;
	{8'd47,8'd28} : s = 75;
	{8'd47,8'd29} : s = 76;
	{8'd47,8'd30} : s = 77;
	{8'd47,8'd31} : s = 78;
	{8'd47,8'd32} : s = 79;
	{8'd47,8'd33} : s = 80;
	{8'd47,8'd34} : s = 81;
	{8'd47,8'd35} : s = 82;
	{8'd47,8'd36} : s = 83;
	{8'd47,8'd37} : s = 84;
	{8'd47,8'd38} : s = 85;
	{8'd47,8'd39} : s = 86;
	{8'd47,8'd40} : s = 87;
	{8'd47,8'd41} : s = 88;
	{8'd47,8'd42} : s = 89;
	{8'd47,8'd43} : s = 90;
	{8'd47,8'd44} : s = 91;
	{8'd47,8'd45} : s = 92;
	{8'd47,8'd46} : s = 93;
	{8'd47,8'd47} : s = 94;
	{8'd47,8'd48} : s = 95;
	{8'd47,8'd49} : s = 96;
	{8'd47,8'd50} : s = 97;
	{8'd47,8'd51} : s = 98;
	{8'd47,8'd52} : s = 99;
	{8'd47,8'd53} : s = 100;
	{8'd47,8'd54} : s = 101;
	{8'd47,8'd55} : s = 102;
	{8'd47,8'd56} : s = 103;
	{8'd47,8'd57} : s = 104;
	{8'd47,8'd58} : s = 105;
	{8'd47,8'd59} : s = 106;
	{8'd47,8'd60} : s = 107;
	{8'd47,8'd61} : s = 108;
	{8'd47,8'd62} : s = 109;
	{8'd47,8'd63} : s = 110;
	{8'd47,8'd64} : s = 111;
	{8'd47,8'd65} : s = 112;
	{8'd47,8'd66} : s = 113;
	{8'd47,8'd67} : s = 114;
	{8'd47,8'd68} : s = 115;
	{8'd47,8'd69} : s = 116;
	{8'd47,8'd70} : s = 117;
	{8'd47,8'd71} : s = 118;
	{8'd47,8'd72} : s = 119;
	{8'd47,8'd73} : s = 120;
	{8'd47,8'd74} : s = 121;
	{8'd47,8'd75} : s = 122;
	{8'd47,8'd76} : s = 123;
	{8'd47,8'd77} : s = 124;
	{8'd47,8'd78} : s = 125;
	{8'd47,8'd79} : s = 126;
	{8'd47,8'd80} : s = 127;
	{8'd47,8'd81} : s = 128;
	{8'd47,8'd82} : s = 129;
	{8'd47,8'd83} : s = 130;
	{8'd47,8'd84} : s = 131;
	{8'd47,8'd85} : s = 132;
	{8'd47,8'd86} : s = 133;
	{8'd47,8'd87} : s = 134;
	{8'd47,8'd88} : s = 135;
	{8'd47,8'd89} : s = 136;
	{8'd47,8'd90} : s = 137;
	{8'd47,8'd91} : s = 138;
	{8'd47,8'd92} : s = 139;
	{8'd47,8'd93} : s = 140;
	{8'd47,8'd94} : s = 141;
	{8'd47,8'd95} : s = 142;
	{8'd47,8'd96} : s = 143;
	{8'd47,8'd97} : s = 144;
	{8'd47,8'd98} : s = 145;
	{8'd47,8'd99} : s = 146;
	{8'd47,8'd100} : s = 147;
	{8'd47,8'd101} : s = 148;
	{8'd47,8'd102} : s = 149;
	{8'd47,8'd103} : s = 150;
	{8'd47,8'd104} : s = 151;
	{8'd47,8'd105} : s = 152;
	{8'd47,8'd106} : s = 153;
	{8'd47,8'd107} : s = 154;
	{8'd47,8'd108} : s = 155;
	{8'd47,8'd109} : s = 156;
	{8'd47,8'd110} : s = 157;
	{8'd47,8'd111} : s = 158;
	{8'd47,8'd112} : s = 159;
	{8'd47,8'd113} : s = 160;
	{8'd47,8'd114} : s = 161;
	{8'd47,8'd115} : s = 162;
	{8'd47,8'd116} : s = 163;
	{8'd47,8'd117} : s = 164;
	{8'd47,8'd118} : s = 165;
	{8'd47,8'd119} : s = 166;
	{8'd47,8'd120} : s = 167;
	{8'd47,8'd121} : s = 168;
	{8'd47,8'd122} : s = 169;
	{8'd47,8'd123} : s = 170;
	{8'd47,8'd124} : s = 171;
	{8'd47,8'd125} : s = 172;
	{8'd47,8'd126} : s = 173;
	{8'd47,8'd127} : s = 174;
	{8'd47,8'd128} : s = 175;
	{8'd47,8'd129} : s = 176;
	{8'd47,8'd130} : s = 177;
	{8'd47,8'd131} : s = 178;
	{8'd47,8'd132} : s = 179;
	{8'd47,8'd133} : s = 180;
	{8'd47,8'd134} : s = 181;
	{8'd47,8'd135} : s = 182;
	{8'd47,8'd136} : s = 183;
	{8'd47,8'd137} : s = 184;
	{8'd47,8'd138} : s = 185;
	{8'd47,8'd139} : s = 186;
	{8'd47,8'd140} : s = 187;
	{8'd47,8'd141} : s = 188;
	{8'd47,8'd142} : s = 189;
	{8'd47,8'd143} : s = 190;
	{8'd47,8'd144} : s = 191;
	{8'd47,8'd145} : s = 192;
	{8'd47,8'd146} : s = 193;
	{8'd47,8'd147} : s = 194;
	{8'd47,8'd148} : s = 195;
	{8'd47,8'd149} : s = 196;
	{8'd47,8'd150} : s = 197;
	{8'd47,8'd151} : s = 198;
	{8'd47,8'd152} : s = 199;
	{8'd47,8'd153} : s = 200;
	{8'd47,8'd154} : s = 201;
	{8'd47,8'd155} : s = 202;
	{8'd47,8'd156} : s = 203;
	{8'd47,8'd157} : s = 204;
	{8'd47,8'd158} : s = 205;
	{8'd47,8'd159} : s = 206;
	{8'd47,8'd160} : s = 207;
	{8'd47,8'd161} : s = 208;
	{8'd47,8'd162} : s = 209;
	{8'd47,8'd163} : s = 210;
	{8'd47,8'd164} : s = 211;
	{8'd47,8'd165} : s = 212;
	{8'd47,8'd166} : s = 213;
	{8'd47,8'd167} : s = 214;
	{8'd47,8'd168} : s = 215;
	{8'd47,8'd169} : s = 216;
	{8'd47,8'd170} : s = 217;
	{8'd47,8'd171} : s = 218;
	{8'd47,8'd172} : s = 219;
	{8'd47,8'd173} : s = 220;
	{8'd47,8'd174} : s = 221;
	{8'd47,8'd175} : s = 222;
	{8'd47,8'd176} : s = 223;
	{8'd47,8'd177} : s = 224;
	{8'd47,8'd178} : s = 225;
	{8'd47,8'd179} : s = 226;
	{8'd47,8'd180} : s = 227;
	{8'd47,8'd181} : s = 228;
	{8'd47,8'd182} : s = 229;
	{8'd47,8'd183} : s = 230;
	{8'd47,8'd184} : s = 231;
	{8'd47,8'd185} : s = 232;
	{8'd47,8'd186} : s = 233;
	{8'd47,8'd187} : s = 234;
	{8'd47,8'd188} : s = 235;
	{8'd47,8'd189} : s = 236;
	{8'd47,8'd190} : s = 237;
	{8'd47,8'd191} : s = 238;
	{8'd47,8'd192} : s = 239;
	{8'd47,8'd193} : s = 240;
	{8'd47,8'd194} : s = 241;
	{8'd47,8'd195} : s = 242;
	{8'd47,8'd196} : s = 243;
	{8'd47,8'd197} : s = 244;
	{8'd47,8'd198} : s = 245;
	{8'd47,8'd199} : s = 246;
	{8'd47,8'd200} : s = 247;
	{8'd47,8'd201} : s = 248;
	{8'd47,8'd202} : s = 249;
	{8'd47,8'd203} : s = 250;
	{8'd47,8'd204} : s = 251;
	{8'd47,8'd205} : s = 252;
	{8'd47,8'd206} : s = 253;
	{8'd47,8'd207} : s = 254;
	{8'd47,8'd208} : s = 255;
	{8'd47,8'd209} : s = 256;
	{8'd47,8'd210} : s = 257;
	{8'd47,8'd211} : s = 258;
	{8'd47,8'd212} : s = 259;
	{8'd47,8'd213} : s = 260;
	{8'd47,8'd214} : s = 261;
	{8'd47,8'd215} : s = 262;
	{8'd47,8'd216} : s = 263;
	{8'd47,8'd217} : s = 264;
	{8'd47,8'd218} : s = 265;
	{8'd47,8'd219} : s = 266;
	{8'd47,8'd220} : s = 267;
	{8'd47,8'd221} : s = 268;
	{8'd47,8'd222} : s = 269;
	{8'd47,8'd223} : s = 270;
	{8'd47,8'd224} : s = 271;
	{8'd47,8'd225} : s = 272;
	{8'd47,8'd226} : s = 273;
	{8'd47,8'd227} : s = 274;
	{8'd47,8'd228} : s = 275;
	{8'd47,8'd229} : s = 276;
	{8'd47,8'd230} : s = 277;
	{8'd47,8'd231} : s = 278;
	{8'd47,8'd232} : s = 279;
	{8'd47,8'd233} : s = 280;
	{8'd47,8'd234} : s = 281;
	{8'd47,8'd235} : s = 282;
	{8'd47,8'd236} : s = 283;
	{8'd47,8'd237} : s = 284;
	{8'd47,8'd238} : s = 285;
	{8'd47,8'd239} : s = 286;
	{8'd47,8'd240} : s = 287;
	{8'd47,8'd241} : s = 288;
	{8'd47,8'd242} : s = 289;
	{8'd47,8'd243} : s = 290;
	{8'd47,8'd244} : s = 291;
	{8'd47,8'd245} : s = 292;
	{8'd47,8'd246} : s = 293;
	{8'd47,8'd247} : s = 294;
	{8'd47,8'd248} : s = 295;
	{8'd47,8'd249} : s = 296;
	{8'd47,8'd250} : s = 297;
	{8'd47,8'd251} : s = 298;
	{8'd47,8'd252} : s = 299;
	{8'd47,8'd253} : s = 300;
	{8'd47,8'd254} : s = 301;
	{8'd47,8'd255} : s = 302;
	{8'd48,8'd0} : s = 48;
	{8'd48,8'd1} : s = 49;
	{8'd48,8'd2} : s = 50;
	{8'd48,8'd3} : s = 51;
	{8'd48,8'd4} : s = 52;
	{8'd48,8'd5} : s = 53;
	{8'd48,8'd6} : s = 54;
	{8'd48,8'd7} : s = 55;
	{8'd48,8'd8} : s = 56;
	{8'd48,8'd9} : s = 57;
	{8'd48,8'd10} : s = 58;
	{8'd48,8'd11} : s = 59;
	{8'd48,8'd12} : s = 60;
	{8'd48,8'd13} : s = 61;
	{8'd48,8'd14} : s = 62;
	{8'd48,8'd15} : s = 63;
	{8'd48,8'd16} : s = 64;
	{8'd48,8'd17} : s = 65;
	{8'd48,8'd18} : s = 66;
	{8'd48,8'd19} : s = 67;
	{8'd48,8'd20} : s = 68;
	{8'd48,8'd21} : s = 69;
	{8'd48,8'd22} : s = 70;
	{8'd48,8'd23} : s = 71;
	{8'd48,8'd24} : s = 72;
	{8'd48,8'd25} : s = 73;
	{8'd48,8'd26} : s = 74;
	{8'd48,8'd27} : s = 75;
	{8'd48,8'd28} : s = 76;
	{8'd48,8'd29} : s = 77;
	{8'd48,8'd30} : s = 78;
	{8'd48,8'd31} : s = 79;
	{8'd48,8'd32} : s = 80;
	{8'd48,8'd33} : s = 81;
	{8'd48,8'd34} : s = 82;
	{8'd48,8'd35} : s = 83;
	{8'd48,8'd36} : s = 84;
	{8'd48,8'd37} : s = 85;
	{8'd48,8'd38} : s = 86;
	{8'd48,8'd39} : s = 87;
	{8'd48,8'd40} : s = 88;
	{8'd48,8'd41} : s = 89;
	{8'd48,8'd42} : s = 90;
	{8'd48,8'd43} : s = 91;
	{8'd48,8'd44} : s = 92;
	{8'd48,8'd45} : s = 93;
	{8'd48,8'd46} : s = 94;
	{8'd48,8'd47} : s = 95;
	{8'd48,8'd48} : s = 96;
	{8'd48,8'd49} : s = 97;
	{8'd48,8'd50} : s = 98;
	{8'd48,8'd51} : s = 99;
	{8'd48,8'd52} : s = 100;
	{8'd48,8'd53} : s = 101;
	{8'd48,8'd54} : s = 102;
	{8'd48,8'd55} : s = 103;
	{8'd48,8'd56} : s = 104;
	{8'd48,8'd57} : s = 105;
	{8'd48,8'd58} : s = 106;
	{8'd48,8'd59} : s = 107;
	{8'd48,8'd60} : s = 108;
	{8'd48,8'd61} : s = 109;
	{8'd48,8'd62} : s = 110;
	{8'd48,8'd63} : s = 111;
	{8'd48,8'd64} : s = 112;
	{8'd48,8'd65} : s = 113;
	{8'd48,8'd66} : s = 114;
	{8'd48,8'd67} : s = 115;
	{8'd48,8'd68} : s = 116;
	{8'd48,8'd69} : s = 117;
	{8'd48,8'd70} : s = 118;
	{8'd48,8'd71} : s = 119;
	{8'd48,8'd72} : s = 120;
	{8'd48,8'd73} : s = 121;
	{8'd48,8'd74} : s = 122;
	{8'd48,8'd75} : s = 123;
	{8'd48,8'd76} : s = 124;
	{8'd48,8'd77} : s = 125;
	{8'd48,8'd78} : s = 126;
	{8'd48,8'd79} : s = 127;
	{8'd48,8'd80} : s = 128;
	{8'd48,8'd81} : s = 129;
	{8'd48,8'd82} : s = 130;
	{8'd48,8'd83} : s = 131;
	{8'd48,8'd84} : s = 132;
	{8'd48,8'd85} : s = 133;
	{8'd48,8'd86} : s = 134;
	{8'd48,8'd87} : s = 135;
	{8'd48,8'd88} : s = 136;
	{8'd48,8'd89} : s = 137;
	{8'd48,8'd90} : s = 138;
	{8'd48,8'd91} : s = 139;
	{8'd48,8'd92} : s = 140;
	{8'd48,8'd93} : s = 141;
	{8'd48,8'd94} : s = 142;
	{8'd48,8'd95} : s = 143;
	{8'd48,8'd96} : s = 144;
	{8'd48,8'd97} : s = 145;
	{8'd48,8'd98} : s = 146;
	{8'd48,8'd99} : s = 147;
	{8'd48,8'd100} : s = 148;
	{8'd48,8'd101} : s = 149;
	{8'd48,8'd102} : s = 150;
	{8'd48,8'd103} : s = 151;
	{8'd48,8'd104} : s = 152;
	{8'd48,8'd105} : s = 153;
	{8'd48,8'd106} : s = 154;
	{8'd48,8'd107} : s = 155;
	{8'd48,8'd108} : s = 156;
	{8'd48,8'd109} : s = 157;
	{8'd48,8'd110} : s = 158;
	{8'd48,8'd111} : s = 159;
	{8'd48,8'd112} : s = 160;
	{8'd48,8'd113} : s = 161;
	{8'd48,8'd114} : s = 162;
	{8'd48,8'd115} : s = 163;
	{8'd48,8'd116} : s = 164;
	{8'd48,8'd117} : s = 165;
	{8'd48,8'd118} : s = 166;
	{8'd48,8'd119} : s = 167;
	{8'd48,8'd120} : s = 168;
	{8'd48,8'd121} : s = 169;
	{8'd48,8'd122} : s = 170;
	{8'd48,8'd123} : s = 171;
	{8'd48,8'd124} : s = 172;
	{8'd48,8'd125} : s = 173;
	{8'd48,8'd126} : s = 174;
	{8'd48,8'd127} : s = 175;
	{8'd48,8'd128} : s = 176;
	{8'd48,8'd129} : s = 177;
	{8'd48,8'd130} : s = 178;
	{8'd48,8'd131} : s = 179;
	{8'd48,8'd132} : s = 180;
	{8'd48,8'd133} : s = 181;
	{8'd48,8'd134} : s = 182;
	{8'd48,8'd135} : s = 183;
	{8'd48,8'd136} : s = 184;
	{8'd48,8'd137} : s = 185;
	{8'd48,8'd138} : s = 186;
	{8'd48,8'd139} : s = 187;
	{8'd48,8'd140} : s = 188;
	{8'd48,8'd141} : s = 189;
	{8'd48,8'd142} : s = 190;
	{8'd48,8'd143} : s = 191;
	{8'd48,8'd144} : s = 192;
	{8'd48,8'd145} : s = 193;
	{8'd48,8'd146} : s = 194;
	{8'd48,8'd147} : s = 195;
	{8'd48,8'd148} : s = 196;
	{8'd48,8'd149} : s = 197;
	{8'd48,8'd150} : s = 198;
	{8'd48,8'd151} : s = 199;
	{8'd48,8'd152} : s = 200;
	{8'd48,8'd153} : s = 201;
	{8'd48,8'd154} : s = 202;
	{8'd48,8'd155} : s = 203;
	{8'd48,8'd156} : s = 204;
	{8'd48,8'd157} : s = 205;
	{8'd48,8'd158} : s = 206;
	{8'd48,8'd159} : s = 207;
	{8'd48,8'd160} : s = 208;
	{8'd48,8'd161} : s = 209;
	{8'd48,8'd162} : s = 210;
	{8'd48,8'd163} : s = 211;
	{8'd48,8'd164} : s = 212;
	{8'd48,8'd165} : s = 213;
	{8'd48,8'd166} : s = 214;
	{8'd48,8'd167} : s = 215;
	{8'd48,8'd168} : s = 216;
	{8'd48,8'd169} : s = 217;
	{8'd48,8'd170} : s = 218;
	{8'd48,8'd171} : s = 219;
	{8'd48,8'd172} : s = 220;
	{8'd48,8'd173} : s = 221;
	{8'd48,8'd174} : s = 222;
	{8'd48,8'd175} : s = 223;
	{8'd48,8'd176} : s = 224;
	{8'd48,8'd177} : s = 225;
	{8'd48,8'd178} : s = 226;
	{8'd48,8'd179} : s = 227;
	{8'd48,8'd180} : s = 228;
	{8'd48,8'd181} : s = 229;
	{8'd48,8'd182} : s = 230;
	{8'd48,8'd183} : s = 231;
	{8'd48,8'd184} : s = 232;
	{8'd48,8'd185} : s = 233;
	{8'd48,8'd186} : s = 234;
	{8'd48,8'd187} : s = 235;
	{8'd48,8'd188} : s = 236;
	{8'd48,8'd189} : s = 237;
	{8'd48,8'd190} : s = 238;
	{8'd48,8'd191} : s = 239;
	{8'd48,8'd192} : s = 240;
	{8'd48,8'd193} : s = 241;
	{8'd48,8'd194} : s = 242;
	{8'd48,8'd195} : s = 243;
	{8'd48,8'd196} : s = 244;
	{8'd48,8'd197} : s = 245;
	{8'd48,8'd198} : s = 246;
	{8'd48,8'd199} : s = 247;
	{8'd48,8'd200} : s = 248;
	{8'd48,8'd201} : s = 249;
	{8'd48,8'd202} : s = 250;
	{8'd48,8'd203} : s = 251;
	{8'd48,8'd204} : s = 252;
	{8'd48,8'd205} : s = 253;
	{8'd48,8'd206} : s = 254;
	{8'd48,8'd207} : s = 255;
	{8'd48,8'd208} : s = 256;
	{8'd48,8'd209} : s = 257;
	{8'd48,8'd210} : s = 258;
	{8'd48,8'd211} : s = 259;
	{8'd48,8'd212} : s = 260;
	{8'd48,8'd213} : s = 261;
	{8'd48,8'd214} : s = 262;
	{8'd48,8'd215} : s = 263;
	{8'd48,8'd216} : s = 264;
	{8'd48,8'd217} : s = 265;
	{8'd48,8'd218} : s = 266;
	{8'd48,8'd219} : s = 267;
	{8'd48,8'd220} : s = 268;
	{8'd48,8'd221} : s = 269;
	{8'd48,8'd222} : s = 270;
	{8'd48,8'd223} : s = 271;
	{8'd48,8'd224} : s = 272;
	{8'd48,8'd225} : s = 273;
	{8'd48,8'd226} : s = 274;
	{8'd48,8'd227} : s = 275;
	{8'd48,8'd228} : s = 276;
	{8'd48,8'd229} : s = 277;
	{8'd48,8'd230} : s = 278;
	{8'd48,8'd231} : s = 279;
	{8'd48,8'd232} : s = 280;
	{8'd48,8'd233} : s = 281;
	{8'd48,8'd234} : s = 282;
	{8'd48,8'd235} : s = 283;
	{8'd48,8'd236} : s = 284;
	{8'd48,8'd237} : s = 285;
	{8'd48,8'd238} : s = 286;
	{8'd48,8'd239} : s = 287;
	{8'd48,8'd240} : s = 288;
	{8'd48,8'd241} : s = 289;
	{8'd48,8'd242} : s = 290;
	{8'd48,8'd243} : s = 291;
	{8'd48,8'd244} : s = 292;
	{8'd48,8'd245} : s = 293;
	{8'd48,8'd246} : s = 294;
	{8'd48,8'd247} : s = 295;
	{8'd48,8'd248} : s = 296;
	{8'd48,8'd249} : s = 297;
	{8'd48,8'd250} : s = 298;
	{8'd48,8'd251} : s = 299;
	{8'd48,8'd252} : s = 300;
	{8'd48,8'd253} : s = 301;
	{8'd48,8'd254} : s = 302;
	{8'd48,8'd255} : s = 303;
	{8'd49,8'd0} : s = 49;
	{8'd49,8'd1} : s = 50;
	{8'd49,8'd2} : s = 51;
	{8'd49,8'd3} : s = 52;
	{8'd49,8'd4} : s = 53;
	{8'd49,8'd5} : s = 54;
	{8'd49,8'd6} : s = 55;
	{8'd49,8'd7} : s = 56;
	{8'd49,8'd8} : s = 57;
	{8'd49,8'd9} : s = 58;
	{8'd49,8'd10} : s = 59;
	{8'd49,8'd11} : s = 60;
	{8'd49,8'd12} : s = 61;
	{8'd49,8'd13} : s = 62;
	{8'd49,8'd14} : s = 63;
	{8'd49,8'd15} : s = 64;
	{8'd49,8'd16} : s = 65;
	{8'd49,8'd17} : s = 66;
	{8'd49,8'd18} : s = 67;
	{8'd49,8'd19} : s = 68;
	{8'd49,8'd20} : s = 69;
	{8'd49,8'd21} : s = 70;
	{8'd49,8'd22} : s = 71;
	{8'd49,8'd23} : s = 72;
	{8'd49,8'd24} : s = 73;
	{8'd49,8'd25} : s = 74;
	{8'd49,8'd26} : s = 75;
	{8'd49,8'd27} : s = 76;
	{8'd49,8'd28} : s = 77;
	{8'd49,8'd29} : s = 78;
	{8'd49,8'd30} : s = 79;
	{8'd49,8'd31} : s = 80;
	{8'd49,8'd32} : s = 81;
	{8'd49,8'd33} : s = 82;
	{8'd49,8'd34} : s = 83;
	{8'd49,8'd35} : s = 84;
	{8'd49,8'd36} : s = 85;
	{8'd49,8'd37} : s = 86;
	{8'd49,8'd38} : s = 87;
	{8'd49,8'd39} : s = 88;
	{8'd49,8'd40} : s = 89;
	{8'd49,8'd41} : s = 90;
	{8'd49,8'd42} : s = 91;
	{8'd49,8'd43} : s = 92;
	{8'd49,8'd44} : s = 93;
	{8'd49,8'd45} : s = 94;
	{8'd49,8'd46} : s = 95;
	{8'd49,8'd47} : s = 96;
	{8'd49,8'd48} : s = 97;
	{8'd49,8'd49} : s = 98;
	{8'd49,8'd50} : s = 99;
	{8'd49,8'd51} : s = 100;
	{8'd49,8'd52} : s = 101;
	{8'd49,8'd53} : s = 102;
	{8'd49,8'd54} : s = 103;
	{8'd49,8'd55} : s = 104;
	{8'd49,8'd56} : s = 105;
	{8'd49,8'd57} : s = 106;
	{8'd49,8'd58} : s = 107;
	{8'd49,8'd59} : s = 108;
	{8'd49,8'd60} : s = 109;
	{8'd49,8'd61} : s = 110;
	{8'd49,8'd62} : s = 111;
	{8'd49,8'd63} : s = 112;
	{8'd49,8'd64} : s = 113;
	{8'd49,8'd65} : s = 114;
	{8'd49,8'd66} : s = 115;
	{8'd49,8'd67} : s = 116;
	{8'd49,8'd68} : s = 117;
	{8'd49,8'd69} : s = 118;
	{8'd49,8'd70} : s = 119;
	{8'd49,8'd71} : s = 120;
	{8'd49,8'd72} : s = 121;
	{8'd49,8'd73} : s = 122;
	{8'd49,8'd74} : s = 123;
	{8'd49,8'd75} : s = 124;
	{8'd49,8'd76} : s = 125;
	{8'd49,8'd77} : s = 126;
	{8'd49,8'd78} : s = 127;
	{8'd49,8'd79} : s = 128;
	{8'd49,8'd80} : s = 129;
	{8'd49,8'd81} : s = 130;
	{8'd49,8'd82} : s = 131;
	{8'd49,8'd83} : s = 132;
	{8'd49,8'd84} : s = 133;
	{8'd49,8'd85} : s = 134;
	{8'd49,8'd86} : s = 135;
	{8'd49,8'd87} : s = 136;
	{8'd49,8'd88} : s = 137;
	{8'd49,8'd89} : s = 138;
	{8'd49,8'd90} : s = 139;
	{8'd49,8'd91} : s = 140;
	{8'd49,8'd92} : s = 141;
	{8'd49,8'd93} : s = 142;
	{8'd49,8'd94} : s = 143;
	{8'd49,8'd95} : s = 144;
	{8'd49,8'd96} : s = 145;
	{8'd49,8'd97} : s = 146;
	{8'd49,8'd98} : s = 147;
	{8'd49,8'd99} : s = 148;
	{8'd49,8'd100} : s = 149;
	{8'd49,8'd101} : s = 150;
	{8'd49,8'd102} : s = 151;
	{8'd49,8'd103} : s = 152;
	{8'd49,8'd104} : s = 153;
	{8'd49,8'd105} : s = 154;
	{8'd49,8'd106} : s = 155;
	{8'd49,8'd107} : s = 156;
	{8'd49,8'd108} : s = 157;
	{8'd49,8'd109} : s = 158;
	{8'd49,8'd110} : s = 159;
	{8'd49,8'd111} : s = 160;
	{8'd49,8'd112} : s = 161;
	{8'd49,8'd113} : s = 162;
	{8'd49,8'd114} : s = 163;
	{8'd49,8'd115} : s = 164;
	{8'd49,8'd116} : s = 165;
	{8'd49,8'd117} : s = 166;
	{8'd49,8'd118} : s = 167;
	{8'd49,8'd119} : s = 168;
	{8'd49,8'd120} : s = 169;
	{8'd49,8'd121} : s = 170;
	{8'd49,8'd122} : s = 171;
	{8'd49,8'd123} : s = 172;
	{8'd49,8'd124} : s = 173;
	{8'd49,8'd125} : s = 174;
	{8'd49,8'd126} : s = 175;
	{8'd49,8'd127} : s = 176;
	{8'd49,8'd128} : s = 177;
	{8'd49,8'd129} : s = 178;
	{8'd49,8'd130} : s = 179;
	{8'd49,8'd131} : s = 180;
	{8'd49,8'd132} : s = 181;
	{8'd49,8'd133} : s = 182;
	{8'd49,8'd134} : s = 183;
	{8'd49,8'd135} : s = 184;
	{8'd49,8'd136} : s = 185;
	{8'd49,8'd137} : s = 186;
	{8'd49,8'd138} : s = 187;
	{8'd49,8'd139} : s = 188;
	{8'd49,8'd140} : s = 189;
	{8'd49,8'd141} : s = 190;
	{8'd49,8'd142} : s = 191;
	{8'd49,8'd143} : s = 192;
	{8'd49,8'd144} : s = 193;
	{8'd49,8'd145} : s = 194;
	{8'd49,8'd146} : s = 195;
	{8'd49,8'd147} : s = 196;
	{8'd49,8'd148} : s = 197;
	{8'd49,8'd149} : s = 198;
	{8'd49,8'd150} : s = 199;
	{8'd49,8'd151} : s = 200;
	{8'd49,8'd152} : s = 201;
	{8'd49,8'd153} : s = 202;
	{8'd49,8'd154} : s = 203;
	{8'd49,8'd155} : s = 204;
	{8'd49,8'd156} : s = 205;
	{8'd49,8'd157} : s = 206;
	{8'd49,8'd158} : s = 207;
	{8'd49,8'd159} : s = 208;
	{8'd49,8'd160} : s = 209;
	{8'd49,8'd161} : s = 210;
	{8'd49,8'd162} : s = 211;
	{8'd49,8'd163} : s = 212;
	{8'd49,8'd164} : s = 213;
	{8'd49,8'd165} : s = 214;
	{8'd49,8'd166} : s = 215;
	{8'd49,8'd167} : s = 216;
	{8'd49,8'd168} : s = 217;
	{8'd49,8'd169} : s = 218;
	{8'd49,8'd170} : s = 219;
	{8'd49,8'd171} : s = 220;
	{8'd49,8'd172} : s = 221;
	{8'd49,8'd173} : s = 222;
	{8'd49,8'd174} : s = 223;
	{8'd49,8'd175} : s = 224;
	{8'd49,8'd176} : s = 225;
	{8'd49,8'd177} : s = 226;
	{8'd49,8'd178} : s = 227;
	{8'd49,8'd179} : s = 228;
	{8'd49,8'd180} : s = 229;
	{8'd49,8'd181} : s = 230;
	{8'd49,8'd182} : s = 231;
	{8'd49,8'd183} : s = 232;
	{8'd49,8'd184} : s = 233;
	{8'd49,8'd185} : s = 234;
	{8'd49,8'd186} : s = 235;
	{8'd49,8'd187} : s = 236;
	{8'd49,8'd188} : s = 237;
	{8'd49,8'd189} : s = 238;
	{8'd49,8'd190} : s = 239;
	{8'd49,8'd191} : s = 240;
	{8'd49,8'd192} : s = 241;
	{8'd49,8'd193} : s = 242;
	{8'd49,8'd194} : s = 243;
	{8'd49,8'd195} : s = 244;
	{8'd49,8'd196} : s = 245;
	{8'd49,8'd197} : s = 246;
	{8'd49,8'd198} : s = 247;
	{8'd49,8'd199} : s = 248;
	{8'd49,8'd200} : s = 249;
	{8'd49,8'd201} : s = 250;
	{8'd49,8'd202} : s = 251;
	{8'd49,8'd203} : s = 252;
	{8'd49,8'd204} : s = 253;
	{8'd49,8'd205} : s = 254;
	{8'd49,8'd206} : s = 255;
	{8'd49,8'd207} : s = 256;
	{8'd49,8'd208} : s = 257;
	{8'd49,8'd209} : s = 258;
	{8'd49,8'd210} : s = 259;
	{8'd49,8'd211} : s = 260;
	{8'd49,8'd212} : s = 261;
	{8'd49,8'd213} : s = 262;
	{8'd49,8'd214} : s = 263;
	{8'd49,8'd215} : s = 264;
	{8'd49,8'd216} : s = 265;
	{8'd49,8'd217} : s = 266;
	{8'd49,8'd218} : s = 267;
	{8'd49,8'd219} : s = 268;
	{8'd49,8'd220} : s = 269;
	{8'd49,8'd221} : s = 270;
	{8'd49,8'd222} : s = 271;
	{8'd49,8'd223} : s = 272;
	{8'd49,8'd224} : s = 273;
	{8'd49,8'd225} : s = 274;
	{8'd49,8'd226} : s = 275;
	{8'd49,8'd227} : s = 276;
	{8'd49,8'd228} : s = 277;
	{8'd49,8'd229} : s = 278;
	{8'd49,8'd230} : s = 279;
	{8'd49,8'd231} : s = 280;
	{8'd49,8'd232} : s = 281;
	{8'd49,8'd233} : s = 282;
	{8'd49,8'd234} : s = 283;
	{8'd49,8'd235} : s = 284;
	{8'd49,8'd236} : s = 285;
	{8'd49,8'd237} : s = 286;
	{8'd49,8'd238} : s = 287;
	{8'd49,8'd239} : s = 288;
	{8'd49,8'd240} : s = 289;
	{8'd49,8'd241} : s = 290;
	{8'd49,8'd242} : s = 291;
	{8'd49,8'd243} : s = 292;
	{8'd49,8'd244} : s = 293;
	{8'd49,8'd245} : s = 294;
	{8'd49,8'd246} : s = 295;
	{8'd49,8'd247} : s = 296;
	{8'd49,8'd248} : s = 297;
	{8'd49,8'd249} : s = 298;
	{8'd49,8'd250} : s = 299;
	{8'd49,8'd251} : s = 300;
	{8'd49,8'd252} : s = 301;
	{8'd49,8'd253} : s = 302;
	{8'd49,8'd254} : s = 303;
	{8'd49,8'd255} : s = 304;
	{8'd50,8'd0} : s = 50;
	{8'd50,8'd1} : s = 51;
	{8'd50,8'd2} : s = 52;
	{8'd50,8'd3} : s = 53;
	{8'd50,8'd4} : s = 54;
	{8'd50,8'd5} : s = 55;
	{8'd50,8'd6} : s = 56;
	{8'd50,8'd7} : s = 57;
	{8'd50,8'd8} : s = 58;
	{8'd50,8'd9} : s = 59;
	{8'd50,8'd10} : s = 60;
	{8'd50,8'd11} : s = 61;
	{8'd50,8'd12} : s = 62;
	{8'd50,8'd13} : s = 63;
	{8'd50,8'd14} : s = 64;
	{8'd50,8'd15} : s = 65;
	{8'd50,8'd16} : s = 66;
	{8'd50,8'd17} : s = 67;
	{8'd50,8'd18} : s = 68;
	{8'd50,8'd19} : s = 69;
	{8'd50,8'd20} : s = 70;
	{8'd50,8'd21} : s = 71;
	{8'd50,8'd22} : s = 72;
	{8'd50,8'd23} : s = 73;
	{8'd50,8'd24} : s = 74;
	{8'd50,8'd25} : s = 75;
	{8'd50,8'd26} : s = 76;
	{8'd50,8'd27} : s = 77;
	{8'd50,8'd28} : s = 78;
	{8'd50,8'd29} : s = 79;
	{8'd50,8'd30} : s = 80;
	{8'd50,8'd31} : s = 81;
	{8'd50,8'd32} : s = 82;
	{8'd50,8'd33} : s = 83;
	{8'd50,8'd34} : s = 84;
	{8'd50,8'd35} : s = 85;
	{8'd50,8'd36} : s = 86;
	{8'd50,8'd37} : s = 87;
	{8'd50,8'd38} : s = 88;
	{8'd50,8'd39} : s = 89;
	{8'd50,8'd40} : s = 90;
	{8'd50,8'd41} : s = 91;
	{8'd50,8'd42} : s = 92;
	{8'd50,8'd43} : s = 93;
	{8'd50,8'd44} : s = 94;
	{8'd50,8'd45} : s = 95;
	{8'd50,8'd46} : s = 96;
	{8'd50,8'd47} : s = 97;
	{8'd50,8'd48} : s = 98;
	{8'd50,8'd49} : s = 99;
	{8'd50,8'd50} : s = 100;
	{8'd50,8'd51} : s = 101;
	{8'd50,8'd52} : s = 102;
	{8'd50,8'd53} : s = 103;
	{8'd50,8'd54} : s = 104;
	{8'd50,8'd55} : s = 105;
	{8'd50,8'd56} : s = 106;
	{8'd50,8'd57} : s = 107;
	{8'd50,8'd58} : s = 108;
	{8'd50,8'd59} : s = 109;
	{8'd50,8'd60} : s = 110;
	{8'd50,8'd61} : s = 111;
	{8'd50,8'd62} : s = 112;
	{8'd50,8'd63} : s = 113;
	{8'd50,8'd64} : s = 114;
	{8'd50,8'd65} : s = 115;
	{8'd50,8'd66} : s = 116;
	{8'd50,8'd67} : s = 117;
	{8'd50,8'd68} : s = 118;
	{8'd50,8'd69} : s = 119;
	{8'd50,8'd70} : s = 120;
	{8'd50,8'd71} : s = 121;
	{8'd50,8'd72} : s = 122;
	{8'd50,8'd73} : s = 123;
	{8'd50,8'd74} : s = 124;
	{8'd50,8'd75} : s = 125;
	{8'd50,8'd76} : s = 126;
	{8'd50,8'd77} : s = 127;
	{8'd50,8'd78} : s = 128;
	{8'd50,8'd79} : s = 129;
	{8'd50,8'd80} : s = 130;
	{8'd50,8'd81} : s = 131;
	{8'd50,8'd82} : s = 132;
	{8'd50,8'd83} : s = 133;
	{8'd50,8'd84} : s = 134;
	{8'd50,8'd85} : s = 135;
	{8'd50,8'd86} : s = 136;
	{8'd50,8'd87} : s = 137;
	{8'd50,8'd88} : s = 138;
	{8'd50,8'd89} : s = 139;
	{8'd50,8'd90} : s = 140;
	{8'd50,8'd91} : s = 141;
	{8'd50,8'd92} : s = 142;
	{8'd50,8'd93} : s = 143;
	{8'd50,8'd94} : s = 144;
	{8'd50,8'd95} : s = 145;
	{8'd50,8'd96} : s = 146;
	{8'd50,8'd97} : s = 147;
	{8'd50,8'd98} : s = 148;
	{8'd50,8'd99} : s = 149;
	{8'd50,8'd100} : s = 150;
	{8'd50,8'd101} : s = 151;
	{8'd50,8'd102} : s = 152;
	{8'd50,8'd103} : s = 153;
	{8'd50,8'd104} : s = 154;
	{8'd50,8'd105} : s = 155;
	{8'd50,8'd106} : s = 156;
	{8'd50,8'd107} : s = 157;
	{8'd50,8'd108} : s = 158;
	{8'd50,8'd109} : s = 159;
	{8'd50,8'd110} : s = 160;
	{8'd50,8'd111} : s = 161;
	{8'd50,8'd112} : s = 162;
	{8'd50,8'd113} : s = 163;
	{8'd50,8'd114} : s = 164;
	{8'd50,8'd115} : s = 165;
	{8'd50,8'd116} : s = 166;
	{8'd50,8'd117} : s = 167;
	{8'd50,8'd118} : s = 168;
	{8'd50,8'd119} : s = 169;
	{8'd50,8'd120} : s = 170;
	{8'd50,8'd121} : s = 171;
	{8'd50,8'd122} : s = 172;
	{8'd50,8'd123} : s = 173;
	{8'd50,8'd124} : s = 174;
	{8'd50,8'd125} : s = 175;
	{8'd50,8'd126} : s = 176;
	{8'd50,8'd127} : s = 177;
	{8'd50,8'd128} : s = 178;
	{8'd50,8'd129} : s = 179;
	{8'd50,8'd130} : s = 180;
	{8'd50,8'd131} : s = 181;
	{8'd50,8'd132} : s = 182;
	{8'd50,8'd133} : s = 183;
	{8'd50,8'd134} : s = 184;
	{8'd50,8'd135} : s = 185;
	{8'd50,8'd136} : s = 186;
	{8'd50,8'd137} : s = 187;
	{8'd50,8'd138} : s = 188;
	{8'd50,8'd139} : s = 189;
	{8'd50,8'd140} : s = 190;
	{8'd50,8'd141} : s = 191;
	{8'd50,8'd142} : s = 192;
	{8'd50,8'd143} : s = 193;
	{8'd50,8'd144} : s = 194;
	{8'd50,8'd145} : s = 195;
	{8'd50,8'd146} : s = 196;
	{8'd50,8'd147} : s = 197;
	{8'd50,8'd148} : s = 198;
	{8'd50,8'd149} : s = 199;
	{8'd50,8'd150} : s = 200;
	{8'd50,8'd151} : s = 201;
	{8'd50,8'd152} : s = 202;
	{8'd50,8'd153} : s = 203;
	{8'd50,8'd154} : s = 204;
	{8'd50,8'd155} : s = 205;
	{8'd50,8'd156} : s = 206;
	{8'd50,8'd157} : s = 207;
	{8'd50,8'd158} : s = 208;
	{8'd50,8'd159} : s = 209;
	{8'd50,8'd160} : s = 210;
	{8'd50,8'd161} : s = 211;
	{8'd50,8'd162} : s = 212;
	{8'd50,8'd163} : s = 213;
	{8'd50,8'd164} : s = 214;
	{8'd50,8'd165} : s = 215;
	{8'd50,8'd166} : s = 216;
	{8'd50,8'd167} : s = 217;
	{8'd50,8'd168} : s = 218;
	{8'd50,8'd169} : s = 219;
	{8'd50,8'd170} : s = 220;
	{8'd50,8'd171} : s = 221;
	{8'd50,8'd172} : s = 222;
	{8'd50,8'd173} : s = 223;
	{8'd50,8'd174} : s = 224;
	{8'd50,8'd175} : s = 225;
	{8'd50,8'd176} : s = 226;
	{8'd50,8'd177} : s = 227;
	{8'd50,8'd178} : s = 228;
	{8'd50,8'd179} : s = 229;
	{8'd50,8'd180} : s = 230;
	{8'd50,8'd181} : s = 231;
	{8'd50,8'd182} : s = 232;
	{8'd50,8'd183} : s = 233;
	{8'd50,8'd184} : s = 234;
	{8'd50,8'd185} : s = 235;
	{8'd50,8'd186} : s = 236;
	{8'd50,8'd187} : s = 237;
	{8'd50,8'd188} : s = 238;
	{8'd50,8'd189} : s = 239;
	{8'd50,8'd190} : s = 240;
	{8'd50,8'd191} : s = 241;
	{8'd50,8'd192} : s = 242;
	{8'd50,8'd193} : s = 243;
	{8'd50,8'd194} : s = 244;
	{8'd50,8'd195} : s = 245;
	{8'd50,8'd196} : s = 246;
	{8'd50,8'd197} : s = 247;
	{8'd50,8'd198} : s = 248;
	{8'd50,8'd199} : s = 249;
	{8'd50,8'd200} : s = 250;
	{8'd50,8'd201} : s = 251;
	{8'd50,8'd202} : s = 252;
	{8'd50,8'd203} : s = 253;
	{8'd50,8'd204} : s = 254;
	{8'd50,8'd205} : s = 255;
	{8'd50,8'd206} : s = 256;
	{8'd50,8'd207} : s = 257;
	{8'd50,8'd208} : s = 258;
	{8'd50,8'd209} : s = 259;
	{8'd50,8'd210} : s = 260;
	{8'd50,8'd211} : s = 261;
	{8'd50,8'd212} : s = 262;
	{8'd50,8'd213} : s = 263;
	{8'd50,8'd214} : s = 264;
	{8'd50,8'd215} : s = 265;
	{8'd50,8'd216} : s = 266;
	{8'd50,8'd217} : s = 267;
	{8'd50,8'd218} : s = 268;
	{8'd50,8'd219} : s = 269;
	{8'd50,8'd220} : s = 270;
	{8'd50,8'd221} : s = 271;
	{8'd50,8'd222} : s = 272;
	{8'd50,8'd223} : s = 273;
	{8'd50,8'd224} : s = 274;
	{8'd50,8'd225} : s = 275;
	{8'd50,8'd226} : s = 276;
	{8'd50,8'd227} : s = 277;
	{8'd50,8'd228} : s = 278;
	{8'd50,8'd229} : s = 279;
	{8'd50,8'd230} : s = 280;
	{8'd50,8'd231} : s = 281;
	{8'd50,8'd232} : s = 282;
	{8'd50,8'd233} : s = 283;
	{8'd50,8'd234} : s = 284;
	{8'd50,8'd235} : s = 285;
	{8'd50,8'd236} : s = 286;
	{8'd50,8'd237} : s = 287;
	{8'd50,8'd238} : s = 288;
	{8'd50,8'd239} : s = 289;
	{8'd50,8'd240} : s = 290;
	{8'd50,8'd241} : s = 291;
	{8'd50,8'd242} : s = 292;
	{8'd50,8'd243} : s = 293;
	{8'd50,8'd244} : s = 294;
	{8'd50,8'd245} : s = 295;
	{8'd50,8'd246} : s = 296;
	{8'd50,8'd247} : s = 297;
	{8'd50,8'd248} : s = 298;
	{8'd50,8'd249} : s = 299;
	{8'd50,8'd250} : s = 300;
	{8'd50,8'd251} : s = 301;
	{8'd50,8'd252} : s = 302;
	{8'd50,8'd253} : s = 303;
	{8'd50,8'd254} : s = 304;
	{8'd50,8'd255} : s = 305;
	{8'd51,8'd0} : s = 51;
	{8'd51,8'd1} : s = 52;
	{8'd51,8'd2} : s = 53;
	{8'd51,8'd3} : s = 54;
	{8'd51,8'd4} : s = 55;
	{8'd51,8'd5} : s = 56;
	{8'd51,8'd6} : s = 57;
	{8'd51,8'd7} : s = 58;
	{8'd51,8'd8} : s = 59;
	{8'd51,8'd9} : s = 60;
	{8'd51,8'd10} : s = 61;
	{8'd51,8'd11} : s = 62;
	{8'd51,8'd12} : s = 63;
	{8'd51,8'd13} : s = 64;
	{8'd51,8'd14} : s = 65;
	{8'd51,8'd15} : s = 66;
	{8'd51,8'd16} : s = 67;
	{8'd51,8'd17} : s = 68;
	{8'd51,8'd18} : s = 69;
	{8'd51,8'd19} : s = 70;
	{8'd51,8'd20} : s = 71;
	{8'd51,8'd21} : s = 72;
	{8'd51,8'd22} : s = 73;
	{8'd51,8'd23} : s = 74;
	{8'd51,8'd24} : s = 75;
	{8'd51,8'd25} : s = 76;
	{8'd51,8'd26} : s = 77;
	{8'd51,8'd27} : s = 78;
	{8'd51,8'd28} : s = 79;
	{8'd51,8'd29} : s = 80;
	{8'd51,8'd30} : s = 81;
	{8'd51,8'd31} : s = 82;
	{8'd51,8'd32} : s = 83;
	{8'd51,8'd33} : s = 84;
	{8'd51,8'd34} : s = 85;
	{8'd51,8'd35} : s = 86;
	{8'd51,8'd36} : s = 87;
	{8'd51,8'd37} : s = 88;
	{8'd51,8'd38} : s = 89;
	{8'd51,8'd39} : s = 90;
	{8'd51,8'd40} : s = 91;
	{8'd51,8'd41} : s = 92;
	{8'd51,8'd42} : s = 93;
	{8'd51,8'd43} : s = 94;
	{8'd51,8'd44} : s = 95;
	{8'd51,8'd45} : s = 96;
	{8'd51,8'd46} : s = 97;
	{8'd51,8'd47} : s = 98;
	{8'd51,8'd48} : s = 99;
	{8'd51,8'd49} : s = 100;
	{8'd51,8'd50} : s = 101;
	{8'd51,8'd51} : s = 102;
	{8'd51,8'd52} : s = 103;
	{8'd51,8'd53} : s = 104;
	{8'd51,8'd54} : s = 105;
	{8'd51,8'd55} : s = 106;
	{8'd51,8'd56} : s = 107;
	{8'd51,8'd57} : s = 108;
	{8'd51,8'd58} : s = 109;
	{8'd51,8'd59} : s = 110;
	{8'd51,8'd60} : s = 111;
	{8'd51,8'd61} : s = 112;
	{8'd51,8'd62} : s = 113;
	{8'd51,8'd63} : s = 114;
	{8'd51,8'd64} : s = 115;
	{8'd51,8'd65} : s = 116;
	{8'd51,8'd66} : s = 117;
	{8'd51,8'd67} : s = 118;
	{8'd51,8'd68} : s = 119;
	{8'd51,8'd69} : s = 120;
	{8'd51,8'd70} : s = 121;
	{8'd51,8'd71} : s = 122;
	{8'd51,8'd72} : s = 123;
	{8'd51,8'd73} : s = 124;
	{8'd51,8'd74} : s = 125;
	{8'd51,8'd75} : s = 126;
	{8'd51,8'd76} : s = 127;
	{8'd51,8'd77} : s = 128;
	{8'd51,8'd78} : s = 129;
	{8'd51,8'd79} : s = 130;
	{8'd51,8'd80} : s = 131;
	{8'd51,8'd81} : s = 132;
	{8'd51,8'd82} : s = 133;
	{8'd51,8'd83} : s = 134;
	{8'd51,8'd84} : s = 135;
	{8'd51,8'd85} : s = 136;
	{8'd51,8'd86} : s = 137;
	{8'd51,8'd87} : s = 138;
	{8'd51,8'd88} : s = 139;
	{8'd51,8'd89} : s = 140;
	{8'd51,8'd90} : s = 141;
	{8'd51,8'd91} : s = 142;
	{8'd51,8'd92} : s = 143;
	{8'd51,8'd93} : s = 144;
	{8'd51,8'd94} : s = 145;
	{8'd51,8'd95} : s = 146;
	{8'd51,8'd96} : s = 147;
	{8'd51,8'd97} : s = 148;
	{8'd51,8'd98} : s = 149;
	{8'd51,8'd99} : s = 150;
	{8'd51,8'd100} : s = 151;
	{8'd51,8'd101} : s = 152;
	{8'd51,8'd102} : s = 153;
	{8'd51,8'd103} : s = 154;
	{8'd51,8'd104} : s = 155;
	{8'd51,8'd105} : s = 156;
	{8'd51,8'd106} : s = 157;
	{8'd51,8'd107} : s = 158;
	{8'd51,8'd108} : s = 159;
	{8'd51,8'd109} : s = 160;
	{8'd51,8'd110} : s = 161;
	{8'd51,8'd111} : s = 162;
	{8'd51,8'd112} : s = 163;
	{8'd51,8'd113} : s = 164;
	{8'd51,8'd114} : s = 165;
	{8'd51,8'd115} : s = 166;
	{8'd51,8'd116} : s = 167;
	{8'd51,8'd117} : s = 168;
	{8'd51,8'd118} : s = 169;
	{8'd51,8'd119} : s = 170;
	{8'd51,8'd120} : s = 171;
	{8'd51,8'd121} : s = 172;
	{8'd51,8'd122} : s = 173;
	{8'd51,8'd123} : s = 174;
	{8'd51,8'd124} : s = 175;
	{8'd51,8'd125} : s = 176;
	{8'd51,8'd126} : s = 177;
	{8'd51,8'd127} : s = 178;
	{8'd51,8'd128} : s = 179;
	{8'd51,8'd129} : s = 180;
	{8'd51,8'd130} : s = 181;
	{8'd51,8'd131} : s = 182;
	{8'd51,8'd132} : s = 183;
	{8'd51,8'd133} : s = 184;
	{8'd51,8'd134} : s = 185;
	{8'd51,8'd135} : s = 186;
	{8'd51,8'd136} : s = 187;
	{8'd51,8'd137} : s = 188;
	{8'd51,8'd138} : s = 189;
	{8'd51,8'd139} : s = 190;
	{8'd51,8'd140} : s = 191;
	{8'd51,8'd141} : s = 192;
	{8'd51,8'd142} : s = 193;
	{8'd51,8'd143} : s = 194;
	{8'd51,8'd144} : s = 195;
	{8'd51,8'd145} : s = 196;
	{8'd51,8'd146} : s = 197;
	{8'd51,8'd147} : s = 198;
	{8'd51,8'd148} : s = 199;
	{8'd51,8'd149} : s = 200;
	{8'd51,8'd150} : s = 201;
	{8'd51,8'd151} : s = 202;
	{8'd51,8'd152} : s = 203;
	{8'd51,8'd153} : s = 204;
	{8'd51,8'd154} : s = 205;
	{8'd51,8'd155} : s = 206;
	{8'd51,8'd156} : s = 207;
	{8'd51,8'd157} : s = 208;
	{8'd51,8'd158} : s = 209;
	{8'd51,8'd159} : s = 210;
	{8'd51,8'd160} : s = 211;
	{8'd51,8'd161} : s = 212;
	{8'd51,8'd162} : s = 213;
	{8'd51,8'd163} : s = 214;
	{8'd51,8'd164} : s = 215;
	{8'd51,8'd165} : s = 216;
	{8'd51,8'd166} : s = 217;
	{8'd51,8'd167} : s = 218;
	{8'd51,8'd168} : s = 219;
	{8'd51,8'd169} : s = 220;
	{8'd51,8'd170} : s = 221;
	{8'd51,8'd171} : s = 222;
	{8'd51,8'd172} : s = 223;
	{8'd51,8'd173} : s = 224;
	{8'd51,8'd174} : s = 225;
	{8'd51,8'd175} : s = 226;
	{8'd51,8'd176} : s = 227;
	{8'd51,8'd177} : s = 228;
	{8'd51,8'd178} : s = 229;
	{8'd51,8'd179} : s = 230;
	{8'd51,8'd180} : s = 231;
	{8'd51,8'd181} : s = 232;
	{8'd51,8'd182} : s = 233;
	{8'd51,8'd183} : s = 234;
	{8'd51,8'd184} : s = 235;
	{8'd51,8'd185} : s = 236;
	{8'd51,8'd186} : s = 237;
	{8'd51,8'd187} : s = 238;
	{8'd51,8'd188} : s = 239;
	{8'd51,8'd189} : s = 240;
	{8'd51,8'd190} : s = 241;
	{8'd51,8'd191} : s = 242;
	{8'd51,8'd192} : s = 243;
	{8'd51,8'd193} : s = 244;
	{8'd51,8'd194} : s = 245;
	{8'd51,8'd195} : s = 246;
	{8'd51,8'd196} : s = 247;
	{8'd51,8'd197} : s = 248;
	{8'd51,8'd198} : s = 249;
	{8'd51,8'd199} : s = 250;
	{8'd51,8'd200} : s = 251;
	{8'd51,8'd201} : s = 252;
	{8'd51,8'd202} : s = 253;
	{8'd51,8'd203} : s = 254;
	{8'd51,8'd204} : s = 255;
	{8'd51,8'd205} : s = 256;
	{8'd51,8'd206} : s = 257;
	{8'd51,8'd207} : s = 258;
	{8'd51,8'd208} : s = 259;
	{8'd51,8'd209} : s = 260;
	{8'd51,8'd210} : s = 261;
	{8'd51,8'd211} : s = 262;
	{8'd51,8'd212} : s = 263;
	{8'd51,8'd213} : s = 264;
	{8'd51,8'd214} : s = 265;
	{8'd51,8'd215} : s = 266;
	{8'd51,8'd216} : s = 267;
	{8'd51,8'd217} : s = 268;
	{8'd51,8'd218} : s = 269;
	{8'd51,8'd219} : s = 270;
	{8'd51,8'd220} : s = 271;
	{8'd51,8'd221} : s = 272;
	{8'd51,8'd222} : s = 273;
	{8'd51,8'd223} : s = 274;
	{8'd51,8'd224} : s = 275;
	{8'd51,8'd225} : s = 276;
	{8'd51,8'd226} : s = 277;
	{8'd51,8'd227} : s = 278;
	{8'd51,8'd228} : s = 279;
	{8'd51,8'd229} : s = 280;
	{8'd51,8'd230} : s = 281;
	{8'd51,8'd231} : s = 282;
	{8'd51,8'd232} : s = 283;
	{8'd51,8'd233} : s = 284;
	{8'd51,8'd234} : s = 285;
	{8'd51,8'd235} : s = 286;
	{8'd51,8'd236} : s = 287;
	{8'd51,8'd237} : s = 288;
	{8'd51,8'd238} : s = 289;
	{8'd51,8'd239} : s = 290;
	{8'd51,8'd240} : s = 291;
	{8'd51,8'd241} : s = 292;
	{8'd51,8'd242} : s = 293;
	{8'd51,8'd243} : s = 294;
	{8'd51,8'd244} : s = 295;
	{8'd51,8'd245} : s = 296;
	{8'd51,8'd246} : s = 297;
	{8'd51,8'd247} : s = 298;
	{8'd51,8'd248} : s = 299;
	{8'd51,8'd249} : s = 300;
	{8'd51,8'd250} : s = 301;
	{8'd51,8'd251} : s = 302;
	{8'd51,8'd252} : s = 303;
	{8'd51,8'd253} : s = 304;
	{8'd51,8'd254} : s = 305;
	{8'd51,8'd255} : s = 306;
	{8'd52,8'd0} : s = 52;
	{8'd52,8'd1} : s = 53;
	{8'd52,8'd2} : s = 54;
	{8'd52,8'd3} : s = 55;
	{8'd52,8'd4} : s = 56;
	{8'd52,8'd5} : s = 57;
	{8'd52,8'd6} : s = 58;
	{8'd52,8'd7} : s = 59;
	{8'd52,8'd8} : s = 60;
	{8'd52,8'd9} : s = 61;
	{8'd52,8'd10} : s = 62;
	{8'd52,8'd11} : s = 63;
	{8'd52,8'd12} : s = 64;
	{8'd52,8'd13} : s = 65;
	{8'd52,8'd14} : s = 66;
	{8'd52,8'd15} : s = 67;
	{8'd52,8'd16} : s = 68;
	{8'd52,8'd17} : s = 69;
	{8'd52,8'd18} : s = 70;
	{8'd52,8'd19} : s = 71;
	{8'd52,8'd20} : s = 72;
	{8'd52,8'd21} : s = 73;
	{8'd52,8'd22} : s = 74;
	{8'd52,8'd23} : s = 75;
	{8'd52,8'd24} : s = 76;
	{8'd52,8'd25} : s = 77;
	{8'd52,8'd26} : s = 78;
	{8'd52,8'd27} : s = 79;
	{8'd52,8'd28} : s = 80;
	{8'd52,8'd29} : s = 81;
	{8'd52,8'd30} : s = 82;
	{8'd52,8'd31} : s = 83;
	{8'd52,8'd32} : s = 84;
	{8'd52,8'd33} : s = 85;
	{8'd52,8'd34} : s = 86;
	{8'd52,8'd35} : s = 87;
	{8'd52,8'd36} : s = 88;
	{8'd52,8'd37} : s = 89;
	{8'd52,8'd38} : s = 90;
	{8'd52,8'd39} : s = 91;
	{8'd52,8'd40} : s = 92;
	{8'd52,8'd41} : s = 93;
	{8'd52,8'd42} : s = 94;
	{8'd52,8'd43} : s = 95;
	{8'd52,8'd44} : s = 96;
	{8'd52,8'd45} : s = 97;
	{8'd52,8'd46} : s = 98;
	{8'd52,8'd47} : s = 99;
	{8'd52,8'd48} : s = 100;
	{8'd52,8'd49} : s = 101;
	{8'd52,8'd50} : s = 102;
	{8'd52,8'd51} : s = 103;
	{8'd52,8'd52} : s = 104;
	{8'd52,8'd53} : s = 105;
	{8'd52,8'd54} : s = 106;
	{8'd52,8'd55} : s = 107;
	{8'd52,8'd56} : s = 108;
	{8'd52,8'd57} : s = 109;
	{8'd52,8'd58} : s = 110;
	{8'd52,8'd59} : s = 111;
	{8'd52,8'd60} : s = 112;
	{8'd52,8'd61} : s = 113;
	{8'd52,8'd62} : s = 114;
	{8'd52,8'd63} : s = 115;
	{8'd52,8'd64} : s = 116;
	{8'd52,8'd65} : s = 117;
	{8'd52,8'd66} : s = 118;
	{8'd52,8'd67} : s = 119;
	{8'd52,8'd68} : s = 120;
	{8'd52,8'd69} : s = 121;
	{8'd52,8'd70} : s = 122;
	{8'd52,8'd71} : s = 123;
	{8'd52,8'd72} : s = 124;
	{8'd52,8'd73} : s = 125;
	{8'd52,8'd74} : s = 126;
	{8'd52,8'd75} : s = 127;
	{8'd52,8'd76} : s = 128;
	{8'd52,8'd77} : s = 129;
	{8'd52,8'd78} : s = 130;
	{8'd52,8'd79} : s = 131;
	{8'd52,8'd80} : s = 132;
	{8'd52,8'd81} : s = 133;
	{8'd52,8'd82} : s = 134;
	{8'd52,8'd83} : s = 135;
	{8'd52,8'd84} : s = 136;
	{8'd52,8'd85} : s = 137;
	{8'd52,8'd86} : s = 138;
	{8'd52,8'd87} : s = 139;
	{8'd52,8'd88} : s = 140;
	{8'd52,8'd89} : s = 141;
	{8'd52,8'd90} : s = 142;
	{8'd52,8'd91} : s = 143;
	{8'd52,8'd92} : s = 144;
	{8'd52,8'd93} : s = 145;
	{8'd52,8'd94} : s = 146;
	{8'd52,8'd95} : s = 147;
	{8'd52,8'd96} : s = 148;
	{8'd52,8'd97} : s = 149;
	{8'd52,8'd98} : s = 150;
	{8'd52,8'd99} : s = 151;
	{8'd52,8'd100} : s = 152;
	{8'd52,8'd101} : s = 153;
	{8'd52,8'd102} : s = 154;
	{8'd52,8'd103} : s = 155;
	{8'd52,8'd104} : s = 156;
	{8'd52,8'd105} : s = 157;
	{8'd52,8'd106} : s = 158;
	{8'd52,8'd107} : s = 159;
	{8'd52,8'd108} : s = 160;
	{8'd52,8'd109} : s = 161;
	{8'd52,8'd110} : s = 162;
	{8'd52,8'd111} : s = 163;
	{8'd52,8'd112} : s = 164;
	{8'd52,8'd113} : s = 165;
	{8'd52,8'd114} : s = 166;
	{8'd52,8'd115} : s = 167;
	{8'd52,8'd116} : s = 168;
	{8'd52,8'd117} : s = 169;
	{8'd52,8'd118} : s = 170;
	{8'd52,8'd119} : s = 171;
	{8'd52,8'd120} : s = 172;
	{8'd52,8'd121} : s = 173;
	{8'd52,8'd122} : s = 174;
	{8'd52,8'd123} : s = 175;
	{8'd52,8'd124} : s = 176;
	{8'd52,8'd125} : s = 177;
	{8'd52,8'd126} : s = 178;
	{8'd52,8'd127} : s = 179;
	{8'd52,8'd128} : s = 180;
	{8'd52,8'd129} : s = 181;
	{8'd52,8'd130} : s = 182;
	{8'd52,8'd131} : s = 183;
	{8'd52,8'd132} : s = 184;
	{8'd52,8'd133} : s = 185;
	{8'd52,8'd134} : s = 186;
	{8'd52,8'd135} : s = 187;
	{8'd52,8'd136} : s = 188;
	{8'd52,8'd137} : s = 189;
	{8'd52,8'd138} : s = 190;
	{8'd52,8'd139} : s = 191;
	{8'd52,8'd140} : s = 192;
	{8'd52,8'd141} : s = 193;
	{8'd52,8'd142} : s = 194;
	{8'd52,8'd143} : s = 195;
	{8'd52,8'd144} : s = 196;
	{8'd52,8'd145} : s = 197;
	{8'd52,8'd146} : s = 198;
	{8'd52,8'd147} : s = 199;
	{8'd52,8'd148} : s = 200;
	{8'd52,8'd149} : s = 201;
	{8'd52,8'd150} : s = 202;
	{8'd52,8'd151} : s = 203;
	{8'd52,8'd152} : s = 204;
	{8'd52,8'd153} : s = 205;
	{8'd52,8'd154} : s = 206;
	{8'd52,8'd155} : s = 207;
	{8'd52,8'd156} : s = 208;
	{8'd52,8'd157} : s = 209;
	{8'd52,8'd158} : s = 210;
	{8'd52,8'd159} : s = 211;
	{8'd52,8'd160} : s = 212;
	{8'd52,8'd161} : s = 213;
	{8'd52,8'd162} : s = 214;
	{8'd52,8'd163} : s = 215;
	{8'd52,8'd164} : s = 216;
	{8'd52,8'd165} : s = 217;
	{8'd52,8'd166} : s = 218;
	{8'd52,8'd167} : s = 219;
	{8'd52,8'd168} : s = 220;
	{8'd52,8'd169} : s = 221;
	{8'd52,8'd170} : s = 222;
	{8'd52,8'd171} : s = 223;
	{8'd52,8'd172} : s = 224;
	{8'd52,8'd173} : s = 225;
	{8'd52,8'd174} : s = 226;
	{8'd52,8'd175} : s = 227;
	{8'd52,8'd176} : s = 228;
	{8'd52,8'd177} : s = 229;
	{8'd52,8'd178} : s = 230;
	{8'd52,8'd179} : s = 231;
	{8'd52,8'd180} : s = 232;
	{8'd52,8'd181} : s = 233;
	{8'd52,8'd182} : s = 234;
	{8'd52,8'd183} : s = 235;
	{8'd52,8'd184} : s = 236;
	{8'd52,8'd185} : s = 237;
	{8'd52,8'd186} : s = 238;
	{8'd52,8'd187} : s = 239;
	{8'd52,8'd188} : s = 240;
	{8'd52,8'd189} : s = 241;
	{8'd52,8'd190} : s = 242;
	{8'd52,8'd191} : s = 243;
	{8'd52,8'd192} : s = 244;
	{8'd52,8'd193} : s = 245;
	{8'd52,8'd194} : s = 246;
	{8'd52,8'd195} : s = 247;
	{8'd52,8'd196} : s = 248;
	{8'd52,8'd197} : s = 249;
	{8'd52,8'd198} : s = 250;
	{8'd52,8'd199} : s = 251;
	{8'd52,8'd200} : s = 252;
	{8'd52,8'd201} : s = 253;
	{8'd52,8'd202} : s = 254;
	{8'd52,8'd203} : s = 255;
	{8'd52,8'd204} : s = 256;
	{8'd52,8'd205} : s = 257;
	{8'd52,8'd206} : s = 258;
	{8'd52,8'd207} : s = 259;
	{8'd52,8'd208} : s = 260;
	{8'd52,8'd209} : s = 261;
	{8'd52,8'd210} : s = 262;
	{8'd52,8'd211} : s = 263;
	{8'd52,8'd212} : s = 264;
	{8'd52,8'd213} : s = 265;
	{8'd52,8'd214} : s = 266;
	{8'd52,8'd215} : s = 267;
	{8'd52,8'd216} : s = 268;
	{8'd52,8'd217} : s = 269;
	{8'd52,8'd218} : s = 270;
	{8'd52,8'd219} : s = 271;
	{8'd52,8'd220} : s = 272;
	{8'd52,8'd221} : s = 273;
	{8'd52,8'd222} : s = 274;
	{8'd52,8'd223} : s = 275;
	{8'd52,8'd224} : s = 276;
	{8'd52,8'd225} : s = 277;
	{8'd52,8'd226} : s = 278;
	{8'd52,8'd227} : s = 279;
	{8'd52,8'd228} : s = 280;
	{8'd52,8'd229} : s = 281;
	{8'd52,8'd230} : s = 282;
	{8'd52,8'd231} : s = 283;
	{8'd52,8'd232} : s = 284;
	{8'd52,8'd233} : s = 285;
	{8'd52,8'd234} : s = 286;
	{8'd52,8'd235} : s = 287;
	{8'd52,8'd236} : s = 288;
	{8'd52,8'd237} : s = 289;
	{8'd52,8'd238} : s = 290;
	{8'd52,8'd239} : s = 291;
	{8'd52,8'd240} : s = 292;
	{8'd52,8'd241} : s = 293;
	{8'd52,8'd242} : s = 294;
	{8'd52,8'd243} : s = 295;
	{8'd52,8'd244} : s = 296;
	{8'd52,8'd245} : s = 297;
	{8'd52,8'd246} : s = 298;
	{8'd52,8'd247} : s = 299;
	{8'd52,8'd248} : s = 300;
	{8'd52,8'd249} : s = 301;
	{8'd52,8'd250} : s = 302;
	{8'd52,8'd251} : s = 303;
	{8'd52,8'd252} : s = 304;
	{8'd52,8'd253} : s = 305;
	{8'd52,8'd254} : s = 306;
	{8'd52,8'd255} : s = 307;
	{8'd53,8'd0} : s = 53;
	{8'd53,8'd1} : s = 54;
	{8'd53,8'd2} : s = 55;
	{8'd53,8'd3} : s = 56;
	{8'd53,8'd4} : s = 57;
	{8'd53,8'd5} : s = 58;
	{8'd53,8'd6} : s = 59;
	{8'd53,8'd7} : s = 60;
	{8'd53,8'd8} : s = 61;
	{8'd53,8'd9} : s = 62;
	{8'd53,8'd10} : s = 63;
	{8'd53,8'd11} : s = 64;
	{8'd53,8'd12} : s = 65;
	{8'd53,8'd13} : s = 66;
	{8'd53,8'd14} : s = 67;
	{8'd53,8'd15} : s = 68;
	{8'd53,8'd16} : s = 69;
	{8'd53,8'd17} : s = 70;
	{8'd53,8'd18} : s = 71;
	{8'd53,8'd19} : s = 72;
	{8'd53,8'd20} : s = 73;
	{8'd53,8'd21} : s = 74;
	{8'd53,8'd22} : s = 75;
	{8'd53,8'd23} : s = 76;
	{8'd53,8'd24} : s = 77;
	{8'd53,8'd25} : s = 78;
	{8'd53,8'd26} : s = 79;
	{8'd53,8'd27} : s = 80;
	{8'd53,8'd28} : s = 81;
	{8'd53,8'd29} : s = 82;
	{8'd53,8'd30} : s = 83;
	{8'd53,8'd31} : s = 84;
	{8'd53,8'd32} : s = 85;
	{8'd53,8'd33} : s = 86;
	{8'd53,8'd34} : s = 87;
	{8'd53,8'd35} : s = 88;
	{8'd53,8'd36} : s = 89;
	{8'd53,8'd37} : s = 90;
	{8'd53,8'd38} : s = 91;
	{8'd53,8'd39} : s = 92;
	{8'd53,8'd40} : s = 93;
	{8'd53,8'd41} : s = 94;
	{8'd53,8'd42} : s = 95;
	{8'd53,8'd43} : s = 96;
	{8'd53,8'd44} : s = 97;
	{8'd53,8'd45} : s = 98;
	{8'd53,8'd46} : s = 99;
	{8'd53,8'd47} : s = 100;
	{8'd53,8'd48} : s = 101;
	{8'd53,8'd49} : s = 102;
	{8'd53,8'd50} : s = 103;
	{8'd53,8'd51} : s = 104;
	{8'd53,8'd52} : s = 105;
	{8'd53,8'd53} : s = 106;
	{8'd53,8'd54} : s = 107;
	{8'd53,8'd55} : s = 108;
	{8'd53,8'd56} : s = 109;
	{8'd53,8'd57} : s = 110;
	{8'd53,8'd58} : s = 111;
	{8'd53,8'd59} : s = 112;
	{8'd53,8'd60} : s = 113;
	{8'd53,8'd61} : s = 114;
	{8'd53,8'd62} : s = 115;
	{8'd53,8'd63} : s = 116;
	{8'd53,8'd64} : s = 117;
	{8'd53,8'd65} : s = 118;
	{8'd53,8'd66} : s = 119;
	{8'd53,8'd67} : s = 120;
	{8'd53,8'd68} : s = 121;
	{8'd53,8'd69} : s = 122;
	{8'd53,8'd70} : s = 123;
	{8'd53,8'd71} : s = 124;
	{8'd53,8'd72} : s = 125;
	{8'd53,8'd73} : s = 126;
	{8'd53,8'd74} : s = 127;
	{8'd53,8'd75} : s = 128;
	{8'd53,8'd76} : s = 129;
	{8'd53,8'd77} : s = 130;
	{8'd53,8'd78} : s = 131;
	{8'd53,8'd79} : s = 132;
	{8'd53,8'd80} : s = 133;
	{8'd53,8'd81} : s = 134;
	{8'd53,8'd82} : s = 135;
	{8'd53,8'd83} : s = 136;
	{8'd53,8'd84} : s = 137;
	{8'd53,8'd85} : s = 138;
	{8'd53,8'd86} : s = 139;
	{8'd53,8'd87} : s = 140;
	{8'd53,8'd88} : s = 141;
	{8'd53,8'd89} : s = 142;
	{8'd53,8'd90} : s = 143;
	{8'd53,8'd91} : s = 144;
	{8'd53,8'd92} : s = 145;
	{8'd53,8'd93} : s = 146;
	{8'd53,8'd94} : s = 147;
	{8'd53,8'd95} : s = 148;
	{8'd53,8'd96} : s = 149;
	{8'd53,8'd97} : s = 150;
	{8'd53,8'd98} : s = 151;
	{8'd53,8'd99} : s = 152;
	{8'd53,8'd100} : s = 153;
	{8'd53,8'd101} : s = 154;
	{8'd53,8'd102} : s = 155;
	{8'd53,8'd103} : s = 156;
	{8'd53,8'd104} : s = 157;
	{8'd53,8'd105} : s = 158;
	{8'd53,8'd106} : s = 159;
	{8'd53,8'd107} : s = 160;
	{8'd53,8'd108} : s = 161;
	{8'd53,8'd109} : s = 162;
	{8'd53,8'd110} : s = 163;
	{8'd53,8'd111} : s = 164;
	{8'd53,8'd112} : s = 165;
	{8'd53,8'd113} : s = 166;
	{8'd53,8'd114} : s = 167;
	{8'd53,8'd115} : s = 168;
	{8'd53,8'd116} : s = 169;
	{8'd53,8'd117} : s = 170;
	{8'd53,8'd118} : s = 171;
	{8'd53,8'd119} : s = 172;
	{8'd53,8'd120} : s = 173;
	{8'd53,8'd121} : s = 174;
	{8'd53,8'd122} : s = 175;
	{8'd53,8'd123} : s = 176;
	{8'd53,8'd124} : s = 177;
	{8'd53,8'd125} : s = 178;
	{8'd53,8'd126} : s = 179;
	{8'd53,8'd127} : s = 180;
	{8'd53,8'd128} : s = 181;
	{8'd53,8'd129} : s = 182;
	{8'd53,8'd130} : s = 183;
	{8'd53,8'd131} : s = 184;
	{8'd53,8'd132} : s = 185;
	{8'd53,8'd133} : s = 186;
	{8'd53,8'd134} : s = 187;
	{8'd53,8'd135} : s = 188;
	{8'd53,8'd136} : s = 189;
	{8'd53,8'd137} : s = 190;
	{8'd53,8'd138} : s = 191;
	{8'd53,8'd139} : s = 192;
	{8'd53,8'd140} : s = 193;
	{8'd53,8'd141} : s = 194;
	{8'd53,8'd142} : s = 195;
	{8'd53,8'd143} : s = 196;
	{8'd53,8'd144} : s = 197;
	{8'd53,8'd145} : s = 198;
	{8'd53,8'd146} : s = 199;
	{8'd53,8'd147} : s = 200;
	{8'd53,8'd148} : s = 201;
	{8'd53,8'd149} : s = 202;
	{8'd53,8'd150} : s = 203;
	{8'd53,8'd151} : s = 204;
	{8'd53,8'd152} : s = 205;
	{8'd53,8'd153} : s = 206;
	{8'd53,8'd154} : s = 207;
	{8'd53,8'd155} : s = 208;
	{8'd53,8'd156} : s = 209;
	{8'd53,8'd157} : s = 210;
	{8'd53,8'd158} : s = 211;
	{8'd53,8'd159} : s = 212;
	{8'd53,8'd160} : s = 213;
	{8'd53,8'd161} : s = 214;
	{8'd53,8'd162} : s = 215;
	{8'd53,8'd163} : s = 216;
	{8'd53,8'd164} : s = 217;
	{8'd53,8'd165} : s = 218;
	{8'd53,8'd166} : s = 219;
	{8'd53,8'd167} : s = 220;
	{8'd53,8'd168} : s = 221;
	{8'd53,8'd169} : s = 222;
	{8'd53,8'd170} : s = 223;
	{8'd53,8'd171} : s = 224;
	{8'd53,8'd172} : s = 225;
	{8'd53,8'd173} : s = 226;
	{8'd53,8'd174} : s = 227;
	{8'd53,8'd175} : s = 228;
	{8'd53,8'd176} : s = 229;
	{8'd53,8'd177} : s = 230;
	{8'd53,8'd178} : s = 231;
	{8'd53,8'd179} : s = 232;
	{8'd53,8'd180} : s = 233;
	{8'd53,8'd181} : s = 234;
	{8'd53,8'd182} : s = 235;
	{8'd53,8'd183} : s = 236;
	{8'd53,8'd184} : s = 237;
	{8'd53,8'd185} : s = 238;
	{8'd53,8'd186} : s = 239;
	{8'd53,8'd187} : s = 240;
	{8'd53,8'd188} : s = 241;
	{8'd53,8'd189} : s = 242;
	{8'd53,8'd190} : s = 243;
	{8'd53,8'd191} : s = 244;
	{8'd53,8'd192} : s = 245;
	{8'd53,8'd193} : s = 246;
	{8'd53,8'd194} : s = 247;
	{8'd53,8'd195} : s = 248;
	{8'd53,8'd196} : s = 249;
	{8'd53,8'd197} : s = 250;
	{8'd53,8'd198} : s = 251;
	{8'd53,8'd199} : s = 252;
	{8'd53,8'd200} : s = 253;
	{8'd53,8'd201} : s = 254;
	{8'd53,8'd202} : s = 255;
	{8'd53,8'd203} : s = 256;
	{8'd53,8'd204} : s = 257;
	{8'd53,8'd205} : s = 258;
	{8'd53,8'd206} : s = 259;
	{8'd53,8'd207} : s = 260;
	{8'd53,8'd208} : s = 261;
	{8'd53,8'd209} : s = 262;
	{8'd53,8'd210} : s = 263;
	{8'd53,8'd211} : s = 264;
	{8'd53,8'd212} : s = 265;
	{8'd53,8'd213} : s = 266;
	{8'd53,8'd214} : s = 267;
	{8'd53,8'd215} : s = 268;
	{8'd53,8'd216} : s = 269;
	{8'd53,8'd217} : s = 270;
	{8'd53,8'd218} : s = 271;
	{8'd53,8'd219} : s = 272;
	{8'd53,8'd220} : s = 273;
	{8'd53,8'd221} : s = 274;
	{8'd53,8'd222} : s = 275;
	{8'd53,8'd223} : s = 276;
	{8'd53,8'd224} : s = 277;
	{8'd53,8'd225} : s = 278;
	{8'd53,8'd226} : s = 279;
	{8'd53,8'd227} : s = 280;
	{8'd53,8'd228} : s = 281;
	{8'd53,8'd229} : s = 282;
	{8'd53,8'd230} : s = 283;
	{8'd53,8'd231} : s = 284;
	{8'd53,8'd232} : s = 285;
	{8'd53,8'd233} : s = 286;
	{8'd53,8'd234} : s = 287;
	{8'd53,8'd235} : s = 288;
	{8'd53,8'd236} : s = 289;
	{8'd53,8'd237} : s = 290;
	{8'd53,8'd238} : s = 291;
	{8'd53,8'd239} : s = 292;
	{8'd53,8'd240} : s = 293;
	{8'd53,8'd241} : s = 294;
	{8'd53,8'd242} : s = 295;
	{8'd53,8'd243} : s = 296;
	{8'd53,8'd244} : s = 297;
	{8'd53,8'd245} : s = 298;
	{8'd53,8'd246} : s = 299;
	{8'd53,8'd247} : s = 300;
	{8'd53,8'd248} : s = 301;
	{8'd53,8'd249} : s = 302;
	{8'd53,8'd250} : s = 303;
	{8'd53,8'd251} : s = 304;
	{8'd53,8'd252} : s = 305;
	{8'd53,8'd253} : s = 306;
	{8'd53,8'd254} : s = 307;
	{8'd53,8'd255} : s = 308;
	{8'd54,8'd0} : s = 54;
	{8'd54,8'd1} : s = 55;
	{8'd54,8'd2} : s = 56;
	{8'd54,8'd3} : s = 57;
	{8'd54,8'd4} : s = 58;
	{8'd54,8'd5} : s = 59;
	{8'd54,8'd6} : s = 60;
	{8'd54,8'd7} : s = 61;
	{8'd54,8'd8} : s = 62;
	{8'd54,8'd9} : s = 63;
	{8'd54,8'd10} : s = 64;
	{8'd54,8'd11} : s = 65;
	{8'd54,8'd12} : s = 66;
	{8'd54,8'd13} : s = 67;
	{8'd54,8'd14} : s = 68;
	{8'd54,8'd15} : s = 69;
	{8'd54,8'd16} : s = 70;
	{8'd54,8'd17} : s = 71;
	{8'd54,8'd18} : s = 72;
	{8'd54,8'd19} : s = 73;
	{8'd54,8'd20} : s = 74;
	{8'd54,8'd21} : s = 75;
	{8'd54,8'd22} : s = 76;
	{8'd54,8'd23} : s = 77;
	{8'd54,8'd24} : s = 78;
	{8'd54,8'd25} : s = 79;
	{8'd54,8'd26} : s = 80;
	{8'd54,8'd27} : s = 81;
	{8'd54,8'd28} : s = 82;
	{8'd54,8'd29} : s = 83;
	{8'd54,8'd30} : s = 84;
	{8'd54,8'd31} : s = 85;
	{8'd54,8'd32} : s = 86;
	{8'd54,8'd33} : s = 87;
	{8'd54,8'd34} : s = 88;
	{8'd54,8'd35} : s = 89;
	{8'd54,8'd36} : s = 90;
	{8'd54,8'd37} : s = 91;
	{8'd54,8'd38} : s = 92;
	{8'd54,8'd39} : s = 93;
	{8'd54,8'd40} : s = 94;
	{8'd54,8'd41} : s = 95;
	{8'd54,8'd42} : s = 96;
	{8'd54,8'd43} : s = 97;
	{8'd54,8'd44} : s = 98;
	{8'd54,8'd45} : s = 99;
	{8'd54,8'd46} : s = 100;
	{8'd54,8'd47} : s = 101;
	{8'd54,8'd48} : s = 102;
	{8'd54,8'd49} : s = 103;
	{8'd54,8'd50} : s = 104;
	{8'd54,8'd51} : s = 105;
	{8'd54,8'd52} : s = 106;
	{8'd54,8'd53} : s = 107;
	{8'd54,8'd54} : s = 108;
	{8'd54,8'd55} : s = 109;
	{8'd54,8'd56} : s = 110;
	{8'd54,8'd57} : s = 111;
	{8'd54,8'd58} : s = 112;
	{8'd54,8'd59} : s = 113;
	{8'd54,8'd60} : s = 114;
	{8'd54,8'd61} : s = 115;
	{8'd54,8'd62} : s = 116;
	{8'd54,8'd63} : s = 117;
	{8'd54,8'd64} : s = 118;
	{8'd54,8'd65} : s = 119;
	{8'd54,8'd66} : s = 120;
	{8'd54,8'd67} : s = 121;
	{8'd54,8'd68} : s = 122;
	{8'd54,8'd69} : s = 123;
	{8'd54,8'd70} : s = 124;
	{8'd54,8'd71} : s = 125;
	{8'd54,8'd72} : s = 126;
	{8'd54,8'd73} : s = 127;
	{8'd54,8'd74} : s = 128;
	{8'd54,8'd75} : s = 129;
	{8'd54,8'd76} : s = 130;
	{8'd54,8'd77} : s = 131;
	{8'd54,8'd78} : s = 132;
	{8'd54,8'd79} : s = 133;
	{8'd54,8'd80} : s = 134;
	{8'd54,8'd81} : s = 135;
	{8'd54,8'd82} : s = 136;
	{8'd54,8'd83} : s = 137;
	{8'd54,8'd84} : s = 138;
	{8'd54,8'd85} : s = 139;
	{8'd54,8'd86} : s = 140;
	{8'd54,8'd87} : s = 141;
	{8'd54,8'd88} : s = 142;
	{8'd54,8'd89} : s = 143;
	{8'd54,8'd90} : s = 144;
	{8'd54,8'd91} : s = 145;
	{8'd54,8'd92} : s = 146;
	{8'd54,8'd93} : s = 147;
	{8'd54,8'd94} : s = 148;
	{8'd54,8'd95} : s = 149;
	{8'd54,8'd96} : s = 150;
	{8'd54,8'd97} : s = 151;
	{8'd54,8'd98} : s = 152;
	{8'd54,8'd99} : s = 153;
	{8'd54,8'd100} : s = 154;
	{8'd54,8'd101} : s = 155;
	{8'd54,8'd102} : s = 156;
	{8'd54,8'd103} : s = 157;
	{8'd54,8'd104} : s = 158;
	{8'd54,8'd105} : s = 159;
	{8'd54,8'd106} : s = 160;
	{8'd54,8'd107} : s = 161;
	{8'd54,8'd108} : s = 162;
	{8'd54,8'd109} : s = 163;
	{8'd54,8'd110} : s = 164;
	{8'd54,8'd111} : s = 165;
	{8'd54,8'd112} : s = 166;
	{8'd54,8'd113} : s = 167;
	{8'd54,8'd114} : s = 168;
	{8'd54,8'd115} : s = 169;
	{8'd54,8'd116} : s = 170;
	{8'd54,8'd117} : s = 171;
	{8'd54,8'd118} : s = 172;
	{8'd54,8'd119} : s = 173;
	{8'd54,8'd120} : s = 174;
	{8'd54,8'd121} : s = 175;
	{8'd54,8'd122} : s = 176;
	{8'd54,8'd123} : s = 177;
	{8'd54,8'd124} : s = 178;
	{8'd54,8'd125} : s = 179;
	{8'd54,8'd126} : s = 180;
	{8'd54,8'd127} : s = 181;
	{8'd54,8'd128} : s = 182;
	{8'd54,8'd129} : s = 183;
	{8'd54,8'd130} : s = 184;
	{8'd54,8'd131} : s = 185;
	{8'd54,8'd132} : s = 186;
	{8'd54,8'd133} : s = 187;
	{8'd54,8'd134} : s = 188;
	{8'd54,8'd135} : s = 189;
	{8'd54,8'd136} : s = 190;
	{8'd54,8'd137} : s = 191;
	{8'd54,8'd138} : s = 192;
	{8'd54,8'd139} : s = 193;
	{8'd54,8'd140} : s = 194;
	{8'd54,8'd141} : s = 195;
	{8'd54,8'd142} : s = 196;
	{8'd54,8'd143} : s = 197;
	{8'd54,8'd144} : s = 198;
	{8'd54,8'd145} : s = 199;
	{8'd54,8'd146} : s = 200;
	{8'd54,8'd147} : s = 201;
	{8'd54,8'd148} : s = 202;
	{8'd54,8'd149} : s = 203;
	{8'd54,8'd150} : s = 204;
	{8'd54,8'd151} : s = 205;
	{8'd54,8'd152} : s = 206;
	{8'd54,8'd153} : s = 207;
	{8'd54,8'd154} : s = 208;
	{8'd54,8'd155} : s = 209;
	{8'd54,8'd156} : s = 210;
	{8'd54,8'd157} : s = 211;
	{8'd54,8'd158} : s = 212;
	{8'd54,8'd159} : s = 213;
	{8'd54,8'd160} : s = 214;
	{8'd54,8'd161} : s = 215;
	{8'd54,8'd162} : s = 216;
	{8'd54,8'd163} : s = 217;
	{8'd54,8'd164} : s = 218;
	{8'd54,8'd165} : s = 219;
	{8'd54,8'd166} : s = 220;
	{8'd54,8'd167} : s = 221;
	{8'd54,8'd168} : s = 222;
	{8'd54,8'd169} : s = 223;
	{8'd54,8'd170} : s = 224;
	{8'd54,8'd171} : s = 225;
	{8'd54,8'd172} : s = 226;
	{8'd54,8'd173} : s = 227;
	{8'd54,8'd174} : s = 228;
	{8'd54,8'd175} : s = 229;
	{8'd54,8'd176} : s = 230;
	{8'd54,8'd177} : s = 231;
	{8'd54,8'd178} : s = 232;
	{8'd54,8'd179} : s = 233;
	{8'd54,8'd180} : s = 234;
	{8'd54,8'd181} : s = 235;
	{8'd54,8'd182} : s = 236;
	{8'd54,8'd183} : s = 237;
	{8'd54,8'd184} : s = 238;
	{8'd54,8'd185} : s = 239;
	{8'd54,8'd186} : s = 240;
	{8'd54,8'd187} : s = 241;
	{8'd54,8'd188} : s = 242;
	{8'd54,8'd189} : s = 243;
	{8'd54,8'd190} : s = 244;
	{8'd54,8'd191} : s = 245;
	{8'd54,8'd192} : s = 246;
	{8'd54,8'd193} : s = 247;
	{8'd54,8'd194} : s = 248;
	{8'd54,8'd195} : s = 249;
	{8'd54,8'd196} : s = 250;
	{8'd54,8'd197} : s = 251;
	{8'd54,8'd198} : s = 252;
	{8'd54,8'd199} : s = 253;
	{8'd54,8'd200} : s = 254;
	{8'd54,8'd201} : s = 255;
	{8'd54,8'd202} : s = 256;
	{8'd54,8'd203} : s = 257;
	{8'd54,8'd204} : s = 258;
	{8'd54,8'd205} : s = 259;
	{8'd54,8'd206} : s = 260;
	{8'd54,8'd207} : s = 261;
	{8'd54,8'd208} : s = 262;
	{8'd54,8'd209} : s = 263;
	{8'd54,8'd210} : s = 264;
	{8'd54,8'd211} : s = 265;
	{8'd54,8'd212} : s = 266;
	{8'd54,8'd213} : s = 267;
	{8'd54,8'd214} : s = 268;
	{8'd54,8'd215} : s = 269;
	{8'd54,8'd216} : s = 270;
	{8'd54,8'd217} : s = 271;
	{8'd54,8'd218} : s = 272;
	{8'd54,8'd219} : s = 273;
	{8'd54,8'd220} : s = 274;
	{8'd54,8'd221} : s = 275;
	{8'd54,8'd222} : s = 276;
	{8'd54,8'd223} : s = 277;
	{8'd54,8'd224} : s = 278;
	{8'd54,8'd225} : s = 279;
	{8'd54,8'd226} : s = 280;
	{8'd54,8'd227} : s = 281;
	{8'd54,8'd228} : s = 282;
	{8'd54,8'd229} : s = 283;
	{8'd54,8'd230} : s = 284;
	{8'd54,8'd231} : s = 285;
	{8'd54,8'd232} : s = 286;
	{8'd54,8'd233} : s = 287;
	{8'd54,8'd234} : s = 288;
	{8'd54,8'd235} : s = 289;
	{8'd54,8'd236} : s = 290;
	{8'd54,8'd237} : s = 291;
	{8'd54,8'd238} : s = 292;
	{8'd54,8'd239} : s = 293;
	{8'd54,8'd240} : s = 294;
	{8'd54,8'd241} : s = 295;
	{8'd54,8'd242} : s = 296;
	{8'd54,8'd243} : s = 297;
	{8'd54,8'd244} : s = 298;
	{8'd54,8'd245} : s = 299;
	{8'd54,8'd246} : s = 300;
	{8'd54,8'd247} : s = 301;
	{8'd54,8'd248} : s = 302;
	{8'd54,8'd249} : s = 303;
	{8'd54,8'd250} : s = 304;
	{8'd54,8'd251} : s = 305;
	{8'd54,8'd252} : s = 306;
	{8'd54,8'd253} : s = 307;
	{8'd54,8'd254} : s = 308;
	{8'd54,8'd255} : s = 309;
	{8'd55,8'd0} : s = 55;
	{8'd55,8'd1} : s = 56;
	{8'd55,8'd2} : s = 57;
	{8'd55,8'd3} : s = 58;
	{8'd55,8'd4} : s = 59;
	{8'd55,8'd5} : s = 60;
	{8'd55,8'd6} : s = 61;
	{8'd55,8'd7} : s = 62;
	{8'd55,8'd8} : s = 63;
	{8'd55,8'd9} : s = 64;
	{8'd55,8'd10} : s = 65;
	{8'd55,8'd11} : s = 66;
	{8'd55,8'd12} : s = 67;
	{8'd55,8'd13} : s = 68;
	{8'd55,8'd14} : s = 69;
	{8'd55,8'd15} : s = 70;
	{8'd55,8'd16} : s = 71;
	{8'd55,8'd17} : s = 72;
	{8'd55,8'd18} : s = 73;
	{8'd55,8'd19} : s = 74;
	{8'd55,8'd20} : s = 75;
	{8'd55,8'd21} : s = 76;
	{8'd55,8'd22} : s = 77;
	{8'd55,8'd23} : s = 78;
	{8'd55,8'd24} : s = 79;
	{8'd55,8'd25} : s = 80;
	{8'd55,8'd26} : s = 81;
	{8'd55,8'd27} : s = 82;
	{8'd55,8'd28} : s = 83;
	{8'd55,8'd29} : s = 84;
	{8'd55,8'd30} : s = 85;
	{8'd55,8'd31} : s = 86;
	{8'd55,8'd32} : s = 87;
	{8'd55,8'd33} : s = 88;
	{8'd55,8'd34} : s = 89;
	{8'd55,8'd35} : s = 90;
	{8'd55,8'd36} : s = 91;
	{8'd55,8'd37} : s = 92;
	{8'd55,8'd38} : s = 93;
	{8'd55,8'd39} : s = 94;
	{8'd55,8'd40} : s = 95;
	{8'd55,8'd41} : s = 96;
	{8'd55,8'd42} : s = 97;
	{8'd55,8'd43} : s = 98;
	{8'd55,8'd44} : s = 99;
	{8'd55,8'd45} : s = 100;
	{8'd55,8'd46} : s = 101;
	{8'd55,8'd47} : s = 102;
	{8'd55,8'd48} : s = 103;
	{8'd55,8'd49} : s = 104;
	{8'd55,8'd50} : s = 105;
	{8'd55,8'd51} : s = 106;
	{8'd55,8'd52} : s = 107;
	{8'd55,8'd53} : s = 108;
	{8'd55,8'd54} : s = 109;
	{8'd55,8'd55} : s = 110;
	{8'd55,8'd56} : s = 111;
	{8'd55,8'd57} : s = 112;
	{8'd55,8'd58} : s = 113;
	{8'd55,8'd59} : s = 114;
	{8'd55,8'd60} : s = 115;
	{8'd55,8'd61} : s = 116;
	{8'd55,8'd62} : s = 117;
	{8'd55,8'd63} : s = 118;
	{8'd55,8'd64} : s = 119;
	{8'd55,8'd65} : s = 120;
	{8'd55,8'd66} : s = 121;
	{8'd55,8'd67} : s = 122;
	{8'd55,8'd68} : s = 123;
	{8'd55,8'd69} : s = 124;
	{8'd55,8'd70} : s = 125;
	{8'd55,8'd71} : s = 126;
	{8'd55,8'd72} : s = 127;
	{8'd55,8'd73} : s = 128;
	{8'd55,8'd74} : s = 129;
	{8'd55,8'd75} : s = 130;
	{8'd55,8'd76} : s = 131;
	{8'd55,8'd77} : s = 132;
	{8'd55,8'd78} : s = 133;
	{8'd55,8'd79} : s = 134;
	{8'd55,8'd80} : s = 135;
	{8'd55,8'd81} : s = 136;
	{8'd55,8'd82} : s = 137;
	{8'd55,8'd83} : s = 138;
	{8'd55,8'd84} : s = 139;
	{8'd55,8'd85} : s = 140;
	{8'd55,8'd86} : s = 141;
	{8'd55,8'd87} : s = 142;
	{8'd55,8'd88} : s = 143;
	{8'd55,8'd89} : s = 144;
	{8'd55,8'd90} : s = 145;
	{8'd55,8'd91} : s = 146;
	{8'd55,8'd92} : s = 147;
	{8'd55,8'd93} : s = 148;
	{8'd55,8'd94} : s = 149;
	{8'd55,8'd95} : s = 150;
	{8'd55,8'd96} : s = 151;
	{8'd55,8'd97} : s = 152;
	{8'd55,8'd98} : s = 153;
	{8'd55,8'd99} : s = 154;
	{8'd55,8'd100} : s = 155;
	{8'd55,8'd101} : s = 156;
	{8'd55,8'd102} : s = 157;
	{8'd55,8'd103} : s = 158;
	{8'd55,8'd104} : s = 159;
	{8'd55,8'd105} : s = 160;
	{8'd55,8'd106} : s = 161;
	{8'd55,8'd107} : s = 162;
	{8'd55,8'd108} : s = 163;
	{8'd55,8'd109} : s = 164;
	{8'd55,8'd110} : s = 165;
	{8'd55,8'd111} : s = 166;
	{8'd55,8'd112} : s = 167;
	{8'd55,8'd113} : s = 168;
	{8'd55,8'd114} : s = 169;
	{8'd55,8'd115} : s = 170;
	{8'd55,8'd116} : s = 171;
	{8'd55,8'd117} : s = 172;
	{8'd55,8'd118} : s = 173;
	{8'd55,8'd119} : s = 174;
	{8'd55,8'd120} : s = 175;
	{8'd55,8'd121} : s = 176;
	{8'd55,8'd122} : s = 177;
	{8'd55,8'd123} : s = 178;
	{8'd55,8'd124} : s = 179;
	{8'd55,8'd125} : s = 180;
	{8'd55,8'd126} : s = 181;
	{8'd55,8'd127} : s = 182;
	{8'd55,8'd128} : s = 183;
	{8'd55,8'd129} : s = 184;
	{8'd55,8'd130} : s = 185;
	{8'd55,8'd131} : s = 186;
	{8'd55,8'd132} : s = 187;
	{8'd55,8'd133} : s = 188;
	{8'd55,8'd134} : s = 189;
	{8'd55,8'd135} : s = 190;
	{8'd55,8'd136} : s = 191;
	{8'd55,8'd137} : s = 192;
	{8'd55,8'd138} : s = 193;
	{8'd55,8'd139} : s = 194;
	{8'd55,8'd140} : s = 195;
	{8'd55,8'd141} : s = 196;
	{8'd55,8'd142} : s = 197;
	{8'd55,8'd143} : s = 198;
	{8'd55,8'd144} : s = 199;
	{8'd55,8'd145} : s = 200;
	{8'd55,8'd146} : s = 201;
	{8'd55,8'd147} : s = 202;
	{8'd55,8'd148} : s = 203;
	{8'd55,8'd149} : s = 204;
	{8'd55,8'd150} : s = 205;
	{8'd55,8'd151} : s = 206;
	{8'd55,8'd152} : s = 207;
	{8'd55,8'd153} : s = 208;
	{8'd55,8'd154} : s = 209;
	{8'd55,8'd155} : s = 210;
	{8'd55,8'd156} : s = 211;
	{8'd55,8'd157} : s = 212;
	{8'd55,8'd158} : s = 213;
	{8'd55,8'd159} : s = 214;
	{8'd55,8'd160} : s = 215;
	{8'd55,8'd161} : s = 216;
	{8'd55,8'd162} : s = 217;
	{8'd55,8'd163} : s = 218;
	{8'd55,8'd164} : s = 219;
	{8'd55,8'd165} : s = 220;
	{8'd55,8'd166} : s = 221;
	{8'd55,8'd167} : s = 222;
	{8'd55,8'd168} : s = 223;
	{8'd55,8'd169} : s = 224;
	{8'd55,8'd170} : s = 225;
	{8'd55,8'd171} : s = 226;
	{8'd55,8'd172} : s = 227;
	{8'd55,8'd173} : s = 228;
	{8'd55,8'd174} : s = 229;
	{8'd55,8'd175} : s = 230;
	{8'd55,8'd176} : s = 231;
	{8'd55,8'd177} : s = 232;
	{8'd55,8'd178} : s = 233;
	{8'd55,8'd179} : s = 234;
	{8'd55,8'd180} : s = 235;
	{8'd55,8'd181} : s = 236;
	{8'd55,8'd182} : s = 237;
	{8'd55,8'd183} : s = 238;
	{8'd55,8'd184} : s = 239;
	{8'd55,8'd185} : s = 240;
	{8'd55,8'd186} : s = 241;
	{8'd55,8'd187} : s = 242;
	{8'd55,8'd188} : s = 243;
	{8'd55,8'd189} : s = 244;
	{8'd55,8'd190} : s = 245;
	{8'd55,8'd191} : s = 246;
	{8'd55,8'd192} : s = 247;
	{8'd55,8'd193} : s = 248;
	{8'd55,8'd194} : s = 249;
	{8'd55,8'd195} : s = 250;
	{8'd55,8'd196} : s = 251;
	{8'd55,8'd197} : s = 252;
	{8'd55,8'd198} : s = 253;
	{8'd55,8'd199} : s = 254;
	{8'd55,8'd200} : s = 255;
	{8'd55,8'd201} : s = 256;
	{8'd55,8'd202} : s = 257;
	{8'd55,8'd203} : s = 258;
	{8'd55,8'd204} : s = 259;
	{8'd55,8'd205} : s = 260;
	{8'd55,8'd206} : s = 261;
	{8'd55,8'd207} : s = 262;
	{8'd55,8'd208} : s = 263;
	{8'd55,8'd209} : s = 264;
	{8'd55,8'd210} : s = 265;
	{8'd55,8'd211} : s = 266;
	{8'd55,8'd212} : s = 267;
	{8'd55,8'd213} : s = 268;
	{8'd55,8'd214} : s = 269;
	{8'd55,8'd215} : s = 270;
	{8'd55,8'd216} : s = 271;
	{8'd55,8'd217} : s = 272;
	{8'd55,8'd218} : s = 273;
	{8'd55,8'd219} : s = 274;
	{8'd55,8'd220} : s = 275;
	{8'd55,8'd221} : s = 276;
	{8'd55,8'd222} : s = 277;
	{8'd55,8'd223} : s = 278;
	{8'd55,8'd224} : s = 279;
	{8'd55,8'd225} : s = 280;
	{8'd55,8'd226} : s = 281;
	{8'd55,8'd227} : s = 282;
	{8'd55,8'd228} : s = 283;
	{8'd55,8'd229} : s = 284;
	{8'd55,8'd230} : s = 285;
	{8'd55,8'd231} : s = 286;
	{8'd55,8'd232} : s = 287;
	{8'd55,8'd233} : s = 288;
	{8'd55,8'd234} : s = 289;
	{8'd55,8'd235} : s = 290;
	{8'd55,8'd236} : s = 291;
	{8'd55,8'd237} : s = 292;
	{8'd55,8'd238} : s = 293;
	{8'd55,8'd239} : s = 294;
	{8'd55,8'd240} : s = 295;
	{8'd55,8'd241} : s = 296;
	{8'd55,8'd242} : s = 297;
	{8'd55,8'd243} : s = 298;
	{8'd55,8'd244} : s = 299;
	{8'd55,8'd245} : s = 300;
	{8'd55,8'd246} : s = 301;
	{8'd55,8'd247} : s = 302;
	{8'd55,8'd248} : s = 303;
	{8'd55,8'd249} : s = 304;
	{8'd55,8'd250} : s = 305;
	{8'd55,8'd251} : s = 306;
	{8'd55,8'd252} : s = 307;
	{8'd55,8'd253} : s = 308;
	{8'd55,8'd254} : s = 309;
	{8'd55,8'd255} : s = 310;
	{8'd56,8'd0} : s = 56;
	{8'd56,8'd1} : s = 57;
	{8'd56,8'd2} : s = 58;
	{8'd56,8'd3} : s = 59;
	{8'd56,8'd4} : s = 60;
	{8'd56,8'd5} : s = 61;
	{8'd56,8'd6} : s = 62;
	{8'd56,8'd7} : s = 63;
	{8'd56,8'd8} : s = 64;
	{8'd56,8'd9} : s = 65;
	{8'd56,8'd10} : s = 66;
	{8'd56,8'd11} : s = 67;
	{8'd56,8'd12} : s = 68;
	{8'd56,8'd13} : s = 69;
	{8'd56,8'd14} : s = 70;
	{8'd56,8'd15} : s = 71;
	{8'd56,8'd16} : s = 72;
	{8'd56,8'd17} : s = 73;
	{8'd56,8'd18} : s = 74;
	{8'd56,8'd19} : s = 75;
	{8'd56,8'd20} : s = 76;
	{8'd56,8'd21} : s = 77;
	{8'd56,8'd22} : s = 78;
	{8'd56,8'd23} : s = 79;
	{8'd56,8'd24} : s = 80;
	{8'd56,8'd25} : s = 81;
	{8'd56,8'd26} : s = 82;
	{8'd56,8'd27} : s = 83;
	{8'd56,8'd28} : s = 84;
	{8'd56,8'd29} : s = 85;
	{8'd56,8'd30} : s = 86;
	{8'd56,8'd31} : s = 87;
	{8'd56,8'd32} : s = 88;
	{8'd56,8'd33} : s = 89;
	{8'd56,8'd34} : s = 90;
	{8'd56,8'd35} : s = 91;
	{8'd56,8'd36} : s = 92;
	{8'd56,8'd37} : s = 93;
	{8'd56,8'd38} : s = 94;
	{8'd56,8'd39} : s = 95;
	{8'd56,8'd40} : s = 96;
	{8'd56,8'd41} : s = 97;
	{8'd56,8'd42} : s = 98;
	{8'd56,8'd43} : s = 99;
	{8'd56,8'd44} : s = 100;
	{8'd56,8'd45} : s = 101;
	{8'd56,8'd46} : s = 102;
	{8'd56,8'd47} : s = 103;
	{8'd56,8'd48} : s = 104;
	{8'd56,8'd49} : s = 105;
	{8'd56,8'd50} : s = 106;
	{8'd56,8'd51} : s = 107;
	{8'd56,8'd52} : s = 108;
	{8'd56,8'd53} : s = 109;
	{8'd56,8'd54} : s = 110;
	{8'd56,8'd55} : s = 111;
	{8'd56,8'd56} : s = 112;
	{8'd56,8'd57} : s = 113;
	{8'd56,8'd58} : s = 114;
	{8'd56,8'd59} : s = 115;
	{8'd56,8'd60} : s = 116;
	{8'd56,8'd61} : s = 117;
	{8'd56,8'd62} : s = 118;
	{8'd56,8'd63} : s = 119;
	{8'd56,8'd64} : s = 120;
	{8'd56,8'd65} : s = 121;
	{8'd56,8'd66} : s = 122;
	{8'd56,8'd67} : s = 123;
	{8'd56,8'd68} : s = 124;
	{8'd56,8'd69} : s = 125;
	{8'd56,8'd70} : s = 126;
	{8'd56,8'd71} : s = 127;
	{8'd56,8'd72} : s = 128;
	{8'd56,8'd73} : s = 129;
	{8'd56,8'd74} : s = 130;
	{8'd56,8'd75} : s = 131;
	{8'd56,8'd76} : s = 132;
	{8'd56,8'd77} : s = 133;
	{8'd56,8'd78} : s = 134;
	{8'd56,8'd79} : s = 135;
	{8'd56,8'd80} : s = 136;
	{8'd56,8'd81} : s = 137;
	{8'd56,8'd82} : s = 138;
	{8'd56,8'd83} : s = 139;
	{8'd56,8'd84} : s = 140;
	{8'd56,8'd85} : s = 141;
	{8'd56,8'd86} : s = 142;
	{8'd56,8'd87} : s = 143;
	{8'd56,8'd88} : s = 144;
	{8'd56,8'd89} : s = 145;
	{8'd56,8'd90} : s = 146;
	{8'd56,8'd91} : s = 147;
	{8'd56,8'd92} : s = 148;
	{8'd56,8'd93} : s = 149;
	{8'd56,8'd94} : s = 150;
	{8'd56,8'd95} : s = 151;
	{8'd56,8'd96} : s = 152;
	{8'd56,8'd97} : s = 153;
	{8'd56,8'd98} : s = 154;
	{8'd56,8'd99} : s = 155;
	{8'd56,8'd100} : s = 156;
	{8'd56,8'd101} : s = 157;
	{8'd56,8'd102} : s = 158;
	{8'd56,8'd103} : s = 159;
	{8'd56,8'd104} : s = 160;
	{8'd56,8'd105} : s = 161;
	{8'd56,8'd106} : s = 162;
	{8'd56,8'd107} : s = 163;
	{8'd56,8'd108} : s = 164;
	{8'd56,8'd109} : s = 165;
	{8'd56,8'd110} : s = 166;
	{8'd56,8'd111} : s = 167;
	{8'd56,8'd112} : s = 168;
	{8'd56,8'd113} : s = 169;
	{8'd56,8'd114} : s = 170;
	{8'd56,8'd115} : s = 171;
	{8'd56,8'd116} : s = 172;
	{8'd56,8'd117} : s = 173;
	{8'd56,8'd118} : s = 174;
	{8'd56,8'd119} : s = 175;
	{8'd56,8'd120} : s = 176;
	{8'd56,8'd121} : s = 177;
	{8'd56,8'd122} : s = 178;
	{8'd56,8'd123} : s = 179;
	{8'd56,8'd124} : s = 180;
	{8'd56,8'd125} : s = 181;
	{8'd56,8'd126} : s = 182;
	{8'd56,8'd127} : s = 183;
	{8'd56,8'd128} : s = 184;
	{8'd56,8'd129} : s = 185;
	{8'd56,8'd130} : s = 186;
	{8'd56,8'd131} : s = 187;
	{8'd56,8'd132} : s = 188;
	{8'd56,8'd133} : s = 189;
	{8'd56,8'd134} : s = 190;
	{8'd56,8'd135} : s = 191;
	{8'd56,8'd136} : s = 192;
	{8'd56,8'd137} : s = 193;
	{8'd56,8'd138} : s = 194;
	{8'd56,8'd139} : s = 195;
	{8'd56,8'd140} : s = 196;
	{8'd56,8'd141} : s = 197;
	{8'd56,8'd142} : s = 198;
	{8'd56,8'd143} : s = 199;
	{8'd56,8'd144} : s = 200;
	{8'd56,8'd145} : s = 201;
	{8'd56,8'd146} : s = 202;
	{8'd56,8'd147} : s = 203;
	{8'd56,8'd148} : s = 204;
	{8'd56,8'd149} : s = 205;
	{8'd56,8'd150} : s = 206;
	{8'd56,8'd151} : s = 207;
	{8'd56,8'd152} : s = 208;
	{8'd56,8'd153} : s = 209;
	{8'd56,8'd154} : s = 210;
	{8'd56,8'd155} : s = 211;
	{8'd56,8'd156} : s = 212;
	{8'd56,8'd157} : s = 213;
	{8'd56,8'd158} : s = 214;
	{8'd56,8'd159} : s = 215;
	{8'd56,8'd160} : s = 216;
	{8'd56,8'd161} : s = 217;
	{8'd56,8'd162} : s = 218;
	{8'd56,8'd163} : s = 219;
	{8'd56,8'd164} : s = 220;
	{8'd56,8'd165} : s = 221;
	{8'd56,8'd166} : s = 222;
	{8'd56,8'd167} : s = 223;
	{8'd56,8'd168} : s = 224;
	{8'd56,8'd169} : s = 225;
	{8'd56,8'd170} : s = 226;
	{8'd56,8'd171} : s = 227;
	{8'd56,8'd172} : s = 228;
	{8'd56,8'd173} : s = 229;
	{8'd56,8'd174} : s = 230;
	{8'd56,8'd175} : s = 231;
	{8'd56,8'd176} : s = 232;
	{8'd56,8'd177} : s = 233;
	{8'd56,8'd178} : s = 234;
	{8'd56,8'd179} : s = 235;
	{8'd56,8'd180} : s = 236;
	{8'd56,8'd181} : s = 237;
	{8'd56,8'd182} : s = 238;
	{8'd56,8'd183} : s = 239;
	{8'd56,8'd184} : s = 240;
	{8'd56,8'd185} : s = 241;
	{8'd56,8'd186} : s = 242;
	{8'd56,8'd187} : s = 243;
	{8'd56,8'd188} : s = 244;
	{8'd56,8'd189} : s = 245;
	{8'd56,8'd190} : s = 246;
	{8'd56,8'd191} : s = 247;
	{8'd56,8'd192} : s = 248;
	{8'd56,8'd193} : s = 249;
	{8'd56,8'd194} : s = 250;
	{8'd56,8'd195} : s = 251;
	{8'd56,8'd196} : s = 252;
	{8'd56,8'd197} : s = 253;
	{8'd56,8'd198} : s = 254;
	{8'd56,8'd199} : s = 255;
	{8'd56,8'd200} : s = 256;
	{8'd56,8'd201} : s = 257;
	{8'd56,8'd202} : s = 258;
	{8'd56,8'd203} : s = 259;
	{8'd56,8'd204} : s = 260;
	{8'd56,8'd205} : s = 261;
	{8'd56,8'd206} : s = 262;
	{8'd56,8'd207} : s = 263;
	{8'd56,8'd208} : s = 264;
	{8'd56,8'd209} : s = 265;
	{8'd56,8'd210} : s = 266;
	{8'd56,8'd211} : s = 267;
	{8'd56,8'd212} : s = 268;
	{8'd56,8'd213} : s = 269;
	{8'd56,8'd214} : s = 270;
	{8'd56,8'd215} : s = 271;
	{8'd56,8'd216} : s = 272;
	{8'd56,8'd217} : s = 273;
	{8'd56,8'd218} : s = 274;
	{8'd56,8'd219} : s = 275;
	{8'd56,8'd220} : s = 276;
	{8'd56,8'd221} : s = 277;
	{8'd56,8'd222} : s = 278;
	{8'd56,8'd223} : s = 279;
	{8'd56,8'd224} : s = 280;
	{8'd56,8'd225} : s = 281;
	{8'd56,8'd226} : s = 282;
	{8'd56,8'd227} : s = 283;
	{8'd56,8'd228} : s = 284;
	{8'd56,8'd229} : s = 285;
	{8'd56,8'd230} : s = 286;
	{8'd56,8'd231} : s = 287;
	{8'd56,8'd232} : s = 288;
	{8'd56,8'd233} : s = 289;
	{8'd56,8'd234} : s = 290;
	{8'd56,8'd235} : s = 291;
	{8'd56,8'd236} : s = 292;
	{8'd56,8'd237} : s = 293;
	{8'd56,8'd238} : s = 294;
	{8'd56,8'd239} : s = 295;
	{8'd56,8'd240} : s = 296;
	{8'd56,8'd241} : s = 297;
	{8'd56,8'd242} : s = 298;
	{8'd56,8'd243} : s = 299;
	{8'd56,8'd244} : s = 300;
	{8'd56,8'd245} : s = 301;
	{8'd56,8'd246} : s = 302;
	{8'd56,8'd247} : s = 303;
	{8'd56,8'd248} : s = 304;
	{8'd56,8'd249} : s = 305;
	{8'd56,8'd250} : s = 306;
	{8'd56,8'd251} : s = 307;
	{8'd56,8'd252} : s = 308;
	{8'd56,8'd253} : s = 309;
	{8'd56,8'd254} : s = 310;
	{8'd56,8'd255} : s = 311;
	{8'd57,8'd0} : s = 57;
	{8'd57,8'd1} : s = 58;
	{8'd57,8'd2} : s = 59;
	{8'd57,8'd3} : s = 60;
	{8'd57,8'd4} : s = 61;
	{8'd57,8'd5} : s = 62;
	{8'd57,8'd6} : s = 63;
	{8'd57,8'd7} : s = 64;
	{8'd57,8'd8} : s = 65;
	{8'd57,8'd9} : s = 66;
	{8'd57,8'd10} : s = 67;
	{8'd57,8'd11} : s = 68;
	{8'd57,8'd12} : s = 69;
	{8'd57,8'd13} : s = 70;
	{8'd57,8'd14} : s = 71;
	{8'd57,8'd15} : s = 72;
	{8'd57,8'd16} : s = 73;
	{8'd57,8'd17} : s = 74;
	{8'd57,8'd18} : s = 75;
	{8'd57,8'd19} : s = 76;
	{8'd57,8'd20} : s = 77;
	{8'd57,8'd21} : s = 78;
	{8'd57,8'd22} : s = 79;
	{8'd57,8'd23} : s = 80;
	{8'd57,8'd24} : s = 81;
	{8'd57,8'd25} : s = 82;
	{8'd57,8'd26} : s = 83;
	{8'd57,8'd27} : s = 84;
	{8'd57,8'd28} : s = 85;
	{8'd57,8'd29} : s = 86;
	{8'd57,8'd30} : s = 87;
	{8'd57,8'd31} : s = 88;
	{8'd57,8'd32} : s = 89;
	{8'd57,8'd33} : s = 90;
	{8'd57,8'd34} : s = 91;
	{8'd57,8'd35} : s = 92;
	{8'd57,8'd36} : s = 93;
	{8'd57,8'd37} : s = 94;
	{8'd57,8'd38} : s = 95;
	{8'd57,8'd39} : s = 96;
	{8'd57,8'd40} : s = 97;
	{8'd57,8'd41} : s = 98;
	{8'd57,8'd42} : s = 99;
	{8'd57,8'd43} : s = 100;
	{8'd57,8'd44} : s = 101;
	{8'd57,8'd45} : s = 102;
	{8'd57,8'd46} : s = 103;
	{8'd57,8'd47} : s = 104;
	{8'd57,8'd48} : s = 105;
	{8'd57,8'd49} : s = 106;
	{8'd57,8'd50} : s = 107;
	{8'd57,8'd51} : s = 108;
	{8'd57,8'd52} : s = 109;
	{8'd57,8'd53} : s = 110;
	{8'd57,8'd54} : s = 111;
	{8'd57,8'd55} : s = 112;
	{8'd57,8'd56} : s = 113;
	{8'd57,8'd57} : s = 114;
	{8'd57,8'd58} : s = 115;
	{8'd57,8'd59} : s = 116;
	{8'd57,8'd60} : s = 117;
	{8'd57,8'd61} : s = 118;
	{8'd57,8'd62} : s = 119;
	{8'd57,8'd63} : s = 120;
	{8'd57,8'd64} : s = 121;
	{8'd57,8'd65} : s = 122;
	{8'd57,8'd66} : s = 123;
	{8'd57,8'd67} : s = 124;
	{8'd57,8'd68} : s = 125;
	{8'd57,8'd69} : s = 126;
	{8'd57,8'd70} : s = 127;
	{8'd57,8'd71} : s = 128;
	{8'd57,8'd72} : s = 129;
	{8'd57,8'd73} : s = 130;
	{8'd57,8'd74} : s = 131;
	{8'd57,8'd75} : s = 132;
	{8'd57,8'd76} : s = 133;
	{8'd57,8'd77} : s = 134;
	{8'd57,8'd78} : s = 135;
	{8'd57,8'd79} : s = 136;
	{8'd57,8'd80} : s = 137;
	{8'd57,8'd81} : s = 138;
	{8'd57,8'd82} : s = 139;
	{8'd57,8'd83} : s = 140;
	{8'd57,8'd84} : s = 141;
	{8'd57,8'd85} : s = 142;
	{8'd57,8'd86} : s = 143;
	{8'd57,8'd87} : s = 144;
	{8'd57,8'd88} : s = 145;
	{8'd57,8'd89} : s = 146;
	{8'd57,8'd90} : s = 147;
	{8'd57,8'd91} : s = 148;
	{8'd57,8'd92} : s = 149;
	{8'd57,8'd93} : s = 150;
	{8'd57,8'd94} : s = 151;
	{8'd57,8'd95} : s = 152;
	{8'd57,8'd96} : s = 153;
	{8'd57,8'd97} : s = 154;
	{8'd57,8'd98} : s = 155;
	{8'd57,8'd99} : s = 156;
	{8'd57,8'd100} : s = 157;
	{8'd57,8'd101} : s = 158;
	{8'd57,8'd102} : s = 159;
	{8'd57,8'd103} : s = 160;
	{8'd57,8'd104} : s = 161;
	{8'd57,8'd105} : s = 162;
	{8'd57,8'd106} : s = 163;
	{8'd57,8'd107} : s = 164;
	{8'd57,8'd108} : s = 165;
	{8'd57,8'd109} : s = 166;
	{8'd57,8'd110} : s = 167;
	{8'd57,8'd111} : s = 168;
	{8'd57,8'd112} : s = 169;
	{8'd57,8'd113} : s = 170;
	{8'd57,8'd114} : s = 171;
	{8'd57,8'd115} : s = 172;
	{8'd57,8'd116} : s = 173;
	{8'd57,8'd117} : s = 174;
	{8'd57,8'd118} : s = 175;
	{8'd57,8'd119} : s = 176;
	{8'd57,8'd120} : s = 177;
	{8'd57,8'd121} : s = 178;
	{8'd57,8'd122} : s = 179;
	{8'd57,8'd123} : s = 180;
	{8'd57,8'd124} : s = 181;
	{8'd57,8'd125} : s = 182;
	{8'd57,8'd126} : s = 183;
	{8'd57,8'd127} : s = 184;
	{8'd57,8'd128} : s = 185;
	{8'd57,8'd129} : s = 186;
	{8'd57,8'd130} : s = 187;
	{8'd57,8'd131} : s = 188;
	{8'd57,8'd132} : s = 189;
	{8'd57,8'd133} : s = 190;
	{8'd57,8'd134} : s = 191;
	{8'd57,8'd135} : s = 192;
	{8'd57,8'd136} : s = 193;
	{8'd57,8'd137} : s = 194;
	{8'd57,8'd138} : s = 195;
	{8'd57,8'd139} : s = 196;
	{8'd57,8'd140} : s = 197;
	{8'd57,8'd141} : s = 198;
	{8'd57,8'd142} : s = 199;
	{8'd57,8'd143} : s = 200;
	{8'd57,8'd144} : s = 201;
	{8'd57,8'd145} : s = 202;
	{8'd57,8'd146} : s = 203;
	{8'd57,8'd147} : s = 204;
	{8'd57,8'd148} : s = 205;
	{8'd57,8'd149} : s = 206;
	{8'd57,8'd150} : s = 207;
	{8'd57,8'd151} : s = 208;
	{8'd57,8'd152} : s = 209;
	{8'd57,8'd153} : s = 210;
	{8'd57,8'd154} : s = 211;
	{8'd57,8'd155} : s = 212;
	{8'd57,8'd156} : s = 213;
	{8'd57,8'd157} : s = 214;
	{8'd57,8'd158} : s = 215;
	{8'd57,8'd159} : s = 216;
	{8'd57,8'd160} : s = 217;
	{8'd57,8'd161} : s = 218;
	{8'd57,8'd162} : s = 219;
	{8'd57,8'd163} : s = 220;
	{8'd57,8'd164} : s = 221;
	{8'd57,8'd165} : s = 222;
	{8'd57,8'd166} : s = 223;
	{8'd57,8'd167} : s = 224;
	{8'd57,8'd168} : s = 225;
	{8'd57,8'd169} : s = 226;
	{8'd57,8'd170} : s = 227;
	{8'd57,8'd171} : s = 228;
	{8'd57,8'd172} : s = 229;
	{8'd57,8'd173} : s = 230;
	{8'd57,8'd174} : s = 231;
	{8'd57,8'd175} : s = 232;
	{8'd57,8'd176} : s = 233;
	{8'd57,8'd177} : s = 234;
	{8'd57,8'd178} : s = 235;
	{8'd57,8'd179} : s = 236;
	{8'd57,8'd180} : s = 237;
	{8'd57,8'd181} : s = 238;
	{8'd57,8'd182} : s = 239;
	{8'd57,8'd183} : s = 240;
	{8'd57,8'd184} : s = 241;
	{8'd57,8'd185} : s = 242;
	{8'd57,8'd186} : s = 243;
	{8'd57,8'd187} : s = 244;
	{8'd57,8'd188} : s = 245;
	{8'd57,8'd189} : s = 246;
	{8'd57,8'd190} : s = 247;
	{8'd57,8'd191} : s = 248;
	{8'd57,8'd192} : s = 249;
	{8'd57,8'd193} : s = 250;
	{8'd57,8'd194} : s = 251;
	{8'd57,8'd195} : s = 252;
	{8'd57,8'd196} : s = 253;
	{8'd57,8'd197} : s = 254;
	{8'd57,8'd198} : s = 255;
	{8'd57,8'd199} : s = 256;
	{8'd57,8'd200} : s = 257;
	{8'd57,8'd201} : s = 258;
	{8'd57,8'd202} : s = 259;
	{8'd57,8'd203} : s = 260;
	{8'd57,8'd204} : s = 261;
	{8'd57,8'd205} : s = 262;
	{8'd57,8'd206} : s = 263;
	{8'd57,8'd207} : s = 264;
	{8'd57,8'd208} : s = 265;
	{8'd57,8'd209} : s = 266;
	{8'd57,8'd210} : s = 267;
	{8'd57,8'd211} : s = 268;
	{8'd57,8'd212} : s = 269;
	{8'd57,8'd213} : s = 270;
	{8'd57,8'd214} : s = 271;
	{8'd57,8'd215} : s = 272;
	{8'd57,8'd216} : s = 273;
	{8'd57,8'd217} : s = 274;
	{8'd57,8'd218} : s = 275;
	{8'd57,8'd219} : s = 276;
	{8'd57,8'd220} : s = 277;
	{8'd57,8'd221} : s = 278;
	{8'd57,8'd222} : s = 279;
	{8'd57,8'd223} : s = 280;
	{8'd57,8'd224} : s = 281;
	{8'd57,8'd225} : s = 282;
	{8'd57,8'd226} : s = 283;
	{8'd57,8'd227} : s = 284;
	{8'd57,8'd228} : s = 285;
	{8'd57,8'd229} : s = 286;
	{8'd57,8'd230} : s = 287;
	{8'd57,8'd231} : s = 288;
	{8'd57,8'd232} : s = 289;
	{8'd57,8'd233} : s = 290;
	{8'd57,8'd234} : s = 291;
	{8'd57,8'd235} : s = 292;
	{8'd57,8'd236} : s = 293;
	{8'd57,8'd237} : s = 294;
	{8'd57,8'd238} : s = 295;
	{8'd57,8'd239} : s = 296;
	{8'd57,8'd240} : s = 297;
	{8'd57,8'd241} : s = 298;
	{8'd57,8'd242} : s = 299;
	{8'd57,8'd243} : s = 300;
	{8'd57,8'd244} : s = 301;
	{8'd57,8'd245} : s = 302;
	{8'd57,8'd246} : s = 303;
	{8'd57,8'd247} : s = 304;
	{8'd57,8'd248} : s = 305;
	{8'd57,8'd249} : s = 306;
	{8'd57,8'd250} : s = 307;
	{8'd57,8'd251} : s = 308;
	{8'd57,8'd252} : s = 309;
	{8'd57,8'd253} : s = 310;
	{8'd57,8'd254} : s = 311;
	{8'd57,8'd255} : s = 312;
	{8'd58,8'd0} : s = 58;
	{8'd58,8'd1} : s = 59;
	{8'd58,8'd2} : s = 60;
	{8'd58,8'd3} : s = 61;
	{8'd58,8'd4} : s = 62;
	{8'd58,8'd5} : s = 63;
	{8'd58,8'd6} : s = 64;
	{8'd58,8'd7} : s = 65;
	{8'd58,8'd8} : s = 66;
	{8'd58,8'd9} : s = 67;
	{8'd58,8'd10} : s = 68;
	{8'd58,8'd11} : s = 69;
	{8'd58,8'd12} : s = 70;
	{8'd58,8'd13} : s = 71;
	{8'd58,8'd14} : s = 72;
	{8'd58,8'd15} : s = 73;
	{8'd58,8'd16} : s = 74;
	{8'd58,8'd17} : s = 75;
	{8'd58,8'd18} : s = 76;
	{8'd58,8'd19} : s = 77;
	{8'd58,8'd20} : s = 78;
	{8'd58,8'd21} : s = 79;
	{8'd58,8'd22} : s = 80;
	{8'd58,8'd23} : s = 81;
	{8'd58,8'd24} : s = 82;
	{8'd58,8'd25} : s = 83;
	{8'd58,8'd26} : s = 84;
	{8'd58,8'd27} : s = 85;
	{8'd58,8'd28} : s = 86;
	{8'd58,8'd29} : s = 87;
	{8'd58,8'd30} : s = 88;
	{8'd58,8'd31} : s = 89;
	{8'd58,8'd32} : s = 90;
	{8'd58,8'd33} : s = 91;
	{8'd58,8'd34} : s = 92;
	{8'd58,8'd35} : s = 93;
	{8'd58,8'd36} : s = 94;
	{8'd58,8'd37} : s = 95;
	{8'd58,8'd38} : s = 96;
	{8'd58,8'd39} : s = 97;
	{8'd58,8'd40} : s = 98;
	{8'd58,8'd41} : s = 99;
	{8'd58,8'd42} : s = 100;
	{8'd58,8'd43} : s = 101;
	{8'd58,8'd44} : s = 102;
	{8'd58,8'd45} : s = 103;
	{8'd58,8'd46} : s = 104;
	{8'd58,8'd47} : s = 105;
	{8'd58,8'd48} : s = 106;
	{8'd58,8'd49} : s = 107;
	{8'd58,8'd50} : s = 108;
	{8'd58,8'd51} : s = 109;
	{8'd58,8'd52} : s = 110;
	{8'd58,8'd53} : s = 111;
	{8'd58,8'd54} : s = 112;
	{8'd58,8'd55} : s = 113;
	{8'd58,8'd56} : s = 114;
	{8'd58,8'd57} : s = 115;
	{8'd58,8'd58} : s = 116;
	{8'd58,8'd59} : s = 117;
	{8'd58,8'd60} : s = 118;
	{8'd58,8'd61} : s = 119;
	{8'd58,8'd62} : s = 120;
	{8'd58,8'd63} : s = 121;
	{8'd58,8'd64} : s = 122;
	{8'd58,8'd65} : s = 123;
	{8'd58,8'd66} : s = 124;
	{8'd58,8'd67} : s = 125;
	{8'd58,8'd68} : s = 126;
	{8'd58,8'd69} : s = 127;
	{8'd58,8'd70} : s = 128;
	{8'd58,8'd71} : s = 129;
	{8'd58,8'd72} : s = 130;
	{8'd58,8'd73} : s = 131;
	{8'd58,8'd74} : s = 132;
	{8'd58,8'd75} : s = 133;
	{8'd58,8'd76} : s = 134;
	{8'd58,8'd77} : s = 135;
	{8'd58,8'd78} : s = 136;
	{8'd58,8'd79} : s = 137;
	{8'd58,8'd80} : s = 138;
	{8'd58,8'd81} : s = 139;
	{8'd58,8'd82} : s = 140;
	{8'd58,8'd83} : s = 141;
	{8'd58,8'd84} : s = 142;
	{8'd58,8'd85} : s = 143;
	{8'd58,8'd86} : s = 144;
	{8'd58,8'd87} : s = 145;
	{8'd58,8'd88} : s = 146;
	{8'd58,8'd89} : s = 147;
	{8'd58,8'd90} : s = 148;
	{8'd58,8'd91} : s = 149;
	{8'd58,8'd92} : s = 150;
	{8'd58,8'd93} : s = 151;
	{8'd58,8'd94} : s = 152;
	{8'd58,8'd95} : s = 153;
	{8'd58,8'd96} : s = 154;
	{8'd58,8'd97} : s = 155;
	{8'd58,8'd98} : s = 156;
	{8'd58,8'd99} : s = 157;
	{8'd58,8'd100} : s = 158;
	{8'd58,8'd101} : s = 159;
	{8'd58,8'd102} : s = 160;
	{8'd58,8'd103} : s = 161;
	{8'd58,8'd104} : s = 162;
	{8'd58,8'd105} : s = 163;
	{8'd58,8'd106} : s = 164;
	{8'd58,8'd107} : s = 165;
	{8'd58,8'd108} : s = 166;
	{8'd58,8'd109} : s = 167;
	{8'd58,8'd110} : s = 168;
	{8'd58,8'd111} : s = 169;
	{8'd58,8'd112} : s = 170;
	{8'd58,8'd113} : s = 171;
	{8'd58,8'd114} : s = 172;
	{8'd58,8'd115} : s = 173;
	{8'd58,8'd116} : s = 174;
	{8'd58,8'd117} : s = 175;
	{8'd58,8'd118} : s = 176;
	{8'd58,8'd119} : s = 177;
	{8'd58,8'd120} : s = 178;
	{8'd58,8'd121} : s = 179;
	{8'd58,8'd122} : s = 180;
	{8'd58,8'd123} : s = 181;
	{8'd58,8'd124} : s = 182;
	{8'd58,8'd125} : s = 183;
	{8'd58,8'd126} : s = 184;
	{8'd58,8'd127} : s = 185;
	{8'd58,8'd128} : s = 186;
	{8'd58,8'd129} : s = 187;
	{8'd58,8'd130} : s = 188;
	{8'd58,8'd131} : s = 189;
	{8'd58,8'd132} : s = 190;
	{8'd58,8'd133} : s = 191;
	{8'd58,8'd134} : s = 192;
	{8'd58,8'd135} : s = 193;
	{8'd58,8'd136} : s = 194;
	{8'd58,8'd137} : s = 195;
	{8'd58,8'd138} : s = 196;
	{8'd58,8'd139} : s = 197;
	{8'd58,8'd140} : s = 198;
	{8'd58,8'd141} : s = 199;
	{8'd58,8'd142} : s = 200;
	{8'd58,8'd143} : s = 201;
	{8'd58,8'd144} : s = 202;
	{8'd58,8'd145} : s = 203;
	{8'd58,8'd146} : s = 204;
	{8'd58,8'd147} : s = 205;
	{8'd58,8'd148} : s = 206;
	{8'd58,8'd149} : s = 207;
	{8'd58,8'd150} : s = 208;
	{8'd58,8'd151} : s = 209;
	{8'd58,8'd152} : s = 210;
	{8'd58,8'd153} : s = 211;
	{8'd58,8'd154} : s = 212;
	{8'd58,8'd155} : s = 213;
	{8'd58,8'd156} : s = 214;
	{8'd58,8'd157} : s = 215;
	{8'd58,8'd158} : s = 216;
	{8'd58,8'd159} : s = 217;
	{8'd58,8'd160} : s = 218;
	{8'd58,8'd161} : s = 219;
	{8'd58,8'd162} : s = 220;
	{8'd58,8'd163} : s = 221;
	{8'd58,8'd164} : s = 222;
	{8'd58,8'd165} : s = 223;
	{8'd58,8'd166} : s = 224;
	{8'd58,8'd167} : s = 225;
	{8'd58,8'd168} : s = 226;
	{8'd58,8'd169} : s = 227;
	{8'd58,8'd170} : s = 228;
	{8'd58,8'd171} : s = 229;
	{8'd58,8'd172} : s = 230;
	{8'd58,8'd173} : s = 231;
	{8'd58,8'd174} : s = 232;
	{8'd58,8'd175} : s = 233;
	{8'd58,8'd176} : s = 234;
	{8'd58,8'd177} : s = 235;
	{8'd58,8'd178} : s = 236;
	{8'd58,8'd179} : s = 237;
	{8'd58,8'd180} : s = 238;
	{8'd58,8'd181} : s = 239;
	{8'd58,8'd182} : s = 240;
	{8'd58,8'd183} : s = 241;
	{8'd58,8'd184} : s = 242;
	{8'd58,8'd185} : s = 243;
	{8'd58,8'd186} : s = 244;
	{8'd58,8'd187} : s = 245;
	{8'd58,8'd188} : s = 246;
	{8'd58,8'd189} : s = 247;
	{8'd58,8'd190} : s = 248;
	{8'd58,8'd191} : s = 249;
	{8'd58,8'd192} : s = 250;
	{8'd58,8'd193} : s = 251;
	{8'd58,8'd194} : s = 252;
	{8'd58,8'd195} : s = 253;
	{8'd58,8'd196} : s = 254;
	{8'd58,8'd197} : s = 255;
	{8'd58,8'd198} : s = 256;
	{8'd58,8'd199} : s = 257;
	{8'd58,8'd200} : s = 258;
	{8'd58,8'd201} : s = 259;
	{8'd58,8'd202} : s = 260;
	{8'd58,8'd203} : s = 261;
	{8'd58,8'd204} : s = 262;
	{8'd58,8'd205} : s = 263;
	{8'd58,8'd206} : s = 264;
	{8'd58,8'd207} : s = 265;
	{8'd58,8'd208} : s = 266;
	{8'd58,8'd209} : s = 267;
	{8'd58,8'd210} : s = 268;
	{8'd58,8'd211} : s = 269;
	{8'd58,8'd212} : s = 270;
	{8'd58,8'd213} : s = 271;
	{8'd58,8'd214} : s = 272;
	{8'd58,8'd215} : s = 273;
	{8'd58,8'd216} : s = 274;
	{8'd58,8'd217} : s = 275;
	{8'd58,8'd218} : s = 276;
	{8'd58,8'd219} : s = 277;
	{8'd58,8'd220} : s = 278;
	{8'd58,8'd221} : s = 279;
	{8'd58,8'd222} : s = 280;
	{8'd58,8'd223} : s = 281;
	{8'd58,8'd224} : s = 282;
	{8'd58,8'd225} : s = 283;
	{8'd58,8'd226} : s = 284;
	{8'd58,8'd227} : s = 285;
	{8'd58,8'd228} : s = 286;
	{8'd58,8'd229} : s = 287;
	{8'd58,8'd230} : s = 288;
	{8'd58,8'd231} : s = 289;
	{8'd58,8'd232} : s = 290;
	{8'd58,8'd233} : s = 291;
	{8'd58,8'd234} : s = 292;
	{8'd58,8'd235} : s = 293;
	{8'd58,8'd236} : s = 294;
	{8'd58,8'd237} : s = 295;
	{8'd58,8'd238} : s = 296;
	{8'd58,8'd239} : s = 297;
	{8'd58,8'd240} : s = 298;
	{8'd58,8'd241} : s = 299;
	{8'd58,8'd242} : s = 300;
	{8'd58,8'd243} : s = 301;
	{8'd58,8'd244} : s = 302;
	{8'd58,8'd245} : s = 303;
	{8'd58,8'd246} : s = 304;
	{8'd58,8'd247} : s = 305;
	{8'd58,8'd248} : s = 306;
	{8'd58,8'd249} : s = 307;
	{8'd58,8'd250} : s = 308;
	{8'd58,8'd251} : s = 309;
	{8'd58,8'd252} : s = 310;
	{8'd58,8'd253} : s = 311;
	{8'd58,8'd254} : s = 312;
	{8'd58,8'd255} : s = 313;
	{8'd59,8'd0} : s = 59;
	{8'd59,8'd1} : s = 60;
	{8'd59,8'd2} : s = 61;
	{8'd59,8'd3} : s = 62;
	{8'd59,8'd4} : s = 63;
	{8'd59,8'd5} : s = 64;
	{8'd59,8'd6} : s = 65;
	{8'd59,8'd7} : s = 66;
	{8'd59,8'd8} : s = 67;
	{8'd59,8'd9} : s = 68;
	{8'd59,8'd10} : s = 69;
	{8'd59,8'd11} : s = 70;
	{8'd59,8'd12} : s = 71;
	{8'd59,8'd13} : s = 72;
	{8'd59,8'd14} : s = 73;
	{8'd59,8'd15} : s = 74;
	{8'd59,8'd16} : s = 75;
	{8'd59,8'd17} : s = 76;
	{8'd59,8'd18} : s = 77;
	{8'd59,8'd19} : s = 78;
	{8'd59,8'd20} : s = 79;
	{8'd59,8'd21} : s = 80;
	{8'd59,8'd22} : s = 81;
	{8'd59,8'd23} : s = 82;
	{8'd59,8'd24} : s = 83;
	{8'd59,8'd25} : s = 84;
	{8'd59,8'd26} : s = 85;
	{8'd59,8'd27} : s = 86;
	{8'd59,8'd28} : s = 87;
	{8'd59,8'd29} : s = 88;
	{8'd59,8'd30} : s = 89;
	{8'd59,8'd31} : s = 90;
	{8'd59,8'd32} : s = 91;
	{8'd59,8'd33} : s = 92;
	{8'd59,8'd34} : s = 93;
	{8'd59,8'd35} : s = 94;
	{8'd59,8'd36} : s = 95;
	{8'd59,8'd37} : s = 96;
	{8'd59,8'd38} : s = 97;
	{8'd59,8'd39} : s = 98;
	{8'd59,8'd40} : s = 99;
	{8'd59,8'd41} : s = 100;
	{8'd59,8'd42} : s = 101;
	{8'd59,8'd43} : s = 102;
	{8'd59,8'd44} : s = 103;
	{8'd59,8'd45} : s = 104;
	{8'd59,8'd46} : s = 105;
	{8'd59,8'd47} : s = 106;
	{8'd59,8'd48} : s = 107;
	{8'd59,8'd49} : s = 108;
	{8'd59,8'd50} : s = 109;
	{8'd59,8'd51} : s = 110;
	{8'd59,8'd52} : s = 111;
	{8'd59,8'd53} : s = 112;
	{8'd59,8'd54} : s = 113;
	{8'd59,8'd55} : s = 114;
	{8'd59,8'd56} : s = 115;
	{8'd59,8'd57} : s = 116;
	{8'd59,8'd58} : s = 117;
	{8'd59,8'd59} : s = 118;
	{8'd59,8'd60} : s = 119;
	{8'd59,8'd61} : s = 120;
	{8'd59,8'd62} : s = 121;
	{8'd59,8'd63} : s = 122;
	{8'd59,8'd64} : s = 123;
	{8'd59,8'd65} : s = 124;
	{8'd59,8'd66} : s = 125;
	{8'd59,8'd67} : s = 126;
	{8'd59,8'd68} : s = 127;
	{8'd59,8'd69} : s = 128;
	{8'd59,8'd70} : s = 129;
	{8'd59,8'd71} : s = 130;
	{8'd59,8'd72} : s = 131;
	{8'd59,8'd73} : s = 132;
	{8'd59,8'd74} : s = 133;
	{8'd59,8'd75} : s = 134;
	{8'd59,8'd76} : s = 135;
	{8'd59,8'd77} : s = 136;
	{8'd59,8'd78} : s = 137;
	{8'd59,8'd79} : s = 138;
	{8'd59,8'd80} : s = 139;
	{8'd59,8'd81} : s = 140;
	{8'd59,8'd82} : s = 141;
	{8'd59,8'd83} : s = 142;
	{8'd59,8'd84} : s = 143;
	{8'd59,8'd85} : s = 144;
	{8'd59,8'd86} : s = 145;
	{8'd59,8'd87} : s = 146;
	{8'd59,8'd88} : s = 147;
	{8'd59,8'd89} : s = 148;
	{8'd59,8'd90} : s = 149;
	{8'd59,8'd91} : s = 150;
	{8'd59,8'd92} : s = 151;
	{8'd59,8'd93} : s = 152;
	{8'd59,8'd94} : s = 153;
	{8'd59,8'd95} : s = 154;
	{8'd59,8'd96} : s = 155;
	{8'd59,8'd97} : s = 156;
	{8'd59,8'd98} : s = 157;
	{8'd59,8'd99} : s = 158;
	{8'd59,8'd100} : s = 159;
	{8'd59,8'd101} : s = 160;
	{8'd59,8'd102} : s = 161;
	{8'd59,8'd103} : s = 162;
	{8'd59,8'd104} : s = 163;
	{8'd59,8'd105} : s = 164;
	{8'd59,8'd106} : s = 165;
	{8'd59,8'd107} : s = 166;
	{8'd59,8'd108} : s = 167;
	{8'd59,8'd109} : s = 168;
	{8'd59,8'd110} : s = 169;
	{8'd59,8'd111} : s = 170;
	{8'd59,8'd112} : s = 171;
	{8'd59,8'd113} : s = 172;
	{8'd59,8'd114} : s = 173;
	{8'd59,8'd115} : s = 174;
	{8'd59,8'd116} : s = 175;
	{8'd59,8'd117} : s = 176;
	{8'd59,8'd118} : s = 177;
	{8'd59,8'd119} : s = 178;
	{8'd59,8'd120} : s = 179;
	{8'd59,8'd121} : s = 180;
	{8'd59,8'd122} : s = 181;
	{8'd59,8'd123} : s = 182;
	{8'd59,8'd124} : s = 183;
	{8'd59,8'd125} : s = 184;
	{8'd59,8'd126} : s = 185;
	{8'd59,8'd127} : s = 186;
	{8'd59,8'd128} : s = 187;
	{8'd59,8'd129} : s = 188;
	{8'd59,8'd130} : s = 189;
	{8'd59,8'd131} : s = 190;
	{8'd59,8'd132} : s = 191;
	{8'd59,8'd133} : s = 192;
	{8'd59,8'd134} : s = 193;
	{8'd59,8'd135} : s = 194;
	{8'd59,8'd136} : s = 195;
	{8'd59,8'd137} : s = 196;
	{8'd59,8'd138} : s = 197;
	{8'd59,8'd139} : s = 198;
	{8'd59,8'd140} : s = 199;
	{8'd59,8'd141} : s = 200;
	{8'd59,8'd142} : s = 201;
	{8'd59,8'd143} : s = 202;
	{8'd59,8'd144} : s = 203;
	{8'd59,8'd145} : s = 204;
	{8'd59,8'd146} : s = 205;
	{8'd59,8'd147} : s = 206;
	{8'd59,8'd148} : s = 207;
	{8'd59,8'd149} : s = 208;
	{8'd59,8'd150} : s = 209;
	{8'd59,8'd151} : s = 210;
	{8'd59,8'd152} : s = 211;
	{8'd59,8'd153} : s = 212;
	{8'd59,8'd154} : s = 213;
	{8'd59,8'd155} : s = 214;
	{8'd59,8'd156} : s = 215;
	{8'd59,8'd157} : s = 216;
	{8'd59,8'd158} : s = 217;
	{8'd59,8'd159} : s = 218;
	{8'd59,8'd160} : s = 219;
	{8'd59,8'd161} : s = 220;
	{8'd59,8'd162} : s = 221;
	{8'd59,8'd163} : s = 222;
	{8'd59,8'd164} : s = 223;
	{8'd59,8'd165} : s = 224;
	{8'd59,8'd166} : s = 225;
	{8'd59,8'd167} : s = 226;
	{8'd59,8'd168} : s = 227;
	{8'd59,8'd169} : s = 228;
	{8'd59,8'd170} : s = 229;
	{8'd59,8'd171} : s = 230;
	{8'd59,8'd172} : s = 231;
	{8'd59,8'd173} : s = 232;
	{8'd59,8'd174} : s = 233;
	{8'd59,8'd175} : s = 234;
	{8'd59,8'd176} : s = 235;
	{8'd59,8'd177} : s = 236;
	{8'd59,8'd178} : s = 237;
	{8'd59,8'd179} : s = 238;
	{8'd59,8'd180} : s = 239;
	{8'd59,8'd181} : s = 240;
	{8'd59,8'd182} : s = 241;
	{8'd59,8'd183} : s = 242;
	{8'd59,8'd184} : s = 243;
	{8'd59,8'd185} : s = 244;
	{8'd59,8'd186} : s = 245;
	{8'd59,8'd187} : s = 246;
	{8'd59,8'd188} : s = 247;
	{8'd59,8'd189} : s = 248;
	{8'd59,8'd190} : s = 249;
	{8'd59,8'd191} : s = 250;
	{8'd59,8'd192} : s = 251;
	{8'd59,8'd193} : s = 252;
	{8'd59,8'd194} : s = 253;
	{8'd59,8'd195} : s = 254;
	{8'd59,8'd196} : s = 255;
	{8'd59,8'd197} : s = 256;
	{8'd59,8'd198} : s = 257;
	{8'd59,8'd199} : s = 258;
	{8'd59,8'd200} : s = 259;
	{8'd59,8'd201} : s = 260;
	{8'd59,8'd202} : s = 261;
	{8'd59,8'd203} : s = 262;
	{8'd59,8'd204} : s = 263;
	{8'd59,8'd205} : s = 264;
	{8'd59,8'd206} : s = 265;
	{8'd59,8'd207} : s = 266;
	{8'd59,8'd208} : s = 267;
	{8'd59,8'd209} : s = 268;
	{8'd59,8'd210} : s = 269;
	{8'd59,8'd211} : s = 270;
	{8'd59,8'd212} : s = 271;
	{8'd59,8'd213} : s = 272;
	{8'd59,8'd214} : s = 273;
	{8'd59,8'd215} : s = 274;
	{8'd59,8'd216} : s = 275;
	{8'd59,8'd217} : s = 276;
	{8'd59,8'd218} : s = 277;
	{8'd59,8'd219} : s = 278;
	{8'd59,8'd220} : s = 279;
	{8'd59,8'd221} : s = 280;
	{8'd59,8'd222} : s = 281;
	{8'd59,8'd223} : s = 282;
	{8'd59,8'd224} : s = 283;
	{8'd59,8'd225} : s = 284;
	{8'd59,8'd226} : s = 285;
	{8'd59,8'd227} : s = 286;
	{8'd59,8'd228} : s = 287;
	{8'd59,8'd229} : s = 288;
	{8'd59,8'd230} : s = 289;
	{8'd59,8'd231} : s = 290;
	{8'd59,8'd232} : s = 291;
	{8'd59,8'd233} : s = 292;
	{8'd59,8'd234} : s = 293;
	{8'd59,8'd235} : s = 294;
	{8'd59,8'd236} : s = 295;
	{8'd59,8'd237} : s = 296;
	{8'd59,8'd238} : s = 297;
	{8'd59,8'd239} : s = 298;
	{8'd59,8'd240} : s = 299;
	{8'd59,8'd241} : s = 300;
	{8'd59,8'd242} : s = 301;
	{8'd59,8'd243} : s = 302;
	{8'd59,8'd244} : s = 303;
	{8'd59,8'd245} : s = 304;
	{8'd59,8'd246} : s = 305;
	{8'd59,8'd247} : s = 306;
	{8'd59,8'd248} : s = 307;
	{8'd59,8'd249} : s = 308;
	{8'd59,8'd250} : s = 309;
	{8'd59,8'd251} : s = 310;
	{8'd59,8'd252} : s = 311;
	{8'd59,8'd253} : s = 312;
	{8'd59,8'd254} : s = 313;
	{8'd59,8'd255} : s = 314;
	{8'd60,8'd0} : s = 60;
	{8'd60,8'd1} : s = 61;
	{8'd60,8'd2} : s = 62;
	{8'd60,8'd3} : s = 63;
	{8'd60,8'd4} : s = 64;
	{8'd60,8'd5} : s = 65;
	{8'd60,8'd6} : s = 66;
	{8'd60,8'd7} : s = 67;
	{8'd60,8'd8} : s = 68;
	{8'd60,8'd9} : s = 69;
	{8'd60,8'd10} : s = 70;
	{8'd60,8'd11} : s = 71;
	{8'd60,8'd12} : s = 72;
	{8'd60,8'd13} : s = 73;
	{8'd60,8'd14} : s = 74;
	{8'd60,8'd15} : s = 75;
	{8'd60,8'd16} : s = 76;
	{8'd60,8'd17} : s = 77;
	{8'd60,8'd18} : s = 78;
	{8'd60,8'd19} : s = 79;
	{8'd60,8'd20} : s = 80;
	{8'd60,8'd21} : s = 81;
	{8'd60,8'd22} : s = 82;
	{8'd60,8'd23} : s = 83;
	{8'd60,8'd24} : s = 84;
	{8'd60,8'd25} : s = 85;
	{8'd60,8'd26} : s = 86;
	{8'd60,8'd27} : s = 87;
	{8'd60,8'd28} : s = 88;
	{8'd60,8'd29} : s = 89;
	{8'd60,8'd30} : s = 90;
	{8'd60,8'd31} : s = 91;
	{8'd60,8'd32} : s = 92;
	{8'd60,8'd33} : s = 93;
	{8'd60,8'd34} : s = 94;
	{8'd60,8'd35} : s = 95;
	{8'd60,8'd36} : s = 96;
	{8'd60,8'd37} : s = 97;
	{8'd60,8'd38} : s = 98;
	{8'd60,8'd39} : s = 99;
	{8'd60,8'd40} : s = 100;
	{8'd60,8'd41} : s = 101;
	{8'd60,8'd42} : s = 102;
	{8'd60,8'd43} : s = 103;
	{8'd60,8'd44} : s = 104;
	{8'd60,8'd45} : s = 105;
	{8'd60,8'd46} : s = 106;
	{8'd60,8'd47} : s = 107;
	{8'd60,8'd48} : s = 108;
	{8'd60,8'd49} : s = 109;
	{8'd60,8'd50} : s = 110;
	{8'd60,8'd51} : s = 111;
	{8'd60,8'd52} : s = 112;
	{8'd60,8'd53} : s = 113;
	{8'd60,8'd54} : s = 114;
	{8'd60,8'd55} : s = 115;
	{8'd60,8'd56} : s = 116;
	{8'd60,8'd57} : s = 117;
	{8'd60,8'd58} : s = 118;
	{8'd60,8'd59} : s = 119;
	{8'd60,8'd60} : s = 120;
	{8'd60,8'd61} : s = 121;
	{8'd60,8'd62} : s = 122;
	{8'd60,8'd63} : s = 123;
	{8'd60,8'd64} : s = 124;
	{8'd60,8'd65} : s = 125;
	{8'd60,8'd66} : s = 126;
	{8'd60,8'd67} : s = 127;
	{8'd60,8'd68} : s = 128;
	{8'd60,8'd69} : s = 129;
	{8'd60,8'd70} : s = 130;
	{8'd60,8'd71} : s = 131;
	{8'd60,8'd72} : s = 132;
	{8'd60,8'd73} : s = 133;
	{8'd60,8'd74} : s = 134;
	{8'd60,8'd75} : s = 135;
	{8'd60,8'd76} : s = 136;
	{8'd60,8'd77} : s = 137;
	{8'd60,8'd78} : s = 138;
	{8'd60,8'd79} : s = 139;
	{8'd60,8'd80} : s = 140;
	{8'd60,8'd81} : s = 141;
	{8'd60,8'd82} : s = 142;
	{8'd60,8'd83} : s = 143;
	{8'd60,8'd84} : s = 144;
	{8'd60,8'd85} : s = 145;
	{8'd60,8'd86} : s = 146;
	{8'd60,8'd87} : s = 147;
	{8'd60,8'd88} : s = 148;
	{8'd60,8'd89} : s = 149;
	{8'd60,8'd90} : s = 150;
	{8'd60,8'd91} : s = 151;
	{8'd60,8'd92} : s = 152;
	{8'd60,8'd93} : s = 153;
	{8'd60,8'd94} : s = 154;
	{8'd60,8'd95} : s = 155;
	{8'd60,8'd96} : s = 156;
	{8'd60,8'd97} : s = 157;
	{8'd60,8'd98} : s = 158;
	{8'd60,8'd99} : s = 159;
	{8'd60,8'd100} : s = 160;
	{8'd60,8'd101} : s = 161;
	{8'd60,8'd102} : s = 162;
	{8'd60,8'd103} : s = 163;
	{8'd60,8'd104} : s = 164;
	{8'd60,8'd105} : s = 165;
	{8'd60,8'd106} : s = 166;
	{8'd60,8'd107} : s = 167;
	{8'd60,8'd108} : s = 168;
	{8'd60,8'd109} : s = 169;
	{8'd60,8'd110} : s = 170;
	{8'd60,8'd111} : s = 171;
	{8'd60,8'd112} : s = 172;
	{8'd60,8'd113} : s = 173;
	{8'd60,8'd114} : s = 174;
	{8'd60,8'd115} : s = 175;
	{8'd60,8'd116} : s = 176;
	{8'd60,8'd117} : s = 177;
	{8'd60,8'd118} : s = 178;
	{8'd60,8'd119} : s = 179;
	{8'd60,8'd120} : s = 180;
	{8'd60,8'd121} : s = 181;
	{8'd60,8'd122} : s = 182;
	{8'd60,8'd123} : s = 183;
	{8'd60,8'd124} : s = 184;
	{8'd60,8'd125} : s = 185;
	{8'd60,8'd126} : s = 186;
	{8'd60,8'd127} : s = 187;
	{8'd60,8'd128} : s = 188;
	{8'd60,8'd129} : s = 189;
	{8'd60,8'd130} : s = 190;
	{8'd60,8'd131} : s = 191;
	{8'd60,8'd132} : s = 192;
	{8'd60,8'd133} : s = 193;
	{8'd60,8'd134} : s = 194;
	{8'd60,8'd135} : s = 195;
	{8'd60,8'd136} : s = 196;
	{8'd60,8'd137} : s = 197;
	{8'd60,8'd138} : s = 198;
	{8'd60,8'd139} : s = 199;
	{8'd60,8'd140} : s = 200;
	{8'd60,8'd141} : s = 201;
	{8'd60,8'd142} : s = 202;
	{8'd60,8'd143} : s = 203;
	{8'd60,8'd144} : s = 204;
	{8'd60,8'd145} : s = 205;
	{8'd60,8'd146} : s = 206;
	{8'd60,8'd147} : s = 207;
	{8'd60,8'd148} : s = 208;
	{8'd60,8'd149} : s = 209;
	{8'd60,8'd150} : s = 210;
	{8'd60,8'd151} : s = 211;
	{8'd60,8'd152} : s = 212;
	{8'd60,8'd153} : s = 213;
	{8'd60,8'd154} : s = 214;
	{8'd60,8'd155} : s = 215;
	{8'd60,8'd156} : s = 216;
	{8'd60,8'd157} : s = 217;
	{8'd60,8'd158} : s = 218;
	{8'd60,8'd159} : s = 219;
	{8'd60,8'd160} : s = 220;
	{8'd60,8'd161} : s = 221;
	{8'd60,8'd162} : s = 222;
	{8'd60,8'd163} : s = 223;
	{8'd60,8'd164} : s = 224;
	{8'd60,8'd165} : s = 225;
	{8'd60,8'd166} : s = 226;
	{8'd60,8'd167} : s = 227;
	{8'd60,8'd168} : s = 228;
	{8'd60,8'd169} : s = 229;
	{8'd60,8'd170} : s = 230;
	{8'd60,8'd171} : s = 231;
	{8'd60,8'd172} : s = 232;
	{8'd60,8'd173} : s = 233;
	{8'd60,8'd174} : s = 234;
	{8'd60,8'd175} : s = 235;
	{8'd60,8'd176} : s = 236;
	{8'd60,8'd177} : s = 237;
	{8'd60,8'd178} : s = 238;
	{8'd60,8'd179} : s = 239;
	{8'd60,8'd180} : s = 240;
	{8'd60,8'd181} : s = 241;
	{8'd60,8'd182} : s = 242;
	{8'd60,8'd183} : s = 243;
	{8'd60,8'd184} : s = 244;
	{8'd60,8'd185} : s = 245;
	{8'd60,8'd186} : s = 246;
	{8'd60,8'd187} : s = 247;
	{8'd60,8'd188} : s = 248;
	{8'd60,8'd189} : s = 249;
	{8'd60,8'd190} : s = 250;
	{8'd60,8'd191} : s = 251;
	{8'd60,8'd192} : s = 252;
	{8'd60,8'd193} : s = 253;
	{8'd60,8'd194} : s = 254;
	{8'd60,8'd195} : s = 255;
	{8'd60,8'd196} : s = 256;
	{8'd60,8'd197} : s = 257;
	{8'd60,8'd198} : s = 258;
	{8'd60,8'd199} : s = 259;
	{8'd60,8'd200} : s = 260;
	{8'd60,8'd201} : s = 261;
	{8'd60,8'd202} : s = 262;
	{8'd60,8'd203} : s = 263;
	{8'd60,8'd204} : s = 264;
	{8'd60,8'd205} : s = 265;
	{8'd60,8'd206} : s = 266;
	{8'd60,8'd207} : s = 267;
	{8'd60,8'd208} : s = 268;
	{8'd60,8'd209} : s = 269;
	{8'd60,8'd210} : s = 270;
	{8'd60,8'd211} : s = 271;
	{8'd60,8'd212} : s = 272;
	{8'd60,8'd213} : s = 273;
	{8'd60,8'd214} : s = 274;
	{8'd60,8'd215} : s = 275;
	{8'd60,8'd216} : s = 276;
	{8'd60,8'd217} : s = 277;
	{8'd60,8'd218} : s = 278;
	{8'd60,8'd219} : s = 279;
	{8'd60,8'd220} : s = 280;
	{8'd60,8'd221} : s = 281;
	{8'd60,8'd222} : s = 282;
	{8'd60,8'd223} : s = 283;
	{8'd60,8'd224} : s = 284;
	{8'd60,8'd225} : s = 285;
	{8'd60,8'd226} : s = 286;
	{8'd60,8'd227} : s = 287;
	{8'd60,8'd228} : s = 288;
	{8'd60,8'd229} : s = 289;
	{8'd60,8'd230} : s = 290;
	{8'd60,8'd231} : s = 291;
	{8'd60,8'd232} : s = 292;
	{8'd60,8'd233} : s = 293;
	{8'd60,8'd234} : s = 294;
	{8'd60,8'd235} : s = 295;
	{8'd60,8'd236} : s = 296;
	{8'd60,8'd237} : s = 297;
	{8'd60,8'd238} : s = 298;
	{8'd60,8'd239} : s = 299;
	{8'd60,8'd240} : s = 300;
	{8'd60,8'd241} : s = 301;
	{8'd60,8'd242} : s = 302;
	{8'd60,8'd243} : s = 303;
	{8'd60,8'd244} : s = 304;
	{8'd60,8'd245} : s = 305;
	{8'd60,8'd246} : s = 306;
	{8'd60,8'd247} : s = 307;
	{8'd60,8'd248} : s = 308;
	{8'd60,8'd249} : s = 309;
	{8'd60,8'd250} : s = 310;
	{8'd60,8'd251} : s = 311;
	{8'd60,8'd252} : s = 312;
	{8'd60,8'd253} : s = 313;
	{8'd60,8'd254} : s = 314;
	{8'd60,8'd255} : s = 315;
	{8'd61,8'd0} : s = 61;
	{8'd61,8'd1} : s = 62;
	{8'd61,8'd2} : s = 63;
	{8'd61,8'd3} : s = 64;
	{8'd61,8'd4} : s = 65;
	{8'd61,8'd5} : s = 66;
	{8'd61,8'd6} : s = 67;
	{8'd61,8'd7} : s = 68;
	{8'd61,8'd8} : s = 69;
	{8'd61,8'd9} : s = 70;
	{8'd61,8'd10} : s = 71;
	{8'd61,8'd11} : s = 72;
	{8'd61,8'd12} : s = 73;
	{8'd61,8'd13} : s = 74;
	{8'd61,8'd14} : s = 75;
	{8'd61,8'd15} : s = 76;
	{8'd61,8'd16} : s = 77;
	{8'd61,8'd17} : s = 78;
	{8'd61,8'd18} : s = 79;
	{8'd61,8'd19} : s = 80;
	{8'd61,8'd20} : s = 81;
	{8'd61,8'd21} : s = 82;
	{8'd61,8'd22} : s = 83;
	{8'd61,8'd23} : s = 84;
	{8'd61,8'd24} : s = 85;
	{8'd61,8'd25} : s = 86;
	{8'd61,8'd26} : s = 87;
	{8'd61,8'd27} : s = 88;
	{8'd61,8'd28} : s = 89;
	{8'd61,8'd29} : s = 90;
	{8'd61,8'd30} : s = 91;
	{8'd61,8'd31} : s = 92;
	{8'd61,8'd32} : s = 93;
	{8'd61,8'd33} : s = 94;
	{8'd61,8'd34} : s = 95;
	{8'd61,8'd35} : s = 96;
	{8'd61,8'd36} : s = 97;
	{8'd61,8'd37} : s = 98;
	{8'd61,8'd38} : s = 99;
	{8'd61,8'd39} : s = 100;
	{8'd61,8'd40} : s = 101;
	{8'd61,8'd41} : s = 102;
	{8'd61,8'd42} : s = 103;
	{8'd61,8'd43} : s = 104;
	{8'd61,8'd44} : s = 105;
	{8'd61,8'd45} : s = 106;
	{8'd61,8'd46} : s = 107;
	{8'd61,8'd47} : s = 108;
	{8'd61,8'd48} : s = 109;
	{8'd61,8'd49} : s = 110;
	{8'd61,8'd50} : s = 111;
	{8'd61,8'd51} : s = 112;
	{8'd61,8'd52} : s = 113;
	{8'd61,8'd53} : s = 114;
	{8'd61,8'd54} : s = 115;
	{8'd61,8'd55} : s = 116;
	{8'd61,8'd56} : s = 117;
	{8'd61,8'd57} : s = 118;
	{8'd61,8'd58} : s = 119;
	{8'd61,8'd59} : s = 120;
	{8'd61,8'd60} : s = 121;
	{8'd61,8'd61} : s = 122;
	{8'd61,8'd62} : s = 123;
	{8'd61,8'd63} : s = 124;
	{8'd61,8'd64} : s = 125;
	{8'd61,8'd65} : s = 126;
	{8'd61,8'd66} : s = 127;
	{8'd61,8'd67} : s = 128;
	{8'd61,8'd68} : s = 129;
	{8'd61,8'd69} : s = 130;
	{8'd61,8'd70} : s = 131;
	{8'd61,8'd71} : s = 132;
	{8'd61,8'd72} : s = 133;
	{8'd61,8'd73} : s = 134;
	{8'd61,8'd74} : s = 135;
	{8'd61,8'd75} : s = 136;
	{8'd61,8'd76} : s = 137;
	{8'd61,8'd77} : s = 138;
	{8'd61,8'd78} : s = 139;
	{8'd61,8'd79} : s = 140;
	{8'd61,8'd80} : s = 141;
	{8'd61,8'd81} : s = 142;
	{8'd61,8'd82} : s = 143;
	{8'd61,8'd83} : s = 144;
	{8'd61,8'd84} : s = 145;
	{8'd61,8'd85} : s = 146;
	{8'd61,8'd86} : s = 147;
	{8'd61,8'd87} : s = 148;
	{8'd61,8'd88} : s = 149;
	{8'd61,8'd89} : s = 150;
	{8'd61,8'd90} : s = 151;
	{8'd61,8'd91} : s = 152;
	{8'd61,8'd92} : s = 153;
	{8'd61,8'd93} : s = 154;
	{8'd61,8'd94} : s = 155;
	{8'd61,8'd95} : s = 156;
	{8'd61,8'd96} : s = 157;
	{8'd61,8'd97} : s = 158;
	{8'd61,8'd98} : s = 159;
	{8'd61,8'd99} : s = 160;
	{8'd61,8'd100} : s = 161;
	{8'd61,8'd101} : s = 162;
	{8'd61,8'd102} : s = 163;
	{8'd61,8'd103} : s = 164;
	{8'd61,8'd104} : s = 165;
	{8'd61,8'd105} : s = 166;
	{8'd61,8'd106} : s = 167;
	{8'd61,8'd107} : s = 168;
	{8'd61,8'd108} : s = 169;
	{8'd61,8'd109} : s = 170;
	{8'd61,8'd110} : s = 171;
	{8'd61,8'd111} : s = 172;
	{8'd61,8'd112} : s = 173;
	{8'd61,8'd113} : s = 174;
	{8'd61,8'd114} : s = 175;
	{8'd61,8'd115} : s = 176;
	{8'd61,8'd116} : s = 177;
	{8'd61,8'd117} : s = 178;
	{8'd61,8'd118} : s = 179;
	{8'd61,8'd119} : s = 180;
	{8'd61,8'd120} : s = 181;
	{8'd61,8'd121} : s = 182;
	{8'd61,8'd122} : s = 183;
	{8'd61,8'd123} : s = 184;
	{8'd61,8'd124} : s = 185;
	{8'd61,8'd125} : s = 186;
	{8'd61,8'd126} : s = 187;
	{8'd61,8'd127} : s = 188;
	{8'd61,8'd128} : s = 189;
	{8'd61,8'd129} : s = 190;
	{8'd61,8'd130} : s = 191;
	{8'd61,8'd131} : s = 192;
	{8'd61,8'd132} : s = 193;
	{8'd61,8'd133} : s = 194;
	{8'd61,8'd134} : s = 195;
	{8'd61,8'd135} : s = 196;
	{8'd61,8'd136} : s = 197;
	{8'd61,8'd137} : s = 198;
	{8'd61,8'd138} : s = 199;
	{8'd61,8'd139} : s = 200;
	{8'd61,8'd140} : s = 201;
	{8'd61,8'd141} : s = 202;
	{8'd61,8'd142} : s = 203;
	{8'd61,8'd143} : s = 204;
	{8'd61,8'd144} : s = 205;
	{8'd61,8'd145} : s = 206;
	{8'd61,8'd146} : s = 207;
	{8'd61,8'd147} : s = 208;
	{8'd61,8'd148} : s = 209;
	{8'd61,8'd149} : s = 210;
	{8'd61,8'd150} : s = 211;
	{8'd61,8'd151} : s = 212;
	{8'd61,8'd152} : s = 213;
	{8'd61,8'd153} : s = 214;
	{8'd61,8'd154} : s = 215;
	{8'd61,8'd155} : s = 216;
	{8'd61,8'd156} : s = 217;
	{8'd61,8'd157} : s = 218;
	{8'd61,8'd158} : s = 219;
	{8'd61,8'd159} : s = 220;
	{8'd61,8'd160} : s = 221;
	{8'd61,8'd161} : s = 222;
	{8'd61,8'd162} : s = 223;
	{8'd61,8'd163} : s = 224;
	{8'd61,8'd164} : s = 225;
	{8'd61,8'd165} : s = 226;
	{8'd61,8'd166} : s = 227;
	{8'd61,8'd167} : s = 228;
	{8'd61,8'd168} : s = 229;
	{8'd61,8'd169} : s = 230;
	{8'd61,8'd170} : s = 231;
	{8'd61,8'd171} : s = 232;
	{8'd61,8'd172} : s = 233;
	{8'd61,8'd173} : s = 234;
	{8'd61,8'd174} : s = 235;
	{8'd61,8'd175} : s = 236;
	{8'd61,8'd176} : s = 237;
	{8'd61,8'd177} : s = 238;
	{8'd61,8'd178} : s = 239;
	{8'd61,8'd179} : s = 240;
	{8'd61,8'd180} : s = 241;
	{8'd61,8'd181} : s = 242;
	{8'd61,8'd182} : s = 243;
	{8'd61,8'd183} : s = 244;
	{8'd61,8'd184} : s = 245;
	{8'd61,8'd185} : s = 246;
	{8'd61,8'd186} : s = 247;
	{8'd61,8'd187} : s = 248;
	{8'd61,8'd188} : s = 249;
	{8'd61,8'd189} : s = 250;
	{8'd61,8'd190} : s = 251;
	{8'd61,8'd191} : s = 252;
	{8'd61,8'd192} : s = 253;
	{8'd61,8'd193} : s = 254;
	{8'd61,8'd194} : s = 255;
	{8'd61,8'd195} : s = 256;
	{8'd61,8'd196} : s = 257;
	{8'd61,8'd197} : s = 258;
	{8'd61,8'd198} : s = 259;
	{8'd61,8'd199} : s = 260;
	{8'd61,8'd200} : s = 261;
	{8'd61,8'd201} : s = 262;
	{8'd61,8'd202} : s = 263;
	{8'd61,8'd203} : s = 264;
	{8'd61,8'd204} : s = 265;
	{8'd61,8'd205} : s = 266;
	{8'd61,8'd206} : s = 267;
	{8'd61,8'd207} : s = 268;
	{8'd61,8'd208} : s = 269;
	{8'd61,8'd209} : s = 270;
	{8'd61,8'd210} : s = 271;
	{8'd61,8'd211} : s = 272;
	{8'd61,8'd212} : s = 273;
	{8'd61,8'd213} : s = 274;
	{8'd61,8'd214} : s = 275;
	{8'd61,8'd215} : s = 276;
	{8'd61,8'd216} : s = 277;
	{8'd61,8'd217} : s = 278;
	{8'd61,8'd218} : s = 279;
	{8'd61,8'd219} : s = 280;
	{8'd61,8'd220} : s = 281;
	{8'd61,8'd221} : s = 282;
	{8'd61,8'd222} : s = 283;
	{8'd61,8'd223} : s = 284;
	{8'd61,8'd224} : s = 285;
	{8'd61,8'd225} : s = 286;
	{8'd61,8'd226} : s = 287;
	{8'd61,8'd227} : s = 288;
	{8'd61,8'd228} : s = 289;
	{8'd61,8'd229} : s = 290;
	{8'd61,8'd230} : s = 291;
	{8'd61,8'd231} : s = 292;
	{8'd61,8'd232} : s = 293;
	{8'd61,8'd233} : s = 294;
	{8'd61,8'd234} : s = 295;
	{8'd61,8'd235} : s = 296;
	{8'd61,8'd236} : s = 297;
	{8'd61,8'd237} : s = 298;
	{8'd61,8'd238} : s = 299;
	{8'd61,8'd239} : s = 300;
	{8'd61,8'd240} : s = 301;
	{8'd61,8'd241} : s = 302;
	{8'd61,8'd242} : s = 303;
	{8'd61,8'd243} : s = 304;
	{8'd61,8'd244} : s = 305;
	{8'd61,8'd245} : s = 306;
	{8'd61,8'd246} : s = 307;
	{8'd61,8'd247} : s = 308;
	{8'd61,8'd248} : s = 309;
	{8'd61,8'd249} : s = 310;
	{8'd61,8'd250} : s = 311;
	{8'd61,8'd251} : s = 312;
	{8'd61,8'd252} : s = 313;
	{8'd61,8'd253} : s = 314;
	{8'd61,8'd254} : s = 315;
	{8'd61,8'd255} : s = 316;
	{8'd62,8'd0} : s = 62;
	{8'd62,8'd1} : s = 63;
	{8'd62,8'd2} : s = 64;
	{8'd62,8'd3} : s = 65;
	{8'd62,8'd4} : s = 66;
	{8'd62,8'd5} : s = 67;
	{8'd62,8'd6} : s = 68;
	{8'd62,8'd7} : s = 69;
	{8'd62,8'd8} : s = 70;
	{8'd62,8'd9} : s = 71;
	{8'd62,8'd10} : s = 72;
	{8'd62,8'd11} : s = 73;
	{8'd62,8'd12} : s = 74;
	{8'd62,8'd13} : s = 75;
	{8'd62,8'd14} : s = 76;
	{8'd62,8'd15} : s = 77;
	{8'd62,8'd16} : s = 78;
	{8'd62,8'd17} : s = 79;
	{8'd62,8'd18} : s = 80;
	{8'd62,8'd19} : s = 81;
	{8'd62,8'd20} : s = 82;
	{8'd62,8'd21} : s = 83;
	{8'd62,8'd22} : s = 84;
	{8'd62,8'd23} : s = 85;
	{8'd62,8'd24} : s = 86;
	{8'd62,8'd25} : s = 87;
	{8'd62,8'd26} : s = 88;
	{8'd62,8'd27} : s = 89;
	{8'd62,8'd28} : s = 90;
	{8'd62,8'd29} : s = 91;
	{8'd62,8'd30} : s = 92;
	{8'd62,8'd31} : s = 93;
	{8'd62,8'd32} : s = 94;
	{8'd62,8'd33} : s = 95;
	{8'd62,8'd34} : s = 96;
	{8'd62,8'd35} : s = 97;
	{8'd62,8'd36} : s = 98;
	{8'd62,8'd37} : s = 99;
	{8'd62,8'd38} : s = 100;
	{8'd62,8'd39} : s = 101;
	{8'd62,8'd40} : s = 102;
	{8'd62,8'd41} : s = 103;
	{8'd62,8'd42} : s = 104;
	{8'd62,8'd43} : s = 105;
	{8'd62,8'd44} : s = 106;
	{8'd62,8'd45} : s = 107;
	{8'd62,8'd46} : s = 108;
	{8'd62,8'd47} : s = 109;
	{8'd62,8'd48} : s = 110;
	{8'd62,8'd49} : s = 111;
	{8'd62,8'd50} : s = 112;
	{8'd62,8'd51} : s = 113;
	{8'd62,8'd52} : s = 114;
	{8'd62,8'd53} : s = 115;
	{8'd62,8'd54} : s = 116;
	{8'd62,8'd55} : s = 117;
	{8'd62,8'd56} : s = 118;
	{8'd62,8'd57} : s = 119;
	{8'd62,8'd58} : s = 120;
	{8'd62,8'd59} : s = 121;
	{8'd62,8'd60} : s = 122;
	{8'd62,8'd61} : s = 123;
	{8'd62,8'd62} : s = 124;
	{8'd62,8'd63} : s = 125;
	{8'd62,8'd64} : s = 126;
	{8'd62,8'd65} : s = 127;
	{8'd62,8'd66} : s = 128;
	{8'd62,8'd67} : s = 129;
	{8'd62,8'd68} : s = 130;
	{8'd62,8'd69} : s = 131;
	{8'd62,8'd70} : s = 132;
	{8'd62,8'd71} : s = 133;
	{8'd62,8'd72} : s = 134;
	{8'd62,8'd73} : s = 135;
	{8'd62,8'd74} : s = 136;
	{8'd62,8'd75} : s = 137;
	{8'd62,8'd76} : s = 138;
	{8'd62,8'd77} : s = 139;
	{8'd62,8'd78} : s = 140;
	{8'd62,8'd79} : s = 141;
	{8'd62,8'd80} : s = 142;
	{8'd62,8'd81} : s = 143;
	{8'd62,8'd82} : s = 144;
	{8'd62,8'd83} : s = 145;
	{8'd62,8'd84} : s = 146;
	{8'd62,8'd85} : s = 147;
	{8'd62,8'd86} : s = 148;
	{8'd62,8'd87} : s = 149;
	{8'd62,8'd88} : s = 150;
	{8'd62,8'd89} : s = 151;
	{8'd62,8'd90} : s = 152;
	{8'd62,8'd91} : s = 153;
	{8'd62,8'd92} : s = 154;
	{8'd62,8'd93} : s = 155;
	{8'd62,8'd94} : s = 156;
	{8'd62,8'd95} : s = 157;
	{8'd62,8'd96} : s = 158;
	{8'd62,8'd97} : s = 159;
	{8'd62,8'd98} : s = 160;
	{8'd62,8'd99} : s = 161;
	{8'd62,8'd100} : s = 162;
	{8'd62,8'd101} : s = 163;
	{8'd62,8'd102} : s = 164;
	{8'd62,8'd103} : s = 165;
	{8'd62,8'd104} : s = 166;
	{8'd62,8'd105} : s = 167;
	{8'd62,8'd106} : s = 168;
	{8'd62,8'd107} : s = 169;
	{8'd62,8'd108} : s = 170;
	{8'd62,8'd109} : s = 171;
	{8'd62,8'd110} : s = 172;
	{8'd62,8'd111} : s = 173;
	{8'd62,8'd112} : s = 174;
	{8'd62,8'd113} : s = 175;
	{8'd62,8'd114} : s = 176;
	{8'd62,8'd115} : s = 177;
	{8'd62,8'd116} : s = 178;
	{8'd62,8'd117} : s = 179;
	{8'd62,8'd118} : s = 180;
	{8'd62,8'd119} : s = 181;
	{8'd62,8'd120} : s = 182;
	{8'd62,8'd121} : s = 183;
	{8'd62,8'd122} : s = 184;
	{8'd62,8'd123} : s = 185;
	{8'd62,8'd124} : s = 186;
	{8'd62,8'd125} : s = 187;
	{8'd62,8'd126} : s = 188;
	{8'd62,8'd127} : s = 189;
	{8'd62,8'd128} : s = 190;
	{8'd62,8'd129} : s = 191;
	{8'd62,8'd130} : s = 192;
	{8'd62,8'd131} : s = 193;
	{8'd62,8'd132} : s = 194;
	{8'd62,8'd133} : s = 195;
	{8'd62,8'd134} : s = 196;
	{8'd62,8'd135} : s = 197;
	{8'd62,8'd136} : s = 198;
	{8'd62,8'd137} : s = 199;
	{8'd62,8'd138} : s = 200;
	{8'd62,8'd139} : s = 201;
	{8'd62,8'd140} : s = 202;
	{8'd62,8'd141} : s = 203;
	{8'd62,8'd142} : s = 204;
	{8'd62,8'd143} : s = 205;
	{8'd62,8'd144} : s = 206;
	{8'd62,8'd145} : s = 207;
	{8'd62,8'd146} : s = 208;
	{8'd62,8'd147} : s = 209;
	{8'd62,8'd148} : s = 210;
	{8'd62,8'd149} : s = 211;
	{8'd62,8'd150} : s = 212;
	{8'd62,8'd151} : s = 213;
	{8'd62,8'd152} : s = 214;
	{8'd62,8'd153} : s = 215;
	{8'd62,8'd154} : s = 216;
	{8'd62,8'd155} : s = 217;
	{8'd62,8'd156} : s = 218;
	{8'd62,8'd157} : s = 219;
	{8'd62,8'd158} : s = 220;
	{8'd62,8'd159} : s = 221;
	{8'd62,8'd160} : s = 222;
	{8'd62,8'd161} : s = 223;
	{8'd62,8'd162} : s = 224;
	{8'd62,8'd163} : s = 225;
	{8'd62,8'd164} : s = 226;
	{8'd62,8'd165} : s = 227;
	{8'd62,8'd166} : s = 228;
	{8'd62,8'd167} : s = 229;
	{8'd62,8'd168} : s = 230;
	{8'd62,8'd169} : s = 231;
	{8'd62,8'd170} : s = 232;
	{8'd62,8'd171} : s = 233;
	{8'd62,8'd172} : s = 234;
	{8'd62,8'd173} : s = 235;
	{8'd62,8'd174} : s = 236;
	{8'd62,8'd175} : s = 237;
	{8'd62,8'd176} : s = 238;
	{8'd62,8'd177} : s = 239;
	{8'd62,8'd178} : s = 240;
	{8'd62,8'd179} : s = 241;
	{8'd62,8'd180} : s = 242;
	{8'd62,8'd181} : s = 243;
	{8'd62,8'd182} : s = 244;
	{8'd62,8'd183} : s = 245;
	{8'd62,8'd184} : s = 246;
	{8'd62,8'd185} : s = 247;
	{8'd62,8'd186} : s = 248;
	{8'd62,8'd187} : s = 249;
	{8'd62,8'd188} : s = 250;
	{8'd62,8'd189} : s = 251;
	{8'd62,8'd190} : s = 252;
	{8'd62,8'd191} : s = 253;
	{8'd62,8'd192} : s = 254;
	{8'd62,8'd193} : s = 255;
	{8'd62,8'd194} : s = 256;
	{8'd62,8'd195} : s = 257;
	{8'd62,8'd196} : s = 258;
	{8'd62,8'd197} : s = 259;
	{8'd62,8'd198} : s = 260;
	{8'd62,8'd199} : s = 261;
	{8'd62,8'd200} : s = 262;
	{8'd62,8'd201} : s = 263;
	{8'd62,8'd202} : s = 264;
	{8'd62,8'd203} : s = 265;
	{8'd62,8'd204} : s = 266;
	{8'd62,8'd205} : s = 267;
	{8'd62,8'd206} : s = 268;
	{8'd62,8'd207} : s = 269;
	{8'd62,8'd208} : s = 270;
	{8'd62,8'd209} : s = 271;
	{8'd62,8'd210} : s = 272;
	{8'd62,8'd211} : s = 273;
	{8'd62,8'd212} : s = 274;
	{8'd62,8'd213} : s = 275;
	{8'd62,8'd214} : s = 276;
	{8'd62,8'd215} : s = 277;
	{8'd62,8'd216} : s = 278;
	{8'd62,8'd217} : s = 279;
	{8'd62,8'd218} : s = 280;
	{8'd62,8'd219} : s = 281;
	{8'd62,8'd220} : s = 282;
	{8'd62,8'd221} : s = 283;
	{8'd62,8'd222} : s = 284;
	{8'd62,8'd223} : s = 285;
	{8'd62,8'd224} : s = 286;
	{8'd62,8'd225} : s = 287;
	{8'd62,8'd226} : s = 288;
	{8'd62,8'd227} : s = 289;
	{8'd62,8'd228} : s = 290;
	{8'd62,8'd229} : s = 291;
	{8'd62,8'd230} : s = 292;
	{8'd62,8'd231} : s = 293;
	{8'd62,8'd232} : s = 294;
	{8'd62,8'd233} : s = 295;
	{8'd62,8'd234} : s = 296;
	{8'd62,8'd235} : s = 297;
	{8'd62,8'd236} : s = 298;
	{8'd62,8'd237} : s = 299;
	{8'd62,8'd238} : s = 300;
	{8'd62,8'd239} : s = 301;
	{8'd62,8'd240} : s = 302;
	{8'd62,8'd241} : s = 303;
	{8'd62,8'd242} : s = 304;
	{8'd62,8'd243} : s = 305;
	{8'd62,8'd244} : s = 306;
	{8'd62,8'd245} : s = 307;
	{8'd62,8'd246} : s = 308;
	{8'd62,8'd247} : s = 309;
	{8'd62,8'd248} : s = 310;
	{8'd62,8'd249} : s = 311;
	{8'd62,8'd250} : s = 312;
	{8'd62,8'd251} : s = 313;
	{8'd62,8'd252} : s = 314;
	{8'd62,8'd253} : s = 315;
	{8'd62,8'd254} : s = 316;
	{8'd62,8'd255} : s = 317;
	{8'd63,8'd0} : s = 63;
	{8'd63,8'd1} : s = 64;
	{8'd63,8'd2} : s = 65;
	{8'd63,8'd3} : s = 66;
	{8'd63,8'd4} : s = 67;
	{8'd63,8'd5} : s = 68;
	{8'd63,8'd6} : s = 69;
	{8'd63,8'd7} : s = 70;
	{8'd63,8'd8} : s = 71;
	{8'd63,8'd9} : s = 72;
	{8'd63,8'd10} : s = 73;
	{8'd63,8'd11} : s = 74;
	{8'd63,8'd12} : s = 75;
	{8'd63,8'd13} : s = 76;
	{8'd63,8'd14} : s = 77;
	{8'd63,8'd15} : s = 78;
	{8'd63,8'd16} : s = 79;
	{8'd63,8'd17} : s = 80;
	{8'd63,8'd18} : s = 81;
	{8'd63,8'd19} : s = 82;
	{8'd63,8'd20} : s = 83;
	{8'd63,8'd21} : s = 84;
	{8'd63,8'd22} : s = 85;
	{8'd63,8'd23} : s = 86;
	{8'd63,8'd24} : s = 87;
	{8'd63,8'd25} : s = 88;
	{8'd63,8'd26} : s = 89;
	{8'd63,8'd27} : s = 90;
	{8'd63,8'd28} : s = 91;
	{8'd63,8'd29} : s = 92;
	{8'd63,8'd30} : s = 93;
	{8'd63,8'd31} : s = 94;
	{8'd63,8'd32} : s = 95;
	{8'd63,8'd33} : s = 96;
	{8'd63,8'd34} : s = 97;
	{8'd63,8'd35} : s = 98;
	{8'd63,8'd36} : s = 99;
	{8'd63,8'd37} : s = 100;
	{8'd63,8'd38} : s = 101;
	{8'd63,8'd39} : s = 102;
	{8'd63,8'd40} : s = 103;
	{8'd63,8'd41} : s = 104;
	{8'd63,8'd42} : s = 105;
	{8'd63,8'd43} : s = 106;
	{8'd63,8'd44} : s = 107;
	{8'd63,8'd45} : s = 108;
	{8'd63,8'd46} : s = 109;
	{8'd63,8'd47} : s = 110;
	{8'd63,8'd48} : s = 111;
	{8'd63,8'd49} : s = 112;
	{8'd63,8'd50} : s = 113;
	{8'd63,8'd51} : s = 114;
	{8'd63,8'd52} : s = 115;
	{8'd63,8'd53} : s = 116;
	{8'd63,8'd54} : s = 117;
	{8'd63,8'd55} : s = 118;
	{8'd63,8'd56} : s = 119;
	{8'd63,8'd57} : s = 120;
	{8'd63,8'd58} : s = 121;
	{8'd63,8'd59} : s = 122;
	{8'd63,8'd60} : s = 123;
	{8'd63,8'd61} : s = 124;
	{8'd63,8'd62} : s = 125;
	{8'd63,8'd63} : s = 126;
	{8'd63,8'd64} : s = 127;
	{8'd63,8'd65} : s = 128;
	{8'd63,8'd66} : s = 129;
	{8'd63,8'd67} : s = 130;
	{8'd63,8'd68} : s = 131;
	{8'd63,8'd69} : s = 132;
	{8'd63,8'd70} : s = 133;
	{8'd63,8'd71} : s = 134;
	{8'd63,8'd72} : s = 135;
	{8'd63,8'd73} : s = 136;
	{8'd63,8'd74} : s = 137;
	{8'd63,8'd75} : s = 138;
	{8'd63,8'd76} : s = 139;
	{8'd63,8'd77} : s = 140;
	{8'd63,8'd78} : s = 141;
	{8'd63,8'd79} : s = 142;
	{8'd63,8'd80} : s = 143;
	{8'd63,8'd81} : s = 144;
	{8'd63,8'd82} : s = 145;
	{8'd63,8'd83} : s = 146;
	{8'd63,8'd84} : s = 147;
	{8'd63,8'd85} : s = 148;
	{8'd63,8'd86} : s = 149;
	{8'd63,8'd87} : s = 150;
	{8'd63,8'd88} : s = 151;
	{8'd63,8'd89} : s = 152;
	{8'd63,8'd90} : s = 153;
	{8'd63,8'd91} : s = 154;
	{8'd63,8'd92} : s = 155;
	{8'd63,8'd93} : s = 156;
	{8'd63,8'd94} : s = 157;
	{8'd63,8'd95} : s = 158;
	{8'd63,8'd96} : s = 159;
	{8'd63,8'd97} : s = 160;
	{8'd63,8'd98} : s = 161;
	{8'd63,8'd99} : s = 162;
	{8'd63,8'd100} : s = 163;
	{8'd63,8'd101} : s = 164;
	{8'd63,8'd102} : s = 165;
	{8'd63,8'd103} : s = 166;
	{8'd63,8'd104} : s = 167;
	{8'd63,8'd105} : s = 168;
	{8'd63,8'd106} : s = 169;
	{8'd63,8'd107} : s = 170;
	{8'd63,8'd108} : s = 171;
	{8'd63,8'd109} : s = 172;
	{8'd63,8'd110} : s = 173;
	{8'd63,8'd111} : s = 174;
	{8'd63,8'd112} : s = 175;
	{8'd63,8'd113} : s = 176;
	{8'd63,8'd114} : s = 177;
	{8'd63,8'd115} : s = 178;
	{8'd63,8'd116} : s = 179;
	{8'd63,8'd117} : s = 180;
	{8'd63,8'd118} : s = 181;
	{8'd63,8'd119} : s = 182;
	{8'd63,8'd120} : s = 183;
	{8'd63,8'd121} : s = 184;
	{8'd63,8'd122} : s = 185;
	{8'd63,8'd123} : s = 186;
	{8'd63,8'd124} : s = 187;
	{8'd63,8'd125} : s = 188;
	{8'd63,8'd126} : s = 189;
	{8'd63,8'd127} : s = 190;
	{8'd63,8'd128} : s = 191;
	{8'd63,8'd129} : s = 192;
	{8'd63,8'd130} : s = 193;
	{8'd63,8'd131} : s = 194;
	{8'd63,8'd132} : s = 195;
	{8'd63,8'd133} : s = 196;
	{8'd63,8'd134} : s = 197;
	{8'd63,8'd135} : s = 198;
	{8'd63,8'd136} : s = 199;
	{8'd63,8'd137} : s = 200;
	{8'd63,8'd138} : s = 201;
	{8'd63,8'd139} : s = 202;
	{8'd63,8'd140} : s = 203;
	{8'd63,8'd141} : s = 204;
	{8'd63,8'd142} : s = 205;
	{8'd63,8'd143} : s = 206;
	{8'd63,8'd144} : s = 207;
	{8'd63,8'd145} : s = 208;
	{8'd63,8'd146} : s = 209;
	{8'd63,8'd147} : s = 210;
	{8'd63,8'd148} : s = 211;
	{8'd63,8'd149} : s = 212;
	{8'd63,8'd150} : s = 213;
	{8'd63,8'd151} : s = 214;
	{8'd63,8'd152} : s = 215;
	{8'd63,8'd153} : s = 216;
	{8'd63,8'd154} : s = 217;
	{8'd63,8'd155} : s = 218;
	{8'd63,8'd156} : s = 219;
	{8'd63,8'd157} : s = 220;
	{8'd63,8'd158} : s = 221;
	{8'd63,8'd159} : s = 222;
	{8'd63,8'd160} : s = 223;
	{8'd63,8'd161} : s = 224;
	{8'd63,8'd162} : s = 225;
	{8'd63,8'd163} : s = 226;
	{8'd63,8'd164} : s = 227;
	{8'd63,8'd165} : s = 228;
	{8'd63,8'd166} : s = 229;
	{8'd63,8'd167} : s = 230;
	{8'd63,8'd168} : s = 231;
	{8'd63,8'd169} : s = 232;
	{8'd63,8'd170} : s = 233;
	{8'd63,8'd171} : s = 234;
	{8'd63,8'd172} : s = 235;
	{8'd63,8'd173} : s = 236;
	{8'd63,8'd174} : s = 237;
	{8'd63,8'd175} : s = 238;
	{8'd63,8'd176} : s = 239;
	{8'd63,8'd177} : s = 240;
	{8'd63,8'd178} : s = 241;
	{8'd63,8'd179} : s = 242;
	{8'd63,8'd180} : s = 243;
	{8'd63,8'd181} : s = 244;
	{8'd63,8'd182} : s = 245;
	{8'd63,8'd183} : s = 246;
	{8'd63,8'd184} : s = 247;
	{8'd63,8'd185} : s = 248;
	{8'd63,8'd186} : s = 249;
	{8'd63,8'd187} : s = 250;
	{8'd63,8'd188} : s = 251;
	{8'd63,8'd189} : s = 252;
	{8'd63,8'd190} : s = 253;
	{8'd63,8'd191} : s = 254;
	{8'd63,8'd192} : s = 255;
	{8'd63,8'd193} : s = 256;
	{8'd63,8'd194} : s = 257;
	{8'd63,8'd195} : s = 258;
	{8'd63,8'd196} : s = 259;
	{8'd63,8'd197} : s = 260;
	{8'd63,8'd198} : s = 261;
	{8'd63,8'd199} : s = 262;
	{8'd63,8'd200} : s = 263;
	{8'd63,8'd201} : s = 264;
	{8'd63,8'd202} : s = 265;
	{8'd63,8'd203} : s = 266;
	{8'd63,8'd204} : s = 267;
	{8'd63,8'd205} : s = 268;
	{8'd63,8'd206} : s = 269;
	{8'd63,8'd207} : s = 270;
	{8'd63,8'd208} : s = 271;
	{8'd63,8'd209} : s = 272;
	{8'd63,8'd210} : s = 273;
	{8'd63,8'd211} : s = 274;
	{8'd63,8'd212} : s = 275;
	{8'd63,8'd213} : s = 276;
	{8'd63,8'd214} : s = 277;
	{8'd63,8'd215} : s = 278;
	{8'd63,8'd216} : s = 279;
	{8'd63,8'd217} : s = 280;
	{8'd63,8'd218} : s = 281;
	{8'd63,8'd219} : s = 282;
	{8'd63,8'd220} : s = 283;
	{8'd63,8'd221} : s = 284;
	{8'd63,8'd222} : s = 285;
	{8'd63,8'd223} : s = 286;
	{8'd63,8'd224} : s = 287;
	{8'd63,8'd225} : s = 288;
	{8'd63,8'd226} : s = 289;
	{8'd63,8'd227} : s = 290;
	{8'd63,8'd228} : s = 291;
	{8'd63,8'd229} : s = 292;
	{8'd63,8'd230} : s = 293;
	{8'd63,8'd231} : s = 294;
	{8'd63,8'd232} : s = 295;
	{8'd63,8'd233} : s = 296;
	{8'd63,8'd234} : s = 297;
	{8'd63,8'd235} : s = 298;
	{8'd63,8'd236} : s = 299;
	{8'd63,8'd237} : s = 300;
	{8'd63,8'd238} : s = 301;
	{8'd63,8'd239} : s = 302;
	{8'd63,8'd240} : s = 303;
	{8'd63,8'd241} : s = 304;
	{8'd63,8'd242} : s = 305;
	{8'd63,8'd243} : s = 306;
	{8'd63,8'd244} : s = 307;
	{8'd63,8'd245} : s = 308;
	{8'd63,8'd246} : s = 309;
	{8'd63,8'd247} : s = 310;
	{8'd63,8'd248} : s = 311;
	{8'd63,8'd249} : s = 312;
	{8'd63,8'd250} : s = 313;
	{8'd63,8'd251} : s = 314;
	{8'd63,8'd252} : s = 315;
	{8'd63,8'd253} : s = 316;
	{8'd63,8'd254} : s = 317;
	{8'd63,8'd255} : s = 318;
	{8'd64,8'd0} : s = 64;
	{8'd64,8'd1} : s = 65;
	{8'd64,8'd2} : s = 66;
	{8'd64,8'd3} : s = 67;
	{8'd64,8'd4} : s = 68;
	{8'd64,8'd5} : s = 69;
	{8'd64,8'd6} : s = 70;
	{8'd64,8'd7} : s = 71;
	{8'd64,8'd8} : s = 72;
	{8'd64,8'd9} : s = 73;
	{8'd64,8'd10} : s = 74;
	{8'd64,8'd11} : s = 75;
	{8'd64,8'd12} : s = 76;
	{8'd64,8'd13} : s = 77;
	{8'd64,8'd14} : s = 78;
	{8'd64,8'd15} : s = 79;
	{8'd64,8'd16} : s = 80;
	{8'd64,8'd17} : s = 81;
	{8'd64,8'd18} : s = 82;
	{8'd64,8'd19} : s = 83;
	{8'd64,8'd20} : s = 84;
	{8'd64,8'd21} : s = 85;
	{8'd64,8'd22} : s = 86;
	{8'd64,8'd23} : s = 87;
	{8'd64,8'd24} : s = 88;
	{8'd64,8'd25} : s = 89;
	{8'd64,8'd26} : s = 90;
	{8'd64,8'd27} : s = 91;
	{8'd64,8'd28} : s = 92;
	{8'd64,8'd29} : s = 93;
	{8'd64,8'd30} : s = 94;
	{8'd64,8'd31} : s = 95;
	{8'd64,8'd32} : s = 96;
	{8'd64,8'd33} : s = 97;
	{8'd64,8'd34} : s = 98;
	{8'd64,8'd35} : s = 99;
	{8'd64,8'd36} : s = 100;
	{8'd64,8'd37} : s = 101;
	{8'd64,8'd38} : s = 102;
	{8'd64,8'd39} : s = 103;
	{8'd64,8'd40} : s = 104;
	{8'd64,8'd41} : s = 105;
	{8'd64,8'd42} : s = 106;
	{8'd64,8'd43} : s = 107;
	{8'd64,8'd44} : s = 108;
	{8'd64,8'd45} : s = 109;
	{8'd64,8'd46} : s = 110;
	{8'd64,8'd47} : s = 111;
	{8'd64,8'd48} : s = 112;
	{8'd64,8'd49} : s = 113;
	{8'd64,8'd50} : s = 114;
	{8'd64,8'd51} : s = 115;
	{8'd64,8'd52} : s = 116;
	{8'd64,8'd53} : s = 117;
	{8'd64,8'd54} : s = 118;
	{8'd64,8'd55} : s = 119;
	{8'd64,8'd56} : s = 120;
	{8'd64,8'd57} : s = 121;
	{8'd64,8'd58} : s = 122;
	{8'd64,8'd59} : s = 123;
	{8'd64,8'd60} : s = 124;
	{8'd64,8'd61} : s = 125;
	{8'd64,8'd62} : s = 126;
	{8'd64,8'd63} : s = 127;
	{8'd64,8'd64} : s = 128;
	{8'd64,8'd65} : s = 129;
	{8'd64,8'd66} : s = 130;
	{8'd64,8'd67} : s = 131;
	{8'd64,8'd68} : s = 132;
	{8'd64,8'd69} : s = 133;
	{8'd64,8'd70} : s = 134;
	{8'd64,8'd71} : s = 135;
	{8'd64,8'd72} : s = 136;
	{8'd64,8'd73} : s = 137;
	{8'd64,8'd74} : s = 138;
	{8'd64,8'd75} : s = 139;
	{8'd64,8'd76} : s = 140;
	{8'd64,8'd77} : s = 141;
	{8'd64,8'd78} : s = 142;
	{8'd64,8'd79} : s = 143;
	{8'd64,8'd80} : s = 144;
	{8'd64,8'd81} : s = 145;
	{8'd64,8'd82} : s = 146;
	{8'd64,8'd83} : s = 147;
	{8'd64,8'd84} : s = 148;
	{8'd64,8'd85} : s = 149;
	{8'd64,8'd86} : s = 150;
	{8'd64,8'd87} : s = 151;
	{8'd64,8'd88} : s = 152;
	{8'd64,8'd89} : s = 153;
	{8'd64,8'd90} : s = 154;
	{8'd64,8'd91} : s = 155;
	{8'd64,8'd92} : s = 156;
	{8'd64,8'd93} : s = 157;
	{8'd64,8'd94} : s = 158;
	{8'd64,8'd95} : s = 159;
	{8'd64,8'd96} : s = 160;
	{8'd64,8'd97} : s = 161;
	{8'd64,8'd98} : s = 162;
	{8'd64,8'd99} : s = 163;
	{8'd64,8'd100} : s = 164;
	{8'd64,8'd101} : s = 165;
	{8'd64,8'd102} : s = 166;
	{8'd64,8'd103} : s = 167;
	{8'd64,8'd104} : s = 168;
	{8'd64,8'd105} : s = 169;
	{8'd64,8'd106} : s = 170;
	{8'd64,8'd107} : s = 171;
	{8'd64,8'd108} : s = 172;
	{8'd64,8'd109} : s = 173;
	{8'd64,8'd110} : s = 174;
	{8'd64,8'd111} : s = 175;
	{8'd64,8'd112} : s = 176;
	{8'd64,8'd113} : s = 177;
	{8'd64,8'd114} : s = 178;
	{8'd64,8'd115} : s = 179;
	{8'd64,8'd116} : s = 180;
	{8'd64,8'd117} : s = 181;
	{8'd64,8'd118} : s = 182;
	{8'd64,8'd119} : s = 183;
	{8'd64,8'd120} : s = 184;
	{8'd64,8'd121} : s = 185;
	{8'd64,8'd122} : s = 186;
	{8'd64,8'd123} : s = 187;
	{8'd64,8'd124} : s = 188;
	{8'd64,8'd125} : s = 189;
	{8'd64,8'd126} : s = 190;
	{8'd64,8'd127} : s = 191;
	{8'd64,8'd128} : s = 192;
	{8'd64,8'd129} : s = 193;
	{8'd64,8'd130} : s = 194;
	{8'd64,8'd131} : s = 195;
	{8'd64,8'd132} : s = 196;
	{8'd64,8'd133} : s = 197;
	{8'd64,8'd134} : s = 198;
	{8'd64,8'd135} : s = 199;
	{8'd64,8'd136} : s = 200;
	{8'd64,8'd137} : s = 201;
	{8'd64,8'd138} : s = 202;
	{8'd64,8'd139} : s = 203;
	{8'd64,8'd140} : s = 204;
	{8'd64,8'd141} : s = 205;
	{8'd64,8'd142} : s = 206;
	{8'd64,8'd143} : s = 207;
	{8'd64,8'd144} : s = 208;
	{8'd64,8'd145} : s = 209;
	{8'd64,8'd146} : s = 210;
	{8'd64,8'd147} : s = 211;
	{8'd64,8'd148} : s = 212;
	{8'd64,8'd149} : s = 213;
	{8'd64,8'd150} : s = 214;
	{8'd64,8'd151} : s = 215;
	{8'd64,8'd152} : s = 216;
	{8'd64,8'd153} : s = 217;
	{8'd64,8'd154} : s = 218;
	{8'd64,8'd155} : s = 219;
	{8'd64,8'd156} : s = 220;
	{8'd64,8'd157} : s = 221;
	{8'd64,8'd158} : s = 222;
	{8'd64,8'd159} : s = 223;
	{8'd64,8'd160} : s = 224;
	{8'd64,8'd161} : s = 225;
	{8'd64,8'd162} : s = 226;
	{8'd64,8'd163} : s = 227;
	{8'd64,8'd164} : s = 228;
	{8'd64,8'd165} : s = 229;
	{8'd64,8'd166} : s = 230;
	{8'd64,8'd167} : s = 231;
	{8'd64,8'd168} : s = 232;
	{8'd64,8'd169} : s = 233;
	{8'd64,8'd170} : s = 234;
	{8'd64,8'd171} : s = 235;
	{8'd64,8'd172} : s = 236;
	{8'd64,8'd173} : s = 237;
	{8'd64,8'd174} : s = 238;
	{8'd64,8'd175} : s = 239;
	{8'd64,8'd176} : s = 240;
	{8'd64,8'd177} : s = 241;
	{8'd64,8'd178} : s = 242;
	{8'd64,8'd179} : s = 243;
	{8'd64,8'd180} : s = 244;
	{8'd64,8'd181} : s = 245;
	{8'd64,8'd182} : s = 246;
	{8'd64,8'd183} : s = 247;
	{8'd64,8'd184} : s = 248;
	{8'd64,8'd185} : s = 249;
	{8'd64,8'd186} : s = 250;
	{8'd64,8'd187} : s = 251;
	{8'd64,8'd188} : s = 252;
	{8'd64,8'd189} : s = 253;
	{8'd64,8'd190} : s = 254;
	{8'd64,8'd191} : s = 255;
	{8'd64,8'd192} : s = 256;
	{8'd64,8'd193} : s = 257;
	{8'd64,8'd194} : s = 258;
	{8'd64,8'd195} : s = 259;
	{8'd64,8'd196} : s = 260;
	{8'd64,8'd197} : s = 261;
	{8'd64,8'd198} : s = 262;
	{8'd64,8'd199} : s = 263;
	{8'd64,8'd200} : s = 264;
	{8'd64,8'd201} : s = 265;
	{8'd64,8'd202} : s = 266;
	{8'd64,8'd203} : s = 267;
	{8'd64,8'd204} : s = 268;
	{8'd64,8'd205} : s = 269;
	{8'd64,8'd206} : s = 270;
	{8'd64,8'd207} : s = 271;
	{8'd64,8'd208} : s = 272;
	{8'd64,8'd209} : s = 273;
	{8'd64,8'd210} : s = 274;
	{8'd64,8'd211} : s = 275;
	{8'd64,8'd212} : s = 276;
	{8'd64,8'd213} : s = 277;
	{8'd64,8'd214} : s = 278;
	{8'd64,8'd215} : s = 279;
	{8'd64,8'd216} : s = 280;
	{8'd64,8'd217} : s = 281;
	{8'd64,8'd218} : s = 282;
	{8'd64,8'd219} : s = 283;
	{8'd64,8'd220} : s = 284;
	{8'd64,8'd221} : s = 285;
	{8'd64,8'd222} : s = 286;
	{8'd64,8'd223} : s = 287;
	{8'd64,8'd224} : s = 288;
	{8'd64,8'd225} : s = 289;
	{8'd64,8'd226} : s = 290;
	{8'd64,8'd227} : s = 291;
	{8'd64,8'd228} : s = 292;
	{8'd64,8'd229} : s = 293;
	{8'd64,8'd230} : s = 294;
	{8'd64,8'd231} : s = 295;
	{8'd64,8'd232} : s = 296;
	{8'd64,8'd233} : s = 297;
	{8'd64,8'd234} : s = 298;
	{8'd64,8'd235} : s = 299;
	{8'd64,8'd236} : s = 300;
	{8'd64,8'd237} : s = 301;
	{8'd64,8'd238} : s = 302;
	{8'd64,8'd239} : s = 303;
	{8'd64,8'd240} : s = 304;
	{8'd64,8'd241} : s = 305;
	{8'd64,8'd242} : s = 306;
	{8'd64,8'd243} : s = 307;
	{8'd64,8'd244} : s = 308;
	{8'd64,8'd245} : s = 309;
	{8'd64,8'd246} : s = 310;
	{8'd64,8'd247} : s = 311;
	{8'd64,8'd248} : s = 312;
	{8'd64,8'd249} : s = 313;
	{8'd64,8'd250} : s = 314;
	{8'd64,8'd251} : s = 315;
	{8'd64,8'd252} : s = 316;
	{8'd64,8'd253} : s = 317;
	{8'd64,8'd254} : s = 318;
	{8'd64,8'd255} : s = 319;
	{8'd65,8'd0} : s = 65;
	{8'd65,8'd1} : s = 66;
	{8'd65,8'd2} : s = 67;
	{8'd65,8'd3} : s = 68;
	{8'd65,8'd4} : s = 69;
	{8'd65,8'd5} : s = 70;
	{8'd65,8'd6} : s = 71;
	{8'd65,8'd7} : s = 72;
	{8'd65,8'd8} : s = 73;
	{8'd65,8'd9} : s = 74;
	{8'd65,8'd10} : s = 75;
	{8'd65,8'd11} : s = 76;
	{8'd65,8'd12} : s = 77;
	{8'd65,8'd13} : s = 78;
	{8'd65,8'd14} : s = 79;
	{8'd65,8'd15} : s = 80;
	{8'd65,8'd16} : s = 81;
	{8'd65,8'd17} : s = 82;
	{8'd65,8'd18} : s = 83;
	{8'd65,8'd19} : s = 84;
	{8'd65,8'd20} : s = 85;
	{8'd65,8'd21} : s = 86;
	{8'd65,8'd22} : s = 87;
	{8'd65,8'd23} : s = 88;
	{8'd65,8'd24} : s = 89;
	{8'd65,8'd25} : s = 90;
	{8'd65,8'd26} : s = 91;
	{8'd65,8'd27} : s = 92;
	{8'd65,8'd28} : s = 93;
	{8'd65,8'd29} : s = 94;
	{8'd65,8'd30} : s = 95;
	{8'd65,8'd31} : s = 96;
	{8'd65,8'd32} : s = 97;
	{8'd65,8'd33} : s = 98;
	{8'd65,8'd34} : s = 99;
	{8'd65,8'd35} : s = 100;
	{8'd65,8'd36} : s = 101;
	{8'd65,8'd37} : s = 102;
	{8'd65,8'd38} : s = 103;
	{8'd65,8'd39} : s = 104;
	{8'd65,8'd40} : s = 105;
	{8'd65,8'd41} : s = 106;
	{8'd65,8'd42} : s = 107;
	{8'd65,8'd43} : s = 108;
	{8'd65,8'd44} : s = 109;
	{8'd65,8'd45} : s = 110;
	{8'd65,8'd46} : s = 111;
	{8'd65,8'd47} : s = 112;
	{8'd65,8'd48} : s = 113;
	{8'd65,8'd49} : s = 114;
	{8'd65,8'd50} : s = 115;
	{8'd65,8'd51} : s = 116;
	{8'd65,8'd52} : s = 117;
	{8'd65,8'd53} : s = 118;
	{8'd65,8'd54} : s = 119;
	{8'd65,8'd55} : s = 120;
	{8'd65,8'd56} : s = 121;
	{8'd65,8'd57} : s = 122;
	{8'd65,8'd58} : s = 123;
	{8'd65,8'd59} : s = 124;
	{8'd65,8'd60} : s = 125;
	{8'd65,8'd61} : s = 126;
	{8'd65,8'd62} : s = 127;
	{8'd65,8'd63} : s = 128;
	{8'd65,8'd64} : s = 129;
	{8'd65,8'd65} : s = 130;
	{8'd65,8'd66} : s = 131;
	{8'd65,8'd67} : s = 132;
	{8'd65,8'd68} : s = 133;
	{8'd65,8'd69} : s = 134;
	{8'd65,8'd70} : s = 135;
	{8'd65,8'd71} : s = 136;
	{8'd65,8'd72} : s = 137;
	{8'd65,8'd73} : s = 138;
	{8'd65,8'd74} : s = 139;
	{8'd65,8'd75} : s = 140;
	{8'd65,8'd76} : s = 141;
	{8'd65,8'd77} : s = 142;
	{8'd65,8'd78} : s = 143;
	{8'd65,8'd79} : s = 144;
	{8'd65,8'd80} : s = 145;
	{8'd65,8'd81} : s = 146;
	{8'd65,8'd82} : s = 147;
	{8'd65,8'd83} : s = 148;
	{8'd65,8'd84} : s = 149;
	{8'd65,8'd85} : s = 150;
	{8'd65,8'd86} : s = 151;
	{8'd65,8'd87} : s = 152;
	{8'd65,8'd88} : s = 153;
	{8'd65,8'd89} : s = 154;
	{8'd65,8'd90} : s = 155;
	{8'd65,8'd91} : s = 156;
	{8'd65,8'd92} : s = 157;
	{8'd65,8'd93} : s = 158;
	{8'd65,8'd94} : s = 159;
	{8'd65,8'd95} : s = 160;
	{8'd65,8'd96} : s = 161;
	{8'd65,8'd97} : s = 162;
	{8'd65,8'd98} : s = 163;
	{8'd65,8'd99} : s = 164;
	{8'd65,8'd100} : s = 165;
	{8'd65,8'd101} : s = 166;
	{8'd65,8'd102} : s = 167;
	{8'd65,8'd103} : s = 168;
	{8'd65,8'd104} : s = 169;
	{8'd65,8'd105} : s = 170;
	{8'd65,8'd106} : s = 171;
	{8'd65,8'd107} : s = 172;
	{8'd65,8'd108} : s = 173;
	{8'd65,8'd109} : s = 174;
	{8'd65,8'd110} : s = 175;
	{8'd65,8'd111} : s = 176;
	{8'd65,8'd112} : s = 177;
	{8'd65,8'd113} : s = 178;
	{8'd65,8'd114} : s = 179;
	{8'd65,8'd115} : s = 180;
	{8'd65,8'd116} : s = 181;
	{8'd65,8'd117} : s = 182;
	{8'd65,8'd118} : s = 183;
	{8'd65,8'd119} : s = 184;
	{8'd65,8'd120} : s = 185;
	{8'd65,8'd121} : s = 186;
	{8'd65,8'd122} : s = 187;
	{8'd65,8'd123} : s = 188;
	{8'd65,8'd124} : s = 189;
	{8'd65,8'd125} : s = 190;
	{8'd65,8'd126} : s = 191;
	{8'd65,8'd127} : s = 192;
	{8'd65,8'd128} : s = 193;
	{8'd65,8'd129} : s = 194;
	{8'd65,8'd130} : s = 195;
	{8'd65,8'd131} : s = 196;
	{8'd65,8'd132} : s = 197;
	{8'd65,8'd133} : s = 198;
	{8'd65,8'd134} : s = 199;
	{8'd65,8'd135} : s = 200;
	{8'd65,8'd136} : s = 201;
	{8'd65,8'd137} : s = 202;
	{8'd65,8'd138} : s = 203;
	{8'd65,8'd139} : s = 204;
	{8'd65,8'd140} : s = 205;
	{8'd65,8'd141} : s = 206;
	{8'd65,8'd142} : s = 207;
	{8'd65,8'd143} : s = 208;
	{8'd65,8'd144} : s = 209;
	{8'd65,8'd145} : s = 210;
	{8'd65,8'd146} : s = 211;
	{8'd65,8'd147} : s = 212;
	{8'd65,8'd148} : s = 213;
	{8'd65,8'd149} : s = 214;
	{8'd65,8'd150} : s = 215;
	{8'd65,8'd151} : s = 216;
	{8'd65,8'd152} : s = 217;
	{8'd65,8'd153} : s = 218;
	{8'd65,8'd154} : s = 219;
	{8'd65,8'd155} : s = 220;
	{8'd65,8'd156} : s = 221;
	{8'd65,8'd157} : s = 222;
	{8'd65,8'd158} : s = 223;
	{8'd65,8'd159} : s = 224;
	{8'd65,8'd160} : s = 225;
	{8'd65,8'd161} : s = 226;
	{8'd65,8'd162} : s = 227;
	{8'd65,8'd163} : s = 228;
	{8'd65,8'd164} : s = 229;
	{8'd65,8'd165} : s = 230;
	{8'd65,8'd166} : s = 231;
	{8'd65,8'd167} : s = 232;
	{8'd65,8'd168} : s = 233;
	{8'd65,8'd169} : s = 234;
	{8'd65,8'd170} : s = 235;
	{8'd65,8'd171} : s = 236;
	{8'd65,8'd172} : s = 237;
	{8'd65,8'd173} : s = 238;
	{8'd65,8'd174} : s = 239;
	{8'd65,8'd175} : s = 240;
	{8'd65,8'd176} : s = 241;
	{8'd65,8'd177} : s = 242;
	{8'd65,8'd178} : s = 243;
	{8'd65,8'd179} : s = 244;
	{8'd65,8'd180} : s = 245;
	{8'd65,8'd181} : s = 246;
	{8'd65,8'd182} : s = 247;
	{8'd65,8'd183} : s = 248;
	{8'd65,8'd184} : s = 249;
	{8'd65,8'd185} : s = 250;
	{8'd65,8'd186} : s = 251;
	{8'd65,8'd187} : s = 252;
	{8'd65,8'd188} : s = 253;
	{8'd65,8'd189} : s = 254;
	{8'd65,8'd190} : s = 255;
	{8'd65,8'd191} : s = 256;
	{8'd65,8'd192} : s = 257;
	{8'd65,8'd193} : s = 258;
	{8'd65,8'd194} : s = 259;
	{8'd65,8'd195} : s = 260;
	{8'd65,8'd196} : s = 261;
	{8'd65,8'd197} : s = 262;
	{8'd65,8'd198} : s = 263;
	{8'd65,8'd199} : s = 264;
	{8'd65,8'd200} : s = 265;
	{8'd65,8'd201} : s = 266;
	{8'd65,8'd202} : s = 267;
	{8'd65,8'd203} : s = 268;
	{8'd65,8'd204} : s = 269;
	{8'd65,8'd205} : s = 270;
	{8'd65,8'd206} : s = 271;
	{8'd65,8'd207} : s = 272;
	{8'd65,8'd208} : s = 273;
	{8'd65,8'd209} : s = 274;
	{8'd65,8'd210} : s = 275;
	{8'd65,8'd211} : s = 276;
	{8'd65,8'd212} : s = 277;
	{8'd65,8'd213} : s = 278;
	{8'd65,8'd214} : s = 279;
	{8'd65,8'd215} : s = 280;
	{8'd65,8'd216} : s = 281;
	{8'd65,8'd217} : s = 282;
	{8'd65,8'd218} : s = 283;
	{8'd65,8'd219} : s = 284;
	{8'd65,8'd220} : s = 285;
	{8'd65,8'd221} : s = 286;
	{8'd65,8'd222} : s = 287;
	{8'd65,8'd223} : s = 288;
	{8'd65,8'd224} : s = 289;
	{8'd65,8'd225} : s = 290;
	{8'd65,8'd226} : s = 291;
	{8'd65,8'd227} : s = 292;
	{8'd65,8'd228} : s = 293;
	{8'd65,8'd229} : s = 294;
	{8'd65,8'd230} : s = 295;
	{8'd65,8'd231} : s = 296;
	{8'd65,8'd232} : s = 297;
	{8'd65,8'd233} : s = 298;
	{8'd65,8'd234} : s = 299;
	{8'd65,8'd235} : s = 300;
	{8'd65,8'd236} : s = 301;
	{8'd65,8'd237} : s = 302;
	{8'd65,8'd238} : s = 303;
	{8'd65,8'd239} : s = 304;
	{8'd65,8'd240} : s = 305;
	{8'd65,8'd241} : s = 306;
	{8'd65,8'd242} : s = 307;
	{8'd65,8'd243} : s = 308;
	{8'd65,8'd244} : s = 309;
	{8'd65,8'd245} : s = 310;
	{8'd65,8'd246} : s = 311;
	{8'd65,8'd247} : s = 312;
	{8'd65,8'd248} : s = 313;
	{8'd65,8'd249} : s = 314;
	{8'd65,8'd250} : s = 315;
	{8'd65,8'd251} : s = 316;
	{8'd65,8'd252} : s = 317;
	{8'd65,8'd253} : s = 318;
	{8'd65,8'd254} : s = 319;
	{8'd65,8'd255} : s = 320;
	{8'd66,8'd0} : s = 66;
	{8'd66,8'd1} : s = 67;
	{8'd66,8'd2} : s = 68;
	{8'd66,8'd3} : s = 69;
	{8'd66,8'd4} : s = 70;
	{8'd66,8'd5} : s = 71;
	{8'd66,8'd6} : s = 72;
	{8'd66,8'd7} : s = 73;
	{8'd66,8'd8} : s = 74;
	{8'd66,8'd9} : s = 75;
	{8'd66,8'd10} : s = 76;
	{8'd66,8'd11} : s = 77;
	{8'd66,8'd12} : s = 78;
	{8'd66,8'd13} : s = 79;
	{8'd66,8'd14} : s = 80;
	{8'd66,8'd15} : s = 81;
	{8'd66,8'd16} : s = 82;
	{8'd66,8'd17} : s = 83;
	{8'd66,8'd18} : s = 84;
	{8'd66,8'd19} : s = 85;
	{8'd66,8'd20} : s = 86;
	{8'd66,8'd21} : s = 87;
	{8'd66,8'd22} : s = 88;
	{8'd66,8'd23} : s = 89;
	{8'd66,8'd24} : s = 90;
	{8'd66,8'd25} : s = 91;
	{8'd66,8'd26} : s = 92;
	{8'd66,8'd27} : s = 93;
	{8'd66,8'd28} : s = 94;
	{8'd66,8'd29} : s = 95;
	{8'd66,8'd30} : s = 96;
	{8'd66,8'd31} : s = 97;
	{8'd66,8'd32} : s = 98;
	{8'd66,8'd33} : s = 99;
	{8'd66,8'd34} : s = 100;
	{8'd66,8'd35} : s = 101;
	{8'd66,8'd36} : s = 102;
	{8'd66,8'd37} : s = 103;
	{8'd66,8'd38} : s = 104;
	{8'd66,8'd39} : s = 105;
	{8'd66,8'd40} : s = 106;
	{8'd66,8'd41} : s = 107;
	{8'd66,8'd42} : s = 108;
	{8'd66,8'd43} : s = 109;
	{8'd66,8'd44} : s = 110;
	{8'd66,8'd45} : s = 111;
	{8'd66,8'd46} : s = 112;
	{8'd66,8'd47} : s = 113;
	{8'd66,8'd48} : s = 114;
	{8'd66,8'd49} : s = 115;
	{8'd66,8'd50} : s = 116;
	{8'd66,8'd51} : s = 117;
	{8'd66,8'd52} : s = 118;
	{8'd66,8'd53} : s = 119;
	{8'd66,8'd54} : s = 120;
	{8'd66,8'd55} : s = 121;
	{8'd66,8'd56} : s = 122;
	{8'd66,8'd57} : s = 123;
	{8'd66,8'd58} : s = 124;
	{8'd66,8'd59} : s = 125;
	{8'd66,8'd60} : s = 126;
	{8'd66,8'd61} : s = 127;
	{8'd66,8'd62} : s = 128;
	{8'd66,8'd63} : s = 129;
	{8'd66,8'd64} : s = 130;
	{8'd66,8'd65} : s = 131;
	{8'd66,8'd66} : s = 132;
	{8'd66,8'd67} : s = 133;
	{8'd66,8'd68} : s = 134;
	{8'd66,8'd69} : s = 135;
	{8'd66,8'd70} : s = 136;
	{8'd66,8'd71} : s = 137;
	{8'd66,8'd72} : s = 138;
	{8'd66,8'd73} : s = 139;
	{8'd66,8'd74} : s = 140;
	{8'd66,8'd75} : s = 141;
	{8'd66,8'd76} : s = 142;
	{8'd66,8'd77} : s = 143;
	{8'd66,8'd78} : s = 144;
	{8'd66,8'd79} : s = 145;
	{8'd66,8'd80} : s = 146;
	{8'd66,8'd81} : s = 147;
	{8'd66,8'd82} : s = 148;
	{8'd66,8'd83} : s = 149;
	{8'd66,8'd84} : s = 150;
	{8'd66,8'd85} : s = 151;
	{8'd66,8'd86} : s = 152;
	{8'd66,8'd87} : s = 153;
	{8'd66,8'd88} : s = 154;
	{8'd66,8'd89} : s = 155;
	{8'd66,8'd90} : s = 156;
	{8'd66,8'd91} : s = 157;
	{8'd66,8'd92} : s = 158;
	{8'd66,8'd93} : s = 159;
	{8'd66,8'd94} : s = 160;
	{8'd66,8'd95} : s = 161;
	{8'd66,8'd96} : s = 162;
	{8'd66,8'd97} : s = 163;
	{8'd66,8'd98} : s = 164;
	{8'd66,8'd99} : s = 165;
	{8'd66,8'd100} : s = 166;
	{8'd66,8'd101} : s = 167;
	{8'd66,8'd102} : s = 168;
	{8'd66,8'd103} : s = 169;
	{8'd66,8'd104} : s = 170;
	{8'd66,8'd105} : s = 171;
	{8'd66,8'd106} : s = 172;
	{8'd66,8'd107} : s = 173;
	{8'd66,8'd108} : s = 174;
	{8'd66,8'd109} : s = 175;
	{8'd66,8'd110} : s = 176;
	{8'd66,8'd111} : s = 177;
	{8'd66,8'd112} : s = 178;
	{8'd66,8'd113} : s = 179;
	{8'd66,8'd114} : s = 180;
	{8'd66,8'd115} : s = 181;
	{8'd66,8'd116} : s = 182;
	{8'd66,8'd117} : s = 183;
	{8'd66,8'd118} : s = 184;
	{8'd66,8'd119} : s = 185;
	{8'd66,8'd120} : s = 186;
	{8'd66,8'd121} : s = 187;
	{8'd66,8'd122} : s = 188;
	{8'd66,8'd123} : s = 189;
	{8'd66,8'd124} : s = 190;
	{8'd66,8'd125} : s = 191;
	{8'd66,8'd126} : s = 192;
	{8'd66,8'd127} : s = 193;
	{8'd66,8'd128} : s = 194;
	{8'd66,8'd129} : s = 195;
	{8'd66,8'd130} : s = 196;
	{8'd66,8'd131} : s = 197;
	{8'd66,8'd132} : s = 198;
	{8'd66,8'd133} : s = 199;
	{8'd66,8'd134} : s = 200;
	{8'd66,8'd135} : s = 201;
	{8'd66,8'd136} : s = 202;
	{8'd66,8'd137} : s = 203;
	{8'd66,8'd138} : s = 204;
	{8'd66,8'd139} : s = 205;
	{8'd66,8'd140} : s = 206;
	{8'd66,8'd141} : s = 207;
	{8'd66,8'd142} : s = 208;
	{8'd66,8'd143} : s = 209;
	{8'd66,8'd144} : s = 210;
	{8'd66,8'd145} : s = 211;
	{8'd66,8'd146} : s = 212;
	{8'd66,8'd147} : s = 213;
	{8'd66,8'd148} : s = 214;
	{8'd66,8'd149} : s = 215;
	{8'd66,8'd150} : s = 216;
	{8'd66,8'd151} : s = 217;
	{8'd66,8'd152} : s = 218;
	{8'd66,8'd153} : s = 219;
	{8'd66,8'd154} : s = 220;
	{8'd66,8'd155} : s = 221;
	{8'd66,8'd156} : s = 222;
	{8'd66,8'd157} : s = 223;
	{8'd66,8'd158} : s = 224;
	{8'd66,8'd159} : s = 225;
	{8'd66,8'd160} : s = 226;
	{8'd66,8'd161} : s = 227;
	{8'd66,8'd162} : s = 228;
	{8'd66,8'd163} : s = 229;
	{8'd66,8'd164} : s = 230;
	{8'd66,8'd165} : s = 231;
	{8'd66,8'd166} : s = 232;
	{8'd66,8'd167} : s = 233;
	{8'd66,8'd168} : s = 234;
	{8'd66,8'd169} : s = 235;
	{8'd66,8'd170} : s = 236;
	{8'd66,8'd171} : s = 237;
	{8'd66,8'd172} : s = 238;
	{8'd66,8'd173} : s = 239;
	{8'd66,8'd174} : s = 240;
	{8'd66,8'd175} : s = 241;
	{8'd66,8'd176} : s = 242;
	{8'd66,8'd177} : s = 243;
	{8'd66,8'd178} : s = 244;
	{8'd66,8'd179} : s = 245;
	{8'd66,8'd180} : s = 246;
	{8'd66,8'd181} : s = 247;
	{8'd66,8'd182} : s = 248;
	{8'd66,8'd183} : s = 249;
	{8'd66,8'd184} : s = 250;
	{8'd66,8'd185} : s = 251;
	{8'd66,8'd186} : s = 252;
	{8'd66,8'd187} : s = 253;
	{8'd66,8'd188} : s = 254;
	{8'd66,8'd189} : s = 255;
	{8'd66,8'd190} : s = 256;
	{8'd66,8'd191} : s = 257;
	{8'd66,8'd192} : s = 258;
	{8'd66,8'd193} : s = 259;
	{8'd66,8'd194} : s = 260;
	{8'd66,8'd195} : s = 261;
	{8'd66,8'd196} : s = 262;
	{8'd66,8'd197} : s = 263;
	{8'd66,8'd198} : s = 264;
	{8'd66,8'd199} : s = 265;
	{8'd66,8'd200} : s = 266;
	{8'd66,8'd201} : s = 267;
	{8'd66,8'd202} : s = 268;
	{8'd66,8'd203} : s = 269;
	{8'd66,8'd204} : s = 270;
	{8'd66,8'd205} : s = 271;
	{8'd66,8'd206} : s = 272;
	{8'd66,8'd207} : s = 273;
	{8'd66,8'd208} : s = 274;
	{8'd66,8'd209} : s = 275;
	{8'd66,8'd210} : s = 276;
	{8'd66,8'd211} : s = 277;
	{8'd66,8'd212} : s = 278;
	{8'd66,8'd213} : s = 279;
	{8'd66,8'd214} : s = 280;
	{8'd66,8'd215} : s = 281;
	{8'd66,8'd216} : s = 282;
	{8'd66,8'd217} : s = 283;
	{8'd66,8'd218} : s = 284;
	{8'd66,8'd219} : s = 285;
	{8'd66,8'd220} : s = 286;
	{8'd66,8'd221} : s = 287;
	{8'd66,8'd222} : s = 288;
	{8'd66,8'd223} : s = 289;
	{8'd66,8'd224} : s = 290;
	{8'd66,8'd225} : s = 291;
	{8'd66,8'd226} : s = 292;
	{8'd66,8'd227} : s = 293;
	{8'd66,8'd228} : s = 294;
	{8'd66,8'd229} : s = 295;
	{8'd66,8'd230} : s = 296;
	{8'd66,8'd231} : s = 297;
	{8'd66,8'd232} : s = 298;
	{8'd66,8'd233} : s = 299;
	{8'd66,8'd234} : s = 300;
	{8'd66,8'd235} : s = 301;
	{8'd66,8'd236} : s = 302;
	{8'd66,8'd237} : s = 303;
	{8'd66,8'd238} : s = 304;
	{8'd66,8'd239} : s = 305;
	{8'd66,8'd240} : s = 306;
	{8'd66,8'd241} : s = 307;
	{8'd66,8'd242} : s = 308;
	{8'd66,8'd243} : s = 309;
	{8'd66,8'd244} : s = 310;
	{8'd66,8'd245} : s = 311;
	{8'd66,8'd246} : s = 312;
	{8'd66,8'd247} : s = 313;
	{8'd66,8'd248} : s = 314;
	{8'd66,8'd249} : s = 315;
	{8'd66,8'd250} : s = 316;
	{8'd66,8'd251} : s = 317;
	{8'd66,8'd252} : s = 318;
	{8'd66,8'd253} : s = 319;
	{8'd66,8'd254} : s = 320;
	{8'd66,8'd255} : s = 321;
	{8'd67,8'd0} : s = 67;
	{8'd67,8'd1} : s = 68;
	{8'd67,8'd2} : s = 69;
	{8'd67,8'd3} : s = 70;
	{8'd67,8'd4} : s = 71;
	{8'd67,8'd5} : s = 72;
	{8'd67,8'd6} : s = 73;
	{8'd67,8'd7} : s = 74;
	{8'd67,8'd8} : s = 75;
	{8'd67,8'd9} : s = 76;
	{8'd67,8'd10} : s = 77;
	{8'd67,8'd11} : s = 78;
	{8'd67,8'd12} : s = 79;
	{8'd67,8'd13} : s = 80;
	{8'd67,8'd14} : s = 81;
	{8'd67,8'd15} : s = 82;
	{8'd67,8'd16} : s = 83;
	{8'd67,8'd17} : s = 84;
	{8'd67,8'd18} : s = 85;
	{8'd67,8'd19} : s = 86;
	{8'd67,8'd20} : s = 87;
	{8'd67,8'd21} : s = 88;
	{8'd67,8'd22} : s = 89;
	{8'd67,8'd23} : s = 90;
	{8'd67,8'd24} : s = 91;
	{8'd67,8'd25} : s = 92;
	{8'd67,8'd26} : s = 93;
	{8'd67,8'd27} : s = 94;
	{8'd67,8'd28} : s = 95;
	{8'd67,8'd29} : s = 96;
	{8'd67,8'd30} : s = 97;
	{8'd67,8'd31} : s = 98;
	{8'd67,8'd32} : s = 99;
	{8'd67,8'd33} : s = 100;
	{8'd67,8'd34} : s = 101;
	{8'd67,8'd35} : s = 102;
	{8'd67,8'd36} : s = 103;
	{8'd67,8'd37} : s = 104;
	{8'd67,8'd38} : s = 105;
	{8'd67,8'd39} : s = 106;
	{8'd67,8'd40} : s = 107;
	{8'd67,8'd41} : s = 108;
	{8'd67,8'd42} : s = 109;
	{8'd67,8'd43} : s = 110;
	{8'd67,8'd44} : s = 111;
	{8'd67,8'd45} : s = 112;
	{8'd67,8'd46} : s = 113;
	{8'd67,8'd47} : s = 114;
	{8'd67,8'd48} : s = 115;
	{8'd67,8'd49} : s = 116;
	{8'd67,8'd50} : s = 117;
	{8'd67,8'd51} : s = 118;
	{8'd67,8'd52} : s = 119;
	{8'd67,8'd53} : s = 120;
	{8'd67,8'd54} : s = 121;
	{8'd67,8'd55} : s = 122;
	{8'd67,8'd56} : s = 123;
	{8'd67,8'd57} : s = 124;
	{8'd67,8'd58} : s = 125;
	{8'd67,8'd59} : s = 126;
	{8'd67,8'd60} : s = 127;
	{8'd67,8'd61} : s = 128;
	{8'd67,8'd62} : s = 129;
	{8'd67,8'd63} : s = 130;
	{8'd67,8'd64} : s = 131;
	{8'd67,8'd65} : s = 132;
	{8'd67,8'd66} : s = 133;
	{8'd67,8'd67} : s = 134;
	{8'd67,8'd68} : s = 135;
	{8'd67,8'd69} : s = 136;
	{8'd67,8'd70} : s = 137;
	{8'd67,8'd71} : s = 138;
	{8'd67,8'd72} : s = 139;
	{8'd67,8'd73} : s = 140;
	{8'd67,8'd74} : s = 141;
	{8'd67,8'd75} : s = 142;
	{8'd67,8'd76} : s = 143;
	{8'd67,8'd77} : s = 144;
	{8'd67,8'd78} : s = 145;
	{8'd67,8'd79} : s = 146;
	{8'd67,8'd80} : s = 147;
	{8'd67,8'd81} : s = 148;
	{8'd67,8'd82} : s = 149;
	{8'd67,8'd83} : s = 150;
	{8'd67,8'd84} : s = 151;
	{8'd67,8'd85} : s = 152;
	{8'd67,8'd86} : s = 153;
	{8'd67,8'd87} : s = 154;
	{8'd67,8'd88} : s = 155;
	{8'd67,8'd89} : s = 156;
	{8'd67,8'd90} : s = 157;
	{8'd67,8'd91} : s = 158;
	{8'd67,8'd92} : s = 159;
	{8'd67,8'd93} : s = 160;
	{8'd67,8'd94} : s = 161;
	{8'd67,8'd95} : s = 162;
	{8'd67,8'd96} : s = 163;
	{8'd67,8'd97} : s = 164;
	{8'd67,8'd98} : s = 165;
	{8'd67,8'd99} : s = 166;
	{8'd67,8'd100} : s = 167;
	{8'd67,8'd101} : s = 168;
	{8'd67,8'd102} : s = 169;
	{8'd67,8'd103} : s = 170;
	{8'd67,8'd104} : s = 171;
	{8'd67,8'd105} : s = 172;
	{8'd67,8'd106} : s = 173;
	{8'd67,8'd107} : s = 174;
	{8'd67,8'd108} : s = 175;
	{8'd67,8'd109} : s = 176;
	{8'd67,8'd110} : s = 177;
	{8'd67,8'd111} : s = 178;
	{8'd67,8'd112} : s = 179;
	{8'd67,8'd113} : s = 180;
	{8'd67,8'd114} : s = 181;
	{8'd67,8'd115} : s = 182;
	{8'd67,8'd116} : s = 183;
	{8'd67,8'd117} : s = 184;
	{8'd67,8'd118} : s = 185;
	{8'd67,8'd119} : s = 186;
	{8'd67,8'd120} : s = 187;
	{8'd67,8'd121} : s = 188;
	{8'd67,8'd122} : s = 189;
	{8'd67,8'd123} : s = 190;
	{8'd67,8'd124} : s = 191;
	{8'd67,8'd125} : s = 192;
	{8'd67,8'd126} : s = 193;
	{8'd67,8'd127} : s = 194;
	{8'd67,8'd128} : s = 195;
	{8'd67,8'd129} : s = 196;
	{8'd67,8'd130} : s = 197;
	{8'd67,8'd131} : s = 198;
	{8'd67,8'd132} : s = 199;
	{8'd67,8'd133} : s = 200;
	{8'd67,8'd134} : s = 201;
	{8'd67,8'd135} : s = 202;
	{8'd67,8'd136} : s = 203;
	{8'd67,8'd137} : s = 204;
	{8'd67,8'd138} : s = 205;
	{8'd67,8'd139} : s = 206;
	{8'd67,8'd140} : s = 207;
	{8'd67,8'd141} : s = 208;
	{8'd67,8'd142} : s = 209;
	{8'd67,8'd143} : s = 210;
	{8'd67,8'd144} : s = 211;
	{8'd67,8'd145} : s = 212;
	{8'd67,8'd146} : s = 213;
	{8'd67,8'd147} : s = 214;
	{8'd67,8'd148} : s = 215;
	{8'd67,8'd149} : s = 216;
	{8'd67,8'd150} : s = 217;
	{8'd67,8'd151} : s = 218;
	{8'd67,8'd152} : s = 219;
	{8'd67,8'd153} : s = 220;
	{8'd67,8'd154} : s = 221;
	{8'd67,8'd155} : s = 222;
	{8'd67,8'd156} : s = 223;
	{8'd67,8'd157} : s = 224;
	{8'd67,8'd158} : s = 225;
	{8'd67,8'd159} : s = 226;
	{8'd67,8'd160} : s = 227;
	{8'd67,8'd161} : s = 228;
	{8'd67,8'd162} : s = 229;
	{8'd67,8'd163} : s = 230;
	{8'd67,8'd164} : s = 231;
	{8'd67,8'd165} : s = 232;
	{8'd67,8'd166} : s = 233;
	{8'd67,8'd167} : s = 234;
	{8'd67,8'd168} : s = 235;
	{8'd67,8'd169} : s = 236;
	{8'd67,8'd170} : s = 237;
	{8'd67,8'd171} : s = 238;
	{8'd67,8'd172} : s = 239;
	{8'd67,8'd173} : s = 240;
	{8'd67,8'd174} : s = 241;
	{8'd67,8'd175} : s = 242;
	{8'd67,8'd176} : s = 243;
	{8'd67,8'd177} : s = 244;
	{8'd67,8'd178} : s = 245;
	{8'd67,8'd179} : s = 246;
	{8'd67,8'd180} : s = 247;
	{8'd67,8'd181} : s = 248;
	{8'd67,8'd182} : s = 249;
	{8'd67,8'd183} : s = 250;
	{8'd67,8'd184} : s = 251;
	{8'd67,8'd185} : s = 252;
	{8'd67,8'd186} : s = 253;
	{8'd67,8'd187} : s = 254;
	{8'd67,8'd188} : s = 255;
	{8'd67,8'd189} : s = 256;
	{8'd67,8'd190} : s = 257;
	{8'd67,8'd191} : s = 258;
	{8'd67,8'd192} : s = 259;
	{8'd67,8'd193} : s = 260;
	{8'd67,8'd194} : s = 261;
	{8'd67,8'd195} : s = 262;
	{8'd67,8'd196} : s = 263;
	{8'd67,8'd197} : s = 264;
	{8'd67,8'd198} : s = 265;
	{8'd67,8'd199} : s = 266;
	{8'd67,8'd200} : s = 267;
	{8'd67,8'd201} : s = 268;
	{8'd67,8'd202} : s = 269;
	{8'd67,8'd203} : s = 270;
	{8'd67,8'd204} : s = 271;
	{8'd67,8'd205} : s = 272;
	{8'd67,8'd206} : s = 273;
	{8'd67,8'd207} : s = 274;
	{8'd67,8'd208} : s = 275;
	{8'd67,8'd209} : s = 276;
	{8'd67,8'd210} : s = 277;
	{8'd67,8'd211} : s = 278;
	{8'd67,8'd212} : s = 279;
	{8'd67,8'd213} : s = 280;
	{8'd67,8'd214} : s = 281;
	{8'd67,8'd215} : s = 282;
	{8'd67,8'd216} : s = 283;
	{8'd67,8'd217} : s = 284;
	{8'd67,8'd218} : s = 285;
	{8'd67,8'd219} : s = 286;
	{8'd67,8'd220} : s = 287;
	{8'd67,8'd221} : s = 288;
	{8'd67,8'd222} : s = 289;
	{8'd67,8'd223} : s = 290;
	{8'd67,8'd224} : s = 291;
	{8'd67,8'd225} : s = 292;
	{8'd67,8'd226} : s = 293;
	{8'd67,8'd227} : s = 294;
	{8'd67,8'd228} : s = 295;
	{8'd67,8'd229} : s = 296;
	{8'd67,8'd230} : s = 297;
	{8'd67,8'd231} : s = 298;
	{8'd67,8'd232} : s = 299;
	{8'd67,8'd233} : s = 300;
	{8'd67,8'd234} : s = 301;
	{8'd67,8'd235} : s = 302;
	{8'd67,8'd236} : s = 303;
	{8'd67,8'd237} : s = 304;
	{8'd67,8'd238} : s = 305;
	{8'd67,8'd239} : s = 306;
	{8'd67,8'd240} : s = 307;
	{8'd67,8'd241} : s = 308;
	{8'd67,8'd242} : s = 309;
	{8'd67,8'd243} : s = 310;
	{8'd67,8'd244} : s = 311;
	{8'd67,8'd245} : s = 312;
	{8'd67,8'd246} : s = 313;
	{8'd67,8'd247} : s = 314;
	{8'd67,8'd248} : s = 315;
	{8'd67,8'd249} : s = 316;
	{8'd67,8'd250} : s = 317;
	{8'd67,8'd251} : s = 318;
	{8'd67,8'd252} : s = 319;
	{8'd67,8'd253} : s = 320;
	{8'd67,8'd254} : s = 321;
	{8'd67,8'd255} : s = 322;
	{8'd68,8'd0} : s = 68;
	{8'd68,8'd1} : s = 69;
	{8'd68,8'd2} : s = 70;
	{8'd68,8'd3} : s = 71;
	{8'd68,8'd4} : s = 72;
	{8'd68,8'd5} : s = 73;
	{8'd68,8'd6} : s = 74;
	{8'd68,8'd7} : s = 75;
	{8'd68,8'd8} : s = 76;
	{8'd68,8'd9} : s = 77;
	{8'd68,8'd10} : s = 78;
	{8'd68,8'd11} : s = 79;
	{8'd68,8'd12} : s = 80;
	{8'd68,8'd13} : s = 81;
	{8'd68,8'd14} : s = 82;
	{8'd68,8'd15} : s = 83;
	{8'd68,8'd16} : s = 84;
	{8'd68,8'd17} : s = 85;
	{8'd68,8'd18} : s = 86;
	{8'd68,8'd19} : s = 87;
	{8'd68,8'd20} : s = 88;
	{8'd68,8'd21} : s = 89;
	{8'd68,8'd22} : s = 90;
	{8'd68,8'd23} : s = 91;
	{8'd68,8'd24} : s = 92;
	{8'd68,8'd25} : s = 93;
	{8'd68,8'd26} : s = 94;
	{8'd68,8'd27} : s = 95;
	{8'd68,8'd28} : s = 96;
	{8'd68,8'd29} : s = 97;
	{8'd68,8'd30} : s = 98;
	{8'd68,8'd31} : s = 99;
	{8'd68,8'd32} : s = 100;
	{8'd68,8'd33} : s = 101;
	{8'd68,8'd34} : s = 102;
	{8'd68,8'd35} : s = 103;
	{8'd68,8'd36} : s = 104;
	{8'd68,8'd37} : s = 105;
	{8'd68,8'd38} : s = 106;
	{8'd68,8'd39} : s = 107;
	{8'd68,8'd40} : s = 108;
	{8'd68,8'd41} : s = 109;
	{8'd68,8'd42} : s = 110;
	{8'd68,8'd43} : s = 111;
	{8'd68,8'd44} : s = 112;
	{8'd68,8'd45} : s = 113;
	{8'd68,8'd46} : s = 114;
	{8'd68,8'd47} : s = 115;
	{8'd68,8'd48} : s = 116;
	{8'd68,8'd49} : s = 117;
	{8'd68,8'd50} : s = 118;
	{8'd68,8'd51} : s = 119;
	{8'd68,8'd52} : s = 120;
	{8'd68,8'd53} : s = 121;
	{8'd68,8'd54} : s = 122;
	{8'd68,8'd55} : s = 123;
	{8'd68,8'd56} : s = 124;
	{8'd68,8'd57} : s = 125;
	{8'd68,8'd58} : s = 126;
	{8'd68,8'd59} : s = 127;
	{8'd68,8'd60} : s = 128;
	{8'd68,8'd61} : s = 129;
	{8'd68,8'd62} : s = 130;
	{8'd68,8'd63} : s = 131;
	{8'd68,8'd64} : s = 132;
	{8'd68,8'd65} : s = 133;
	{8'd68,8'd66} : s = 134;
	{8'd68,8'd67} : s = 135;
	{8'd68,8'd68} : s = 136;
	{8'd68,8'd69} : s = 137;
	{8'd68,8'd70} : s = 138;
	{8'd68,8'd71} : s = 139;
	{8'd68,8'd72} : s = 140;
	{8'd68,8'd73} : s = 141;
	{8'd68,8'd74} : s = 142;
	{8'd68,8'd75} : s = 143;
	{8'd68,8'd76} : s = 144;
	{8'd68,8'd77} : s = 145;
	{8'd68,8'd78} : s = 146;
	{8'd68,8'd79} : s = 147;
	{8'd68,8'd80} : s = 148;
	{8'd68,8'd81} : s = 149;
	{8'd68,8'd82} : s = 150;
	{8'd68,8'd83} : s = 151;
	{8'd68,8'd84} : s = 152;
	{8'd68,8'd85} : s = 153;
	{8'd68,8'd86} : s = 154;
	{8'd68,8'd87} : s = 155;
	{8'd68,8'd88} : s = 156;
	{8'd68,8'd89} : s = 157;
	{8'd68,8'd90} : s = 158;
	{8'd68,8'd91} : s = 159;
	{8'd68,8'd92} : s = 160;
	{8'd68,8'd93} : s = 161;
	{8'd68,8'd94} : s = 162;
	{8'd68,8'd95} : s = 163;
	{8'd68,8'd96} : s = 164;
	{8'd68,8'd97} : s = 165;
	{8'd68,8'd98} : s = 166;
	{8'd68,8'd99} : s = 167;
	{8'd68,8'd100} : s = 168;
	{8'd68,8'd101} : s = 169;
	{8'd68,8'd102} : s = 170;
	{8'd68,8'd103} : s = 171;
	{8'd68,8'd104} : s = 172;
	{8'd68,8'd105} : s = 173;
	{8'd68,8'd106} : s = 174;
	{8'd68,8'd107} : s = 175;
	{8'd68,8'd108} : s = 176;
	{8'd68,8'd109} : s = 177;
	{8'd68,8'd110} : s = 178;
	{8'd68,8'd111} : s = 179;
	{8'd68,8'd112} : s = 180;
	{8'd68,8'd113} : s = 181;
	{8'd68,8'd114} : s = 182;
	{8'd68,8'd115} : s = 183;
	{8'd68,8'd116} : s = 184;
	{8'd68,8'd117} : s = 185;
	{8'd68,8'd118} : s = 186;
	{8'd68,8'd119} : s = 187;
	{8'd68,8'd120} : s = 188;
	{8'd68,8'd121} : s = 189;
	{8'd68,8'd122} : s = 190;
	{8'd68,8'd123} : s = 191;
	{8'd68,8'd124} : s = 192;
	{8'd68,8'd125} : s = 193;
	{8'd68,8'd126} : s = 194;
	{8'd68,8'd127} : s = 195;
	{8'd68,8'd128} : s = 196;
	{8'd68,8'd129} : s = 197;
	{8'd68,8'd130} : s = 198;
	{8'd68,8'd131} : s = 199;
	{8'd68,8'd132} : s = 200;
	{8'd68,8'd133} : s = 201;
	{8'd68,8'd134} : s = 202;
	{8'd68,8'd135} : s = 203;
	{8'd68,8'd136} : s = 204;
	{8'd68,8'd137} : s = 205;
	{8'd68,8'd138} : s = 206;
	{8'd68,8'd139} : s = 207;
	{8'd68,8'd140} : s = 208;
	{8'd68,8'd141} : s = 209;
	{8'd68,8'd142} : s = 210;
	{8'd68,8'd143} : s = 211;
	{8'd68,8'd144} : s = 212;
	{8'd68,8'd145} : s = 213;
	{8'd68,8'd146} : s = 214;
	{8'd68,8'd147} : s = 215;
	{8'd68,8'd148} : s = 216;
	{8'd68,8'd149} : s = 217;
	{8'd68,8'd150} : s = 218;
	{8'd68,8'd151} : s = 219;
	{8'd68,8'd152} : s = 220;
	{8'd68,8'd153} : s = 221;
	{8'd68,8'd154} : s = 222;
	{8'd68,8'd155} : s = 223;
	{8'd68,8'd156} : s = 224;
	{8'd68,8'd157} : s = 225;
	{8'd68,8'd158} : s = 226;
	{8'd68,8'd159} : s = 227;
	{8'd68,8'd160} : s = 228;
	{8'd68,8'd161} : s = 229;
	{8'd68,8'd162} : s = 230;
	{8'd68,8'd163} : s = 231;
	{8'd68,8'd164} : s = 232;
	{8'd68,8'd165} : s = 233;
	{8'd68,8'd166} : s = 234;
	{8'd68,8'd167} : s = 235;
	{8'd68,8'd168} : s = 236;
	{8'd68,8'd169} : s = 237;
	{8'd68,8'd170} : s = 238;
	{8'd68,8'd171} : s = 239;
	{8'd68,8'd172} : s = 240;
	{8'd68,8'd173} : s = 241;
	{8'd68,8'd174} : s = 242;
	{8'd68,8'd175} : s = 243;
	{8'd68,8'd176} : s = 244;
	{8'd68,8'd177} : s = 245;
	{8'd68,8'd178} : s = 246;
	{8'd68,8'd179} : s = 247;
	{8'd68,8'd180} : s = 248;
	{8'd68,8'd181} : s = 249;
	{8'd68,8'd182} : s = 250;
	{8'd68,8'd183} : s = 251;
	{8'd68,8'd184} : s = 252;
	{8'd68,8'd185} : s = 253;
	{8'd68,8'd186} : s = 254;
	{8'd68,8'd187} : s = 255;
	{8'd68,8'd188} : s = 256;
	{8'd68,8'd189} : s = 257;
	{8'd68,8'd190} : s = 258;
	{8'd68,8'd191} : s = 259;
	{8'd68,8'd192} : s = 260;
	{8'd68,8'd193} : s = 261;
	{8'd68,8'd194} : s = 262;
	{8'd68,8'd195} : s = 263;
	{8'd68,8'd196} : s = 264;
	{8'd68,8'd197} : s = 265;
	{8'd68,8'd198} : s = 266;
	{8'd68,8'd199} : s = 267;
	{8'd68,8'd200} : s = 268;
	{8'd68,8'd201} : s = 269;
	{8'd68,8'd202} : s = 270;
	{8'd68,8'd203} : s = 271;
	{8'd68,8'd204} : s = 272;
	{8'd68,8'd205} : s = 273;
	{8'd68,8'd206} : s = 274;
	{8'd68,8'd207} : s = 275;
	{8'd68,8'd208} : s = 276;
	{8'd68,8'd209} : s = 277;
	{8'd68,8'd210} : s = 278;
	{8'd68,8'd211} : s = 279;
	{8'd68,8'd212} : s = 280;
	{8'd68,8'd213} : s = 281;
	{8'd68,8'd214} : s = 282;
	{8'd68,8'd215} : s = 283;
	{8'd68,8'd216} : s = 284;
	{8'd68,8'd217} : s = 285;
	{8'd68,8'd218} : s = 286;
	{8'd68,8'd219} : s = 287;
	{8'd68,8'd220} : s = 288;
	{8'd68,8'd221} : s = 289;
	{8'd68,8'd222} : s = 290;
	{8'd68,8'd223} : s = 291;
	{8'd68,8'd224} : s = 292;
	{8'd68,8'd225} : s = 293;
	{8'd68,8'd226} : s = 294;
	{8'd68,8'd227} : s = 295;
	{8'd68,8'd228} : s = 296;
	{8'd68,8'd229} : s = 297;
	{8'd68,8'd230} : s = 298;
	{8'd68,8'd231} : s = 299;
	{8'd68,8'd232} : s = 300;
	{8'd68,8'd233} : s = 301;
	{8'd68,8'd234} : s = 302;
	{8'd68,8'd235} : s = 303;
	{8'd68,8'd236} : s = 304;
	{8'd68,8'd237} : s = 305;
	{8'd68,8'd238} : s = 306;
	{8'd68,8'd239} : s = 307;
	{8'd68,8'd240} : s = 308;
	{8'd68,8'd241} : s = 309;
	{8'd68,8'd242} : s = 310;
	{8'd68,8'd243} : s = 311;
	{8'd68,8'd244} : s = 312;
	{8'd68,8'd245} : s = 313;
	{8'd68,8'd246} : s = 314;
	{8'd68,8'd247} : s = 315;
	{8'd68,8'd248} : s = 316;
	{8'd68,8'd249} : s = 317;
	{8'd68,8'd250} : s = 318;
	{8'd68,8'd251} : s = 319;
	{8'd68,8'd252} : s = 320;
	{8'd68,8'd253} : s = 321;
	{8'd68,8'd254} : s = 322;
	{8'd68,8'd255} : s = 323;
	{8'd69,8'd0} : s = 69;
	{8'd69,8'd1} : s = 70;
	{8'd69,8'd2} : s = 71;
	{8'd69,8'd3} : s = 72;
	{8'd69,8'd4} : s = 73;
	{8'd69,8'd5} : s = 74;
	{8'd69,8'd6} : s = 75;
	{8'd69,8'd7} : s = 76;
	{8'd69,8'd8} : s = 77;
	{8'd69,8'd9} : s = 78;
	{8'd69,8'd10} : s = 79;
	{8'd69,8'd11} : s = 80;
	{8'd69,8'd12} : s = 81;
	{8'd69,8'd13} : s = 82;
	{8'd69,8'd14} : s = 83;
	{8'd69,8'd15} : s = 84;
	{8'd69,8'd16} : s = 85;
	{8'd69,8'd17} : s = 86;
	{8'd69,8'd18} : s = 87;
	{8'd69,8'd19} : s = 88;
	{8'd69,8'd20} : s = 89;
	{8'd69,8'd21} : s = 90;
	{8'd69,8'd22} : s = 91;
	{8'd69,8'd23} : s = 92;
	{8'd69,8'd24} : s = 93;
	{8'd69,8'd25} : s = 94;
	{8'd69,8'd26} : s = 95;
	{8'd69,8'd27} : s = 96;
	{8'd69,8'd28} : s = 97;
	{8'd69,8'd29} : s = 98;
	{8'd69,8'd30} : s = 99;
	{8'd69,8'd31} : s = 100;
	{8'd69,8'd32} : s = 101;
	{8'd69,8'd33} : s = 102;
	{8'd69,8'd34} : s = 103;
	{8'd69,8'd35} : s = 104;
	{8'd69,8'd36} : s = 105;
	{8'd69,8'd37} : s = 106;
	{8'd69,8'd38} : s = 107;
	{8'd69,8'd39} : s = 108;
	{8'd69,8'd40} : s = 109;
	{8'd69,8'd41} : s = 110;
	{8'd69,8'd42} : s = 111;
	{8'd69,8'd43} : s = 112;
	{8'd69,8'd44} : s = 113;
	{8'd69,8'd45} : s = 114;
	{8'd69,8'd46} : s = 115;
	{8'd69,8'd47} : s = 116;
	{8'd69,8'd48} : s = 117;
	{8'd69,8'd49} : s = 118;
	{8'd69,8'd50} : s = 119;
	{8'd69,8'd51} : s = 120;
	{8'd69,8'd52} : s = 121;
	{8'd69,8'd53} : s = 122;
	{8'd69,8'd54} : s = 123;
	{8'd69,8'd55} : s = 124;
	{8'd69,8'd56} : s = 125;
	{8'd69,8'd57} : s = 126;
	{8'd69,8'd58} : s = 127;
	{8'd69,8'd59} : s = 128;
	{8'd69,8'd60} : s = 129;
	{8'd69,8'd61} : s = 130;
	{8'd69,8'd62} : s = 131;
	{8'd69,8'd63} : s = 132;
	{8'd69,8'd64} : s = 133;
	{8'd69,8'd65} : s = 134;
	{8'd69,8'd66} : s = 135;
	{8'd69,8'd67} : s = 136;
	{8'd69,8'd68} : s = 137;
	{8'd69,8'd69} : s = 138;
	{8'd69,8'd70} : s = 139;
	{8'd69,8'd71} : s = 140;
	{8'd69,8'd72} : s = 141;
	{8'd69,8'd73} : s = 142;
	{8'd69,8'd74} : s = 143;
	{8'd69,8'd75} : s = 144;
	{8'd69,8'd76} : s = 145;
	{8'd69,8'd77} : s = 146;
	{8'd69,8'd78} : s = 147;
	{8'd69,8'd79} : s = 148;
	{8'd69,8'd80} : s = 149;
	{8'd69,8'd81} : s = 150;
	{8'd69,8'd82} : s = 151;
	{8'd69,8'd83} : s = 152;
	{8'd69,8'd84} : s = 153;
	{8'd69,8'd85} : s = 154;
	{8'd69,8'd86} : s = 155;
	{8'd69,8'd87} : s = 156;
	{8'd69,8'd88} : s = 157;
	{8'd69,8'd89} : s = 158;
	{8'd69,8'd90} : s = 159;
	{8'd69,8'd91} : s = 160;
	{8'd69,8'd92} : s = 161;
	{8'd69,8'd93} : s = 162;
	{8'd69,8'd94} : s = 163;
	{8'd69,8'd95} : s = 164;
	{8'd69,8'd96} : s = 165;
	{8'd69,8'd97} : s = 166;
	{8'd69,8'd98} : s = 167;
	{8'd69,8'd99} : s = 168;
	{8'd69,8'd100} : s = 169;
	{8'd69,8'd101} : s = 170;
	{8'd69,8'd102} : s = 171;
	{8'd69,8'd103} : s = 172;
	{8'd69,8'd104} : s = 173;
	{8'd69,8'd105} : s = 174;
	{8'd69,8'd106} : s = 175;
	{8'd69,8'd107} : s = 176;
	{8'd69,8'd108} : s = 177;
	{8'd69,8'd109} : s = 178;
	{8'd69,8'd110} : s = 179;
	{8'd69,8'd111} : s = 180;
	{8'd69,8'd112} : s = 181;
	{8'd69,8'd113} : s = 182;
	{8'd69,8'd114} : s = 183;
	{8'd69,8'd115} : s = 184;
	{8'd69,8'd116} : s = 185;
	{8'd69,8'd117} : s = 186;
	{8'd69,8'd118} : s = 187;
	{8'd69,8'd119} : s = 188;
	{8'd69,8'd120} : s = 189;
	{8'd69,8'd121} : s = 190;
	{8'd69,8'd122} : s = 191;
	{8'd69,8'd123} : s = 192;
	{8'd69,8'd124} : s = 193;
	{8'd69,8'd125} : s = 194;
	{8'd69,8'd126} : s = 195;
	{8'd69,8'd127} : s = 196;
	{8'd69,8'd128} : s = 197;
	{8'd69,8'd129} : s = 198;
	{8'd69,8'd130} : s = 199;
	{8'd69,8'd131} : s = 200;
	{8'd69,8'd132} : s = 201;
	{8'd69,8'd133} : s = 202;
	{8'd69,8'd134} : s = 203;
	{8'd69,8'd135} : s = 204;
	{8'd69,8'd136} : s = 205;
	{8'd69,8'd137} : s = 206;
	{8'd69,8'd138} : s = 207;
	{8'd69,8'd139} : s = 208;
	{8'd69,8'd140} : s = 209;
	{8'd69,8'd141} : s = 210;
	{8'd69,8'd142} : s = 211;
	{8'd69,8'd143} : s = 212;
	{8'd69,8'd144} : s = 213;
	{8'd69,8'd145} : s = 214;
	{8'd69,8'd146} : s = 215;
	{8'd69,8'd147} : s = 216;
	{8'd69,8'd148} : s = 217;
	{8'd69,8'd149} : s = 218;
	{8'd69,8'd150} : s = 219;
	{8'd69,8'd151} : s = 220;
	{8'd69,8'd152} : s = 221;
	{8'd69,8'd153} : s = 222;
	{8'd69,8'd154} : s = 223;
	{8'd69,8'd155} : s = 224;
	{8'd69,8'd156} : s = 225;
	{8'd69,8'd157} : s = 226;
	{8'd69,8'd158} : s = 227;
	{8'd69,8'd159} : s = 228;
	{8'd69,8'd160} : s = 229;
	{8'd69,8'd161} : s = 230;
	{8'd69,8'd162} : s = 231;
	{8'd69,8'd163} : s = 232;
	{8'd69,8'd164} : s = 233;
	{8'd69,8'd165} : s = 234;
	{8'd69,8'd166} : s = 235;
	{8'd69,8'd167} : s = 236;
	{8'd69,8'd168} : s = 237;
	{8'd69,8'd169} : s = 238;
	{8'd69,8'd170} : s = 239;
	{8'd69,8'd171} : s = 240;
	{8'd69,8'd172} : s = 241;
	{8'd69,8'd173} : s = 242;
	{8'd69,8'd174} : s = 243;
	{8'd69,8'd175} : s = 244;
	{8'd69,8'd176} : s = 245;
	{8'd69,8'd177} : s = 246;
	{8'd69,8'd178} : s = 247;
	{8'd69,8'd179} : s = 248;
	{8'd69,8'd180} : s = 249;
	{8'd69,8'd181} : s = 250;
	{8'd69,8'd182} : s = 251;
	{8'd69,8'd183} : s = 252;
	{8'd69,8'd184} : s = 253;
	{8'd69,8'd185} : s = 254;
	{8'd69,8'd186} : s = 255;
	{8'd69,8'd187} : s = 256;
	{8'd69,8'd188} : s = 257;
	{8'd69,8'd189} : s = 258;
	{8'd69,8'd190} : s = 259;
	{8'd69,8'd191} : s = 260;
	{8'd69,8'd192} : s = 261;
	{8'd69,8'd193} : s = 262;
	{8'd69,8'd194} : s = 263;
	{8'd69,8'd195} : s = 264;
	{8'd69,8'd196} : s = 265;
	{8'd69,8'd197} : s = 266;
	{8'd69,8'd198} : s = 267;
	{8'd69,8'd199} : s = 268;
	{8'd69,8'd200} : s = 269;
	{8'd69,8'd201} : s = 270;
	{8'd69,8'd202} : s = 271;
	{8'd69,8'd203} : s = 272;
	{8'd69,8'd204} : s = 273;
	{8'd69,8'd205} : s = 274;
	{8'd69,8'd206} : s = 275;
	{8'd69,8'd207} : s = 276;
	{8'd69,8'd208} : s = 277;
	{8'd69,8'd209} : s = 278;
	{8'd69,8'd210} : s = 279;
	{8'd69,8'd211} : s = 280;
	{8'd69,8'd212} : s = 281;
	{8'd69,8'd213} : s = 282;
	{8'd69,8'd214} : s = 283;
	{8'd69,8'd215} : s = 284;
	{8'd69,8'd216} : s = 285;
	{8'd69,8'd217} : s = 286;
	{8'd69,8'd218} : s = 287;
	{8'd69,8'd219} : s = 288;
	{8'd69,8'd220} : s = 289;
	{8'd69,8'd221} : s = 290;
	{8'd69,8'd222} : s = 291;
	{8'd69,8'd223} : s = 292;
	{8'd69,8'd224} : s = 293;
	{8'd69,8'd225} : s = 294;
	{8'd69,8'd226} : s = 295;
	{8'd69,8'd227} : s = 296;
	{8'd69,8'd228} : s = 297;
	{8'd69,8'd229} : s = 298;
	{8'd69,8'd230} : s = 299;
	{8'd69,8'd231} : s = 300;
	{8'd69,8'd232} : s = 301;
	{8'd69,8'd233} : s = 302;
	{8'd69,8'd234} : s = 303;
	{8'd69,8'd235} : s = 304;
	{8'd69,8'd236} : s = 305;
	{8'd69,8'd237} : s = 306;
	{8'd69,8'd238} : s = 307;
	{8'd69,8'd239} : s = 308;
	{8'd69,8'd240} : s = 309;
	{8'd69,8'd241} : s = 310;
	{8'd69,8'd242} : s = 311;
	{8'd69,8'd243} : s = 312;
	{8'd69,8'd244} : s = 313;
	{8'd69,8'd245} : s = 314;
	{8'd69,8'd246} : s = 315;
	{8'd69,8'd247} : s = 316;
	{8'd69,8'd248} : s = 317;
	{8'd69,8'd249} : s = 318;
	{8'd69,8'd250} : s = 319;
	{8'd69,8'd251} : s = 320;
	{8'd69,8'd252} : s = 321;
	{8'd69,8'd253} : s = 322;
	{8'd69,8'd254} : s = 323;
	{8'd69,8'd255} : s = 324;
	{8'd70,8'd0} : s = 70;
	{8'd70,8'd1} : s = 71;
	{8'd70,8'd2} : s = 72;
	{8'd70,8'd3} : s = 73;
	{8'd70,8'd4} : s = 74;
	{8'd70,8'd5} : s = 75;
	{8'd70,8'd6} : s = 76;
	{8'd70,8'd7} : s = 77;
	{8'd70,8'd8} : s = 78;
	{8'd70,8'd9} : s = 79;
	{8'd70,8'd10} : s = 80;
	{8'd70,8'd11} : s = 81;
	{8'd70,8'd12} : s = 82;
	{8'd70,8'd13} : s = 83;
	{8'd70,8'd14} : s = 84;
	{8'd70,8'd15} : s = 85;
	{8'd70,8'd16} : s = 86;
	{8'd70,8'd17} : s = 87;
	{8'd70,8'd18} : s = 88;
	{8'd70,8'd19} : s = 89;
	{8'd70,8'd20} : s = 90;
	{8'd70,8'd21} : s = 91;
	{8'd70,8'd22} : s = 92;
	{8'd70,8'd23} : s = 93;
	{8'd70,8'd24} : s = 94;
	{8'd70,8'd25} : s = 95;
	{8'd70,8'd26} : s = 96;
	{8'd70,8'd27} : s = 97;
	{8'd70,8'd28} : s = 98;
	{8'd70,8'd29} : s = 99;
	{8'd70,8'd30} : s = 100;
	{8'd70,8'd31} : s = 101;
	{8'd70,8'd32} : s = 102;
	{8'd70,8'd33} : s = 103;
	{8'd70,8'd34} : s = 104;
	{8'd70,8'd35} : s = 105;
	{8'd70,8'd36} : s = 106;
	{8'd70,8'd37} : s = 107;
	{8'd70,8'd38} : s = 108;
	{8'd70,8'd39} : s = 109;
	{8'd70,8'd40} : s = 110;
	{8'd70,8'd41} : s = 111;
	{8'd70,8'd42} : s = 112;
	{8'd70,8'd43} : s = 113;
	{8'd70,8'd44} : s = 114;
	{8'd70,8'd45} : s = 115;
	{8'd70,8'd46} : s = 116;
	{8'd70,8'd47} : s = 117;
	{8'd70,8'd48} : s = 118;
	{8'd70,8'd49} : s = 119;
	{8'd70,8'd50} : s = 120;
	{8'd70,8'd51} : s = 121;
	{8'd70,8'd52} : s = 122;
	{8'd70,8'd53} : s = 123;
	{8'd70,8'd54} : s = 124;
	{8'd70,8'd55} : s = 125;
	{8'd70,8'd56} : s = 126;
	{8'd70,8'd57} : s = 127;
	{8'd70,8'd58} : s = 128;
	{8'd70,8'd59} : s = 129;
	{8'd70,8'd60} : s = 130;
	{8'd70,8'd61} : s = 131;
	{8'd70,8'd62} : s = 132;
	{8'd70,8'd63} : s = 133;
	{8'd70,8'd64} : s = 134;
	{8'd70,8'd65} : s = 135;
	{8'd70,8'd66} : s = 136;
	{8'd70,8'd67} : s = 137;
	{8'd70,8'd68} : s = 138;
	{8'd70,8'd69} : s = 139;
	{8'd70,8'd70} : s = 140;
	{8'd70,8'd71} : s = 141;
	{8'd70,8'd72} : s = 142;
	{8'd70,8'd73} : s = 143;
	{8'd70,8'd74} : s = 144;
	{8'd70,8'd75} : s = 145;
	{8'd70,8'd76} : s = 146;
	{8'd70,8'd77} : s = 147;
	{8'd70,8'd78} : s = 148;
	{8'd70,8'd79} : s = 149;
	{8'd70,8'd80} : s = 150;
	{8'd70,8'd81} : s = 151;
	{8'd70,8'd82} : s = 152;
	{8'd70,8'd83} : s = 153;
	{8'd70,8'd84} : s = 154;
	{8'd70,8'd85} : s = 155;
	{8'd70,8'd86} : s = 156;
	{8'd70,8'd87} : s = 157;
	{8'd70,8'd88} : s = 158;
	{8'd70,8'd89} : s = 159;
	{8'd70,8'd90} : s = 160;
	{8'd70,8'd91} : s = 161;
	{8'd70,8'd92} : s = 162;
	{8'd70,8'd93} : s = 163;
	{8'd70,8'd94} : s = 164;
	{8'd70,8'd95} : s = 165;
	{8'd70,8'd96} : s = 166;
	{8'd70,8'd97} : s = 167;
	{8'd70,8'd98} : s = 168;
	{8'd70,8'd99} : s = 169;
	{8'd70,8'd100} : s = 170;
	{8'd70,8'd101} : s = 171;
	{8'd70,8'd102} : s = 172;
	{8'd70,8'd103} : s = 173;
	{8'd70,8'd104} : s = 174;
	{8'd70,8'd105} : s = 175;
	{8'd70,8'd106} : s = 176;
	{8'd70,8'd107} : s = 177;
	{8'd70,8'd108} : s = 178;
	{8'd70,8'd109} : s = 179;
	{8'd70,8'd110} : s = 180;
	{8'd70,8'd111} : s = 181;
	{8'd70,8'd112} : s = 182;
	{8'd70,8'd113} : s = 183;
	{8'd70,8'd114} : s = 184;
	{8'd70,8'd115} : s = 185;
	{8'd70,8'd116} : s = 186;
	{8'd70,8'd117} : s = 187;
	{8'd70,8'd118} : s = 188;
	{8'd70,8'd119} : s = 189;
	{8'd70,8'd120} : s = 190;
	{8'd70,8'd121} : s = 191;
	{8'd70,8'd122} : s = 192;
	{8'd70,8'd123} : s = 193;
	{8'd70,8'd124} : s = 194;
	{8'd70,8'd125} : s = 195;
	{8'd70,8'd126} : s = 196;
	{8'd70,8'd127} : s = 197;
	{8'd70,8'd128} : s = 198;
	{8'd70,8'd129} : s = 199;
	{8'd70,8'd130} : s = 200;
	{8'd70,8'd131} : s = 201;
	{8'd70,8'd132} : s = 202;
	{8'd70,8'd133} : s = 203;
	{8'd70,8'd134} : s = 204;
	{8'd70,8'd135} : s = 205;
	{8'd70,8'd136} : s = 206;
	{8'd70,8'd137} : s = 207;
	{8'd70,8'd138} : s = 208;
	{8'd70,8'd139} : s = 209;
	{8'd70,8'd140} : s = 210;
	{8'd70,8'd141} : s = 211;
	{8'd70,8'd142} : s = 212;
	{8'd70,8'd143} : s = 213;
	{8'd70,8'd144} : s = 214;
	{8'd70,8'd145} : s = 215;
	{8'd70,8'd146} : s = 216;
	{8'd70,8'd147} : s = 217;
	{8'd70,8'd148} : s = 218;
	{8'd70,8'd149} : s = 219;
	{8'd70,8'd150} : s = 220;
	{8'd70,8'd151} : s = 221;
	{8'd70,8'd152} : s = 222;
	{8'd70,8'd153} : s = 223;
	{8'd70,8'd154} : s = 224;
	{8'd70,8'd155} : s = 225;
	{8'd70,8'd156} : s = 226;
	{8'd70,8'd157} : s = 227;
	{8'd70,8'd158} : s = 228;
	{8'd70,8'd159} : s = 229;
	{8'd70,8'd160} : s = 230;
	{8'd70,8'd161} : s = 231;
	{8'd70,8'd162} : s = 232;
	{8'd70,8'd163} : s = 233;
	{8'd70,8'd164} : s = 234;
	{8'd70,8'd165} : s = 235;
	{8'd70,8'd166} : s = 236;
	{8'd70,8'd167} : s = 237;
	{8'd70,8'd168} : s = 238;
	{8'd70,8'd169} : s = 239;
	{8'd70,8'd170} : s = 240;
	{8'd70,8'd171} : s = 241;
	{8'd70,8'd172} : s = 242;
	{8'd70,8'd173} : s = 243;
	{8'd70,8'd174} : s = 244;
	{8'd70,8'd175} : s = 245;
	{8'd70,8'd176} : s = 246;
	{8'd70,8'd177} : s = 247;
	{8'd70,8'd178} : s = 248;
	{8'd70,8'd179} : s = 249;
	{8'd70,8'd180} : s = 250;
	{8'd70,8'd181} : s = 251;
	{8'd70,8'd182} : s = 252;
	{8'd70,8'd183} : s = 253;
	{8'd70,8'd184} : s = 254;
	{8'd70,8'd185} : s = 255;
	{8'd70,8'd186} : s = 256;
	{8'd70,8'd187} : s = 257;
	{8'd70,8'd188} : s = 258;
	{8'd70,8'd189} : s = 259;
	{8'd70,8'd190} : s = 260;
	{8'd70,8'd191} : s = 261;
	{8'd70,8'd192} : s = 262;
	{8'd70,8'd193} : s = 263;
	{8'd70,8'd194} : s = 264;
	{8'd70,8'd195} : s = 265;
	{8'd70,8'd196} : s = 266;
	{8'd70,8'd197} : s = 267;
	{8'd70,8'd198} : s = 268;
	{8'd70,8'd199} : s = 269;
	{8'd70,8'd200} : s = 270;
	{8'd70,8'd201} : s = 271;
	{8'd70,8'd202} : s = 272;
	{8'd70,8'd203} : s = 273;
	{8'd70,8'd204} : s = 274;
	{8'd70,8'd205} : s = 275;
	{8'd70,8'd206} : s = 276;
	{8'd70,8'd207} : s = 277;
	{8'd70,8'd208} : s = 278;
	{8'd70,8'd209} : s = 279;
	{8'd70,8'd210} : s = 280;
	{8'd70,8'd211} : s = 281;
	{8'd70,8'd212} : s = 282;
	{8'd70,8'd213} : s = 283;
	{8'd70,8'd214} : s = 284;
	{8'd70,8'd215} : s = 285;
	{8'd70,8'd216} : s = 286;
	{8'd70,8'd217} : s = 287;
	{8'd70,8'd218} : s = 288;
	{8'd70,8'd219} : s = 289;
	{8'd70,8'd220} : s = 290;
	{8'd70,8'd221} : s = 291;
	{8'd70,8'd222} : s = 292;
	{8'd70,8'd223} : s = 293;
	{8'd70,8'd224} : s = 294;
	{8'd70,8'd225} : s = 295;
	{8'd70,8'd226} : s = 296;
	{8'd70,8'd227} : s = 297;
	{8'd70,8'd228} : s = 298;
	{8'd70,8'd229} : s = 299;
	{8'd70,8'd230} : s = 300;
	{8'd70,8'd231} : s = 301;
	{8'd70,8'd232} : s = 302;
	{8'd70,8'd233} : s = 303;
	{8'd70,8'd234} : s = 304;
	{8'd70,8'd235} : s = 305;
	{8'd70,8'd236} : s = 306;
	{8'd70,8'd237} : s = 307;
	{8'd70,8'd238} : s = 308;
	{8'd70,8'd239} : s = 309;
	{8'd70,8'd240} : s = 310;
	{8'd70,8'd241} : s = 311;
	{8'd70,8'd242} : s = 312;
	{8'd70,8'd243} : s = 313;
	{8'd70,8'd244} : s = 314;
	{8'd70,8'd245} : s = 315;
	{8'd70,8'd246} : s = 316;
	{8'd70,8'd247} : s = 317;
	{8'd70,8'd248} : s = 318;
	{8'd70,8'd249} : s = 319;
	{8'd70,8'd250} : s = 320;
	{8'd70,8'd251} : s = 321;
	{8'd70,8'd252} : s = 322;
	{8'd70,8'd253} : s = 323;
	{8'd70,8'd254} : s = 324;
	{8'd70,8'd255} : s = 325;
	{8'd71,8'd0} : s = 71;
	{8'd71,8'd1} : s = 72;
	{8'd71,8'd2} : s = 73;
	{8'd71,8'd3} : s = 74;
	{8'd71,8'd4} : s = 75;
	{8'd71,8'd5} : s = 76;
	{8'd71,8'd6} : s = 77;
	{8'd71,8'd7} : s = 78;
	{8'd71,8'd8} : s = 79;
	{8'd71,8'd9} : s = 80;
	{8'd71,8'd10} : s = 81;
	{8'd71,8'd11} : s = 82;
	{8'd71,8'd12} : s = 83;
	{8'd71,8'd13} : s = 84;
	{8'd71,8'd14} : s = 85;
	{8'd71,8'd15} : s = 86;
	{8'd71,8'd16} : s = 87;
	{8'd71,8'd17} : s = 88;
	{8'd71,8'd18} : s = 89;
	{8'd71,8'd19} : s = 90;
	{8'd71,8'd20} : s = 91;
	{8'd71,8'd21} : s = 92;
	{8'd71,8'd22} : s = 93;
	{8'd71,8'd23} : s = 94;
	{8'd71,8'd24} : s = 95;
	{8'd71,8'd25} : s = 96;
	{8'd71,8'd26} : s = 97;
	{8'd71,8'd27} : s = 98;
	{8'd71,8'd28} : s = 99;
	{8'd71,8'd29} : s = 100;
	{8'd71,8'd30} : s = 101;
	{8'd71,8'd31} : s = 102;
	{8'd71,8'd32} : s = 103;
	{8'd71,8'd33} : s = 104;
	{8'd71,8'd34} : s = 105;
	{8'd71,8'd35} : s = 106;
	{8'd71,8'd36} : s = 107;
	{8'd71,8'd37} : s = 108;
	{8'd71,8'd38} : s = 109;
	{8'd71,8'd39} : s = 110;
	{8'd71,8'd40} : s = 111;
	{8'd71,8'd41} : s = 112;
	{8'd71,8'd42} : s = 113;
	{8'd71,8'd43} : s = 114;
	{8'd71,8'd44} : s = 115;
	{8'd71,8'd45} : s = 116;
	{8'd71,8'd46} : s = 117;
	{8'd71,8'd47} : s = 118;
	{8'd71,8'd48} : s = 119;
	{8'd71,8'd49} : s = 120;
	{8'd71,8'd50} : s = 121;
	{8'd71,8'd51} : s = 122;
	{8'd71,8'd52} : s = 123;
	{8'd71,8'd53} : s = 124;
	{8'd71,8'd54} : s = 125;
	{8'd71,8'd55} : s = 126;
	{8'd71,8'd56} : s = 127;
	{8'd71,8'd57} : s = 128;
	{8'd71,8'd58} : s = 129;
	{8'd71,8'd59} : s = 130;
	{8'd71,8'd60} : s = 131;
	{8'd71,8'd61} : s = 132;
	{8'd71,8'd62} : s = 133;
	{8'd71,8'd63} : s = 134;
	{8'd71,8'd64} : s = 135;
	{8'd71,8'd65} : s = 136;
	{8'd71,8'd66} : s = 137;
	{8'd71,8'd67} : s = 138;
	{8'd71,8'd68} : s = 139;
	{8'd71,8'd69} : s = 140;
	{8'd71,8'd70} : s = 141;
	{8'd71,8'd71} : s = 142;
	{8'd71,8'd72} : s = 143;
	{8'd71,8'd73} : s = 144;
	{8'd71,8'd74} : s = 145;
	{8'd71,8'd75} : s = 146;
	{8'd71,8'd76} : s = 147;
	{8'd71,8'd77} : s = 148;
	{8'd71,8'd78} : s = 149;
	{8'd71,8'd79} : s = 150;
	{8'd71,8'd80} : s = 151;
	{8'd71,8'd81} : s = 152;
	{8'd71,8'd82} : s = 153;
	{8'd71,8'd83} : s = 154;
	{8'd71,8'd84} : s = 155;
	{8'd71,8'd85} : s = 156;
	{8'd71,8'd86} : s = 157;
	{8'd71,8'd87} : s = 158;
	{8'd71,8'd88} : s = 159;
	{8'd71,8'd89} : s = 160;
	{8'd71,8'd90} : s = 161;
	{8'd71,8'd91} : s = 162;
	{8'd71,8'd92} : s = 163;
	{8'd71,8'd93} : s = 164;
	{8'd71,8'd94} : s = 165;
	{8'd71,8'd95} : s = 166;
	{8'd71,8'd96} : s = 167;
	{8'd71,8'd97} : s = 168;
	{8'd71,8'd98} : s = 169;
	{8'd71,8'd99} : s = 170;
	{8'd71,8'd100} : s = 171;
	{8'd71,8'd101} : s = 172;
	{8'd71,8'd102} : s = 173;
	{8'd71,8'd103} : s = 174;
	{8'd71,8'd104} : s = 175;
	{8'd71,8'd105} : s = 176;
	{8'd71,8'd106} : s = 177;
	{8'd71,8'd107} : s = 178;
	{8'd71,8'd108} : s = 179;
	{8'd71,8'd109} : s = 180;
	{8'd71,8'd110} : s = 181;
	{8'd71,8'd111} : s = 182;
	{8'd71,8'd112} : s = 183;
	{8'd71,8'd113} : s = 184;
	{8'd71,8'd114} : s = 185;
	{8'd71,8'd115} : s = 186;
	{8'd71,8'd116} : s = 187;
	{8'd71,8'd117} : s = 188;
	{8'd71,8'd118} : s = 189;
	{8'd71,8'd119} : s = 190;
	{8'd71,8'd120} : s = 191;
	{8'd71,8'd121} : s = 192;
	{8'd71,8'd122} : s = 193;
	{8'd71,8'd123} : s = 194;
	{8'd71,8'd124} : s = 195;
	{8'd71,8'd125} : s = 196;
	{8'd71,8'd126} : s = 197;
	{8'd71,8'd127} : s = 198;
	{8'd71,8'd128} : s = 199;
	{8'd71,8'd129} : s = 200;
	{8'd71,8'd130} : s = 201;
	{8'd71,8'd131} : s = 202;
	{8'd71,8'd132} : s = 203;
	{8'd71,8'd133} : s = 204;
	{8'd71,8'd134} : s = 205;
	{8'd71,8'd135} : s = 206;
	{8'd71,8'd136} : s = 207;
	{8'd71,8'd137} : s = 208;
	{8'd71,8'd138} : s = 209;
	{8'd71,8'd139} : s = 210;
	{8'd71,8'd140} : s = 211;
	{8'd71,8'd141} : s = 212;
	{8'd71,8'd142} : s = 213;
	{8'd71,8'd143} : s = 214;
	{8'd71,8'd144} : s = 215;
	{8'd71,8'd145} : s = 216;
	{8'd71,8'd146} : s = 217;
	{8'd71,8'd147} : s = 218;
	{8'd71,8'd148} : s = 219;
	{8'd71,8'd149} : s = 220;
	{8'd71,8'd150} : s = 221;
	{8'd71,8'd151} : s = 222;
	{8'd71,8'd152} : s = 223;
	{8'd71,8'd153} : s = 224;
	{8'd71,8'd154} : s = 225;
	{8'd71,8'd155} : s = 226;
	{8'd71,8'd156} : s = 227;
	{8'd71,8'd157} : s = 228;
	{8'd71,8'd158} : s = 229;
	{8'd71,8'd159} : s = 230;
	{8'd71,8'd160} : s = 231;
	{8'd71,8'd161} : s = 232;
	{8'd71,8'd162} : s = 233;
	{8'd71,8'd163} : s = 234;
	{8'd71,8'd164} : s = 235;
	{8'd71,8'd165} : s = 236;
	{8'd71,8'd166} : s = 237;
	{8'd71,8'd167} : s = 238;
	{8'd71,8'd168} : s = 239;
	{8'd71,8'd169} : s = 240;
	{8'd71,8'd170} : s = 241;
	{8'd71,8'd171} : s = 242;
	{8'd71,8'd172} : s = 243;
	{8'd71,8'd173} : s = 244;
	{8'd71,8'd174} : s = 245;
	{8'd71,8'd175} : s = 246;
	{8'd71,8'd176} : s = 247;
	{8'd71,8'd177} : s = 248;
	{8'd71,8'd178} : s = 249;
	{8'd71,8'd179} : s = 250;
	{8'd71,8'd180} : s = 251;
	{8'd71,8'd181} : s = 252;
	{8'd71,8'd182} : s = 253;
	{8'd71,8'd183} : s = 254;
	{8'd71,8'd184} : s = 255;
	{8'd71,8'd185} : s = 256;
	{8'd71,8'd186} : s = 257;
	{8'd71,8'd187} : s = 258;
	{8'd71,8'd188} : s = 259;
	{8'd71,8'd189} : s = 260;
	{8'd71,8'd190} : s = 261;
	{8'd71,8'd191} : s = 262;
	{8'd71,8'd192} : s = 263;
	{8'd71,8'd193} : s = 264;
	{8'd71,8'd194} : s = 265;
	{8'd71,8'd195} : s = 266;
	{8'd71,8'd196} : s = 267;
	{8'd71,8'd197} : s = 268;
	{8'd71,8'd198} : s = 269;
	{8'd71,8'd199} : s = 270;
	{8'd71,8'd200} : s = 271;
	{8'd71,8'd201} : s = 272;
	{8'd71,8'd202} : s = 273;
	{8'd71,8'd203} : s = 274;
	{8'd71,8'd204} : s = 275;
	{8'd71,8'd205} : s = 276;
	{8'd71,8'd206} : s = 277;
	{8'd71,8'd207} : s = 278;
	{8'd71,8'd208} : s = 279;
	{8'd71,8'd209} : s = 280;
	{8'd71,8'd210} : s = 281;
	{8'd71,8'd211} : s = 282;
	{8'd71,8'd212} : s = 283;
	{8'd71,8'd213} : s = 284;
	{8'd71,8'd214} : s = 285;
	{8'd71,8'd215} : s = 286;
	{8'd71,8'd216} : s = 287;
	{8'd71,8'd217} : s = 288;
	{8'd71,8'd218} : s = 289;
	{8'd71,8'd219} : s = 290;
	{8'd71,8'd220} : s = 291;
	{8'd71,8'd221} : s = 292;
	{8'd71,8'd222} : s = 293;
	{8'd71,8'd223} : s = 294;
	{8'd71,8'd224} : s = 295;
	{8'd71,8'd225} : s = 296;
	{8'd71,8'd226} : s = 297;
	{8'd71,8'd227} : s = 298;
	{8'd71,8'd228} : s = 299;
	{8'd71,8'd229} : s = 300;
	{8'd71,8'd230} : s = 301;
	{8'd71,8'd231} : s = 302;
	{8'd71,8'd232} : s = 303;
	{8'd71,8'd233} : s = 304;
	{8'd71,8'd234} : s = 305;
	{8'd71,8'd235} : s = 306;
	{8'd71,8'd236} : s = 307;
	{8'd71,8'd237} : s = 308;
	{8'd71,8'd238} : s = 309;
	{8'd71,8'd239} : s = 310;
	{8'd71,8'd240} : s = 311;
	{8'd71,8'd241} : s = 312;
	{8'd71,8'd242} : s = 313;
	{8'd71,8'd243} : s = 314;
	{8'd71,8'd244} : s = 315;
	{8'd71,8'd245} : s = 316;
	{8'd71,8'd246} : s = 317;
	{8'd71,8'd247} : s = 318;
	{8'd71,8'd248} : s = 319;
	{8'd71,8'd249} : s = 320;
	{8'd71,8'd250} : s = 321;
	{8'd71,8'd251} : s = 322;
	{8'd71,8'd252} : s = 323;
	{8'd71,8'd253} : s = 324;
	{8'd71,8'd254} : s = 325;
	{8'd71,8'd255} : s = 326;
	{8'd72,8'd0} : s = 72;
	{8'd72,8'd1} : s = 73;
	{8'd72,8'd2} : s = 74;
	{8'd72,8'd3} : s = 75;
	{8'd72,8'd4} : s = 76;
	{8'd72,8'd5} : s = 77;
	{8'd72,8'd6} : s = 78;
	{8'd72,8'd7} : s = 79;
	{8'd72,8'd8} : s = 80;
	{8'd72,8'd9} : s = 81;
	{8'd72,8'd10} : s = 82;
	{8'd72,8'd11} : s = 83;
	{8'd72,8'd12} : s = 84;
	{8'd72,8'd13} : s = 85;
	{8'd72,8'd14} : s = 86;
	{8'd72,8'd15} : s = 87;
	{8'd72,8'd16} : s = 88;
	{8'd72,8'd17} : s = 89;
	{8'd72,8'd18} : s = 90;
	{8'd72,8'd19} : s = 91;
	{8'd72,8'd20} : s = 92;
	{8'd72,8'd21} : s = 93;
	{8'd72,8'd22} : s = 94;
	{8'd72,8'd23} : s = 95;
	{8'd72,8'd24} : s = 96;
	{8'd72,8'd25} : s = 97;
	{8'd72,8'd26} : s = 98;
	{8'd72,8'd27} : s = 99;
	{8'd72,8'd28} : s = 100;
	{8'd72,8'd29} : s = 101;
	{8'd72,8'd30} : s = 102;
	{8'd72,8'd31} : s = 103;
	{8'd72,8'd32} : s = 104;
	{8'd72,8'd33} : s = 105;
	{8'd72,8'd34} : s = 106;
	{8'd72,8'd35} : s = 107;
	{8'd72,8'd36} : s = 108;
	{8'd72,8'd37} : s = 109;
	{8'd72,8'd38} : s = 110;
	{8'd72,8'd39} : s = 111;
	{8'd72,8'd40} : s = 112;
	{8'd72,8'd41} : s = 113;
	{8'd72,8'd42} : s = 114;
	{8'd72,8'd43} : s = 115;
	{8'd72,8'd44} : s = 116;
	{8'd72,8'd45} : s = 117;
	{8'd72,8'd46} : s = 118;
	{8'd72,8'd47} : s = 119;
	{8'd72,8'd48} : s = 120;
	{8'd72,8'd49} : s = 121;
	{8'd72,8'd50} : s = 122;
	{8'd72,8'd51} : s = 123;
	{8'd72,8'd52} : s = 124;
	{8'd72,8'd53} : s = 125;
	{8'd72,8'd54} : s = 126;
	{8'd72,8'd55} : s = 127;
	{8'd72,8'd56} : s = 128;
	{8'd72,8'd57} : s = 129;
	{8'd72,8'd58} : s = 130;
	{8'd72,8'd59} : s = 131;
	{8'd72,8'd60} : s = 132;
	{8'd72,8'd61} : s = 133;
	{8'd72,8'd62} : s = 134;
	{8'd72,8'd63} : s = 135;
	{8'd72,8'd64} : s = 136;
	{8'd72,8'd65} : s = 137;
	{8'd72,8'd66} : s = 138;
	{8'd72,8'd67} : s = 139;
	{8'd72,8'd68} : s = 140;
	{8'd72,8'd69} : s = 141;
	{8'd72,8'd70} : s = 142;
	{8'd72,8'd71} : s = 143;
	{8'd72,8'd72} : s = 144;
	{8'd72,8'd73} : s = 145;
	{8'd72,8'd74} : s = 146;
	{8'd72,8'd75} : s = 147;
	{8'd72,8'd76} : s = 148;
	{8'd72,8'd77} : s = 149;
	{8'd72,8'd78} : s = 150;
	{8'd72,8'd79} : s = 151;
	{8'd72,8'd80} : s = 152;
	{8'd72,8'd81} : s = 153;
	{8'd72,8'd82} : s = 154;
	{8'd72,8'd83} : s = 155;
	{8'd72,8'd84} : s = 156;
	{8'd72,8'd85} : s = 157;
	{8'd72,8'd86} : s = 158;
	{8'd72,8'd87} : s = 159;
	{8'd72,8'd88} : s = 160;
	{8'd72,8'd89} : s = 161;
	{8'd72,8'd90} : s = 162;
	{8'd72,8'd91} : s = 163;
	{8'd72,8'd92} : s = 164;
	{8'd72,8'd93} : s = 165;
	{8'd72,8'd94} : s = 166;
	{8'd72,8'd95} : s = 167;
	{8'd72,8'd96} : s = 168;
	{8'd72,8'd97} : s = 169;
	{8'd72,8'd98} : s = 170;
	{8'd72,8'd99} : s = 171;
	{8'd72,8'd100} : s = 172;
	{8'd72,8'd101} : s = 173;
	{8'd72,8'd102} : s = 174;
	{8'd72,8'd103} : s = 175;
	{8'd72,8'd104} : s = 176;
	{8'd72,8'd105} : s = 177;
	{8'd72,8'd106} : s = 178;
	{8'd72,8'd107} : s = 179;
	{8'd72,8'd108} : s = 180;
	{8'd72,8'd109} : s = 181;
	{8'd72,8'd110} : s = 182;
	{8'd72,8'd111} : s = 183;
	{8'd72,8'd112} : s = 184;
	{8'd72,8'd113} : s = 185;
	{8'd72,8'd114} : s = 186;
	{8'd72,8'd115} : s = 187;
	{8'd72,8'd116} : s = 188;
	{8'd72,8'd117} : s = 189;
	{8'd72,8'd118} : s = 190;
	{8'd72,8'd119} : s = 191;
	{8'd72,8'd120} : s = 192;
	{8'd72,8'd121} : s = 193;
	{8'd72,8'd122} : s = 194;
	{8'd72,8'd123} : s = 195;
	{8'd72,8'd124} : s = 196;
	{8'd72,8'd125} : s = 197;
	{8'd72,8'd126} : s = 198;
	{8'd72,8'd127} : s = 199;
	{8'd72,8'd128} : s = 200;
	{8'd72,8'd129} : s = 201;
	{8'd72,8'd130} : s = 202;
	{8'd72,8'd131} : s = 203;
	{8'd72,8'd132} : s = 204;
	{8'd72,8'd133} : s = 205;
	{8'd72,8'd134} : s = 206;
	{8'd72,8'd135} : s = 207;
	{8'd72,8'd136} : s = 208;
	{8'd72,8'd137} : s = 209;
	{8'd72,8'd138} : s = 210;
	{8'd72,8'd139} : s = 211;
	{8'd72,8'd140} : s = 212;
	{8'd72,8'd141} : s = 213;
	{8'd72,8'd142} : s = 214;
	{8'd72,8'd143} : s = 215;
	{8'd72,8'd144} : s = 216;
	{8'd72,8'd145} : s = 217;
	{8'd72,8'd146} : s = 218;
	{8'd72,8'd147} : s = 219;
	{8'd72,8'd148} : s = 220;
	{8'd72,8'd149} : s = 221;
	{8'd72,8'd150} : s = 222;
	{8'd72,8'd151} : s = 223;
	{8'd72,8'd152} : s = 224;
	{8'd72,8'd153} : s = 225;
	{8'd72,8'd154} : s = 226;
	{8'd72,8'd155} : s = 227;
	{8'd72,8'd156} : s = 228;
	{8'd72,8'd157} : s = 229;
	{8'd72,8'd158} : s = 230;
	{8'd72,8'd159} : s = 231;
	{8'd72,8'd160} : s = 232;
	{8'd72,8'd161} : s = 233;
	{8'd72,8'd162} : s = 234;
	{8'd72,8'd163} : s = 235;
	{8'd72,8'd164} : s = 236;
	{8'd72,8'd165} : s = 237;
	{8'd72,8'd166} : s = 238;
	{8'd72,8'd167} : s = 239;
	{8'd72,8'd168} : s = 240;
	{8'd72,8'd169} : s = 241;
	{8'd72,8'd170} : s = 242;
	{8'd72,8'd171} : s = 243;
	{8'd72,8'd172} : s = 244;
	{8'd72,8'd173} : s = 245;
	{8'd72,8'd174} : s = 246;
	{8'd72,8'd175} : s = 247;
	{8'd72,8'd176} : s = 248;
	{8'd72,8'd177} : s = 249;
	{8'd72,8'd178} : s = 250;
	{8'd72,8'd179} : s = 251;
	{8'd72,8'd180} : s = 252;
	{8'd72,8'd181} : s = 253;
	{8'd72,8'd182} : s = 254;
	{8'd72,8'd183} : s = 255;
	{8'd72,8'd184} : s = 256;
	{8'd72,8'd185} : s = 257;
	{8'd72,8'd186} : s = 258;
	{8'd72,8'd187} : s = 259;
	{8'd72,8'd188} : s = 260;
	{8'd72,8'd189} : s = 261;
	{8'd72,8'd190} : s = 262;
	{8'd72,8'd191} : s = 263;
	{8'd72,8'd192} : s = 264;
	{8'd72,8'd193} : s = 265;
	{8'd72,8'd194} : s = 266;
	{8'd72,8'd195} : s = 267;
	{8'd72,8'd196} : s = 268;
	{8'd72,8'd197} : s = 269;
	{8'd72,8'd198} : s = 270;
	{8'd72,8'd199} : s = 271;
	{8'd72,8'd200} : s = 272;
	{8'd72,8'd201} : s = 273;
	{8'd72,8'd202} : s = 274;
	{8'd72,8'd203} : s = 275;
	{8'd72,8'd204} : s = 276;
	{8'd72,8'd205} : s = 277;
	{8'd72,8'd206} : s = 278;
	{8'd72,8'd207} : s = 279;
	{8'd72,8'd208} : s = 280;
	{8'd72,8'd209} : s = 281;
	{8'd72,8'd210} : s = 282;
	{8'd72,8'd211} : s = 283;
	{8'd72,8'd212} : s = 284;
	{8'd72,8'd213} : s = 285;
	{8'd72,8'd214} : s = 286;
	{8'd72,8'd215} : s = 287;
	{8'd72,8'd216} : s = 288;
	{8'd72,8'd217} : s = 289;
	{8'd72,8'd218} : s = 290;
	{8'd72,8'd219} : s = 291;
	{8'd72,8'd220} : s = 292;
	{8'd72,8'd221} : s = 293;
	{8'd72,8'd222} : s = 294;
	{8'd72,8'd223} : s = 295;
	{8'd72,8'd224} : s = 296;
	{8'd72,8'd225} : s = 297;
	{8'd72,8'd226} : s = 298;
	{8'd72,8'd227} : s = 299;
	{8'd72,8'd228} : s = 300;
	{8'd72,8'd229} : s = 301;
	{8'd72,8'd230} : s = 302;
	{8'd72,8'd231} : s = 303;
	{8'd72,8'd232} : s = 304;
	{8'd72,8'd233} : s = 305;
	{8'd72,8'd234} : s = 306;
	{8'd72,8'd235} : s = 307;
	{8'd72,8'd236} : s = 308;
	{8'd72,8'd237} : s = 309;
	{8'd72,8'd238} : s = 310;
	{8'd72,8'd239} : s = 311;
	{8'd72,8'd240} : s = 312;
	{8'd72,8'd241} : s = 313;
	{8'd72,8'd242} : s = 314;
	{8'd72,8'd243} : s = 315;
	{8'd72,8'd244} : s = 316;
	{8'd72,8'd245} : s = 317;
	{8'd72,8'd246} : s = 318;
	{8'd72,8'd247} : s = 319;
	{8'd72,8'd248} : s = 320;
	{8'd72,8'd249} : s = 321;
	{8'd72,8'd250} : s = 322;
	{8'd72,8'd251} : s = 323;
	{8'd72,8'd252} : s = 324;
	{8'd72,8'd253} : s = 325;
	{8'd72,8'd254} : s = 326;
	{8'd72,8'd255} : s = 327;
	{8'd73,8'd0} : s = 73;
	{8'd73,8'd1} : s = 74;
	{8'd73,8'd2} : s = 75;
	{8'd73,8'd3} : s = 76;
	{8'd73,8'd4} : s = 77;
	{8'd73,8'd5} : s = 78;
	{8'd73,8'd6} : s = 79;
	{8'd73,8'd7} : s = 80;
	{8'd73,8'd8} : s = 81;
	{8'd73,8'd9} : s = 82;
	{8'd73,8'd10} : s = 83;
	{8'd73,8'd11} : s = 84;
	{8'd73,8'd12} : s = 85;
	{8'd73,8'd13} : s = 86;
	{8'd73,8'd14} : s = 87;
	{8'd73,8'd15} : s = 88;
	{8'd73,8'd16} : s = 89;
	{8'd73,8'd17} : s = 90;
	{8'd73,8'd18} : s = 91;
	{8'd73,8'd19} : s = 92;
	{8'd73,8'd20} : s = 93;
	{8'd73,8'd21} : s = 94;
	{8'd73,8'd22} : s = 95;
	{8'd73,8'd23} : s = 96;
	{8'd73,8'd24} : s = 97;
	{8'd73,8'd25} : s = 98;
	{8'd73,8'd26} : s = 99;
	{8'd73,8'd27} : s = 100;
	{8'd73,8'd28} : s = 101;
	{8'd73,8'd29} : s = 102;
	{8'd73,8'd30} : s = 103;
	{8'd73,8'd31} : s = 104;
	{8'd73,8'd32} : s = 105;
	{8'd73,8'd33} : s = 106;
	{8'd73,8'd34} : s = 107;
	{8'd73,8'd35} : s = 108;
	{8'd73,8'd36} : s = 109;
	{8'd73,8'd37} : s = 110;
	{8'd73,8'd38} : s = 111;
	{8'd73,8'd39} : s = 112;
	{8'd73,8'd40} : s = 113;
	{8'd73,8'd41} : s = 114;
	{8'd73,8'd42} : s = 115;
	{8'd73,8'd43} : s = 116;
	{8'd73,8'd44} : s = 117;
	{8'd73,8'd45} : s = 118;
	{8'd73,8'd46} : s = 119;
	{8'd73,8'd47} : s = 120;
	{8'd73,8'd48} : s = 121;
	{8'd73,8'd49} : s = 122;
	{8'd73,8'd50} : s = 123;
	{8'd73,8'd51} : s = 124;
	{8'd73,8'd52} : s = 125;
	{8'd73,8'd53} : s = 126;
	{8'd73,8'd54} : s = 127;
	{8'd73,8'd55} : s = 128;
	{8'd73,8'd56} : s = 129;
	{8'd73,8'd57} : s = 130;
	{8'd73,8'd58} : s = 131;
	{8'd73,8'd59} : s = 132;
	{8'd73,8'd60} : s = 133;
	{8'd73,8'd61} : s = 134;
	{8'd73,8'd62} : s = 135;
	{8'd73,8'd63} : s = 136;
	{8'd73,8'd64} : s = 137;
	{8'd73,8'd65} : s = 138;
	{8'd73,8'd66} : s = 139;
	{8'd73,8'd67} : s = 140;
	{8'd73,8'd68} : s = 141;
	{8'd73,8'd69} : s = 142;
	{8'd73,8'd70} : s = 143;
	{8'd73,8'd71} : s = 144;
	{8'd73,8'd72} : s = 145;
	{8'd73,8'd73} : s = 146;
	{8'd73,8'd74} : s = 147;
	{8'd73,8'd75} : s = 148;
	{8'd73,8'd76} : s = 149;
	{8'd73,8'd77} : s = 150;
	{8'd73,8'd78} : s = 151;
	{8'd73,8'd79} : s = 152;
	{8'd73,8'd80} : s = 153;
	{8'd73,8'd81} : s = 154;
	{8'd73,8'd82} : s = 155;
	{8'd73,8'd83} : s = 156;
	{8'd73,8'd84} : s = 157;
	{8'd73,8'd85} : s = 158;
	{8'd73,8'd86} : s = 159;
	{8'd73,8'd87} : s = 160;
	{8'd73,8'd88} : s = 161;
	{8'd73,8'd89} : s = 162;
	{8'd73,8'd90} : s = 163;
	{8'd73,8'd91} : s = 164;
	{8'd73,8'd92} : s = 165;
	{8'd73,8'd93} : s = 166;
	{8'd73,8'd94} : s = 167;
	{8'd73,8'd95} : s = 168;
	{8'd73,8'd96} : s = 169;
	{8'd73,8'd97} : s = 170;
	{8'd73,8'd98} : s = 171;
	{8'd73,8'd99} : s = 172;
	{8'd73,8'd100} : s = 173;
	{8'd73,8'd101} : s = 174;
	{8'd73,8'd102} : s = 175;
	{8'd73,8'd103} : s = 176;
	{8'd73,8'd104} : s = 177;
	{8'd73,8'd105} : s = 178;
	{8'd73,8'd106} : s = 179;
	{8'd73,8'd107} : s = 180;
	{8'd73,8'd108} : s = 181;
	{8'd73,8'd109} : s = 182;
	{8'd73,8'd110} : s = 183;
	{8'd73,8'd111} : s = 184;
	{8'd73,8'd112} : s = 185;
	{8'd73,8'd113} : s = 186;
	{8'd73,8'd114} : s = 187;
	{8'd73,8'd115} : s = 188;
	{8'd73,8'd116} : s = 189;
	{8'd73,8'd117} : s = 190;
	{8'd73,8'd118} : s = 191;
	{8'd73,8'd119} : s = 192;
	{8'd73,8'd120} : s = 193;
	{8'd73,8'd121} : s = 194;
	{8'd73,8'd122} : s = 195;
	{8'd73,8'd123} : s = 196;
	{8'd73,8'd124} : s = 197;
	{8'd73,8'd125} : s = 198;
	{8'd73,8'd126} : s = 199;
	{8'd73,8'd127} : s = 200;
	{8'd73,8'd128} : s = 201;
	{8'd73,8'd129} : s = 202;
	{8'd73,8'd130} : s = 203;
	{8'd73,8'd131} : s = 204;
	{8'd73,8'd132} : s = 205;
	{8'd73,8'd133} : s = 206;
	{8'd73,8'd134} : s = 207;
	{8'd73,8'd135} : s = 208;
	{8'd73,8'd136} : s = 209;
	{8'd73,8'd137} : s = 210;
	{8'd73,8'd138} : s = 211;
	{8'd73,8'd139} : s = 212;
	{8'd73,8'd140} : s = 213;
	{8'd73,8'd141} : s = 214;
	{8'd73,8'd142} : s = 215;
	{8'd73,8'd143} : s = 216;
	{8'd73,8'd144} : s = 217;
	{8'd73,8'd145} : s = 218;
	{8'd73,8'd146} : s = 219;
	{8'd73,8'd147} : s = 220;
	{8'd73,8'd148} : s = 221;
	{8'd73,8'd149} : s = 222;
	{8'd73,8'd150} : s = 223;
	{8'd73,8'd151} : s = 224;
	{8'd73,8'd152} : s = 225;
	{8'd73,8'd153} : s = 226;
	{8'd73,8'd154} : s = 227;
	{8'd73,8'd155} : s = 228;
	{8'd73,8'd156} : s = 229;
	{8'd73,8'd157} : s = 230;
	{8'd73,8'd158} : s = 231;
	{8'd73,8'd159} : s = 232;
	{8'd73,8'd160} : s = 233;
	{8'd73,8'd161} : s = 234;
	{8'd73,8'd162} : s = 235;
	{8'd73,8'd163} : s = 236;
	{8'd73,8'd164} : s = 237;
	{8'd73,8'd165} : s = 238;
	{8'd73,8'd166} : s = 239;
	{8'd73,8'd167} : s = 240;
	{8'd73,8'd168} : s = 241;
	{8'd73,8'd169} : s = 242;
	{8'd73,8'd170} : s = 243;
	{8'd73,8'd171} : s = 244;
	{8'd73,8'd172} : s = 245;
	{8'd73,8'd173} : s = 246;
	{8'd73,8'd174} : s = 247;
	{8'd73,8'd175} : s = 248;
	{8'd73,8'd176} : s = 249;
	{8'd73,8'd177} : s = 250;
	{8'd73,8'd178} : s = 251;
	{8'd73,8'd179} : s = 252;
	{8'd73,8'd180} : s = 253;
	{8'd73,8'd181} : s = 254;
	{8'd73,8'd182} : s = 255;
	{8'd73,8'd183} : s = 256;
	{8'd73,8'd184} : s = 257;
	{8'd73,8'd185} : s = 258;
	{8'd73,8'd186} : s = 259;
	{8'd73,8'd187} : s = 260;
	{8'd73,8'd188} : s = 261;
	{8'd73,8'd189} : s = 262;
	{8'd73,8'd190} : s = 263;
	{8'd73,8'd191} : s = 264;
	{8'd73,8'd192} : s = 265;
	{8'd73,8'd193} : s = 266;
	{8'd73,8'd194} : s = 267;
	{8'd73,8'd195} : s = 268;
	{8'd73,8'd196} : s = 269;
	{8'd73,8'd197} : s = 270;
	{8'd73,8'd198} : s = 271;
	{8'd73,8'd199} : s = 272;
	{8'd73,8'd200} : s = 273;
	{8'd73,8'd201} : s = 274;
	{8'd73,8'd202} : s = 275;
	{8'd73,8'd203} : s = 276;
	{8'd73,8'd204} : s = 277;
	{8'd73,8'd205} : s = 278;
	{8'd73,8'd206} : s = 279;
	{8'd73,8'd207} : s = 280;
	{8'd73,8'd208} : s = 281;
	{8'd73,8'd209} : s = 282;
	{8'd73,8'd210} : s = 283;
	{8'd73,8'd211} : s = 284;
	{8'd73,8'd212} : s = 285;
	{8'd73,8'd213} : s = 286;
	{8'd73,8'd214} : s = 287;
	{8'd73,8'd215} : s = 288;
	{8'd73,8'd216} : s = 289;
	{8'd73,8'd217} : s = 290;
	{8'd73,8'd218} : s = 291;
	{8'd73,8'd219} : s = 292;
	{8'd73,8'd220} : s = 293;
	{8'd73,8'd221} : s = 294;
	{8'd73,8'd222} : s = 295;
	{8'd73,8'd223} : s = 296;
	{8'd73,8'd224} : s = 297;
	{8'd73,8'd225} : s = 298;
	{8'd73,8'd226} : s = 299;
	{8'd73,8'd227} : s = 300;
	{8'd73,8'd228} : s = 301;
	{8'd73,8'd229} : s = 302;
	{8'd73,8'd230} : s = 303;
	{8'd73,8'd231} : s = 304;
	{8'd73,8'd232} : s = 305;
	{8'd73,8'd233} : s = 306;
	{8'd73,8'd234} : s = 307;
	{8'd73,8'd235} : s = 308;
	{8'd73,8'd236} : s = 309;
	{8'd73,8'd237} : s = 310;
	{8'd73,8'd238} : s = 311;
	{8'd73,8'd239} : s = 312;
	{8'd73,8'd240} : s = 313;
	{8'd73,8'd241} : s = 314;
	{8'd73,8'd242} : s = 315;
	{8'd73,8'd243} : s = 316;
	{8'd73,8'd244} : s = 317;
	{8'd73,8'd245} : s = 318;
	{8'd73,8'd246} : s = 319;
	{8'd73,8'd247} : s = 320;
	{8'd73,8'd248} : s = 321;
	{8'd73,8'd249} : s = 322;
	{8'd73,8'd250} : s = 323;
	{8'd73,8'd251} : s = 324;
	{8'd73,8'd252} : s = 325;
	{8'd73,8'd253} : s = 326;
	{8'd73,8'd254} : s = 327;
	{8'd73,8'd255} : s = 328;
	{8'd74,8'd0} : s = 74;
	{8'd74,8'd1} : s = 75;
	{8'd74,8'd2} : s = 76;
	{8'd74,8'd3} : s = 77;
	{8'd74,8'd4} : s = 78;
	{8'd74,8'd5} : s = 79;
	{8'd74,8'd6} : s = 80;
	{8'd74,8'd7} : s = 81;
	{8'd74,8'd8} : s = 82;
	{8'd74,8'd9} : s = 83;
	{8'd74,8'd10} : s = 84;
	{8'd74,8'd11} : s = 85;
	{8'd74,8'd12} : s = 86;
	{8'd74,8'd13} : s = 87;
	{8'd74,8'd14} : s = 88;
	{8'd74,8'd15} : s = 89;
	{8'd74,8'd16} : s = 90;
	{8'd74,8'd17} : s = 91;
	{8'd74,8'd18} : s = 92;
	{8'd74,8'd19} : s = 93;
	{8'd74,8'd20} : s = 94;
	{8'd74,8'd21} : s = 95;
	{8'd74,8'd22} : s = 96;
	{8'd74,8'd23} : s = 97;
	{8'd74,8'd24} : s = 98;
	{8'd74,8'd25} : s = 99;
	{8'd74,8'd26} : s = 100;
	{8'd74,8'd27} : s = 101;
	{8'd74,8'd28} : s = 102;
	{8'd74,8'd29} : s = 103;
	{8'd74,8'd30} : s = 104;
	{8'd74,8'd31} : s = 105;
	{8'd74,8'd32} : s = 106;
	{8'd74,8'd33} : s = 107;
	{8'd74,8'd34} : s = 108;
	{8'd74,8'd35} : s = 109;
	{8'd74,8'd36} : s = 110;
	{8'd74,8'd37} : s = 111;
	{8'd74,8'd38} : s = 112;
	{8'd74,8'd39} : s = 113;
	{8'd74,8'd40} : s = 114;
	{8'd74,8'd41} : s = 115;
	{8'd74,8'd42} : s = 116;
	{8'd74,8'd43} : s = 117;
	{8'd74,8'd44} : s = 118;
	{8'd74,8'd45} : s = 119;
	{8'd74,8'd46} : s = 120;
	{8'd74,8'd47} : s = 121;
	{8'd74,8'd48} : s = 122;
	{8'd74,8'd49} : s = 123;
	{8'd74,8'd50} : s = 124;
	{8'd74,8'd51} : s = 125;
	{8'd74,8'd52} : s = 126;
	{8'd74,8'd53} : s = 127;
	{8'd74,8'd54} : s = 128;
	{8'd74,8'd55} : s = 129;
	{8'd74,8'd56} : s = 130;
	{8'd74,8'd57} : s = 131;
	{8'd74,8'd58} : s = 132;
	{8'd74,8'd59} : s = 133;
	{8'd74,8'd60} : s = 134;
	{8'd74,8'd61} : s = 135;
	{8'd74,8'd62} : s = 136;
	{8'd74,8'd63} : s = 137;
	{8'd74,8'd64} : s = 138;
	{8'd74,8'd65} : s = 139;
	{8'd74,8'd66} : s = 140;
	{8'd74,8'd67} : s = 141;
	{8'd74,8'd68} : s = 142;
	{8'd74,8'd69} : s = 143;
	{8'd74,8'd70} : s = 144;
	{8'd74,8'd71} : s = 145;
	{8'd74,8'd72} : s = 146;
	{8'd74,8'd73} : s = 147;
	{8'd74,8'd74} : s = 148;
	{8'd74,8'd75} : s = 149;
	{8'd74,8'd76} : s = 150;
	{8'd74,8'd77} : s = 151;
	{8'd74,8'd78} : s = 152;
	{8'd74,8'd79} : s = 153;
	{8'd74,8'd80} : s = 154;
	{8'd74,8'd81} : s = 155;
	{8'd74,8'd82} : s = 156;
	{8'd74,8'd83} : s = 157;
	{8'd74,8'd84} : s = 158;
	{8'd74,8'd85} : s = 159;
	{8'd74,8'd86} : s = 160;
	{8'd74,8'd87} : s = 161;
	{8'd74,8'd88} : s = 162;
	{8'd74,8'd89} : s = 163;
	{8'd74,8'd90} : s = 164;
	{8'd74,8'd91} : s = 165;
	{8'd74,8'd92} : s = 166;
	{8'd74,8'd93} : s = 167;
	{8'd74,8'd94} : s = 168;
	{8'd74,8'd95} : s = 169;
	{8'd74,8'd96} : s = 170;
	{8'd74,8'd97} : s = 171;
	{8'd74,8'd98} : s = 172;
	{8'd74,8'd99} : s = 173;
	{8'd74,8'd100} : s = 174;
	{8'd74,8'd101} : s = 175;
	{8'd74,8'd102} : s = 176;
	{8'd74,8'd103} : s = 177;
	{8'd74,8'd104} : s = 178;
	{8'd74,8'd105} : s = 179;
	{8'd74,8'd106} : s = 180;
	{8'd74,8'd107} : s = 181;
	{8'd74,8'd108} : s = 182;
	{8'd74,8'd109} : s = 183;
	{8'd74,8'd110} : s = 184;
	{8'd74,8'd111} : s = 185;
	{8'd74,8'd112} : s = 186;
	{8'd74,8'd113} : s = 187;
	{8'd74,8'd114} : s = 188;
	{8'd74,8'd115} : s = 189;
	{8'd74,8'd116} : s = 190;
	{8'd74,8'd117} : s = 191;
	{8'd74,8'd118} : s = 192;
	{8'd74,8'd119} : s = 193;
	{8'd74,8'd120} : s = 194;
	{8'd74,8'd121} : s = 195;
	{8'd74,8'd122} : s = 196;
	{8'd74,8'd123} : s = 197;
	{8'd74,8'd124} : s = 198;
	{8'd74,8'd125} : s = 199;
	{8'd74,8'd126} : s = 200;
	{8'd74,8'd127} : s = 201;
	{8'd74,8'd128} : s = 202;
	{8'd74,8'd129} : s = 203;
	{8'd74,8'd130} : s = 204;
	{8'd74,8'd131} : s = 205;
	{8'd74,8'd132} : s = 206;
	{8'd74,8'd133} : s = 207;
	{8'd74,8'd134} : s = 208;
	{8'd74,8'd135} : s = 209;
	{8'd74,8'd136} : s = 210;
	{8'd74,8'd137} : s = 211;
	{8'd74,8'd138} : s = 212;
	{8'd74,8'd139} : s = 213;
	{8'd74,8'd140} : s = 214;
	{8'd74,8'd141} : s = 215;
	{8'd74,8'd142} : s = 216;
	{8'd74,8'd143} : s = 217;
	{8'd74,8'd144} : s = 218;
	{8'd74,8'd145} : s = 219;
	{8'd74,8'd146} : s = 220;
	{8'd74,8'd147} : s = 221;
	{8'd74,8'd148} : s = 222;
	{8'd74,8'd149} : s = 223;
	{8'd74,8'd150} : s = 224;
	{8'd74,8'd151} : s = 225;
	{8'd74,8'd152} : s = 226;
	{8'd74,8'd153} : s = 227;
	{8'd74,8'd154} : s = 228;
	{8'd74,8'd155} : s = 229;
	{8'd74,8'd156} : s = 230;
	{8'd74,8'd157} : s = 231;
	{8'd74,8'd158} : s = 232;
	{8'd74,8'd159} : s = 233;
	{8'd74,8'd160} : s = 234;
	{8'd74,8'd161} : s = 235;
	{8'd74,8'd162} : s = 236;
	{8'd74,8'd163} : s = 237;
	{8'd74,8'd164} : s = 238;
	{8'd74,8'd165} : s = 239;
	{8'd74,8'd166} : s = 240;
	{8'd74,8'd167} : s = 241;
	{8'd74,8'd168} : s = 242;
	{8'd74,8'd169} : s = 243;
	{8'd74,8'd170} : s = 244;
	{8'd74,8'd171} : s = 245;
	{8'd74,8'd172} : s = 246;
	{8'd74,8'd173} : s = 247;
	{8'd74,8'd174} : s = 248;
	{8'd74,8'd175} : s = 249;
	{8'd74,8'd176} : s = 250;
	{8'd74,8'd177} : s = 251;
	{8'd74,8'd178} : s = 252;
	{8'd74,8'd179} : s = 253;
	{8'd74,8'd180} : s = 254;
	{8'd74,8'd181} : s = 255;
	{8'd74,8'd182} : s = 256;
	{8'd74,8'd183} : s = 257;
	{8'd74,8'd184} : s = 258;
	{8'd74,8'd185} : s = 259;
	{8'd74,8'd186} : s = 260;
	{8'd74,8'd187} : s = 261;
	{8'd74,8'd188} : s = 262;
	{8'd74,8'd189} : s = 263;
	{8'd74,8'd190} : s = 264;
	{8'd74,8'd191} : s = 265;
	{8'd74,8'd192} : s = 266;
	{8'd74,8'd193} : s = 267;
	{8'd74,8'd194} : s = 268;
	{8'd74,8'd195} : s = 269;
	{8'd74,8'd196} : s = 270;
	{8'd74,8'd197} : s = 271;
	{8'd74,8'd198} : s = 272;
	{8'd74,8'd199} : s = 273;
	{8'd74,8'd200} : s = 274;
	{8'd74,8'd201} : s = 275;
	{8'd74,8'd202} : s = 276;
	{8'd74,8'd203} : s = 277;
	{8'd74,8'd204} : s = 278;
	{8'd74,8'd205} : s = 279;
	{8'd74,8'd206} : s = 280;
	{8'd74,8'd207} : s = 281;
	{8'd74,8'd208} : s = 282;
	{8'd74,8'd209} : s = 283;
	{8'd74,8'd210} : s = 284;
	{8'd74,8'd211} : s = 285;
	{8'd74,8'd212} : s = 286;
	{8'd74,8'd213} : s = 287;
	{8'd74,8'd214} : s = 288;
	{8'd74,8'd215} : s = 289;
	{8'd74,8'd216} : s = 290;
	{8'd74,8'd217} : s = 291;
	{8'd74,8'd218} : s = 292;
	{8'd74,8'd219} : s = 293;
	{8'd74,8'd220} : s = 294;
	{8'd74,8'd221} : s = 295;
	{8'd74,8'd222} : s = 296;
	{8'd74,8'd223} : s = 297;
	{8'd74,8'd224} : s = 298;
	{8'd74,8'd225} : s = 299;
	{8'd74,8'd226} : s = 300;
	{8'd74,8'd227} : s = 301;
	{8'd74,8'd228} : s = 302;
	{8'd74,8'd229} : s = 303;
	{8'd74,8'd230} : s = 304;
	{8'd74,8'd231} : s = 305;
	{8'd74,8'd232} : s = 306;
	{8'd74,8'd233} : s = 307;
	{8'd74,8'd234} : s = 308;
	{8'd74,8'd235} : s = 309;
	{8'd74,8'd236} : s = 310;
	{8'd74,8'd237} : s = 311;
	{8'd74,8'd238} : s = 312;
	{8'd74,8'd239} : s = 313;
	{8'd74,8'd240} : s = 314;
	{8'd74,8'd241} : s = 315;
	{8'd74,8'd242} : s = 316;
	{8'd74,8'd243} : s = 317;
	{8'd74,8'd244} : s = 318;
	{8'd74,8'd245} : s = 319;
	{8'd74,8'd246} : s = 320;
	{8'd74,8'd247} : s = 321;
	{8'd74,8'd248} : s = 322;
	{8'd74,8'd249} : s = 323;
	{8'd74,8'd250} : s = 324;
	{8'd74,8'd251} : s = 325;
	{8'd74,8'd252} : s = 326;
	{8'd74,8'd253} : s = 327;
	{8'd74,8'd254} : s = 328;
	{8'd74,8'd255} : s = 329;
	{8'd75,8'd0} : s = 75;
	{8'd75,8'd1} : s = 76;
	{8'd75,8'd2} : s = 77;
	{8'd75,8'd3} : s = 78;
	{8'd75,8'd4} : s = 79;
	{8'd75,8'd5} : s = 80;
	{8'd75,8'd6} : s = 81;
	{8'd75,8'd7} : s = 82;
	{8'd75,8'd8} : s = 83;
	{8'd75,8'd9} : s = 84;
	{8'd75,8'd10} : s = 85;
	{8'd75,8'd11} : s = 86;
	{8'd75,8'd12} : s = 87;
	{8'd75,8'd13} : s = 88;
	{8'd75,8'd14} : s = 89;
	{8'd75,8'd15} : s = 90;
	{8'd75,8'd16} : s = 91;
	{8'd75,8'd17} : s = 92;
	{8'd75,8'd18} : s = 93;
	{8'd75,8'd19} : s = 94;
	{8'd75,8'd20} : s = 95;
	{8'd75,8'd21} : s = 96;
	{8'd75,8'd22} : s = 97;
	{8'd75,8'd23} : s = 98;
	{8'd75,8'd24} : s = 99;
	{8'd75,8'd25} : s = 100;
	{8'd75,8'd26} : s = 101;
	{8'd75,8'd27} : s = 102;
	{8'd75,8'd28} : s = 103;
	{8'd75,8'd29} : s = 104;
	{8'd75,8'd30} : s = 105;
	{8'd75,8'd31} : s = 106;
	{8'd75,8'd32} : s = 107;
	{8'd75,8'd33} : s = 108;
	{8'd75,8'd34} : s = 109;
	{8'd75,8'd35} : s = 110;
	{8'd75,8'd36} : s = 111;
	{8'd75,8'd37} : s = 112;
	{8'd75,8'd38} : s = 113;
	{8'd75,8'd39} : s = 114;
	{8'd75,8'd40} : s = 115;
	{8'd75,8'd41} : s = 116;
	{8'd75,8'd42} : s = 117;
	{8'd75,8'd43} : s = 118;
	{8'd75,8'd44} : s = 119;
	{8'd75,8'd45} : s = 120;
	{8'd75,8'd46} : s = 121;
	{8'd75,8'd47} : s = 122;
	{8'd75,8'd48} : s = 123;
	{8'd75,8'd49} : s = 124;
	{8'd75,8'd50} : s = 125;
	{8'd75,8'd51} : s = 126;
	{8'd75,8'd52} : s = 127;
	{8'd75,8'd53} : s = 128;
	{8'd75,8'd54} : s = 129;
	{8'd75,8'd55} : s = 130;
	{8'd75,8'd56} : s = 131;
	{8'd75,8'd57} : s = 132;
	{8'd75,8'd58} : s = 133;
	{8'd75,8'd59} : s = 134;
	{8'd75,8'd60} : s = 135;
	{8'd75,8'd61} : s = 136;
	{8'd75,8'd62} : s = 137;
	{8'd75,8'd63} : s = 138;
	{8'd75,8'd64} : s = 139;
	{8'd75,8'd65} : s = 140;
	{8'd75,8'd66} : s = 141;
	{8'd75,8'd67} : s = 142;
	{8'd75,8'd68} : s = 143;
	{8'd75,8'd69} : s = 144;
	{8'd75,8'd70} : s = 145;
	{8'd75,8'd71} : s = 146;
	{8'd75,8'd72} : s = 147;
	{8'd75,8'd73} : s = 148;
	{8'd75,8'd74} : s = 149;
	{8'd75,8'd75} : s = 150;
	{8'd75,8'd76} : s = 151;
	{8'd75,8'd77} : s = 152;
	{8'd75,8'd78} : s = 153;
	{8'd75,8'd79} : s = 154;
	{8'd75,8'd80} : s = 155;
	{8'd75,8'd81} : s = 156;
	{8'd75,8'd82} : s = 157;
	{8'd75,8'd83} : s = 158;
	{8'd75,8'd84} : s = 159;
	{8'd75,8'd85} : s = 160;
	{8'd75,8'd86} : s = 161;
	{8'd75,8'd87} : s = 162;
	{8'd75,8'd88} : s = 163;
	{8'd75,8'd89} : s = 164;
	{8'd75,8'd90} : s = 165;
	{8'd75,8'd91} : s = 166;
	{8'd75,8'd92} : s = 167;
	{8'd75,8'd93} : s = 168;
	{8'd75,8'd94} : s = 169;
	{8'd75,8'd95} : s = 170;
	{8'd75,8'd96} : s = 171;
	{8'd75,8'd97} : s = 172;
	{8'd75,8'd98} : s = 173;
	{8'd75,8'd99} : s = 174;
	{8'd75,8'd100} : s = 175;
	{8'd75,8'd101} : s = 176;
	{8'd75,8'd102} : s = 177;
	{8'd75,8'd103} : s = 178;
	{8'd75,8'd104} : s = 179;
	{8'd75,8'd105} : s = 180;
	{8'd75,8'd106} : s = 181;
	{8'd75,8'd107} : s = 182;
	{8'd75,8'd108} : s = 183;
	{8'd75,8'd109} : s = 184;
	{8'd75,8'd110} : s = 185;
	{8'd75,8'd111} : s = 186;
	{8'd75,8'd112} : s = 187;
	{8'd75,8'd113} : s = 188;
	{8'd75,8'd114} : s = 189;
	{8'd75,8'd115} : s = 190;
	{8'd75,8'd116} : s = 191;
	{8'd75,8'd117} : s = 192;
	{8'd75,8'd118} : s = 193;
	{8'd75,8'd119} : s = 194;
	{8'd75,8'd120} : s = 195;
	{8'd75,8'd121} : s = 196;
	{8'd75,8'd122} : s = 197;
	{8'd75,8'd123} : s = 198;
	{8'd75,8'd124} : s = 199;
	{8'd75,8'd125} : s = 200;
	{8'd75,8'd126} : s = 201;
	{8'd75,8'd127} : s = 202;
	{8'd75,8'd128} : s = 203;
	{8'd75,8'd129} : s = 204;
	{8'd75,8'd130} : s = 205;
	{8'd75,8'd131} : s = 206;
	{8'd75,8'd132} : s = 207;
	{8'd75,8'd133} : s = 208;
	{8'd75,8'd134} : s = 209;
	{8'd75,8'd135} : s = 210;
	{8'd75,8'd136} : s = 211;
	{8'd75,8'd137} : s = 212;
	{8'd75,8'd138} : s = 213;
	{8'd75,8'd139} : s = 214;
	{8'd75,8'd140} : s = 215;
	{8'd75,8'd141} : s = 216;
	{8'd75,8'd142} : s = 217;
	{8'd75,8'd143} : s = 218;
	{8'd75,8'd144} : s = 219;
	{8'd75,8'd145} : s = 220;
	{8'd75,8'd146} : s = 221;
	{8'd75,8'd147} : s = 222;
	{8'd75,8'd148} : s = 223;
	{8'd75,8'd149} : s = 224;
	{8'd75,8'd150} : s = 225;
	{8'd75,8'd151} : s = 226;
	{8'd75,8'd152} : s = 227;
	{8'd75,8'd153} : s = 228;
	{8'd75,8'd154} : s = 229;
	{8'd75,8'd155} : s = 230;
	{8'd75,8'd156} : s = 231;
	{8'd75,8'd157} : s = 232;
	{8'd75,8'd158} : s = 233;
	{8'd75,8'd159} : s = 234;
	{8'd75,8'd160} : s = 235;
	{8'd75,8'd161} : s = 236;
	{8'd75,8'd162} : s = 237;
	{8'd75,8'd163} : s = 238;
	{8'd75,8'd164} : s = 239;
	{8'd75,8'd165} : s = 240;
	{8'd75,8'd166} : s = 241;
	{8'd75,8'd167} : s = 242;
	{8'd75,8'd168} : s = 243;
	{8'd75,8'd169} : s = 244;
	{8'd75,8'd170} : s = 245;
	{8'd75,8'd171} : s = 246;
	{8'd75,8'd172} : s = 247;
	{8'd75,8'd173} : s = 248;
	{8'd75,8'd174} : s = 249;
	{8'd75,8'd175} : s = 250;
	{8'd75,8'd176} : s = 251;
	{8'd75,8'd177} : s = 252;
	{8'd75,8'd178} : s = 253;
	{8'd75,8'd179} : s = 254;
	{8'd75,8'd180} : s = 255;
	{8'd75,8'd181} : s = 256;
	{8'd75,8'd182} : s = 257;
	{8'd75,8'd183} : s = 258;
	{8'd75,8'd184} : s = 259;
	{8'd75,8'd185} : s = 260;
	{8'd75,8'd186} : s = 261;
	{8'd75,8'd187} : s = 262;
	{8'd75,8'd188} : s = 263;
	{8'd75,8'd189} : s = 264;
	{8'd75,8'd190} : s = 265;
	{8'd75,8'd191} : s = 266;
	{8'd75,8'd192} : s = 267;
	{8'd75,8'd193} : s = 268;
	{8'd75,8'd194} : s = 269;
	{8'd75,8'd195} : s = 270;
	{8'd75,8'd196} : s = 271;
	{8'd75,8'd197} : s = 272;
	{8'd75,8'd198} : s = 273;
	{8'd75,8'd199} : s = 274;
	{8'd75,8'd200} : s = 275;
	{8'd75,8'd201} : s = 276;
	{8'd75,8'd202} : s = 277;
	{8'd75,8'd203} : s = 278;
	{8'd75,8'd204} : s = 279;
	{8'd75,8'd205} : s = 280;
	{8'd75,8'd206} : s = 281;
	{8'd75,8'd207} : s = 282;
	{8'd75,8'd208} : s = 283;
	{8'd75,8'd209} : s = 284;
	{8'd75,8'd210} : s = 285;
	{8'd75,8'd211} : s = 286;
	{8'd75,8'd212} : s = 287;
	{8'd75,8'd213} : s = 288;
	{8'd75,8'd214} : s = 289;
	{8'd75,8'd215} : s = 290;
	{8'd75,8'd216} : s = 291;
	{8'd75,8'd217} : s = 292;
	{8'd75,8'd218} : s = 293;
	{8'd75,8'd219} : s = 294;
	{8'd75,8'd220} : s = 295;
	{8'd75,8'd221} : s = 296;
	{8'd75,8'd222} : s = 297;
	{8'd75,8'd223} : s = 298;
	{8'd75,8'd224} : s = 299;
	{8'd75,8'd225} : s = 300;
	{8'd75,8'd226} : s = 301;
	{8'd75,8'd227} : s = 302;
	{8'd75,8'd228} : s = 303;
	{8'd75,8'd229} : s = 304;
	{8'd75,8'd230} : s = 305;
	{8'd75,8'd231} : s = 306;
	{8'd75,8'd232} : s = 307;
	{8'd75,8'd233} : s = 308;
	{8'd75,8'd234} : s = 309;
	{8'd75,8'd235} : s = 310;
	{8'd75,8'd236} : s = 311;
	{8'd75,8'd237} : s = 312;
	{8'd75,8'd238} : s = 313;
	{8'd75,8'd239} : s = 314;
	{8'd75,8'd240} : s = 315;
	{8'd75,8'd241} : s = 316;
	{8'd75,8'd242} : s = 317;
	{8'd75,8'd243} : s = 318;
	{8'd75,8'd244} : s = 319;
	{8'd75,8'd245} : s = 320;
	{8'd75,8'd246} : s = 321;
	{8'd75,8'd247} : s = 322;
	{8'd75,8'd248} : s = 323;
	{8'd75,8'd249} : s = 324;
	{8'd75,8'd250} : s = 325;
	{8'd75,8'd251} : s = 326;
	{8'd75,8'd252} : s = 327;
	{8'd75,8'd253} : s = 328;
	{8'd75,8'd254} : s = 329;
	{8'd75,8'd255} : s = 330;
	{8'd76,8'd0} : s = 76;
	{8'd76,8'd1} : s = 77;
	{8'd76,8'd2} : s = 78;
	{8'd76,8'd3} : s = 79;
	{8'd76,8'd4} : s = 80;
	{8'd76,8'd5} : s = 81;
	{8'd76,8'd6} : s = 82;
	{8'd76,8'd7} : s = 83;
	{8'd76,8'd8} : s = 84;
	{8'd76,8'd9} : s = 85;
	{8'd76,8'd10} : s = 86;
	{8'd76,8'd11} : s = 87;
	{8'd76,8'd12} : s = 88;
	{8'd76,8'd13} : s = 89;
	{8'd76,8'd14} : s = 90;
	{8'd76,8'd15} : s = 91;
	{8'd76,8'd16} : s = 92;
	{8'd76,8'd17} : s = 93;
	{8'd76,8'd18} : s = 94;
	{8'd76,8'd19} : s = 95;
	{8'd76,8'd20} : s = 96;
	{8'd76,8'd21} : s = 97;
	{8'd76,8'd22} : s = 98;
	{8'd76,8'd23} : s = 99;
	{8'd76,8'd24} : s = 100;
	{8'd76,8'd25} : s = 101;
	{8'd76,8'd26} : s = 102;
	{8'd76,8'd27} : s = 103;
	{8'd76,8'd28} : s = 104;
	{8'd76,8'd29} : s = 105;
	{8'd76,8'd30} : s = 106;
	{8'd76,8'd31} : s = 107;
	{8'd76,8'd32} : s = 108;
	{8'd76,8'd33} : s = 109;
	{8'd76,8'd34} : s = 110;
	{8'd76,8'd35} : s = 111;
	{8'd76,8'd36} : s = 112;
	{8'd76,8'd37} : s = 113;
	{8'd76,8'd38} : s = 114;
	{8'd76,8'd39} : s = 115;
	{8'd76,8'd40} : s = 116;
	{8'd76,8'd41} : s = 117;
	{8'd76,8'd42} : s = 118;
	{8'd76,8'd43} : s = 119;
	{8'd76,8'd44} : s = 120;
	{8'd76,8'd45} : s = 121;
	{8'd76,8'd46} : s = 122;
	{8'd76,8'd47} : s = 123;
	{8'd76,8'd48} : s = 124;
	{8'd76,8'd49} : s = 125;
	{8'd76,8'd50} : s = 126;
	{8'd76,8'd51} : s = 127;
	{8'd76,8'd52} : s = 128;
	{8'd76,8'd53} : s = 129;
	{8'd76,8'd54} : s = 130;
	{8'd76,8'd55} : s = 131;
	{8'd76,8'd56} : s = 132;
	{8'd76,8'd57} : s = 133;
	{8'd76,8'd58} : s = 134;
	{8'd76,8'd59} : s = 135;
	{8'd76,8'd60} : s = 136;
	{8'd76,8'd61} : s = 137;
	{8'd76,8'd62} : s = 138;
	{8'd76,8'd63} : s = 139;
	{8'd76,8'd64} : s = 140;
	{8'd76,8'd65} : s = 141;
	{8'd76,8'd66} : s = 142;
	{8'd76,8'd67} : s = 143;
	{8'd76,8'd68} : s = 144;
	{8'd76,8'd69} : s = 145;
	{8'd76,8'd70} : s = 146;
	{8'd76,8'd71} : s = 147;
	{8'd76,8'd72} : s = 148;
	{8'd76,8'd73} : s = 149;
	{8'd76,8'd74} : s = 150;
	{8'd76,8'd75} : s = 151;
	{8'd76,8'd76} : s = 152;
	{8'd76,8'd77} : s = 153;
	{8'd76,8'd78} : s = 154;
	{8'd76,8'd79} : s = 155;
	{8'd76,8'd80} : s = 156;
	{8'd76,8'd81} : s = 157;
	{8'd76,8'd82} : s = 158;
	{8'd76,8'd83} : s = 159;
	{8'd76,8'd84} : s = 160;
	{8'd76,8'd85} : s = 161;
	{8'd76,8'd86} : s = 162;
	{8'd76,8'd87} : s = 163;
	{8'd76,8'd88} : s = 164;
	{8'd76,8'd89} : s = 165;
	{8'd76,8'd90} : s = 166;
	{8'd76,8'd91} : s = 167;
	{8'd76,8'd92} : s = 168;
	{8'd76,8'd93} : s = 169;
	{8'd76,8'd94} : s = 170;
	{8'd76,8'd95} : s = 171;
	{8'd76,8'd96} : s = 172;
	{8'd76,8'd97} : s = 173;
	{8'd76,8'd98} : s = 174;
	{8'd76,8'd99} : s = 175;
	{8'd76,8'd100} : s = 176;
	{8'd76,8'd101} : s = 177;
	{8'd76,8'd102} : s = 178;
	{8'd76,8'd103} : s = 179;
	{8'd76,8'd104} : s = 180;
	{8'd76,8'd105} : s = 181;
	{8'd76,8'd106} : s = 182;
	{8'd76,8'd107} : s = 183;
	{8'd76,8'd108} : s = 184;
	{8'd76,8'd109} : s = 185;
	{8'd76,8'd110} : s = 186;
	{8'd76,8'd111} : s = 187;
	{8'd76,8'd112} : s = 188;
	{8'd76,8'd113} : s = 189;
	{8'd76,8'd114} : s = 190;
	{8'd76,8'd115} : s = 191;
	{8'd76,8'd116} : s = 192;
	{8'd76,8'd117} : s = 193;
	{8'd76,8'd118} : s = 194;
	{8'd76,8'd119} : s = 195;
	{8'd76,8'd120} : s = 196;
	{8'd76,8'd121} : s = 197;
	{8'd76,8'd122} : s = 198;
	{8'd76,8'd123} : s = 199;
	{8'd76,8'd124} : s = 200;
	{8'd76,8'd125} : s = 201;
	{8'd76,8'd126} : s = 202;
	{8'd76,8'd127} : s = 203;
	{8'd76,8'd128} : s = 204;
	{8'd76,8'd129} : s = 205;
	{8'd76,8'd130} : s = 206;
	{8'd76,8'd131} : s = 207;
	{8'd76,8'd132} : s = 208;
	{8'd76,8'd133} : s = 209;
	{8'd76,8'd134} : s = 210;
	{8'd76,8'd135} : s = 211;
	{8'd76,8'd136} : s = 212;
	{8'd76,8'd137} : s = 213;
	{8'd76,8'd138} : s = 214;
	{8'd76,8'd139} : s = 215;
	{8'd76,8'd140} : s = 216;
	{8'd76,8'd141} : s = 217;
	{8'd76,8'd142} : s = 218;
	{8'd76,8'd143} : s = 219;
	{8'd76,8'd144} : s = 220;
	{8'd76,8'd145} : s = 221;
	{8'd76,8'd146} : s = 222;
	{8'd76,8'd147} : s = 223;
	{8'd76,8'd148} : s = 224;
	{8'd76,8'd149} : s = 225;
	{8'd76,8'd150} : s = 226;
	{8'd76,8'd151} : s = 227;
	{8'd76,8'd152} : s = 228;
	{8'd76,8'd153} : s = 229;
	{8'd76,8'd154} : s = 230;
	{8'd76,8'd155} : s = 231;
	{8'd76,8'd156} : s = 232;
	{8'd76,8'd157} : s = 233;
	{8'd76,8'd158} : s = 234;
	{8'd76,8'd159} : s = 235;
	{8'd76,8'd160} : s = 236;
	{8'd76,8'd161} : s = 237;
	{8'd76,8'd162} : s = 238;
	{8'd76,8'd163} : s = 239;
	{8'd76,8'd164} : s = 240;
	{8'd76,8'd165} : s = 241;
	{8'd76,8'd166} : s = 242;
	{8'd76,8'd167} : s = 243;
	{8'd76,8'd168} : s = 244;
	{8'd76,8'd169} : s = 245;
	{8'd76,8'd170} : s = 246;
	{8'd76,8'd171} : s = 247;
	{8'd76,8'd172} : s = 248;
	{8'd76,8'd173} : s = 249;
	{8'd76,8'd174} : s = 250;
	{8'd76,8'd175} : s = 251;
	{8'd76,8'd176} : s = 252;
	{8'd76,8'd177} : s = 253;
	{8'd76,8'd178} : s = 254;
	{8'd76,8'd179} : s = 255;
	{8'd76,8'd180} : s = 256;
	{8'd76,8'd181} : s = 257;
	{8'd76,8'd182} : s = 258;
	{8'd76,8'd183} : s = 259;
	{8'd76,8'd184} : s = 260;
	{8'd76,8'd185} : s = 261;
	{8'd76,8'd186} : s = 262;
	{8'd76,8'd187} : s = 263;
	{8'd76,8'd188} : s = 264;
	{8'd76,8'd189} : s = 265;
	{8'd76,8'd190} : s = 266;
	{8'd76,8'd191} : s = 267;
	{8'd76,8'd192} : s = 268;
	{8'd76,8'd193} : s = 269;
	{8'd76,8'd194} : s = 270;
	{8'd76,8'd195} : s = 271;
	{8'd76,8'd196} : s = 272;
	{8'd76,8'd197} : s = 273;
	{8'd76,8'd198} : s = 274;
	{8'd76,8'd199} : s = 275;
	{8'd76,8'd200} : s = 276;
	{8'd76,8'd201} : s = 277;
	{8'd76,8'd202} : s = 278;
	{8'd76,8'd203} : s = 279;
	{8'd76,8'd204} : s = 280;
	{8'd76,8'd205} : s = 281;
	{8'd76,8'd206} : s = 282;
	{8'd76,8'd207} : s = 283;
	{8'd76,8'd208} : s = 284;
	{8'd76,8'd209} : s = 285;
	{8'd76,8'd210} : s = 286;
	{8'd76,8'd211} : s = 287;
	{8'd76,8'd212} : s = 288;
	{8'd76,8'd213} : s = 289;
	{8'd76,8'd214} : s = 290;
	{8'd76,8'd215} : s = 291;
	{8'd76,8'd216} : s = 292;
	{8'd76,8'd217} : s = 293;
	{8'd76,8'd218} : s = 294;
	{8'd76,8'd219} : s = 295;
	{8'd76,8'd220} : s = 296;
	{8'd76,8'd221} : s = 297;
	{8'd76,8'd222} : s = 298;
	{8'd76,8'd223} : s = 299;
	{8'd76,8'd224} : s = 300;
	{8'd76,8'd225} : s = 301;
	{8'd76,8'd226} : s = 302;
	{8'd76,8'd227} : s = 303;
	{8'd76,8'd228} : s = 304;
	{8'd76,8'd229} : s = 305;
	{8'd76,8'd230} : s = 306;
	{8'd76,8'd231} : s = 307;
	{8'd76,8'd232} : s = 308;
	{8'd76,8'd233} : s = 309;
	{8'd76,8'd234} : s = 310;
	{8'd76,8'd235} : s = 311;
	{8'd76,8'd236} : s = 312;
	{8'd76,8'd237} : s = 313;
	{8'd76,8'd238} : s = 314;
	{8'd76,8'd239} : s = 315;
	{8'd76,8'd240} : s = 316;
	{8'd76,8'd241} : s = 317;
	{8'd76,8'd242} : s = 318;
	{8'd76,8'd243} : s = 319;
	{8'd76,8'd244} : s = 320;
	{8'd76,8'd245} : s = 321;
	{8'd76,8'd246} : s = 322;
	{8'd76,8'd247} : s = 323;
	{8'd76,8'd248} : s = 324;
	{8'd76,8'd249} : s = 325;
	{8'd76,8'd250} : s = 326;
	{8'd76,8'd251} : s = 327;
	{8'd76,8'd252} : s = 328;
	{8'd76,8'd253} : s = 329;
	{8'd76,8'd254} : s = 330;
	{8'd76,8'd255} : s = 331;
	{8'd77,8'd0} : s = 77;
	{8'd77,8'd1} : s = 78;
	{8'd77,8'd2} : s = 79;
	{8'd77,8'd3} : s = 80;
	{8'd77,8'd4} : s = 81;
	{8'd77,8'd5} : s = 82;
	{8'd77,8'd6} : s = 83;
	{8'd77,8'd7} : s = 84;
	{8'd77,8'd8} : s = 85;
	{8'd77,8'd9} : s = 86;
	{8'd77,8'd10} : s = 87;
	{8'd77,8'd11} : s = 88;
	{8'd77,8'd12} : s = 89;
	{8'd77,8'd13} : s = 90;
	{8'd77,8'd14} : s = 91;
	{8'd77,8'd15} : s = 92;
	{8'd77,8'd16} : s = 93;
	{8'd77,8'd17} : s = 94;
	{8'd77,8'd18} : s = 95;
	{8'd77,8'd19} : s = 96;
	{8'd77,8'd20} : s = 97;
	{8'd77,8'd21} : s = 98;
	{8'd77,8'd22} : s = 99;
	{8'd77,8'd23} : s = 100;
	{8'd77,8'd24} : s = 101;
	{8'd77,8'd25} : s = 102;
	{8'd77,8'd26} : s = 103;
	{8'd77,8'd27} : s = 104;
	{8'd77,8'd28} : s = 105;
	{8'd77,8'd29} : s = 106;
	{8'd77,8'd30} : s = 107;
	{8'd77,8'd31} : s = 108;
	{8'd77,8'd32} : s = 109;
	{8'd77,8'd33} : s = 110;
	{8'd77,8'd34} : s = 111;
	{8'd77,8'd35} : s = 112;
	{8'd77,8'd36} : s = 113;
	{8'd77,8'd37} : s = 114;
	{8'd77,8'd38} : s = 115;
	{8'd77,8'd39} : s = 116;
	{8'd77,8'd40} : s = 117;
	{8'd77,8'd41} : s = 118;
	{8'd77,8'd42} : s = 119;
	{8'd77,8'd43} : s = 120;
	{8'd77,8'd44} : s = 121;
	{8'd77,8'd45} : s = 122;
	{8'd77,8'd46} : s = 123;
	{8'd77,8'd47} : s = 124;
	{8'd77,8'd48} : s = 125;
	{8'd77,8'd49} : s = 126;
	{8'd77,8'd50} : s = 127;
	{8'd77,8'd51} : s = 128;
	{8'd77,8'd52} : s = 129;
	{8'd77,8'd53} : s = 130;
	{8'd77,8'd54} : s = 131;
	{8'd77,8'd55} : s = 132;
	{8'd77,8'd56} : s = 133;
	{8'd77,8'd57} : s = 134;
	{8'd77,8'd58} : s = 135;
	{8'd77,8'd59} : s = 136;
	{8'd77,8'd60} : s = 137;
	{8'd77,8'd61} : s = 138;
	{8'd77,8'd62} : s = 139;
	{8'd77,8'd63} : s = 140;
	{8'd77,8'd64} : s = 141;
	{8'd77,8'd65} : s = 142;
	{8'd77,8'd66} : s = 143;
	{8'd77,8'd67} : s = 144;
	{8'd77,8'd68} : s = 145;
	{8'd77,8'd69} : s = 146;
	{8'd77,8'd70} : s = 147;
	{8'd77,8'd71} : s = 148;
	{8'd77,8'd72} : s = 149;
	{8'd77,8'd73} : s = 150;
	{8'd77,8'd74} : s = 151;
	{8'd77,8'd75} : s = 152;
	{8'd77,8'd76} : s = 153;
	{8'd77,8'd77} : s = 154;
	{8'd77,8'd78} : s = 155;
	{8'd77,8'd79} : s = 156;
	{8'd77,8'd80} : s = 157;
	{8'd77,8'd81} : s = 158;
	{8'd77,8'd82} : s = 159;
	{8'd77,8'd83} : s = 160;
	{8'd77,8'd84} : s = 161;
	{8'd77,8'd85} : s = 162;
	{8'd77,8'd86} : s = 163;
	{8'd77,8'd87} : s = 164;
	{8'd77,8'd88} : s = 165;
	{8'd77,8'd89} : s = 166;
	{8'd77,8'd90} : s = 167;
	{8'd77,8'd91} : s = 168;
	{8'd77,8'd92} : s = 169;
	{8'd77,8'd93} : s = 170;
	{8'd77,8'd94} : s = 171;
	{8'd77,8'd95} : s = 172;
	{8'd77,8'd96} : s = 173;
	{8'd77,8'd97} : s = 174;
	{8'd77,8'd98} : s = 175;
	{8'd77,8'd99} : s = 176;
	{8'd77,8'd100} : s = 177;
	{8'd77,8'd101} : s = 178;
	{8'd77,8'd102} : s = 179;
	{8'd77,8'd103} : s = 180;
	{8'd77,8'd104} : s = 181;
	{8'd77,8'd105} : s = 182;
	{8'd77,8'd106} : s = 183;
	{8'd77,8'd107} : s = 184;
	{8'd77,8'd108} : s = 185;
	{8'd77,8'd109} : s = 186;
	{8'd77,8'd110} : s = 187;
	{8'd77,8'd111} : s = 188;
	{8'd77,8'd112} : s = 189;
	{8'd77,8'd113} : s = 190;
	{8'd77,8'd114} : s = 191;
	{8'd77,8'd115} : s = 192;
	{8'd77,8'd116} : s = 193;
	{8'd77,8'd117} : s = 194;
	{8'd77,8'd118} : s = 195;
	{8'd77,8'd119} : s = 196;
	{8'd77,8'd120} : s = 197;
	{8'd77,8'd121} : s = 198;
	{8'd77,8'd122} : s = 199;
	{8'd77,8'd123} : s = 200;
	{8'd77,8'd124} : s = 201;
	{8'd77,8'd125} : s = 202;
	{8'd77,8'd126} : s = 203;
	{8'd77,8'd127} : s = 204;
	{8'd77,8'd128} : s = 205;
	{8'd77,8'd129} : s = 206;
	{8'd77,8'd130} : s = 207;
	{8'd77,8'd131} : s = 208;
	{8'd77,8'd132} : s = 209;
	{8'd77,8'd133} : s = 210;
	{8'd77,8'd134} : s = 211;
	{8'd77,8'd135} : s = 212;
	{8'd77,8'd136} : s = 213;
	{8'd77,8'd137} : s = 214;
	{8'd77,8'd138} : s = 215;
	{8'd77,8'd139} : s = 216;
	{8'd77,8'd140} : s = 217;
	{8'd77,8'd141} : s = 218;
	{8'd77,8'd142} : s = 219;
	{8'd77,8'd143} : s = 220;
	{8'd77,8'd144} : s = 221;
	{8'd77,8'd145} : s = 222;
	{8'd77,8'd146} : s = 223;
	{8'd77,8'd147} : s = 224;
	{8'd77,8'd148} : s = 225;
	{8'd77,8'd149} : s = 226;
	{8'd77,8'd150} : s = 227;
	{8'd77,8'd151} : s = 228;
	{8'd77,8'd152} : s = 229;
	{8'd77,8'd153} : s = 230;
	{8'd77,8'd154} : s = 231;
	{8'd77,8'd155} : s = 232;
	{8'd77,8'd156} : s = 233;
	{8'd77,8'd157} : s = 234;
	{8'd77,8'd158} : s = 235;
	{8'd77,8'd159} : s = 236;
	{8'd77,8'd160} : s = 237;
	{8'd77,8'd161} : s = 238;
	{8'd77,8'd162} : s = 239;
	{8'd77,8'd163} : s = 240;
	{8'd77,8'd164} : s = 241;
	{8'd77,8'd165} : s = 242;
	{8'd77,8'd166} : s = 243;
	{8'd77,8'd167} : s = 244;
	{8'd77,8'd168} : s = 245;
	{8'd77,8'd169} : s = 246;
	{8'd77,8'd170} : s = 247;
	{8'd77,8'd171} : s = 248;
	{8'd77,8'd172} : s = 249;
	{8'd77,8'd173} : s = 250;
	{8'd77,8'd174} : s = 251;
	{8'd77,8'd175} : s = 252;
	{8'd77,8'd176} : s = 253;
	{8'd77,8'd177} : s = 254;
	{8'd77,8'd178} : s = 255;
	{8'd77,8'd179} : s = 256;
	{8'd77,8'd180} : s = 257;
	{8'd77,8'd181} : s = 258;
	{8'd77,8'd182} : s = 259;
	{8'd77,8'd183} : s = 260;
	{8'd77,8'd184} : s = 261;
	{8'd77,8'd185} : s = 262;
	{8'd77,8'd186} : s = 263;
	{8'd77,8'd187} : s = 264;
	{8'd77,8'd188} : s = 265;
	{8'd77,8'd189} : s = 266;
	{8'd77,8'd190} : s = 267;
	{8'd77,8'd191} : s = 268;
	{8'd77,8'd192} : s = 269;
	{8'd77,8'd193} : s = 270;
	{8'd77,8'd194} : s = 271;
	{8'd77,8'd195} : s = 272;
	{8'd77,8'd196} : s = 273;
	{8'd77,8'd197} : s = 274;
	{8'd77,8'd198} : s = 275;
	{8'd77,8'd199} : s = 276;
	{8'd77,8'd200} : s = 277;
	{8'd77,8'd201} : s = 278;
	{8'd77,8'd202} : s = 279;
	{8'd77,8'd203} : s = 280;
	{8'd77,8'd204} : s = 281;
	{8'd77,8'd205} : s = 282;
	{8'd77,8'd206} : s = 283;
	{8'd77,8'd207} : s = 284;
	{8'd77,8'd208} : s = 285;
	{8'd77,8'd209} : s = 286;
	{8'd77,8'd210} : s = 287;
	{8'd77,8'd211} : s = 288;
	{8'd77,8'd212} : s = 289;
	{8'd77,8'd213} : s = 290;
	{8'd77,8'd214} : s = 291;
	{8'd77,8'd215} : s = 292;
	{8'd77,8'd216} : s = 293;
	{8'd77,8'd217} : s = 294;
	{8'd77,8'd218} : s = 295;
	{8'd77,8'd219} : s = 296;
	{8'd77,8'd220} : s = 297;
	{8'd77,8'd221} : s = 298;
	{8'd77,8'd222} : s = 299;
	{8'd77,8'd223} : s = 300;
	{8'd77,8'd224} : s = 301;
	{8'd77,8'd225} : s = 302;
	{8'd77,8'd226} : s = 303;
	{8'd77,8'd227} : s = 304;
	{8'd77,8'd228} : s = 305;
	{8'd77,8'd229} : s = 306;
	{8'd77,8'd230} : s = 307;
	{8'd77,8'd231} : s = 308;
	{8'd77,8'd232} : s = 309;
	{8'd77,8'd233} : s = 310;
	{8'd77,8'd234} : s = 311;
	{8'd77,8'd235} : s = 312;
	{8'd77,8'd236} : s = 313;
	{8'd77,8'd237} : s = 314;
	{8'd77,8'd238} : s = 315;
	{8'd77,8'd239} : s = 316;
	{8'd77,8'd240} : s = 317;
	{8'd77,8'd241} : s = 318;
	{8'd77,8'd242} : s = 319;
	{8'd77,8'd243} : s = 320;
	{8'd77,8'd244} : s = 321;
	{8'd77,8'd245} : s = 322;
	{8'd77,8'd246} : s = 323;
	{8'd77,8'd247} : s = 324;
	{8'd77,8'd248} : s = 325;
	{8'd77,8'd249} : s = 326;
	{8'd77,8'd250} : s = 327;
	{8'd77,8'd251} : s = 328;
	{8'd77,8'd252} : s = 329;
	{8'd77,8'd253} : s = 330;
	{8'd77,8'd254} : s = 331;
	{8'd77,8'd255} : s = 332;
	{8'd78,8'd0} : s = 78;
	{8'd78,8'd1} : s = 79;
	{8'd78,8'd2} : s = 80;
	{8'd78,8'd3} : s = 81;
	{8'd78,8'd4} : s = 82;
	{8'd78,8'd5} : s = 83;
	{8'd78,8'd6} : s = 84;
	{8'd78,8'd7} : s = 85;
	{8'd78,8'd8} : s = 86;
	{8'd78,8'd9} : s = 87;
	{8'd78,8'd10} : s = 88;
	{8'd78,8'd11} : s = 89;
	{8'd78,8'd12} : s = 90;
	{8'd78,8'd13} : s = 91;
	{8'd78,8'd14} : s = 92;
	{8'd78,8'd15} : s = 93;
	{8'd78,8'd16} : s = 94;
	{8'd78,8'd17} : s = 95;
	{8'd78,8'd18} : s = 96;
	{8'd78,8'd19} : s = 97;
	{8'd78,8'd20} : s = 98;
	{8'd78,8'd21} : s = 99;
	{8'd78,8'd22} : s = 100;
	{8'd78,8'd23} : s = 101;
	{8'd78,8'd24} : s = 102;
	{8'd78,8'd25} : s = 103;
	{8'd78,8'd26} : s = 104;
	{8'd78,8'd27} : s = 105;
	{8'd78,8'd28} : s = 106;
	{8'd78,8'd29} : s = 107;
	{8'd78,8'd30} : s = 108;
	{8'd78,8'd31} : s = 109;
	{8'd78,8'd32} : s = 110;
	{8'd78,8'd33} : s = 111;
	{8'd78,8'd34} : s = 112;
	{8'd78,8'd35} : s = 113;
	{8'd78,8'd36} : s = 114;
	{8'd78,8'd37} : s = 115;
	{8'd78,8'd38} : s = 116;
	{8'd78,8'd39} : s = 117;
	{8'd78,8'd40} : s = 118;
	{8'd78,8'd41} : s = 119;
	{8'd78,8'd42} : s = 120;
	{8'd78,8'd43} : s = 121;
	{8'd78,8'd44} : s = 122;
	{8'd78,8'd45} : s = 123;
	{8'd78,8'd46} : s = 124;
	{8'd78,8'd47} : s = 125;
	{8'd78,8'd48} : s = 126;
	{8'd78,8'd49} : s = 127;
	{8'd78,8'd50} : s = 128;
	{8'd78,8'd51} : s = 129;
	{8'd78,8'd52} : s = 130;
	{8'd78,8'd53} : s = 131;
	{8'd78,8'd54} : s = 132;
	{8'd78,8'd55} : s = 133;
	{8'd78,8'd56} : s = 134;
	{8'd78,8'd57} : s = 135;
	{8'd78,8'd58} : s = 136;
	{8'd78,8'd59} : s = 137;
	{8'd78,8'd60} : s = 138;
	{8'd78,8'd61} : s = 139;
	{8'd78,8'd62} : s = 140;
	{8'd78,8'd63} : s = 141;
	{8'd78,8'd64} : s = 142;
	{8'd78,8'd65} : s = 143;
	{8'd78,8'd66} : s = 144;
	{8'd78,8'd67} : s = 145;
	{8'd78,8'd68} : s = 146;
	{8'd78,8'd69} : s = 147;
	{8'd78,8'd70} : s = 148;
	{8'd78,8'd71} : s = 149;
	{8'd78,8'd72} : s = 150;
	{8'd78,8'd73} : s = 151;
	{8'd78,8'd74} : s = 152;
	{8'd78,8'd75} : s = 153;
	{8'd78,8'd76} : s = 154;
	{8'd78,8'd77} : s = 155;
	{8'd78,8'd78} : s = 156;
	{8'd78,8'd79} : s = 157;
	{8'd78,8'd80} : s = 158;
	{8'd78,8'd81} : s = 159;
	{8'd78,8'd82} : s = 160;
	{8'd78,8'd83} : s = 161;
	{8'd78,8'd84} : s = 162;
	{8'd78,8'd85} : s = 163;
	{8'd78,8'd86} : s = 164;
	{8'd78,8'd87} : s = 165;
	{8'd78,8'd88} : s = 166;
	{8'd78,8'd89} : s = 167;
	{8'd78,8'd90} : s = 168;
	{8'd78,8'd91} : s = 169;
	{8'd78,8'd92} : s = 170;
	{8'd78,8'd93} : s = 171;
	{8'd78,8'd94} : s = 172;
	{8'd78,8'd95} : s = 173;
	{8'd78,8'd96} : s = 174;
	{8'd78,8'd97} : s = 175;
	{8'd78,8'd98} : s = 176;
	{8'd78,8'd99} : s = 177;
	{8'd78,8'd100} : s = 178;
	{8'd78,8'd101} : s = 179;
	{8'd78,8'd102} : s = 180;
	{8'd78,8'd103} : s = 181;
	{8'd78,8'd104} : s = 182;
	{8'd78,8'd105} : s = 183;
	{8'd78,8'd106} : s = 184;
	{8'd78,8'd107} : s = 185;
	{8'd78,8'd108} : s = 186;
	{8'd78,8'd109} : s = 187;
	{8'd78,8'd110} : s = 188;
	{8'd78,8'd111} : s = 189;
	{8'd78,8'd112} : s = 190;
	{8'd78,8'd113} : s = 191;
	{8'd78,8'd114} : s = 192;
	{8'd78,8'd115} : s = 193;
	{8'd78,8'd116} : s = 194;
	{8'd78,8'd117} : s = 195;
	{8'd78,8'd118} : s = 196;
	{8'd78,8'd119} : s = 197;
	{8'd78,8'd120} : s = 198;
	{8'd78,8'd121} : s = 199;
	{8'd78,8'd122} : s = 200;
	{8'd78,8'd123} : s = 201;
	{8'd78,8'd124} : s = 202;
	{8'd78,8'd125} : s = 203;
	{8'd78,8'd126} : s = 204;
	{8'd78,8'd127} : s = 205;
	{8'd78,8'd128} : s = 206;
	{8'd78,8'd129} : s = 207;
	{8'd78,8'd130} : s = 208;
	{8'd78,8'd131} : s = 209;
	{8'd78,8'd132} : s = 210;
	{8'd78,8'd133} : s = 211;
	{8'd78,8'd134} : s = 212;
	{8'd78,8'd135} : s = 213;
	{8'd78,8'd136} : s = 214;
	{8'd78,8'd137} : s = 215;
	{8'd78,8'd138} : s = 216;
	{8'd78,8'd139} : s = 217;
	{8'd78,8'd140} : s = 218;
	{8'd78,8'd141} : s = 219;
	{8'd78,8'd142} : s = 220;
	{8'd78,8'd143} : s = 221;
	{8'd78,8'd144} : s = 222;
	{8'd78,8'd145} : s = 223;
	{8'd78,8'd146} : s = 224;
	{8'd78,8'd147} : s = 225;
	{8'd78,8'd148} : s = 226;
	{8'd78,8'd149} : s = 227;
	{8'd78,8'd150} : s = 228;
	{8'd78,8'd151} : s = 229;
	{8'd78,8'd152} : s = 230;
	{8'd78,8'd153} : s = 231;
	{8'd78,8'd154} : s = 232;
	{8'd78,8'd155} : s = 233;
	{8'd78,8'd156} : s = 234;
	{8'd78,8'd157} : s = 235;
	{8'd78,8'd158} : s = 236;
	{8'd78,8'd159} : s = 237;
	{8'd78,8'd160} : s = 238;
	{8'd78,8'd161} : s = 239;
	{8'd78,8'd162} : s = 240;
	{8'd78,8'd163} : s = 241;
	{8'd78,8'd164} : s = 242;
	{8'd78,8'd165} : s = 243;
	{8'd78,8'd166} : s = 244;
	{8'd78,8'd167} : s = 245;
	{8'd78,8'd168} : s = 246;
	{8'd78,8'd169} : s = 247;
	{8'd78,8'd170} : s = 248;
	{8'd78,8'd171} : s = 249;
	{8'd78,8'd172} : s = 250;
	{8'd78,8'd173} : s = 251;
	{8'd78,8'd174} : s = 252;
	{8'd78,8'd175} : s = 253;
	{8'd78,8'd176} : s = 254;
	{8'd78,8'd177} : s = 255;
	{8'd78,8'd178} : s = 256;
	{8'd78,8'd179} : s = 257;
	{8'd78,8'd180} : s = 258;
	{8'd78,8'd181} : s = 259;
	{8'd78,8'd182} : s = 260;
	{8'd78,8'd183} : s = 261;
	{8'd78,8'd184} : s = 262;
	{8'd78,8'd185} : s = 263;
	{8'd78,8'd186} : s = 264;
	{8'd78,8'd187} : s = 265;
	{8'd78,8'd188} : s = 266;
	{8'd78,8'd189} : s = 267;
	{8'd78,8'd190} : s = 268;
	{8'd78,8'd191} : s = 269;
	{8'd78,8'd192} : s = 270;
	{8'd78,8'd193} : s = 271;
	{8'd78,8'd194} : s = 272;
	{8'd78,8'd195} : s = 273;
	{8'd78,8'd196} : s = 274;
	{8'd78,8'd197} : s = 275;
	{8'd78,8'd198} : s = 276;
	{8'd78,8'd199} : s = 277;
	{8'd78,8'd200} : s = 278;
	{8'd78,8'd201} : s = 279;
	{8'd78,8'd202} : s = 280;
	{8'd78,8'd203} : s = 281;
	{8'd78,8'd204} : s = 282;
	{8'd78,8'd205} : s = 283;
	{8'd78,8'd206} : s = 284;
	{8'd78,8'd207} : s = 285;
	{8'd78,8'd208} : s = 286;
	{8'd78,8'd209} : s = 287;
	{8'd78,8'd210} : s = 288;
	{8'd78,8'd211} : s = 289;
	{8'd78,8'd212} : s = 290;
	{8'd78,8'd213} : s = 291;
	{8'd78,8'd214} : s = 292;
	{8'd78,8'd215} : s = 293;
	{8'd78,8'd216} : s = 294;
	{8'd78,8'd217} : s = 295;
	{8'd78,8'd218} : s = 296;
	{8'd78,8'd219} : s = 297;
	{8'd78,8'd220} : s = 298;
	{8'd78,8'd221} : s = 299;
	{8'd78,8'd222} : s = 300;
	{8'd78,8'd223} : s = 301;
	{8'd78,8'd224} : s = 302;
	{8'd78,8'd225} : s = 303;
	{8'd78,8'd226} : s = 304;
	{8'd78,8'd227} : s = 305;
	{8'd78,8'd228} : s = 306;
	{8'd78,8'd229} : s = 307;
	{8'd78,8'd230} : s = 308;
	{8'd78,8'd231} : s = 309;
	{8'd78,8'd232} : s = 310;
	{8'd78,8'd233} : s = 311;
	{8'd78,8'd234} : s = 312;
	{8'd78,8'd235} : s = 313;
	{8'd78,8'd236} : s = 314;
	{8'd78,8'd237} : s = 315;
	{8'd78,8'd238} : s = 316;
	{8'd78,8'd239} : s = 317;
	{8'd78,8'd240} : s = 318;
	{8'd78,8'd241} : s = 319;
	{8'd78,8'd242} : s = 320;
	{8'd78,8'd243} : s = 321;
	{8'd78,8'd244} : s = 322;
	{8'd78,8'd245} : s = 323;
	{8'd78,8'd246} : s = 324;
	{8'd78,8'd247} : s = 325;
	{8'd78,8'd248} : s = 326;
	{8'd78,8'd249} : s = 327;
	{8'd78,8'd250} : s = 328;
	{8'd78,8'd251} : s = 329;
	{8'd78,8'd252} : s = 330;
	{8'd78,8'd253} : s = 331;
	{8'd78,8'd254} : s = 332;
	{8'd78,8'd255} : s = 333;
	{8'd79,8'd0} : s = 79;
	{8'd79,8'd1} : s = 80;
	{8'd79,8'd2} : s = 81;
	{8'd79,8'd3} : s = 82;
	{8'd79,8'd4} : s = 83;
	{8'd79,8'd5} : s = 84;
	{8'd79,8'd6} : s = 85;
	{8'd79,8'd7} : s = 86;
	{8'd79,8'd8} : s = 87;
	{8'd79,8'd9} : s = 88;
	{8'd79,8'd10} : s = 89;
	{8'd79,8'd11} : s = 90;
	{8'd79,8'd12} : s = 91;
	{8'd79,8'd13} : s = 92;
	{8'd79,8'd14} : s = 93;
	{8'd79,8'd15} : s = 94;
	{8'd79,8'd16} : s = 95;
	{8'd79,8'd17} : s = 96;
	{8'd79,8'd18} : s = 97;
	{8'd79,8'd19} : s = 98;
	{8'd79,8'd20} : s = 99;
	{8'd79,8'd21} : s = 100;
	{8'd79,8'd22} : s = 101;
	{8'd79,8'd23} : s = 102;
	{8'd79,8'd24} : s = 103;
	{8'd79,8'd25} : s = 104;
	{8'd79,8'd26} : s = 105;
	{8'd79,8'd27} : s = 106;
	{8'd79,8'd28} : s = 107;
	{8'd79,8'd29} : s = 108;
	{8'd79,8'd30} : s = 109;
	{8'd79,8'd31} : s = 110;
	{8'd79,8'd32} : s = 111;
	{8'd79,8'd33} : s = 112;
	{8'd79,8'd34} : s = 113;
	{8'd79,8'd35} : s = 114;
	{8'd79,8'd36} : s = 115;
	{8'd79,8'd37} : s = 116;
	{8'd79,8'd38} : s = 117;
	{8'd79,8'd39} : s = 118;
	{8'd79,8'd40} : s = 119;
	{8'd79,8'd41} : s = 120;
	{8'd79,8'd42} : s = 121;
	{8'd79,8'd43} : s = 122;
	{8'd79,8'd44} : s = 123;
	{8'd79,8'd45} : s = 124;
	{8'd79,8'd46} : s = 125;
	{8'd79,8'd47} : s = 126;
	{8'd79,8'd48} : s = 127;
	{8'd79,8'd49} : s = 128;
	{8'd79,8'd50} : s = 129;
	{8'd79,8'd51} : s = 130;
	{8'd79,8'd52} : s = 131;
	{8'd79,8'd53} : s = 132;
	{8'd79,8'd54} : s = 133;
	{8'd79,8'd55} : s = 134;
	{8'd79,8'd56} : s = 135;
	{8'd79,8'd57} : s = 136;
	{8'd79,8'd58} : s = 137;
	{8'd79,8'd59} : s = 138;
	{8'd79,8'd60} : s = 139;
	{8'd79,8'd61} : s = 140;
	{8'd79,8'd62} : s = 141;
	{8'd79,8'd63} : s = 142;
	{8'd79,8'd64} : s = 143;
	{8'd79,8'd65} : s = 144;
	{8'd79,8'd66} : s = 145;
	{8'd79,8'd67} : s = 146;
	{8'd79,8'd68} : s = 147;
	{8'd79,8'd69} : s = 148;
	{8'd79,8'd70} : s = 149;
	{8'd79,8'd71} : s = 150;
	{8'd79,8'd72} : s = 151;
	{8'd79,8'd73} : s = 152;
	{8'd79,8'd74} : s = 153;
	{8'd79,8'd75} : s = 154;
	{8'd79,8'd76} : s = 155;
	{8'd79,8'd77} : s = 156;
	{8'd79,8'd78} : s = 157;
	{8'd79,8'd79} : s = 158;
	{8'd79,8'd80} : s = 159;
	{8'd79,8'd81} : s = 160;
	{8'd79,8'd82} : s = 161;
	{8'd79,8'd83} : s = 162;
	{8'd79,8'd84} : s = 163;
	{8'd79,8'd85} : s = 164;
	{8'd79,8'd86} : s = 165;
	{8'd79,8'd87} : s = 166;
	{8'd79,8'd88} : s = 167;
	{8'd79,8'd89} : s = 168;
	{8'd79,8'd90} : s = 169;
	{8'd79,8'd91} : s = 170;
	{8'd79,8'd92} : s = 171;
	{8'd79,8'd93} : s = 172;
	{8'd79,8'd94} : s = 173;
	{8'd79,8'd95} : s = 174;
	{8'd79,8'd96} : s = 175;
	{8'd79,8'd97} : s = 176;
	{8'd79,8'd98} : s = 177;
	{8'd79,8'd99} : s = 178;
	{8'd79,8'd100} : s = 179;
	{8'd79,8'd101} : s = 180;
	{8'd79,8'd102} : s = 181;
	{8'd79,8'd103} : s = 182;
	{8'd79,8'd104} : s = 183;
	{8'd79,8'd105} : s = 184;
	{8'd79,8'd106} : s = 185;
	{8'd79,8'd107} : s = 186;
	{8'd79,8'd108} : s = 187;
	{8'd79,8'd109} : s = 188;
	{8'd79,8'd110} : s = 189;
	{8'd79,8'd111} : s = 190;
	{8'd79,8'd112} : s = 191;
	{8'd79,8'd113} : s = 192;
	{8'd79,8'd114} : s = 193;
	{8'd79,8'd115} : s = 194;
	{8'd79,8'd116} : s = 195;
	{8'd79,8'd117} : s = 196;
	{8'd79,8'd118} : s = 197;
	{8'd79,8'd119} : s = 198;
	{8'd79,8'd120} : s = 199;
	{8'd79,8'd121} : s = 200;
	{8'd79,8'd122} : s = 201;
	{8'd79,8'd123} : s = 202;
	{8'd79,8'd124} : s = 203;
	{8'd79,8'd125} : s = 204;
	{8'd79,8'd126} : s = 205;
	{8'd79,8'd127} : s = 206;
	{8'd79,8'd128} : s = 207;
	{8'd79,8'd129} : s = 208;
	{8'd79,8'd130} : s = 209;
	{8'd79,8'd131} : s = 210;
	{8'd79,8'd132} : s = 211;
	{8'd79,8'd133} : s = 212;
	{8'd79,8'd134} : s = 213;
	{8'd79,8'd135} : s = 214;
	{8'd79,8'd136} : s = 215;
	{8'd79,8'd137} : s = 216;
	{8'd79,8'd138} : s = 217;
	{8'd79,8'd139} : s = 218;
	{8'd79,8'd140} : s = 219;
	{8'd79,8'd141} : s = 220;
	{8'd79,8'd142} : s = 221;
	{8'd79,8'd143} : s = 222;
	{8'd79,8'd144} : s = 223;
	{8'd79,8'd145} : s = 224;
	{8'd79,8'd146} : s = 225;
	{8'd79,8'd147} : s = 226;
	{8'd79,8'd148} : s = 227;
	{8'd79,8'd149} : s = 228;
	{8'd79,8'd150} : s = 229;
	{8'd79,8'd151} : s = 230;
	{8'd79,8'd152} : s = 231;
	{8'd79,8'd153} : s = 232;
	{8'd79,8'd154} : s = 233;
	{8'd79,8'd155} : s = 234;
	{8'd79,8'd156} : s = 235;
	{8'd79,8'd157} : s = 236;
	{8'd79,8'd158} : s = 237;
	{8'd79,8'd159} : s = 238;
	{8'd79,8'd160} : s = 239;
	{8'd79,8'd161} : s = 240;
	{8'd79,8'd162} : s = 241;
	{8'd79,8'd163} : s = 242;
	{8'd79,8'd164} : s = 243;
	{8'd79,8'd165} : s = 244;
	{8'd79,8'd166} : s = 245;
	{8'd79,8'd167} : s = 246;
	{8'd79,8'd168} : s = 247;
	{8'd79,8'd169} : s = 248;
	{8'd79,8'd170} : s = 249;
	{8'd79,8'd171} : s = 250;
	{8'd79,8'd172} : s = 251;
	{8'd79,8'd173} : s = 252;
	{8'd79,8'd174} : s = 253;
	{8'd79,8'd175} : s = 254;
	{8'd79,8'd176} : s = 255;
	{8'd79,8'd177} : s = 256;
	{8'd79,8'd178} : s = 257;
	{8'd79,8'd179} : s = 258;
	{8'd79,8'd180} : s = 259;
	{8'd79,8'd181} : s = 260;
	{8'd79,8'd182} : s = 261;
	{8'd79,8'd183} : s = 262;
	{8'd79,8'd184} : s = 263;
	{8'd79,8'd185} : s = 264;
	{8'd79,8'd186} : s = 265;
	{8'd79,8'd187} : s = 266;
	{8'd79,8'd188} : s = 267;
	{8'd79,8'd189} : s = 268;
	{8'd79,8'd190} : s = 269;
	{8'd79,8'd191} : s = 270;
	{8'd79,8'd192} : s = 271;
	{8'd79,8'd193} : s = 272;
	{8'd79,8'd194} : s = 273;
	{8'd79,8'd195} : s = 274;
	{8'd79,8'd196} : s = 275;
	{8'd79,8'd197} : s = 276;
	{8'd79,8'd198} : s = 277;
	{8'd79,8'd199} : s = 278;
	{8'd79,8'd200} : s = 279;
	{8'd79,8'd201} : s = 280;
	{8'd79,8'd202} : s = 281;
	{8'd79,8'd203} : s = 282;
	{8'd79,8'd204} : s = 283;
	{8'd79,8'd205} : s = 284;
	{8'd79,8'd206} : s = 285;
	{8'd79,8'd207} : s = 286;
	{8'd79,8'd208} : s = 287;
	{8'd79,8'd209} : s = 288;
	{8'd79,8'd210} : s = 289;
	{8'd79,8'd211} : s = 290;
	{8'd79,8'd212} : s = 291;
	{8'd79,8'd213} : s = 292;
	{8'd79,8'd214} : s = 293;
	{8'd79,8'd215} : s = 294;
	{8'd79,8'd216} : s = 295;
	{8'd79,8'd217} : s = 296;
	{8'd79,8'd218} : s = 297;
	{8'd79,8'd219} : s = 298;
	{8'd79,8'd220} : s = 299;
	{8'd79,8'd221} : s = 300;
	{8'd79,8'd222} : s = 301;
	{8'd79,8'd223} : s = 302;
	{8'd79,8'd224} : s = 303;
	{8'd79,8'd225} : s = 304;
	{8'd79,8'd226} : s = 305;
	{8'd79,8'd227} : s = 306;
	{8'd79,8'd228} : s = 307;
	{8'd79,8'd229} : s = 308;
	{8'd79,8'd230} : s = 309;
	{8'd79,8'd231} : s = 310;
	{8'd79,8'd232} : s = 311;
	{8'd79,8'd233} : s = 312;
	{8'd79,8'd234} : s = 313;
	{8'd79,8'd235} : s = 314;
	{8'd79,8'd236} : s = 315;
	{8'd79,8'd237} : s = 316;
	{8'd79,8'd238} : s = 317;
	{8'd79,8'd239} : s = 318;
	{8'd79,8'd240} : s = 319;
	{8'd79,8'd241} : s = 320;
	{8'd79,8'd242} : s = 321;
	{8'd79,8'd243} : s = 322;
	{8'd79,8'd244} : s = 323;
	{8'd79,8'd245} : s = 324;
	{8'd79,8'd246} : s = 325;
	{8'd79,8'd247} : s = 326;
	{8'd79,8'd248} : s = 327;
	{8'd79,8'd249} : s = 328;
	{8'd79,8'd250} : s = 329;
	{8'd79,8'd251} : s = 330;
	{8'd79,8'd252} : s = 331;
	{8'd79,8'd253} : s = 332;
	{8'd79,8'd254} : s = 333;
	{8'd79,8'd255} : s = 334;
	{8'd80,8'd0} : s = 80;
	{8'd80,8'd1} : s = 81;
	{8'd80,8'd2} : s = 82;
	{8'd80,8'd3} : s = 83;
	{8'd80,8'd4} : s = 84;
	{8'd80,8'd5} : s = 85;
	{8'd80,8'd6} : s = 86;
	{8'd80,8'd7} : s = 87;
	{8'd80,8'd8} : s = 88;
	{8'd80,8'd9} : s = 89;
	{8'd80,8'd10} : s = 90;
	{8'd80,8'd11} : s = 91;
	{8'd80,8'd12} : s = 92;
	{8'd80,8'd13} : s = 93;
	{8'd80,8'd14} : s = 94;
	{8'd80,8'd15} : s = 95;
	{8'd80,8'd16} : s = 96;
	{8'd80,8'd17} : s = 97;
	{8'd80,8'd18} : s = 98;
	{8'd80,8'd19} : s = 99;
	{8'd80,8'd20} : s = 100;
	{8'd80,8'd21} : s = 101;
	{8'd80,8'd22} : s = 102;
	{8'd80,8'd23} : s = 103;
	{8'd80,8'd24} : s = 104;
	{8'd80,8'd25} : s = 105;
	{8'd80,8'd26} : s = 106;
	{8'd80,8'd27} : s = 107;
	{8'd80,8'd28} : s = 108;
	{8'd80,8'd29} : s = 109;
	{8'd80,8'd30} : s = 110;
	{8'd80,8'd31} : s = 111;
	{8'd80,8'd32} : s = 112;
	{8'd80,8'd33} : s = 113;
	{8'd80,8'd34} : s = 114;
	{8'd80,8'd35} : s = 115;
	{8'd80,8'd36} : s = 116;
	{8'd80,8'd37} : s = 117;
	{8'd80,8'd38} : s = 118;
	{8'd80,8'd39} : s = 119;
	{8'd80,8'd40} : s = 120;
	{8'd80,8'd41} : s = 121;
	{8'd80,8'd42} : s = 122;
	{8'd80,8'd43} : s = 123;
	{8'd80,8'd44} : s = 124;
	{8'd80,8'd45} : s = 125;
	{8'd80,8'd46} : s = 126;
	{8'd80,8'd47} : s = 127;
	{8'd80,8'd48} : s = 128;
	{8'd80,8'd49} : s = 129;
	{8'd80,8'd50} : s = 130;
	{8'd80,8'd51} : s = 131;
	{8'd80,8'd52} : s = 132;
	{8'd80,8'd53} : s = 133;
	{8'd80,8'd54} : s = 134;
	{8'd80,8'd55} : s = 135;
	{8'd80,8'd56} : s = 136;
	{8'd80,8'd57} : s = 137;
	{8'd80,8'd58} : s = 138;
	{8'd80,8'd59} : s = 139;
	{8'd80,8'd60} : s = 140;
	{8'd80,8'd61} : s = 141;
	{8'd80,8'd62} : s = 142;
	{8'd80,8'd63} : s = 143;
	{8'd80,8'd64} : s = 144;
	{8'd80,8'd65} : s = 145;
	{8'd80,8'd66} : s = 146;
	{8'd80,8'd67} : s = 147;
	{8'd80,8'd68} : s = 148;
	{8'd80,8'd69} : s = 149;
	{8'd80,8'd70} : s = 150;
	{8'd80,8'd71} : s = 151;
	{8'd80,8'd72} : s = 152;
	{8'd80,8'd73} : s = 153;
	{8'd80,8'd74} : s = 154;
	{8'd80,8'd75} : s = 155;
	{8'd80,8'd76} : s = 156;
	{8'd80,8'd77} : s = 157;
	{8'd80,8'd78} : s = 158;
	{8'd80,8'd79} : s = 159;
	{8'd80,8'd80} : s = 160;
	{8'd80,8'd81} : s = 161;
	{8'd80,8'd82} : s = 162;
	{8'd80,8'd83} : s = 163;
	{8'd80,8'd84} : s = 164;
	{8'd80,8'd85} : s = 165;
	{8'd80,8'd86} : s = 166;
	{8'd80,8'd87} : s = 167;
	{8'd80,8'd88} : s = 168;
	{8'd80,8'd89} : s = 169;
	{8'd80,8'd90} : s = 170;
	{8'd80,8'd91} : s = 171;
	{8'd80,8'd92} : s = 172;
	{8'd80,8'd93} : s = 173;
	{8'd80,8'd94} : s = 174;
	{8'd80,8'd95} : s = 175;
	{8'd80,8'd96} : s = 176;
	{8'd80,8'd97} : s = 177;
	{8'd80,8'd98} : s = 178;
	{8'd80,8'd99} : s = 179;
	{8'd80,8'd100} : s = 180;
	{8'd80,8'd101} : s = 181;
	{8'd80,8'd102} : s = 182;
	{8'd80,8'd103} : s = 183;
	{8'd80,8'd104} : s = 184;
	{8'd80,8'd105} : s = 185;
	{8'd80,8'd106} : s = 186;
	{8'd80,8'd107} : s = 187;
	{8'd80,8'd108} : s = 188;
	{8'd80,8'd109} : s = 189;
	{8'd80,8'd110} : s = 190;
	{8'd80,8'd111} : s = 191;
	{8'd80,8'd112} : s = 192;
	{8'd80,8'd113} : s = 193;
	{8'd80,8'd114} : s = 194;
	{8'd80,8'd115} : s = 195;
	{8'd80,8'd116} : s = 196;
	{8'd80,8'd117} : s = 197;
	{8'd80,8'd118} : s = 198;
	{8'd80,8'd119} : s = 199;
	{8'd80,8'd120} : s = 200;
	{8'd80,8'd121} : s = 201;
	{8'd80,8'd122} : s = 202;
	{8'd80,8'd123} : s = 203;
	{8'd80,8'd124} : s = 204;
	{8'd80,8'd125} : s = 205;
	{8'd80,8'd126} : s = 206;
	{8'd80,8'd127} : s = 207;
	{8'd80,8'd128} : s = 208;
	{8'd80,8'd129} : s = 209;
	{8'd80,8'd130} : s = 210;
	{8'd80,8'd131} : s = 211;
	{8'd80,8'd132} : s = 212;
	{8'd80,8'd133} : s = 213;
	{8'd80,8'd134} : s = 214;
	{8'd80,8'd135} : s = 215;
	{8'd80,8'd136} : s = 216;
	{8'd80,8'd137} : s = 217;
	{8'd80,8'd138} : s = 218;
	{8'd80,8'd139} : s = 219;
	{8'd80,8'd140} : s = 220;
	{8'd80,8'd141} : s = 221;
	{8'd80,8'd142} : s = 222;
	{8'd80,8'd143} : s = 223;
	{8'd80,8'd144} : s = 224;
	{8'd80,8'd145} : s = 225;
	{8'd80,8'd146} : s = 226;
	{8'd80,8'd147} : s = 227;
	{8'd80,8'd148} : s = 228;
	{8'd80,8'd149} : s = 229;
	{8'd80,8'd150} : s = 230;
	{8'd80,8'd151} : s = 231;
	{8'd80,8'd152} : s = 232;
	{8'd80,8'd153} : s = 233;
	{8'd80,8'd154} : s = 234;
	{8'd80,8'd155} : s = 235;
	{8'd80,8'd156} : s = 236;
	{8'd80,8'd157} : s = 237;
	{8'd80,8'd158} : s = 238;
	{8'd80,8'd159} : s = 239;
	{8'd80,8'd160} : s = 240;
	{8'd80,8'd161} : s = 241;
	{8'd80,8'd162} : s = 242;
	{8'd80,8'd163} : s = 243;
	{8'd80,8'd164} : s = 244;
	{8'd80,8'd165} : s = 245;
	{8'd80,8'd166} : s = 246;
	{8'd80,8'd167} : s = 247;
	{8'd80,8'd168} : s = 248;
	{8'd80,8'd169} : s = 249;
	{8'd80,8'd170} : s = 250;
	{8'd80,8'd171} : s = 251;
	{8'd80,8'd172} : s = 252;
	{8'd80,8'd173} : s = 253;
	{8'd80,8'd174} : s = 254;
	{8'd80,8'd175} : s = 255;
	{8'd80,8'd176} : s = 256;
	{8'd80,8'd177} : s = 257;
	{8'd80,8'd178} : s = 258;
	{8'd80,8'd179} : s = 259;
	{8'd80,8'd180} : s = 260;
	{8'd80,8'd181} : s = 261;
	{8'd80,8'd182} : s = 262;
	{8'd80,8'd183} : s = 263;
	{8'd80,8'd184} : s = 264;
	{8'd80,8'd185} : s = 265;
	{8'd80,8'd186} : s = 266;
	{8'd80,8'd187} : s = 267;
	{8'd80,8'd188} : s = 268;
	{8'd80,8'd189} : s = 269;
	{8'd80,8'd190} : s = 270;
	{8'd80,8'd191} : s = 271;
	{8'd80,8'd192} : s = 272;
	{8'd80,8'd193} : s = 273;
	{8'd80,8'd194} : s = 274;
	{8'd80,8'd195} : s = 275;
	{8'd80,8'd196} : s = 276;
	{8'd80,8'd197} : s = 277;
	{8'd80,8'd198} : s = 278;
	{8'd80,8'd199} : s = 279;
	{8'd80,8'd200} : s = 280;
	{8'd80,8'd201} : s = 281;
	{8'd80,8'd202} : s = 282;
	{8'd80,8'd203} : s = 283;
	{8'd80,8'd204} : s = 284;
	{8'd80,8'd205} : s = 285;
	{8'd80,8'd206} : s = 286;
	{8'd80,8'd207} : s = 287;
	{8'd80,8'd208} : s = 288;
	{8'd80,8'd209} : s = 289;
	{8'd80,8'd210} : s = 290;
	{8'd80,8'd211} : s = 291;
	{8'd80,8'd212} : s = 292;
	{8'd80,8'd213} : s = 293;
	{8'd80,8'd214} : s = 294;
	{8'd80,8'd215} : s = 295;
	{8'd80,8'd216} : s = 296;
	{8'd80,8'd217} : s = 297;
	{8'd80,8'd218} : s = 298;
	{8'd80,8'd219} : s = 299;
	{8'd80,8'd220} : s = 300;
	{8'd80,8'd221} : s = 301;
	{8'd80,8'd222} : s = 302;
	{8'd80,8'd223} : s = 303;
	{8'd80,8'd224} : s = 304;
	{8'd80,8'd225} : s = 305;
	{8'd80,8'd226} : s = 306;
	{8'd80,8'd227} : s = 307;
	{8'd80,8'd228} : s = 308;
	{8'd80,8'd229} : s = 309;
	{8'd80,8'd230} : s = 310;
	{8'd80,8'd231} : s = 311;
	{8'd80,8'd232} : s = 312;
	{8'd80,8'd233} : s = 313;
	{8'd80,8'd234} : s = 314;
	{8'd80,8'd235} : s = 315;
	{8'd80,8'd236} : s = 316;
	{8'd80,8'd237} : s = 317;
	{8'd80,8'd238} : s = 318;
	{8'd80,8'd239} : s = 319;
	{8'd80,8'd240} : s = 320;
	{8'd80,8'd241} : s = 321;
	{8'd80,8'd242} : s = 322;
	{8'd80,8'd243} : s = 323;
	{8'd80,8'd244} : s = 324;
	{8'd80,8'd245} : s = 325;
	{8'd80,8'd246} : s = 326;
	{8'd80,8'd247} : s = 327;
	{8'd80,8'd248} : s = 328;
	{8'd80,8'd249} : s = 329;
	{8'd80,8'd250} : s = 330;
	{8'd80,8'd251} : s = 331;
	{8'd80,8'd252} : s = 332;
	{8'd80,8'd253} : s = 333;
	{8'd80,8'd254} : s = 334;
	{8'd80,8'd255} : s = 335;
	{8'd81,8'd0} : s = 81;
	{8'd81,8'd1} : s = 82;
	{8'd81,8'd2} : s = 83;
	{8'd81,8'd3} : s = 84;
	{8'd81,8'd4} : s = 85;
	{8'd81,8'd5} : s = 86;
	{8'd81,8'd6} : s = 87;
	{8'd81,8'd7} : s = 88;
	{8'd81,8'd8} : s = 89;
	{8'd81,8'd9} : s = 90;
	{8'd81,8'd10} : s = 91;
	{8'd81,8'd11} : s = 92;
	{8'd81,8'd12} : s = 93;
	{8'd81,8'd13} : s = 94;
	{8'd81,8'd14} : s = 95;
	{8'd81,8'd15} : s = 96;
	{8'd81,8'd16} : s = 97;
	{8'd81,8'd17} : s = 98;
	{8'd81,8'd18} : s = 99;
	{8'd81,8'd19} : s = 100;
	{8'd81,8'd20} : s = 101;
	{8'd81,8'd21} : s = 102;
	{8'd81,8'd22} : s = 103;
	{8'd81,8'd23} : s = 104;
	{8'd81,8'd24} : s = 105;
	{8'd81,8'd25} : s = 106;
	{8'd81,8'd26} : s = 107;
	{8'd81,8'd27} : s = 108;
	{8'd81,8'd28} : s = 109;
	{8'd81,8'd29} : s = 110;
	{8'd81,8'd30} : s = 111;
	{8'd81,8'd31} : s = 112;
	{8'd81,8'd32} : s = 113;
	{8'd81,8'd33} : s = 114;
	{8'd81,8'd34} : s = 115;
	{8'd81,8'd35} : s = 116;
	{8'd81,8'd36} : s = 117;
	{8'd81,8'd37} : s = 118;
	{8'd81,8'd38} : s = 119;
	{8'd81,8'd39} : s = 120;
	{8'd81,8'd40} : s = 121;
	{8'd81,8'd41} : s = 122;
	{8'd81,8'd42} : s = 123;
	{8'd81,8'd43} : s = 124;
	{8'd81,8'd44} : s = 125;
	{8'd81,8'd45} : s = 126;
	{8'd81,8'd46} : s = 127;
	{8'd81,8'd47} : s = 128;
	{8'd81,8'd48} : s = 129;
	{8'd81,8'd49} : s = 130;
	{8'd81,8'd50} : s = 131;
	{8'd81,8'd51} : s = 132;
	{8'd81,8'd52} : s = 133;
	{8'd81,8'd53} : s = 134;
	{8'd81,8'd54} : s = 135;
	{8'd81,8'd55} : s = 136;
	{8'd81,8'd56} : s = 137;
	{8'd81,8'd57} : s = 138;
	{8'd81,8'd58} : s = 139;
	{8'd81,8'd59} : s = 140;
	{8'd81,8'd60} : s = 141;
	{8'd81,8'd61} : s = 142;
	{8'd81,8'd62} : s = 143;
	{8'd81,8'd63} : s = 144;
	{8'd81,8'd64} : s = 145;
	{8'd81,8'd65} : s = 146;
	{8'd81,8'd66} : s = 147;
	{8'd81,8'd67} : s = 148;
	{8'd81,8'd68} : s = 149;
	{8'd81,8'd69} : s = 150;
	{8'd81,8'd70} : s = 151;
	{8'd81,8'd71} : s = 152;
	{8'd81,8'd72} : s = 153;
	{8'd81,8'd73} : s = 154;
	{8'd81,8'd74} : s = 155;
	{8'd81,8'd75} : s = 156;
	{8'd81,8'd76} : s = 157;
	{8'd81,8'd77} : s = 158;
	{8'd81,8'd78} : s = 159;
	{8'd81,8'd79} : s = 160;
	{8'd81,8'd80} : s = 161;
	{8'd81,8'd81} : s = 162;
	{8'd81,8'd82} : s = 163;
	{8'd81,8'd83} : s = 164;
	{8'd81,8'd84} : s = 165;
	{8'd81,8'd85} : s = 166;
	{8'd81,8'd86} : s = 167;
	{8'd81,8'd87} : s = 168;
	{8'd81,8'd88} : s = 169;
	{8'd81,8'd89} : s = 170;
	{8'd81,8'd90} : s = 171;
	{8'd81,8'd91} : s = 172;
	{8'd81,8'd92} : s = 173;
	{8'd81,8'd93} : s = 174;
	{8'd81,8'd94} : s = 175;
	{8'd81,8'd95} : s = 176;
	{8'd81,8'd96} : s = 177;
	{8'd81,8'd97} : s = 178;
	{8'd81,8'd98} : s = 179;
	{8'd81,8'd99} : s = 180;
	{8'd81,8'd100} : s = 181;
	{8'd81,8'd101} : s = 182;
	{8'd81,8'd102} : s = 183;
	{8'd81,8'd103} : s = 184;
	{8'd81,8'd104} : s = 185;
	{8'd81,8'd105} : s = 186;
	{8'd81,8'd106} : s = 187;
	{8'd81,8'd107} : s = 188;
	{8'd81,8'd108} : s = 189;
	{8'd81,8'd109} : s = 190;
	{8'd81,8'd110} : s = 191;
	{8'd81,8'd111} : s = 192;
	{8'd81,8'd112} : s = 193;
	{8'd81,8'd113} : s = 194;
	{8'd81,8'd114} : s = 195;
	{8'd81,8'd115} : s = 196;
	{8'd81,8'd116} : s = 197;
	{8'd81,8'd117} : s = 198;
	{8'd81,8'd118} : s = 199;
	{8'd81,8'd119} : s = 200;
	{8'd81,8'd120} : s = 201;
	{8'd81,8'd121} : s = 202;
	{8'd81,8'd122} : s = 203;
	{8'd81,8'd123} : s = 204;
	{8'd81,8'd124} : s = 205;
	{8'd81,8'd125} : s = 206;
	{8'd81,8'd126} : s = 207;
	{8'd81,8'd127} : s = 208;
	{8'd81,8'd128} : s = 209;
	{8'd81,8'd129} : s = 210;
	{8'd81,8'd130} : s = 211;
	{8'd81,8'd131} : s = 212;
	{8'd81,8'd132} : s = 213;
	{8'd81,8'd133} : s = 214;
	{8'd81,8'd134} : s = 215;
	{8'd81,8'd135} : s = 216;
	{8'd81,8'd136} : s = 217;
	{8'd81,8'd137} : s = 218;
	{8'd81,8'd138} : s = 219;
	{8'd81,8'd139} : s = 220;
	{8'd81,8'd140} : s = 221;
	{8'd81,8'd141} : s = 222;
	{8'd81,8'd142} : s = 223;
	{8'd81,8'd143} : s = 224;
	{8'd81,8'd144} : s = 225;
	{8'd81,8'd145} : s = 226;
	{8'd81,8'd146} : s = 227;
	{8'd81,8'd147} : s = 228;
	{8'd81,8'd148} : s = 229;
	{8'd81,8'd149} : s = 230;
	{8'd81,8'd150} : s = 231;
	{8'd81,8'd151} : s = 232;
	{8'd81,8'd152} : s = 233;
	{8'd81,8'd153} : s = 234;
	{8'd81,8'd154} : s = 235;
	{8'd81,8'd155} : s = 236;
	{8'd81,8'd156} : s = 237;
	{8'd81,8'd157} : s = 238;
	{8'd81,8'd158} : s = 239;
	{8'd81,8'd159} : s = 240;
	{8'd81,8'd160} : s = 241;
	{8'd81,8'd161} : s = 242;
	{8'd81,8'd162} : s = 243;
	{8'd81,8'd163} : s = 244;
	{8'd81,8'd164} : s = 245;
	{8'd81,8'd165} : s = 246;
	{8'd81,8'd166} : s = 247;
	{8'd81,8'd167} : s = 248;
	{8'd81,8'd168} : s = 249;
	{8'd81,8'd169} : s = 250;
	{8'd81,8'd170} : s = 251;
	{8'd81,8'd171} : s = 252;
	{8'd81,8'd172} : s = 253;
	{8'd81,8'd173} : s = 254;
	{8'd81,8'd174} : s = 255;
	{8'd81,8'd175} : s = 256;
	{8'd81,8'd176} : s = 257;
	{8'd81,8'd177} : s = 258;
	{8'd81,8'd178} : s = 259;
	{8'd81,8'd179} : s = 260;
	{8'd81,8'd180} : s = 261;
	{8'd81,8'd181} : s = 262;
	{8'd81,8'd182} : s = 263;
	{8'd81,8'd183} : s = 264;
	{8'd81,8'd184} : s = 265;
	{8'd81,8'd185} : s = 266;
	{8'd81,8'd186} : s = 267;
	{8'd81,8'd187} : s = 268;
	{8'd81,8'd188} : s = 269;
	{8'd81,8'd189} : s = 270;
	{8'd81,8'd190} : s = 271;
	{8'd81,8'd191} : s = 272;
	{8'd81,8'd192} : s = 273;
	{8'd81,8'd193} : s = 274;
	{8'd81,8'd194} : s = 275;
	{8'd81,8'd195} : s = 276;
	{8'd81,8'd196} : s = 277;
	{8'd81,8'd197} : s = 278;
	{8'd81,8'd198} : s = 279;
	{8'd81,8'd199} : s = 280;
	{8'd81,8'd200} : s = 281;
	{8'd81,8'd201} : s = 282;
	{8'd81,8'd202} : s = 283;
	{8'd81,8'd203} : s = 284;
	{8'd81,8'd204} : s = 285;
	{8'd81,8'd205} : s = 286;
	{8'd81,8'd206} : s = 287;
	{8'd81,8'd207} : s = 288;
	{8'd81,8'd208} : s = 289;
	{8'd81,8'd209} : s = 290;
	{8'd81,8'd210} : s = 291;
	{8'd81,8'd211} : s = 292;
	{8'd81,8'd212} : s = 293;
	{8'd81,8'd213} : s = 294;
	{8'd81,8'd214} : s = 295;
	{8'd81,8'd215} : s = 296;
	{8'd81,8'd216} : s = 297;
	{8'd81,8'd217} : s = 298;
	{8'd81,8'd218} : s = 299;
	{8'd81,8'd219} : s = 300;
	{8'd81,8'd220} : s = 301;
	{8'd81,8'd221} : s = 302;
	{8'd81,8'd222} : s = 303;
	{8'd81,8'd223} : s = 304;
	{8'd81,8'd224} : s = 305;
	{8'd81,8'd225} : s = 306;
	{8'd81,8'd226} : s = 307;
	{8'd81,8'd227} : s = 308;
	{8'd81,8'd228} : s = 309;
	{8'd81,8'd229} : s = 310;
	{8'd81,8'd230} : s = 311;
	{8'd81,8'd231} : s = 312;
	{8'd81,8'd232} : s = 313;
	{8'd81,8'd233} : s = 314;
	{8'd81,8'd234} : s = 315;
	{8'd81,8'd235} : s = 316;
	{8'd81,8'd236} : s = 317;
	{8'd81,8'd237} : s = 318;
	{8'd81,8'd238} : s = 319;
	{8'd81,8'd239} : s = 320;
	{8'd81,8'd240} : s = 321;
	{8'd81,8'd241} : s = 322;
	{8'd81,8'd242} : s = 323;
	{8'd81,8'd243} : s = 324;
	{8'd81,8'd244} : s = 325;
	{8'd81,8'd245} : s = 326;
	{8'd81,8'd246} : s = 327;
	{8'd81,8'd247} : s = 328;
	{8'd81,8'd248} : s = 329;
	{8'd81,8'd249} : s = 330;
	{8'd81,8'd250} : s = 331;
	{8'd81,8'd251} : s = 332;
	{8'd81,8'd252} : s = 333;
	{8'd81,8'd253} : s = 334;
	{8'd81,8'd254} : s = 335;
	{8'd81,8'd255} : s = 336;
	{8'd82,8'd0} : s = 82;
	{8'd82,8'd1} : s = 83;
	{8'd82,8'd2} : s = 84;
	{8'd82,8'd3} : s = 85;
	{8'd82,8'd4} : s = 86;
	{8'd82,8'd5} : s = 87;
	{8'd82,8'd6} : s = 88;
	{8'd82,8'd7} : s = 89;
	{8'd82,8'd8} : s = 90;
	{8'd82,8'd9} : s = 91;
	{8'd82,8'd10} : s = 92;
	{8'd82,8'd11} : s = 93;
	{8'd82,8'd12} : s = 94;
	{8'd82,8'd13} : s = 95;
	{8'd82,8'd14} : s = 96;
	{8'd82,8'd15} : s = 97;
	{8'd82,8'd16} : s = 98;
	{8'd82,8'd17} : s = 99;
	{8'd82,8'd18} : s = 100;
	{8'd82,8'd19} : s = 101;
	{8'd82,8'd20} : s = 102;
	{8'd82,8'd21} : s = 103;
	{8'd82,8'd22} : s = 104;
	{8'd82,8'd23} : s = 105;
	{8'd82,8'd24} : s = 106;
	{8'd82,8'd25} : s = 107;
	{8'd82,8'd26} : s = 108;
	{8'd82,8'd27} : s = 109;
	{8'd82,8'd28} : s = 110;
	{8'd82,8'd29} : s = 111;
	{8'd82,8'd30} : s = 112;
	{8'd82,8'd31} : s = 113;
	{8'd82,8'd32} : s = 114;
	{8'd82,8'd33} : s = 115;
	{8'd82,8'd34} : s = 116;
	{8'd82,8'd35} : s = 117;
	{8'd82,8'd36} : s = 118;
	{8'd82,8'd37} : s = 119;
	{8'd82,8'd38} : s = 120;
	{8'd82,8'd39} : s = 121;
	{8'd82,8'd40} : s = 122;
	{8'd82,8'd41} : s = 123;
	{8'd82,8'd42} : s = 124;
	{8'd82,8'd43} : s = 125;
	{8'd82,8'd44} : s = 126;
	{8'd82,8'd45} : s = 127;
	{8'd82,8'd46} : s = 128;
	{8'd82,8'd47} : s = 129;
	{8'd82,8'd48} : s = 130;
	{8'd82,8'd49} : s = 131;
	{8'd82,8'd50} : s = 132;
	{8'd82,8'd51} : s = 133;
	{8'd82,8'd52} : s = 134;
	{8'd82,8'd53} : s = 135;
	{8'd82,8'd54} : s = 136;
	{8'd82,8'd55} : s = 137;
	{8'd82,8'd56} : s = 138;
	{8'd82,8'd57} : s = 139;
	{8'd82,8'd58} : s = 140;
	{8'd82,8'd59} : s = 141;
	{8'd82,8'd60} : s = 142;
	{8'd82,8'd61} : s = 143;
	{8'd82,8'd62} : s = 144;
	{8'd82,8'd63} : s = 145;
	{8'd82,8'd64} : s = 146;
	{8'd82,8'd65} : s = 147;
	{8'd82,8'd66} : s = 148;
	{8'd82,8'd67} : s = 149;
	{8'd82,8'd68} : s = 150;
	{8'd82,8'd69} : s = 151;
	{8'd82,8'd70} : s = 152;
	{8'd82,8'd71} : s = 153;
	{8'd82,8'd72} : s = 154;
	{8'd82,8'd73} : s = 155;
	{8'd82,8'd74} : s = 156;
	{8'd82,8'd75} : s = 157;
	{8'd82,8'd76} : s = 158;
	{8'd82,8'd77} : s = 159;
	{8'd82,8'd78} : s = 160;
	{8'd82,8'd79} : s = 161;
	{8'd82,8'd80} : s = 162;
	{8'd82,8'd81} : s = 163;
	{8'd82,8'd82} : s = 164;
	{8'd82,8'd83} : s = 165;
	{8'd82,8'd84} : s = 166;
	{8'd82,8'd85} : s = 167;
	{8'd82,8'd86} : s = 168;
	{8'd82,8'd87} : s = 169;
	{8'd82,8'd88} : s = 170;
	{8'd82,8'd89} : s = 171;
	{8'd82,8'd90} : s = 172;
	{8'd82,8'd91} : s = 173;
	{8'd82,8'd92} : s = 174;
	{8'd82,8'd93} : s = 175;
	{8'd82,8'd94} : s = 176;
	{8'd82,8'd95} : s = 177;
	{8'd82,8'd96} : s = 178;
	{8'd82,8'd97} : s = 179;
	{8'd82,8'd98} : s = 180;
	{8'd82,8'd99} : s = 181;
	{8'd82,8'd100} : s = 182;
	{8'd82,8'd101} : s = 183;
	{8'd82,8'd102} : s = 184;
	{8'd82,8'd103} : s = 185;
	{8'd82,8'd104} : s = 186;
	{8'd82,8'd105} : s = 187;
	{8'd82,8'd106} : s = 188;
	{8'd82,8'd107} : s = 189;
	{8'd82,8'd108} : s = 190;
	{8'd82,8'd109} : s = 191;
	{8'd82,8'd110} : s = 192;
	{8'd82,8'd111} : s = 193;
	{8'd82,8'd112} : s = 194;
	{8'd82,8'd113} : s = 195;
	{8'd82,8'd114} : s = 196;
	{8'd82,8'd115} : s = 197;
	{8'd82,8'd116} : s = 198;
	{8'd82,8'd117} : s = 199;
	{8'd82,8'd118} : s = 200;
	{8'd82,8'd119} : s = 201;
	{8'd82,8'd120} : s = 202;
	{8'd82,8'd121} : s = 203;
	{8'd82,8'd122} : s = 204;
	{8'd82,8'd123} : s = 205;
	{8'd82,8'd124} : s = 206;
	{8'd82,8'd125} : s = 207;
	{8'd82,8'd126} : s = 208;
	{8'd82,8'd127} : s = 209;
	{8'd82,8'd128} : s = 210;
	{8'd82,8'd129} : s = 211;
	{8'd82,8'd130} : s = 212;
	{8'd82,8'd131} : s = 213;
	{8'd82,8'd132} : s = 214;
	{8'd82,8'd133} : s = 215;
	{8'd82,8'd134} : s = 216;
	{8'd82,8'd135} : s = 217;
	{8'd82,8'd136} : s = 218;
	{8'd82,8'd137} : s = 219;
	{8'd82,8'd138} : s = 220;
	{8'd82,8'd139} : s = 221;
	{8'd82,8'd140} : s = 222;
	{8'd82,8'd141} : s = 223;
	{8'd82,8'd142} : s = 224;
	{8'd82,8'd143} : s = 225;
	{8'd82,8'd144} : s = 226;
	{8'd82,8'd145} : s = 227;
	{8'd82,8'd146} : s = 228;
	{8'd82,8'd147} : s = 229;
	{8'd82,8'd148} : s = 230;
	{8'd82,8'd149} : s = 231;
	{8'd82,8'd150} : s = 232;
	{8'd82,8'd151} : s = 233;
	{8'd82,8'd152} : s = 234;
	{8'd82,8'd153} : s = 235;
	{8'd82,8'd154} : s = 236;
	{8'd82,8'd155} : s = 237;
	{8'd82,8'd156} : s = 238;
	{8'd82,8'd157} : s = 239;
	{8'd82,8'd158} : s = 240;
	{8'd82,8'd159} : s = 241;
	{8'd82,8'd160} : s = 242;
	{8'd82,8'd161} : s = 243;
	{8'd82,8'd162} : s = 244;
	{8'd82,8'd163} : s = 245;
	{8'd82,8'd164} : s = 246;
	{8'd82,8'd165} : s = 247;
	{8'd82,8'd166} : s = 248;
	{8'd82,8'd167} : s = 249;
	{8'd82,8'd168} : s = 250;
	{8'd82,8'd169} : s = 251;
	{8'd82,8'd170} : s = 252;
	{8'd82,8'd171} : s = 253;
	{8'd82,8'd172} : s = 254;
	{8'd82,8'd173} : s = 255;
	{8'd82,8'd174} : s = 256;
	{8'd82,8'd175} : s = 257;
	{8'd82,8'd176} : s = 258;
	{8'd82,8'd177} : s = 259;
	{8'd82,8'd178} : s = 260;
	{8'd82,8'd179} : s = 261;
	{8'd82,8'd180} : s = 262;
	{8'd82,8'd181} : s = 263;
	{8'd82,8'd182} : s = 264;
	{8'd82,8'd183} : s = 265;
	{8'd82,8'd184} : s = 266;
	{8'd82,8'd185} : s = 267;
	{8'd82,8'd186} : s = 268;
	{8'd82,8'd187} : s = 269;
	{8'd82,8'd188} : s = 270;
	{8'd82,8'd189} : s = 271;
	{8'd82,8'd190} : s = 272;
	{8'd82,8'd191} : s = 273;
	{8'd82,8'd192} : s = 274;
	{8'd82,8'd193} : s = 275;
	{8'd82,8'd194} : s = 276;
	{8'd82,8'd195} : s = 277;
	{8'd82,8'd196} : s = 278;
	{8'd82,8'd197} : s = 279;
	{8'd82,8'd198} : s = 280;
	{8'd82,8'd199} : s = 281;
	{8'd82,8'd200} : s = 282;
	{8'd82,8'd201} : s = 283;
	{8'd82,8'd202} : s = 284;
	{8'd82,8'd203} : s = 285;
	{8'd82,8'd204} : s = 286;
	{8'd82,8'd205} : s = 287;
	{8'd82,8'd206} : s = 288;
	{8'd82,8'd207} : s = 289;
	{8'd82,8'd208} : s = 290;
	{8'd82,8'd209} : s = 291;
	{8'd82,8'd210} : s = 292;
	{8'd82,8'd211} : s = 293;
	{8'd82,8'd212} : s = 294;
	{8'd82,8'd213} : s = 295;
	{8'd82,8'd214} : s = 296;
	{8'd82,8'd215} : s = 297;
	{8'd82,8'd216} : s = 298;
	{8'd82,8'd217} : s = 299;
	{8'd82,8'd218} : s = 300;
	{8'd82,8'd219} : s = 301;
	{8'd82,8'd220} : s = 302;
	{8'd82,8'd221} : s = 303;
	{8'd82,8'd222} : s = 304;
	{8'd82,8'd223} : s = 305;
	{8'd82,8'd224} : s = 306;
	{8'd82,8'd225} : s = 307;
	{8'd82,8'd226} : s = 308;
	{8'd82,8'd227} : s = 309;
	{8'd82,8'd228} : s = 310;
	{8'd82,8'd229} : s = 311;
	{8'd82,8'd230} : s = 312;
	{8'd82,8'd231} : s = 313;
	{8'd82,8'd232} : s = 314;
	{8'd82,8'd233} : s = 315;
	{8'd82,8'd234} : s = 316;
	{8'd82,8'd235} : s = 317;
	{8'd82,8'd236} : s = 318;
	{8'd82,8'd237} : s = 319;
	{8'd82,8'd238} : s = 320;
	{8'd82,8'd239} : s = 321;
	{8'd82,8'd240} : s = 322;
	{8'd82,8'd241} : s = 323;
	{8'd82,8'd242} : s = 324;
	{8'd82,8'd243} : s = 325;
	{8'd82,8'd244} : s = 326;
	{8'd82,8'd245} : s = 327;
	{8'd82,8'd246} : s = 328;
	{8'd82,8'd247} : s = 329;
	{8'd82,8'd248} : s = 330;
	{8'd82,8'd249} : s = 331;
	{8'd82,8'd250} : s = 332;
	{8'd82,8'd251} : s = 333;
	{8'd82,8'd252} : s = 334;
	{8'd82,8'd253} : s = 335;
	{8'd82,8'd254} : s = 336;
	{8'd82,8'd255} : s = 337;
	{8'd83,8'd0} : s = 83;
	{8'd83,8'd1} : s = 84;
	{8'd83,8'd2} : s = 85;
	{8'd83,8'd3} : s = 86;
	{8'd83,8'd4} : s = 87;
	{8'd83,8'd5} : s = 88;
	{8'd83,8'd6} : s = 89;
	{8'd83,8'd7} : s = 90;
	{8'd83,8'd8} : s = 91;
	{8'd83,8'd9} : s = 92;
	{8'd83,8'd10} : s = 93;
	{8'd83,8'd11} : s = 94;
	{8'd83,8'd12} : s = 95;
	{8'd83,8'd13} : s = 96;
	{8'd83,8'd14} : s = 97;
	{8'd83,8'd15} : s = 98;
	{8'd83,8'd16} : s = 99;
	{8'd83,8'd17} : s = 100;
	{8'd83,8'd18} : s = 101;
	{8'd83,8'd19} : s = 102;
	{8'd83,8'd20} : s = 103;
	{8'd83,8'd21} : s = 104;
	{8'd83,8'd22} : s = 105;
	{8'd83,8'd23} : s = 106;
	{8'd83,8'd24} : s = 107;
	{8'd83,8'd25} : s = 108;
	{8'd83,8'd26} : s = 109;
	{8'd83,8'd27} : s = 110;
	{8'd83,8'd28} : s = 111;
	{8'd83,8'd29} : s = 112;
	{8'd83,8'd30} : s = 113;
	{8'd83,8'd31} : s = 114;
	{8'd83,8'd32} : s = 115;
	{8'd83,8'd33} : s = 116;
	{8'd83,8'd34} : s = 117;
	{8'd83,8'd35} : s = 118;
	{8'd83,8'd36} : s = 119;
	{8'd83,8'd37} : s = 120;
	{8'd83,8'd38} : s = 121;
	{8'd83,8'd39} : s = 122;
	{8'd83,8'd40} : s = 123;
	{8'd83,8'd41} : s = 124;
	{8'd83,8'd42} : s = 125;
	{8'd83,8'd43} : s = 126;
	{8'd83,8'd44} : s = 127;
	{8'd83,8'd45} : s = 128;
	{8'd83,8'd46} : s = 129;
	{8'd83,8'd47} : s = 130;
	{8'd83,8'd48} : s = 131;
	{8'd83,8'd49} : s = 132;
	{8'd83,8'd50} : s = 133;
	{8'd83,8'd51} : s = 134;
	{8'd83,8'd52} : s = 135;
	{8'd83,8'd53} : s = 136;
	{8'd83,8'd54} : s = 137;
	{8'd83,8'd55} : s = 138;
	{8'd83,8'd56} : s = 139;
	{8'd83,8'd57} : s = 140;
	{8'd83,8'd58} : s = 141;
	{8'd83,8'd59} : s = 142;
	{8'd83,8'd60} : s = 143;
	{8'd83,8'd61} : s = 144;
	{8'd83,8'd62} : s = 145;
	{8'd83,8'd63} : s = 146;
	{8'd83,8'd64} : s = 147;
	{8'd83,8'd65} : s = 148;
	{8'd83,8'd66} : s = 149;
	{8'd83,8'd67} : s = 150;
	{8'd83,8'd68} : s = 151;
	{8'd83,8'd69} : s = 152;
	{8'd83,8'd70} : s = 153;
	{8'd83,8'd71} : s = 154;
	{8'd83,8'd72} : s = 155;
	{8'd83,8'd73} : s = 156;
	{8'd83,8'd74} : s = 157;
	{8'd83,8'd75} : s = 158;
	{8'd83,8'd76} : s = 159;
	{8'd83,8'd77} : s = 160;
	{8'd83,8'd78} : s = 161;
	{8'd83,8'd79} : s = 162;
	{8'd83,8'd80} : s = 163;
	{8'd83,8'd81} : s = 164;
	{8'd83,8'd82} : s = 165;
	{8'd83,8'd83} : s = 166;
	{8'd83,8'd84} : s = 167;
	{8'd83,8'd85} : s = 168;
	{8'd83,8'd86} : s = 169;
	{8'd83,8'd87} : s = 170;
	{8'd83,8'd88} : s = 171;
	{8'd83,8'd89} : s = 172;
	{8'd83,8'd90} : s = 173;
	{8'd83,8'd91} : s = 174;
	{8'd83,8'd92} : s = 175;
	{8'd83,8'd93} : s = 176;
	{8'd83,8'd94} : s = 177;
	{8'd83,8'd95} : s = 178;
	{8'd83,8'd96} : s = 179;
	{8'd83,8'd97} : s = 180;
	{8'd83,8'd98} : s = 181;
	{8'd83,8'd99} : s = 182;
	{8'd83,8'd100} : s = 183;
	{8'd83,8'd101} : s = 184;
	{8'd83,8'd102} : s = 185;
	{8'd83,8'd103} : s = 186;
	{8'd83,8'd104} : s = 187;
	{8'd83,8'd105} : s = 188;
	{8'd83,8'd106} : s = 189;
	{8'd83,8'd107} : s = 190;
	{8'd83,8'd108} : s = 191;
	{8'd83,8'd109} : s = 192;
	{8'd83,8'd110} : s = 193;
	{8'd83,8'd111} : s = 194;
	{8'd83,8'd112} : s = 195;
	{8'd83,8'd113} : s = 196;
	{8'd83,8'd114} : s = 197;
	{8'd83,8'd115} : s = 198;
	{8'd83,8'd116} : s = 199;
	{8'd83,8'd117} : s = 200;
	{8'd83,8'd118} : s = 201;
	{8'd83,8'd119} : s = 202;
	{8'd83,8'd120} : s = 203;
	{8'd83,8'd121} : s = 204;
	{8'd83,8'd122} : s = 205;
	{8'd83,8'd123} : s = 206;
	{8'd83,8'd124} : s = 207;
	{8'd83,8'd125} : s = 208;
	{8'd83,8'd126} : s = 209;
	{8'd83,8'd127} : s = 210;
	{8'd83,8'd128} : s = 211;
	{8'd83,8'd129} : s = 212;
	{8'd83,8'd130} : s = 213;
	{8'd83,8'd131} : s = 214;
	{8'd83,8'd132} : s = 215;
	{8'd83,8'd133} : s = 216;
	{8'd83,8'd134} : s = 217;
	{8'd83,8'd135} : s = 218;
	{8'd83,8'd136} : s = 219;
	{8'd83,8'd137} : s = 220;
	{8'd83,8'd138} : s = 221;
	{8'd83,8'd139} : s = 222;
	{8'd83,8'd140} : s = 223;
	{8'd83,8'd141} : s = 224;
	{8'd83,8'd142} : s = 225;
	{8'd83,8'd143} : s = 226;
	{8'd83,8'd144} : s = 227;
	{8'd83,8'd145} : s = 228;
	{8'd83,8'd146} : s = 229;
	{8'd83,8'd147} : s = 230;
	{8'd83,8'd148} : s = 231;
	{8'd83,8'd149} : s = 232;
	{8'd83,8'd150} : s = 233;
	{8'd83,8'd151} : s = 234;
	{8'd83,8'd152} : s = 235;
	{8'd83,8'd153} : s = 236;
	{8'd83,8'd154} : s = 237;
	{8'd83,8'd155} : s = 238;
	{8'd83,8'd156} : s = 239;
	{8'd83,8'd157} : s = 240;
	{8'd83,8'd158} : s = 241;
	{8'd83,8'd159} : s = 242;
	{8'd83,8'd160} : s = 243;
	{8'd83,8'd161} : s = 244;
	{8'd83,8'd162} : s = 245;
	{8'd83,8'd163} : s = 246;
	{8'd83,8'd164} : s = 247;
	{8'd83,8'd165} : s = 248;
	{8'd83,8'd166} : s = 249;
	{8'd83,8'd167} : s = 250;
	{8'd83,8'd168} : s = 251;
	{8'd83,8'd169} : s = 252;
	{8'd83,8'd170} : s = 253;
	{8'd83,8'd171} : s = 254;
	{8'd83,8'd172} : s = 255;
	{8'd83,8'd173} : s = 256;
	{8'd83,8'd174} : s = 257;
	{8'd83,8'd175} : s = 258;
	{8'd83,8'd176} : s = 259;
	{8'd83,8'd177} : s = 260;
	{8'd83,8'd178} : s = 261;
	{8'd83,8'd179} : s = 262;
	{8'd83,8'd180} : s = 263;
	{8'd83,8'd181} : s = 264;
	{8'd83,8'd182} : s = 265;
	{8'd83,8'd183} : s = 266;
	{8'd83,8'd184} : s = 267;
	{8'd83,8'd185} : s = 268;
	{8'd83,8'd186} : s = 269;
	{8'd83,8'd187} : s = 270;
	{8'd83,8'd188} : s = 271;
	{8'd83,8'd189} : s = 272;
	{8'd83,8'd190} : s = 273;
	{8'd83,8'd191} : s = 274;
	{8'd83,8'd192} : s = 275;
	{8'd83,8'd193} : s = 276;
	{8'd83,8'd194} : s = 277;
	{8'd83,8'd195} : s = 278;
	{8'd83,8'd196} : s = 279;
	{8'd83,8'd197} : s = 280;
	{8'd83,8'd198} : s = 281;
	{8'd83,8'd199} : s = 282;
	{8'd83,8'd200} : s = 283;
	{8'd83,8'd201} : s = 284;
	{8'd83,8'd202} : s = 285;
	{8'd83,8'd203} : s = 286;
	{8'd83,8'd204} : s = 287;
	{8'd83,8'd205} : s = 288;
	{8'd83,8'd206} : s = 289;
	{8'd83,8'd207} : s = 290;
	{8'd83,8'd208} : s = 291;
	{8'd83,8'd209} : s = 292;
	{8'd83,8'd210} : s = 293;
	{8'd83,8'd211} : s = 294;
	{8'd83,8'd212} : s = 295;
	{8'd83,8'd213} : s = 296;
	{8'd83,8'd214} : s = 297;
	{8'd83,8'd215} : s = 298;
	{8'd83,8'd216} : s = 299;
	{8'd83,8'd217} : s = 300;
	{8'd83,8'd218} : s = 301;
	{8'd83,8'd219} : s = 302;
	{8'd83,8'd220} : s = 303;
	{8'd83,8'd221} : s = 304;
	{8'd83,8'd222} : s = 305;
	{8'd83,8'd223} : s = 306;
	{8'd83,8'd224} : s = 307;
	{8'd83,8'd225} : s = 308;
	{8'd83,8'd226} : s = 309;
	{8'd83,8'd227} : s = 310;
	{8'd83,8'd228} : s = 311;
	{8'd83,8'd229} : s = 312;
	{8'd83,8'd230} : s = 313;
	{8'd83,8'd231} : s = 314;
	{8'd83,8'd232} : s = 315;
	{8'd83,8'd233} : s = 316;
	{8'd83,8'd234} : s = 317;
	{8'd83,8'd235} : s = 318;
	{8'd83,8'd236} : s = 319;
	{8'd83,8'd237} : s = 320;
	{8'd83,8'd238} : s = 321;
	{8'd83,8'd239} : s = 322;
	{8'd83,8'd240} : s = 323;
	{8'd83,8'd241} : s = 324;
	{8'd83,8'd242} : s = 325;
	{8'd83,8'd243} : s = 326;
	{8'd83,8'd244} : s = 327;
	{8'd83,8'd245} : s = 328;
	{8'd83,8'd246} : s = 329;
	{8'd83,8'd247} : s = 330;
	{8'd83,8'd248} : s = 331;
	{8'd83,8'd249} : s = 332;
	{8'd83,8'd250} : s = 333;
	{8'd83,8'd251} : s = 334;
	{8'd83,8'd252} : s = 335;
	{8'd83,8'd253} : s = 336;
	{8'd83,8'd254} : s = 337;
	{8'd83,8'd255} : s = 338;
	{8'd84,8'd0} : s = 84;
	{8'd84,8'd1} : s = 85;
	{8'd84,8'd2} : s = 86;
	{8'd84,8'd3} : s = 87;
	{8'd84,8'd4} : s = 88;
	{8'd84,8'd5} : s = 89;
	{8'd84,8'd6} : s = 90;
	{8'd84,8'd7} : s = 91;
	{8'd84,8'd8} : s = 92;
	{8'd84,8'd9} : s = 93;
	{8'd84,8'd10} : s = 94;
	{8'd84,8'd11} : s = 95;
	{8'd84,8'd12} : s = 96;
	{8'd84,8'd13} : s = 97;
	{8'd84,8'd14} : s = 98;
	{8'd84,8'd15} : s = 99;
	{8'd84,8'd16} : s = 100;
	{8'd84,8'd17} : s = 101;
	{8'd84,8'd18} : s = 102;
	{8'd84,8'd19} : s = 103;
	{8'd84,8'd20} : s = 104;
	{8'd84,8'd21} : s = 105;
	{8'd84,8'd22} : s = 106;
	{8'd84,8'd23} : s = 107;
	{8'd84,8'd24} : s = 108;
	{8'd84,8'd25} : s = 109;
	{8'd84,8'd26} : s = 110;
	{8'd84,8'd27} : s = 111;
	{8'd84,8'd28} : s = 112;
	{8'd84,8'd29} : s = 113;
	{8'd84,8'd30} : s = 114;
	{8'd84,8'd31} : s = 115;
	{8'd84,8'd32} : s = 116;
	{8'd84,8'd33} : s = 117;
	{8'd84,8'd34} : s = 118;
	{8'd84,8'd35} : s = 119;
	{8'd84,8'd36} : s = 120;
	{8'd84,8'd37} : s = 121;
	{8'd84,8'd38} : s = 122;
	{8'd84,8'd39} : s = 123;
	{8'd84,8'd40} : s = 124;
	{8'd84,8'd41} : s = 125;
	{8'd84,8'd42} : s = 126;
	{8'd84,8'd43} : s = 127;
	{8'd84,8'd44} : s = 128;
	{8'd84,8'd45} : s = 129;
	{8'd84,8'd46} : s = 130;
	{8'd84,8'd47} : s = 131;
	{8'd84,8'd48} : s = 132;
	{8'd84,8'd49} : s = 133;
	{8'd84,8'd50} : s = 134;
	{8'd84,8'd51} : s = 135;
	{8'd84,8'd52} : s = 136;
	{8'd84,8'd53} : s = 137;
	{8'd84,8'd54} : s = 138;
	{8'd84,8'd55} : s = 139;
	{8'd84,8'd56} : s = 140;
	{8'd84,8'd57} : s = 141;
	{8'd84,8'd58} : s = 142;
	{8'd84,8'd59} : s = 143;
	{8'd84,8'd60} : s = 144;
	{8'd84,8'd61} : s = 145;
	{8'd84,8'd62} : s = 146;
	{8'd84,8'd63} : s = 147;
	{8'd84,8'd64} : s = 148;
	{8'd84,8'd65} : s = 149;
	{8'd84,8'd66} : s = 150;
	{8'd84,8'd67} : s = 151;
	{8'd84,8'd68} : s = 152;
	{8'd84,8'd69} : s = 153;
	{8'd84,8'd70} : s = 154;
	{8'd84,8'd71} : s = 155;
	{8'd84,8'd72} : s = 156;
	{8'd84,8'd73} : s = 157;
	{8'd84,8'd74} : s = 158;
	{8'd84,8'd75} : s = 159;
	{8'd84,8'd76} : s = 160;
	{8'd84,8'd77} : s = 161;
	{8'd84,8'd78} : s = 162;
	{8'd84,8'd79} : s = 163;
	{8'd84,8'd80} : s = 164;
	{8'd84,8'd81} : s = 165;
	{8'd84,8'd82} : s = 166;
	{8'd84,8'd83} : s = 167;
	{8'd84,8'd84} : s = 168;
	{8'd84,8'd85} : s = 169;
	{8'd84,8'd86} : s = 170;
	{8'd84,8'd87} : s = 171;
	{8'd84,8'd88} : s = 172;
	{8'd84,8'd89} : s = 173;
	{8'd84,8'd90} : s = 174;
	{8'd84,8'd91} : s = 175;
	{8'd84,8'd92} : s = 176;
	{8'd84,8'd93} : s = 177;
	{8'd84,8'd94} : s = 178;
	{8'd84,8'd95} : s = 179;
	{8'd84,8'd96} : s = 180;
	{8'd84,8'd97} : s = 181;
	{8'd84,8'd98} : s = 182;
	{8'd84,8'd99} : s = 183;
	{8'd84,8'd100} : s = 184;
	{8'd84,8'd101} : s = 185;
	{8'd84,8'd102} : s = 186;
	{8'd84,8'd103} : s = 187;
	{8'd84,8'd104} : s = 188;
	{8'd84,8'd105} : s = 189;
	{8'd84,8'd106} : s = 190;
	{8'd84,8'd107} : s = 191;
	{8'd84,8'd108} : s = 192;
	{8'd84,8'd109} : s = 193;
	{8'd84,8'd110} : s = 194;
	{8'd84,8'd111} : s = 195;
	{8'd84,8'd112} : s = 196;
	{8'd84,8'd113} : s = 197;
	{8'd84,8'd114} : s = 198;
	{8'd84,8'd115} : s = 199;
	{8'd84,8'd116} : s = 200;
	{8'd84,8'd117} : s = 201;
	{8'd84,8'd118} : s = 202;
	{8'd84,8'd119} : s = 203;
	{8'd84,8'd120} : s = 204;
	{8'd84,8'd121} : s = 205;
	{8'd84,8'd122} : s = 206;
	{8'd84,8'd123} : s = 207;
	{8'd84,8'd124} : s = 208;
	{8'd84,8'd125} : s = 209;
	{8'd84,8'd126} : s = 210;
	{8'd84,8'd127} : s = 211;
	{8'd84,8'd128} : s = 212;
	{8'd84,8'd129} : s = 213;
	{8'd84,8'd130} : s = 214;
	{8'd84,8'd131} : s = 215;
	{8'd84,8'd132} : s = 216;
	{8'd84,8'd133} : s = 217;
	{8'd84,8'd134} : s = 218;
	{8'd84,8'd135} : s = 219;
	{8'd84,8'd136} : s = 220;
	{8'd84,8'd137} : s = 221;
	{8'd84,8'd138} : s = 222;
	{8'd84,8'd139} : s = 223;
	{8'd84,8'd140} : s = 224;
	{8'd84,8'd141} : s = 225;
	{8'd84,8'd142} : s = 226;
	{8'd84,8'd143} : s = 227;
	{8'd84,8'd144} : s = 228;
	{8'd84,8'd145} : s = 229;
	{8'd84,8'd146} : s = 230;
	{8'd84,8'd147} : s = 231;
	{8'd84,8'd148} : s = 232;
	{8'd84,8'd149} : s = 233;
	{8'd84,8'd150} : s = 234;
	{8'd84,8'd151} : s = 235;
	{8'd84,8'd152} : s = 236;
	{8'd84,8'd153} : s = 237;
	{8'd84,8'd154} : s = 238;
	{8'd84,8'd155} : s = 239;
	{8'd84,8'd156} : s = 240;
	{8'd84,8'd157} : s = 241;
	{8'd84,8'd158} : s = 242;
	{8'd84,8'd159} : s = 243;
	{8'd84,8'd160} : s = 244;
	{8'd84,8'd161} : s = 245;
	{8'd84,8'd162} : s = 246;
	{8'd84,8'd163} : s = 247;
	{8'd84,8'd164} : s = 248;
	{8'd84,8'd165} : s = 249;
	{8'd84,8'd166} : s = 250;
	{8'd84,8'd167} : s = 251;
	{8'd84,8'd168} : s = 252;
	{8'd84,8'd169} : s = 253;
	{8'd84,8'd170} : s = 254;
	{8'd84,8'd171} : s = 255;
	{8'd84,8'd172} : s = 256;
	{8'd84,8'd173} : s = 257;
	{8'd84,8'd174} : s = 258;
	{8'd84,8'd175} : s = 259;
	{8'd84,8'd176} : s = 260;
	{8'd84,8'd177} : s = 261;
	{8'd84,8'd178} : s = 262;
	{8'd84,8'd179} : s = 263;
	{8'd84,8'd180} : s = 264;
	{8'd84,8'd181} : s = 265;
	{8'd84,8'd182} : s = 266;
	{8'd84,8'd183} : s = 267;
	{8'd84,8'd184} : s = 268;
	{8'd84,8'd185} : s = 269;
	{8'd84,8'd186} : s = 270;
	{8'd84,8'd187} : s = 271;
	{8'd84,8'd188} : s = 272;
	{8'd84,8'd189} : s = 273;
	{8'd84,8'd190} : s = 274;
	{8'd84,8'd191} : s = 275;
	{8'd84,8'd192} : s = 276;
	{8'd84,8'd193} : s = 277;
	{8'd84,8'd194} : s = 278;
	{8'd84,8'd195} : s = 279;
	{8'd84,8'd196} : s = 280;
	{8'd84,8'd197} : s = 281;
	{8'd84,8'd198} : s = 282;
	{8'd84,8'd199} : s = 283;
	{8'd84,8'd200} : s = 284;
	{8'd84,8'd201} : s = 285;
	{8'd84,8'd202} : s = 286;
	{8'd84,8'd203} : s = 287;
	{8'd84,8'd204} : s = 288;
	{8'd84,8'd205} : s = 289;
	{8'd84,8'd206} : s = 290;
	{8'd84,8'd207} : s = 291;
	{8'd84,8'd208} : s = 292;
	{8'd84,8'd209} : s = 293;
	{8'd84,8'd210} : s = 294;
	{8'd84,8'd211} : s = 295;
	{8'd84,8'd212} : s = 296;
	{8'd84,8'd213} : s = 297;
	{8'd84,8'd214} : s = 298;
	{8'd84,8'd215} : s = 299;
	{8'd84,8'd216} : s = 300;
	{8'd84,8'd217} : s = 301;
	{8'd84,8'd218} : s = 302;
	{8'd84,8'd219} : s = 303;
	{8'd84,8'd220} : s = 304;
	{8'd84,8'd221} : s = 305;
	{8'd84,8'd222} : s = 306;
	{8'd84,8'd223} : s = 307;
	{8'd84,8'd224} : s = 308;
	{8'd84,8'd225} : s = 309;
	{8'd84,8'd226} : s = 310;
	{8'd84,8'd227} : s = 311;
	{8'd84,8'd228} : s = 312;
	{8'd84,8'd229} : s = 313;
	{8'd84,8'd230} : s = 314;
	{8'd84,8'd231} : s = 315;
	{8'd84,8'd232} : s = 316;
	{8'd84,8'd233} : s = 317;
	{8'd84,8'd234} : s = 318;
	{8'd84,8'd235} : s = 319;
	{8'd84,8'd236} : s = 320;
	{8'd84,8'd237} : s = 321;
	{8'd84,8'd238} : s = 322;
	{8'd84,8'd239} : s = 323;
	{8'd84,8'd240} : s = 324;
	{8'd84,8'd241} : s = 325;
	{8'd84,8'd242} : s = 326;
	{8'd84,8'd243} : s = 327;
	{8'd84,8'd244} : s = 328;
	{8'd84,8'd245} : s = 329;
	{8'd84,8'd246} : s = 330;
	{8'd84,8'd247} : s = 331;
	{8'd84,8'd248} : s = 332;
	{8'd84,8'd249} : s = 333;
	{8'd84,8'd250} : s = 334;
	{8'd84,8'd251} : s = 335;
	{8'd84,8'd252} : s = 336;
	{8'd84,8'd253} : s = 337;
	{8'd84,8'd254} : s = 338;
	{8'd84,8'd255} : s = 339;
	{8'd85,8'd0} : s = 85;
	{8'd85,8'd1} : s = 86;
	{8'd85,8'd2} : s = 87;
	{8'd85,8'd3} : s = 88;
	{8'd85,8'd4} : s = 89;
	{8'd85,8'd5} : s = 90;
	{8'd85,8'd6} : s = 91;
	{8'd85,8'd7} : s = 92;
	{8'd85,8'd8} : s = 93;
	{8'd85,8'd9} : s = 94;
	{8'd85,8'd10} : s = 95;
	{8'd85,8'd11} : s = 96;
	{8'd85,8'd12} : s = 97;
	{8'd85,8'd13} : s = 98;
	{8'd85,8'd14} : s = 99;
	{8'd85,8'd15} : s = 100;
	{8'd85,8'd16} : s = 101;
	{8'd85,8'd17} : s = 102;
	{8'd85,8'd18} : s = 103;
	{8'd85,8'd19} : s = 104;
	{8'd85,8'd20} : s = 105;
	{8'd85,8'd21} : s = 106;
	{8'd85,8'd22} : s = 107;
	{8'd85,8'd23} : s = 108;
	{8'd85,8'd24} : s = 109;
	{8'd85,8'd25} : s = 110;
	{8'd85,8'd26} : s = 111;
	{8'd85,8'd27} : s = 112;
	{8'd85,8'd28} : s = 113;
	{8'd85,8'd29} : s = 114;
	{8'd85,8'd30} : s = 115;
	{8'd85,8'd31} : s = 116;
	{8'd85,8'd32} : s = 117;
	{8'd85,8'd33} : s = 118;
	{8'd85,8'd34} : s = 119;
	{8'd85,8'd35} : s = 120;
	{8'd85,8'd36} : s = 121;
	{8'd85,8'd37} : s = 122;
	{8'd85,8'd38} : s = 123;
	{8'd85,8'd39} : s = 124;
	{8'd85,8'd40} : s = 125;
	{8'd85,8'd41} : s = 126;
	{8'd85,8'd42} : s = 127;
	{8'd85,8'd43} : s = 128;
	{8'd85,8'd44} : s = 129;
	{8'd85,8'd45} : s = 130;
	{8'd85,8'd46} : s = 131;
	{8'd85,8'd47} : s = 132;
	{8'd85,8'd48} : s = 133;
	{8'd85,8'd49} : s = 134;
	{8'd85,8'd50} : s = 135;
	{8'd85,8'd51} : s = 136;
	{8'd85,8'd52} : s = 137;
	{8'd85,8'd53} : s = 138;
	{8'd85,8'd54} : s = 139;
	{8'd85,8'd55} : s = 140;
	{8'd85,8'd56} : s = 141;
	{8'd85,8'd57} : s = 142;
	{8'd85,8'd58} : s = 143;
	{8'd85,8'd59} : s = 144;
	{8'd85,8'd60} : s = 145;
	{8'd85,8'd61} : s = 146;
	{8'd85,8'd62} : s = 147;
	{8'd85,8'd63} : s = 148;
	{8'd85,8'd64} : s = 149;
	{8'd85,8'd65} : s = 150;
	{8'd85,8'd66} : s = 151;
	{8'd85,8'd67} : s = 152;
	{8'd85,8'd68} : s = 153;
	{8'd85,8'd69} : s = 154;
	{8'd85,8'd70} : s = 155;
	{8'd85,8'd71} : s = 156;
	{8'd85,8'd72} : s = 157;
	{8'd85,8'd73} : s = 158;
	{8'd85,8'd74} : s = 159;
	{8'd85,8'd75} : s = 160;
	{8'd85,8'd76} : s = 161;
	{8'd85,8'd77} : s = 162;
	{8'd85,8'd78} : s = 163;
	{8'd85,8'd79} : s = 164;
	{8'd85,8'd80} : s = 165;
	{8'd85,8'd81} : s = 166;
	{8'd85,8'd82} : s = 167;
	{8'd85,8'd83} : s = 168;
	{8'd85,8'd84} : s = 169;
	{8'd85,8'd85} : s = 170;
	{8'd85,8'd86} : s = 171;
	{8'd85,8'd87} : s = 172;
	{8'd85,8'd88} : s = 173;
	{8'd85,8'd89} : s = 174;
	{8'd85,8'd90} : s = 175;
	{8'd85,8'd91} : s = 176;
	{8'd85,8'd92} : s = 177;
	{8'd85,8'd93} : s = 178;
	{8'd85,8'd94} : s = 179;
	{8'd85,8'd95} : s = 180;
	{8'd85,8'd96} : s = 181;
	{8'd85,8'd97} : s = 182;
	{8'd85,8'd98} : s = 183;
	{8'd85,8'd99} : s = 184;
	{8'd85,8'd100} : s = 185;
	{8'd85,8'd101} : s = 186;
	{8'd85,8'd102} : s = 187;
	{8'd85,8'd103} : s = 188;
	{8'd85,8'd104} : s = 189;
	{8'd85,8'd105} : s = 190;
	{8'd85,8'd106} : s = 191;
	{8'd85,8'd107} : s = 192;
	{8'd85,8'd108} : s = 193;
	{8'd85,8'd109} : s = 194;
	{8'd85,8'd110} : s = 195;
	{8'd85,8'd111} : s = 196;
	{8'd85,8'd112} : s = 197;
	{8'd85,8'd113} : s = 198;
	{8'd85,8'd114} : s = 199;
	{8'd85,8'd115} : s = 200;
	{8'd85,8'd116} : s = 201;
	{8'd85,8'd117} : s = 202;
	{8'd85,8'd118} : s = 203;
	{8'd85,8'd119} : s = 204;
	{8'd85,8'd120} : s = 205;
	{8'd85,8'd121} : s = 206;
	{8'd85,8'd122} : s = 207;
	{8'd85,8'd123} : s = 208;
	{8'd85,8'd124} : s = 209;
	{8'd85,8'd125} : s = 210;
	{8'd85,8'd126} : s = 211;
	{8'd85,8'd127} : s = 212;
	{8'd85,8'd128} : s = 213;
	{8'd85,8'd129} : s = 214;
	{8'd85,8'd130} : s = 215;
	{8'd85,8'd131} : s = 216;
	{8'd85,8'd132} : s = 217;
	{8'd85,8'd133} : s = 218;
	{8'd85,8'd134} : s = 219;
	{8'd85,8'd135} : s = 220;
	{8'd85,8'd136} : s = 221;
	{8'd85,8'd137} : s = 222;
	{8'd85,8'd138} : s = 223;
	{8'd85,8'd139} : s = 224;
	{8'd85,8'd140} : s = 225;
	{8'd85,8'd141} : s = 226;
	{8'd85,8'd142} : s = 227;
	{8'd85,8'd143} : s = 228;
	{8'd85,8'd144} : s = 229;
	{8'd85,8'd145} : s = 230;
	{8'd85,8'd146} : s = 231;
	{8'd85,8'd147} : s = 232;
	{8'd85,8'd148} : s = 233;
	{8'd85,8'd149} : s = 234;
	{8'd85,8'd150} : s = 235;
	{8'd85,8'd151} : s = 236;
	{8'd85,8'd152} : s = 237;
	{8'd85,8'd153} : s = 238;
	{8'd85,8'd154} : s = 239;
	{8'd85,8'd155} : s = 240;
	{8'd85,8'd156} : s = 241;
	{8'd85,8'd157} : s = 242;
	{8'd85,8'd158} : s = 243;
	{8'd85,8'd159} : s = 244;
	{8'd85,8'd160} : s = 245;
	{8'd85,8'd161} : s = 246;
	{8'd85,8'd162} : s = 247;
	{8'd85,8'd163} : s = 248;
	{8'd85,8'd164} : s = 249;
	{8'd85,8'd165} : s = 250;
	{8'd85,8'd166} : s = 251;
	{8'd85,8'd167} : s = 252;
	{8'd85,8'd168} : s = 253;
	{8'd85,8'd169} : s = 254;
	{8'd85,8'd170} : s = 255;
	{8'd85,8'd171} : s = 256;
	{8'd85,8'd172} : s = 257;
	{8'd85,8'd173} : s = 258;
	{8'd85,8'd174} : s = 259;
	{8'd85,8'd175} : s = 260;
	{8'd85,8'd176} : s = 261;
	{8'd85,8'd177} : s = 262;
	{8'd85,8'd178} : s = 263;
	{8'd85,8'd179} : s = 264;
	{8'd85,8'd180} : s = 265;
	{8'd85,8'd181} : s = 266;
	{8'd85,8'd182} : s = 267;
	{8'd85,8'd183} : s = 268;
	{8'd85,8'd184} : s = 269;
	{8'd85,8'd185} : s = 270;
	{8'd85,8'd186} : s = 271;
	{8'd85,8'd187} : s = 272;
	{8'd85,8'd188} : s = 273;
	{8'd85,8'd189} : s = 274;
	{8'd85,8'd190} : s = 275;
	{8'd85,8'd191} : s = 276;
	{8'd85,8'd192} : s = 277;
	{8'd85,8'd193} : s = 278;
	{8'd85,8'd194} : s = 279;
	{8'd85,8'd195} : s = 280;
	{8'd85,8'd196} : s = 281;
	{8'd85,8'd197} : s = 282;
	{8'd85,8'd198} : s = 283;
	{8'd85,8'd199} : s = 284;
	{8'd85,8'd200} : s = 285;
	{8'd85,8'd201} : s = 286;
	{8'd85,8'd202} : s = 287;
	{8'd85,8'd203} : s = 288;
	{8'd85,8'd204} : s = 289;
	{8'd85,8'd205} : s = 290;
	{8'd85,8'd206} : s = 291;
	{8'd85,8'd207} : s = 292;
	{8'd85,8'd208} : s = 293;
	{8'd85,8'd209} : s = 294;
	{8'd85,8'd210} : s = 295;
	{8'd85,8'd211} : s = 296;
	{8'd85,8'd212} : s = 297;
	{8'd85,8'd213} : s = 298;
	{8'd85,8'd214} : s = 299;
	{8'd85,8'd215} : s = 300;
	{8'd85,8'd216} : s = 301;
	{8'd85,8'd217} : s = 302;
	{8'd85,8'd218} : s = 303;
	{8'd85,8'd219} : s = 304;
	{8'd85,8'd220} : s = 305;
	{8'd85,8'd221} : s = 306;
	{8'd85,8'd222} : s = 307;
	{8'd85,8'd223} : s = 308;
	{8'd85,8'd224} : s = 309;
	{8'd85,8'd225} : s = 310;
	{8'd85,8'd226} : s = 311;
	{8'd85,8'd227} : s = 312;
	{8'd85,8'd228} : s = 313;
	{8'd85,8'd229} : s = 314;
	{8'd85,8'd230} : s = 315;
	{8'd85,8'd231} : s = 316;
	{8'd85,8'd232} : s = 317;
	{8'd85,8'd233} : s = 318;
	{8'd85,8'd234} : s = 319;
	{8'd85,8'd235} : s = 320;
	{8'd85,8'd236} : s = 321;
	{8'd85,8'd237} : s = 322;
	{8'd85,8'd238} : s = 323;
	{8'd85,8'd239} : s = 324;
	{8'd85,8'd240} : s = 325;
	{8'd85,8'd241} : s = 326;
	{8'd85,8'd242} : s = 327;
	{8'd85,8'd243} : s = 328;
	{8'd85,8'd244} : s = 329;
	{8'd85,8'd245} : s = 330;
	{8'd85,8'd246} : s = 331;
	{8'd85,8'd247} : s = 332;
	{8'd85,8'd248} : s = 333;
	{8'd85,8'd249} : s = 334;
	{8'd85,8'd250} : s = 335;
	{8'd85,8'd251} : s = 336;
	{8'd85,8'd252} : s = 337;
	{8'd85,8'd253} : s = 338;
	{8'd85,8'd254} : s = 339;
	{8'd85,8'd255} : s = 340;
	{8'd86,8'd0} : s = 86;
	{8'd86,8'd1} : s = 87;
	{8'd86,8'd2} : s = 88;
	{8'd86,8'd3} : s = 89;
	{8'd86,8'd4} : s = 90;
	{8'd86,8'd5} : s = 91;
	{8'd86,8'd6} : s = 92;
	{8'd86,8'd7} : s = 93;
	{8'd86,8'd8} : s = 94;
	{8'd86,8'd9} : s = 95;
	{8'd86,8'd10} : s = 96;
	{8'd86,8'd11} : s = 97;
	{8'd86,8'd12} : s = 98;
	{8'd86,8'd13} : s = 99;
	{8'd86,8'd14} : s = 100;
	{8'd86,8'd15} : s = 101;
	{8'd86,8'd16} : s = 102;
	{8'd86,8'd17} : s = 103;
	{8'd86,8'd18} : s = 104;
	{8'd86,8'd19} : s = 105;
	{8'd86,8'd20} : s = 106;
	{8'd86,8'd21} : s = 107;
	{8'd86,8'd22} : s = 108;
	{8'd86,8'd23} : s = 109;
	{8'd86,8'd24} : s = 110;
	{8'd86,8'd25} : s = 111;
	{8'd86,8'd26} : s = 112;
	{8'd86,8'd27} : s = 113;
	{8'd86,8'd28} : s = 114;
	{8'd86,8'd29} : s = 115;
	{8'd86,8'd30} : s = 116;
	{8'd86,8'd31} : s = 117;
	{8'd86,8'd32} : s = 118;
	{8'd86,8'd33} : s = 119;
	{8'd86,8'd34} : s = 120;
	{8'd86,8'd35} : s = 121;
	{8'd86,8'd36} : s = 122;
	{8'd86,8'd37} : s = 123;
	{8'd86,8'd38} : s = 124;
	{8'd86,8'd39} : s = 125;
	{8'd86,8'd40} : s = 126;
	{8'd86,8'd41} : s = 127;
	{8'd86,8'd42} : s = 128;
	{8'd86,8'd43} : s = 129;
	{8'd86,8'd44} : s = 130;
	{8'd86,8'd45} : s = 131;
	{8'd86,8'd46} : s = 132;
	{8'd86,8'd47} : s = 133;
	{8'd86,8'd48} : s = 134;
	{8'd86,8'd49} : s = 135;
	{8'd86,8'd50} : s = 136;
	{8'd86,8'd51} : s = 137;
	{8'd86,8'd52} : s = 138;
	{8'd86,8'd53} : s = 139;
	{8'd86,8'd54} : s = 140;
	{8'd86,8'd55} : s = 141;
	{8'd86,8'd56} : s = 142;
	{8'd86,8'd57} : s = 143;
	{8'd86,8'd58} : s = 144;
	{8'd86,8'd59} : s = 145;
	{8'd86,8'd60} : s = 146;
	{8'd86,8'd61} : s = 147;
	{8'd86,8'd62} : s = 148;
	{8'd86,8'd63} : s = 149;
	{8'd86,8'd64} : s = 150;
	{8'd86,8'd65} : s = 151;
	{8'd86,8'd66} : s = 152;
	{8'd86,8'd67} : s = 153;
	{8'd86,8'd68} : s = 154;
	{8'd86,8'd69} : s = 155;
	{8'd86,8'd70} : s = 156;
	{8'd86,8'd71} : s = 157;
	{8'd86,8'd72} : s = 158;
	{8'd86,8'd73} : s = 159;
	{8'd86,8'd74} : s = 160;
	{8'd86,8'd75} : s = 161;
	{8'd86,8'd76} : s = 162;
	{8'd86,8'd77} : s = 163;
	{8'd86,8'd78} : s = 164;
	{8'd86,8'd79} : s = 165;
	{8'd86,8'd80} : s = 166;
	{8'd86,8'd81} : s = 167;
	{8'd86,8'd82} : s = 168;
	{8'd86,8'd83} : s = 169;
	{8'd86,8'd84} : s = 170;
	{8'd86,8'd85} : s = 171;
	{8'd86,8'd86} : s = 172;
	{8'd86,8'd87} : s = 173;
	{8'd86,8'd88} : s = 174;
	{8'd86,8'd89} : s = 175;
	{8'd86,8'd90} : s = 176;
	{8'd86,8'd91} : s = 177;
	{8'd86,8'd92} : s = 178;
	{8'd86,8'd93} : s = 179;
	{8'd86,8'd94} : s = 180;
	{8'd86,8'd95} : s = 181;
	{8'd86,8'd96} : s = 182;
	{8'd86,8'd97} : s = 183;
	{8'd86,8'd98} : s = 184;
	{8'd86,8'd99} : s = 185;
	{8'd86,8'd100} : s = 186;
	{8'd86,8'd101} : s = 187;
	{8'd86,8'd102} : s = 188;
	{8'd86,8'd103} : s = 189;
	{8'd86,8'd104} : s = 190;
	{8'd86,8'd105} : s = 191;
	{8'd86,8'd106} : s = 192;
	{8'd86,8'd107} : s = 193;
	{8'd86,8'd108} : s = 194;
	{8'd86,8'd109} : s = 195;
	{8'd86,8'd110} : s = 196;
	{8'd86,8'd111} : s = 197;
	{8'd86,8'd112} : s = 198;
	{8'd86,8'd113} : s = 199;
	{8'd86,8'd114} : s = 200;
	{8'd86,8'd115} : s = 201;
	{8'd86,8'd116} : s = 202;
	{8'd86,8'd117} : s = 203;
	{8'd86,8'd118} : s = 204;
	{8'd86,8'd119} : s = 205;
	{8'd86,8'd120} : s = 206;
	{8'd86,8'd121} : s = 207;
	{8'd86,8'd122} : s = 208;
	{8'd86,8'd123} : s = 209;
	{8'd86,8'd124} : s = 210;
	{8'd86,8'd125} : s = 211;
	{8'd86,8'd126} : s = 212;
	{8'd86,8'd127} : s = 213;
	{8'd86,8'd128} : s = 214;
	{8'd86,8'd129} : s = 215;
	{8'd86,8'd130} : s = 216;
	{8'd86,8'd131} : s = 217;
	{8'd86,8'd132} : s = 218;
	{8'd86,8'd133} : s = 219;
	{8'd86,8'd134} : s = 220;
	{8'd86,8'd135} : s = 221;
	{8'd86,8'd136} : s = 222;
	{8'd86,8'd137} : s = 223;
	{8'd86,8'd138} : s = 224;
	{8'd86,8'd139} : s = 225;
	{8'd86,8'd140} : s = 226;
	{8'd86,8'd141} : s = 227;
	{8'd86,8'd142} : s = 228;
	{8'd86,8'd143} : s = 229;
	{8'd86,8'd144} : s = 230;
	{8'd86,8'd145} : s = 231;
	{8'd86,8'd146} : s = 232;
	{8'd86,8'd147} : s = 233;
	{8'd86,8'd148} : s = 234;
	{8'd86,8'd149} : s = 235;
	{8'd86,8'd150} : s = 236;
	{8'd86,8'd151} : s = 237;
	{8'd86,8'd152} : s = 238;
	{8'd86,8'd153} : s = 239;
	{8'd86,8'd154} : s = 240;
	{8'd86,8'd155} : s = 241;
	{8'd86,8'd156} : s = 242;
	{8'd86,8'd157} : s = 243;
	{8'd86,8'd158} : s = 244;
	{8'd86,8'd159} : s = 245;
	{8'd86,8'd160} : s = 246;
	{8'd86,8'd161} : s = 247;
	{8'd86,8'd162} : s = 248;
	{8'd86,8'd163} : s = 249;
	{8'd86,8'd164} : s = 250;
	{8'd86,8'd165} : s = 251;
	{8'd86,8'd166} : s = 252;
	{8'd86,8'd167} : s = 253;
	{8'd86,8'd168} : s = 254;
	{8'd86,8'd169} : s = 255;
	{8'd86,8'd170} : s = 256;
	{8'd86,8'd171} : s = 257;
	{8'd86,8'd172} : s = 258;
	{8'd86,8'd173} : s = 259;
	{8'd86,8'd174} : s = 260;
	{8'd86,8'd175} : s = 261;
	{8'd86,8'd176} : s = 262;
	{8'd86,8'd177} : s = 263;
	{8'd86,8'd178} : s = 264;
	{8'd86,8'd179} : s = 265;
	{8'd86,8'd180} : s = 266;
	{8'd86,8'd181} : s = 267;
	{8'd86,8'd182} : s = 268;
	{8'd86,8'd183} : s = 269;
	{8'd86,8'd184} : s = 270;
	{8'd86,8'd185} : s = 271;
	{8'd86,8'd186} : s = 272;
	{8'd86,8'd187} : s = 273;
	{8'd86,8'd188} : s = 274;
	{8'd86,8'd189} : s = 275;
	{8'd86,8'd190} : s = 276;
	{8'd86,8'd191} : s = 277;
	{8'd86,8'd192} : s = 278;
	{8'd86,8'd193} : s = 279;
	{8'd86,8'd194} : s = 280;
	{8'd86,8'd195} : s = 281;
	{8'd86,8'd196} : s = 282;
	{8'd86,8'd197} : s = 283;
	{8'd86,8'd198} : s = 284;
	{8'd86,8'd199} : s = 285;
	{8'd86,8'd200} : s = 286;
	{8'd86,8'd201} : s = 287;
	{8'd86,8'd202} : s = 288;
	{8'd86,8'd203} : s = 289;
	{8'd86,8'd204} : s = 290;
	{8'd86,8'd205} : s = 291;
	{8'd86,8'd206} : s = 292;
	{8'd86,8'd207} : s = 293;
	{8'd86,8'd208} : s = 294;
	{8'd86,8'd209} : s = 295;
	{8'd86,8'd210} : s = 296;
	{8'd86,8'd211} : s = 297;
	{8'd86,8'd212} : s = 298;
	{8'd86,8'd213} : s = 299;
	{8'd86,8'd214} : s = 300;
	{8'd86,8'd215} : s = 301;
	{8'd86,8'd216} : s = 302;
	{8'd86,8'd217} : s = 303;
	{8'd86,8'd218} : s = 304;
	{8'd86,8'd219} : s = 305;
	{8'd86,8'd220} : s = 306;
	{8'd86,8'd221} : s = 307;
	{8'd86,8'd222} : s = 308;
	{8'd86,8'd223} : s = 309;
	{8'd86,8'd224} : s = 310;
	{8'd86,8'd225} : s = 311;
	{8'd86,8'd226} : s = 312;
	{8'd86,8'd227} : s = 313;
	{8'd86,8'd228} : s = 314;
	{8'd86,8'd229} : s = 315;
	{8'd86,8'd230} : s = 316;
	{8'd86,8'd231} : s = 317;
	{8'd86,8'd232} : s = 318;
	{8'd86,8'd233} : s = 319;
	{8'd86,8'd234} : s = 320;
	{8'd86,8'd235} : s = 321;
	{8'd86,8'd236} : s = 322;
	{8'd86,8'd237} : s = 323;
	{8'd86,8'd238} : s = 324;
	{8'd86,8'd239} : s = 325;
	{8'd86,8'd240} : s = 326;
	{8'd86,8'd241} : s = 327;
	{8'd86,8'd242} : s = 328;
	{8'd86,8'd243} : s = 329;
	{8'd86,8'd244} : s = 330;
	{8'd86,8'd245} : s = 331;
	{8'd86,8'd246} : s = 332;
	{8'd86,8'd247} : s = 333;
	{8'd86,8'd248} : s = 334;
	{8'd86,8'd249} : s = 335;
	{8'd86,8'd250} : s = 336;
	{8'd86,8'd251} : s = 337;
	{8'd86,8'd252} : s = 338;
	{8'd86,8'd253} : s = 339;
	{8'd86,8'd254} : s = 340;
	{8'd86,8'd255} : s = 341;
	{8'd87,8'd0} : s = 87;
	{8'd87,8'd1} : s = 88;
	{8'd87,8'd2} : s = 89;
	{8'd87,8'd3} : s = 90;
	{8'd87,8'd4} : s = 91;
	{8'd87,8'd5} : s = 92;
	{8'd87,8'd6} : s = 93;
	{8'd87,8'd7} : s = 94;
	{8'd87,8'd8} : s = 95;
	{8'd87,8'd9} : s = 96;
	{8'd87,8'd10} : s = 97;
	{8'd87,8'd11} : s = 98;
	{8'd87,8'd12} : s = 99;
	{8'd87,8'd13} : s = 100;
	{8'd87,8'd14} : s = 101;
	{8'd87,8'd15} : s = 102;
	{8'd87,8'd16} : s = 103;
	{8'd87,8'd17} : s = 104;
	{8'd87,8'd18} : s = 105;
	{8'd87,8'd19} : s = 106;
	{8'd87,8'd20} : s = 107;
	{8'd87,8'd21} : s = 108;
	{8'd87,8'd22} : s = 109;
	{8'd87,8'd23} : s = 110;
	{8'd87,8'd24} : s = 111;
	{8'd87,8'd25} : s = 112;
	{8'd87,8'd26} : s = 113;
	{8'd87,8'd27} : s = 114;
	{8'd87,8'd28} : s = 115;
	{8'd87,8'd29} : s = 116;
	{8'd87,8'd30} : s = 117;
	{8'd87,8'd31} : s = 118;
	{8'd87,8'd32} : s = 119;
	{8'd87,8'd33} : s = 120;
	{8'd87,8'd34} : s = 121;
	{8'd87,8'd35} : s = 122;
	{8'd87,8'd36} : s = 123;
	{8'd87,8'd37} : s = 124;
	{8'd87,8'd38} : s = 125;
	{8'd87,8'd39} : s = 126;
	{8'd87,8'd40} : s = 127;
	{8'd87,8'd41} : s = 128;
	{8'd87,8'd42} : s = 129;
	{8'd87,8'd43} : s = 130;
	{8'd87,8'd44} : s = 131;
	{8'd87,8'd45} : s = 132;
	{8'd87,8'd46} : s = 133;
	{8'd87,8'd47} : s = 134;
	{8'd87,8'd48} : s = 135;
	{8'd87,8'd49} : s = 136;
	{8'd87,8'd50} : s = 137;
	{8'd87,8'd51} : s = 138;
	{8'd87,8'd52} : s = 139;
	{8'd87,8'd53} : s = 140;
	{8'd87,8'd54} : s = 141;
	{8'd87,8'd55} : s = 142;
	{8'd87,8'd56} : s = 143;
	{8'd87,8'd57} : s = 144;
	{8'd87,8'd58} : s = 145;
	{8'd87,8'd59} : s = 146;
	{8'd87,8'd60} : s = 147;
	{8'd87,8'd61} : s = 148;
	{8'd87,8'd62} : s = 149;
	{8'd87,8'd63} : s = 150;
	{8'd87,8'd64} : s = 151;
	{8'd87,8'd65} : s = 152;
	{8'd87,8'd66} : s = 153;
	{8'd87,8'd67} : s = 154;
	{8'd87,8'd68} : s = 155;
	{8'd87,8'd69} : s = 156;
	{8'd87,8'd70} : s = 157;
	{8'd87,8'd71} : s = 158;
	{8'd87,8'd72} : s = 159;
	{8'd87,8'd73} : s = 160;
	{8'd87,8'd74} : s = 161;
	{8'd87,8'd75} : s = 162;
	{8'd87,8'd76} : s = 163;
	{8'd87,8'd77} : s = 164;
	{8'd87,8'd78} : s = 165;
	{8'd87,8'd79} : s = 166;
	{8'd87,8'd80} : s = 167;
	{8'd87,8'd81} : s = 168;
	{8'd87,8'd82} : s = 169;
	{8'd87,8'd83} : s = 170;
	{8'd87,8'd84} : s = 171;
	{8'd87,8'd85} : s = 172;
	{8'd87,8'd86} : s = 173;
	{8'd87,8'd87} : s = 174;
	{8'd87,8'd88} : s = 175;
	{8'd87,8'd89} : s = 176;
	{8'd87,8'd90} : s = 177;
	{8'd87,8'd91} : s = 178;
	{8'd87,8'd92} : s = 179;
	{8'd87,8'd93} : s = 180;
	{8'd87,8'd94} : s = 181;
	{8'd87,8'd95} : s = 182;
	{8'd87,8'd96} : s = 183;
	{8'd87,8'd97} : s = 184;
	{8'd87,8'd98} : s = 185;
	{8'd87,8'd99} : s = 186;
	{8'd87,8'd100} : s = 187;
	{8'd87,8'd101} : s = 188;
	{8'd87,8'd102} : s = 189;
	{8'd87,8'd103} : s = 190;
	{8'd87,8'd104} : s = 191;
	{8'd87,8'd105} : s = 192;
	{8'd87,8'd106} : s = 193;
	{8'd87,8'd107} : s = 194;
	{8'd87,8'd108} : s = 195;
	{8'd87,8'd109} : s = 196;
	{8'd87,8'd110} : s = 197;
	{8'd87,8'd111} : s = 198;
	{8'd87,8'd112} : s = 199;
	{8'd87,8'd113} : s = 200;
	{8'd87,8'd114} : s = 201;
	{8'd87,8'd115} : s = 202;
	{8'd87,8'd116} : s = 203;
	{8'd87,8'd117} : s = 204;
	{8'd87,8'd118} : s = 205;
	{8'd87,8'd119} : s = 206;
	{8'd87,8'd120} : s = 207;
	{8'd87,8'd121} : s = 208;
	{8'd87,8'd122} : s = 209;
	{8'd87,8'd123} : s = 210;
	{8'd87,8'd124} : s = 211;
	{8'd87,8'd125} : s = 212;
	{8'd87,8'd126} : s = 213;
	{8'd87,8'd127} : s = 214;
	{8'd87,8'd128} : s = 215;
	{8'd87,8'd129} : s = 216;
	{8'd87,8'd130} : s = 217;
	{8'd87,8'd131} : s = 218;
	{8'd87,8'd132} : s = 219;
	{8'd87,8'd133} : s = 220;
	{8'd87,8'd134} : s = 221;
	{8'd87,8'd135} : s = 222;
	{8'd87,8'd136} : s = 223;
	{8'd87,8'd137} : s = 224;
	{8'd87,8'd138} : s = 225;
	{8'd87,8'd139} : s = 226;
	{8'd87,8'd140} : s = 227;
	{8'd87,8'd141} : s = 228;
	{8'd87,8'd142} : s = 229;
	{8'd87,8'd143} : s = 230;
	{8'd87,8'd144} : s = 231;
	{8'd87,8'd145} : s = 232;
	{8'd87,8'd146} : s = 233;
	{8'd87,8'd147} : s = 234;
	{8'd87,8'd148} : s = 235;
	{8'd87,8'd149} : s = 236;
	{8'd87,8'd150} : s = 237;
	{8'd87,8'd151} : s = 238;
	{8'd87,8'd152} : s = 239;
	{8'd87,8'd153} : s = 240;
	{8'd87,8'd154} : s = 241;
	{8'd87,8'd155} : s = 242;
	{8'd87,8'd156} : s = 243;
	{8'd87,8'd157} : s = 244;
	{8'd87,8'd158} : s = 245;
	{8'd87,8'd159} : s = 246;
	{8'd87,8'd160} : s = 247;
	{8'd87,8'd161} : s = 248;
	{8'd87,8'd162} : s = 249;
	{8'd87,8'd163} : s = 250;
	{8'd87,8'd164} : s = 251;
	{8'd87,8'd165} : s = 252;
	{8'd87,8'd166} : s = 253;
	{8'd87,8'd167} : s = 254;
	{8'd87,8'd168} : s = 255;
	{8'd87,8'd169} : s = 256;
	{8'd87,8'd170} : s = 257;
	{8'd87,8'd171} : s = 258;
	{8'd87,8'd172} : s = 259;
	{8'd87,8'd173} : s = 260;
	{8'd87,8'd174} : s = 261;
	{8'd87,8'd175} : s = 262;
	{8'd87,8'd176} : s = 263;
	{8'd87,8'd177} : s = 264;
	{8'd87,8'd178} : s = 265;
	{8'd87,8'd179} : s = 266;
	{8'd87,8'd180} : s = 267;
	{8'd87,8'd181} : s = 268;
	{8'd87,8'd182} : s = 269;
	{8'd87,8'd183} : s = 270;
	{8'd87,8'd184} : s = 271;
	{8'd87,8'd185} : s = 272;
	{8'd87,8'd186} : s = 273;
	{8'd87,8'd187} : s = 274;
	{8'd87,8'd188} : s = 275;
	{8'd87,8'd189} : s = 276;
	{8'd87,8'd190} : s = 277;
	{8'd87,8'd191} : s = 278;
	{8'd87,8'd192} : s = 279;
	{8'd87,8'd193} : s = 280;
	{8'd87,8'd194} : s = 281;
	{8'd87,8'd195} : s = 282;
	{8'd87,8'd196} : s = 283;
	{8'd87,8'd197} : s = 284;
	{8'd87,8'd198} : s = 285;
	{8'd87,8'd199} : s = 286;
	{8'd87,8'd200} : s = 287;
	{8'd87,8'd201} : s = 288;
	{8'd87,8'd202} : s = 289;
	{8'd87,8'd203} : s = 290;
	{8'd87,8'd204} : s = 291;
	{8'd87,8'd205} : s = 292;
	{8'd87,8'd206} : s = 293;
	{8'd87,8'd207} : s = 294;
	{8'd87,8'd208} : s = 295;
	{8'd87,8'd209} : s = 296;
	{8'd87,8'd210} : s = 297;
	{8'd87,8'd211} : s = 298;
	{8'd87,8'd212} : s = 299;
	{8'd87,8'd213} : s = 300;
	{8'd87,8'd214} : s = 301;
	{8'd87,8'd215} : s = 302;
	{8'd87,8'd216} : s = 303;
	{8'd87,8'd217} : s = 304;
	{8'd87,8'd218} : s = 305;
	{8'd87,8'd219} : s = 306;
	{8'd87,8'd220} : s = 307;
	{8'd87,8'd221} : s = 308;
	{8'd87,8'd222} : s = 309;
	{8'd87,8'd223} : s = 310;
	{8'd87,8'd224} : s = 311;
	{8'd87,8'd225} : s = 312;
	{8'd87,8'd226} : s = 313;
	{8'd87,8'd227} : s = 314;
	{8'd87,8'd228} : s = 315;
	{8'd87,8'd229} : s = 316;
	{8'd87,8'd230} : s = 317;
	{8'd87,8'd231} : s = 318;
	{8'd87,8'd232} : s = 319;
	{8'd87,8'd233} : s = 320;
	{8'd87,8'd234} : s = 321;
	{8'd87,8'd235} : s = 322;
	{8'd87,8'd236} : s = 323;
	{8'd87,8'd237} : s = 324;
	{8'd87,8'd238} : s = 325;
	{8'd87,8'd239} : s = 326;
	{8'd87,8'd240} : s = 327;
	{8'd87,8'd241} : s = 328;
	{8'd87,8'd242} : s = 329;
	{8'd87,8'd243} : s = 330;
	{8'd87,8'd244} : s = 331;
	{8'd87,8'd245} : s = 332;
	{8'd87,8'd246} : s = 333;
	{8'd87,8'd247} : s = 334;
	{8'd87,8'd248} : s = 335;
	{8'd87,8'd249} : s = 336;
	{8'd87,8'd250} : s = 337;
	{8'd87,8'd251} : s = 338;
	{8'd87,8'd252} : s = 339;
	{8'd87,8'd253} : s = 340;
	{8'd87,8'd254} : s = 341;
	{8'd87,8'd255} : s = 342;
	{8'd88,8'd0} : s = 88;
	{8'd88,8'd1} : s = 89;
	{8'd88,8'd2} : s = 90;
	{8'd88,8'd3} : s = 91;
	{8'd88,8'd4} : s = 92;
	{8'd88,8'd5} : s = 93;
	{8'd88,8'd6} : s = 94;
	{8'd88,8'd7} : s = 95;
	{8'd88,8'd8} : s = 96;
	{8'd88,8'd9} : s = 97;
	{8'd88,8'd10} : s = 98;
	{8'd88,8'd11} : s = 99;
	{8'd88,8'd12} : s = 100;
	{8'd88,8'd13} : s = 101;
	{8'd88,8'd14} : s = 102;
	{8'd88,8'd15} : s = 103;
	{8'd88,8'd16} : s = 104;
	{8'd88,8'd17} : s = 105;
	{8'd88,8'd18} : s = 106;
	{8'd88,8'd19} : s = 107;
	{8'd88,8'd20} : s = 108;
	{8'd88,8'd21} : s = 109;
	{8'd88,8'd22} : s = 110;
	{8'd88,8'd23} : s = 111;
	{8'd88,8'd24} : s = 112;
	{8'd88,8'd25} : s = 113;
	{8'd88,8'd26} : s = 114;
	{8'd88,8'd27} : s = 115;
	{8'd88,8'd28} : s = 116;
	{8'd88,8'd29} : s = 117;
	{8'd88,8'd30} : s = 118;
	{8'd88,8'd31} : s = 119;
	{8'd88,8'd32} : s = 120;
	{8'd88,8'd33} : s = 121;
	{8'd88,8'd34} : s = 122;
	{8'd88,8'd35} : s = 123;
	{8'd88,8'd36} : s = 124;
	{8'd88,8'd37} : s = 125;
	{8'd88,8'd38} : s = 126;
	{8'd88,8'd39} : s = 127;
	{8'd88,8'd40} : s = 128;
	{8'd88,8'd41} : s = 129;
	{8'd88,8'd42} : s = 130;
	{8'd88,8'd43} : s = 131;
	{8'd88,8'd44} : s = 132;
	{8'd88,8'd45} : s = 133;
	{8'd88,8'd46} : s = 134;
	{8'd88,8'd47} : s = 135;
	{8'd88,8'd48} : s = 136;
	{8'd88,8'd49} : s = 137;
	{8'd88,8'd50} : s = 138;
	{8'd88,8'd51} : s = 139;
	{8'd88,8'd52} : s = 140;
	{8'd88,8'd53} : s = 141;
	{8'd88,8'd54} : s = 142;
	{8'd88,8'd55} : s = 143;
	{8'd88,8'd56} : s = 144;
	{8'd88,8'd57} : s = 145;
	{8'd88,8'd58} : s = 146;
	{8'd88,8'd59} : s = 147;
	{8'd88,8'd60} : s = 148;
	{8'd88,8'd61} : s = 149;
	{8'd88,8'd62} : s = 150;
	{8'd88,8'd63} : s = 151;
	{8'd88,8'd64} : s = 152;
	{8'd88,8'd65} : s = 153;
	{8'd88,8'd66} : s = 154;
	{8'd88,8'd67} : s = 155;
	{8'd88,8'd68} : s = 156;
	{8'd88,8'd69} : s = 157;
	{8'd88,8'd70} : s = 158;
	{8'd88,8'd71} : s = 159;
	{8'd88,8'd72} : s = 160;
	{8'd88,8'd73} : s = 161;
	{8'd88,8'd74} : s = 162;
	{8'd88,8'd75} : s = 163;
	{8'd88,8'd76} : s = 164;
	{8'd88,8'd77} : s = 165;
	{8'd88,8'd78} : s = 166;
	{8'd88,8'd79} : s = 167;
	{8'd88,8'd80} : s = 168;
	{8'd88,8'd81} : s = 169;
	{8'd88,8'd82} : s = 170;
	{8'd88,8'd83} : s = 171;
	{8'd88,8'd84} : s = 172;
	{8'd88,8'd85} : s = 173;
	{8'd88,8'd86} : s = 174;
	{8'd88,8'd87} : s = 175;
	{8'd88,8'd88} : s = 176;
	{8'd88,8'd89} : s = 177;
	{8'd88,8'd90} : s = 178;
	{8'd88,8'd91} : s = 179;
	{8'd88,8'd92} : s = 180;
	{8'd88,8'd93} : s = 181;
	{8'd88,8'd94} : s = 182;
	{8'd88,8'd95} : s = 183;
	{8'd88,8'd96} : s = 184;
	{8'd88,8'd97} : s = 185;
	{8'd88,8'd98} : s = 186;
	{8'd88,8'd99} : s = 187;
	{8'd88,8'd100} : s = 188;
	{8'd88,8'd101} : s = 189;
	{8'd88,8'd102} : s = 190;
	{8'd88,8'd103} : s = 191;
	{8'd88,8'd104} : s = 192;
	{8'd88,8'd105} : s = 193;
	{8'd88,8'd106} : s = 194;
	{8'd88,8'd107} : s = 195;
	{8'd88,8'd108} : s = 196;
	{8'd88,8'd109} : s = 197;
	{8'd88,8'd110} : s = 198;
	{8'd88,8'd111} : s = 199;
	{8'd88,8'd112} : s = 200;
	{8'd88,8'd113} : s = 201;
	{8'd88,8'd114} : s = 202;
	{8'd88,8'd115} : s = 203;
	{8'd88,8'd116} : s = 204;
	{8'd88,8'd117} : s = 205;
	{8'd88,8'd118} : s = 206;
	{8'd88,8'd119} : s = 207;
	{8'd88,8'd120} : s = 208;
	{8'd88,8'd121} : s = 209;
	{8'd88,8'd122} : s = 210;
	{8'd88,8'd123} : s = 211;
	{8'd88,8'd124} : s = 212;
	{8'd88,8'd125} : s = 213;
	{8'd88,8'd126} : s = 214;
	{8'd88,8'd127} : s = 215;
	{8'd88,8'd128} : s = 216;
	{8'd88,8'd129} : s = 217;
	{8'd88,8'd130} : s = 218;
	{8'd88,8'd131} : s = 219;
	{8'd88,8'd132} : s = 220;
	{8'd88,8'd133} : s = 221;
	{8'd88,8'd134} : s = 222;
	{8'd88,8'd135} : s = 223;
	{8'd88,8'd136} : s = 224;
	{8'd88,8'd137} : s = 225;
	{8'd88,8'd138} : s = 226;
	{8'd88,8'd139} : s = 227;
	{8'd88,8'd140} : s = 228;
	{8'd88,8'd141} : s = 229;
	{8'd88,8'd142} : s = 230;
	{8'd88,8'd143} : s = 231;
	{8'd88,8'd144} : s = 232;
	{8'd88,8'd145} : s = 233;
	{8'd88,8'd146} : s = 234;
	{8'd88,8'd147} : s = 235;
	{8'd88,8'd148} : s = 236;
	{8'd88,8'd149} : s = 237;
	{8'd88,8'd150} : s = 238;
	{8'd88,8'd151} : s = 239;
	{8'd88,8'd152} : s = 240;
	{8'd88,8'd153} : s = 241;
	{8'd88,8'd154} : s = 242;
	{8'd88,8'd155} : s = 243;
	{8'd88,8'd156} : s = 244;
	{8'd88,8'd157} : s = 245;
	{8'd88,8'd158} : s = 246;
	{8'd88,8'd159} : s = 247;
	{8'd88,8'd160} : s = 248;
	{8'd88,8'd161} : s = 249;
	{8'd88,8'd162} : s = 250;
	{8'd88,8'd163} : s = 251;
	{8'd88,8'd164} : s = 252;
	{8'd88,8'd165} : s = 253;
	{8'd88,8'd166} : s = 254;
	{8'd88,8'd167} : s = 255;
	{8'd88,8'd168} : s = 256;
	{8'd88,8'd169} : s = 257;
	{8'd88,8'd170} : s = 258;
	{8'd88,8'd171} : s = 259;
	{8'd88,8'd172} : s = 260;
	{8'd88,8'd173} : s = 261;
	{8'd88,8'd174} : s = 262;
	{8'd88,8'd175} : s = 263;
	{8'd88,8'd176} : s = 264;
	{8'd88,8'd177} : s = 265;
	{8'd88,8'd178} : s = 266;
	{8'd88,8'd179} : s = 267;
	{8'd88,8'd180} : s = 268;
	{8'd88,8'd181} : s = 269;
	{8'd88,8'd182} : s = 270;
	{8'd88,8'd183} : s = 271;
	{8'd88,8'd184} : s = 272;
	{8'd88,8'd185} : s = 273;
	{8'd88,8'd186} : s = 274;
	{8'd88,8'd187} : s = 275;
	{8'd88,8'd188} : s = 276;
	{8'd88,8'd189} : s = 277;
	{8'd88,8'd190} : s = 278;
	{8'd88,8'd191} : s = 279;
	{8'd88,8'd192} : s = 280;
	{8'd88,8'd193} : s = 281;
	{8'd88,8'd194} : s = 282;
	{8'd88,8'd195} : s = 283;
	{8'd88,8'd196} : s = 284;
	{8'd88,8'd197} : s = 285;
	{8'd88,8'd198} : s = 286;
	{8'd88,8'd199} : s = 287;
	{8'd88,8'd200} : s = 288;
	{8'd88,8'd201} : s = 289;
	{8'd88,8'd202} : s = 290;
	{8'd88,8'd203} : s = 291;
	{8'd88,8'd204} : s = 292;
	{8'd88,8'd205} : s = 293;
	{8'd88,8'd206} : s = 294;
	{8'd88,8'd207} : s = 295;
	{8'd88,8'd208} : s = 296;
	{8'd88,8'd209} : s = 297;
	{8'd88,8'd210} : s = 298;
	{8'd88,8'd211} : s = 299;
	{8'd88,8'd212} : s = 300;
	{8'd88,8'd213} : s = 301;
	{8'd88,8'd214} : s = 302;
	{8'd88,8'd215} : s = 303;
	{8'd88,8'd216} : s = 304;
	{8'd88,8'd217} : s = 305;
	{8'd88,8'd218} : s = 306;
	{8'd88,8'd219} : s = 307;
	{8'd88,8'd220} : s = 308;
	{8'd88,8'd221} : s = 309;
	{8'd88,8'd222} : s = 310;
	{8'd88,8'd223} : s = 311;
	{8'd88,8'd224} : s = 312;
	{8'd88,8'd225} : s = 313;
	{8'd88,8'd226} : s = 314;
	{8'd88,8'd227} : s = 315;
	{8'd88,8'd228} : s = 316;
	{8'd88,8'd229} : s = 317;
	{8'd88,8'd230} : s = 318;
	{8'd88,8'd231} : s = 319;
	{8'd88,8'd232} : s = 320;
	{8'd88,8'd233} : s = 321;
	{8'd88,8'd234} : s = 322;
	{8'd88,8'd235} : s = 323;
	{8'd88,8'd236} : s = 324;
	{8'd88,8'd237} : s = 325;
	{8'd88,8'd238} : s = 326;
	{8'd88,8'd239} : s = 327;
	{8'd88,8'd240} : s = 328;
	{8'd88,8'd241} : s = 329;
	{8'd88,8'd242} : s = 330;
	{8'd88,8'd243} : s = 331;
	{8'd88,8'd244} : s = 332;
	{8'd88,8'd245} : s = 333;
	{8'd88,8'd246} : s = 334;
	{8'd88,8'd247} : s = 335;
	{8'd88,8'd248} : s = 336;
	{8'd88,8'd249} : s = 337;
	{8'd88,8'd250} : s = 338;
	{8'd88,8'd251} : s = 339;
	{8'd88,8'd252} : s = 340;
	{8'd88,8'd253} : s = 341;
	{8'd88,8'd254} : s = 342;
	{8'd88,8'd255} : s = 343;
	{8'd89,8'd0} : s = 89;
	{8'd89,8'd1} : s = 90;
	{8'd89,8'd2} : s = 91;
	{8'd89,8'd3} : s = 92;
	{8'd89,8'd4} : s = 93;
	{8'd89,8'd5} : s = 94;
	{8'd89,8'd6} : s = 95;
	{8'd89,8'd7} : s = 96;
	{8'd89,8'd8} : s = 97;
	{8'd89,8'd9} : s = 98;
	{8'd89,8'd10} : s = 99;
	{8'd89,8'd11} : s = 100;
	{8'd89,8'd12} : s = 101;
	{8'd89,8'd13} : s = 102;
	{8'd89,8'd14} : s = 103;
	{8'd89,8'd15} : s = 104;
	{8'd89,8'd16} : s = 105;
	{8'd89,8'd17} : s = 106;
	{8'd89,8'd18} : s = 107;
	{8'd89,8'd19} : s = 108;
	{8'd89,8'd20} : s = 109;
	{8'd89,8'd21} : s = 110;
	{8'd89,8'd22} : s = 111;
	{8'd89,8'd23} : s = 112;
	{8'd89,8'd24} : s = 113;
	{8'd89,8'd25} : s = 114;
	{8'd89,8'd26} : s = 115;
	{8'd89,8'd27} : s = 116;
	{8'd89,8'd28} : s = 117;
	{8'd89,8'd29} : s = 118;
	{8'd89,8'd30} : s = 119;
	{8'd89,8'd31} : s = 120;
	{8'd89,8'd32} : s = 121;
	{8'd89,8'd33} : s = 122;
	{8'd89,8'd34} : s = 123;
	{8'd89,8'd35} : s = 124;
	{8'd89,8'd36} : s = 125;
	{8'd89,8'd37} : s = 126;
	{8'd89,8'd38} : s = 127;
	{8'd89,8'd39} : s = 128;
	{8'd89,8'd40} : s = 129;
	{8'd89,8'd41} : s = 130;
	{8'd89,8'd42} : s = 131;
	{8'd89,8'd43} : s = 132;
	{8'd89,8'd44} : s = 133;
	{8'd89,8'd45} : s = 134;
	{8'd89,8'd46} : s = 135;
	{8'd89,8'd47} : s = 136;
	{8'd89,8'd48} : s = 137;
	{8'd89,8'd49} : s = 138;
	{8'd89,8'd50} : s = 139;
	{8'd89,8'd51} : s = 140;
	{8'd89,8'd52} : s = 141;
	{8'd89,8'd53} : s = 142;
	{8'd89,8'd54} : s = 143;
	{8'd89,8'd55} : s = 144;
	{8'd89,8'd56} : s = 145;
	{8'd89,8'd57} : s = 146;
	{8'd89,8'd58} : s = 147;
	{8'd89,8'd59} : s = 148;
	{8'd89,8'd60} : s = 149;
	{8'd89,8'd61} : s = 150;
	{8'd89,8'd62} : s = 151;
	{8'd89,8'd63} : s = 152;
	{8'd89,8'd64} : s = 153;
	{8'd89,8'd65} : s = 154;
	{8'd89,8'd66} : s = 155;
	{8'd89,8'd67} : s = 156;
	{8'd89,8'd68} : s = 157;
	{8'd89,8'd69} : s = 158;
	{8'd89,8'd70} : s = 159;
	{8'd89,8'd71} : s = 160;
	{8'd89,8'd72} : s = 161;
	{8'd89,8'd73} : s = 162;
	{8'd89,8'd74} : s = 163;
	{8'd89,8'd75} : s = 164;
	{8'd89,8'd76} : s = 165;
	{8'd89,8'd77} : s = 166;
	{8'd89,8'd78} : s = 167;
	{8'd89,8'd79} : s = 168;
	{8'd89,8'd80} : s = 169;
	{8'd89,8'd81} : s = 170;
	{8'd89,8'd82} : s = 171;
	{8'd89,8'd83} : s = 172;
	{8'd89,8'd84} : s = 173;
	{8'd89,8'd85} : s = 174;
	{8'd89,8'd86} : s = 175;
	{8'd89,8'd87} : s = 176;
	{8'd89,8'd88} : s = 177;
	{8'd89,8'd89} : s = 178;
	{8'd89,8'd90} : s = 179;
	{8'd89,8'd91} : s = 180;
	{8'd89,8'd92} : s = 181;
	{8'd89,8'd93} : s = 182;
	{8'd89,8'd94} : s = 183;
	{8'd89,8'd95} : s = 184;
	{8'd89,8'd96} : s = 185;
	{8'd89,8'd97} : s = 186;
	{8'd89,8'd98} : s = 187;
	{8'd89,8'd99} : s = 188;
	{8'd89,8'd100} : s = 189;
	{8'd89,8'd101} : s = 190;
	{8'd89,8'd102} : s = 191;
	{8'd89,8'd103} : s = 192;
	{8'd89,8'd104} : s = 193;
	{8'd89,8'd105} : s = 194;
	{8'd89,8'd106} : s = 195;
	{8'd89,8'd107} : s = 196;
	{8'd89,8'd108} : s = 197;
	{8'd89,8'd109} : s = 198;
	{8'd89,8'd110} : s = 199;
	{8'd89,8'd111} : s = 200;
	{8'd89,8'd112} : s = 201;
	{8'd89,8'd113} : s = 202;
	{8'd89,8'd114} : s = 203;
	{8'd89,8'd115} : s = 204;
	{8'd89,8'd116} : s = 205;
	{8'd89,8'd117} : s = 206;
	{8'd89,8'd118} : s = 207;
	{8'd89,8'd119} : s = 208;
	{8'd89,8'd120} : s = 209;
	{8'd89,8'd121} : s = 210;
	{8'd89,8'd122} : s = 211;
	{8'd89,8'd123} : s = 212;
	{8'd89,8'd124} : s = 213;
	{8'd89,8'd125} : s = 214;
	{8'd89,8'd126} : s = 215;
	{8'd89,8'd127} : s = 216;
	{8'd89,8'd128} : s = 217;
	{8'd89,8'd129} : s = 218;
	{8'd89,8'd130} : s = 219;
	{8'd89,8'd131} : s = 220;
	{8'd89,8'd132} : s = 221;
	{8'd89,8'd133} : s = 222;
	{8'd89,8'd134} : s = 223;
	{8'd89,8'd135} : s = 224;
	{8'd89,8'd136} : s = 225;
	{8'd89,8'd137} : s = 226;
	{8'd89,8'd138} : s = 227;
	{8'd89,8'd139} : s = 228;
	{8'd89,8'd140} : s = 229;
	{8'd89,8'd141} : s = 230;
	{8'd89,8'd142} : s = 231;
	{8'd89,8'd143} : s = 232;
	{8'd89,8'd144} : s = 233;
	{8'd89,8'd145} : s = 234;
	{8'd89,8'd146} : s = 235;
	{8'd89,8'd147} : s = 236;
	{8'd89,8'd148} : s = 237;
	{8'd89,8'd149} : s = 238;
	{8'd89,8'd150} : s = 239;
	{8'd89,8'd151} : s = 240;
	{8'd89,8'd152} : s = 241;
	{8'd89,8'd153} : s = 242;
	{8'd89,8'd154} : s = 243;
	{8'd89,8'd155} : s = 244;
	{8'd89,8'd156} : s = 245;
	{8'd89,8'd157} : s = 246;
	{8'd89,8'd158} : s = 247;
	{8'd89,8'd159} : s = 248;
	{8'd89,8'd160} : s = 249;
	{8'd89,8'd161} : s = 250;
	{8'd89,8'd162} : s = 251;
	{8'd89,8'd163} : s = 252;
	{8'd89,8'd164} : s = 253;
	{8'd89,8'd165} : s = 254;
	{8'd89,8'd166} : s = 255;
	{8'd89,8'd167} : s = 256;
	{8'd89,8'd168} : s = 257;
	{8'd89,8'd169} : s = 258;
	{8'd89,8'd170} : s = 259;
	{8'd89,8'd171} : s = 260;
	{8'd89,8'd172} : s = 261;
	{8'd89,8'd173} : s = 262;
	{8'd89,8'd174} : s = 263;
	{8'd89,8'd175} : s = 264;
	{8'd89,8'd176} : s = 265;
	{8'd89,8'd177} : s = 266;
	{8'd89,8'd178} : s = 267;
	{8'd89,8'd179} : s = 268;
	{8'd89,8'd180} : s = 269;
	{8'd89,8'd181} : s = 270;
	{8'd89,8'd182} : s = 271;
	{8'd89,8'd183} : s = 272;
	{8'd89,8'd184} : s = 273;
	{8'd89,8'd185} : s = 274;
	{8'd89,8'd186} : s = 275;
	{8'd89,8'd187} : s = 276;
	{8'd89,8'd188} : s = 277;
	{8'd89,8'd189} : s = 278;
	{8'd89,8'd190} : s = 279;
	{8'd89,8'd191} : s = 280;
	{8'd89,8'd192} : s = 281;
	{8'd89,8'd193} : s = 282;
	{8'd89,8'd194} : s = 283;
	{8'd89,8'd195} : s = 284;
	{8'd89,8'd196} : s = 285;
	{8'd89,8'd197} : s = 286;
	{8'd89,8'd198} : s = 287;
	{8'd89,8'd199} : s = 288;
	{8'd89,8'd200} : s = 289;
	{8'd89,8'd201} : s = 290;
	{8'd89,8'd202} : s = 291;
	{8'd89,8'd203} : s = 292;
	{8'd89,8'd204} : s = 293;
	{8'd89,8'd205} : s = 294;
	{8'd89,8'd206} : s = 295;
	{8'd89,8'd207} : s = 296;
	{8'd89,8'd208} : s = 297;
	{8'd89,8'd209} : s = 298;
	{8'd89,8'd210} : s = 299;
	{8'd89,8'd211} : s = 300;
	{8'd89,8'd212} : s = 301;
	{8'd89,8'd213} : s = 302;
	{8'd89,8'd214} : s = 303;
	{8'd89,8'd215} : s = 304;
	{8'd89,8'd216} : s = 305;
	{8'd89,8'd217} : s = 306;
	{8'd89,8'd218} : s = 307;
	{8'd89,8'd219} : s = 308;
	{8'd89,8'd220} : s = 309;
	{8'd89,8'd221} : s = 310;
	{8'd89,8'd222} : s = 311;
	{8'd89,8'd223} : s = 312;
	{8'd89,8'd224} : s = 313;
	{8'd89,8'd225} : s = 314;
	{8'd89,8'd226} : s = 315;
	{8'd89,8'd227} : s = 316;
	{8'd89,8'd228} : s = 317;
	{8'd89,8'd229} : s = 318;
	{8'd89,8'd230} : s = 319;
	{8'd89,8'd231} : s = 320;
	{8'd89,8'd232} : s = 321;
	{8'd89,8'd233} : s = 322;
	{8'd89,8'd234} : s = 323;
	{8'd89,8'd235} : s = 324;
	{8'd89,8'd236} : s = 325;
	{8'd89,8'd237} : s = 326;
	{8'd89,8'd238} : s = 327;
	{8'd89,8'd239} : s = 328;
	{8'd89,8'd240} : s = 329;
	{8'd89,8'd241} : s = 330;
	{8'd89,8'd242} : s = 331;
	{8'd89,8'd243} : s = 332;
	{8'd89,8'd244} : s = 333;
	{8'd89,8'd245} : s = 334;
	{8'd89,8'd246} : s = 335;
	{8'd89,8'd247} : s = 336;
	{8'd89,8'd248} : s = 337;
	{8'd89,8'd249} : s = 338;
	{8'd89,8'd250} : s = 339;
	{8'd89,8'd251} : s = 340;
	{8'd89,8'd252} : s = 341;
	{8'd89,8'd253} : s = 342;
	{8'd89,8'd254} : s = 343;
	{8'd89,8'd255} : s = 344;
	{8'd90,8'd0} : s = 90;
	{8'd90,8'd1} : s = 91;
	{8'd90,8'd2} : s = 92;
	{8'd90,8'd3} : s = 93;
	{8'd90,8'd4} : s = 94;
	{8'd90,8'd5} : s = 95;
	{8'd90,8'd6} : s = 96;
	{8'd90,8'd7} : s = 97;
	{8'd90,8'd8} : s = 98;
	{8'd90,8'd9} : s = 99;
	{8'd90,8'd10} : s = 100;
	{8'd90,8'd11} : s = 101;
	{8'd90,8'd12} : s = 102;
	{8'd90,8'd13} : s = 103;
	{8'd90,8'd14} : s = 104;
	{8'd90,8'd15} : s = 105;
	{8'd90,8'd16} : s = 106;
	{8'd90,8'd17} : s = 107;
	{8'd90,8'd18} : s = 108;
	{8'd90,8'd19} : s = 109;
	{8'd90,8'd20} : s = 110;
	{8'd90,8'd21} : s = 111;
	{8'd90,8'd22} : s = 112;
	{8'd90,8'd23} : s = 113;
	{8'd90,8'd24} : s = 114;
	{8'd90,8'd25} : s = 115;
	{8'd90,8'd26} : s = 116;
	{8'd90,8'd27} : s = 117;
	{8'd90,8'd28} : s = 118;
	{8'd90,8'd29} : s = 119;
	{8'd90,8'd30} : s = 120;
	{8'd90,8'd31} : s = 121;
	{8'd90,8'd32} : s = 122;
	{8'd90,8'd33} : s = 123;
	{8'd90,8'd34} : s = 124;
	{8'd90,8'd35} : s = 125;
	{8'd90,8'd36} : s = 126;
	{8'd90,8'd37} : s = 127;
	{8'd90,8'd38} : s = 128;
	{8'd90,8'd39} : s = 129;
	{8'd90,8'd40} : s = 130;
	{8'd90,8'd41} : s = 131;
	{8'd90,8'd42} : s = 132;
	{8'd90,8'd43} : s = 133;
	{8'd90,8'd44} : s = 134;
	{8'd90,8'd45} : s = 135;
	{8'd90,8'd46} : s = 136;
	{8'd90,8'd47} : s = 137;
	{8'd90,8'd48} : s = 138;
	{8'd90,8'd49} : s = 139;
	{8'd90,8'd50} : s = 140;
	{8'd90,8'd51} : s = 141;
	{8'd90,8'd52} : s = 142;
	{8'd90,8'd53} : s = 143;
	{8'd90,8'd54} : s = 144;
	{8'd90,8'd55} : s = 145;
	{8'd90,8'd56} : s = 146;
	{8'd90,8'd57} : s = 147;
	{8'd90,8'd58} : s = 148;
	{8'd90,8'd59} : s = 149;
	{8'd90,8'd60} : s = 150;
	{8'd90,8'd61} : s = 151;
	{8'd90,8'd62} : s = 152;
	{8'd90,8'd63} : s = 153;
	{8'd90,8'd64} : s = 154;
	{8'd90,8'd65} : s = 155;
	{8'd90,8'd66} : s = 156;
	{8'd90,8'd67} : s = 157;
	{8'd90,8'd68} : s = 158;
	{8'd90,8'd69} : s = 159;
	{8'd90,8'd70} : s = 160;
	{8'd90,8'd71} : s = 161;
	{8'd90,8'd72} : s = 162;
	{8'd90,8'd73} : s = 163;
	{8'd90,8'd74} : s = 164;
	{8'd90,8'd75} : s = 165;
	{8'd90,8'd76} : s = 166;
	{8'd90,8'd77} : s = 167;
	{8'd90,8'd78} : s = 168;
	{8'd90,8'd79} : s = 169;
	{8'd90,8'd80} : s = 170;
	{8'd90,8'd81} : s = 171;
	{8'd90,8'd82} : s = 172;
	{8'd90,8'd83} : s = 173;
	{8'd90,8'd84} : s = 174;
	{8'd90,8'd85} : s = 175;
	{8'd90,8'd86} : s = 176;
	{8'd90,8'd87} : s = 177;
	{8'd90,8'd88} : s = 178;
	{8'd90,8'd89} : s = 179;
	{8'd90,8'd90} : s = 180;
	{8'd90,8'd91} : s = 181;
	{8'd90,8'd92} : s = 182;
	{8'd90,8'd93} : s = 183;
	{8'd90,8'd94} : s = 184;
	{8'd90,8'd95} : s = 185;
	{8'd90,8'd96} : s = 186;
	{8'd90,8'd97} : s = 187;
	{8'd90,8'd98} : s = 188;
	{8'd90,8'd99} : s = 189;
	{8'd90,8'd100} : s = 190;
	{8'd90,8'd101} : s = 191;
	{8'd90,8'd102} : s = 192;
	{8'd90,8'd103} : s = 193;
	{8'd90,8'd104} : s = 194;
	{8'd90,8'd105} : s = 195;
	{8'd90,8'd106} : s = 196;
	{8'd90,8'd107} : s = 197;
	{8'd90,8'd108} : s = 198;
	{8'd90,8'd109} : s = 199;
	{8'd90,8'd110} : s = 200;
	{8'd90,8'd111} : s = 201;
	{8'd90,8'd112} : s = 202;
	{8'd90,8'd113} : s = 203;
	{8'd90,8'd114} : s = 204;
	{8'd90,8'd115} : s = 205;
	{8'd90,8'd116} : s = 206;
	{8'd90,8'd117} : s = 207;
	{8'd90,8'd118} : s = 208;
	{8'd90,8'd119} : s = 209;
	{8'd90,8'd120} : s = 210;
	{8'd90,8'd121} : s = 211;
	{8'd90,8'd122} : s = 212;
	{8'd90,8'd123} : s = 213;
	{8'd90,8'd124} : s = 214;
	{8'd90,8'd125} : s = 215;
	{8'd90,8'd126} : s = 216;
	{8'd90,8'd127} : s = 217;
	{8'd90,8'd128} : s = 218;
	{8'd90,8'd129} : s = 219;
	{8'd90,8'd130} : s = 220;
	{8'd90,8'd131} : s = 221;
	{8'd90,8'd132} : s = 222;
	{8'd90,8'd133} : s = 223;
	{8'd90,8'd134} : s = 224;
	{8'd90,8'd135} : s = 225;
	{8'd90,8'd136} : s = 226;
	{8'd90,8'd137} : s = 227;
	{8'd90,8'd138} : s = 228;
	{8'd90,8'd139} : s = 229;
	{8'd90,8'd140} : s = 230;
	{8'd90,8'd141} : s = 231;
	{8'd90,8'd142} : s = 232;
	{8'd90,8'd143} : s = 233;
	{8'd90,8'd144} : s = 234;
	{8'd90,8'd145} : s = 235;
	{8'd90,8'd146} : s = 236;
	{8'd90,8'd147} : s = 237;
	{8'd90,8'd148} : s = 238;
	{8'd90,8'd149} : s = 239;
	{8'd90,8'd150} : s = 240;
	{8'd90,8'd151} : s = 241;
	{8'd90,8'd152} : s = 242;
	{8'd90,8'd153} : s = 243;
	{8'd90,8'd154} : s = 244;
	{8'd90,8'd155} : s = 245;
	{8'd90,8'd156} : s = 246;
	{8'd90,8'd157} : s = 247;
	{8'd90,8'd158} : s = 248;
	{8'd90,8'd159} : s = 249;
	{8'd90,8'd160} : s = 250;
	{8'd90,8'd161} : s = 251;
	{8'd90,8'd162} : s = 252;
	{8'd90,8'd163} : s = 253;
	{8'd90,8'd164} : s = 254;
	{8'd90,8'd165} : s = 255;
	{8'd90,8'd166} : s = 256;
	{8'd90,8'd167} : s = 257;
	{8'd90,8'd168} : s = 258;
	{8'd90,8'd169} : s = 259;
	{8'd90,8'd170} : s = 260;
	{8'd90,8'd171} : s = 261;
	{8'd90,8'd172} : s = 262;
	{8'd90,8'd173} : s = 263;
	{8'd90,8'd174} : s = 264;
	{8'd90,8'd175} : s = 265;
	{8'd90,8'd176} : s = 266;
	{8'd90,8'd177} : s = 267;
	{8'd90,8'd178} : s = 268;
	{8'd90,8'd179} : s = 269;
	{8'd90,8'd180} : s = 270;
	{8'd90,8'd181} : s = 271;
	{8'd90,8'd182} : s = 272;
	{8'd90,8'd183} : s = 273;
	{8'd90,8'd184} : s = 274;
	{8'd90,8'd185} : s = 275;
	{8'd90,8'd186} : s = 276;
	{8'd90,8'd187} : s = 277;
	{8'd90,8'd188} : s = 278;
	{8'd90,8'd189} : s = 279;
	{8'd90,8'd190} : s = 280;
	{8'd90,8'd191} : s = 281;
	{8'd90,8'd192} : s = 282;
	{8'd90,8'd193} : s = 283;
	{8'd90,8'd194} : s = 284;
	{8'd90,8'd195} : s = 285;
	{8'd90,8'd196} : s = 286;
	{8'd90,8'd197} : s = 287;
	{8'd90,8'd198} : s = 288;
	{8'd90,8'd199} : s = 289;
	{8'd90,8'd200} : s = 290;
	{8'd90,8'd201} : s = 291;
	{8'd90,8'd202} : s = 292;
	{8'd90,8'd203} : s = 293;
	{8'd90,8'd204} : s = 294;
	{8'd90,8'd205} : s = 295;
	{8'd90,8'd206} : s = 296;
	{8'd90,8'd207} : s = 297;
	{8'd90,8'd208} : s = 298;
	{8'd90,8'd209} : s = 299;
	{8'd90,8'd210} : s = 300;
	{8'd90,8'd211} : s = 301;
	{8'd90,8'd212} : s = 302;
	{8'd90,8'd213} : s = 303;
	{8'd90,8'd214} : s = 304;
	{8'd90,8'd215} : s = 305;
	{8'd90,8'd216} : s = 306;
	{8'd90,8'd217} : s = 307;
	{8'd90,8'd218} : s = 308;
	{8'd90,8'd219} : s = 309;
	{8'd90,8'd220} : s = 310;
	{8'd90,8'd221} : s = 311;
	{8'd90,8'd222} : s = 312;
	{8'd90,8'd223} : s = 313;
	{8'd90,8'd224} : s = 314;
	{8'd90,8'd225} : s = 315;
	{8'd90,8'd226} : s = 316;
	{8'd90,8'd227} : s = 317;
	{8'd90,8'd228} : s = 318;
	{8'd90,8'd229} : s = 319;
	{8'd90,8'd230} : s = 320;
	{8'd90,8'd231} : s = 321;
	{8'd90,8'd232} : s = 322;
	{8'd90,8'd233} : s = 323;
	{8'd90,8'd234} : s = 324;
	{8'd90,8'd235} : s = 325;
	{8'd90,8'd236} : s = 326;
	{8'd90,8'd237} : s = 327;
	{8'd90,8'd238} : s = 328;
	{8'd90,8'd239} : s = 329;
	{8'd90,8'd240} : s = 330;
	{8'd90,8'd241} : s = 331;
	{8'd90,8'd242} : s = 332;
	{8'd90,8'd243} : s = 333;
	{8'd90,8'd244} : s = 334;
	{8'd90,8'd245} : s = 335;
	{8'd90,8'd246} : s = 336;
	{8'd90,8'd247} : s = 337;
	{8'd90,8'd248} : s = 338;
	{8'd90,8'd249} : s = 339;
	{8'd90,8'd250} : s = 340;
	{8'd90,8'd251} : s = 341;
	{8'd90,8'd252} : s = 342;
	{8'd90,8'd253} : s = 343;
	{8'd90,8'd254} : s = 344;
	{8'd90,8'd255} : s = 345;
	{8'd91,8'd0} : s = 91;
	{8'd91,8'd1} : s = 92;
	{8'd91,8'd2} : s = 93;
	{8'd91,8'd3} : s = 94;
	{8'd91,8'd4} : s = 95;
	{8'd91,8'd5} : s = 96;
	{8'd91,8'd6} : s = 97;
	{8'd91,8'd7} : s = 98;
	{8'd91,8'd8} : s = 99;
	{8'd91,8'd9} : s = 100;
	{8'd91,8'd10} : s = 101;
	{8'd91,8'd11} : s = 102;
	{8'd91,8'd12} : s = 103;
	{8'd91,8'd13} : s = 104;
	{8'd91,8'd14} : s = 105;
	{8'd91,8'd15} : s = 106;
	{8'd91,8'd16} : s = 107;
	{8'd91,8'd17} : s = 108;
	{8'd91,8'd18} : s = 109;
	{8'd91,8'd19} : s = 110;
	{8'd91,8'd20} : s = 111;
	{8'd91,8'd21} : s = 112;
	{8'd91,8'd22} : s = 113;
	{8'd91,8'd23} : s = 114;
	{8'd91,8'd24} : s = 115;
	{8'd91,8'd25} : s = 116;
	{8'd91,8'd26} : s = 117;
	{8'd91,8'd27} : s = 118;
	{8'd91,8'd28} : s = 119;
	{8'd91,8'd29} : s = 120;
	{8'd91,8'd30} : s = 121;
	{8'd91,8'd31} : s = 122;
	{8'd91,8'd32} : s = 123;
	{8'd91,8'd33} : s = 124;
	{8'd91,8'd34} : s = 125;
	{8'd91,8'd35} : s = 126;
	{8'd91,8'd36} : s = 127;
	{8'd91,8'd37} : s = 128;
	{8'd91,8'd38} : s = 129;
	{8'd91,8'd39} : s = 130;
	{8'd91,8'd40} : s = 131;
	{8'd91,8'd41} : s = 132;
	{8'd91,8'd42} : s = 133;
	{8'd91,8'd43} : s = 134;
	{8'd91,8'd44} : s = 135;
	{8'd91,8'd45} : s = 136;
	{8'd91,8'd46} : s = 137;
	{8'd91,8'd47} : s = 138;
	{8'd91,8'd48} : s = 139;
	{8'd91,8'd49} : s = 140;
	{8'd91,8'd50} : s = 141;
	{8'd91,8'd51} : s = 142;
	{8'd91,8'd52} : s = 143;
	{8'd91,8'd53} : s = 144;
	{8'd91,8'd54} : s = 145;
	{8'd91,8'd55} : s = 146;
	{8'd91,8'd56} : s = 147;
	{8'd91,8'd57} : s = 148;
	{8'd91,8'd58} : s = 149;
	{8'd91,8'd59} : s = 150;
	{8'd91,8'd60} : s = 151;
	{8'd91,8'd61} : s = 152;
	{8'd91,8'd62} : s = 153;
	{8'd91,8'd63} : s = 154;
	{8'd91,8'd64} : s = 155;
	{8'd91,8'd65} : s = 156;
	{8'd91,8'd66} : s = 157;
	{8'd91,8'd67} : s = 158;
	{8'd91,8'd68} : s = 159;
	{8'd91,8'd69} : s = 160;
	{8'd91,8'd70} : s = 161;
	{8'd91,8'd71} : s = 162;
	{8'd91,8'd72} : s = 163;
	{8'd91,8'd73} : s = 164;
	{8'd91,8'd74} : s = 165;
	{8'd91,8'd75} : s = 166;
	{8'd91,8'd76} : s = 167;
	{8'd91,8'd77} : s = 168;
	{8'd91,8'd78} : s = 169;
	{8'd91,8'd79} : s = 170;
	{8'd91,8'd80} : s = 171;
	{8'd91,8'd81} : s = 172;
	{8'd91,8'd82} : s = 173;
	{8'd91,8'd83} : s = 174;
	{8'd91,8'd84} : s = 175;
	{8'd91,8'd85} : s = 176;
	{8'd91,8'd86} : s = 177;
	{8'd91,8'd87} : s = 178;
	{8'd91,8'd88} : s = 179;
	{8'd91,8'd89} : s = 180;
	{8'd91,8'd90} : s = 181;
	{8'd91,8'd91} : s = 182;
	{8'd91,8'd92} : s = 183;
	{8'd91,8'd93} : s = 184;
	{8'd91,8'd94} : s = 185;
	{8'd91,8'd95} : s = 186;
	{8'd91,8'd96} : s = 187;
	{8'd91,8'd97} : s = 188;
	{8'd91,8'd98} : s = 189;
	{8'd91,8'd99} : s = 190;
	{8'd91,8'd100} : s = 191;
	{8'd91,8'd101} : s = 192;
	{8'd91,8'd102} : s = 193;
	{8'd91,8'd103} : s = 194;
	{8'd91,8'd104} : s = 195;
	{8'd91,8'd105} : s = 196;
	{8'd91,8'd106} : s = 197;
	{8'd91,8'd107} : s = 198;
	{8'd91,8'd108} : s = 199;
	{8'd91,8'd109} : s = 200;
	{8'd91,8'd110} : s = 201;
	{8'd91,8'd111} : s = 202;
	{8'd91,8'd112} : s = 203;
	{8'd91,8'd113} : s = 204;
	{8'd91,8'd114} : s = 205;
	{8'd91,8'd115} : s = 206;
	{8'd91,8'd116} : s = 207;
	{8'd91,8'd117} : s = 208;
	{8'd91,8'd118} : s = 209;
	{8'd91,8'd119} : s = 210;
	{8'd91,8'd120} : s = 211;
	{8'd91,8'd121} : s = 212;
	{8'd91,8'd122} : s = 213;
	{8'd91,8'd123} : s = 214;
	{8'd91,8'd124} : s = 215;
	{8'd91,8'd125} : s = 216;
	{8'd91,8'd126} : s = 217;
	{8'd91,8'd127} : s = 218;
	{8'd91,8'd128} : s = 219;
	{8'd91,8'd129} : s = 220;
	{8'd91,8'd130} : s = 221;
	{8'd91,8'd131} : s = 222;
	{8'd91,8'd132} : s = 223;
	{8'd91,8'd133} : s = 224;
	{8'd91,8'd134} : s = 225;
	{8'd91,8'd135} : s = 226;
	{8'd91,8'd136} : s = 227;
	{8'd91,8'd137} : s = 228;
	{8'd91,8'd138} : s = 229;
	{8'd91,8'd139} : s = 230;
	{8'd91,8'd140} : s = 231;
	{8'd91,8'd141} : s = 232;
	{8'd91,8'd142} : s = 233;
	{8'd91,8'd143} : s = 234;
	{8'd91,8'd144} : s = 235;
	{8'd91,8'd145} : s = 236;
	{8'd91,8'd146} : s = 237;
	{8'd91,8'd147} : s = 238;
	{8'd91,8'd148} : s = 239;
	{8'd91,8'd149} : s = 240;
	{8'd91,8'd150} : s = 241;
	{8'd91,8'd151} : s = 242;
	{8'd91,8'd152} : s = 243;
	{8'd91,8'd153} : s = 244;
	{8'd91,8'd154} : s = 245;
	{8'd91,8'd155} : s = 246;
	{8'd91,8'd156} : s = 247;
	{8'd91,8'd157} : s = 248;
	{8'd91,8'd158} : s = 249;
	{8'd91,8'd159} : s = 250;
	{8'd91,8'd160} : s = 251;
	{8'd91,8'd161} : s = 252;
	{8'd91,8'd162} : s = 253;
	{8'd91,8'd163} : s = 254;
	{8'd91,8'd164} : s = 255;
	{8'd91,8'd165} : s = 256;
	{8'd91,8'd166} : s = 257;
	{8'd91,8'd167} : s = 258;
	{8'd91,8'd168} : s = 259;
	{8'd91,8'd169} : s = 260;
	{8'd91,8'd170} : s = 261;
	{8'd91,8'd171} : s = 262;
	{8'd91,8'd172} : s = 263;
	{8'd91,8'd173} : s = 264;
	{8'd91,8'd174} : s = 265;
	{8'd91,8'd175} : s = 266;
	{8'd91,8'd176} : s = 267;
	{8'd91,8'd177} : s = 268;
	{8'd91,8'd178} : s = 269;
	{8'd91,8'd179} : s = 270;
	{8'd91,8'd180} : s = 271;
	{8'd91,8'd181} : s = 272;
	{8'd91,8'd182} : s = 273;
	{8'd91,8'd183} : s = 274;
	{8'd91,8'd184} : s = 275;
	{8'd91,8'd185} : s = 276;
	{8'd91,8'd186} : s = 277;
	{8'd91,8'd187} : s = 278;
	{8'd91,8'd188} : s = 279;
	{8'd91,8'd189} : s = 280;
	{8'd91,8'd190} : s = 281;
	{8'd91,8'd191} : s = 282;
	{8'd91,8'd192} : s = 283;
	{8'd91,8'd193} : s = 284;
	{8'd91,8'd194} : s = 285;
	{8'd91,8'd195} : s = 286;
	{8'd91,8'd196} : s = 287;
	{8'd91,8'd197} : s = 288;
	{8'd91,8'd198} : s = 289;
	{8'd91,8'd199} : s = 290;
	{8'd91,8'd200} : s = 291;
	{8'd91,8'd201} : s = 292;
	{8'd91,8'd202} : s = 293;
	{8'd91,8'd203} : s = 294;
	{8'd91,8'd204} : s = 295;
	{8'd91,8'd205} : s = 296;
	{8'd91,8'd206} : s = 297;
	{8'd91,8'd207} : s = 298;
	{8'd91,8'd208} : s = 299;
	{8'd91,8'd209} : s = 300;
	{8'd91,8'd210} : s = 301;
	{8'd91,8'd211} : s = 302;
	{8'd91,8'd212} : s = 303;
	{8'd91,8'd213} : s = 304;
	{8'd91,8'd214} : s = 305;
	{8'd91,8'd215} : s = 306;
	{8'd91,8'd216} : s = 307;
	{8'd91,8'd217} : s = 308;
	{8'd91,8'd218} : s = 309;
	{8'd91,8'd219} : s = 310;
	{8'd91,8'd220} : s = 311;
	{8'd91,8'd221} : s = 312;
	{8'd91,8'd222} : s = 313;
	{8'd91,8'd223} : s = 314;
	{8'd91,8'd224} : s = 315;
	{8'd91,8'd225} : s = 316;
	{8'd91,8'd226} : s = 317;
	{8'd91,8'd227} : s = 318;
	{8'd91,8'd228} : s = 319;
	{8'd91,8'd229} : s = 320;
	{8'd91,8'd230} : s = 321;
	{8'd91,8'd231} : s = 322;
	{8'd91,8'd232} : s = 323;
	{8'd91,8'd233} : s = 324;
	{8'd91,8'd234} : s = 325;
	{8'd91,8'd235} : s = 326;
	{8'd91,8'd236} : s = 327;
	{8'd91,8'd237} : s = 328;
	{8'd91,8'd238} : s = 329;
	{8'd91,8'd239} : s = 330;
	{8'd91,8'd240} : s = 331;
	{8'd91,8'd241} : s = 332;
	{8'd91,8'd242} : s = 333;
	{8'd91,8'd243} : s = 334;
	{8'd91,8'd244} : s = 335;
	{8'd91,8'd245} : s = 336;
	{8'd91,8'd246} : s = 337;
	{8'd91,8'd247} : s = 338;
	{8'd91,8'd248} : s = 339;
	{8'd91,8'd249} : s = 340;
	{8'd91,8'd250} : s = 341;
	{8'd91,8'd251} : s = 342;
	{8'd91,8'd252} : s = 343;
	{8'd91,8'd253} : s = 344;
	{8'd91,8'd254} : s = 345;
	{8'd91,8'd255} : s = 346;
	{8'd92,8'd0} : s = 92;
	{8'd92,8'd1} : s = 93;
	{8'd92,8'd2} : s = 94;
	{8'd92,8'd3} : s = 95;
	{8'd92,8'd4} : s = 96;
	{8'd92,8'd5} : s = 97;
	{8'd92,8'd6} : s = 98;
	{8'd92,8'd7} : s = 99;
	{8'd92,8'd8} : s = 100;
	{8'd92,8'd9} : s = 101;
	{8'd92,8'd10} : s = 102;
	{8'd92,8'd11} : s = 103;
	{8'd92,8'd12} : s = 104;
	{8'd92,8'd13} : s = 105;
	{8'd92,8'd14} : s = 106;
	{8'd92,8'd15} : s = 107;
	{8'd92,8'd16} : s = 108;
	{8'd92,8'd17} : s = 109;
	{8'd92,8'd18} : s = 110;
	{8'd92,8'd19} : s = 111;
	{8'd92,8'd20} : s = 112;
	{8'd92,8'd21} : s = 113;
	{8'd92,8'd22} : s = 114;
	{8'd92,8'd23} : s = 115;
	{8'd92,8'd24} : s = 116;
	{8'd92,8'd25} : s = 117;
	{8'd92,8'd26} : s = 118;
	{8'd92,8'd27} : s = 119;
	{8'd92,8'd28} : s = 120;
	{8'd92,8'd29} : s = 121;
	{8'd92,8'd30} : s = 122;
	{8'd92,8'd31} : s = 123;
	{8'd92,8'd32} : s = 124;
	{8'd92,8'd33} : s = 125;
	{8'd92,8'd34} : s = 126;
	{8'd92,8'd35} : s = 127;
	{8'd92,8'd36} : s = 128;
	{8'd92,8'd37} : s = 129;
	{8'd92,8'd38} : s = 130;
	{8'd92,8'd39} : s = 131;
	{8'd92,8'd40} : s = 132;
	{8'd92,8'd41} : s = 133;
	{8'd92,8'd42} : s = 134;
	{8'd92,8'd43} : s = 135;
	{8'd92,8'd44} : s = 136;
	{8'd92,8'd45} : s = 137;
	{8'd92,8'd46} : s = 138;
	{8'd92,8'd47} : s = 139;
	{8'd92,8'd48} : s = 140;
	{8'd92,8'd49} : s = 141;
	{8'd92,8'd50} : s = 142;
	{8'd92,8'd51} : s = 143;
	{8'd92,8'd52} : s = 144;
	{8'd92,8'd53} : s = 145;
	{8'd92,8'd54} : s = 146;
	{8'd92,8'd55} : s = 147;
	{8'd92,8'd56} : s = 148;
	{8'd92,8'd57} : s = 149;
	{8'd92,8'd58} : s = 150;
	{8'd92,8'd59} : s = 151;
	{8'd92,8'd60} : s = 152;
	{8'd92,8'd61} : s = 153;
	{8'd92,8'd62} : s = 154;
	{8'd92,8'd63} : s = 155;
	{8'd92,8'd64} : s = 156;
	{8'd92,8'd65} : s = 157;
	{8'd92,8'd66} : s = 158;
	{8'd92,8'd67} : s = 159;
	{8'd92,8'd68} : s = 160;
	{8'd92,8'd69} : s = 161;
	{8'd92,8'd70} : s = 162;
	{8'd92,8'd71} : s = 163;
	{8'd92,8'd72} : s = 164;
	{8'd92,8'd73} : s = 165;
	{8'd92,8'd74} : s = 166;
	{8'd92,8'd75} : s = 167;
	{8'd92,8'd76} : s = 168;
	{8'd92,8'd77} : s = 169;
	{8'd92,8'd78} : s = 170;
	{8'd92,8'd79} : s = 171;
	{8'd92,8'd80} : s = 172;
	{8'd92,8'd81} : s = 173;
	{8'd92,8'd82} : s = 174;
	{8'd92,8'd83} : s = 175;
	{8'd92,8'd84} : s = 176;
	{8'd92,8'd85} : s = 177;
	{8'd92,8'd86} : s = 178;
	{8'd92,8'd87} : s = 179;
	{8'd92,8'd88} : s = 180;
	{8'd92,8'd89} : s = 181;
	{8'd92,8'd90} : s = 182;
	{8'd92,8'd91} : s = 183;
	{8'd92,8'd92} : s = 184;
	{8'd92,8'd93} : s = 185;
	{8'd92,8'd94} : s = 186;
	{8'd92,8'd95} : s = 187;
	{8'd92,8'd96} : s = 188;
	{8'd92,8'd97} : s = 189;
	{8'd92,8'd98} : s = 190;
	{8'd92,8'd99} : s = 191;
	{8'd92,8'd100} : s = 192;
	{8'd92,8'd101} : s = 193;
	{8'd92,8'd102} : s = 194;
	{8'd92,8'd103} : s = 195;
	{8'd92,8'd104} : s = 196;
	{8'd92,8'd105} : s = 197;
	{8'd92,8'd106} : s = 198;
	{8'd92,8'd107} : s = 199;
	{8'd92,8'd108} : s = 200;
	{8'd92,8'd109} : s = 201;
	{8'd92,8'd110} : s = 202;
	{8'd92,8'd111} : s = 203;
	{8'd92,8'd112} : s = 204;
	{8'd92,8'd113} : s = 205;
	{8'd92,8'd114} : s = 206;
	{8'd92,8'd115} : s = 207;
	{8'd92,8'd116} : s = 208;
	{8'd92,8'd117} : s = 209;
	{8'd92,8'd118} : s = 210;
	{8'd92,8'd119} : s = 211;
	{8'd92,8'd120} : s = 212;
	{8'd92,8'd121} : s = 213;
	{8'd92,8'd122} : s = 214;
	{8'd92,8'd123} : s = 215;
	{8'd92,8'd124} : s = 216;
	{8'd92,8'd125} : s = 217;
	{8'd92,8'd126} : s = 218;
	{8'd92,8'd127} : s = 219;
	{8'd92,8'd128} : s = 220;
	{8'd92,8'd129} : s = 221;
	{8'd92,8'd130} : s = 222;
	{8'd92,8'd131} : s = 223;
	{8'd92,8'd132} : s = 224;
	{8'd92,8'd133} : s = 225;
	{8'd92,8'd134} : s = 226;
	{8'd92,8'd135} : s = 227;
	{8'd92,8'd136} : s = 228;
	{8'd92,8'd137} : s = 229;
	{8'd92,8'd138} : s = 230;
	{8'd92,8'd139} : s = 231;
	{8'd92,8'd140} : s = 232;
	{8'd92,8'd141} : s = 233;
	{8'd92,8'd142} : s = 234;
	{8'd92,8'd143} : s = 235;
	{8'd92,8'd144} : s = 236;
	{8'd92,8'd145} : s = 237;
	{8'd92,8'd146} : s = 238;
	{8'd92,8'd147} : s = 239;
	{8'd92,8'd148} : s = 240;
	{8'd92,8'd149} : s = 241;
	{8'd92,8'd150} : s = 242;
	{8'd92,8'd151} : s = 243;
	{8'd92,8'd152} : s = 244;
	{8'd92,8'd153} : s = 245;
	{8'd92,8'd154} : s = 246;
	{8'd92,8'd155} : s = 247;
	{8'd92,8'd156} : s = 248;
	{8'd92,8'd157} : s = 249;
	{8'd92,8'd158} : s = 250;
	{8'd92,8'd159} : s = 251;
	{8'd92,8'd160} : s = 252;
	{8'd92,8'd161} : s = 253;
	{8'd92,8'd162} : s = 254;
	{8'd92,8'd163} : s = 255;
	{8'd92,8'd164} : s = 256;
	{8'd92,8'd165} : s = 257;
	{8'd92,8'd166} : s = 258;
	{8'd92,8'd167} : s = 259;
	{8'd92,8'd168} : s = 260;
	{8'd92,8'd169} : s = 261;
	{8'd92,8'd170} : s = 262;
	{8'd92,8'd171} : s = 263;
	{8'd92,8'd172} : s = 264;
	{8'd92,8'd173} : s = 265;
	{8'd92,8'd174} : s = 266;
	{8'd92,8'd175} : s = 267;
	{8'd92,8'd176} : s = 268;
	{8'd92,8'd177} : s = 269;
	{8'd92,8'd178} : s = 270;
	{8'd92,8'd179} : s = 271;
	{8'd92,8'd180} : s = 272;
	{8'd92,8'd181} : s = 273;
	{8'd92,8'd182} : s = 274;
	{8'd92,8'd183} : s = 275;
	{8'd92,8'd184} : s = 276;
	{8'd92,8'd185} : s = 277;
	{8'd92,8'd186} : s = 278;
	{8'd92,8'd187} : s = 279;
	{8'd92,8'd188} : s = 280;
	{8'd92,8'd189} : s = 281;
	{8'd92,8'd190} : s = 282;
	{8'd92,8'd191} : s = 283;
	{8'd92,8'd192} : s = 284;
	{8'd92,8'd193} : s = 285;
	{8'd92,8'd194} : s = 286;
	{8'd92,8'd195} : s = 287;
	{8'd92,8'd196} : s = 288;
	{8'd92,8'd197} : s = 289;
	{8'd92,8'd198} : s = 290;
	{8'd92,8'd199} : s = 291;
	{8'd92,8'd200} : s = 292;
	{8'd92,8'd201} : s = 293;
	{8'd92,8'd202} : s = 294;
	{8'd92,8'd203} : s = 295;
	{8'd92,8'd204} : s = 296;
	{8'd92,8'd205} : s = 297;
	{8'd92,8'd206} : s = 298;
	{8'd92,8'd207} : s = 299;
	{8'd92,8'd208} : s = 300;
	{8'd92,8'd209} : s = 301;
	{8'd92,8'd210} : s = 302;
	{8'd92,8'd211} : s = 303;
	{8'd92,8'd212} : s = 304;
	{8'd92,8'd213} : s = 305;
	{8'd92,8'd214} : s = 306;
	{8'd92,8'd215} : s = 307;
	{8'd92,8'd216} : s = 308;
	{8'd92,8'd217} : s = 309;
	{8'd92,8'd218} : s = 310;
	{8'd92,8'd219} : s = 311;
	{8'd92,8'd220} : s = 312;
	{8'd92,8'd221} : s = 313;
	{8'd92,8'd222} : s = 314;
	{8'd92,8'd223} : s = 315;
	{8'd92,8'd224} : s = 316;
	{8'd92,8'd225} : s = 317;
	{8'd92,8'd226} : s = 318;
	{8'd92,8'd227} : s = 319;
	{8'd92,8'd228} : s = 320;
	{8'd92,8'd229} : s = 321;
	{8'd92,8'd230} : s = 322;
	{8'd92,8'd231} : s = 323;
	{8'd92,8'd232} : s = 324;
	{8'd92,8'd233} : s = 325;
	{8'd92,8'd234} : s = 326;
	{8'd92,8'd235} : s = 327;
	{8'd92,8'd236} : s = 328;
	{8'd92,8'd237} : s = 329;
	{8'd92,8'd238} : s = 330;
	{8'd92,8'd239} : s = 331;
	{8'd92,8'd240} : s = 332;
	{8'd92,8'd241} : s = 333;
	{8'd92,8'd242} : s = 334;
	{8'd92,8'd243} : s = 335;
	{8'd92,8'd244} : s = 336;
	{8'd92,8'd245} : s = 337;
	{8'd92,8'd246} : s = 338;
	{8'd92,8'd247} : s = 339;
	{8'd92,8'd248} : s = 340;
	{8'd92,8'd249} : s = 341;
	{8'd92,8'd250} : s = 342;
	{8'd92,8'd251} : s = 343;
	{8'd92,8'd252} : s = 344;
	{8'd92,8'd253} : s = 345;
	{8'd92,8'd254} : s = 346;
	{8'd92,8'd255} : s = 347;
	{8'd93,8'd0} : s = 93;
	{8'd93,8'd1} : s = 94;
	{8'd93,8'd2} : s = 95;
	{8'd93,8'd3} : s = 96;
	{8'd93,8'd4} : s = 97;
	{8'd93,8'd5} : s = 98;
	{8'd93,8'd6} : s = 99;
	{8'd93,8'd7} : s = 100;
	{8'd93,8'd8} : s = 101;
	{8'd93,8'd9} : s = 102;
	{8'd93,8'd10} : s = 103;
	{8'd93,8'd11} : s = 104;
	{8'd93,8'd12} : s = 105;
	{8'd93,8'd13} : s = 106;
	{8'd93,8'd14} : s = 107;
	{8'd93,8'd15} : s = 108;
	{8'd93,8'd16} : s = 109;
	{8'd93,8'd17} : s = 110;
	{8'd93,8'd18} : s = 111;
	{8'd93,8'd19} : s = 112;
	{8'd93,8'd20} : s = 113;
	{8'd93,8'd21} : s = 114;
	{8'd93,8'd22} : s = 115;
	{8'd93,8'd23} : s = 116;
	{8'd93,8'd24} : s = 117;
	{8'd93,8'd25} : s = 118;
	{8'd93,8'd26} : s = 119;
	{8'd93,8'd27} : s = 120;
	{8'd93,8'd28} : s = 121;
	{8'd93,8'd29} : s = 122;
	{8'd93,8'd30} : s = 123;
	{8'd93,8'd31} : s = 124;
	{8'd93,8'd32} : s = 125;
	{8'd93,8'd33} : s = 126;
	{8'd93,8'd34} : s = 127;
	{8'd93,8'd35} : s = 128;
	{8'd93,8'd36} : s = 129;
	{8'd93,8'd37} : s = 130;
	{8'd93,8'd38} : s = 131;
	{8'd93,8'd39} : s = 132;
	{8'd93,8'd40} : s = 133;
	{8'd93,8'd41} : s = 134;
	{8'd93,8'd42} : s = 135;
	{8'd93,8'd43} : s = 136;
	{8'd93,8'd44} : s = 137;
	{8'd93,8'd45} : s = 138;
	{8'd93,8'd46} : s = 139;
	{8'd93,8'd47} : s = 140;
	{8'd93,8'd48} : s = 141;
	{8'd93,8'd49} : s = 142;
	{8'd93,8'd50} : s = 143;
	{8'd93,8'd51} : s = 144;
	{8'd93,8'd52} : s = 145;
	{8'd93,8'd53} : s = 146;
	{8'd93,8'd54} : s = 147;
	{8'd93,8'd55} : s = 148;
	{8'd93,8'd56} : s = 149;
	{8'd93,8'd57} : s = 150;
	{8'd93,8'd58} : s = 151;
	{8'd93,8'd59} : s = 152;
	{8'd93,8'd60} : s = 153;
	{8'd93,8'd61} : s = 154;
	{8'd93,8'd62} : s = 155;
	{8'd93,8'd63} : s = 156;
	{8'd93,8'd64} : s = 157;
	{8'd93,8'd65} : s = 158;
	{8'd93,8'd66} : s = 159;
	{8'd93,8'd67} : s = 160;
	{8'd93,8'd68} : s = 161;
	{8'd93,8'd69} : s = 162;
	{8'd93,8'd70} : s = 163;
	{8'd93,8'd71} : s = 164;
	{8'd93,8'd72} : s = 165;
	{8'd93,8'd73} : s = 166;
	{8'd93,8'd74} : s = 167;
	{8'd93,8'd75} : s = 168;
	{8'd93,8'd76} : s = 169;
	{8'd93,8'd77} : s = 170;
	{8'd93,8'd78} : s = 171;
	{8'd93,8'd79} : s = 172;
	{8'd93,8'd80} : s = 173;
	{8'd93,8'd81} : s = 174;
	{8'd93,8'd82} : s = 175;
	{8'd93,8'd83} : s = 176;
	{8'd93,8'd84} : s = 177;
	{8'd93,8'd85} : s = 178;
	{8'd93,8'd86} : s = 179;
	{8'd93,8'd87} : s = 180;
	{8'd93,8'd88} : s = 181;
	{8'd93,8'd89} : s = 182;
	{8'd93,8'd90} : s = 183;
	{8'd93,8'd91} : s = 184;
	{8'd93,8'd92} : s = 185;
	{8'd93,8'd93} : s = 186;
	{8'd93,8'd94} : s = 187;
	{8'd93,8'd95} : s = 188;
	{8'd93,8'd96} : s = 189;
	{8'd93,8'd97} : s = 190;
	{8'd93,8'd98} : s = 191;
	{8'd93,8'd99} : s = 192;
	{8'd93,8'd100} : s = 193;
	{8'd93,8'd101} : s = 194;
	{8'd93,8'd102} : s = 195;
	{8'd93,8'd103} : s = 196;
	{8'd93,8'd104} : s = 197;
	{8'd93,8'd105} : s = 198;
	{8'd93,8'd106} : s = 199;
	{8'd93,8'd107} : s = 200;
	{8'd93,8'd108} : s = 201;
	{8'd93,8'd109} : s = 202;
	{8'd93,8'd110} : s = 203;
	{8'd93,8'd111} : s = 204;
	{8'd93,8'd112} : s = 205;
	{8'd93,8'd113} : s = 206;
	{8'd93,8'd114} : s = 207;
	{8'd93,8'd115} : s = 208;
	{8'd93,8'd116} : s = 209;
	{8'd93,8'd117} : s = 210;
	{8'd93,8'd118} : s = 211;
	{8'd93,8'd119} : s = 212;
	{8'd93,8'd120} : s = 213;
	{8'd93,8'd121} : s = 214;
	{8'd93,8'd122} : s = 215;
	{8'd93,8'd123} : s = 216;
	{8'd93,8'd124} : s = 217;
	{8'd93,8'd125} : s = 218;
	{8'd93,8'd126} : s = 219;
	{8'd93,8'd127} : s = 220;
	{8'd93,8'd128} : s = 221;
	{8'd93,8'd129} : s = 222;
	{8'd93,8'd130} : s = 223;
	{8'd93,8'd131} : s = 224;
	{8'd93,8'd132} : s = 225;
	{8'd93,8'd133} : s = 226;
	{8'd93,8'd134} : s = 227;
	{8'd93,8'd135} : s = 228;
	{8'd93,8'd136} : s = 229;
	{8'd93,8'd137} : s = 230;
	{8'd93,8'd138} : s = 231;
	{8'd93,8'd139} : s = 232;
	{8'd93,8'd140} : s = 233;
	{8'd93,8'd141} : s = 234;
	{8'd93,8'd142} : s = 235;
	{8'd93,8'd143} : s = 236;
	{8'd93,8'd144} : s = 237;
	{8'd93,8'd145} : s = 238;
	{8'd93,8'd146} : s = 239;
	{8'd93,8'd147} : s = 240;
	{8'd93,8'd148} : s = 241;
	{8'd93,8'd149} : s = 242;
	{8'd93,8'd150} : s = 243;
	{8'd93,8'd151} : s = 244;
	{8'd93,8'd152} : s = 245;
	{8'd93,8'd153} : s = 246;
	{8'd93,8'd154} : s = 247;
	{8'd93,8'd155} : s = 248;
	{8'd93,8'd156} : s = 249;
	{8'd93,8'd157} : s = 250;
	{8'd93,8'd158} : s = 251;
	{8'd93,8'd159} : s = 252;
	{8'd93,8'd160} : s = 253;
	{8'd93,8'd161} : s = 254;
	{8'd93,8'd162} : s = 255;
	{8'd93,8'd163} : s = 256;
	{8'd93,8'd164} : s = 257;
	{8'd93,8'd165} : s = 258;
	{8'd93,8'd166} : s = 259;
	{8'd93,8'd167} : s = 260;
	{8'd93,8'd168} : s = 261;
	{8'd93,8'd169} : s = 262;
	{8'd93,8'd170} : s = 263;
	{8'd93,8'd171} : s = 264;
	{8'd93,8'd172} : s = 265;
	{8'd93,8'd173} : s = 266;
	{8'd93,8'd174} : s = 267;
	{8'd93,8'd175} : s = 268;
	{8'd93,8'd176} : s = 269;
	{8'd93,8'd177} : s = 270;
	{8'd93,8'd178} : s = 271;
	{8'd93,8'd179} : s = 272;
	{8'd93,8'd180} : s = 273;
	{8'd93,8'd181} : s = 274;
	{8'd93,8'd182} : s = 275;
	{8'd93,8'd183} : s = 276;
	{8'd93,8'd184} : s = 277;
	{8'd93,8'd185} : s = 278;
	{8'd93,8'd186} : s = 279;
	{8'd93,8'd187} : s = 280;
	{8'd93,8'd188} : s = 281;
	{8'd93,8'd189} : s = 282;
	{8'd93,8'd190} : s = 283;
	{8'd93,8'd191} : s = 284;
	{8'd93,8'd192} : s = 285;
	{8'd93,8'd193} : s = 286;
	{8'd93,8'd194} : s = 287;
	{8'd93,8'd195} : s = 288;
	{8'd93,8'd196} : s = 289;
	{8'd93,8'd197} : s = 290;
	{8'd93,8'd198} : s = 291;
	{8'd93,8'd199} : s = 292;
	{8'd93,8'd200} : s = 293;
	{8'd93,8'd201} : s = 294;
	{8'd93,8'd202} : s = 295;
	{8'd93,8'd203} : s = 296;
	{8'd93,8'd204} : s = 297;
	{8'd93,8'd205} : s = 298;
	{8'd93,8'd206} : s = 299;
	{8'd93,8'd207} : s = 300;
	{8'd93,8'd208} : s = 301;
	{8'd93,8'd209} : s = 302;
	{8'd93,8'd210} : s = 303;
	{8'd93,8'd211} : s = 304;
	{8'd93,8'd212} : s = 305;
	{8'd93,8'd213} : s = 306;
	{8'd93,8'd214} : s = 307;
	{8'd93,8'd215} : s = 308;
	{8'd93,8'd216} : s = 309;
	{8'd93,8'd217} : s = 310;
	{8'd93,8'd218} : s = 311;
	{8'd93,8'd219} : s = 312;
	{8'd93,8'd220} : s = 313;
	{8'd93,8'd221} : s = 314;
	{8'd93,8'd222} : s = 315;
	{8'd93,8'd223} : s = 316;
	{8'd93,8'd224} : s = 317;
	{8'd93,8'd225} : s = 318;
	{8'd93,8'd226} : s = 319;
	{8'd93,8'd227} : s = 320;
	{8'd93,8'd228} : s = 321;
	{8'd93,8'd229} : s = 322;
	{8'd93,8'd230} : s = 323;
	{8'd93,8'd231} : s = 324;
	{8'd93,8'd232} : s = 325;
	{8'd93,8'd233} : s = 326;
	{8'd93,8'd234} : s = 327;
	{8'd93,8'd235} : s = 328;
	{8'd93,8'd236} : s = 329;
	{8'd93,8'd237} : s = 330;
	{8'd93,8'd238} : s = 331;
	{8'd93,8'd239} : s = 332;
	{8'd93,8'd240} : s = 333;
	{8'd93,8'd241} : s = 334;
	{8'd93,8'd242} : s = 335;
	{8'd93,8'd243} : s = 336;
	{8'd93,8'd244} : s = 337;
	{8'd93,8'd245} : s = 338;
	{8'd93,8'd246} : s = 339;
	{8'd93,8'd247} : s = 340;
	{8'd93,8'd248} : s = 341;
	{8'd93,8'd249} : s = 342;
	{8'd93,8'd250} : s = 343;
	{8'd93,8'd251} : s = 344;
	{8'd93,8'd252} : s = 345;
	{8'd93,8'd253} : s = 346;
	{8'd93,8'd254} : s = 347;
	{8'd93,8'd255} : s = 348;
	{8'd94,8'd0} : s = 94;
	{8'd94,8'd1} : s = 95;
	{8'd94,8'd2} : s = 96;
	{8'd94,8'd3} : s = 97;
	{8'd94,8'd4} : s = 98;
	{8'd94,8'd5} : s = 99;
	{8'd94,8'd6} : s = 100;
	{8'd94,8'd7} : s = 101;
	{8'd94,8'd8} : s = 102;
	{8'd94,8'd9} : s = 103;
	{8'd94,8'd10} : s = 104;
	{8'd94,8'd11} : s = 105;
	{8'd94,8'd12} : s = 106;
	{8'd94,8'd13} : s = 107;
	{8'd94,8'd14} : s = 108;
	{8'd94,8'd15} : s = 109;
	{8'd94,8'd16} : s = 110;
	{8'd94,8'd17} : s = 111;
	{8'd94,8'd18} : s = 112;
	{8'd94,8'd19} : s = 113;
	{8'd94,8'd20} : s = 114;
	{8'd94,8'd21} : s = 115;
	{8'd94,8'd22} : s = 116;
	{8'd94,8'd23} : s = 117;
	{8'd94,8'd24} : s = 118;
	{8'd94,8'd25} : s = 119;
	{8'd94,8'd26} : s = 120;
	{8'd94,8'd27} : s = 121;
	{8'd94,8'd28} : s = 122;
	{8'd94,8'd29} : s = 123;
	{8'd94,8'd30} : s = 124;
	{8'd94,8'd31} : s = 125;
	{8'd94,8'd32} : s = 126;
	{8'd94,8'd33} : s = 127;
	{8'd94,8'd34} : s = 128;
	{8'd94,8'd35} : s = 129;
	{8'd94,8'd36} : s = 130;
	{8'd94,8'd37} : s = 131;
	{8'd94,8'd38} : s = 132;
	{8'd94,8'd39} : s = 133;
	{8'd94,8'd40} : s = 134;
	{8'd94,8'd41} : s = 135;
	{8'd94,8'd42} : s = 136;
	{8'd94,8'd43} : s = 137;
	{8'd94,8'd44} : s = 138;
	{8'd94,8'd45} : s = 139;
	{8'd94,8'd46} : s = 140;
	{8'd94,8'd47} : s = 141;
	{8'd94,8'd48} : s = 142;
	{8'd94,8'd49} : s = 143;
	{8'd94,8'd50} : s = 144;
	{8'd94,8'd51} : s = 145;
	{8'd94,8'd52} : s = 146;
	{8'd94,8'd53} : s = 147;
	{8'd94,8'd54} : s = 148;
	{8'd94,8'd55} : s = 149;
	{8'd94,8'd56} : s = 150;
	{8'd94,8'd57} : s = 151;
	{8'd94,8'd58} : s = 152;
	{8'd94,8'd59} : s = 153;
	{8'd94,8'd60} : s = 154;
	{8'd94,8'd61} : s = 155;
	{8'd94,8'd62} : s = 156;
	{8'd94,8'd63} : s = 157;
	{8'd94,8'd64} : s = 158;
	{8'd94,8'd65} : s = 159;
	{8'd94,8'd66} : s = 160;
	{8'd94,8'd67} : s = 161;
	{8'd94,8'd68} : s = 162;
	{8'd94,8'd69} : s = 163;
	{8'd94,8'd70} : s = 164;
	{8'd94,8'd71} : s = 165;
	{8'd94,8'd72} : s = 166;
	{8'd94,8'd73} : s = 167;
	{8'd94,8'd74} : s = 168;
	{8'd94,8'd75} : s = 169;
	{8'd94,8'd76} : s = 170;
	{8'd94,8'd77} : s = 171;
	{8'd94,8'd78} : s = 172;
	{8'd94,8'd79} : s = 173;
	{8'd94,8'd80} : s = 174;
	{8'd94,8'd81} : s = 175;
	{8'd94,8'd82} : s = 176;
	{8'd94,8'd83} : s = 177;
	{8'd94,8'd84} : s = 178;
	{8'd94,8'd85} : s = 179;
	{8'd94,8'd86} : s = 180;
	{8'd94,8'd87} : s = 181;
	{8'd94,8'd88} : s = 182;
	{8'd94,8'd89} : s = 183;
	{8'd94,8'd90} : s = 184;
	{8'd94,8'd91} : s = 185;
	{8'd94,8'd92} : s = 186;
	{8'd94,8'd93} : s = 187;
	{8'd94,8'd94} : s = 188;
	{8'd94,8'd95} : s = 189;
	{8'd94,8'd96} : s = 190;
	{8'd94,8'd97} : s = 191;
	{8'd94,8'd98} : s = 192;
	{8'd94,8'd99} : s = 193;
	{8'd94,8'd100} : s = 194;
	{8'd94,8'd101} : s = 195;
	{8'd94,8'd102} : s = 196;
	{8'd94,8'd103} : s = 197;
	{8'd94,8'd104} : s = 198;
	{8'd94,8'd105} : s = 199;
	{8'd94,8'd106} : s = 200;
	{8'd94,8'd107} : s = 201;
	{8'd94,8'd108} : s = 202;
	{8'd94,8'd109} : s = 203;
	{8'd94,8'd110} : s = 204;
	{8'd94,8'd111} : s = 205;
	{8'd94,8'd112} : s = 206;
	{8'd94,8'd113} : s = 207;
	{8'd94,8'd114} : s = 208;
	{8'd94,8'd115} : s = 209;
	{8'd94,8'd116} : s = 210;
	{8'd94,8'd117} : s = 211;
	{8'd94,8'd118} : s = 212;
	{8'd94,8'd119} : s = 213;
	{8'd94,8'd120} : s = 214;
	{8'd94,8'd121} : s = 215;
	{8'd94,8'd122} : s = 216;
	{8'd94,8'd123} : s = 217;
	{8'd94,8'd124} : s = 218;
	{8'd94,8'd125} : s = 219;
	{8'd94,8'd126} : s = 220;
	{8'd94,8'd127} : s = 221;
	{8'd94,8'd128} : s = 222;
	{8'd94,8'd129} : s = 223;
	{8'd94,8'd130} : s = 224;
	{8'd94,8'd131} : s = 225;
	{8'd94,8'd132} : s = 226;
	{8'd94,8'd133} : s = 227;
	{8'd94,8'd134} : s = 228;
	{8'd94,8'd135} : s = 229;
	{8'd94,8'd136} : s = 230;
	{8'd94,8'd137} : s = 231;
	{8'd94,8'd138} : s = 232;
	{8'd94,8'd139} : s = 233;
	{8'd94,8'd140} : s = 234;
	{8'd94,8'd141} : s = 235;
	{8'd94,8'd142} : s = 236;
	{8'd94,8'd143} : s = 237;
	{8'd94,8'd144} : s = 238;
	{8'd94,8'd145} : s = 239;
	{8'd94,8'd146} : s = 240;
	{8'd94,8'd147} : s = 241;
	{8'd94,8'd148} : s = 242;
	{8'd94,8'd149} : s = 243;
	{8'd94,8'd150} : s = 244;
	{8'd94,8'd151} : s = 245;
	{8'd94,8'd152} : s = 246;
	{8'd94,8'd153} : s = 247;
	{8'd94,8'd154} : s = 248;
	{8'd94,8'd155} : s = 249;
	{8'd94,8'd156} : s = 250;
	{8'd94,8'd157} : s = 251;
	{8'd94,8'd158} : s = 252;
	{8'd94,8'd159} : s = 253;
	{8'd94,8'd160} : s = 254;
	{8'd94,8'd161} : s = 255;
	{8'd94,8'd162} : s = 256;
	{8'd94,8'd163} : s = 257;
	{8'd94,8'd164} : s = 258;
	{8'd94,8'd165} : s = 259;
	{8'd94,8'd166} : s = 260;
	{8'd94,8'd167} : s = 261;
	{8'd94,8'd168} : s = 262;
	{8'd94,8'd169} : s = 263;
	{8'd94,8'd170} : s = 264;
	{8'd94,8'd171} : s = 265;
	{8'd94,8'd172} : s = 266;
	{8'd94,8'd173} : s = 267;
	{8'd94,8'd174} : s = 268;
	{8'd94,8'd175} : s = 269;
	{8'd94,8'd176} : s = 270;
	{8'd94,8'd177} : s = 271;
	{8'd94,8'd178} : s = 272;
	{8'd94,8'd179} : s = 273;
	{8'd94,8'd180} : s = 274;
	{8'd94,8'd181} : s = 275;
	{8'd94,8'd182} : s = 276;
	{8'd94,8'd183} : s = 277;
	{8'd94,8'd184} : s = 278;
	{8'd94,8'd185} : s = 279;
	{8'd94,8'd186} : s = 280;
	{8'd94,8'd187} : s = 281;
	{8'd94,8'd188} : s = 282;
	{8'd94,8'd189} : s = 283;
	{8'd94,8'd190} : s = 284;
	{8'd94,8'd191} : s = 285;
	{8'd94,8'd192} : s = 286;
	{8'd94,8'd193} : s = 287;
	{8'd94,8'd194} : s = 288;
	{8'd94,8'd195} : s = 289;
	{8'd94,8'd196} : s = 290;
	{8'd94,8'd197} : s = 291;
	{8'd94,8'd198} : s = 292;
	{8'd94,8'd199} : s = 293;
	{8'd94,8'd200} : s = 294;
	{8'd94,8'd201} : s = 295;
	{8'd94,8'd202} : s = 296;
	{8'd94,8'd203} : s = 297;
	{8'd94,8'd204} : s = 298;
	{8'd94,8'd205} : s = 299;
	{8'd94,8'd206} : s = 300;
	{8'd94,8'd207} : s = 301;
	{8'd94,8'd208} : s = 302;
	{8'd94,8'd209} : s = 303;
	{8'd94,8'd210} : s = 304;
	{8'd94,8'd211} : s = 305;
	{8'd94,8'd212} : s = 306;
	{8'd94,8'd213} : s = 307;
	{8'd94,8'd214} : s = 308;
	{8'd94,8'd215} : s = 309;
	{8'd94,8'd216} : s = 310;
	{8'd94,8'd217} : s = 311;
	{8'd94,8'd218} : s = 312;
	{8'd94,8'd219} : s = 313;
	{8'd94,8'd220} : s = 314;
	{8'd94,8'd221} : s = 315;
	{8'd94,8'd222} : s = 316;
	{8'd94,8'd223} : s = 317;
	{8'd94,8'd224} : s = 318;
	{8'd94,8'd225} : s = 319;
	{8'd94,8'd226} : s = 320;
	{8'd94,8'd227} : s = 321;
	{8'd94,8'd228} : s = 322;
	{8'd94,8'd229} : s = 323;
	{8'd94,8'd230} : s = 324;
	{8'd94,8'd231} : s = 325;
	{8'd94,8'd232} : s = 326;
	{8'd94,8'd233} : s = 327;
	{8'd94,8'd234} : s = 328;
	{8'd94,8'd235} : s = 329;
	{8'd94,8'd236} : s = 330;
	{8'd94,8'd237} : s = 331;
	{8'd94,8'd238} : s = 332;
	{8'd94,8'd239} : s = 333;
	{8'd94,8'd240} : s = 334;
	{8'd94,8'd241} : s = 335;
	{8'd94,8'd242} : s = 336;
	{8'd94,8'd243} : s = 337;
	{8'd94,8'd244} : s = 338;
	{8'd94,8'd245} : s = 339;
	{8'd94,8'd246} : s = 340;
	{8'd94,8'd247} : s = 341;
	{8'd94,8'd248} : s = 342;
	{8'd94,8'd249} : s = 343;
	{8'd94,8'd250} : s = 344;
	{8'd94,8'd251} : s = 345;
	{8'd94,8'd252} : s = 346;
	{8'd94,8'd253} : s = 347;
	{8'd94,8'd254} : s = 348;
	{8'd94,8'd255} : s = 349;
	{8'd95,8'd0} : s = 95;
	{8'd95,8'd1} : s = 96;
	{8'd95,8'd2} : s = 97;
	{8'd95,8'd3} : s = 98;
	{8'd95,8'd4} : s = 99;
	{8'd95,8'd5} : s = 100;
	{8'd95,8'd6} : s = 101;
	{8'd95,8'd7} : s = 102;
	{8'd95,8'd8} : s = 103;
	{8'd95,8'd9} : s = 104;
	{8'd95,8'd10} : s = 105;
	{8'd95,8'd11} : s = 106;
	{8'd95,8'd12} : s = 107;
	{8'd95,8'd13} : s = 108;
	{8'd95,8'd14} : s = 109;
	{8'd95,8'd15} : s = 110;
	{8'd95,8'd16} : s = 111;
	{8'd95,8'd17} : s = 112;
	{8'd95,8'd18} : s = 113;
	{8'd95,8'd19} : s = 114;
	{8'd95,8'd20} : s = 115;
	{8'd95,8'd21} : s = 116;
	{8'd95,8'd22} : s = 117;
	{8'd95,8'd23} : s = 118;
	{8'd95,8'd24} : s = 119;
	{8'd95,8'd25} : s = 120;
	{8'd95,8'd26} : s = 121;
	{8'd95,8'd27} : s = 122;
	{8'd95,8'd28} : s = 123;
	{8'd95,8'd29} : s = 124;
	{8'd95,8'd30} : s = 125;
	{8'd95,8'd31} : s = 126;
	{8'd95,8'd32} : s = 127;
	{8'd95,8'd33} : s = 128;
	{8'd95,8'd34} : s = 129;
	{8'd95,8'd35} : s = 130;
	{8'd95,8'd36} : s = 131;
	{8'd95,8'd37} : s = 132;
	{8'd95,8'd38} : s = 133;
	{8'd95,8'd39} : s = 134;
	{8'd95,8'd40} : s = 135;
	{8'd95,8'd41} : s = 136;
	{8'd95,8'd42} : s = 137;
	{8'd95,8'd43} : s = 138;
	{8'd95,8'd44} : s = 139;
	{8'd95,8'd45} : s = 140;
	{8'd95,8'd46} : s = 141;
	{8'd95,8'd47} : s = 142;
	{8'd95,8'd48} : s = 143;
	{8'd95,8'd49} : s = 144;
	{8'd95,8'd50} : s = 145;
	{8'd95,8'd51} : s = 146;
	{8'd95,8'd52} : s = 147;
	{8'd95,8'd53} : s = 148;
	{8'd95,8'd54} : s = 149;
	{8'd95,8'd55} : s = 150;
	{8'd95,8'd56} : s = 151;
	{8'd95,8'd57} : s = 152;
	{8'd95,8'd58} : s = 153;
	{8'd95,8'd59} : s = 154;
	{8'd95,8'd60} : s = 155;
	{8'd95,8'd61} : s = 156;
	{8'd95,8'd62} : s = 157;
	{8'd95,8'd63} : s = 158;
	{8'd95,8'd64} : s = 159;
	{8'd95,8'd65} : s = 160;
	{8'd95,8'd66} : s = 161;
	{8'd95,8'd67} : s = 162;
	{8'd95,8'd68} : s = 163;
	{8'd95,8'd69} : s = 164;
	{8'd95,8'd70} : s = 165;
	{8'd95,8'd71} : s = 166;
	{8'd95,8'd72} : s = 167;
	{8'd95,8'd73} : s = 168;
	{8'd95,8'd74} : s = 169;
	{8'd95,8'd75} : s = 170;
	{8'd95,8'd76} : s = 171;
	{8'd95,8'd77} : s = 172;
	{8'd95,8'd78} : s = 173;
	{8'd95,8'd79} : s = 174;
	{8'd95,8'd80} : s = 175;
	{8'd95,8'd81} : s = 176;
	{8'd95,8'd82} : s = 177;
	{8'd95,8'd83} : s = 178;
	{8'd95,8'd84} : s = 179;
	{8'd95,8'd85} : s = 180;
	{8'd95,8'd86} : s = 181;
	{8'd95,8'd87} : s = 182;
	{8'd95,8'd88} : s = 183;
	{8'd95,8'd89} : s = 184;
	{8'd95,8'd90} : s = 185;
	{8'd95,8'd91} : s = 186;
	{8'd95,8'd92} : s = 187;
	{8'd95,8'd93} : s = 188;
	{8'd95,8'd94} : s = 189;
	{8'd95,8'd95} : s = 190;
	{8'd95,8'd96} : s = 191;
	{8'd95,8'd97} : s = 192;
	{8'd95,8'd98} : s = 193;
	{8'd95,8'd99} : s = 194;
	{8'd95,8'd100} : s = 195;
	{8'd95,8'd101} : s = 196;
	{8'd95,8'd102} : s = 197;
	{8'd95,8'd103} : s = 198;
	{8'd95,8'd104} : s = 199;
	{8'd95,8'd105} : s = 200;
	{8'd95,8'd106} : s = 201;
	{8'd95,8'd107} : s = 202;
	{8'd95,8'd108} : s = 203;
	{8'd95,8'd109} : s = 204;
	{8'd95,8'd110} : s = 205;
	{8'd95,8'd111} : s = 206;
	{8'd95,8'd112} : s = 207;
	{8'd95,8'd113} : s = 208;
	{8'd95,8'd114} : s = 209;
	{8'd95,8'd115} : s = 210;
	{8'd95,8'd116} : s = 211;
	{8'd95,8'd117} : s = 212;
	{8'd95,8'd118} : s = 213;
	{8'd95,8'd119} : s = 214;
	{8'd95,8'd120} : s = 215;
	{8'd95,8'd121} : s = 216;
	{8'd95,8'd122} : s = 217;
	{8'd95,8'd123} : s = 218;
	{8'd95,8'd124} : s = 219;
	{8'd95,8'd125} : s = 220;
	{8'd95,8'd126} : s = 221;
	{8'd95,8'd127} : s = 222;
	{8'd95,8'd128} : s = 223;
	{8'd95,8'd129} : s = 224;
	{8'd95,8'd130} : s = 225;
	{8'd95,8'd131} : s = 226;
	{8'd95,8'd132} : s = 227;
	{8'd95,8'd133} : s = 228;
	{8'd95,8'd134} : s = 229;
	{8'd95,8'd135} : s = 230;
	{8'd95,8'd136} : s = 231;
	{8'd95,8'd137} : s = 232;
	{8'd95,8'd138} : s = 233;
	{8'd95,8'd139} : s = 234;
	{8'd95,8'd140} : s = 235;
	{8'd95,8'd141} : s = 236;
	{8'd95,8'd142} : s = 237;
	{8'd95,8'd143} : s = 238;
	{8'd95,8'd144} : s = 239;
	{8'd95,8'd145} : s = 240;
	{8'd95,8'd146} : s = 241;
	{8'd95,8'd147} : s = 242;
	{8'd95,8'd148} : s = 243;
	{8'd95,8'd149} : s = 244;
	{8'd95,8'd150} : s = 245;
	{8'd95,8'd151} : s = 246;
	{8'd95,8'd152} : s = 247;
	{8'd95,8'd153} : s = 248;
	{8'd95,8'd154} : s = 249;
	{8'd95,8'd155} : s = 250;
	{8'd95,8'd156} : s = 251;
	{8'd95,8'd157} : s = 252;
	{8'd95,8'd158} : s = 253;
	{8'd95,8'd159} : s = 254;
	{8'd95,8'd160} : s = 255;
	{8'd95,8'd161} : s = 256;
	{8'd95,8'd162} : s = 257;
	{8'd95,8'd163} : s = 258;
	{8'd95,8'd164} : s = 259;
	{8'd95,8'd165} : s = 260;
	{8'd95,8'd166} : s = 261;
	{8'd95,8'd167} : s = 262;
	{8'd95,8'd168} : s = 263;
	{8'd95,8'd169} : s = 264;
	{8'd95,8'd170} : s = 265;
	{8'd95,8'd171} : s = 266;
	{8'd95,8'd172} : s = 267;
	{8'd95,8'd173} : s = 268;
	{8'd95,8'd174} : s = 269;
	{8'd95,8'd175} : s = 270;
	{8'd95,8'd176} : s = 271;
	{8'd95,8'd177} : s = 272;
	{8'd95,8'd178} : s = 273;
	{8'd95,8'd179} : s = 274;
	{8'd95,8'd180} : s = 275;
	{8'd95,8'd181} : s = 276;
	{8'd95,8'd182} : s = 277;
	{8'd95,8'd183} : s = 278;
	{8'd95,8'd184} : s = 279;
	{8'd95,8'd185} : s = 280;
	{8'd95,8'd186} : s = 281;
	{8'd95,8'd187} : s = 282;
	{8'd95,8'd188} : s = 283;
	{8'd95,8'd189} : s = 284;
	{8'd95,8'd190} : s = 285;
	{8'd95,8'd191} : s = 286;
	{8'd95,8'd192} : s = 287;
	{8'd95,8'd193} : s = 288;
	{8'd95,8'd194} : s = 289;
	{8'd95,8'd195} : s = 290;
	{8'd95,8'd196} : s = 291;
	{8'd95,8'd197} : s = 292;
	{8'd95,8'd198} : s = 293;
	{8'd95,8'd199} : s = 294;
	{8'd95,8'd200} : s = 295;
	{8'd95,8'd201} : s = 296;
	{8'd95,8'd202} : s = 297;
	{8'd95,8'd203} : s = 298;
	{8'd95,8'd204} : s = 299;
	{8'd95,8'd205} : s = 300;
	{8'd95,8'd206} : s = 301;
	{8'd95,8'd207} : s = 302;
	{8'd95,8'd208} : s = 303;
	{8'd95,8'd209} : s = 304;
	{8'd95,8'd210} : s = 305;
	{8'd95,8'd211} : s = 306;
	{8'd95,8'd212} : s = 307;
	{8'd95,8'd213} : s = 308;
	{8'd95,8'd214} : s = 309;
	{8'd95,8'd215} : s = 310;
	{8'd95,8'd216} : s = 311;
	{8'd95,8'd217} : s = 312;
	{8'd95,8'd218} : s = 313;
	{8'd95,8'd219} : s = 314;
	{8'd95,8'd220} : s = 315;
	{8'd95,8'd221} : s = 316;
	{8'd95,8'd222} : s = 317;
	{8'd95,8'd223} : s = 318;
	{8'd95,8'd224} : s = 319;
	{8'd95,8'd225} : s = 320;
	{8'd95,8'd226} : s = 321;
	{8'd95,8'd227} : s = 322;
	{8'd95,8'd228} : s = 323;
	{8'd95,8'd229} : s = 324;
	{8'd95,8'd230} : s = 325;
	{8'd95,8'd231} : s = 326;
	{8'd95,8'd232} : s = 327;
	{8'd95,8'd233} : s = 328;
	{8'd95,8'd234} : s = 329;
	{8'd95,8'd235} : s = 330;
	{8'd95,8'd236} : s = 331;
	{8'd95,8'd237} : s = 332;
	{8'd95,8'd238} : s = 333;
	{8'd95,8'd239} : s = 334;
	{8'd95,8'd240} : s = 335;
	{8'd95,8'd241} : s = 336;
	{8'd95,8'd242} : s = 337;
	{8'd95,8'd243} : s = 338;
	{8'd95,8'd244} : s = 339;
	{8'd95,8'd245} : s = 340;
	{8'd95,8'd246} : s = 341;
	{8'd95,8'd247} : s = 342;
	{8'd95,8'd248} : s = 343;
	{8'd95,8'd249} : s = 344;
	{8'd95,8'd250} : s = 345;
	{8'd95,8'd251} : s = 346;
	{8'd95,8'd252} : s = 347;
	{8'd95,8'd253} : s = 348;
	{8'd95,8'd254} : s = 349;
	{8'd95,8'd255} : s = 350;
	{8'd96,8'd0} : s = 96;
	{8'd96,8'd1} : s = 97;
	{8'd96,8'd2} : s = 98;
	{8'd96,8'd3} : s = 99;
	{8'd96,8'd4} : s = 100;
	{8'd96,8'd5} : s = 101;
	{8'd96,8'd6} : s = 102;
	{8'd96,8'd7} : s = 103;
	{8'd96,8'd8} : s = 104;
	{8'd96,8'd9} : s = 105;
	{8'd96,8'd10} : s = 106;
	{8'd96,8'd11} : s = 107;
	{8'd96,8'd12} : s = 108;
	{8'd96,8'd13} : s = 109;
	{8'd96,8'd14} : s = 110;
	{8'd96,8'd15} : s = 111;
	{8'd96,8'd16} : s = 112;
	{8'd96,8'd17} : s = 113;
	{8'd96,8'd18} : s = 114;
	{8'd96,8'd19} : s = 115;
	{8'd96,8'd20} : s = 116;
	{8'd96,8'd21} : s = 117;
	{8'd96,8'd22} : s = 118;
	{8'd96,8'd23} : s = 119;
	{8'd96,8'd24} : s = 120;
	{8'd96,8'd25} : s = 121;
	{8'd96,8'd26} : s = 122;
	{8'd96,8'd27} : s = 123;
	{8'd96,8'd28} : s = 124;
	{8'd96,8'd29} : s = 125;
	{8'd96,8'd30} : s = 126;
	{8'd96,8'd31} : s = 127;
	{8'd96,8'd32} : s = 128;
	{8'd96,8'd33} : s = 129;
	{8'd96,8'd34} : s = 130;
	{8'd96,8'd35} : s = 131;
	{8'd96,8'd36} : s = 132;
	{8'd96,8'd37} : s = 133;
	{8'd96,8'd38} : s = 134;
	{8'd96,8'd39} : s = 135;
	{8'd96,8'd40} : s = 136;
	{8'd96,8'd41} : s = 137;
	{8'd96,8'd42} : s = 138;
	{8'd96,8'd43} : s = 139;
	{8'd96,8'd44} : s = 140;
	{8'd96,8'd45} : s = 141;
	{8'd96,8'd46} : s = 142;
	{8'd96,8'd47} : s = 143;
	{8'd96,8'd48} : s = 144;
	{8'd96,8'd49} : s = 145;
	{8'd96,8'd50} : s = 146;
	{8'd96,8'd51} : s = 147;
	{8'd96,8'd52} : s = 148;
	{8'd96,8'd53} : s = 149;
	{8'd96,8'd54} : s = 150;
	{8'd96,8'd55} : s = 151;
	{8'd96,8'd56} : s = 152;
	{8'd96,8'd57} : s = 153;
	{8'd96,8'd58} : s = 154;
	{8'd96,8'd59} : s = 155;
	{8'd96,8'd60} : s = 156;
	{8'd96,8'd61} : s = 157;
	{8'd96,8'd62} : s = 158;
	{8'd96,8'd63} : s = 159;
	{8'd96,8'd64} : s = 160;
	{8'd96,8'd65} : s = 161;
	{8'd96,8'd66} : s = 162;
	{8'd96,8'd67} : s = 163;
	{8'd96,8'd68} : s = 164;
	{8'd96,8'd69} : s = 165;
	{8'd96,8'd70} : s = 166;
	{8'd96,8'd71} : s = 167;
	{8'd96,8'd72} : s = 168;
	{8'd96,8'd73} : s = 169;
	{8'd96,8'd74} : s = 170;
	{8'd96,8'd75} : s = 171;
	{8'd96,8'd76} : s = 172;
	{8'd96,8'd77} : s = 173;
	{8'd96,8'd78} : s = 174;
	{8'd96,8'd79} : s = 175;
	{8'd96,8'd80} : s = 176;
	{8'd96,8'd81} : s = 177;
	{8'd96,8'd82} : s = 178;
	{8'd96,8'd83} : s = 179;
	{8'd96,8'd84} : s = 180;
	{8'd96,8'd85} : s = 181;
	{8'd96,8'd86} : s = 182;
	{8'd96,8'd87} : s = 183;
	{8'd96,8'd88} : s = 184;
	{8'd96,8'd89} : s = 185;
	{8'd96,8'd90} : s = 186;
	{8'd96,8'd91} : s = 187;
	{8'd96,8'd92} : s = 188;
	{8'd96,8'd93} : s = 189;
	{8'd96,8'd94} : s = 190;
	{8'd96,8'd95} : s = 191;
	{8'd96,8'd96} : s = 192;
	{8'd96,8'd97} : s = 193;
	{8'd96,8'd98} : s = 194;
	{8'd96,8'd99} : s = 195;
	{8'd96,8'd100} : s = 196;
	{8'd96,8'd101} : s = 197;
	{8'd96,8'd102} : s = 198;
	{8'd96,8'd103} : s = 199;
	{8'd96,8'd104} : s = 200;
	{8'd96,8'd105} : s = 201;
	{8'd96,8'd106} : s = 202;
	{8'd96,8'd107} : s = 203;
	{8'd96,8'd108} : s = 204;
	{8'd96,8'd109} : s = 205;
	{8'd96,8'd110} : s = 206;
	{8'd96,8'd111} : s = 207;
	{8'd96,8'd112} : s = 208;
	{8'd96,8'd113} : s = 209;
	{8'd96,8'd114} : s = 210;
	{8'd96,8'd115} : s = 211;
	{8'd96,8'd116} : s = 212;
	{8'd96,8'd117} : s = 213;
	{8'd96,8'd118} : s = 214;
	{8'd96,8'd119} : s = 215;
	{8'd96,8'd120} : s = 216;
	{8'd96,8'd121} : s = 217;
	{8'd96,8'd122} : s = 218;
	{8'd96,8'd123} : s = 219;
	{8'd96,8'd124} : s = 220;
	{8'd96,8'd125} : s = 221;
	{8'd96,8'd126} : s = 222;
	{8'd96,8'd127} : s = 223;
	{8'd96,8'd128} : s = 224;
	{8'd96,8'd129} : s = 225;
	{8'd96,8'd130} : s = 226;
	{8'd96,8'd131} : s = 227;
	{8'd96,8'd132} : s = 228;
	{8'd96,8'd133} : s = 229;
	{8'd96,8'd134} : s = 230;
	{8'd96,8'd135} : s = 231;
	{8'd96,8'd136} : s = 232;
	{8'd96,8'd137} : s = 233;
	{8'd96,8'd138} : s = 234;
	{8'd96,8'd139} : s = 235;
	{8'd96,8'd140} : s = 236;
	{8'd96,8'd141} : s = 237;
	{8'd96,8'd142} : s = 238;
	{8'd96,8'd143} : s = 239;
	{8'd96,8'd144} : s = 240;
	{8'd96,8'd145} : s = 241;
	{8'd96,8'd146} : s = 242;
	{8'd96,8'd147} : s = 243;
	{8'd96,8'd148} : s = 244;
	{8'd96,8'd149} : s = 245;
	{8'd96,8'd150} : s = 246;
	{8'd96,8'd151} : s = 247;
	{8'd96,8'd152} : s = 248;
	{8'd96,8'd153} : s = 249;
	{8'd96,8'd154} : s = 250;
	{8'd96,8'd155} : s = 251;
	{8'd96,8'd156} : s = 252;
	{8'd96,8'd157} : s = 253;
	{8'd96,8'd158} : s = 254;
	{8'd96,8'd159} : s = 255;
	{8'd96,8'd160} : s = 256;
	{8'd96,8'd161} : s = 257;
	{8'd96,8'd162} : s = 258;
	{8'd96,8'd163} : s = 259;
	{8'd96,8'd164} : s = 260;
	{8'd96,8'd165} : s = 261;
	{8'd96,8'd166} : s = 262;
	{8'd96,8'd167} : s = 263;
	{8'd96,8'd168} : s = 264;
	{8'd96,8'd169} : s = 265;
	{8'd96,8'd170} : s = 266;
	{8'd96,8'd171} : s = 267;
	{8'd96,8'd172} : s = 268;
	{8'd96,8'd173} : s = 269;
	{8'd96,8'd174} : s = 270;
	{8'd96,8'd175} : s = 271;
	{8'd96,8'd176} : s = 272;
	{8'd96,8'd177} : s = 273;
	{8'd96,8'd178} : s = 274;
	{8'd96,8'd179} : s = 275;
	{8'd96,8'd180} : s = 276;
	{8'd96,8'd181} : s = 277;
	{8'd96,8'd182} : s = 278;
	{8'd96,8'd183} : s = 279;
	{8'd96,8'd184} : s = 280;
	{8'd96,8'd185} : s = 281;
	{8'd96,8'd186} : s = 282;
	{8'd96,8'd187} : s = 283;
	{8'd96,8'd188} : s = 284;
	{8'd96,8'd189} : s = 285;
	{8'd96,8'd190} : s = 286;
	{8'd96,8'd191} : s = 287;
	{8'd96,8'd192} : s = 288;
	{8'd96,8'd193} : s = 289;
	{8'd96,8'd194} : s = 290;
	{8'd96,8'd195} : s = 291;
	{8'd96,8'd196} : s = 292;
	{8'd96,8'd197} : s = 293;
	{8'd96,8'd198} : s = 294;
	{8'd96,8'd199} : s = 295;
	{8'd96,8'd200} : s = 296;
	{8'd96,8'd201} : s = 297;
	{8'd96,8'd202} : s = 298;
	{8'd96,8'd203} : s = 299;
	{8'd96,8'd204} : s = 300;
	{8'd96,8'd205} : s = 301;
	{8'd96,8'd206} : s = 302;
	{8'd96,8'd207} : s = 303;
	{8'd96,8'd208} : s = 304;
	{8'd96,8'd209} : s = 305;
	{8'd96,8'd210} : s = 306;
	{8'd96,8'd211} : s = 307;
	{8'd96,8'd212} : s = 308;
	{8'd96,8'd213} : s = 309;
	{8'd96,8'd214} : s = 310;
	{8'd96,8'd215} : s = 311;
	{8'd96,8'd216} : s = 312;
	{8'd96,8'd217} : s = 313;
	{8'd96,8'd218} : s = 314;
	{8'd96,8'd219} : s = 315;
	{8'd96,8'd220} : s = 316;
	{8'd96,8'd221} : s = 317;
	{8'd96,8'd222} : s = 318;
	{8'd96,8'd223} : s = 319;
	{8'd96,8'd224} : s = 320;
	{8'd96,8'd225} : s = 321;
	{8'd96,8'd226} : s = 322;
	{8'd96,8'd227} : s = 323;
	{8'd96,8'd228} : s = 324;
	{8'd96,8'd229} : s = 325;
	{8'd96,8'd230} : s = 326;
	{8'd96,8'd231} : s = 327;
	{8'd96,8'd232} : s = 328;
	{8'd96,8'd233} : s = 329;
	{8'd96,8'd234} : s = 330;
	{8'd96,8'd235} : s = 331;
	{8'd96,8'd236} : s = 332;
	{8'd96,8'd237} : s = 333;
	{8'd96,8'd238} : s = 334;
	{8'd96,8'd239} : s = 335;
	{8'd96,8'd240} : s = 336;
	{8'd96,8'd241} : s = 337;
	{8'd96,8'd242} : s = 338;
	{8'd96,8'd243} : s = 339;
	{8'd96,8'd244} : s = 340;
	{8'd96,8'd245} : s = 341;
	{8'd96,8'd246} : s = 342;
	{8'd96,8'd247} : s = 343;
	{8'd96,8'd248} : s = 344;
	{8'd96,8'd249} : s = 345;
	{8'd96,8'd250} : s = 346;
	{8'd96,8'd251} : s = 347;
	{8'd96,8'd252} : s = 348;
	{8'd96,8'd253} : s = 349;
	{8'd96,8'd254} : s = 350;
	{8'd96,8'd255} : s = 351;
	{8'd97,8'd0} : s = 97;
	{8'd97,8'd1} : s = 98;
	{8'd97,8'd2} : s = 99;
	{8'd97,8'd3} : s = 100;
	{8'd97,8'd4} : s = 101;
	{8'd97,8'd5} : s = 102;
	{8'd97,8'd6} : s = 103;
	{8'd97,8'd7} : s = 104;
	{8'd97,8'd8} : s = 105;
	{8'd97,8'd9} : s = 106;
	{8'd97,8'd10} : s = 107;
	{8'd97,8'd11} : s = 108;
	{8'd97,8'd12} : s = 109;
	{8'd97,8'd13} : s = 110;
	{8'd97,8'd14} : s = 111;
	{8'd97,8'd15} : s = 112;
	{8'd97,8'd16} : s = 113;
	{8'd97,8'd17} : s = 114;
	{8'd97,8'd18} : s = 115;
	{8'd97,8'd19} : s = 116;
	{8'd97,8'd20} : s = 117;
	{8'd97,8'd21} : s = 118;
	{8'd97,8'd22} : s = 119;
	{8'd97,8'd23} : s = 120;
	{8'd97,8'd24} : s = 121;
	{8'd97,8'd25} : s = 122;
	{8'd97,8'd26} : s = 123;
	{8'd97,8'd27} : s = 124;
	{8'd97,8'd28} : s = 125;
	{8'd97,8'd29} : s = 126;
	{8'd97,8'd30} : s = 127;
	{8'd97,8'd31} : s = 128;
	{8'd97,8'd32} : s = 129;
	{8'd97,8'd33} : s = 130;
	{8'd97,8'd34} : s = 131;
	{8'd97,8'd35} : s = 132;
	{8'd97,8'd36} : s = 133;
	{8'd97,8'd37} : s = 134;
	{8'd97,8'd38} : s = 135;
	{8'd97,8'd39} : s = 136;
	{8'd97,8'd40} : s = 137;
	{8'd97,8'd41} : s = 138;
	{8'd97,8'd42} : s = 139;
	{8'd97,8'd43} : s = 140;
	{8'd97,8'd44} : s = 141;
	{8'd97,8'd45} : s = 142;
	{8'd97,8'd46} : s = 143;
	{8'd97,8'd47} : s = 144;
	{8'd97,8'd48} : s = 145;
	{8'd97,8'd49} : s = 146;
	{8'd97,8'd50} : s = 147;
	{8'd97,8'd51} : s = 148;
	{8'd97,8'd52} : s = 149;
	{8'd97,8'd53} : s = 150;
	{8'd97,8'd54} : s = 151;
	{8'd97,8'd55} : s = 152;
	{8'd97,8'd56} : s = 153;
	{8'd97,8'd57} : s = 154;
	{8'd97,8'd58} : s = 155;
	{8'd97,8'd59} : s = 156;
	{8'd97,8'd60} : s = 157;
	{8'd97,8'd61} : s = 158;
	{8'd97,8'd62} : s = 159;
	{8'd97,8'd63} : s = 160;
	{8'd97,8'd64} : s = 161;
	{8'd97,8'd65} : s = 162;
	{8'd97,8'd66} : s = 163;
	{8'd97,8'd67} : s = 164;
	{8'd97,8'd68} : s = 165;
	{8'd97,8'd69} : s = 166;
	{8'd97,8'd70} : s = 167;
	{8'd97,8'd71} : s = 168;
	{8'd97,8'd72} : s = 169;
	{8'd97,8'd73} : s = 170;
	{8'd97,8'd74} : s = 171;
	{8'd97,8'd75} : s = 172;
	{8'd97,8'd76} : s = 173;
	{8'd97,8'd77} : s = 174;
	{8'd97,8'd78} : s = 175;
	{8'd97,8'd79} : s = 176;
	{8'd97,8'd80} : s = 177;
	{8'd97,8'd81} : s = 178;
	{8'd97,8'd82} : s = 179;
	{8'd97,8'd83} : s = 180;
	{8'd97,8'd84} : s = 181;
	{8'd97,8'd85} : s = 182;
	{8'd97,8'd86} : s = 183;
	{8'd97,8'd87} : s = 184;
	{8'd97,8'd88} : s = 185;
	{8'd97,8'd89} : s = 186;
	{8'd97,8'd90} : s = 187;
	{8'd97,8'd91} : s = 188;
	{8'd97,8'd92} : s = 189;
	{8'd97,8'd93} : s = 190;
	{8'd97,8'd94} : s = 191;
	{8'd97,8'd95} : s = 192;
	{8'd97,8'd96} : s = 193;
	{8'd97,8'd97} : s = 194;
	{8'd97,8'd98} : s = 195;
	{8'd97,8'd99} : s = 196;
	{8'd97,8'd100} : s = 197;
	{8'd97,8'd101} : s = 198;
	{8'd97,8'd102} : s = 199;
	{8'd97,8'd103} : s = 200;
	{8'd97,8'd104} : s = 201;
	{8'd97,8'd105} : s = 202;
	{8'd97,8'd106} : s = 203;
	{8'd97,8'd107} : s = 204;
	{8'd97,8'd108} : s = 205;
	{8'd97,8'd109} : s = 206;
	{8'd97,8'd110} : s = 207;
	{8'd97,8'd111} : s = 208;
	{8'd97,8'd112} : s = 209;
	{8'd97,8'd113} : s = 210;
	{8'd97,8'd114} : s = 211;
	{8'd97,8'd115} : s = 212;
	{8'd97,8'd116} : s = 213;
	{8'd97,8'd117} : s = 214;
	{8'd97,8'd118} : s = 215;
	{8'd97,8'd119} : s = 216;
	{8'd97,8'd120} : s = 217;
	{8'd97,8'd121} : s = 218;
	{8'd97,8'd122} : s = 219;
	{8'd97,8'd123} : s = 220;
	{8'd97,8'd124} : s = 221;
	{8'd97,8'd125} : s = 222;
	{8'd97,8'd126} : s = 223;
	{8'd97,8'd127} : s = 224;
	{8'd97,8'd128} : s = 225;
	{8'd97,8'd129} : s = 226;
	{8'd97,8'd130} : s = 227;
	{8'd97,8'd131} : s = 228;
	{8'd97,8'd132} : s = 229;
	{8'd97,8'd133} : s = 230;
	{8'd97,8'd134} : s = 231;
	{8'd97,8'd135} : s = 232;
	{8'd97,8'd136} : s = 233;
	{8'd97,8'd137} : s = 234;
	{8'd97,8'd138} : s = 235;
	{8'd97,8'd139} : s = 236;
	{8'd97,8'd140} : s = 237;
	{8'd97,8'd141} : s = 238;
	{8'd97,8'd142} : s = 239;
	{8'd97,8'd143} : s = 240;
	{8'd97,8'd144} : s = 241;
	{8'd97,8'd145} : s = 242;
	{8'd97,8'd146} : s = 243;
	{8'd97,8'd147} : s = 244;
	{8'd97,8'd148} : s = 245;
	{8'd97,8'd149} : s = 246;
	{8'd97,8'd150} : s = 247;
	{8'd97,8'd151} : s = 248;
	{8'd97,8'd152} : s = 249;
	{8'd97,8'd153} : s = 250;
	{8'd97,8'd154} : s = 251;
	{8'd97,8'd155} : s = 252;
	{8'd97,8'd156} : s = 253;
	{8'd97,8'd157} : s = 254;
	{8'd97,8'd158} : s = 255;
	{8'd97,8'd159} : s = 256;
	{8'd97,8'd160} : s = 257;
	{8'd97,8'd161} : s = 258;
	{8'd97,8'd162} : s = 259;
	{8'd97,8'd163} : s = 260;
	{8'd97,8'd164} : s = 261;
	{8'd97,8'd165} : s = 262;
	{8'd97,8'd166} : s = 263;
	{8'd97,8'd167} : s = 264;
	{8'd97,8'd168} : s = 265;
	{8'd97,8'd169} : s = 266;
	{8'd97,8'd170} : s = 267;
	{8'd97,8'd171} : s = 268;
	{8'd97,8'd172} : s = 269;
	{8'd97,8'd173} : s = 270;
	{8'd97,8'd174} : s = 271;
	{8'd97,8'd175} : s = 272;
	{8'd97,8'd176} : s = 273;
	{8'd97,8'd177} : s = 274;
	{8'd97,8'd178} : s = 275;
	{8'd97,8'd179} : s = 276;
	{8'd97,8'd180} : s = 277;
	{8'd97,8'd181} : s = 278;
	{8'd97,8'd182} : s = 279;
	{8'd97,8'd183} : s = 280;
	{8'd97,8'd184} : s = 281;
	{8'd97,8'd185} : s = 282;
	{8'd97,8'd186} : s = 283;
	{8'd97,8'd187} : s = 284;
	{8'd97,8'd188} : s = 285;
	{8'd97,8'd189} : s = 286;
	{8'd97,8'd190} : s = 287;
	{8'd97,8'd191} : s = 288;
	{8'd97,8'd192} : s = 289;
	{8'd97,8'd193} : s = 290;
	{8'd97,8'd194} : s = 291;
	{8'd97,8'd195} : s = 292;
	{8'd97,8'd196} : s = 293;
	{8'd97,8'd197} : s = 294;
	{8'd97,8'd198} : s = 295;
	{8'd97,8'd199} : s = 296;
	{8'd97,8'd200} : s = 297;
	{8'd97,8'd201} : s = 298;
	{8'd97,8'd202} : s = 299;
	{8'd97,8'd203} : s = 300;
	{8'd97,8'd204} : s = 301;
	{8'd97,8'd205} : s = 302;
	{8'd97,8'd206} : s = 303;
	{8'd97,8'd207} : s = 304;
	{8'd97,8'd208} : s = 305;
	{8'd97,8'd209} : s = 306;
	{8'd97,8'd210} : s = 307;
	{8'd97,8'd211} : s = 308;
	{8'd97,8'd212} : s = 309;
	{8'd97,8'd213} : s = 310;
	{8'd97,8'd214} : s = 311;
	{8'd97,8'd215} : s = 312;
	{8'd97,8'd216} : s = 313;
	{8'd97,8'd217} : s = 314;
	{8'd97,8'd218} : s = 315;
	{8'd97,8'd219} : s = 316;
	{8'd97,8'd220} : s = 317;
	{8'd97,8'd221} : s = 318;
	{8'd97,8'd222} : s = 319;
	{8'd97,8'd223} : s = 320;
	{8'd97,8'd224} : s = 321;
	{8'd97,8'd225} : s = 322;
	{8'd97,8'd226} : s = 323;
	{8'd97,8'd227} : s = 324;
	{8'd97,8'd228} : s = 325;
	{8'd97,8'd229} : s = 326;
	{8'd97,8'd230} : s = 327;
	{8'd97,8'd231} : s = 328;
	{8'd97,8'd232} : s = 329;
	{8'd97,8'd233} : s = 330;
	{8'd97,8'd234} : s = 331;
	{8'd97,8'd235} : s = 332;
	{8'd97,8'd236} : s = 333;
	{8'd97,8'd237} : s = 334;
	{8'd97,8'd238} : s = 335;
	{8'd97,8'd239} : s = 336;
	{8'd97,8'd240} : s = 337;
	{8'd97,8'd241} : s = 338;
	{8'd97,8'd242} : s = 339;
	{8'd97,8'd243} : s = 340;
	{8'd97,8'd244} : s = 341;
	{8'd97,8'd245} : s = 342;
	{8'd97,8'd246} : s = 343;
	{8'd97,8'd247} : s = 344;
	{8'd97,8'd248} : s = 345;
	{8'd97,8'd249} : s = 346;
	{8'd97,8'd250} : s = 347;
	{8'd97,8'd251} : s = 348;
	{8'd97,8'd252} : s = 349;
	{8'd97,8'd253} : s = 350;
	{8'd97,8'd254} : s = 351;
	{8'd97,8'd255} : s = 352;
	{8'd98,8'd0} : s = 98;
	{8'd98,8'd1} : s = 99;
	{8'd98,8'd2} : s = 100;
	{8'd98,8'd3} : s = 101;
	{8'd98,8'd4} : s = 102;
	{8'd98,8'd5} : s = 103;
	{8'd98,8'd6} : s = 104;
	{8'd98,8'd7} : s = 105;
	{8'd98,8'd8} : s = 106;
	{8'd98,8'd9} : s = 107;
	{8'd98,8'd10} : s = 108;
	{8'd98,8'd11} : s = 109;
	{8'd98,8'd12} : s = 110;
	{8'd98,8'd13} : s = 111;
	{8'd98,8'd14} : s = 112;
	{8'd98,8'd15} : s = 113;
	{8'd98,8'd16} : s = 114;
	{8'd98,8'd17} : s = 115;
	{8'd98,8'd18} : s = 116;
	{8'd98,8'd19} : s = 117;
	{8'd98,8'd20} : s = 118;
	{8'd98,8'd21} : s = 119;
	{8'd98,8'd22} : s = 120;
	{8'd98,8'd23} : s = 121;
	{8'd98,8'd24} : s = 122;
	{8'd98,8'd25} : s = 123;
	{8'd98,8'd26} : s = 124;
	{8'd98,8'd27} : s = 125;
	{8'd98,8'd28} : s = 126;
	{8'd98,8'd29} : s = 127;
	{8'd98,8'd30} : s = 128;
	{8'd98,8'd31} : s = 129;
	{8'd98,8'd32} : s = 130;
	{8'd98,8'd33} : s = 131;
	{8'd98,8'd34} : s = 132;
	{8'd98,8'd35} : s = 133;
	{8'd98,8'd36} : s = 134;
	{8'd98,8'd37} : s = 135;
	{8'd98,8'd38} : s = 136;
	{8'd98,8'd39} : s = 137;
	{8'd98,8'd40} : s = 138;
	{8'd98,8'd41} : s = 139;
	{8'd98,8'd42} : s = 140;
	{8'd98,8'd43} : s = 141;
	{8'd98,8'd44} : s = 142;
	{8'd98,8'd45} : s = 143;
	{8'd98,8'd46} : s = 144;
	{8'd98,8'd47} : s = 145;
	{8'd98,8'd48} : s = 146;
	{8'd98,8'd49} : s = 147;
	{8'd98,8'd50} : s = 148;
	{8'd98,8'd51} : s = 149;
	{8'd98,8'd52} : s = 150;
	{8'd98,8'd53} : s = 151;
	{8'd98,8'd54} : s = 152;
	{8'd98,8'd55} : s = 153;
	{8'd98,8'd56} : s = 154;
	{8'd98,8'd57} : s = 155;
	{8'd98,8'd58} : s = 156;
	{8'd98,8'd59} : s = 157;
	{8'd98,8'd60} : s = 158;
	{8'd98,8'd61} : s = 159;
	{8'd98,8'd62} : s = 160;
	{8'd98,8'd63} : s = 161;
	{8'd98,8'd64} : s = 162;
	{8'd98,8'd65} : s = 163;
	{8'd98,8'd66} : s = 164;
	{8'd98,8'd67} : s = 165;
	{8'd98,8'd68} : s = 166;
	{8'd98,8'd69} : s = 167;
	{8'd98,8'd70} : s = 168;
	{8'd98,8'd71} : s = 169;
	{8'd98,8'd72} : s = 170;
	{8'd98,8'd73} : s = 171;
	{8'd98,8'd74} : s = 172;
	{8'd98,8'd75} : s = 173;
	{8'd98,8'd76} : s = 174;
	{8'd98,8'd77} : s = 175;
	{8'd98,8'd78} : s = 176;
	{8'd98,8'd79} : s = 177;
	{8'd98,8'd80} : s = 178;
	{8'd98,8'd81} : s = 179;
	{8'd98,8'd82} : s = 180;
	{8'd98,8'd83} : s = 181;
	{8'd98,8'd84} : s = 182;
	{8'd98,8'd85} : s = 183;
	{8'd98,8'd86} : s = 184;
	{8'd98,8'd87} : s = 185;
	{8'd98,8'd88} : s = 186;
	{8'd98,8'd89} : s = 187;
	{8'd98,8'd90} : s = 188;
	{8'd98,8'd91} : s = 189;
	{8'd98,8'd92} : s = 190;
	{8'd98,8'd93} : s = 191;
	{8'd98,8'd94} : s = 192;
	{8'd98,8'd95} : s = 193;
	{8'd98,8'd96} : s = 194;
	{8'd98,8'd97} : s = 195;
	{8'd98,8'd98} : s = 196;
	{8'd98,8'd99} : s = 197;
	{8'd98,8'd100} : s = 198;
	{8'd98,8'd101} : s = 199;
	{8'd98,8'd102} : s = 200;
	{8'd98,8'd103} : s = 201;
	{8'd98,8'd104} : s = 202;
	{8'd98,8'd105} : s = 203;
	{8'd98,8'd106} : s = 204;
	{8'd98,8'd107} : s = 205;
	{8'd98,8'd108} : s = 206;
	{8'd98,8'd109} : s = 207;
	{8'd98,8'd110} : s = 208;
	{8'd98,8'd111} : s = 209;
	{8'd98,8'd112} : s = 210;
	{8'd98,8'd113} : s = 211;
	{8'd98,8'd114} : s = 212;
	{8'd98,8'd115} : s = 213;
	{8'd98,8'd116} : s = 214;
	{8'd98,8'd117} : s = 215;
	{8'd98,8'd118} : s = 216;
	{8'd98,8'd119} : s = 217;
	{8'd98,8'd120} : s = 218;
	{8'd98,8'd121} : s = 219;
	{8'd98,8'd122} : s = 220;
	{8'd98,8'd123} : s = 221;
	{8'd98,8'd124} : s = 222;
	{8'd98,8'd125} : s = 223;
	{8'd98,8'd126} : s = 224;
	{8'd98,8'd127} : s = 225;
	{8'd98,8'd128} : s = 226;
	{8'd98,8'd129} : s = 227;
	{8'd98,8'd130} : s = 228;
	{8'd98,8'd131} : s = 229;
	{8'd98,8'd132} : s = 230;
	{8'd98,8'd133} : s = 231;
	{8'd98,8'd134} : s = 232;
	{8'd98,8'd135} : s = 233;
	{8'd98,8'd136} : s = 234;
	{8'd98,8'd137} : s = 235;
	{8'd98,8'd138} : s = 236;
	{8'd98,8'd139} : s = 237;
	{8'd98,8'd140} : s = 238;
	{8'd98,8'd141} : s = 239;
	{8'd98,8'd142} : s = 240;
	{8'd98,8'd143} : s = 241;
	{8'd98,8'd144} : s = 242;
	{8'd98,8'd145} : s = 243;
	{8'd98,8'd146} : s = 244;
	{8'd98,8'd147} : s = 245;
	{8'd98,8'd148} : s = 246;
	{8'd98,8'd149} : s = 247;
	{8'd98,8'd150} : s = 248;
	{8'd98,8'd151} : s = 249;
	{8'd98,8'd152} : s = 250;
	{8'd98,8'd153} : s = 251;
	{8'd98,8'd154} : s = 252;
	{8'd98,8'd155} : s = 253;
	{8'd98,8'd156} : s = 254;
	{8'd98,8'd157} : s = 255;
	{8'd98,8'd158} : s = 256;
	{8'd98,8'd159} : s = 257;
	{8'd98,8'd160} : s = 258;
	{8'd98,8'd161} : s = 259;
	{8'd98,8'd162} : s = 260;
	{8'd98,8'd163} : s = 261;
	{8'd98,8'd164} : s = 262;
	{8'd98,8'd165} : s = 263;
	{8'd98,8'd166} : s = 264;
	{8'd98,8'd167} : s = 265;
	{8'd98,8'd168} : s = 266;
	{8'd98,8'd169} : s = 267;
	{8'd98,8'd170} : s = 268;
	{8'd98,8'd171} : s = 269;
	{8'd98,8'd172} : s = 270;
	{8'd98,8'd173} : s = 271;
	{8'd98,8'd174} : s = 272;
	{8'd98,8'd175} : s = 273;
	{8'd98,8'd176} : s = 274;
	{8'd98,8'd177} : s = 275;
	{8'd98,8'd178} : s = 276;
	{8'd98,8'd179} : s = 277;
	{8'd98,8'd180} : s = 278;
	{8'd98,8'd181} : s = 279;
	{8'd98,8'd182} : s = 280;
	{8'd98,8'd183} : s = 281;
	{8'd98,8'd184} : s = 282;
	{8'd98,8'd185} : s = 283;
	{8'd98,8'd186} : s = 284;
	{8'd98,8'd187} : s = 285;
	{8'd98,8'd188} : s = 286;
	{8'd98,8'd189} : s = 287;
	{8'd98,8'd190} : s = 288;
	{8'd98,8'd191} : s = 289;
	{8'd98,8'd192} : s = 290;
	{8'd98,8'd193} : s = 291;
	{8'd98,8'd194} : s = 292;
	{8'd98,8'd195} : s = 293;
	{8'd98,8'd196} : s = 294;
	{8'd98,8'd197} : s = 295;
	{8'd98,8'd198} : s = 296;
	{8'd98,8'd199} : s = 297;
	{8'd98,8'd200} : s = 298;
	{8'd98,8'd201} : s = 299;
	{8'd98,8'd202} : s = 300;
	{8'd98,8'd203} : s = 301;
	{8'd98,8'd204} : s = 302;
	{8'd98,8'd205} : s = 303;
	{8'd98,8'd206} : s = 304;
	{8'd98,8'd207} : s = 305;
	{8'd98,8'd208} : s = 306;
	{8'd98,8'd209} : s = 307;
	{8'd98,8'd210} : s = 308;
	{8'd98,8'd211} : s = 309;
	{8'd98,8'd212} : s = 310;
	{8'd98,8'd213} : s = 311;
	{8'd98,8'd214} : s = 312;
	{8'd98,8'd215} : s = 313;
	{8'd98,8'd216} : s = 314;
	{8'd98,8'd217} : s = 315;
	{8'd98,8'd218} : s = 316;
	{8'd98,8'd219} : s = 317;
	{8'd98,8'd220} : s = 318;
	{8'd98,8'd221} : s = 319;
	{8'd98,8'd222} : s = 320;
	{8'd98,8'd223} : s = 321;
	{8'd98,8'd224} : s = 322;
	{8'd98,8'd225} : s = 323;
	{8'd98,8'd226} : s = 324;
	{8'd98,8'd227} : s = 325;
	{8'd98,8'd228} : s = 326;
	{8'd98,8'd229} : s = 327;
	{8'd98,8'd230} : s = 328;
	{8'd98,8'd231} : s = 329;
	{8'd98,8'd232} : s = 330;
	{8'd98,8'd233} : s = 331;
	{8'd98,8'd234} : s = 332;
	{8'd98,8'd235} : s = 333;
	{8'd98,8'd236} : s = 334;
	{8'd98,8'd237} : s = 335;
	{8'd98,8'd238} : s = 336;
	{8'd98,8'd239} : s = 337;
	{8'd98,8'd240} : s = 338;
	{8'd98,8'd241} : s = 339;
	{8'd98,8'd242} : s = 340;
	{8'd98,8'd243} : s = 341;
	{8'd98,8'd244} : s = 342;
	{8'd98,8'd245} : s = 343;
	{8'd98,8'd246} : s = 344;
	{8'd98,8'd247} : s = 345;
	{8'd98,8'd248} : s = 346;
	{8'd98,8'd249} : s = 347;
	{8'd98,8'd250} : s = 348;
	{8'd98,8'd251} : s = 349;
	{8'd98,8'd252} : s = 350;
	{8'd98,8'd253} : s = 351;
	{8'd98,8'd254} : s = 352;
	{8'd98,8'd255} : s = 353;
	{8'd99,8'd0} : s = 99;
	{8'd99,8'd1} : s = 100;
	{8'd99,8'd2} : s = 101;
	{8'd99,8'd3} : s = 102;
	{8'd99,8'd4} : s = 103;
	{8'd99,8'd5} : s = 104;
	{8'd99,8'd6} : s = 105;
	{8'd99,8'd7} : s = 106;
	{8'd99,8'd8} : s = 107;
	{8'd99,8'd9} : s = 108;
	{8'd99,8'd10} : s = 109;
	{8'd99,8'd11} : s = 110;
	{8'd99,8'd12} : s = 111;
	{8'd99,8'd13} : s = 112;
	{8'd99,8'd14} : s = 113;
	{8'd99,8'd15} : s = 114;
	{8'd99,8'd16} : s = 115;
	{8'd99,8'd17} : s = 116;
	{8'd99,8'd18} : s = 117;
	{8'd99,8'd19} : s = 118;
	{8'd99,8'd20} : s = 119;
	{8'd99,8'd21} : s = 120;
	{8'd99,8'd22} : s = 121;
	{8'd99,8'd23} : s = 122;
	{8'd99,8'd24} : s = 123;
	{8'd99,8'd25} : s = 124;
	{8'd99,8'd26} : s = 125;
	{8'd99,8'd27} : s = 126;
	{8'd99,8'd28} : s = 127;
	{8'd99,8'd29} : s = 128;
	{8'd99,8'd30} : s = 129;
	{8'd99,8'd31} : s = 130;
	{8'd99,8'd32} : s = 131;
	{8'd99,8'd33} : s = 132;
	{8'd99,8'd34} : s = 133;
	{8'd99,8'd35} : s = 134;
	{8'd99,8'd36} : s = 135;
	{8'd99,8'd37} : s = 136;
	{8'd99,8'd38} : s = 137;
	{8'd99,8'd39} : s = 138;
	{8'd99,8'd40} : s = 139;
	{8'd99,8'd41} : s = 140;
	{8'd99,8'd42} : s = 141;
	{8'd99,8'd43} : s = 142;
	{8'd99,8'd44} : s = 143;
	{8'd99,8'd45} : s = 144;
	{8'd99,8'd46} : s = 145;
	{8'd99,8'd47} : s = 146;
	{8'd99,8'd48} : s = 147;
	{8'd99,8'd49} : s = 148;
	{8'd99,8'd50} : s = 149;
	{8'd99,8'd51} : s = 150;
	{8'd99,8'd52} : s = 151;
	{8'd99,8'd53} : s = 152;
	{8'd99,8'd54} : s = 153;
	{8'd99,8'd55} : s = 154;
	{8'd99,8'd56} : s = 155;
	{8'd99,8'd57} : s = 156;
	{8'd99,8'd58} : s = 157;
	{8'd99,8'd59} : s = 158;
	{8'd99,8'd60} : s = 159;
	{8'd99,8'd61} : s = 160;
	{8'd99,8'd62} : s = 161;
	{8'd99,8'd63} : s = 162;
	{8'd99,8'd64} : s = 163;
	{8'd99,8'd65} : s = 164;
	{8'd99,8'd66} : s = 165;
	{8'd99,8'd67} : s = 166;
	{8'd99,8'd68} : s = 167;
	{8'd99,8'd69} : s = 168;
	{8'd99,8'd70} : s = 169;
	{8'd99,8'd71} : s = 170;
	{8'd99,8'd72} : s = 171;
	{8'd99,8'd73} : s = 172;
	{8'd99,8'd74} : s = 173;
	{8'd99,8'd75} : s = 174;
	{8'd99,8'd76} : s = 175;
	{8'd99,8'd77} : s = 176;
	{8'd99,8'd78} : s = 177;
	{8'd99,8'd79} : s = 178;
	{8'd99,8'd80} : s = 179;
	{8'd99,8'd81} : s = 180;
	{8'd99,8'd82} : s = 181;
	{8'd99,8'd83} : s = 182;
	{8'd99,8'd84} : s = 183;
	{8'd99,8'd85} : s = 184;
	{8'd99,8'd86} : s = 185;
	{8'd99,8'd87} : s = 186;
	{8'd99,8'd88} : s = 187;
	{8'd99,8'd89} : s = 188;
	{8'd99,8'd90} : s = 189;
	{8'd99,8'd91} : s = 190;
	{8'd99,8'd92} : s = 191;
	{8'd99,8'd93} : s = 192;
	{8'd99,8'd94} : s = 193;
	{8'd99,8'd95} : s = 194;
	{8'd99,8'd96} : s = 195;
	{8'd99,8'd97} : s = 196;
	{8'd99,8'd98} : s = 197;
	{8'd99,8'd99} : s = 198;
	{8'd99,8'd100} : s = 199;
	{8'd99,8'd101} : s = 200;
	{8'd99,8'd102} : s = 201;
	{8'd99,8'd103} : s = 202;
	{8'd99,8'd104} : s = 203;
	{8'd99,8'd105} : s = 204;
	{8'd99,8'd106} : s = 205;
	{8'd99,8'd107} : s = 206;
	{8'd99,8'd108} : s = 207;
	{8'd99,8'd109} : s = 208;
	{8'd99,8'd110} : s = 209;
	{8'd99,8'd111} : s = 210;
	{8'd99,8'd112} : s = 211;
	{8'd99,8'd113} : s = 212;
	{8'd99,8'd114} : s = 213;
	{8'd99,8'd115} : s = 214;
	{8'd99,8'd116} : s = 215;
	{8'd99,8'd117} : s = 216;
	{8'd99,8'd118} : s = 217;
	{8'd99,8'd119} : s = 218;
	{8'd99,8'd120} : s = 219;
	{8'd99,8'd121} : s = 220;
	{8'd99,8'd122} : s = 221;
	{8'd99,8'd123} : s = 222;
	{8'd99,8'd124} : s = 223;
	{8'd99,8'd125} : s = 224;
	{8'd99,8'd126} : s = 225;
	{8'd99,8'd127} : s = 226;
	{8'd99,8'd128} : s = 227;
	{8'd99,8'd129} : s = 228;
	{8'd99,8'd130} : s = 229;
	{8'd99,8'd131} : s = 230;
	{8'd99,8'd132} : s = 231;
	{8'd99,8'd133} : s = 232;
	{8'd99,8'd134} : s = 233;
	{8'd99,8'd135} : s = 234;
	{8'd99,8'd136} : s = 235;
	{8'd99,8'd137} : s = 236;
	{8'd99,8'd138} : s = 237;
	{8'd99,8'd139} : s = 238;
	{8'd99,8'd140} : s = 239;
	{8'd99,8'd141} : s = 240;
	{8'd99,8'd142} : s = 241;
	{8'd99,8'd143} : s = 242;
	{8'd99,8'd144} : s = 243;
	{8'd99,8'd145} : s = 244;
	{8'd99,8'd146} : s = 245;
	{8'd99,8'd147} : s = 246;
	{8'd99,8'd148} : s = 247;
	{8'd99,8'd149} : s = 248;
	{8'd99,8'd150} : s = 249;
	{8'd99,8'd151} : s = 250;
	{8'd99,8'd152} : s = 251;
	{8'd99,8'd153} : s = 252;
	{8'd99,8'd154} : s = 253;
	{8'd99,8'd155} : s = 254;
	{8'd99,8'd156} : s = 255;
	{8'd99,8'd157} : s = 256;
	{8'd99,8'd158} : s = 257;
	{8'd99,8'd159} : s = 258;
	{8'd99,8'd160} : s = 259;
	{8'd99,8'd161} : s = 260;
	{8'd99,8'd162} : s = 261;
	{8'd99,8'd163} : s = 262;
	{8'd99,8'd164} : s = 263;
	{8'd99,8'd165} : s = 264;
	{8'd99,8'd166} : s = 265;
	{8'd99,8'd167} : s = 266;
	{8'd99,8'd168} : s = 267;
	{8'd99,8'd169} : s = 268;
	{8'd99,8'd170} : s = 269;
	{8'd99,8'd171} : s = 270;
	{8'd99,8'd172} : s = 271;
	{8'd99,8'd173} : s = 272;
	{8'd99,8'd174} : s = 273;
	{8'd99,8'd175} : s = 274;
	{8'd99,8'd176} : s = 275;
	{8'd99,8'd177} : s = 276;
	{8'd99,8'd178} : s = 277;
	{8'd99,8'd179} : s = 278;
	{8'd99,8'd180} : s = 279;
	{8'd99,8'd181} : s = 280;
	{8'd99,8'd182} : s = 281;
	{8'd99,8'd183} : s = 282;
	{8'd99,8'd184} : s = 283;
	{8'd99,8'd185} : s = 284;
	{8'd99,8'd186} : s = 285;
	{8'd99,8'd187} : s = 286;
	{8'd99,8'd188} : s = 287;
	{8'd99,8'd189} : s = 288;
	{8'd99,8'd190} : s = 289;
	{8'd99,8'd191} : s = 290;
	{8'd99,8'd192} : s = 291;
	{8'd99,8'd193} : s = 292;
	{8'd99,8'd194} : s = 293;
	{8'd99,8'd195} : s = 294;
	{8'd99,8'd196} : s = 295;
	{8'd99,8'd197} : s = 296;
	{8'd99,8'd198} : s = 297;
	{8'd99,8'd199} : s = 298;
	{8'd99,8'd200} : s = 299;
	{8'd99,8'd201} : s = 300;
	{8'd99,8'd202} : s = 301;
	{8'd99,8'd203} : s = 302;
	{8'd99,8'd204} : s = 303;
	{8'd99,8'd205} : s = 304;
	{8'd99,8'd206} : s = 305;
	{8'd99,8'd207} : s = 306;
	{8'd99,8'd208} : s = 307;
	{8'd99,8'd209} : s = 308;
	{8'd99,8'd210} : s = 309;
	{8'd99,8'd211} : s = 310;
	{8'd99,8'd212} : s = 311;
	{8'd99,8'd213} : s = 312;
	{8'd99,8'd214} : s = 313;
	{8'd99,8'd215} : s = 314;
	{8'd99,8'd216} : s = 315;
	{8'd99,8'd217} : s = 316;
	{8'd99,8'd218} : s = 317;
	{8'd99,8'd219} : s = 318;
	{8'd99,8'd220} : s = 319;
	{8'd99,8'd221} : s = 320;
	{8'd99,8'd222} : s = 321;
	{8'd99,8'd223} : s = 322;
	{8'd99,8'd224} : s = 323;
	{8'd99,8'd225} : s = 324;
	{8'd99,8'd226} : s = 325;
	{8'd99,8'd227} : s = 326;
	{8'd99,8'd228} : s = 327;
	{8'd99,8'd229} : s = 328;
	{8'd99,8'd230} : s = 329;
	{8'd99,8'd231} : s = 330;
	{8'd99,8'd232} : s = 331;
	{8'd99,8'd233} : s = 332;
	{8'd99,8'd234} : s = 333;
	{8'd99,8'd235} : s = 334;
	{8'd99,8'd236} : s = 335;
	{8'd99,8'd237} : s = 336;
	{8'd99,8'd238} : s = 337;
	{8'd99,8'd239} : s = 338;
	{8'd99,8'd240} : s = 339;
	{8'd99,8'd241} : s = 340;
	{8'd99,8'd242} : s = 341;
	{8'd99,8'd243} : s = 342;
	{8'd99,8'd244} : s = 343;
	{8'd99,8'd245} : s = 344;
	{8'd99,8'd246} : s = 345;
	{8'd99,8'd247} : s = 346;
	{8'd99,8'd248} : s = 347;
	{8'd99,8'd249} : s = 348;
	{8'd99,8'd250} : s = 349;
	{8'd99,8'd251} : s = 350;
	{8'd99,8'd252} : s = 351;
	{8'd99,8'd253} : s = 352;
	{8'd99,8'd254} : s = 353;
	{8'd99,8'd255} : s = 354;
	{8'd100,8'd0} : s = 100;
	{8'd100,8'd1} : s = 101;
	{8'd100,8'd2} : s = 102;
	{8'd100,8'd3} : s = 103;
	{8'd100,8'd4} : s = 104;
	{8'd100,8'd5} : s = 105;
	{8'd100,8'd6} : s = 106;
	{8'd100,8'd7} : s = 107;
	{8'd100,8'd8} : s = 108;
	{8'd100,8'd9} : s = 109;
	{8'd100,8'd10} : s = 110;
	{8'd100,8'd11} : s = 111;
	{8'd100,8'd12} : s = 112;
	{8'd100,8'd13} : s = 113;
	{8'd100,8'd14} : s = 114;
	{8'd100,8'd15} : s = 115;
	{8'd100,8'd16} : s = 116;
	{8'd100,8'd17} : s = 117;
	{8'd100,8'd18} : s = 118;
	{8'd100,8'd19} : s = 119;
	{8'd100,8'd20} : s = 120;
	{8'd100,8'd21} : s = 121;
	{8'd100,8'd22} : s = 122;
	{8'd100,8'd23} : s = 123;
	{8'd100,8'd24} : s = 124;
	{8'd100,8'd25} : s = 125;
	{8'd100,8'd26} : s = 126;
	{8'd100,8'd27} : s = 127;
	{8'd100,8'd28} : s = 128;
	{8'd100,8'd29} : s = 129;
	{8'd100,8'd30} : s = 130;
	{8'd100,8'd31} : s = 131;
	{8'd100,8'd32} : s = 132;
	{8'd100,8'd33} : s = 133;
	{8'd100,8'd34} : s = 134;
	{8'd100,8'd35} : s = 135;
	{8'd100,8'd36} : s = 136;
	{8'd100,8'd37} : s = 137;
	{8'd100,8'd38} : s = 138;
	{8'd100,8'd39} : s = 139;
	{8'd100,8'd40} : s = 140;
	{8'd100,8'd41} : s = 141;
	{8'd100,8'd42} : s = 142;
	{8'd100,8'd43} : s = 143;
	{8'd100,8'd44} : s = 144;
	{8'd100,8'd45} : s = 145;
	{8'd100,8'd46} : s = 146;
	{8'd100,8'd47} : s = 147;
	{8'd100,8'd48} : s = 148;
	{8'd100,8'd49} : s = 149;
	{8'd100,8'd50} : s = 150;
	{8'd100,8'd51} : s = 151;
	{8'd100,8'd52} : s = 152;
	{8'd100,8'd53} : s = 153;
	{8'd100,8'd54} : s = 154;
	{8'd100,8'd55} : s = 155;
	{8'd100,8'd56} : s = 156;
	{8'd100,8'd57} : s = 157;
	{8'd100,8'd58} : s = 158;
	{8'd100,8'd59} : s = 159;
	{8'd100,8'd60} : s = 160;
	{8'd100,8'd61} : s = 161;
	{8'd100,8'd62} : s = 162;
	{8'd100,8'd63} : s = 163;
	{8'd100,8'd64} : s = 164;
	{8'd100,8'd65} : s = 165;
	{8'd100,8'd66} : s = 166;
	{8'd100,8'd67} : s = 167;
	{8'd100,8'd68} : s = 168;
	{8'd100,8'd69} : s = 169;
	{8'd100,8'd70} : s = 170;
	{8'd100,8'd71} : s = 171;
	{8'd100,8'd72} : s = 172;
	{8'd100,8'd73} : s = 173;
	{8'd100,8'd74} : s = 174;
	{8'd100,8'd75} : s = 175;
	{8'd100,8'd76} : s = 176;
	{8'd100,8'd77} : s = 177;
	{8'd100,8'd78} : s = 178;
	{8'd100,8'd79} : s = 179;
	{8'd100,8'd80} : s = 180;
	{8'd100,8'd81} : s = 181;
	{8'd100,8'd82} : s = 182;
	{8'd100,8'd83} : s = 183;
	{8'd100,8'd84} : s = 184;
	{8'd100,8'd85} : s = 185;
	{8'd100,8'd86} : s = 186;
	{8'd100,8'd87} : s = 187;
	{8'd100,8'd88} : s = 188;
	{8'd100,8'd89} : s = 189;
	{8'd100,8'd90} : s = 190;
	{8'd100,8'd91} : s = 191;
	{8'd100,8'd92} : s = 192;
	{8'd100,8'd93} : s = 193;
	{8'd100,8'd94} : s = 194;
	{8'd100,8'd95} : s = 195;
	{8'd100,8'd96} : s = 196;
	{8'd100,8'd97} : s = 197;
	{8'd100,8'd98} : s = 198;
	{8'd100,8'd99} : s = 199;
	{8'd100,8'd100} : s = 200;
	{8'd100,8'd101} : s = 201;
	{8'd100,8'd102} : s = 202;
	{8'd100,8'd103} : s = 203;
	{8'd100,8'd104} : s = 204;
	{8'd100,8'd105} : s = 205;
	{8'd100,8'd106} : s = 206;
	{8'd100,8'd107} : s = 207;
	{8'd100,8'd108} : s = 208;
	{8'd100,8'd109} : s = 209;
	{8'd100,8'd110} : s = 210;
	{8'd100,8'd111} : s = 211;
	{8'd100,8'd112} : s = 212;
	{8'd100,8'd113} : s = 213;
	{8'd100,8'd114} : s = 214;
	{8'd100,8'd115} : s = 215;
	{8'd100,8'd116} : s = 216;
	{8'd100,8'd117} : s = 217;
	{8'd100,8'd118} : s = 218;
	{8'd100,8'd119} : s = 219;
	{8'd100,8'd120} : s = 220;
	{8'd100,8'd121} : s = 221;
	{8'd100,8'd122} : s = 222;
	{8'd100,8'd123} : s = 223;
	{8'd100,8'd124} : s = 224;
	{8'd100,8'd125} : s = 225;
	{8'd100,8'd126} : s = 226;
	{8'd100,8'd127} : s = 227;
	{8'd100,8'd128} : s = 228;
	{8'd100,8'd129} : s = 229;
	{8'd100,8'd130} : s = 230;
	{8'd100,8'd131} : s = 231;
	{8'd100,8'd132} : s = 232;
	{8'd100,8'd133} : s = 233;
	{8'd100,8'd134} : s = 234;
	{8'd100,8'd135} : s = 235;
	{8'd100,8'd136} : s = 236;
	{8'd100,8'd137} : s = 237;
	{8'd100,8'd138} : s = 238;
	{8'd100,8'd139} : s = 239;
	{8'd100,8'd140} : s = 240;
	{8'd100,8'd141} : s = 241;
	{8'd100,8'd142} : s = 242;
	{8'd100,8'd143} : s = 243;
	{8'd100,8'd144} : s = 244;
	{8'd100,8'd145} : s = 245;
	{8'd100,8'd146} : s = 246;
	{8'd100,8'd147} : s = 247;
	{8'd100,8'd148} : s = 248;
	{8'd100,8'd149} : s = 249;
	{8'd100,8'd150} : s = 250;
	{8'd100,8'd151} : s = 251;
	{8'd100,8'd152} : s = 252;
	{8'd100,8'd153} : s = 253;
	{8'd100,8'd154} : s = 254;
	{8'd100,8'd155} : s = 255;
	{8'd100,8'd156} : s = 256;
	{8'd100,8'd157} : s = 257;
	{8'd100,8'd158} : s = 258;
	{8'd100,8'd159} : s = 259;
	{8'd100,8'd160} : s = 260;
	{8'd100,8'd161} : s = 261;
	{8'd100,8'd162} : s = 262;
	{8'd100,8'd163} : s = 263;
	{8'd100,8'd164} : s = 264;
	{8'd100,8'd165} : s = 265;
	{8'd100,8'd166} : s = 266;
	{8'd100,8'd167} : s = 267;
	{8'd100,8'd168} : s = 268;
	{8'd100,8'd169} : s = 269;
	{8'd100,8'd170} : s = 270;
	{8'd100,8'd171} : s = 271;
	{8'd100,8'd172} : s = 272;
	{8'd100,8'd173} : s = 273;
	{8'd100,8'd174} : s = 274;
	{8'd100,8'd175} : s = 275;
	{8'd100,8'd176} : s = 276;
	{8'd100,8'd177} : s = 277;
	{8'd100,8'd178} : s = 278;
	{8'd100,8'd179} : s = 279;
	{8'd100,8'd180} : s = 280;
	{8'd100,8'd181} : s = 281;
	{8'd100,8'd182} : s = 282;
	{8'd100,8'd183} : s = 283;
	{8'd100,8'd184} : s = 284;
	{8'd100,8'd185} : s = 285;
	{8'd100,8'd186} : s = 286;
	{8'd100,8'd187} : s = 287;
	{8'd100,8'd188} : s = 288;
	{8'd100,8'd189} : s = 289;
	{8'd100,8'd190} : s = 290;
	{8'd100,8'd191} : s = 291;
	{8'd100,8'd192} : s = 292;
	{8'd100,8'd193} : s = 293;
	{8'd100,8'd194} : s = 294;
	{8'd100,8'd195} : s = 295;
	{8'd100,8'd196} : s = 296;
	{8'd100,8'd197} : s = 297;
	{8'd100,8'd198} : s = 298;
	{8'd100,8'd199} : s = 299;
	{8'd100,8'd200} : s = 300;
	{8'd100,8'd201} : s = 301;
	{8'd100,8'd202} : s = 302;
	{8'd100,8'd203} : s = 303;
	{8'd100,8'd204} : s = 304;
	{8'd100,8'd205} : s = 305;
	{8'd100,8'd206} : s = 306;
	{8'd100,8'd207} : s = 307;
	{8'd100,8'd208} : s = 308;
	{8'd100,8'd209} : s = 309;
	{8'd100,8'd210} : s = 310;
	{8'd100,8'd211} : s = 311;
	{8'd100,8'd212} : s = 312;
	{8'd100,8'd213} : s = 313;
	{8'd100,8'd214} : s = 314;
	{8'd100,8'd215} : s = 315;
	{8'd100,8'd216} : s = 316;
	{8'd100,8'd217} : s = 317;
	{8'd100,8'd218} : s = 318;
	{8'd100,8'd219} : s = 319;
	{8'd100,8'd220} : s = 320;
	{8'd100,8'd221} : s = 321;
	{8'd100,8'd222} : s = 322;
	{8'd100,8'd223} : s = 323;
	{8'd100,8'd224} : s = 324;
	{8'd100,8'd225} : s = 325;
	{8'd100,8'd226} : s = 326;
	{8'd100,8'd227} : s = 327;
	{8'd100,8'd228} : s = 328;
	{8'd100,8'd229} : s = 329;
	{8'd100,8'd230} : s = 330;
	{8'd100,8'd231} : s = 331;
	{8'd100,8'd232} : s = 332;
	{8'd100,8'd233} : s = 333;
	{8'd100,8'd234} : s = 334;
	{8'd100,8'd235} : s = 335;
	{8'd100,8'd236} : s = 336;
	{8'd100,8'd237} : s = 337;
	{8'd100,8'd238} : s = 338;
	{8'd100,8'd239} : s = 339;
	{8'd100,8'd240} : s = 340;
	{8'd100,8'd241} : s = 341;
	{8'd100,8'd242} : s = 342;
	{8'd100,8'd243} : s = 343;
	{8'd100,8'd244} : s = 344;
	{8'd100,8'd245} : s = 345;
	{8'd100,8'd246} : s = 346;
	{8'd100,8'd247} : s = 347;
	{8'd100,8'd248} : s = 348;
	{8'd100,8'd249} : s = 349;
	{8'd100,8'd250} : s = 350;
	{8'd100,8'd251} : s = 351;
	{8'd100,8'd252} : s = 352;
	{8'd100,8'd253} : s = 353;
	{8'd100,8'd254} : s = 354;
	{8'd100,8'd255} : s = 355;
	{8'd101,8'd0} : s = 101;
	{8'd101,8'd1} : s = 102;
	{8'd101,8'd2} : s = 103;
	{8'd101,8'd3} : s = 104;
	{8'd101,8'd4} : s = 105;
	{8'd101,8'd5} : s = 106;
	{8'd101,8'd6} : s = 107;
	{8'd101,8'd7} : s = 108;
	{8'd101,8'd8} : s = 109;
	{8'd101,8'd9} : s = 110;
	{8'd101,8'd10} : s = 111;
	{8'd101,8'd11} : s = 112;
	{8'd101,8'd12} : s = 113;
	{8'd101,8'd13} : s = 114;
	{8'd101,8'd14} : s = 115;
	{8'd101,8'd15} : s = 116;
	{8'd101,8'd16} : s = 117;
	{8'd101,8'd17} : s = 118;
	{8'd101,8'd18} : s = 119;
	{8'd101,8'd19} : s = 120;
	{8'd101,8'd20} : s = 121;
	{8'd101,8'd21} : s = 122;
	{8'd101,8'd22} : s = 123;
	{8'd101,8'd23} : s = 124;
	{8'd101,8'd24} : s = 125;
	{8'd101,8'd25} : s = 126;
	{8'd101,8'd26} : s = 127;
	{8'd101,8'd27} : s = 128;
	{8'd101,8'd28} : s = 129;
	{8'd101,8'd29} : s = 130;
	{8'd101,8'd30} : s = 131;
	{8'd101,8'd31} : s = 132;
	{8'd101,8'd32} : s = 133;
	{8'd101,8'd33} : s = 134;
	{8'd101,8'd34} : s = 135;
	{8'd101,8'd35} : s = 136;
	{8'd101,8'd36} : s = 137;
	{8'd101,8'd37} : s = 138;
	{8'd101,8'd38} : s = 139;
	{8'd101,8'd39} : s = 140;
	{8'd101,8'd40} : s = 141;
	{8'd101,8'd41} : s = 142;
	{8'd101,8'd42} : s = 143;
	{8'd101,8'd43} : s = 144;
	{8'd101,8'd44} : s = 145;
	{8'd101,8'd45} : s = 146;
	{8'd101,8'd46} : s = 147;
	{8'd101,8'd47} : s = 148;
	{8'd101,8'd48} : s = 149;
	{8'd101,8'd49} : s = 150;
	{8'd101,8'd50} : s = 151;
	{8'd101,8'd51} : s = 152;
	{8'd101,8'd52} : s = 153;
	{8'd101,8'd53} : s = 154;
	{8'd101,8'd54} : s = 155;
	{8'd101,8'd55} : s = 156;
	{8'd101,8'd56} : s = 157;
	{8'd101,8'd57} : s = 158;
	{8'd101,8'd58} : s = 159;
	{8'd101,8'd59} : s = 160;
	{8'd101,8'd60} : s = 161;
	{8'd101,8'd61} : s = 162;
	{8'd101,8'd62} : s = 163;
	{8'd101,8'd63} : s = 164;
	{8'd101,8'd64} : s = 165;
	{8'd101,8'd65} : s = 166;
	{8'd101,8'd66} : s = 167;
	{8'd101,8'd67} : s = 168;
	{8'd101,8'd68} : s = 169;
	{8'd101,8'd69} : s = 170;
	{8'd101,8'd70} : s = 171;
	{8'd101,8'd71} : s = 172;
	{8'd101,8'd72} : s = 173;
	{8'd101,8'd73} : s = 174;
	{8'd101,8'd74} : s = 175;
	{8'd101,8'd75} : s = 176;
	{8'd101,8'd76} : s = 177;
	{8'd101,8'd77} : s = 178;
	{8'd101,8'd78} : s = 179;
	{8'd101,8'd79} : s = 180;
	{8'd101,8'd80} : s = 181;
	{8'd101,8'd81} : s = 182;
	{8'd101,8'd82} : s = 183;
	{8'd101,8'd83} : s = 184;
	{8'd101,8'd84} : s = 185;
	{8'd101,8'd85} : s = 186;
	{8'd101,8'd86} : s = 187;
	{8'd101,8'd87} : s = 188;
	{8'd101,8'd88} : s = 189;
	{8'd101,8'd89} : s = 190;
	{8'd101,8'd90} : s = 191;
	{8'd101,8'd91} : s = 192;
	{8'd101,8'd92} : s = 193;
	{8'd101,8'd93} : s = 194;
	{8'd101,8'd94} : s = 195;
	{8'd101,8'd95} : s = 196;
	{8'd101,8'd96} : s = 197;
	{8'd101,8'd97} : s = 198;
	{8'd101,8'd98} : s = 199;
	{8'd101,8'd99} : s = 200;
	{8'd101,8'd100} : s = 201;
	{8'd101,8'd101} : s = 202;
	{8'd101,8'd102} : s = 203;
	{8'd101,8'd103} : s = 204;
	{8'd101,8'd104} : s = 205;
	{8'd101,8'd105} : s = 206;
	{8'd101,8'd106} : s = 207;
	{8'd101,8'd107} : s = 208;
	{8'd101,8'd108} : s = 209;
	{8'd101,8'd109} : s = 210;
	{8'd101,8'd110} : s = 211;
	{8'd101,8'd111} : s = 212;
	{8'd101,8'd112} : s = 213;
	{8'd101,8'd113} : s = 214;
	{8'd101,8'd114} : s = 215;
	{8'd101,8'd115} : s = 216;
	{8'd101,8'd116} : s = 217;
	{8'd101,8'd117} : s = 218;
	{8'd101,8'd118} : s = 219;
	{8'd101,8'd119} : s = 220;
	{8'd101,8'd120} : s = 221;
	{8'd101,8'd121} : s = 222;
	{8'd101,8'd122} : s = 223;
	{8'd101,8'd123} : s = 224;
	{8'd101,8'd124} : s = 225;
	{8'd101,8'd125} : s = 226;
	{8'd101,8'd126} : s = 227;
	{8'd101,8'd127} : s = 228;
	{8'd101,8'd128} : s = 229;
	{8'd101,8'd129} : s = 230;
	{8'd101,8'd130} : s = 231;
	{8'd101,8'd131} : s = 232;
	{8'd101,8'd132} : s = 233;
	{8'd101,8'd133} : s = 234;
	{8'd101,8'd134} : s = 235;
	{8'd101,8'd135} : s = 236;
	{8'd101,8'd136} : s = 237;
	{8'd101,8'd137} : s = 238;
	{8'd101,8'd138} : s = 239;
	{8'd101,8'd139} : s = 240;
	{8'd101,8'd140} : s = 241;
	{8'd101,8'd141} : s = 242;
	{8'd101,8'd142} : s = 243;
	{8'd101,8'd143} : s = 244;
	{8'd101,8'd144} : s = 245;
	{8'd101,8'd145} : s = 246;
	{8'd101,8'd146} : s = 247;
	{8'd101,8'd147} : s = 248;
	{8'd101,8'd148} : s = 249;
	{8'd101,8'd149} : s = 250;
	{8'd101,8'd150} : s = 251;
	{8'd101,8'd151} : s = 252;
	{8'd101,8'd152} : s = 253;
	{8'd101,8'd153} : s = 254;
	{8'd101,8'd154} : s = 255;
	{8'd101,8'd155} : s = 256;
	{8'd101,8'd156} : s = 257;
	{8'd101,8'd157} : s = 258;
	{8'd101,8'd158} : s = 259;
	{8'd101,8'd159} : s = 260;
	{8'd101,8'd160} : s = 261;
	{8'd101,8'd161} : s = 262;
	{8'd101,8'd162} : s = 263;
	{8'd101,8'd163} : s = 264;
	{8'd101,8'd164} : s = 265;
	{8'd101,8'd165} : s = 266;
	{8'd101,8'd166} : s = 267;
	{8'd101,8'd167} : s = 268;
	{8'd101,8'd168} : s = 269;
	{8'd101,8'd169} : s = 270;
	{8'd101,8'd170} : s = 271;
	{8'd101,8'd171} : s = 272;
	{8'd101,8'd172} : s = 273;
	{8'd101,8'd173} : s = 274;
	{8'd101,8'd174} : s = 275;
	{8'd101,8'd175} : s = 276;
	{8'd101,8'd176} : s = 277;
	{8'd101,8'd177} : s = 278;
	{8'd101,8'd178} : s = 279;
	{8'd101,8'd179} : s = 280;
	{8'd101,8'd180} : s = 281;
	{8'd101,8'd181} : s = 282;
	{8'd101,8'd182} : s = 283;
	{8'd101,8'd183} : s = 284;
	{8'd101,8'd184} : s = 285;
	{8'd101,8'd185} : s = 286;
	{8'd101,8'd186} : s = 287;
	{8'd101,8'd187} : s = 288;
	{8'd101,8'd188} : s = 289;
	{8'd101,8'd189} : s = 290;
	{8'd101,8'd190} : s = 291;
	{8'd101,8'd191} : s = 292;
	{8'd101,8'd192} : s = 293;
	{8'd101,8'd193} : s = 294;
	{8'd101,8'd194} : s = 295;
	{8'd101,8'd195} : s = 296;
	{8'd101,8'd196} : s = 297;
	{8'd101,8'd197} : s = 298;
	{8'd101,8'd198} : s = 299;
	{8'd101,8'd199} : s = 300;
	{8'd101,8'd200} : s = 301;
	{8'd101,8'd201} : s = 302;
	{8'd101,8'd202} : s = 303;
	{8'd101,8'd203} : s = 304;
	{8'd101,8'd204} : s = 305;
	{8'd101,8'd205} : s = 306;
	{8'd101,8'd206} : s = 307;
	{8'd101,8'd207} : s = 308;
	{8'd101,8'd208} : s = 309;
	{8'd101,8'd209} : s = 310;
	{8'd101,8'd210} : s = 311;
	{8'd101,8'd211} : s = 312;
	{8'd101,8'd212} : s = 313;
	{8'd101,8'd213} : s = 314;
	{8'd101,8'd214} : s = 315;
	{8'd101,8'd215} : s = 316;
	{8'd101,8'd216} : s = 317;
	{8'd101,8'd217} : s = 318;
	{8'd101,8'd218} : s = 319;
	{8'd101,8'd219} : s = 320;
	{8'd101,8'd220} : s = 321;
	{8'd101,8'd221} : s = 322;
	{8'd101,8'd222} : s = 323;
	{8'd101,8'd223} : s = 324;
	{8'd101,8'd224} : s = 325;
	{8'd101,8'd225} : s = 326;
	{8'd101,8'd226} : s = 327;
	{8'd101,8'd227} : s = 328;
	{8'd101,8'd228} : s = 329;
	{8'd101,8'd229} : s = 330;
	{8'd101,8'd230} : s = 331;
	{8'd101,8'd231} : s = 332;
	{8'd101,8'd232} : s = 333;
	{8'd101,8'd233} : s = 334;
	{8'd101,8'd234} : s = 335;
	{8'd101,8'd235} : s = 336;
	{8'd101,8'd236} : s = 337;
	{8'd101,8'd237} : s = 338;
	{8'd101,8'd238} : s = 339;
	{8'd101,8'd239} : s = 340;
	{8'd101,8'd240} : s = 341;
	{8'd101,8'd241} : s = 342;
	{8'd101,8'd242} : s = 343;
	{8'd101,8'd243} : s = 344;
	{8'd101,8'd244} : s = 345;
	{8'd101,8'd245} : s = 346;
	{8'd101,8'd246} : s = 347;
	{8'd101,8'd247} : s = 348;
	{8'd101,8'd248} : s = 349;
	{8'd101,8'd249} : s = 350;
	{8'd101,8'd250} : s = 351;
	{8'd101,8'd251} : s = 352;
	{8'd101,8'd252} : s = 353;
	{8'd101,8'd253} : s = 354;
	{8'd101,8'd254} : s = 355;
	{8'd101,8'd255} : s = 356;
	{8'd102,8'd0} : s = 102;
	{8'd102,8'd1} : s = 103;
	{8'd102,8'd2} : s = 104;
	{8'd102,8'd3} : s = 105;
	{8'd102,8'd4} : s = 106;
	{8'd102,8'd5} : s = 107;
	{8'd102,8'd6} : s = 108;
	{8'd102,8'd7} : s = 109;
	{8'd102,8'd8} : s = 110;
	{8'd102,8'd9} : s = 111;
	{8'd102,8'd10} : s = 112;
	{8'd102,8'd11} : s = 113;
	{8'd102,8'd12} : s = 114;
	{8'd102,8'd13} : s = 115;
	{8'd102,8'd14} : s = 116;
	{8'd102,8'd15} : s = 117;
	{8'd102,8'd16} : s = 118;
	{8'd102,8'd17} : s = 119;
	{8'd102,8'd18} : s = 120;
	{8'd102,8'd19} : s = 121;
	{8'd102,8'd20} : s = 122;
	{8'd102,8'd21} : s = 123;
	{8'd102,8'd22} : s = 124;
	{8'd102,8'd23} : s = 125;
	{8'd102,8'd24} : s = 126;
	{8'd102,8'd25} : s = 127;
	{8'd102,8'd26} : s = 128;
	{8'd102,8'd27} : s = 129;
	{8'd102,8'd28} : s = 130;
	{8'd102,8'd29} : s = 131;
	{8'd102,8'd30} : s = 132;
	{8'd102,8'd31} : s = 133;
	{8'd102,8'd32} : s = 134;
	{8'd102,8'd33} : s = 135;
	{8'd102,8'd34} : s = 136;
	{8'd102,8'd35} : s = 137;
	{8'd102,8'd36} : s = 138;
	{8'd102,8'd37} : s = 139;
	{8'd102,8'd38} : s = 140;
	{8'd102,8'd39} : s = 141;
	{8'd102,8'd40} : s = 142;
	{8'd102,8'd41} : s = 143;
	{8'd102,8'd42} : s = 144;
	{8'd102,8'd43} : s = 145;
	{8'd102,8'd44} : s = 146;
	{8'd102,8'd45} : s = 147;
	{8'd102,8'd46} : s = 148;
	{8'd102,8'd47} : s = 149;
	{8'd102,8'd48} : s = 150;
	{8'd102,8'd49} : s = 151;
	{8'd102,8'd50} : s = 152;
	{8'd102,8'd51} : s = 153;
	{8'd102,8'd52} : s = 154;
	{8'd102,8'd53} : s = 155;
	{8'd102,8'd54} : s = 156;
	{8'd102,8'd55} : s = 157;
	{8'd102,8'd56} : s = 158;
	{8'd102,8'd57} : s = 159;
	{8'd102,8'd58} : s = 160;
	{8'd102,8'd59} : s = 161;
	{8'd102,8'd60} : s = 162;
	{8'd102,8'd61} : s = 163;
	{8'd102,8'd62} : s = 164;
	{8'd102,8'd63} : s = 165;
	{8'd102,8'd64} : s = 166;
	{8'd102,8'd65} : s = 167;
	{8'd102,8'd66} : s = 168;
	{8'd102,8'd67} : s = 169;
	{8'd102,8'd68} : s = 170;
	{8'd102,8'd69} : s = 171;
	{8'd102,8'd70} : s = 172;
	{8'd102,8'd71} : s = 173;
	{8'd102,8'd72} : s = 174;
	{8'd102,8'd73} : s = 175;
	{8'd102,8'd74} : s = 176;
	{8'd102,8'd75} : s = 177;
	{8'd102,8'd76} : s = 178;
	{8'd102,8'd77} : s = 179;
	{8'd102,8'd78} : s = 180;
	{8'd102,8'd79} : s = 181;
	{8'd102,8'd80} : s = 182;
	{8'd102,8'd81} : s = 183;
	{8'd102,8'd82} : s = 184;
	{8'd102,8'd83} : s = 185;
	{8'd102,8'd84} : s = 186;
	{8'd102,8'd85} : s = 187;
	{8'd102,8'd86} : s = 188;
	{8'd102,8'd87} : s = 189;
	{8'd102,8'd88} : s = 190;
	{8'd102,8'd89} : s = 191;
	{8'd102,8'd90} : s = 192;
	{8'd102,8'd91} : s = 193;
	{8'd102,8'd92} : s = 194;
	{8'd102,8'd93} : s = 195;
	{8'd102,8'd94} : s = 196;
	{8'd102,8'd95} : s = 197;
	{8'd102,8'd96} : s = 198;
	{8'd102,8'd97} : s = 199;
	{8'd102,8'd98} : s = 200;
	{8'd102,8'd99} : s = 201;
	{8'd102,8'd100} : s = 202;
	{8'd102,8'd101} : s = 203;
	{8'd102,8'd102} : s = 204;
	{8'd102,8'd103} : s = 205;
	{8'd102,8'd104} : s = 206;
	{8'd102,8'd105} : s = 207;
	{8'd102,8'd106} : s = 208;
	{8'd102,8'd107} : s = 209;
	{8'd102,8'd108} : s = 210;
	{8'd102,8'd109} : s = 211;
	{8'd102,8'd110} : s = 212;
	{8'd102,8'd111} : s = 213;
	{8'd102,8'd112} : s = 214;
	{8'd102,8'd113} : s = 215;
	{8'd102,8'd114} : s = 216;
	{8'd102,8'd115} : s = 217;
	{8'd102,8'd116} : s = 218;
	{8'd102,8'd117} : s = 219;
	{8'd102,8'd118} : s = 220;
	{8'd102,8'd119} : s = 221;
	{8'd102,8'd120} : s = 222;
	{8'd102,8'd121} : s = 223;
	{8'd102,8'd122} : s = 224;
	{8'd102,8'd123} : s = 225;
	{8'd102,8'd124} : s = 226;
	{8'd102,8'd125} : s = 227;
	{8'd102,8'd126} : s = 228;
	{8'd102,8'd127} : s = 229;
	{8'd102,8'd128} : s = 230;
	{8'd102,8'd129} : s = 231;
	{8'd102,8'd130} : s = 232;
	{8'd102,8'd131} : s = 233;
	{8'd102,8'd132} : s = 234;
	{8'd102,8'd133} : s = 235;
	{8'd102,8'd134} : s = 236;
	{8'd102,8'd135} : s = 237;
	{8'd102,8'd136} : s = 238;
	{8'd102,8'd137} : s = 239;
	{8'd102,8'd138} : s = 240;
	{8'd102,8'd139} : s = 241;
	{8'd102,8'd140} : s = 242;
	{8'd102,8'd141} : s = 243;
	{8'd102,8'd142} : s = 244;
	{8'd102,8'd143} : s = 245;
	{8'd102,8'd144} : s = 246;
	{8'd102,8'd145} : s = 247;
	{8'd102,8'd146} : s = 248;
	{8'd102,8'd147} : s = 249;
	{8'd102,8'd148} : s = 250;
	{8'd102,8'd149} : s = 251;
	{8'd102,8'd150} : s = 252;
	{8'd102,8'd151} : s = 253;
	{8'd102,8'd152} : s = 254;
	{8'd102,8'd153} : s = 255;
	{8'd102,8'd154} : s = 256;
	{8'd102,8'd155} : s = 257;
	{8'd102,8'd156} : s = 258;
	{8'd102,8'd157} : s = 259;
	{8'd102,8'd158} : s = 260;
	{8'd102,8'd159} : s = 261;
	{8'd102,8'd160} : s = 262;
	{8'd102,8'd161} : s = 263;
	{8'd102,8'd162} : s = 264;
	{8'd102,8'd163} : s = 265;
	{8'd102,8'd164} : s = 266;
	{8'd102,8'd165} : s = 267;
	{8'd102,8'd166} : s = 268;
	{8'd102,8'd167} : s = 269;
	{8'd102,8'd168} : s = 270;
	{8'd102,8'd169} : s = 271;
	{8'd102,8'd170} : s = 272;
	{8'd102,8'd171} : s = 273;
	{8'd102,8'd172} : s = 274;
	{8'd102,8'd173} : s = 275;
	{8'd102,8'd174} : s = 276;
	{8'd102,8'd175} : s = 277;
	{8'd102,8'd176} : s = 278;
	{8'd102,8'd177} : s = 279;
	{8'd102,8'd178} : s = 280;
	{8'd102,8'd179} : s = 281;
	{8'd102,8'd180} : s = 282;
	{8'd102,8'd181} : s = 283;
	{8'd102,8'd182} : s = 284;
	{8'd102,8'd183} : s = 285;
	{8'd102,8'd184} : s = 286;
	{8'd102,8'd185} : s = 287;
	{8'd102,8'd186} : s = 288;
	{8'd102,8'd187} : s = 289;
	{8'd102,8'd188} : s = 290;
	{8'd102,8'd189} : s = 291;
	{8'd102,8'd190} : s = 292;
	{8'd102,8'd191} : s = 293;
	{8'd102,8'd192} : s = 294;
	{8'd102,8'd193} : s = 295;
	{8'd102,8'd194} : s = 296;
	{8'd102,8'd195} : s = 297;
	{8'd102,8'd196} : s = 298;
	{8'd102,8'd197} : s = 299;
	{8'd102,8'd198} : s = 300;
	{8'd102,8'd199} : s = 301;
	{8'd102,8'd200} : s = 302;
	{8'd102,8'd201} : s = 303;
	{8'd102,8'd202} : s = 304;
	{8'd102,8'd203} : s = 305;
	{8'd102,8'd204} : s = 306;
	{8'd102,8'd205} : s = 307;
	{8'd102,8'd206} : s = 308;
	{8'd102,8'd207} : s = 309;
	{8'd102,8'd208} : s = 310;
	{8'd102,8'd209} : s = 311;
	{8'd102,8'd210} : s = 312;
	{8'd102,8'd211} : s = 313;
	{8'd102,8'd212} : s = 314;
	{8'd102,8'd213} : s = 315;
	{8'd102,8'd214} : s = 316;
	{8'd102,8'd215} : s = 317;
	{8'd102,8'd216} : s = 318;
	{8'd102,8'd217} : s = 319;
	{8'd102,8'd218} : s = 320;
	{8'd102,8'd219} : s = 321;
	{8'd102,8'd220} : s = 322;
	{8'd102,8'd221} : s = 323;
	{8'd102,8'd222} : s = 324;
	{8'd102,8'd223} : s = 325;
	{8'd102,8'd224} : s = 326;
	{8'd102,8'd225} : s = 327;
	{8'd102,8'd226} : s = 328;
	{8'd102,8'd227} : s = 329;
	{8'd102,8'd228} : s = 330;
	{8'd102,8'd229} : s = 331;
	{8'd102,8'd230} : s = 332;
	{8'd102,8'd231} : s = 333;
	{8'd102,8'd232} : s = 334;
	{8'd102,8'd233} : s = 335;
	{8'd102,8'd234} : s = 336;
	{8'd102,8'd235} : s = 337;
	{8'd102,8'd236} : s = 338;
	{8'd102,8'd237} : s = 339;
	{8'd102,8'd238} : s = 340;
	{8'd102,8'd239} : s = 341;
	{8'd102,8'd240} : s = 342;
	{8'd102,8'd241} : s = 343;
	{8'd102,8'd242} : s = 344;
	{8'd102,8'd243} : s = 345;
	{8'd102,8'd244} : s = 346;
	{8'd102,8'd245} : s = 347;
	{8'd102,8'd246} : s = 348;
	{8'd102,8'd247} : s = 349;
	{8'd102,8'd248} : s = 350;
	{8'd102,8'd249} : s = 351;
	{8'd102,8'd250} : s = 352;
	{8'd102,8'd251} : s = 353;
	{8'd102,8'd252} : s = 354;
	{8'd102,8'd253} : s = 355;
	{8'd102,8'd254} : s = 356;
	{8'd102,8'd255} : s = 357;
	{8'd103,8'd0} : s = 103;
	{8'd103,8'd1} : s = 104;
	{8'd103,8'd2} : s = 105;
	{8'd103,8'd3} : s = 106;
	{8'd103,8'd4} : s = 107;
	{8'd103,8'd5} : s = 108;
	{8'd103,8'd6} : s = 109;
	{8'd103,8'd7} : s = 110;
	{8'd103,8'd8} : s = 111;
	{8'd103,8'd9} : s = 112;
	{8'd103,8'd10} : s = 113;
	{8'd103,8'd11} : s = 114;
	{8'd103,8'd12} : s = 115;
	{8'd103,8'd13} : s = 116;
	{8'd103,8'd14} : s = 117;
	{8'd103,8'd15} : s = 118;
	{8'd103,8'd16} : s = 119;
	{8'd103,8'd17} : s = 120;
	{8'd103,8'd18} : s = 121;
	{8'd103,8'd19} : s = 122;
	{8'd103,8'd20} : s = 123;
	{8'd103,8'd21} : s = 124;
	{8'd103,8'd22} : s = 125;
	{8'd103,8'd23} : s = 126;
	{8'd103,8'd24} : s = 127;
	{8'd103,8'd25} : s = 128;
	{8'd103,8'd26} : s = 129;
	{8'd103,8'd27} : s = 130;
	{8'd103,8'd28} : s = 131;
	{8'd103,8'd29} : s = 132;
	{8'd103,8'd30} : s = 133;
	{8'd103,8'd31} : s = 134;
	{8'd103,8'd32} : s = 135;
	{8'd103,8'd33} : s = 136;
	{8'd103,8'd34} : s = 137;
	{8'd103,8'd35} : s = 138;
	{8'd103,8'd36} : s = 139;
	{8'd103,8'd37} : s = 140;
	{8'd103,8'd38} : s = 141;
	{8'd103,8'd39} : s = 142;
	{8'd103,8'd40} : s = 143;
	{8'd103,8'd41} : s = 144;
	{8'd103,8'd42} : s = 145;
	{8'd103,8'd43} : s = 146;
	{8'd103,8'd44} : s = 147;
	{8'd103,8'd45} : s = 148;
	{8'd103,8'd46} : s = 149;
	{8'd103,8'd47} : s = 150;
	{8'd103,8'd48} : s = 151;
	{8'd103,8'd49} : s = 152;
	{8'd103,8'd50} : s = 153;
	{8'd103,8'd51} : s = 154;
	{8'd103,8'd52} : s = 155;
	{8'd103,8'd53} : s = 156;
	{8'd103,8'd54} : s = 157;
	{8'd103,8'd55} : s = 158;
	{8'd103,8'd56} : s = 159;
	{8'd103,8'd57} : s = 160;
	{8'd103,8'd58} : s = 161;
	{8'd103,8'd59} : s = 162;
	{8'd103,8'd60} : s = 163;
	{8'd103,8'd61} : s = 164;
	{8'd103,8'd62} : s = 165;
	{8'd103,8'd63} : s = 166;
	{8'd103,8'd64} : s = 167;
	{8'd103,8'd65} : s = 168;
	{8'd103,8'd66} : s = 169;
	{8'd103,8'd67} : s = 170;
	{8'd103,8'd68} : s = 171;
	{8'd103,8'd69} : s = 172;
	{8'd103,8'd70} : s = 173;
	{8'd103,8'd71} : s = 174;
	{8'd103,8'd72} : s = 175;
	{8'd103,8'd73} : s = 176;
	{8'd103,8'd74} : s = 177;
	{8'd103,8'd75} : s = 178;
	{8'd103,8'd76} : s = 179;
	{8'd103,8'd77} : s = 180;
	{8'd103,8'd78} : s = 181;
	{8'd103,8'd79} : s = 182;
	{8'd103,8'd80} : s = 183;
	{8'd103,8'd81} : s = 184;
	{8'd103,8'd82} : s = 185;
	{8'd103,8'd83} : s = 186;
	{8'd103,8'd84} : s = 187;
	{8'd103,8'd85} : s = 188;
	{8'd103,8'd86} : s = 189;
	{8'd103,8'd87} : s = 190;
	{8'd103,8'd88} : s = 191;
	{8'd103,8'd89} : s = 192;
	{8'd103,8'd90} : s = 193;
	{8'd103,8'd91} : s = 194;
	{8'd103,8'd92} : s = 195;
	{8'd103,8'd93} : s = 196;
	{8'd103,8'd94} : s = 197;
	{8'd103,8'd95} : s = 198;
	{8'd103,8'd96} : s = 199;
	{8'd103,8'd97} : s = 200;
	{8'd103,8'd98} : s = 201;
	{8'd103,8'd99} : s = 202;
	{8'd103,8'd100} : s = 203;
	{8'd103,8'd101} : s = 204;
	{8'd103,8'd102} : s = 205;
	{8'd103,8'd103} : s = 206;
	{8'd103,8'd104} : s = 207;
	{8'd103,8'd105} : s = 208;
	{8'd103,8'd106} : s = 209;
	{8'd103,8'd107} : s = 210;
	{8'd103,8'd108} : s = 211;
	{8'd103,8'd109} : s = 212;
	{8'd103,8'd110} : s = 213;
	{8'd103,8'd111} : s = 214;
	{8'd103,8'd112} : s = 215;
	{8'd103,8'd113} : s = 216;
	{8'd103,8'd114} : s = 217;
	{8'd103,8'd115} : s = 218;
	{8'd103,8'd116} : s = 219;
	{8'd103,8'd117} : s = 220;
	{8'd103,8'd118} : s = 221;
	{8'd103,8'd119} : s = 222;
	{8'd103,8'd120} : s = 223;
	{8'd103,8'd121} : s = 224;
	{8'd103,8'd122} : s = 225;
	{8'd103,8'd123} : s = 226;
	{8'd103,8'd124} : s = 227;
	{8'd103,8'd125} : s = 228;
	{8'd103,8'd126} : s = 229;
	{8'd103,8'd127} : s = 230;
	{8'd103,8'd128} : s = 231;
	{8'd103,8'd129} : s = 232;
	{8'd103,8'd130} : s = 233;
	{8'd103,8'd131} : s = 234;
	{8'd103,8'd132} : s = 235;
	{8'd103,8'd133} : s = 236;
	{8'd103,8'd134} : s = 237;
	{8'd103,8'd135} : s = 238;
	{8'd103,8'd136} : s = 239;
	{8'd103,8'd137} : s = 240;
	{8'd103,8'd138} : s = 241;
	{8'd103,8'd139} : s = 242;
	{8'd103,8'd140} : s = 243;
	{8'd103,8'd141} : s = 244;
	{8'd103,8'd142} : s = 245;
	{8'd103,8'd143} : s = 246;
	{8'd103,8'd144} : s = 247;
	{8'd103,8'd145} : s = 248;
	{8'd103,8'd146} : s = 249;
	{8'd103,8'd147} : s = 250;
	{8'd103,8'd148} : s = 251;
	{8'd103,8'd149} : s = 252;
	{8'd103,8'd150} : s = 253;
	{8'd103,8'd151} : s = 254;
	{8'd103,8'd152} : s = 255;
	{8'd103,8'd153} : s = 256;
	{8'd103,8'd154} : s = 257;
	{8'd103,8'd155} : s = 258;
	{8'd103,8'd156} : s = 259;
	{8'd103,8'd157} : s = 260;
	{8'd103,8'd158} : s = 261;
	{8'd103,8'd159} : s = 262;
	{8'd103,8'd160} : s = 263;
	{8'd103,8'd161} : s = 264;
	{8'd103,8'd162} : s = 265;
	{8'd103,8'd163} : s = 266;
	{8'd103,8'd164} : s = 267;
	{8'd103,8'd165} : s = 268;
	{8'd103,8'd166} : s = 269;
	{8'd103,8'd167} : s = 270;
	{8'd103,8'd168} : s = 271;
	{8'd103,8'd169} : s = 272;
	{8'd103,8'd170} : s = 273;
	{8'd103,8'd171} : s = 274;
	{8'd103,8'd172} : s = 275;
	{8'd103,8'd173} : s = 276;
	{8'd103,8'd174} : s = 277;
	{8'd103,8'd175} : s = 278;
	{8'd103,8'd176} : s = 279;
	{8'd103,8'd177} : s = 280;
	{8'd103,8'd178} : s = 281;
	{8'd103,8'd179} : s = 282;
	{8'd103,8'd180} : s = 283;
	{8'd103,8'd181} : s = 284;
	{8'd103,8'd182} : s = 285;
	{8'd103,8'd183} : s = 286;
	{8'd103,8'd184} : s = 287;
	{8'd103,8'd185} : s = 288;
	{8'd103,8'd186} : s = 289;
	{8'd103,8'd187} : s = 290;
	{8'd103,8'd188} : s = 291;
	{8'd103,8'd189} : s = 292;
	{8'd103,8'd190} : s = 293;
	{8'd103,8'd191} : s = 294;
	{8'd103,8'd192} : s = 295;
	{8'd103,8'd193} : s = 296;
	{8'd103,8'd194} : s = 297;
	{8'd103,8'd195} : s = 298;
	{8'd103,8'd196} : s = 299;
	{8'd103,8'd197} : s = 300;
	{8'd103,8'd198} : s = 301;
	{8'd103,8'd199} : s = 302;
	{8'd103,8'd200} : s = 303;
	{8'd103,8'd201} : s = 304;
	{8'd103,8'd202} : s = 305;
	{8'd103,8'd203} : s = 306;
	{8'd103,8'd204} : s = 307;
	{8'd103,8'd205} : s = 308;
	{8'd103,8'd206} : s = 309;
	{8'd103,8'd207} : s = 310;
	{8'd103,8'd208} : s = 311;
	{8'd103,8'd209} : s = 312;
	{8'd103,8'd210} : s = 313;
	{8'd103,8'd211} : s = 314;
	{8'd103,8'd212} : s = 315;
	{8'd103,8'd213} : s = 316;
	{8'd103,8'd214} : s = 317;
	{8'd103,8'd215} : s = 318;
	{8'd103,8'd216} : s = 319;
	{8'd103,8'd217} : s = 320;
	{8'd103,8'd218} : s = 321;
	{8'd103,8'd219} : s = 322;
	{8'd103,8'd220} : s = 323;
	{8'd103,8'd221} : s = 324;
	{8'd103,8'd222} : s = 325;
	{8'd103,8'd223} : s = 326;
	{8'd103,8'd224} : s = 327;
	{8'd103,8'd225} : s = 328;
	{8'd103,8'd226} : s = 329;
	{8'd103,8'd227} : s = 330;
	{8'd103,8'd228} : s = 331;
	{8'd103,8'd229} : s = 332;
	{8'd103,8'd230} : s = 333;
	{8'd103,8'd231} : s = 334;
	{8'd103,8'd232} : s = 335;
	{8'd103,8'd233} : s = 336;
	{8'd103,8'd234} : s = 337;
	{8'd103,8'd235} : s = 338;
	{8'd103,8'd236} : s = 339;
	{8'd103,8'd237} : s = 340;
	{8'd103,8'd238} : s = 341;
	{8'd103,8'd239} : s = 342;
	{8'd103,8'd240} : s = 343;
	{8'd103,8'd241} : s = 344;
	{8'd103,8'd242} : s = 345;
	{8'd103,8'd243} : s = 346;
	{8'd103,8'd244} : s = 347;
	{8'd103,8'd245} : s = 348;
	{8'd103,8'd246} : s = 349;
	{8'd103,8'd247} : s = 350;
	{8'd103,8'd248} : s = 351;
	{8'd103,8'd249} : s = 352;
	{8'd103,8'd250} : s = 353;
	{8'd103,8'd251} : s = 354;
	{8'd103,8'd252} : s = 355;
	{8'd103,8'd253} : s = 356;
	{8'd103,8'd254} : s = 357;
	{8'd103,8'd255} : s = 358;
	{8'd104,8'd0} : s = 104;
	{8'd104,8'd1} : s = 105;
	{8'd104,8'd2} : s = 106;
	{8'd104,8'd3} : s = 107;
	{8'd104,8'd4} : s = 108;
	{8'd104,8'd5} : s = 109;
	{8'd104,8'd6} : s = 110;
	{8'd104,8'd7} : s = 111;
	{8'd104,8'd8} : s = 112;
	{8'd104,8'd9} : s = 113;
	{8'd104,8'd10} : s = 114;
	{8'd104,8'd11} : s = 115;
	{8'd104,8'd12} : s = 116;
	{8'd104,8'd13} : s = 117;
	{8'd104,8'd14} : s = 118;
	{8'd104,8'd15} : s = 119;
	{8'd104,8'd16} : s = 120;
	{8'd104,8'd17} : s = 121;
	{8'd104,8'd18} : s = 122;
	{8'd104,8'd19} : s = 123;
	{8'd104,8'd20} : s = 124;
	{8'd104,8'd21} : s = 125;
	{8'd104,8'd22} : s = 126;
	{8'd104,8'd23} : s = 127;
	{8'd104,8'd24} : s = 128;
	{8'd104,8'd25} : s = 129;
	{8'd104,8'd26} : s = 130;
	{8'd104,8'd27} : s = 131;
	{8'd104,8'd28} : s = 132;
	{8'd104,8'd29} : s = 133;
	{8'd104,8'd30} : s = 134;
	{8'd104,8'd31} : s = 135;
	{8'd104,8'd32} : s = 136;
	{8'd104,8'd33} : s = 137;
	{8'd104,8'd34} : s = 138;
	{8'd104,8'd35} : s = 139;
	{8'd104,8'd36} : s = 140;
	{8'd104,8'd37} : s = 141;
	{8'd104,8'd38} : s = 142;
	{8'd104,8'd39} : s = 143;
	{8'd104,8'd40} : s = 144;
	{8'd104,8'd41} : s = 145;
	{8'd104,8'd42} : s = 146;
	{8'd104,8'd43} : s = 147;
	{8'd104,8'd44} : s = 148;
	{8'd104,8'd45} : s = 149;
	{8'd104,8'd46} : s = 150;
	{8'd104,8'd47} : s = 151;
	{8'd104,8'd48} : s = 152;
	{8'd104,8'd49} : s = 153;
	{8'd104,8'd50} : s = 154;
	{8'd104,8'd51} : s = 155;
	{8'd104,8'd52} : s = 156;
	{8'd104,8'd53} : s = 157;
	{8'd104,8'd54} : s = 158;
	{8'd104,8'd55} : s = 159;
	{8'd104,8'd56} : s = 160;
	{8'd104,8'd57} : s = 161;
	{8'd104,8'd58} : s = 162;
	{8'd104,8'd59} : s = 163;
	{8'd104,8'd60} : s = 164;
	{8'd104,8'd61} : s = 165;
	{8'd104,8'd62} : s = 166;
	{8'd104,8'd63} : s = 167;
	{8'd104,8'd64} : s = 168;
	{8'd104,8'd65} : s = 169;
	{8'd104,8'd66} : s = 170;
	{8'd104,8'd67} : s = 171;
	{8'd104,8'd68} : s = 172;
	{8'd104,8'd69} : s = 173;
	{8'd104,8'd70} : s = 174;
	{8'd104,8'd71} : s = 175;
	{8'd104,8'd72} : s = 176;
	{8'd104,8'd73} : s = 177;
	{8'd104,8'd74} : s = 178;
	{8'd104,8'd75} : s = 179;
	{8'd104,8'd76} : s = 180;
	{8'd104,8'd77} : s = 181;
	{8'd104,8'd78} : s = 182;
	{8'd104,8'd79} : s = 183;
	{8'd104,8'd80} : s = 184;
	{8'd104,8'd81} : s = 185;
	{8'd104,8'd82} : s = 186;
	{8'd104,8'd83} : s = 187;
	{8'd104,8'd84} : s = 188;
	{8'd104,8'd85} : s = 189;
	{8'd104,8'd86} : s = 190;
	{8'd104,8'd87} : s = 191;
	{8'd104,8'd88} : s = 192;
	{8'd104,8'd89} : s = 193;
	{8'd104,8'd90} : s = 194;
	{8'd104,8'd91} : s = 195;
	{8'd104,8'd92} : s = 196;
	{8'd104,8'd93} : s = 197;
	{8'd104,8'd94} : s = 198;
	{8'd104,8'd95} : s = 199;
	{8'd104,8'd96} : s = 200;
	{8'd104,8'd97} : s = 201;
	{8'd104,8'd98} : s = 202;
	{8'd104,8'd99} : s = 203;
	{8'd104,8'd100} : s = 204;
	{8'd104,8'd101} : s = 205;
	{8'd104,8'd102} : s = 206;
	{8'd104,8'd103} : s = 207;
	{8'd104,8'd104} : s = 208;
	{8'd104,8'd105} : s = 209;
	{8'd104,8'd106} : s = 210;
	{8'd104,8'd107} : s = 211;
	{8'd104,8'd108} : s = 212;
	{8'd104,8'd109} : s = 213;
	{8'd104,8'd110} : s = 214;
	{8'd104,8'd111} : s = 215;
	{8'd104,8'd112} : s = 216;
	{8'd104,8'd113} : s = 217;
	{8'd104,8'd114} : s = 218;
	{8'd104,8'd115} : s = 219;
	{8'd104,8'd116} : s = 220;
	{8'd104,8'd117} : s = 221;
	{8'd104,8'd118} : s = 222;
	{8'd104,8'd119} : s = 223;
	{8'd104,8'd120} : s = 224;
	{8'd104,8'd121} : s = 225;
	{8'd104,8'd122} : s = 226;
	{8'd104,8'd123} : s = 227;
	{8'd104,8'd124} : s = 228;
	{8'd104,8'd125} : s = 229;
	{8'd104,8'd126} : s = 230;
	{8'd104,8'd127} : s = 231;
	{8'd104,8'd128} : s = 232;
	{8'd104,8'd129} : s = 233;
	{8'd104,8'd130} : s = 234;
	{8'd104,8'd131} : s = 235;
	{8'd104,8'd132} : s = 236;
	{8'd104,8'd133} : s = 237;
	{8'd104,8'd134} : s = 238;
	{8'd104,8'd135} : s = 239;
	{8'd104,8'd136} : s = 240;
	{8'd104,8'd137} : s = 241;
	{8'd104,8'd138} : s = 242;
	{8'd104,8'd139} : s = 243;
	{8'd104,8'd140} : s = 244;
	{8'd104,8'd141} : s = 245;
	{8'd104,8'd142} : s = 246;
	{8'd104,8'd143} : s = 247;
	{8'd104,8'd144} : s = 248;
	{8'd104,8'd145} : s = 249;
	{8'd104,8'd146} : s = 250;
	{8'd104,8'd147} : s = 251;
	{8'd104,8'd148} : s = 252;
	{8'd104,8'd149} : s = 253;
	{8'd104,8'd150} : s = 254;
	{8'd104,8'd151} : s = 255;
	{8'd104,8'd152} : s = 256;
	{8'd104,8'd153} : s = 257;
	{8'd104,8'd154} : s = 258;
	{8'd104,8'd155} : s = 259;
	{8'd104,8'd156} : s = 260;
	{8'd104,8'd157} : s = 261;
	{8'd104,8'd158} : s = 262;
	{8'd104,8'd159} : s = 263;
	{8'd104,8'd160} : s = 264;
	{8'd104,8'd161} : s = 265;
	{8'd104,8'd162} : s = 266;
	{8'd104,8'd163} : s = 267;
	{8'd104,8'd164} : s = 268;
	{8'd104,8'd165} : s = 269;
	{8'd104,8'd166} : s = 270;
	{8'd104,8'd167} : s = 271;
	{8'd104,8'd168} : s = 272;
	{8'd104,8'd169} : s = 273;
	{8'd104,8'd170} : s = 274;
	{8'd104,8'd171} : s = 275;
	{8'd104,8'd172} : s = 276;
	{8'd104,8'd173} : s = 277;
	{8'd104,8'd174} : s = 278;
	{8'd104,8'd175} : s = 279;
	{8'd104,8'd176} : s = 280;
	{8'd104,8'd177} : s = 281;
	{8'd104,8'd178} : s = 282;
	{8'd104,8'd179} : s = 283;
	{8'd104,8'd180} : s = 284;
	{8'd104,8'd181} : s = 285;
	{8'd104,8'd182} : s = 286;
	{8'd104,8'd183} : s = 287;
	{8'd104,8'd184} : s = 288;
	{8'd104,8'd185} : s = 289;
	{8'd104,8'd186} : s = 290;
	{8'd104,8'd187} : s = 291;
	{8'd104,8'd188} : s = 292;
	{8'd104,8'd189} : s = 293;
	{8'd104,8'd190} : s = 294;
	{8'd104,8'd191} : s = 295;
	{8'd104,8'd192} : s = 296;
	{8'd104,8'd193} : s = 297;
	{8'd104,8'd194} : s = 298;
	{8'd104,8'd195} : s = 299;
	{8'd104,8'd196} : s = 300;
	{8'd104,8'd197} : s = 301;
	{8'd104,8'd198} : s = 302;
	{8'd104,8'd199} : s = 303;
	{8'd104,8'd200} : s = 304;
	{8'd104,8'd201} : s = 305;
	{8'd104,8'd202} : s = 306;
	{8'd104,8'd203} : s = 307;
	{8'd104,8'd204} : s = 308;
	{8'd104,8'd205} : s = 309;
	{8'd104,8'd206} : s = 310;
	{8'd104,8'd207} : s = 311;
	{8'd104,8'd208} : s = 312;
	{8'd104,8'd209} : s = 313;
	{8'd104,8'd210} : s = 314;
	{8'd104,8'd211} : s = 315;
	{8'd104,8'd212} : s = 316;
	{8'd104,8'd213} : s = 317;
	{8'd104,8'd214} : s = 318;
	{8'd104,8'd215} : s = 319;
	{8'd104,8'd216} : s = 320;
	{8'd104,8'd217} : s = 321;
	{8'd104,8'd218} : s = 322;
	{8'd104,8'd219} : s = 323;
	{8'd104,8'd220} : s = 324;
	{8'd104,8'd221} : s = 325;
	{8'd104,8'd222} : s = 326;
	{8'd104,8'd223} : s = 327;
	{8'd104,8'd224} : s = 328;
	{8'd104,8'd225} : s = 329;
	{8'd104,8'd226} : s = 330;
	{8'd104,8'd227} : s = 331;
	{8'd104,8'd228} : s = 332;
	{8'd104,8'd229} : s = 333;
	{8'd104,8'd230} : s = 334;
	{8'd104,8'd231} : s = 335;
	{8'd104,8'd232} : s = 336;
	{8'd104,8'd233} : s = 337;
	{8'd104,8'd234} : s = 338;
	{8'd104,8'd235} : s = 339;
	{8'd104,8'd236} : s = 340;
	{8'd104,8'd237} : s = 341;
	{8'd104,8'd238} : s = 342;
	{8'd104,8'd239} : s = 343;
	{8'd104,8'd240} : s = 344;
	{8'd104,8'd241} : s = 345;
	{8'd104,8'd242} : s = 346;
	{8'd104,8'd243} : s = 347;
	{8'd104,8'd244} : s = 348;
	{8'd104,8'd245} : s = 349;
	{8'd104,8'd246} : s = 350;
	{8'd104,8'd247} : s = 351;
	{8'd104,8'd248} : s = 352;
	{8'd104,8'd249} : s = 353;
	{8'd104,8'd250} : s = 354;
	{8'd104,8'd251} : s = 355;
	{8'd104,8'd252} : s = 356;
	{8'd104,8'd253} : s = 357;
	{8'd104,8'd254} : s = 358;
	{8'd104,8'd255} : s = 359;
	{8'd105,8'd0} : s = 105;
	{8'd105,8'd1} : s = 106;
	{8'd105,8'd2} : s = 107;
	{8'd105,8'd3} : s = 108;
	{8'd105,8'd4} : s = 109;
	{8'd105,8'd5} : s = 110;
	{8'd105,8'd6} : s = 111;
	{8'd105,8'd7} : s = 112;
	{8'd105,8'd8} : s = 113;
	{8'd105,8'd9} : s = 114;
	{8'd105,8'd10} : s = 115;
	{8'd105,8'd11} : s = 116;
	{8'd105,8'd12} : s = 117;
	{8'd105,8'd13} : s = 118;
	{8'd105,8'd14} : s = 119;
	{8'd105,8'd15} : s = 120;
	{8'd105,8'd16} : s = 121;
	{8'd105,8'd17} : s = 122;
	{8'd105,8'd18} : s = 123;
	{8'd105,8'd19} : s = 124;
	{8'd105,8'd20} : s = 125;
	{8'd105,8'd21} : s = 126;
	{8'd105,8'd22} : s = 127;
	{8'd105,8'd23} : s = 128;
	{8'd105,8'd24} : s = 129;
	{8'd105,8'd25} : s = 130;
	{8'd105,8'd26} : s = 131;
	{8'd105,8'd27} : s = 132;
	{8'd105,8'd28} : s = 133;
	{8'd105,8'd29} : s = 134;
	{8'd105,8'd30} : s = 135;
	{8'd105,8'd31} : s = 136;
	{8'd105,8'd32} : s = 137;
	{8'd105,8'd33} : s = 138;
	{8'd105,8'd34} : s = 139;
	{8'd105,8'd35} : s = 140;
	{8'd105,8'd36} : s = 141;
	{8'd105,8'd37} : s = 142;
	{8'd105,8'd38} : s = 143;
	{8'd105,8'd39} : s = 144;
	{8'd105,8'd40} : s = 145;
	{8'd105,8'd41} : s = 146;
	{8'd105,8'd42} : s = 147;
	{8'd105,8'd43} : s = 148;
	{8'd105,8'd44} : s = 149;
	{8'd105,8'd45} : s = 150;
	{8'd105,8'd46} : s = 151;
	{8'd105,8'd47} : s = 152;
	{8'd105,8'd48} : s = 153;
	{8'd105,8'd49} : s = 154;
	{8'd105,8'd50} : s = 155;
	{8'd105,8'd51} : s = 156;
	{8'd105,8'd52} : s = 157;
	{8'd105,8'd53} : s = 158;
	{8'd105,8'd54} : s = 159;
	{8'd105,8'd55} : s = 160;
	{8'd105,8'd56} : s = 161;
	{8'd105,8'd57} : s = 162;
	{8'd105,8'd58} : s = 163;
	{8'd105,8'd59} : s = 164;
	{8'd105,8'd60} : s = 165;
	{8'd105,8'd61} : s = 166;
	{8'd105,8'd62} : s = 167;
	{8'd105,8'd63} : s = 168;
	{8'd105,8'd64} : s = 169;
	{8'd105,8'd65} : s = 170;
	{8'd105,8'd66} : s = 171;
	{8'd105,8'd67} : s = 172;
	{8'd105,8'd68} : s = 173;
	{8'd105,8'd69} : s = 174;
	{8'd105,8'd70} : s = 175;
	{8'd105,8'd71} : s = 176;
	{8'd105,8'd72} : s = 177;
	{8'd105,8'd73} : s = 178;
	{8'd105,8'd74} : s = 179;
	{8'd105,8'd75} : s = 180;
	{8'd105,8'd76} : s = 181;
	{8'd105,8'd77} : s = 182;
	{8'd105,8'd78} : s = 183;
	{8'd105,8'd79} : s = 184;
	{8'd105,8'd80} : s = 185;
	{8'd105,8'd81} : s = 186;
	{8'd105,8'd82} : s = 187;
	{8'd105,8'd83} : s = 188;
	{8'd105,8'd84} : s = 189;
	{8'd105,8'd85} : s = 190;
	{8'd105,8'd86} : s = 191;
	{8'd105,8'd87} : s = 192;
	{8'd105,8'd88} : s = 193;
	{8'd105,8'd89} : s = 194;
	{8'd105,8'd90} : s = 195;
	{8'd105,8'd91} : s = 196;
	{8'd105,8'd92} : s = 197;
	{8'd105,8'd93} : s = 198;
	{8'd105,8'd94} : s = 199;
	{8'd105,8'd95} : s = 200;
	{8'd105,8'd96} : s = 201;
	{8'd105,8'd97} : s = 202;
	{8'd105,8'd98} : s = 203;
	{8'd105,8'd99} : s = 204;
	{8'd105,8'd100} : s = 205;
	{8'd105,8'd101} : s = 206;
	{8'd105,8'd102} : s = 207;
	{8'd105,8'd103} : s = 208;
	{8'd105,8'd104} : s = 209;
	{8'd105,8'd105} : s = 210;
	{8'd105,8'd106} : s = 211;
	{8'd105,8'd107} : s = 212;
	{8'd105,8'd108} : s = 213;
	{8'd105,8'd109} : s = 214;
	{8'd105,8'd110} : s = 215;
	{8'd105,8'd111} : s = 216;
	{8'd105,8'd112} : s = 217;
	{8'd105,8'd113} : s = 218;
	{8'd105,8'd114} : s = 219;
	{8'd105,8'd115} : s = 220;
	{8'd105,8'd116} : s = 221;
	{8'd105,8'd117} : s = 222;
	{8'd105,8'd118} : s = 223;
	{8'd105,8'd119} : s = 224;
	{8'd105,8'd120} : s = 225;
	{8'd105,8'd121} : s = 226;
	{8'd105,8'd122} : s = 227;
	{8'd105,8'd123} : s = 228;
	{8'd105,8'd124} : s = 229;
	{8'd105,8'd125} : s = 230;
	{8'd105,8'd126} : s = 231;
	{8'd105,8'd127} : s = 232;
	{8'd105,8'd128} : s = 233;
	{8'd105,8'd129} : s = 234;
	{8'd105,8'd130} : s = 235;
	{8'd105,8'd131} : s = 236;
	{8'd105,8'd132} : s = 237;
	{8'd105,8'd133} : s = 238;
	{8'd105,8'd134} : s = 239;
	{8'd105,8'd135} : s = 240;
	{8'd105,8'd136} : s = 241;
	{8'd105,8'd137} : s = 242;
	{8'd105,8'd138} : s = 243;
	{8'd105,8'd139} : s = 244;
	{8'd105,8'd140} : s = 245;
	{8'd105,8'd141} : s = 246;
	{8'd105,8'd142} : s = 247;
	{8'd105,8'd143} : s = 248;
	{8'd105,8'd144} : s = 249;
	{8'd105,8'd145} : s = 250;
	{8'd105,8'd146} : s = 251;
	{8'd105,8'd147} : s = 252;
	{8'd105,8'd148} : s = 253;
	{8'd105,8'd149} : s = 254;
	{8'd105,8'd150} : s = 255;
	{8'd105,8'd151} : s = 256;
	{8'd105,8'd152} : s = 257;
	{8'd105,8'd153} : s = 258;
	{8'd105,8'd154} : s = 259;
	{8'd105,8'd155} : s = 260;
	{8'd105,8'd156} : s = 261;
	{8'd105,8'd157} : s = 262;
	{8'd105,8'd158} : s = 263;
	{8'd105,8'd159} : s = 264;
	{8'd105,8'd160} : s = 265;
	{8'd105,8'd161} : s = 266;
	{8'd105,8'd162} : s = 267;
	{8'd105,8'd163} : s = 268;
	{8'd105,8'd164} : s = 269;
	{8'd105,8'd165} : s = 270;
	{8'd105,8'd166} : s = 271;
	{8'd105,8'd167} : s = 272;
	{8'd105,8'd168} : s = 273;
	{8'd105,8'd169} : s = 274;
	{8'd105,8'd170} : s = 275;
	{8'd105,8'd171} : s = 276;
	{8'd105,8'd172} : s = 277;
	{8'd105,8'd173} : s = 278;
	{8'd105,8'd174} : s = 279;
	{8'd105,8'd175} : s = 280;
	{8'd105,8'd176} : s = 281;
	{8'd105,8'd177} : s = 282;
	{8'd105,8'd178} : s = 283;
	{8'd105,8'd179} : s = 284;
	{8'd105,8'd180} : s = 285;
	{8'd105,8'd181} : s = 286;
	{8'd105,8'd182} : s = 287;
	{8'd105,8'd183} : s = 288;
	{8'd105,8'd184} : s = 289;
	{8'd105,8'd185} : s = 290;
	{8'd105,8'd186} : s = 291;
	{8'd105,8'd187} : s = 292;
	{8'd105,8'd188} : s = 293;
	{8'd105,8'd189} : s = 294;
	{8'd105,8'd190} : s = 295;
	{8'd105,8'd191} : s = 296;
	{8'd105,8'd192} : s = 297;
	{8'd105,8'd193} : s = 298;
	{8'd105,8'd194} : s = 299;
	{8'd105,8'd195} : s = 300;
	{8'd105,8'd196} : s = 301;
	{8'd105,8'd197} : s = 302;
	{8'd105,8'd198} : s = 303;
	{8'd105,8'd199} : s = 304;
	{8'd105,8'd200} : s = 305;
	{8'd105,8'd201} : s = 306;
	{8'd105,8'd202} : s = 307;
	{8'd105,8'd203} : s = 308;
	{8'd105,8'd204} : s = 309;
	{8'd105,8'd205} : s = 310;
	{8'd105,8'd206} : s = 311;
	{8'd105,8'd207} : s = 312;
	{8'd105,8'd208} : s = 313;
	{8'd105,8'd209} : s = 314;
	{8'd105,8'd210} : s = 315;
	{8'd105,8'd211} : s = 316;
	{8'd105,8'd212} : s = 317;
	{8'd105,8'd213} : s = 318;
	{8'd105,8'd214} : s = 319;
	{8'd105,8'd215} : s = 320;
	{8'd105,8'd216} : s = 321;
	{8'd105,8'd217} : s = 322;
	{8'd105,8'd218} : s = 323;
	{8'd105,8'd219} : s = 324;
	{8'd105,8'd220} : s = 325;
	{8'd105,8'd221} : s = 326;
	{8'd105,8'd222} : s = 327;
	{8'd105,8'd223} : s = 328;
	{8'd105,8'd224} : s = 329;
	{8'd105,8'd225} : s = 330;
	{8'd105,8'd226} : s = 331;
	{8'd105,8'd227} : s = 332;
	{8'd105,8'd228} : s = 333;
	{8'd105,8'd229} : s = 334;
	{8'd105,8'd230} : s = 335;
	{8'd105,8'd231} : s = 336;
	{8'd105,8'd232} : s = 337;
	{8'd105,8'd233} : s = 338;
	{8'd105,8'd234} : s = 339;
	{8'd105,8'd235} : s = 340;
	{8'd105,8'd236} : s = 341;
	{8'd105,8'd237} : s = 342;
	{8'd105,8'd238} : s = 343;
	{8'd105,8'd239} : s = 344;
	{8'd105,8'd240} : s = 345;
	{8'd105,8'd241} : s = 346;
	{8'd105,8'd242} : s = 347;
	{8'd105,8'd243} : s = 348;
	{8'd105,8'd244} : s = 349;
	{8'd105,8'd245} : s = 350;
	{8'd105,8'd246} : s = 351;
	{8'd105,8'd247} : s = 352;
	{8'd105,8'd248} : s = 353;
	{8'd105,8'd249} : s = 354;
	{8'd105,8'd250} : s = 355;
	{8'd105,8'd251} : s = 356;
	{8'd105,8'd252} : s = 357;
	{8'd105,8'd253} : s = 358;
	{8'd105,8'd254} : s = 359;
	{8'd105,8'd255} : s = 360;
	{8'd106,8'd0} : s = 106;
	{8'd106,8'd1} : s = 107;
	{8'd106,8'd2} : s = 108;
	{8'd106,8'd3} : s = 109;
	{8'd106,8'd4} : s = 110;
	{8'd106,8'd5} : s = 111;
	{8'd106,8'd6} : s = 112;
	{8'd106,8'd7} : s = 113;
	{8'd106,8'd8} : s = 114;
	{8'd106,8'd9} : s = 115;
	{8'd106,8'd10} : s = 116;
	{8'd106,8'd11} : s = 117;
	{8'd106,8'd12} : s = 118;
	{8'd106,8'd13} : s = 119;
	{8'd106,8'd14} : s = 120;
	{8'd106,8'd15} : s = 121;
	{8'd106,8'd16} : s = 122;
	{8'd106,8'd17} : s = 123;
	{8'd106,8'd18} : s = 124;
	{8'd106,8'd19} : s = 125;
	{8'd106,8'd20} : s = 126;
	{8'd106,8'd21} : s = 127;
	{8'd106,8'd22} : s = 128;
	{8'd106,8'd23} : s = 129;
	{8'd106,8'd24} : s = 130;
	{8'd106,8'd25} : s = 131;
	{8'd106,8'd26} : s = 132;
	{8'd106,8'd27} : s = 133;
	{8'd106,8'd28} : s = 134;
	{8'd106,8'd29} : s = 135;
	{8'd106,8'd30} : s = 136;
	{8'd106,8'd31} : s = 137;
	{8'd106,8'd32} : s = 138;
	{8'd106,8'd33} : s = 139;
	{8'd106,8'd34} : s = 140;
	{8'd106,8'd35} : s = 141;
	{8'd106,8'd36} : s = 142;
	{8'd106,8'd37} : s = 143;
	{8'd106,8'd38} : s = 144;
	{8'd106,8'd39} : s = 145;
	{8'd106,8'd40} : s = 146;
	{8'd106,8'd41} : s = 147;
	{8'd106,8'd42} : s = 148;
	{8'd106,8'd43} : s = 149;
	{8'd106,8'd44} : s = 150;
	{8'd106,8'd45} : s = 151;
	{8'd106,8'd46} : s = 152;
	{8'd106,8'd47} : s = 153;
	{8'd106,8'd48} : s = 154;
	{8'd106,8'd49} : s = 155;
	{8'd106,8'd50} : s = 156;
	{8'd106,8'd51} : s = 157;
	{8'd106,8'd52} : s = 158;
	{8'd106,8'd53} : s = 159;
	{8'd106,8'd54} : s = 160;
	{8'd106,8'd55} : s = 161;
	{8'd106,8'd56} : s = 162;
	{8'd106,8'd57} : s = 163;
	{8'd106,8'd58} : s = 164;
	{8'd106,8'd59} : s = 165;
	{8'd106,8'd60} : s = 166;
	{8'd106,8'd61} : s = 167;
	{8'd106,8'd62} : s = 168;
	{8'd106,8'd63} : s = 169;
	{8'd106,8'd64} : s = 170;
	{8'd106,8'd65} : s = 171;
	{8'd106,8'd66} : s = 172;
	{8'd106,8'd67} : s = 173;
	{8'd106,8'd68} : s = 174;
	{8'd106,8'd69} : s = 175;
	{8'd106,8'd70} : s = 176;
	{8'd106,8'd71} : s = 177;
	{8'd106,8'd72} : s = 178;
	{8'd106,8'd73} : s = 179;
	{8'd106,8'd74} : s = 180;
	{8'd106,8'd75} : s = 181;
	{8'd106,8'd76} : s = 182;
	{8'd106,8'd77} : s = 183;
	{8'd106,8'd78} : s = 184;
	{8'd106,8'd79} : s = 185;
	{8'd106,8'd80} : s = 186;
	{8'd106,8'd81} : s = 187;
	{8'd106,8'd82} : s = 188;
	{8'd106,8'd83} : s = 189;
	{8'd106,8'd84} : s = 190;
	{8'd106,8'd85} : s = 191;
	{8'd106,8'd86} : s = 192;
	{8'd106,8'd87} : s = 193;
	{8'd106,8'd88} : s = 194;
	{8'd106,8'd89} : s = 195;
	{8'd106,8'd90} : s = 196;
	{8'd106,8'd91} : s = 197;
	{8'd106,8'd92} : s = 198;
	{8'd106,8'd93} : s = 199;
	{8'd106,8'd94} : s = 200;
	{8'd106,8'd95} : s = 201;
	{8'd106,8'd96} : s = 202;
	{8'd106,8'd97} : s = 203;
	{8'd106,8'd98} : s = 204;
	{8'd106,8'd99} : s = 205;
	{8'd106,8'd100} : s = 206;
	{8'd106,8'd101} : s = 207;
	{8'd106,8'd102} : s = 208;
	{8'd106,8'd103} : s = 209;
	{8'd106,8'd104} : s = 210;
	{8'd106,8'd105} : s = 211;
	{8'd106,8'd106} : s = 212;
	{8'd106,8'd107} : s = 213;
	{8'd106,8'd108} : s = 214;
	{8'd106,8'd109} : s = 215;
	{8'd106,8'd110} : s = 216;
	{8'd106,8'd111} : s = 217;
	{8'd106,8'd112} : s = 218;
	{8'd106,8'd113} : s = 219;
	{8'd106,8'd114} : s = 220;
	{8'd106,8'd115} : s = 221;
	{8'd106,8'd116} : s = 222;
	{8'd106,8'd117} : s = 223;
	{8'd106,8'd118} : s = 224;
	{8'd106,8'd119} : s = 225;
	{8'd106,8'd120} : s = 226;
	{8'd106,8'd121} : s = 227;
	{8'd106,8'd122} : s = 228;
	{8'd106,8'd123} : s = 229;
	{8'd106,8'd124} : s = 230;
	{8'd106,8'd125} : s = 231;
	{8'd106,8'd126} : s = 232;
	{8'd106,8'd127} : s = 233;
	{8'd106,8'd128} : s = 234;
	{8'd106,8'd129} : s = 235;
	{8'd106,8'd130} : s = 236;
	{8'd106,8'd131} : s = 237;
	{8'd106,8'd132} : s = 238;
	{8'd106,8'd133} : s = 239;
	{8'd106,8'd134} : s = 240;
	{8'd106,8'd135} : s = 241;
	{8'd106,8'd136} : s = 242;
	{8'd106,8'd137} : s = 243;
	{8'd106,8'd138} : s = 244;
	{8'd106,8'd139} : s = 245;
	{8'd106,8'd140} : s = 246;
	{8'd106,8'd141} : s = 247;
	{8'd106,8'd142} : s = 248;
	{8'd106,8'd143} : s = 249;
	{8'd106,8'd144} : s = 250;
	{8'd106,8'd145} : s = 251;
	{8'd106,8'd146} : s = 252;
	{8'd106,8'd147} : s = 253;
	{8'd106,8'd148} : s = 254;
	{8'd106,8'd149} : s = 255;
	{8'd106,8'd150} : s = 256;
	{8'd106,8'd151} : s = 257;
	{8'd106,8'd152} : s = 258;
	{8'd106,8'd153} : s = 259;
	{8'd106,8'd154} : s = 260;
	{8'd106,8'd155} : s = 261;
	{8'd106,8'd156} : s = 262;
	{8'd106,8'd157} : s = 263;
	{8'd106,8'd158} : s = 264;
	{8'd106,8'd159} : s = 265;
	{8'd106,8'd160} : s = 266;
	{8'd106,8'd161} : s = 267;
	{8'd106,8'd162} : s = 268;
	{8'd106,8'd163} : s = 269;
	{8'd106,8'd164} : s = 270;
	{8'd106,8'd165} : s = 271;
	{8'd106,8'd166} : s = 272;
	{8'd106,8'd167} : s = 273;
	{8'd106,8'd168} : s = 274;
	{8'd106,8'd169} : s = 275;
	{8'd106,8'd170} : s = 276;
	{8'd106,8'd171} : s = 277;
	{8'd106,8'd172} : s = 278;
	{8'd106,8'd173} : s = 279;
	{8'd106,8'd174} : s = 280;
	{8'd106,8'd175} : s = 281;
	{8'd106,8'd176} : s = 282;
	{8'd106,8'd177} : s = 283;
	{8'd106,8'd178} : s = 284;
	{8'd106,8'd179} : s = 285;
	{8'd106,8'd180} : s = 286;
	{8'd106,8'd181} : s = 287;
	{8'd106,8'd182} : s = 288;
	{8'd106,8'd183} : s = 289;
	{8'd106,8'd184} : s = 290;
	{8'd106,8'd185} : s = 291;
	{8'd106,8'd186} : s = 292;
	{8'd106,8'd187} : s = 293;
	{8'd106,8'd188} : s = 294;
	{8'd106,8'd189} : s = 295;
	{8'd106,8'd190} : s = 296;
	{8'd106,8'd191} : s = 297;
	{8'd106,8'd192} : s = 298;
	{8'd106,8'd193} : s = 299;
	{8'd106,8'd194} : s = 300;
	{8'd106,8'd195} : s = 301;
	{8'd106,8'd196} : s = 302;
	{8'd106,8'd197} : s = 303;
	{8'd106,8'd198} : s = 304;
	{8'd106,8'd199} : s = 305;
	{8'd106,8'd200} : s = 306;
	{8'd106,8'd201} : s = 307;
	{8'd106,8'd202} : s = 308;
	{8'd106,8'd203} : s = 309;
	{8'd106,8'd204} : s = 310;
	{8'd106,8'd205} : s = 311;
	{8'd106,8'd206} : s = 312;
	{8'd106,8'd207} : s = 313;
	{8'd106,8'd208} : s = 314;
	{8'd106,8'd209} : s = 315;
	{8'd106,8'd210} : s = 316;
	{8'd106,8'd211} : s = 317;
	{8'd106,8'd212} : s = 318;
	{8'd106,8'd213} : s = 319;
	{8'd106,8'd214} : s = 320;
	{8'd106,8'd215} : s = 321;
	{8'd106,8'd216} : s = 322;
	{8'd106,8'd217} : s = 323;
	{8'd106,8'd218} : s = 324;
	{8'd106,8'd219} : s = 325;
	{8'd106,8'd220} : s = 326;
	{8'd106,8'd221} : s = 327;
	{8'd106,8'd222} : s = 328;
	{8'd106,8'd223} : s = 329;
	{8'd106,8'd224} : s = 330;
	{8'd106,8'd225} : s = 331;
	{8'd106,8'd226} : s = 332;
	{8'd106,8'd227} : s = 333;
	{8'd106,8'd228} : s = 334;
	{8'd106,8'd229} : s = 335;
	{8'd106,8'd230} : s = 336;
	{8'd106,8'd231} : s = 337;
	{8'd106,8'd232} : s = 338;
	{8'd106,8'd233} : s = 339;
	{8'd106,8'd234} : s = 340;
	{8'd106,8'd235} : s = 341;
	{8'd106,8'd236} : s = 342;
	{8'd106,8'd237} : s = 343;
	{8'd106,8'd238} : s = 344;
	{8'd106,8'd239} : s = 345;
	{8'd106,8'd240} : s = 346;
	{8'd106,8'd241} : s = 347;
	{8'd106,8'd242} : s = 348;
	{8'd106,8'd243} : s = 349;
	{8'd106,8'd244} : s = 350;
	{8'd106,8'd245} : s = 351;
	{8'd106,8'd246} : s = 352;
	{8'd106,8'd247} : s = 353;
	{8'd106,8'd248} : s = 354;
	{8'd106,8'd249} : s = 355;
	{8'd106,8'd250} : s = 356;
	{8'd106,8'd251} : s = 357;
	{8'd106,8'd252} : s = 358;
	{8'd106,8'd253} : s = 359;
	{8'd106,8'd254} : s = 360;
	{8'd106,8'd255} : s = 361;
	{8'd107,8'd0} : s = 107;
	{8'd107,8'd1} : s = 108;
	{8'd107,8'd2} : s = 109;
	{8'd107,8'd3} : s = 110;
	{8'd107,8'd4} : s = 111;
	{8'd107,8'd5} : s = 112;
	{8'd107,8'd6} : s = 113;
	{8'd107,8'd7} : s = 114;
	{8'd107,8'd8} : s = 115;
	{8'd107,8'd9} : s = 116;
	{8'd107,8'd10} : s = 117;
	{8'd107,8'd11} : s = 118;
	{8'd107,8'd12} : s = 119;
	{8'd107,8'd13} : s = 120;
	{8'd107,8'd14} : s = 121;
	{8'd107,8'd15} : s = 122;
	{8'd107,8'd16} : s = 123;
	{8'd107,8'd17} : s = 124;
	{8'd107,8'd18} : s = 125;
	{8'd107,8'd19} : s = 126;
	{8'd107,8'd20} : s = 127;
	{8'd107,8'd21} : s = 128;
	{8'd107,8'd22} : s = 129;
	{8'd107,8'd23} : s = 130;
	{8'd107,8'd24} : s = 131;
	{8'd107,8'd25} : s = 132;
	{8'd107,8'd26} : s = 133;
	{8'd107,8'd27} : s = 134;
	{8'd107,8'd28} : s = 135;
	{8'd107,8'd29} : s = 136;
	{8'd107,8'd30} : s = 137;
	{8'd107,8'd31} : s = 138;
	{8'd107,8'd32} : s = 139;
	{8'd107,8'd33} : s = 140;
	{8'd107,8'd34} : s = 141;
	{8'd107,8'd35} : s = 142;
	{8'd107,8'd36} : s = 143;
	{8'd107,8'd37} : s = 144;
	{8'd107,8'd38} : s = 145;
	{8'd107,8'd39} : s = 146;
	{8'd107,8'd40} : s = 147;
	{8'd107,8'd41} : s = 148;
	{8'd107,8'd42} : s = 149;
	{8'd107,8'd43} : s = 150;
	{8'd107,8'd44} : s = 151;
	{8'd107,8'd45} : s = 152;
	{8'd107,8'd46} : s = 153;
	{8'd107,8'd47} : s = 154;
	{8'd107,8'd48} : s = 155;
	{8'd107,8'd49} : s = 156;
	{8'd107,8'd50} : s = 157;
	{8'd107,8'd51} : s = 158;
	{8'd107,8'd52} : s = 159;
	{8'd107,8'd53} : s = 160;
	{8'd107,8'd54} : s = 161;
	{8'd107,8'd55} : s = 162;
	{8'd107,8'd56} : s = 163;
	{8'd107,8'd57} : s = 164;
	{8'd107,8'd58} : s = 165;
	{8'd107,8'd59} : s = 166;
	{8'd107,8'd60} : s = 167;
	{8'd107,8'd61} : s = 168;
	{8'd107,8'd62} : s = 169;
	{8'd107,8'd63} : s = 170;
	{8'd107,8'd64} : s = 171;
	{8'd107,8'd65} : s = 172;
	{8'd107,8'd66} : s = 173;
	{8'd107,8'd67} : s = 174;
	{8'd107,8'd68} : s = 175;
	{8'd107,8'd69} : s = 176;
	{8'd107,8'd70} : s = 177;
	{8'd107,8'd71} : s = 178;
	{8'd107,8'd72} : s = 179;
	{8'd107,8'd73} : s = 180;
	{8'd107,8'd74} : s = 181;
	{8'd107,8'd75} : s = 182;
	{8'd107,8'd76} : s = 183;
	{8'd107,8'd77} : s = 184;
	{8'd107,8'd78} : s = 185;
	{8'd107,8'd79} : s = 186;
	{8'd107,8'd80} : s = 187;
	{8'd107,8'd81} : s = 188;
	{8'd107,8'd82} : s = 189;
	{8'd107,8'd83} : s = 190;
	{8'd107,8'd84} : s = 191;
	{8'd107,8'd85} : s = 192;
	{8'd107,8'd86} : s = 193;
	{8'd107,8'd87} : s = 194;
	{8'd107,8'd88} : s = 195;
	{8'd107,8'd89} : s = 196;
	{8'd107,8'd90} : s = 197;
	{8'd107,8'd91} : s = 198;
	{8'd107,8'd92} : s = 199;
	{8'd107,8'd93} : s = 200;
	{8'd107,8'd94} : s = 201;
	{8'd107,8'd95} : s = 202;
	{8'd107,8'd96} : s = 203;
	{8'd107,8'd97} : s = 204;
	{8'd107,8'd98} : s = 205;
	{8'd107,8'd99} : s = 206;
	{8'd107,8'd100} : s = 207;
	{8'd107,8'd101} : s = 208;
	{8'd107,8'd102} : s = 209;
	{8'd107,8'd103} : s = 210;
	{8'd107,8'd104} : s = 211;
	{8'd107,8'd105} : s = 212;
	{8'd107,8'd106} : s = 213;
	{8'd107,8'd107} : s = 214;
	{8'd107,8'd108} : s = 215;
	{8'd107,8'd109} : s = 216;
	{8'd107,8'd110} : s = 217;
	{8'd107,8'd111} : s = 218;
	{8'd107,8'd112} : s = 219;
	{8'd107,8'd113} : s = 220;
	{8'd107,8'd114} : s = 221;
	{8'd107,8'd115} : s = 222;
	{8'd107,8'd116} : s = 223;
	{8'd107,8'd117} : s = 224;
	{8'd107,8'd118} : s = 225;
	{8'd107,8'd119} : s = 226;
	{8'd107,8'd120} : s = 227;
	{8'd107,8'd121} : s = 228;
	{8'd107,8'd122} : s = 229;
	{8'd107,8'd123} : s = 230;
	{8'd107,8'd124} : s = 231;
	{8'd107,8'd125} : s = 232;
	{8'd107,8'd126} : s = 233;
	{8'd107,8'd127} : s = 234;
	{8'd107,8'd128} : s = 235;
	{8'd107,8'd129} : s = 236;
	{8'd107,8'd130} : s = 237;
	{8'd107,8'd131} : s = 238;
	{8'd107,8'd132} : s = 239;
	{8'd107,8'd133} : s = 240;
	{8'd107,8'd134} : s = 241;
	{8'd107,8'd135} : s = 242;
	{8'd107,8'd136} : s = 243;
	{8'd107,8'd137} : s = 244;
	{8'd107,8'd138} : s = 245;
	{8'd107,8'd139} : s = 246;
	{8'd107,8'd140} : s = 247;
	{8'd107,8'd141} : s = 248;
	{8'd107,8'd142} : s = 249;
	{8'd107,8'd143} : s = 250;
	{8'd107,8'd144} : s = 251;
	{8'd107,8'd145} : s = 252;
	{8'd107,8'd146} : s = 253;
	{8'd107,8'd147} : s = 254;
	{8'd107,8'd148} : s = 255;
	{8'd107,8'd149} : s = 256;
	{8'd107,8'd150} : s = 257;
	{8'd107,8'd151} : s = 258;
	{8'd107,8'd152} : s = 259;
	{8'd107,8'd153} : s = 260;
	{8'd107,8'd154} : s = 261;
	{8'd107,8'd155} : s = 262;
	{8'd107,8'd156} : s = 263;
	{8'd107,8'd157} : s = 264;
	{8'd107,8'd158} : s = 265;
	{8'd107,8'd159} : s = 266;
	{8'd107,8'd160} : s = 267;
	{8'd107,8'd161} : s = 268;
	{8'd107,8'd162} : s = 269;
	{8'd107,8'd163} : s = 270;
	{8'd107,8'd164} : s = 271;
	{8'd107,8'd165} : s = 272;
	{8'd107,8'd166} : s = 273;
	{8'd107,8'd167} : s = 274;
	{8'd107,8'd168} : s = 275;
	{8'd107,8'd169} : s = 276;
	{8'd107,8'd170} : s = 277;
	{8'd107,8'd171} : s = 278;
	{8'd107,8'd172} : s = 279;
	{8'd107,8'd173} : s = 280;
	{8'd107,8'd174} : s = 281;
	{8'd107,8'd175} : s = 282;
	{8'd107,8'd176} : s = 283;
	{8'd107,8'd177} : s = 284;
	{8'd107,8'd178} : s = 285;
	{8'd107,8'd179} : s = 286;
	{8'd107,8'd180} : s = 287;
	{8'd107,8'd181} : s = 288;
	{8'd107,8'd182} : s = 289;
	{8'd107,8'd183} : s = 290;
	{8'd107,8'd184} : s = 291;
	{8'd107,8'd185} : s = 292;
	{8'd107,8'd186} : s = 293;
	{8'd107,8'd187} : s = 294;
	{8'd107,8'd188} : s = 295;
	{8'd107,8'd189} : s = 296;
	{8'd107,8'd190} : s = 297;
	{8'd107,8'd191} : s = 298;
	{8'd107,8'd192} : s = 299;
	{8'd107,8'd193} : s = 300;
	{8'd107,8'd194} : s = 301;
	{8'd107,8'd195} : s = 302;
	{8'd107,8'd196} : s = 303;
	{8'd107,8'd197} : s = 304;
	{8'd107,8'd198} : s = 305;
	{8'd107,8'd199} : s = 306;
	{8'd107,8'd200} : s = 307;
	{8'd107,8'd201} : s = 308;
	{8'd107,8'd202} : s = 309;
	{8'd107,8'd203} : s = 310;
	{8'd107,8'd204} : s = 311;
	{8'd107,8'd205} : s = 312;
	{8'd107,8'd206} : s = 313;
	{8'd107,8'd207} : s = 314;
	{8'd107,8'd208} : s = 315;
	{8'd107,8'd209} : s = 316;
	{8'd107,8'd210} : s = 317;
	{8'd107,8'd211} : s = 318;
	{8'd107,8'd212} : s = 319;
	{8'd107,8'd213} : s = 320;
	{8'd107,8'd214} : s = 321;
	{8'd107,8'd215} : s = 322;
	{8'd107,8'd216} : s = 323;
	{8'd107,8'd217} : s = 324;
	{8'd107,8'd218} : s = 325;
	{8'd107,8'd219} : s = 326;
	{8'd107,8'd220} : s = 327;
	{8'd107,8'd221} : s = 328;
	{8'd107,8'd222} : s = 329;
	{8'd107,8'd223} : s = 330;
	{8'd107,8'd224} : s = 331;
	{8'd107,8'd225} : s = 332;
	{8'd107,8'd226} : s = 333;
	{8'd107,8'd227} : s = 334;
	{8'd107,8'd228} : s = 335;
	{8'd107,8'd229} : s = 336;
	{8'd107,8'd230} : s = 337;
	{8'd107,8'd231} : s = 338;
	{8'd107,8'd232} : s = 339;
	{8'd107,8'd233} : s = 340;
	{8'd107,8'd234} : s = 341;
	{8'd107,8'd235} : s = 342;
	{8'd107,8'd236} : s = 343;
	{8'd107,8'd237} : s = 344;
	{8'd107,8'd238} : s = 345;
	{8'd107,8'd239} : s = 346;
	{8'd107,8'd240} : s = 347;
	{8'd107,8'd241} : s = 348;
	{8'd107,8'd242} : s = 349;
	{8'd107,8'd243} : s = 350;
	{8'd107,8'd244} : s = 351;
	{8'd107,8'd245} : s = 352;
	{8'd107,8'd246} : s = 353;
	{8'd107,8'd247} : s = 354;
	{8'd107,8'd248} : s = 355;
	{8'd107,8'd249} : s = 356;
	{8'd107,8'd250} : s = 357;
	{8'd107,8'd251} : s = 358;
	{8'd107,8'd252} : s = 359;
	{8'd107,8'd253} : s = 360;
	{8'd107,8'd254} : s = 361;
	{8'd107,8'd255} : s = 362;
	{8'd108,8'd0} : s = 108;
	{8'd108,8'd1} : s = 109;
	{8'd108,8'd2} : s = 110;
	{8'd108,8'd3} : s = 111;
	{8'd108,8'd4} : s = 112;
	{8'd108,8'd5} : s = 113;
	{8'd108,8'd6} : s = 114;
	{8'd108,8'd7} : s = 115;
	{8'd108,8'd8} : s = 116;
	{8'd108,8'd9} : s = 117;
	{8'd108,8'd10} : s = 118;
	{8'd108,8'd11} : s = 119;
	{8'd108,8'd12} : s = 120;
	{8'd108,8'd13} : s = 121;
	{8'd108,8'd14} : s = 122;
	{8'd108,8'd15} : s = 123;
	{8'd108,8'd16} : s = 124;
	{8'd108,8'd17} : s = 125;
	{8'd108,8'd18} : s = 126;
	{8'd108,8'd19} : s = 127;
	{8'd108,8'd20} : s = 128;
	{8'd108,8'd21} : s = 129;
	{8'd108,8'd22} : s = 130;
	{8'd108,8'd23} : s = 131;
	{8'd108,8'd24} : s = 132;
	{8'd108,8'd25} : s = 133;
	{8'd108,8'd26} : s = 134;
	{8'd108,8'd27} : s = 135;
	{8'd108,8'd28} : s = 136;
	{8'd108,8'd29} : s = 137;
	{8'd108,8'd30} : s = 138;
	{8'd108,8'd31} : s = 139;
	{8'd108,8'd32} : s = 140;
	{8'd108,8'd33} : s = 141;
	{8'd108,8'd34} : s = 142;
	{8'd108,8'd35} : s = 143;
	{8'd108,8'd36} : s = 144;
	{8'd108,8'd37} : s = 145;
	{8'd108,8'd38} : s = 146;
	{8'd108,8'd39} : s = 147;
	{8'd108,8'd40} : s = 148;
	{8'd108,8'd41} : s = 149;
	{8'd108,8'd42} : s = 150;
	{8'd108,8'd43} : s = 151;
	{8'd108,8'd44} : s = 152;
	{8'd108,8'd45} : s = 153;
	{8'd108,8'd46} : s = 154;
	{8'd108,8'd47} : s = 155;
	{8'd108,8'd48} : s = 156;
	{8'd108,8'd49} : s = 157;
	{8'd108,8'd50} : s = 158;
	{8'd108,8'd51} : s = 159;
	{8'd108,8'd52} : s = 160;
	{8'd108,8'd53} : s = 161;
	{8'd108,8'd54} : s = 162;
	{8'd108,8'd55} : s = 163;
	{8'd108,8'd56} : s = 164;
	{8'd108,8'd57} : s = 165;
	{8'd108,8'd58} : s = 166;
	{8'd108,8'd59} : s = 167;
	{8'd108,8'd60} : s = 168;
	{8'd108,8'd61} : s = 169;
	{8'd108,8'd62} : s = 170;
	{8'd108,8'd63} : s = 171;
	{8'd108,8'd64} : s = 172;
	{8'd108,8'd65} : s = 173;
	{8'd108,8'd66} : s = 174;
	{8'd108,8'd67} : s = 175;
	{8'd108,8'd68} : s = 176;
	{8'd108,8'd69} : s = 177;
	{8'd108,8'd70} : s = 178;
	{8'd108,8'd71} : s = 179;
	{8'd108,8'd72} : s = 180;
	{8'd108,8'd73} : s = 181;
	{8'd108,8'd74} : s = 182;
	{8'd108,8'd75} : s = 183;
	{8'd108,8'd76} : s = 184;
	{8'd108,8'd77} : s = 185;
	{8'd108,8'd78} : s = 186;
	{8'd108,8'd79} : s = 187;
	{8'd108,8'd80} : s = 188;
	{8'd108,8'd81} : s = 189;
	{8'd108,8'd82} : s = 190;
	{8'd108,8'd83} : s = 191;
	{8'd108,8'd84} : s = 192;
	{8'd108,8'd85} : s = 193;
	{8'd108,8'd86} : s = 194;
	{8'd108,8'd87} : s = 195;
	{8'd108,8'd88} : s = 196;
	{8'd108,8'd89} : s = 197;
	{8'd108,8'd90} : s = 198;
	{8'd108,8'd91} : s = 199;
	{8'd108,8'd92} : s = 200;
	{8'd108,8'd93} : s = 201;
	{8'd108,8'd94} : s = 202;
	{8'd108,8'd95} : s = 203;
	{8'd108,8'd96} : s = 204;
	{8'd108,8'd97} : s = 205;
	{8'd108,8'd98} : s = 206;
	{8'd108,8'd99} : s = 207;
	{8'd108,8'd100} : s = 208;
	{8'd108,8'd101} : s = 209;
	{8'd108,8'd102} : s = 210;
	{8'd108,8'd103} : s = 211;
	{8'd108,8'd104} : s = 212;
	{8'd108,8'd105} : s = 213;
	{8'd108,8'd106} : s = 214;
	{8'd108,8'd107} : s = 215;
	{8'd108,8'd108} : s = 216;
	{8'd108,8'd109} : s = 217;
	{8'd108,8'd110} : s = 218;
	{8'd108,8'd111} : s = 219;
	{8'd108,8'd112} : s = 220;
	{8'd108,8'd113} : s = 221;
	{8'd108,8'd114} : s = 222;
	{8'd108,8'd115} : s = 223;
	{8'd108,8'd116} : s = 224;
	{8'd108,8'd117} : s = 225;
	{8'd108,8'd118} : s = 226;
	{8'd108,8'd119} : s = 227;
	{8'd108,8'd120} : s = 228;
	{8'd108,8'd121} : s = 229;
	{8'd108,8'd122} : s = 230;
	{8'd108,8'd123} : s = 231;
	{8'd108,8'd124} : s = 232;
	{8'd108,8'd125} : s = 233;
	{8'd108,8'd126} : s = 234;
	{8'd108,8'd127} : s = 235;
	{8'd108,8'd128} : s = 236;
	{8'd108,8'd129} : s = 237;
	{8'd108,8'd130} : s = 238;
	{8'd108,8'd131} : s = 239;
	{8'd108,8'd132} : s = 240;
	{8'd108,8'd133} : s = 241;
	{8'd108,8'd134} : s = 242;
	{8'd108,8'd135} : s = 243;
	{8'd108,8'd136} : s = 244;
	{8'd108,8'd137} : s = 245;
	{8'd108,8'd138} : s = 246;
	{8'd108,8'd139} : s = 247;
	{8'd108,8'd140} : s = 248;
	{8'd108,8'd141} : s = 249;
	{8'd108,8'd142} : s = 250;
	{8'd108,8'd143} : s = 251;
	{8'd108,8'd144} : s = 252;
	{8'd108,8'd145} : s = 253;
	{8'd108,8'd146} : s = 254;
	{8'd108,8'd147} : s = 255;
	{8'd108,8'd148} : s = 256;
	{8'd108,8'd149} : s = 257;
	{8'd108,8'd150} : s = 258;
	{8'd108,8'd151} : s = 259;
	{8'd108,8'd152} : s = 260;
	{8'd108,8'd153} : s = 261;
	{8'd108,8'd154} : s = 262;
	{8'd108,8'd155} : s = 263;
	{8'd108,8'd156} : s = 264;
	{8'd108,8'd157} : s = 265;
	{8'd108,8'd158} : s = 266;
	{8'd108,8'd159} : s = 267;
	{8'd108,8'd160} : s = 268;
	{8'd108,8'd161} : s = 269;
	{8'd108,8'd162} : s = 270;
	{8'd108,8'd163} : s = 271;
	{8'd108,8'd164} : s = 272;
	{8'd108,8'd165} : s = 273;
	{8'd108,8'd166} : s = 274;
	{8'd108,8'd167} : s = 275;
	{8'd108,8'd168} : s = 276;
	{8'd108,8'd169} : s = 277;
	{8'd108,8'd170} : s = 278;
	{8'd108,8'd171} : s = 279;
	{8'd108,8'd172} : s = 280;
	{8'd108,8'd173} : s = 281;
	{8'd108,8'd174} : s = 282;
	{8'd108,8'd175} : s = 283;
	{8'd108,8'd176} : s = 284;
	{8'd108,8'd177} : s = 285;
	{8'd108,8'd178} : s = 286;
	{8'd108,8'd179} : s = 287;
	{8'd108,8'd180} : s = 288;
	{8'd108,8'd181} : s = 289;
	{8'd108,8'd182} : s = 290;
	{8'd108,8'd183} : s = 291;
	{8'd108,8'd184} : s = 292;
	{8'd108,8'd185} : s = 293;
	{8'd108,8'd186} : s = 294;
	{8'd108,8'd187} : s = 295;
	{8'd108,8'd188} : s = 296;
	{8'd108,8'd189} : s = 297;
	{8'd108,8'd190} : s = 298;
	{8'd108,8'd191} : s = 299;
	{8'd108,8'd192} : s = 300;
	{8'd108,8'd193} : s = 301;
	{8'd108,8'd194} : s = 302;
	{8'd108,8'd195} : s = 303;
	{8'd108,8'd196} : s = 304;
	{8'd108,8'd197} : s = 305;
	{8'd108,8'd198} : s = 306;
	{8'd108,8'd199} : s = 307;
	{8'd108,8'd200} : s = 308;
	{8'd108,8'd201} : s = 309;
	{8'd108,8'd202} : s = 310;
	{8'd108,8'd203} : s = 311;
	{8'd108,8'd204} : s = 312;
	{8'd108,8'd205} : s = 313;
	{8'd108,8'd206} : s = 314;
	{8'd108,8'd207} : s = 315;
	{8'd108,8'd208} : s = 316;
	{8'd108,8'd209} : s = 317;
	{8'd108,8'd210} : s = 318;
	{8'd108,8'd211} : s = 319;
	{8'd108,8'd212} : s = 320;
	{8'd108,8'd213} : s = 321;
	{8'd108,8'd214} : s = 322;
	{8'd108,8'd215} : s = 323;
	{8'd108,8'd216} : s = 324;
	{8'd108,8'd217} : s = 325;
	{8'd108,8'd218} : s = 326;
	{8'd108,8'd219} : s = 327;
	{8'd108,8'd220} : s = 328;
	{8'd108,8'd221} : s = 329;
	{8'd108,8'd222} : s = 330;
	{8'd108,8'd223} : s = 331;
	{8'd108,8'd224} : s = 332;
	{8'd108,8'd225} : s = 333;
	{8'd108,8'd226} : s = 334;
	{8'd108,8'd227} : s = 335;
	{8'd108,8'd228} : s = 336;
	{8'd108,8'd229} : s = 337;
	{8'd108,8'd230} : s = 338;
	{8'd108,8'd231} : s = 339;
	{8'd108,8'd232} : s = 340;
	{8'd108,8'd233} : s = 341;
	{8'd108,8'd234} : s = 342;
	{8'd108,8'd235} : s = 343;
	{8'd108,8'd236} : s = 344;
	{8'd108,8'd237} : s = 345;
	{8'd108,8'd238} : s = 346;
	{8'd108,8'd239} : s = 347;
	{8'd108,8'd240} : s = 348;
	{8'd108,8'd241} : s = 349;
	{8'd108,8'd242} : s = 350;
	{8'd108,8'd243} : s = 351;
	{8'd108,8'd244} : s = 352;
	{8'd108,8'd245} : s = 353;
	{8'd108,8'd246} : s = 354;
	{8'd108,8'd247} : s = 355;
	{8'd108,8'd248} : s = 356;
	{8'd108,8'd249} : s = 357;
	{8'd108,8'd250} : s = 358;
	{8'd108,8'd251} : s = 359;
	{8'd108,8'd252} : s = 360;
	{8'd108,8'd253} : s = 361;
	{8'd108,8'd254} : s = 362;
	{8'd108,8'd255} : s = 363;
	{8'd109,8'd0} : s = 109;
	{8'd109,8'd1} : s = 110;
	{8'd109,8'd2} : s = 111;
	{8'd109,8'd3} : s = 112;
	{8'd109,8'd4} : s = 113;
	{8'd109,8'd5} : s = 114;
	{8'd109,8'd6} : s = 115;
	{8'd109,8'd7} : s = 116;
	{8'd109,8'd8} : s = 117;
	{8'd109,8'd9} : s = 118;
	{8'd109,8'd10} : s = 119;
	{8'd109,8'd11} : s = 120;
	{8'd109,8'd12} : s = 121;
	{8'd109,8'd13} : s = 122;
	{8'd109,8'd14} : s = 123;
	{8'd109,8'd15} : s = 124;
	{8'd109,8'd16} : s = 125;
	{8'd109,8'd17} : s = 126;
	{8'd109,8'd18} : s = 127;
	{8'd109,8'd19} : s = 128;
	{8'd109,8'd20} : s = 129;
	{8'd109,8'd21} : s = 130;
	{8'd109,8'd22} : s = 131;
	{8'd109,8'd23} : s = 132;
	{8'd109,8'd24} : s = 133;
	{8'd109,8'd25} : s = 134;
	{8'd109,8'd26} : s = 135;
	{8'd109,8'd27} : s = 136;
	{8'd109,8'd28} : s = 137;
	{8'd109,8'd29} : s = 138;
	{8'd109,8'd30} : s = 139;
	{8'd109,8'd31} : s = 140;
	{8'd109,8'd32} : s = 141;
	{8'd109,8'd33} : s = 142;
	{8'd109,8'd34} : s = 143;
	{8'd109,8'd35} : s = 144;
	{8'd109,8'd36} : s = 145;
	{8'd109,8'd37} : s = 146;
	{8'd109,8'd38} : s = 147;
	{8'd109,8'd39} : s = 148;
	{8'd109,8'd40} : s = 149;
	{8'd109,8'd41} : s = 150;
	{8'd109,8'd42} : s = 151;
	{8'd109,8'd43} : s = 152;
	{8'd109,8'd44} : s = 153;
	{8'd109,8'd45} : s = 154;
	{8'd109,8'd46} : s = 155;
	{8'd109,8'd47} : s = 156;
	{8'd109,8'd48} : s = 157;
	{8'd109,8'd49} : s = 158;
	{8'd109,8'd50} : s = 159;
	{8'd109,8'd51} : s = 160;
	{8'd109,8'd52} : s = 161;
	{8'd109,8'd53} : s = 162;
	{8'd109,8'd54} : s = 163;
	{8'd109,8'd55} : s = 164;
	{8'd109,8'd56} : s = 165;
	{8'd109,8'd57} : s = 166;
	{8'd109,8'd58} : s = 167;
	{8'd109,8'd59} : s = 168;
	{8'd109,8'd60} : s = 169;
	{8'd109,8'd61} : s = 170;
	{8'd109,8'd62} : s = 171;
	{8'd109,8'd63} : s = 172;
	{8'd109,8'd64} : s = 173;
	{8'd109,8'd65} : s = 174;
	{8'd109,8'd66} : s = 175;
	{8'd109,8'd67} : s = 176;
	{8'd109,8'd68} : s = 177;
	{8'd109,8'd69} : s = 178;
	{8'd109,8'd70} : s = 179;
	{8'd109,8'd71} : s = 180;
	{8'd109,8'd72} : s = 181;
	{8'd109,8'd73} : s = 182;
	{8'd109,8'd74} : s = 183;
	{8'd109,8'd75} : s = 184;
	{8'd109,8'd76} : s = 185;
	{8'd109,8'd77} : s = 186;
	{8'd109,8'd78} : s = 187;
	{8'd109,8'd79} : s = 188;
	{8'd109,8'd80} : s = 189;
	{8'd109,8'd81} : s = 190;
	{8'd109,8'd82} : s = 191;
	{8'd109,8'd83} : s = 192;
	{8'd109,8'd84} : s = 193;
	{8'd109,8'd85} : s = 194;
	{8'd109,8'd86} : s = 195;
	{8'd109,8'd87} : s = 196;
	{8'd109,8'd88} : s = 197;
	{8'd109,8'd89} : s = 198;
	{8'd109,8'd90} : s = 199;
	{8'd109,8'd91} : s = 200;
	{8'd109,8'd92} : s = 201;
	{8'd109,8'd93} : s = 202;
	{8'd109,8'd94} : s = 203;
	{8'd109,8'd95} : s = 204;
	{8'd109,8'd96} : s = 205;
	{8'd109,8'd97} : s = 206;
	{8'd109,8'd98} : s = 207;
	{8'd109,8'd99} : s = 208;
	{8'd109,8'd100} : s = 209;
	{8'd109,8'd101} : s = 210;
	{8'd109,8'd102} : s = 211;
	{8'd109,8'd103} : s = 212;
	{8'd109,8'd104} : s = 213;
	{8'd109,8'd105} : s = 214;
	{8'd109,8'd106} : s = 215;
	{8'd109,8'd107} : s = 216;
	{8'd109,8'd108} : s = 217;
	{8'd109,8'd109} : s = 218;
	{8'd109,8'd110} : s = 219;
	{8'd109,8'd111} : s = 220;
	{8'd109,8'd112} : s = 221;
	{8'd109,8'd113} : s = 222;
	{8'd109,8'd114} : s = 223;
	{8'd109,8'd115} : s = 224;
	{8'd109,8'd116} : s = 225;
	{8'd109,8'd117} : s = 226;
	{8'd109,8'd118} : s = 227;
	{8'd109,8'd119} : s = 228;
	{8'd109,8'd120} : s = 229;
	{8'd109,8'd121} : s = 230;
	{8'd109,8'd122} : s = 231;
	{8'd109,8'd123} : s = 232;
	{8'd109,8'd124} : s = 233;
	{8'd109,8'd125} : s = 234;
	{8'd109,8'd126} : s = 235;
	{8'd109,8'd127} : s = 236;
	{8'd109,8'd128} : s = 237;
	{8'd109,8'd129} : s = 238;
	{8'd109,8'd130} : s = 239;
	{8'd109,8'd131} : s = 240;
	{8'd109,8'd132} : s = 241;
	{8'd109,8'd133} : s = 242;
	{8'd109,8'd134} : s = 243;
	{8'd109,8'd135} : s = 244;
	{8'd109,8'd136} : s = 245;
	{8'd109,8'd137} : s = 246;
	{8'd109,8'd138} : s = 247;
	{8'd109,8'd139} : s = 248;
	{8'd109,8'd140} : s = 249;
	{8'd109,8'd141} : s = 250;
	{8'd109,8'd142} : s = 251;
	{8'd109,8'd143} : s = 252;
	{8'd109,8'd144} : s = 253;
	{8'd109,8'd145} : s = 254;
	{8'd109,8'd146} : s = 255;
	{8'd109,8'd147} : s = 256;
	{8'd109,8'd148} : s = 257;
	{8'd109,8'd149} : s = 258;
	{8'd109,8'd150} : s = 259;
	{8'd109,8'd151} : s = 260;
	{8'd109,8'd152} : s = 261;
	{8'd109,8'd153} : s = 262;
	{8'd109,8'd154} : s = 263;
	{8'd109,8'd155} : s = 264;
	{8'd109,8'd156} : s = 265;
	{8'd109,8'd157} : s = 266;
	{8'd109,8'd158} : s = 267;
	{8'd109,8'd159} : s = 268;
	{8'd109,8'd160} : s = 269;
	{8'd109,8'd161} : s = 270;
	{8'd109,8'd162} : s = 271;
	{8'd109,8'd163} : s = 272;
	{8'd109,8'd164} : s = 273;
	{8'd109,8'd165} : s = 274;
	{8'd109,8'd166} : s = 275;
	{8'd109,8'd167} : s = 276;
	{8'd109,8'd168} : s = 277;
	{8'd109,8'd169} : s = 278;
	{8'd109,8'd170} : s = 279;
	{8'd109,8'd171} : s = 280;
	{8'd109,8'd172} : s = 281;
	{8'd109,8'd173} : s = 282;
	{8'd109,8'd174} : s = 283;
	{8'd109,8'd175} : s = 284;
	{8'd109,8'd176} : s = 285;
	{8'd109,8'd177} : s = 286;
	{8'd109,8'd178} : s = 287;
	{8'd109,8'd179} : s = 288;
	{8'd109,8'd180} : s = 289;
	{8'd109,8'd181} : s = 290;
	{8'd109,8'd182} : s = 291;
	{8'd109,8'd183} : s = 292;
	{8'd109,8'd184} : s = 293;
	{8'd109,8'd185} : s = 294;
	{8'd109,8'd186} : s = 295;
	{8'd109,8'd187} : s = 296;
	{8'd109,8'd188} : s = 297;
	{8'd109,8'd189} : s = 298;
	{8'd109,8'd190} : s = 299;
	{8'd109,8'd191} : s = 300;
	{8'd109,8'd192} : s = 301;
	{8'd109,8'd193} : s = 302;
	{8'd109,8'd194} : s = 303;
	{8'd109,8'd195} : s = 304;
	{8'd109,8'd196} : s = 305;
	{8'd109,8'd197} : s = 306;
	{8'd109,8'd198} : s = 307;
	{8'd109,8'd199} : s = 308;
	{8'd109,8'd200} : s = 309;
	{8'd109,8'd201} : s = 310;
	{8'd109,8'd202} : s = 311;
	{8'd109,8'd203} : s = 312;
	{8'd109,8'd204} : s = 313;
	{8'd109,8'd205} : s = 314;
	{8'd109,8'd206} : s = 315;
	{8'd109,8'd207} : s = 316;
	{8'd109,8'd208} : s = 317;
	{8'd109,8'd209} : s = 318;
	{8'd109,8'd210} : s = 319;
	{8'd109,8'd211} : s = 320;
	{8'd109,8'd212} : s = 321;
	{8'd109,8'd213} : s = 322;
	{8'd109,8'd214} : s = 323;
	{8'd109,8'd215} : s = 324;
	{8'd109,8'd216} : s = 325;
	{8'd109,8'd217} : s = 326;
	{8'd109,8'd218} : s = 327;
	{8'd109,8'd219} : s = 328;
	{8'd109,8'd220} : s = 329;
	{8'd109,8'd221} : s = 330;
	{8'd109,8'd222} : s = 331;
	{8'd109,8'd223} : s = 332;
	{8'd109,8'd224} : s = 333;
	{8'd109,8'd225} : s = 334;
	{8'd109,8'd226} : s = 335;
	{8'd109,8'd227} : s = 336;
	{8'd109,8'd228} : s = 337;
	{8'd109,8'd229} : s = 338;
	{8'd109,8'd230} : s = 339;
	{8'd109,8'd231} : s = 340;
	{8'd109,8'd232} : s = 341;
	{8'd109,8'd233} : s = 342;
	{8'd109,8'd234} : s = 343;
	{8'd109,8'd235} : s = 344;
	{8'd109,8'd236} : s = 345;
	{8'd109,8'd237} : s = 346;
	{8'd109,8'd238} : s = 347;
	{8'd109,8'd239} : s = 348;
	{8'd109,8'd240} : s = 349;
	{8'd109,8'd241} : s = 350;
	{8'd109,8'd242} : s = 351;
	{8'd109,8'd243} : s = 352;
	{8'd109,8'd244} : s = 353;
	{8'd109,8'd245} : s = 354;
	{8'd109,8'd246} : s = 355;
	{8'd109,8'd247} : s = 356;
	{8'd109,8'd248} : s = 357;
	{8'd109,8'd249} : s = 358;
	{8'd109,8'd250} : s = 359;
	{8'd109,8'd251} : s = 360;
	{8'd109,8'd252} : s = 361;
	{8'd109,8'd253} : s = 362;
	{8'd109,8'd254} : s = 363;
	{8'd109,8'd255} : s = 364;
	{8'd110,8'd0} : s = 110;
	{8'd110,8'd1} : s = 111;
	{8'd110,8'd2} : s = 112;
	{8'd110,8'd3} : s = 113;
	{8'd110,8'd4} : s = 114;
	{8'd110,8'd5} : s = 115;
	{8'd110,8'd6} : s = 116;
	{8'd110,8'd7} : s = 117;
	{8'd110,8'd8} : s = 118;
	{8'd110,8'd9} : s = 119;
	{8'd110,8'd10} : s = 120;
	{8'd110,8'd11} : s = 121;
	{8'd110,8'd12} : s = 122;
	{8'd110,8'd13} : s = 123;
	{8'd110,8'd14} : s = 124;
	{8'd110,8'd15} : s = 125;
	{8'd110,8'd16} : s = 126;
	{8'd110,8'd17} : s = 127;
	{8'd110,8'd18} : s = 128;
	{8'd110,8'd19} : s = 129;
	{8'd110,8'd20} : s = 130;
	{8'd110,8'd21} : s = 131;
	{8'd110,8'd22} : s = 132;
	{8'd110,8'd23} : s = 133;
	{8'd110,8'd24} : s = 134;
	{8'd110,8'd25} : s = 135;
	{8'd110,8'd26} : s = 136;
	{8'd110,8'd27} : s = 137;
	{8'd110,8'd28} : s = 138;
	{8'd110,8'd29} : s = 139;
	{8'd110,8'd30} : s = 140;
	{8'd110,8'd31} : s = 141;
	{8'd110,8'd32} : s = 142;
	{8'd110,8'd33} : s = 143;
	{8'd110,8'd34} : s = 144;
	{8'd110,8'd35} : s = 145;
	{8'd110,8'd36} : s = 146;
	{8'd110,8'd37} : s = 147;
	{8'd110,8'd38} : s = 148;
	{8'd110,8'd39} : s = 149;
	{8'd110,8'd40} : s = 150;
	{8'd110,8'd41} : s = 151;
	{8'd110,8'd42} : s = 152;
	{8'd110,8'd43} : s = 153;
	{8'd110,8'd44} : s = 154;
	{8'd110,8'd45} : s = 155;
	{8'd110,8'd46} : s = 156;
	{8'd110,8'd47} : s = 157;
	{8'd110,8'd48} : s = 158;
	{8'd110,8'd49} : s = 159;
	{8'd110,8'd50} : s = 160;
	{8'd110,8'd51} : s = 161;
	{8'd110,8'd52} : s = 162;
	{8'd110,8'd53} : s = 163;
	{8'd110,8'd54} : s = 164;
	{8'd110,8'd55} : s = 165;
	{8'd110,8'd56} : s = 166;
	{8'd110,8'd57} : s = 167;
	{8'd110,8'd58} : s = 168;
	{8'd110,8'd59} : s = 169;
	{8'd110,8'd60} : s = 170;
	{8'd110,8'd61} : s = 171;
	{8'd110,8'd62} : s = 172;
	{8'd110,8'd63} : s = 173;
	{8'd110,8'd64} : s = 174;
	{8'd110,8'd65} : s = 175;
	{8'd110,8'd66} : s = 176;
	{8'd110,8'd67} : s = 177;
	{8'd110,8'd68} : s = 178;
	{8'd110,8'd69} : s = 179;
	{8'd110,8'd70} : s = 180;
	{8'd110,8'd71} : s = 181;
	{8'd110,8'd72} : s = 182;
	{8'd110,8'd73} : s = 183;
	{8'd110,8'd74} : s = 184;
	{8'd110,8'd75} : s = 185;
	{8'd110,8'd76} : s = 186;
	{8'd110,8'd77} : s = 187;
	{8'd110,8'd78} : s = 188;
	{8'd110,8'd79} : s = 189;
	{8'd110,8'd80} : s = 190;
	{8'd110,8'd81} : s = 191;
	{8'd110,8'd82} : s = 192;
	{8'd110,8'd83} : s = 193;
	{8'd110,8'd84} : s = 194;
	{8'd110,8'd85} : s = 195;
	{8'd110,8'd86} : s = 196;
	{8'd110,8'd87} : s = 197;
	{8'd110,8'd88} : s = 198;
	{8'd110,8'd89} : s = 199;
	{8'd110,8'd90} : s = 200;
	{8'd110,8'd91} : s = 201;
	{8'd110,8'd92} : s = 202;
	{8'd110,8'd93} : s = 203;
	{8'd110,8'd94} : s = 204;
	{8'd110,8'd95} : s = 205;
	{8'd110,8'd96} : s = 206;
	{8'd110,8'd97} : s = 207;
	{8'd110,8'd98} : s = 208;
	{8'd110,8'd99} : s = 209;
	{8'd110,8'd100} : s = 210;
	{8'd110,8'd101} : s = 211;
	{8'd110,8'd102} : s = 212;
	{8'd110,8'd103} : s = 213;
	{8'd110,8'd104} : s = 214;
	{8'd110,8'd105} : s = 215;
	{8'd110,8'd106} : s = 216;
	{8'd110,8'd107} : s = 217;
	{8'd110,8'd108} : s = 218;
	{8'd110,8'd109} : s = 219;
	{8'd110,8'd110} : s = 220;
	{8'd110,8'd111} : s = 221;
	{8'd110,8'd112} : s = 222;
	{8'd110,8'd113} : s = 223;
	{8'd110,8'd114} : s = 224;
	{8'd110,8'd115} : s = 225;
	{8'd110,8'd116} : s = 226;
	{8'd110,8'd117} : s = 227;
	{8'd110,8'd118} : s = 228;
	{8'd110,8'd119} : s = 229;
	{8'd110,8'd120} : s = 230;
	{8'd110,8'd121} : s = 231;
	{8'd110,8'd122} : s = 232;
	{8'd110,8'd123} : s = 233;
	{8'd110,8'd124} : s = 234;
	{8'd110,8'd125} : s = 235;
	{8'd110,8'd126} : s = 236;
	{8'd110,8'd127} : s = 237;
	{8'd110,8'd128} : s = 238;
	{8'd110,8'd129} : s = 239;
	{8'd110,8'd130} : s = 240;
	{8'd110,8'd131} : s = 241;
	{8'd110,8'd132} : s = 242;
	{8'd110,8'd133} : s = 243;
	{8'd110,8'd134} : s = 244;
	{8'd110,8'd135} : s = 245;
	{8'd110,8'd136} : s = 246;
	{8'd110,8'd137} : s = 247;
	{8'd110,8'd138} : s = 248;
	{8'd110,8'd139} : s = 249;
	{8'd110,8'd140} : s = 250;
	{8'd110,8'd141} : s = 251;
	{8'd110,8'd142} : s = 252;
	{8'd110,8'd143} : s = 253;
	{8'd110,8'd144} : s = 254;
	{8'd110,8'd145} : s = 255;
	{8'd110,8'd146} : s = 256;
	{8'd110,8'd147} : s = 257;
	{8'd110,8'd148} : s = 258;
	{8'd110,8'd149} : s = 259;
	{8'd110,8'd150} : s = 260;
	{8'd110,8'd151} : s = 261;
	{8'd110,8'd152} : s = 262;
	{8'd110,8'd153} : s = 263;
	{8'd110,8'd154} : s = 264;
	{8'd110,8'd155} : s = 265;
	{8'd110,8'd156} : s = 266;
	{8'd110,8'd157} : s = 267;
	{8'd110,8'd158} : s = 268;
	{8'd110,8'd159} : s = 269;
	{8'd110,8'd160} : s = 270;
	{8'd110,8'd161} : s = 271;
	{8'd110,8'd162} : s = 272;
	{8'd110,8'd163} : s = 273;
	{8'd110,8'd164} : s = 274;
	{8'd110,8'd165} : s = 275;
	{8'd110,8'd166} : s = 276;
	{8'd110,8'd167} : s = 277;
	{8'd110,8'd168} : s = 278;
	{8'd110,8'd169} : s = 279;
	{8'd110,8'd170} : s = 280;
	{8'd110,8'd171} : s = 281;
	{8'd110,8'd172} : s = 282;
	{8'd110,8'd173} : s = 283;
	{8'd110,8'd174} : s = 284;
	{8'd110,8'd175} : s = 285;
	{8'd110,8'd176} : s = 286;
	{8'd110,8'd177} : s = 287;
	{8'd110,8'd178} : s = 288;
	{8'd110,8'd179} : s = 289;
	{8'd110,8'd180} : s = 290;
	{8'd110,8'd181} : s = 291;
	{8'd110,8'd182} : s = 292;
	{8'd110,8'd183} : s = 293;
	{8'd110,8'd184} : s = 294;
	{8'd110,8'd185} : s = 295;
	{8'd110,8'd186} : s = 296;
	{8'd110,8'd187} : s = 297;
	{8'd110,8'd188} : s = 298;
	{8'd110,8'd189} : s = 299;
	{8'd110,8'd190} : s = 300;
	{8'd110,8'd191} : s = 301;
	{8'd110,8'd192} : s = 302;
	{8'd110,8'd193} : s = 303;
	{8'd110,8'd194} : s = 304;
	{8'd110,8'd195} : s = 305;
	{8'd110,8'd196} : s = 306;
	{8'd110,8'd197} : s = 307;
	{8'd110,8'd198} : s = 308;
	{8'd110,8'd199} : s = 309;
	{8'd110,8'd200} : s = 310;
	{8'd110,8'd201} : s = 311;
	{8'd110,8'd202} : s = 312;
	{8'd110,8'd203} : s = 313;
	{8'd110,8'd204} : s = 314;
	{8'd110,8'd205} : s = 315;
	{8'd110,8'd206} : s = 316;
	{8'd110,8'd207} : s = 317;
	{8'd110,8'd208} : s = 318;
	{8'd110,8'd209} : s = 319;
	{8'd110,8'd210} : s = 320;
	{8'd110,8'd211} : s = 321;
	{8'd110,8'd212} : s = 322;
	{8'd110,8'd213} : s = 323;
	{8'd110,8'd214} : s = 324;
	{8'd110,8'd215} : s = 325;
	{8'd110,8'd216} : s = 326;
	{8'd110,8'd217} : s = 327;
	{8'd110,8'd218} : s = 328;
	{8'd110,8'd219} : s = 329;
	{8'd110,8'd220} : s = 330;
	{8'd110,8'd221} : s = 331;
	{8'd110,8'd222} : s = 332;
	{8'd110,8'd223} : s = 333;
	{8'd110,8'd224} : s = 334;
	{8'd110,8'd225} : s = 335;
	{8'd110,8'd226} : s = 336;
	{8'd110,8'd227} : s = 337;
	{8'd110,8'd228} : s = 338;
	{8'd110,8'd229} : s = 339;
	{8'd110,8'd230} : s = 340;
	{8'd110,8'd231} : s = 341;
	{8'd110,8'd232} : s = 342;
	{8'd110,8'd233} : s = 343;
	{8'd110,8'd234} : s = 344;
	{8'd110,8'd235} : s = 345;
	{8'd110,8'd236} : s = 346;
	{8'd110,8'd237} : s = 347;
	{8'd110,8'd238} : s = 348;
	{8'd110,8'd239} : s = 349;
	{8'd110,8'd240} : s = 350;
	{8'd110,8'd241} : s = 351;
	{8'd110,8'd242} : s = 352;
	{8'd110,8'd243} : s = 353;
	{8'd110,8'd244} : s = 354;
	{8'd110,8'd245} : s = 355;
	{8'd110,8'd246} : s = 356;
	{8'd110,8'd247} : s = 357;
	{8'd110,8'd248} : s = 358;
	{8'd110,8'd249} : s = 359;
	{8'd110,8'd250} : s = 360;
	{8'd110,8'd251} : s = 361;
	{8'd110,8'd252} : s = 362;
	{8'd110,8'd253} : s = 363;
	{8'd110,8'd254} : s = 364;
	{8'd110,8'd255} : s = 365;
	{8'd111,8'd0} : s = 111;
	{8'd111,8'd1} : s = 112;
	{8'd111,8'd2} : s = 113;
	{8'd111,8'd3} : s = 114;
	{8'd111,8'd4} : s = 115;
	{8'd111,8'd5} : s = 116;
	{8'd111,8'd6} : s = 117;
	{8'd111,8'd7} : s = 118;
	{8'd111,8'd8} : s = 119;
	{8'd111,8'd9} : s = 120;
	{8'd111,8'd10} : s = 121;
	{8'd111,8'd11} : s = 122;
	{8'd111,8'd12} : s = 123;
	{8'd111,8'd13} : s = 124;
	{8'd111,8'd14} : s = 125;
	{8'd111,8'd15} : s = 126;
	{8'd111,8'd16} : s = 127;
	{8'd111,8'd17} : s = 128;
	{8'd111,8'd18} : s = 129;
	{8'd111,8'd19} : s = 130;
	{8'd111,8'd20} : s = 131;
	{8'd111,8'd21} : s = 132;
	{8'd111,8'd22} : s = 133;
	{8'd111,8'd23} : s = 134;
	{8'd111,8'd24} : s = 135;
	{8'd111,8'd25} : s = 136;
	{8'd111,8'd26} : s = 137;
	{8'd111,8'd27} : s = 138;
	{8'd111,8'd28} : s = 139;
	{8'd111,8'd29} : s = 140;
	{8'd111,8'd30} : s = 141;
	{8'd111,8'd31} : s = 142;
	{8'd111,8'd32} : s = 143;
	{8'd111,8'd33} : s = 144;
	{8'd111,8'd34} : s = 145;
	{8'd111,8'd35} : s = 146;
	{8'd111,8'd36} : s = 147;
	{8'd111,8'd37} : s = 148;
	{8'd111,8'd38} : s = 149;
	{8'd111,8'd39} : s = 150;
	{8'd111,8'd40} : s = 151;
	{8'd111,8'd41} : s = 152;
	{8'd111,8'd42} : s = 153;
	{8'd111,8'd43} : s = 154;
	{8'd111,8'd44} : s = 155;
	{8'd111,8'd45} : s = 156;
	{8'd111,8'd46} : s = 157;
	{8'd111,8'd47} : s = 158;
	{8'd111,8'd48} : s = 159;
	{8'd111,8'd49} : s = 160;
	{8'd111,8'd50} : s = 161;
	{8'd111,8'd51} : s = 162;
	{8'd111,8'd52} : s = 163;
	{8'd111,8'd53} : s = 164;
	{8'd111,8'd54} : s = 165;
	{8'd111,8'd55} : s = 166;
	{8'd111,8'd56} : s = 167;
	{8'd111,8'd57} : s = 168;
	{8'd111,8'd58} : s = 169;
	{8'd111,8'd59} : s = 170;
	{8'd111,8'd60} : s = 171;
	{8'd111,8'd61} : s = 172;
	{8'd111,8'd62} : s = 173;
	{8'd111,8'd63} : s = 174;
	{8'd111,8'd64} : s = 175;
	{8'd111,8'd65} : s = 176;
	{8'd111,8'd66} : s = 177;
	{8'd111,8'd67} : s = 178;
	{8'd111,8'd68} : s = 179;
	{8'd111,8'd69} : s = 180;
	{8'd111,8'd70} : s = 181;
	{8'd111,8'd71} : s = 182;
	{8'd111,8'd72} : s = 183;
	{8'd111,8'd73} : s = 184;
	{8'd111,8'd74} : s = 185;
	{8'd111,8'd75} : s = 186;
	{8'd111,8'd76} : s = 187;
	{8'd111,8'd77} : s = 188;
	{8'd111,8'd78} : s = 189;
	{8'd111,8'd79} : s = 190;
	{8'd111,8'd80} : s = 191;
	{8'd111,8'd81} : s = 192;
	{8'd111,8'd82} : s = 193;
	{8'd111,8'd83} : s = 194;
	{8'd111,8'd84} : s = 195;
	{8'd111,8'd85} : s = 196;
	{8'd111,8'd86} : s = 197;
	{8'd111,8'd87} : s = 198;
	{8'd111,8'd88} : s = 199;
	{8'd111,8'd89} : s = 200;
	{8'd111,8'd90} : s = 201;
	{8'd111,8'd91} : s = 202;
	{8'd111,8'd92} : s = 203;
	{8'd111,8'd93} : s = 204;
	{8'd111,8'd94} : s = 205;
	{8'd111,8'd95} : s = 206;
	{8'd111,8'd96} : s = 207;
	{8'd111,8'd97} : s = 208;
	{8'd111,8'd98} : s = 209;
	{8'd111,8'd99} : s = 210;
	{8'd111,8'd100} : s = 211;
	{8'd111,8'd101} : s = 212;
	{8'd111,8'd102} : s = 213;
	{8'd111,8'd103} : s = 214;
	{8'd111,8'd104} : s = 215;
	{8'd111,8'd105} : s = 216;
	{8'd111,8'd106} : s = 217;
	{8'd111,8'd107} : s = 218;
	{8'd111,8'd108} : s = 219;
	{8'd111,8'd109} : s = 220;
	{8'd111,8'd110} : s = 221;
	{8'd111,8'd111} : s = 222;
	{8'd111,8'd112} : s = 223;
	{8'd111,8'd113} : s = 224;
	{8'd111,8'd114} : s = 225;
	{8'd111,8'd115} : s = 226;
	{8'd111,8'd116} : s = 227;
	{8'd111,8'd117} : s = 228;
	{8'd111,8'd118} : s = 229;
	{8'd111,8'd119} : s = 230;
	{8'd111,8'd120} : s = 231;
	{8'd111,8'd121} : s = 232;
	{8'd111,8'd122} : s = 233;
	{8'd111,8'd123} : s = 234;
	{8'd111,8'd124} : s = 235;
	{8'd111,8'd125} : s = 236;
	{8'd111,8'd126} : s = 237;
	{8'd111,8'd127} : s = 238;
	{8'd111,8'd128} : s = 239;
	{8'd111,8'd129} : s = 240;
	{8'd111,8'd130} : s = 241;
	{8'd111,8'd131} : s = 242;
	{8'd111,8'd132} : s = 243;
	{8'd111,8'd133} : s = 244;
	{8'd111,8'd134} : s = 245;
	{8'd111,8'd135} : s = 246;
	{8'd111,8'd136} : s = 247;
	{8'd111,8'd137} : s = 248;
	{8'd111,8'd138} : s = 249;
	{8'd111,8'd139} : s = 250;
	{8'd111,8'd140} : s = 251;
	{8'd111,8'd141} : s = 252;
	{8'd111,8'd142} : s = 253;
	{8'd111,8'd143} : s = 254;
	{8'd111,8'd144} : s = 255;
	{8'd111,8'd145} : s = 256;
	{8'd111,8'd146} : s = 257;
	{8'd111,8'd147} : s = 258;
	{8'd111,8'd148} : s = 259;
	{8'd111,8'd149} : s = 260;
	{8'd111,8'd150} : s = 261;
	{8'd111,8'd151} : s = 262;
	{8'd111,8'd152} : s = 263;
	{8'd111,8'd153} : s = 264;
	{8'd111,8'd154} : s = 265;
	{8'd111,8'd155} : s = 266;
	{8'd111,8'd156} : s = 267;
	{8'd111,8'd157} : s = 268;
	{8'd111,8'd158} : s = 269;
	{8'd111,8'd159} : s = 270;
	{8'd111,8'd160} : s = 271;
	{8'd111,8'd161} : s = 272;
	{8'd111,8'd162} : s = 273;
	{8'd111,8'd163} : s = 274;
	{8'd111,8'd164} : s = 275;
	{8'd111,8'd165} : s = 276;
	{8'd111,8'd166} : s = 277;
	{8'd111,8'd167} : s = 278;
	{8'd111,8'd168} : s = 279;
	{8'd111,8'd169} : s = 280;
	{8'd111,8'd170} : s = 281;
	{8'd111,8'd171} : s = 282;
	{8'd111,8'd172} : s = 283;
	{8'd111,8'd173} : s = 284;
	{8'd111,8'd174} : s = 285;
	{8'd111,8'd175} : s = 286;
	{8'd111,8'd176} : s = 287;
	{8'd111,8'd177} : s = 288;
	{8'd111,8'd178} : s = 289;
	{8'd111,8'd179} : s = 290;
	{8'd111,8'd180} : s = 291;
	{8'd111,8'd181} : s = 292;
	{8'd111,8'd182} : s = 293;
	{8'd111,8'd183} : s = 294;
	{8'd111,8'd184} : s = 295;
	{8'd111,8'd185} : s = 296;
	{8'd111,8'd186} : s = 297;
	{8'd111,8'd187} : s = 298;
	{8'd111,8'd188} : s = 299;
	{8'd111,8'd189} : s = 300;
	{8'd111,8'd190} : s = 301;
	{8'd111,8'd191} : s = 302;
	{8'd111,8'd192} : s = 303;
	{8'd111,8'd193} : s = 304;
	{8'd111,8'd194} : s = 305;
	{8'd111,8'd195} : s = 306;
	{8'd111,8'd196} : s = 307;
	{8'd111,8'd197} : s = 308;
	{8'd111,8'd198} : s = 309;
	{8'd111,8'd199} : s = 310;
	{8'd111,8'd200} : s = 311;
	{8'd111,8'd201} : s = 312;
	{8'd111,8'd202} : s = 313;
	{8'd111,8'd203} : s = 314;
	{8'd111,8'd204} : s = 315;
	{8'd111,8'd205} : s = 316;
	{8'd111,8'd206} : s = 317;
	{8'd111,8'd207} : s = 318;
	{8'd111,8'd208} : s = 319;
	{8'd111,8'd209} : s = 320;
	{8'd111,8'd210} : s = 321;
	{8'd111,8'd211} : s = 322;
	{8'd111,8'd212} : s = 323;
	{8'd111,8'd213} : s = 324;
	{8'd111,8'd214} : s = 325;
	{8'd111,8'd215} : s = 326;
	{8'd111,8'd216} : s = 327;
	{8'd111,8'd217} : s = 328;
	{8'd111,8'd218} : s = 329;
	{8'd111,8'd219} : s = 330;
	{8'd111,8'd220} : s = 331;
	{8'd111,8'd221} : s = 332;
	{8'd111,8'd222} : s = 333;
	{8'd111,8'd223} : s = 334;
	{8'd111,8'd224} : s = 335;
	{8'd111,8'd225} : s = 336;
	{8'd111,8'd226} : s = 337;
	{8'd111,8'd227} : s = 338;
	{8'd111,8'd228} : s = 339;
	{8'd111,8'd229} : s = 340;
	{8'd111,8'd230} : s = 341;
	{8'd111,8'd231} : s = 342;
	{8'd111,8'd232} : s = 343;
	{8'd111,8'd233} : s = 344;
	{8'd111,8'd234} : s = 345;
	{8'd111,8'd235} : s = 346;
	{8'd111,8'd236} : s = 347;
	{8'd111,8'd237} : s = 348;
	{8'd111,8'd238} : s = 349;
	{8'd111,8'd239} : s = 350;
	{8'd111,8'd240} : s = 351;
	{8'd111,8'd241} : s = 352;
	{8'd111,8'd242} : s = 353;
	{8'd111,8'd243} : s = 354;
	{8'd111,8'd244} : s = 355;
	{8'd111,8'd245} : s = 356;
	{8'd111,8'd246} : s = 357;
	{8'd111,8'd247} : s = 358;
	{8'd111,8'd248} : s = 359;
	{8'd111,8'd249} : s = 360;
	{8'd111,8'd250} : s = 361;
	{8'd111,8'd251} : s = 362;
	{8'd111,8'd252} : s = 363;
	{8'd111,8'd253} : s = 364;
	{8'd111,8'd254} : s = 365;
	{8'd111,8'd255} : s = 366;
	{8'd112,8'd0} : s = 112;
	{8'd112,8'd1} : s = 113;
	{8'd112,8'd2} : s = 114;
	{8'd112,8'd3} : s = 115;
	{8'd112,8'd4} : s = 116;
	{8'd112,8'd5} : s = 117;
	{8'd112,8'd6} : s = 118;
	{8'd112,8'd7} : s = 119;
	{8'd112,8'd8} : s = 120;
	{8'd112,8'd9} : s = 121;
	{8'd112,8'd10} : s = 122;
	{8'd112,8'd11} : s = 123;
	{8'd112,8'd12} : s = 124;
	{8'd112,8'd13} : s = 125;
	{8'd112,8'd14} : s = 126;
	{8'd112,8'd15} : s = 127;
	{8'd112,8'd16} : s = 128;
	{8'd112,8'd17} : s = 129;
	{8'd112,8'd18} : s = 130;
	{8'd112,8'd19} : s = 131;
	{8'd112,8'd20} : s = 132;
	{8'd112,8'd21} : s = 133;
	{8'd112,8'd22} : s = 134;
	{8'd112,8'd23} : s = 135;
	{8'd112,8'd24} : s = 136;
	{8'd112,8'd25} : s = 137;
	{8'd112,8'd26} : s = 138;
	{8'd112,8'd27} : s = 139;
	{8'd112,8'd28} : s = 140;
	{8'd112,8'd29} : s = 141;
	{8'd112,8'd30} : s = 142;
	{8'd112,8'd31} : s = 143;
	{8'd112,8'd32} : s = 144;
	{8'd112,8'd33} : s = 145;
	{8'd112,8'd34} : s = 146;
	{8'd112,8'd35} : s = 147;
	{8'd112,8'd36} : s = 148;
	{8'd112,8'd37} : s = 149;
	{8'd112,8'd38} : s = 150;
	{8'd112,8'd39} : s = 151;
	{8'd112,8'd40} : s = 152;
	{8'd112,8'd41} : s = 153;
	{8'd112,8'd42} : s = 154;
	{8'd112,8'd43} : s = 155;
	{8'd112,8'd44} : s = 156;
	{8'd112,8'd45} : s = 157;
	{8'd112,8'd46} : s = 158;
	{8'd112,8'd47} : s = 159;
	{8'd112,8'd48} : s = 160;
	{8'd112,8'd49} : s = 161;
	{8'd112,8'd50} : s = 162;
	{8'd112,8'd51} : s = 163;
	{8'd112,8'd52} : s = 164;
	{8'd112,8'd53} : s = 165;
	{8'd112,8'd54} : s = 166;
	{8'd112,8'd55} : s = 167;
	{8'd112,8'd56} : s = 168;
	{8'd112,8'd57} : s = 169;
	{8'd112,8'd58} : s = 170;
	{8'd112,8'd59} : s = 171;
	{8'd112,8'd60} : s = 172;
	{8'd112,8'd61} : s = 173;
	{8'd112,8'd62} : s = 174;
	{8'd112,8'd63} : s = 175;
	{8'd112,8'd64} : s = 176;
	{8'd112,8'd65} : s = 177;
	{8'd112,8'd66} : s = 178;
	{8'd112,8'd67} : s = 179;
	{8'd112,8'd68} : s = 180;
	{8'd112,8'd69} : s = 181;
	{8'd112,8'd70} : s = 182;
	{8'd112,8'd71} : s = 183;
	{8'd112,8'd72} : s = 184;
	{8'd112,8'd73} : s = 185;
	{8'd112,8'd74} : s = 186;
	{8'd112,8'd75} : s = 187;
	{8'd112,8'd76} : s = 188;
	{8'd112,8'd77} : s = 189;
	{8'd112,8'd78} : s = 190;
	{8'd112,8'd79} : s = 191;
	{8'd112,8'd80} : s = 192;
	{8'd112,8'd81} : s = 193;
	{8'd112,8'd82} : s = 194;
	{8'd112,8'd83} : s = 195;
	{8'd112,8'd84} : s = 196;
	{8'd112,8'd85} : s = 197;
	{8'd112,8'd86} : s = 198;
	{8'd112,8'd87} : s = 199;
	{8'd112,8'd88} : s = 200;
	{8'd112,8'd89} : s = 201;
	{8'd112,8'd90} : s = 202;
	{8'd112,8'd91} : s = 203;
	{8'd112,8'd92} : s = 204;
	{8'd112,8'd93} : s = 205;
	{8'd112,8'd94} : s = 206;
	{8'd112,8'd95} : s = 207;
	{8'd112,8'd96} : s = 208;
	{8'd112,8'd97} : s = 209;
	{8'd112,8'd98} : s = 210;
	{8'd112,8'd99} : s = 211;
	{8'd112,8'd100} : s = 212;
	{8'd112,8'd101} : s = 213;
	{8'd112,8'd102} : s = 214;
	{8'd112,8'd103} : s = 215;
	{8'd112,8'd104} : s = 216;
	{8'd112,8'd105} : s = 217;
	{8'd112,8'd106} : s = 218;
	{8'd112,8'd107} : s = 219;
	{8'd112,8'd108} : s = 220;
	{8'd112,8'd109} : s = 221;
	{8'd112,8'd110} : s = 222;
	{8'd112,8'd111} : s = 223;
	{8'd112,8'd112} : s = 224;
	{8'd112,8'd113} : s = 225;
	{8'd112,8'd114} : s = 226;
	{8'd112,8'd115} : s = 227;
	{8'd112,8'd116} : s = 228;
	{8'd112,8'd117} : s = 229;
	{8'd112,8'd118} : s = 230;
	{8'd112,8'd119} : s = 231;
	{8'd112,8'd120} : s = 232;
	{8'd112,8'd121} : s = 233;
	{8'd112,8'd122} : s = 234;
	{8'd112,8'd123} : s = 235;
	{8'd112,8'd124} : s = 236;
	{8'd112,8'd125} : s = 237;
	{8'd112,8'd126} : s = 238;
	{8'd112,8'd127} : s = 239;
	{8'd112,8'd128} : s = 240;
	{8'd112,8'd129} : s = 241;
	{8'd112,8'd130} : s = 242;
	{8'd112,8'd131} : s = 243;
	{8'd112,8'd132} : s = 244;
	{8'd112,8'd133} : s = 245;
	{8'd112,8'd134} : s = 246;
	{8'd112,8'd135} : s = 247;
	{8'd112,8'd136} : s = 248;
	{8'd112,8'd137} : s = 249;
	{8'd112,8'd138} : s = 250;
	{8'd112,8'd139} : s = 251;
	{8'd112,8'd140} : s = 252;
	{8'd112,8'd141} : s = 253;
	{8'd112,8'd142} : s = 254;
	{8'd112,8'd143} : s = 255;
	{8'd112,8'd144} : s = 256;
	{8'd112,8'd145} : s = 257;
	{8'd112,8'd146} : s = 258;
	{8'd112,8'd147} : s = 259;
	{8'd112,8'd148} : s = 260;
	{8'd112,8'd149} : s = 261;
	{8'd112,8'd150} : s = 262;
	{8'd112,8'd151} : s = 263;
	{8'd112,8'd152} : s = 264;
	{8'd112,8'd153} : s = 265;
	{8'd112,8'd154} : s = 266;
	{8'd112,8'd155} : s = 267;
	{8'd112,8'd156} : s = 268;
	{8'd112,8'd157} : s = 269;
	{8'd112,8'd158} : s = 270;
	{8'd112,8'd159} : s = 271;
	{8'd112,8'd160} : s = 272;
	{8'd112,8'd161} : s = 273;
	{8'd112,8'd162} : s = 274;
	{8'd112,8'd163} : s = 275;
	{8'd112,8'd164} : s = 276;
	{8'd112,8'd165} : s = 277;
	{8'd112,8'd166} : s = 278;
	{8'd112,8'd167} : s = 279;
	{8'd112,8'd168} : s = 280;
	{8'd112,8'd169} : s = 281;
	{8'd112,8'd170} : s = 282;
	{8'd112,8'd171} : s = 283;
	{8'd112,8'd172} : s = 284;
	{8'd112,8'd173} : s = 285;
	{8'd112,8'd174} : s = 286;
	{8'd112,8'd175} : s = 287;
	{8'd112,8'd176} : s = 288;
	{8'd112,8'd177} : s = 289;
	{8'd112,8'd178} : s = 290;
	{8'd112,8'd179} : s = 291;
	{8'd112,8'd180} : s = 292;
	{8'd112,8'd181} : s = 293;
	{8'd112,8'd182} : s = 294;
	{8'd112,8'd183} : s = 295;
	{8'd112,8'd184} : s = 296;
	{8'd112,8'd185} : s = 297;
	{8'd112,8'd186} : s = 298;
	{8'd112,8'd187} : s = 299;
	{8'd112,8'd188} : s = 300;
	{8'd112,8'd189} : s = 301;
	{8'd112,8'd190} : s = 302;
	{8'd112,8'd191} : s = 303;
	{8'd112,8'd192} : s = 304;
	{8'd112,8'd193} : s = 305;
	{8'd112,8'd194} : s = 306;
	{8'd112,8'd195} : s = 307;
	{8'd112,8'd196} : s = 308;
	{8'd112,8'd197} : s = 309;
	{8'd112,8'd198} : s = 310;
	{8'd112,8'd199} : s = 311;
	{8'd112,8'd200} : s = 312;
	{8'd112,8'd201} : s = 313;
	{8'd112,8'd202} : s = 314;
	{8'd112,8'd203} : s = 315;
	{8'd112,8'd204} : s = 316;
	{8'd112,8'd205} : s = 317;
	{8'd112,8'd206} : s = 318;
	{8'd112,8'd207} : s = 319;
	{8'd112,8'd208} : s = 320;
	{8'd112,8'd209} : s = 321;
	{8'd112,8'd210} : s = 322;
	{8'd112,8'd211} : s = 323;
	{8'd112,8'd212} : s = 324;
	{8'd112,8'd213} : s = 325;
	{8'd112,8'd214} : s = 326;
	{8'd112,8'd215} : s = 327;
	{8'd112,8'd216} : s = 328;
	{8'd112,8'd217} : s = 329;
	{8'd112,8'd218} : s = 330;
	{8'd112,8'd219} : s = 331;
	{8'd112,8'd220} : s = 332;
	{8'd112,8'd221} : s = 333;
	{8'd112,8'd222} : s = 334;
	{8'd112,8'd223} : s = 335;
	{8'd112,8'd224} : s = 336;
	{8'd112,8'd225} : s = 337;
	{8'd112,8'd226} : s = 338;
	{8'd112,8'd227} : s = 339;
	{8'd112,8'd228} : s = 340;
	{8'd112,8'd229} : s = 341;
	{8'd112,8'd230} : s = 342;
	{8'd112,8'd231} : s = 343;
	{8'd112,8'd232} : s = 344;
	{8'd112,8'd233} : s = 345;
	{8'd112,8'd234} : s = 346;
	{8'd112,8'd235} : s = 347;
	{8'd112,8'd236} : s = 348;
	{8'd112,8'd237} : s = 349;
	{8'd112,8'd238} : s = 350;
	{8'd112,8'd239} : s = 351;
	{8'd112,8'd240} : s = 352;
	{8'd112,8'd241} : s = 353;
	{8'd112,8'd242} : s = 354;
	{8'd112,8'd243} : s = 355;
	{8'd112,8'd244} : s = 356;
	{8'd112,8'd245} : s = 357;
	{8'd112,8'd246} : s = 358;
	{8'd112,8'd247} : s = 359;
	{8'd112,8'd248} : s = 360;
	{8'd112,8'd249} : s = 361;
	{8'd112,8'd250} : s = 362;
	{8'd112,8'd251} : s = 363;
	{8'd112,8'd252} : s = 364;
	{8'd112,8'd253} : s = 365;
	{8'd112,8'd254} : s = 366;
	{8'd112,8'd255} : s = 367;
	{8'd113,8'd0} : s = 113;
	{8'd113,8'd1} : s = 114;
	{8'd113,8'd2} : s = 115;
	{8'd113,8'd3} : s = 116;
	{8'd113,8'd4} : s = 117;
	{8'd113,8'd5} : s = 118;
	{8'd113,8'd6} : s = 119;
	{8'd113,8'd7} : s = 120;
	{8'd113,8'd8} : s = 121;
	{8'd113,8'd9} : s = 122;
	{8'd113,8'd10} : s = 123;
	{8'd113,8'd11} : s = 124;
	{8'd113,8'd12} : s = 125;
	{8'd113,8'd13} : s = 126;
	{8'd113,8'd14} : s = 127;
	{8'd113,8'd15} : s = 128;
	{8'd113,8'd16} : s = 129;
	{8'd113,8'd17} : s = 130;
	{8'd113,8'd18} : s = 131;
	{8'd113,8'd19} : s = 132;
	{8'd113,8'd20} : s = 133;
	{8'd113,8'd21} : s = 134;
	{8'd113,8'd22} : s = 135;
	{8'd113,8'd23} : s = 136;
	{8'd113,8'd24} : s = 137;
	{8'd113,8'd25} : s = 138;
	{8'd113,8'd26} : s = 139;
	{8'd113,8'd27} : s = 140;
	{8'd113,8'd28} : s = 141;
	{8'd113,8'd29} : s = 142;
	{8'd113,8'd30} : s = 143;
	{8'd113,8'd31} : s = 144;
	{8'd113,8'd32} : s = 145;
	{8'd113,8'd33} : s = 146;
	{8'd113,8'd34} : s = 147;
	{8'd113,8'd35} : s = 148;
	{8'd113,8'd36} : s = 149;
	{8'd113,8'd37} : s = 150;
	{8'd113,8'd38} : s = 151;
	{8'd113,8'd39} : s = 152;
	{8'd113,8'd40} : s = 153;
	{8'd113,8'd41} : s = 154;
	{8'd113,8'd42} : s = 155;
	{8'd113,8'd43} : s = 156;
	{8'd113,8'd44} : s = 157;
	{8'd113,8'd45} : s = 158;
	{8'd113,8'd46} : s = 159;
	{8'd113,8'd47} : s = 160;
	{8'd113,8'd48} : s = 161;
	{8'd113,8'd49} : s = 162;
	{8'd113,8'd50} : s = 163;
	{8'd113,8'd51} : s = 164;
	{8'd113,8'd52} : s = 165;
	{8'd113,8'd53} : s = 166;
	{8'd113,8'd54} : s = 167;
	{8'd113,8'd55} : s = 168;
	{8'd113,8'd56} : s = 169;
	{8'd113,8'd57} : s = 170;
	{8'd113,8'd58} : s = 171;
	{8'd113,8'd59} : s = 172;
	{8'd113,8'd60} : s = 173;
	{8'd113,8'd61} : s = 174;
	{8'd113,8'd62} : s = 175;
	{8'd113,8'd63} : s = 176;
	{8'd113,8'd64} : s = 177;
	{8'd113,8'd65} : s = 178;
	{8'd113,8'd66} : s = 179;
	{8'd113,8'd67} : s = 180;
	{8'd113,8'd68} : s = 181;
	{8'd113,8'd69} : s = 182;
	{8'd113,8'd70} : s = 183;
	{8'd113,8'd71} : s = 184;
	{8'd113,8'd72} : s = 185;
	{8'd113,8'd73} : s = 186;
	{8'd113,8'd74} : s = 187;
	{8'd113,8'd75} : s = 188;
	{8'd113,8'd76} : s = 189;
	{8'd113,8'd77} : s = 190;
	{8'd113,8'd78} : s = 191;
	{8'd113,8'd79} : s = 192;
	{8'd113,8'd80} : s = 193;
	{8'd113,8'd81} : s = 194;
	{8'd113,8'd82} : s = 195;
	{8'd113,8'd83} : s = 196;
	{8'd113,8'd84} : s = 197;
	{8'd113,8'd85} : s = 198;
	{8'd113,8'd86} : s = 199;
	{8'd113,8'd87} : s = 200;
	{8'd113,8'd88} : s = 201;
	{8'd113,8'd89} : s = 202;
	{8'd113,8'd90} : s = 203;
	{8'd113,8'd91} : s = 204;
	{8'd113,8'd92} : s = 205;
	{8'd113,8'd93} : s = 206;
	{8'd113,8'd94} : s = 207;
	{8'd113,8'd95} : s = 208;
	{8'd113,8'd96} : s = 209;
	{8'd113,8'd97} : s = 210;
	{8'd113,8'd98} : s = 211;
	{8'd113,8'd99} : s = 212;
	{8'd113,8'd100} : s = 213;
	{8'd113,8'd101} : s = 214;
	{8'd113,8'd102} : s = 215;
	{8'd113,8'd103} : s = 216;
	{8'd113,8'd104} : s = 217;
	{8'd113,8'd105} : s = 218;
	{8'd113,8'd106} : s = 219;
	{8'd113,8'd107} : s = 220;
	{8'd113,8'd108} : s = 221;
	{8'd113,8'd109} : s = 222;
	{8'd113,8'd110} : s = 223;
	{8'd113,8'd111} : s = 224;
	{8'd113,8'd112} : s = 225;
	{8'd113,8'd113} : s = 226;
	{8'd113,8'd114} : s = 227;
	{8'd113,8'd115} : s = 228;
	{8'd113,8'd116} : s = 229;
	{8'd113,8'd117} : s = 230;
	{8'd113,8'd118} : s = 231;
	{8'd113,8'd119} : s = 232;
	{8'd113,8'd120} : s = 233;
	{8'd113,8'd121} : s = 234;
	{8'd113,8'd122} : s = 235;
	{8'd113,8'd123} : s = 236;
	{8'd113,8'd124} : s = 237;
	{8'd113,8'd125} : s = 238;
	{8'd113,8'd126} : s = 239;
	{8'd113,8'd127} : s = 240;
	{8'd113,8'd128} : s = 241;
	{8'd113,8'd129} : s = 242;
	{8'd113,8'd130} : s = 243;
	{8'd113,8'd131} : s = 244;
	{8'd113,8'd132} : s = 245;
	{8'd113,8'd133} : s = 246;
	{8'd113,8'd134} : s = 247;
	{8'd113,8'd135} : s = 248;
	{8'd113,8'd136} : s = 249;
	{8'd113,8'd137} : s = 250;
	{8'd113,8'd138} : s = 251;
	{8'd113,8'd139} : s = 252;
	{8'd113,8'd140} : s = 253;
	{8'd113,8'd141} : s = 254;
	{8'd113,8'd142} : s = 255;
	{8'd113,8'd143} : s = 256;
	{8'd113,8'd144} : s = 257;
	{8'd113,8'd145} : s = 258;
	{8'd113,8'd146} : s = 259;
	{8'd113,8'd147} : s = 260;
	{8'd113,8'd148} : s = 261;
	{8'd113,8'd149} : s = 262;
	{8'd113,8'd150} : s = 263;
	{8'd113,8'd151} : s = 264;
	{8'd113,8'd152} : s = 265;
	{8'd113,8'd153} : s = 266;
	{8'd113,8'd154} : s = 267;
	{8'd113,8'd155} : s = 268;
	{8'd113,8'd156} : s = 269;
	{8'd113,8'd157} : s = 270;
	{8'd113,8'd158} : s = 271;
	{8'd113,8'd159} : s = 272;
	{8'd113,8'd160} : s = 273;
	{8'd113,8'd161} : s = 274;
	{8'd113,8'd162} : s = 275;
	{8'd113,8'd163} : s = 276;
	{8'd113,8'd164} : s = 277;
	{8'd113,8'd165} : s = 278;
	{8'd113,8'd166} : s = 279;
	{8'd113,8'd167} : s = 280;
	{8'd113,8'd168} : s = 281;
	{8'd113,8'd169} : s = 282;
	{8'd113,8'd170} : s = 283;
	{8'd113,8'd171} : s = 284;
	{8'd113,8'd172} : s = 285;
	{8'd113,8'd173} : s = 286;
	{8'd113,8'd174} : s = 287;
	{8'd113,8'd175} : s = 288;
	{8'd113,8'd176} : s = 289;
	{8'd113,8'd177} : s = 290;
	{8'd113,8'd178} : s = 291;
	{8'd113,8'd179} : s = 292;
	{8'd113,8'd180} : s = 293;
	{8'd113,8'd181} : s = 294;
	{8'd113,8'd182} : s = 295;
	{8'd113,8'd183} : s = 296;
	{8'd113,8'd184} : s = 297;
	{8'd113,8'd185} : s = 298;
	{8'd113,8'd186} : s = 299;
	{8'd113,8'd187} : s = 300;
	{8'd113,8'd188} : s = 301;
	{8'd113,8'd189} : s = 302;
	{8'd113,8'd190} : s = 303;
	{8'd113,8'd191} : s = 304;
	{8'd113,8'd192} : s = 305;
	{8'd113,8'd193} : s = 306;
	{8'd113,8'd194} : s = 307;
	{8'd113,8'd195} : s = 308;
	{8'd113,8'd196} : s = 309;
	{8'd113,8'd197} : s = 310;
	{8'd113,8'd198} : s = 311;
	{8'd113,8'd199} : s = 312;
	{8'd113,8'd200} : s = 313;
	{8'd113,8'd201} : s = 314;
	{8'd113,8'd202} : s = 315;
	{8'd113,8'd203} : s = 316;
	{8'd113,8'd204} : s = 317;
	{8'd113,8'd205} : s = 318;
	{8'd113,8'd206} : s = 319;
	{8'd113,8'd207} : s = 320;
	{8'd113,8'd208} : s = 321;
	{8'd113,8'd209} : s = 322;
	{8'd113,8'd210} : s = 323;
	{8'd113,8'd211} : s = 324;
	{8'd113,8'd212} : s = 325;
	{8'd113,8'd213} : s = 326;
	{8'd113,8'd214} : s = 327;
	{8'd113,8'd215} : s = 328;
	{8'd113,8'd216} : s = 329;
	{8'd113,8'd217} : s = 330;
	{8'd113,8'd218} : s = 331;
	{8'd113,8'd219} : s = 332;
	{8'd113,8'd220} : s = 333;
	{8'd113,8'd221} : s = 334;
	{8'd113,8'd222} : s = 335;
	{8'd113,8'd223} : s = 336;
	{8'd113,8'd224} : s = 337;
	{8'd113,8'd225} : s = 338;
	{8'd113,8'd226} : s = 339;
	{8'd113,8'd227} : s = 340;
	{8'd113,8'd228} : s = 341;
	{8'd113,8'd229} : s = 342;
	{8'd113,8'd230} : s = 343;
	{8'd113,8'd231} : s = 344;
	{8'd113,8'd232} : s = 345;
	{8'd113,8'd233} : s = 346;
	{8'd113,8'd234} : s = 347;
	{8'd113,8'd235} : s = 348;
	{8'd113,8'd236} : s = 349;
	{8'd113,8'd237} : s = 350;
	{8'd113,8'd238} : s = 351;
	{8'd113,8'd239} : s = 352;
	{8'd113,8'd240} : s = 353;
	{8'd113,8'd241} : s = 354;
	{8'd113,8'd242} : s = 355;
	{8'd113,8'd243} : s = 356;
	{8'd113,8'd244} : s = 357;
	{8'd113,8'd245} : s = 358;
	{8'd113,8'd246} : s = 359;
	{8'd113,8'd247} : s = 360;
	{8'd113,8'd248} : s = 361;
	{8'd113,8'd249} : s = 362;
	{8'd113,8'd250} : s = 363;
	{8'd113,8'd251} : s = 364;
	{8'd113,8'd252} : s = 365;
	{8'd113,8'd253} : s = 366;
	{8'd113,8'd254} : s = 367;
	{8'd113,8'd255} : s = 368;
	{8'd114,8'd0} : s = 114;
	{8'd114,8'd1} : s = 115;
	{8'd114,8'd2} : s = 116;
	{8'd114,8'd3} : s = 117;
	{8'd114,8'd4} : s = 118;
	{8'd114,8'd5} : s = 119;
	{8'd114,8'd6} : s = 120;
	{8'd114,8'd7} : s = 121;
	{8'd114,8'd8} : s = 122;
	{8'd114,8'd9} : s = 123;
	{8'd114,8'd10} : s = 124;
	{8'd114,8'd11} : s = 125;
	{8'd114,8'd12} : s = 126;
	{8'd114,8'd13} : s = 127;
	{8'd114,8'd14} : s = 128;
	{8'd114,8'd15} : s = 129;
	{8'd114,8'd16} : s = 130;
	{8'd114,8'd17} : s = 131;
	{8'd114,8'd18} : s = 132;
	{8'd114,8'd19} : s = 133;
	{8'd114,8'd20} : s = 134;
	{8'd114,8'd21} : s = 135;
	{8'd114,8'd22} : s = 136;
	{8'd114,8'd23} : s = 137;
	{8'd114,8'd24} : s = 138;
	{8'd114,8'd25} : s = 139;
	{8'd114,8'd26} : s = 140;
	{8'd114,8'd27} : s = 141;
	{8'd114,8'd28} : s = 142;
	{8'd114,8'd29} : s = 143;
	{8'd114,8'd30} : s = 144;
	{8'd114,8'd31} : s = 145;
	{8'd114,8'd32} : s = 146;
	{8'd114,8'd33} : s = 147;
	{8'd114,8'd34} : s = 148;
	{8'd114,8'd35} : s = 149;
	{8'd114,8'd36} : s = 150;
	{8'd114,8'd37} : s = 151;
	{8'd114,8'd38} : s = 152;
	{8'd114,8'd39} : s = 153;
	{8'd114,8'd40} : s = 154;
	{8'd114,8'd41} : s = 155;
	{8'd114,8'd42} : s = 156;
	{8'd114,8'd43} : s = 157;
	{8'd114,8'd44} : s = 158;
	{8'd114,8'd45} : s = 159;
	{8'd114,8'd46} : s = 160;
	{8'd114,8'd47} : s = 161;
	{8'd114,8'd48} : s = 162;
	{8'd114,8'd49} : s = 163;
	{8'd114,8'd50} : s = 164;
	{8'd114,8'd51} : s = 165;
	{8'd114,8'd52} : s = 166;
	{8'd114,8'd53} : s = 167;
	{8'd114,8'd54} : s = 168;
	{8'd114,8'd55} : s = 169;
	{8'd114,8'd56} : s = 170;
	{8'd114,8'd57} : s = 171;
	{8'd114,8'd58} : s = 172;
	{8'd114,8'd59} : s = 173;
	{8'd114,8'd60} : s = 174;
	{8'd114,8'd61} : s = 175;
	{8'd114,8'd62} : s = 176;
	{8'd114,8'd63} : s = 177;
	{8'd114,8'd64} : s = 178;
	{8'd114,8'd65} : s = 179;
	{8'd114,8'd66} : s = 180;
	{8'd114,8'd67} : s = 181;
	{8'd114,8'd68} : s = 182;
	{8'd114,8'd69} : s = 183;
	{8'd114,8'd70} : s = 184;
	{8'd114,8'd71} : s = 185;
	{8'd114,8'd72} : s = 186;
	{8'd114,8'd73} : s = 187;
	{8'd114,8'd74} : s = 188;
	{8'd114,8'd75} : s = 189;
	{8'd114,8'd76} : s = 190;
	{8'd114,8'd77} : s = 191;
	{8'd114,8'd78} : s = 192;
	{8'd114,8'd79} : s = 193;
	{8'd114,8'd80} : s = 194;
	{8'd114,8'd81} : s = 195;
	{8'd114,8'd82} : s = 196;
	{8'd114,8'd83} : s = 197;
	{8'd114,8'd84} : s = 198;
	{8'd114,8'd85} : s = 199;
	{8'd114,8'd86} : s = 200;
	{8'd114,8'd87} : s = 201;
	{8'd114,8'd88} : s = 202;
	{8'd114,8'd89} : s = 203;
	{8'd114,8'd90} : s = 204;
	{8'd114,8'd91} : s = 205;
	{8'd114,8'd92} : s = 206;
	{8'd114,8'd93} : s = 207;
	{8'd114,8'd94} : s = 208;
	{8'd114,8'd95} : s = 209;
	{8'd114,8'd96} : s = 210;
	{8'd114,8'd97} : s = 211;
	{8'd114,8'd98} : s = 212;
	{8'd114,8'd99} : s = 213;
	{8'd114,8'd100} : s = 214;
	{8'd114,8'd101} : s = 215;
	{8'd114,8'd102} : s = 216;
	{8'd114,8'd103} : s = 217;
	{8'd114,8'd104} : s = 218;
	{8'd114,8'd105} : s = 219;
	{8'd114,8'd106} : s = 220;
	{8'd114,8'd107} : s = 221;
	{8'd114,8'd108} : s = 222;
	{8'd114,8'd109} : s = 223;
	{8'd114,8'd110} : s = 224;
	{8'd114,8'd111} : s = 225;
	{8'd114,8'd112} : s = 226;
	{8'd114,8'd113} : s = 227;
	{8'd114,8'd114} : s = 228;
	{8'd114,8'd115} : s = 229;
	{8'd114,8'd116} : s = 230;
	{8'd114,8'd117} : s = 231;
	{8'd114,8'd118} : s = 232;
	{8'd114,8'd119} : s = 233;
	{8'd114,8'd120} : s = 234;
	{8'd114,8'd121} : s = 235;
	{8'd114,8'd122} : s = 236;
	{8'd114,8'd123} : s = 237;
	{8'd114,8'd124} : s = 238;
	{8'd114,8'd125} : s = 239;
	{8'd114,8'd126} : s = 240;
	{8'd114,8'd127} : s = 241;
	{8'd114,8'd128} : s = 242;
	{8'd114,8'd129} : s = 243;
	{8'd114,8'd130} : s = 244;
	{8'd114,8'd131} : s = 245;
	{8'd114,8'd132} : s = 246;
	{8'd114,8'd133} : s = 247;
	{8'd114,8'd134} : s = 248;
	{8'd114,8'd135} : s = 249;
	{8'd114,8'd136} : s = 250;
	{8'd114,8'd137} : s = 251;
	{8'd114,8'd138} : s = 252;
	{8'd114,8'd139} : s = 253;
	{8'd114,8'd140} : s = 254;
	{8'd114,8'd141} : s = 255;
	{8'd114,8'd142} : s = 256;
	{8'd114,8'd143} : s = 257;
	{8'd114,8'd144} : s = 258;
	{8'd114,8'd145} : s = 259;
	{8'd114,8'd146} : s = 260;
	{8'd114,8'd147} : s = 261;
	{8'd114,8'd148} : s = 262;
	{8'd114,8'd149} : s = 263;
	{8'd114,8'd150} : s = 264;
	{8'd114,8'd151} : s = 265;
	{8'd114,8'd152} : s = 266;
	{8'd114,8'd153} : s = 267;
	{8'd114,8'd154} : s = 268;
	{8'd114,8'd155} : s = 269;
	{8'd114,8'd156} : s = 270;
	{8'd114,8'd157} : s = 271;
	{8'd114,8'd158} : s = 272;
	{8'd114,8'd159} : s = 273;
	{8'd114,8'd160} : s = 274;
	{8'd114,8'd161} : s = 275;
	{8'd114,8'd162} : s = 276;
	{8'd114,8'd163} : s = 277;
	{8'd114,8'd164} : s = 278;
	{8'd114,8'd165} : s = 279;
	{8'd114,8'd166} : s = 280;
	{8'd114,8'd167} : s = 281;
	{8'd114,8'd168} : s = 282;
	{8'd114,8'd169} : s = 283;
	{8'd114,8'd170} : s = 284;
	{8'd114,8'd171} : s = 285;
	{8'd114,8'd172} : s = 286;
	{8'd114,8'd173} : s = 287;
	{8'd114,8'd174} : s = 288;
	{8'd114,8'd175} : s = 289;
	{8'd114,8'd176} : s = 290;
	{8'd114,8'd177} : s = 291;
	{8'd114,8'd178} : s = 292;
	{8'd114,8'd179} : s = 293;
	{8'd114,8'd180} : s = 294;
	{8'd114,8'd181} : s = 295;
	{8'd114,8'd182} : s = 296;
	{8'd114,8'd183} : s = 297;
	{8'd114,8'd184} : s = 298;
	{8'd114,8'd185} : s = 299;
	{8'd114,8'd186} : s = 300;
	{8'd114,8'd187} : s = 301;
	{8'd114,8'd188} : s = 302;
	{8'd114,8'd189} : s = 303;
	{8'd114,8'd190} : s = 304;
	{8'd114,8'd191} : s = 305;
	{8'd114,8'd192} : s = 306;
	{8'd114,8'd193} : s = 307;
	{8'd114,8'd194} : s = 308;
	{8'd114,8'd195} : s = 309;
	{8'd114,8'd196} : s = 310;
	{8'd114,8'd197} : s = 311;
	{8'd114,8'd198} : s = 312;
	{8'd114,8'd199} : s = 313;
	{8'd114,8'd200} : s = 314;
	{8'd114,8'd201} : s = 315;
	{8'd114,8'd202} : s = 316;
	{8'd114,8'd203} : s = 317;
	{8'd114,8'd204} : s = 318;
	{8'd114,8'd205} : s = 319;
	{8'd114,8'd206} : s = 320;
	{8'd114,8'd207} : s = 321;
	{8'd114,8'd208} : s = 322;
	{8'd114,8'd209} : s = 323;
	{8'd114,8'd210} : s = 324;
	{8'd114,8'd211} : s = 325;
	{8'd114,8'd212} : s = 326;
	{8'd114,8'd213} : s = 327;
	{8'd114,8'd214} : s = 328;
	{8'd114,8'd215} : s = 329;
	{8'd114,8'd216} : s = 330;
	{8'd114,8'd217} : s = 331;
	{8'd114,8'd218} : s = 332;
	{8'd114,8'd219} : s = 333;
	{8'd114,8'd220} : s = 334;
	{8'd114,8'd221} : s = 335;
	{8'd114,8'd222} : s = 336;
	{8'd114,8'd223} : s = 337;
	{8'd114,8'd224} : s = 338;
	{8'd114,8'd225} : s = 339;
	{8'd114,8'd226} : s = 340;
	{8'd114,8'd227} : s = 341;
	{8'd114,8'd228} : s = 342;
	{8'd114,8'd229} : s = 343;
	{8'd114,8'd230} : s = 344;
	{8'd114,8'd231} : s = 345;
	{8'd114,8'd232} : s = 346;
	{8'd114,8'd233} : s = 347;
	{8'd114,8'd234} : s = 348;
	{8'd114,8'd235} : s = 349;
	{8'd114,8'd236} : s = 350;
	{8'd114,8'd237} : s = 351;
	{8'd114,8'd238} : s = 352;
	{8'd114,8'd239} : s = 353;
	{8'd114,8'd240} : s = 354;
	{8'd114,8'd241} : s = 355;
	{8'd114,8'd242} : s = 356;
	{8'd114,8'd243} : s = 357;
	{8'd114,8'd244} : s = 358;
	{8'd114,8'd245} : s = 359;
	{8'd114,8'd246} : s = 360;
	{8'd114,8'd247} : s = 361;
	{8'd114,8'd248} : s = 362;
	{8'd114,8'd249} : s = 363;
	{8'd114,8'd250} : s = 364;
	{8'd114,8'd251} : s = 365;
	{8'd114,8'd252} : s = 366;
	{8'd114,8'd253} : s = 367;
	{8'd114,8'd254} : s = 368;
	{8'd114,8'd255} : s = 369;
	{8'd115,8'd0} : s = 115;
	{8'd115,8'd1} : s = 116;
	{8'd115,8'd2} : s = 117;
	{8'd115,8'd3} : s = 118;
	{8'd115,8'd4} : s = 119;
	{8'd115,8'd5} : s = 120;
	{8'd115,8'd6} : s = 121;
	{8'd115,8'd7} : s = 122;
	{8'd115,8'd8} : s = 123;
	{8'd115,8'd9} : s = 124;
	{8'd115,8'd10} : s = 125;
	{8'd115,8'd11} : s = 126;
	{8'd115,8'd12} : s = 127;
	{8'd115,8'd13} : s = 128;
	{8'd115,8'd14} : s = 129;
	{8'd115,8'd15} : s = 130;
	{8'd115,8'd16} : s = 131;
	{8'd115,8'd17} : s = 132;
	{8'd115,8'd18} : s = 133;
	{8'd115,8'd19} : s = 134;
	{8'd115,8'd20} : s = 135;
	{8'd115,8'd21} : s = 136;
	{8'd115,8'd22} : s = 137;
	{8'd115,8'd23} : s = 138;
	{8'd115,8'd24} : s = 139;
	{8'd115,8'd25} : s = 140;
	{8'd115,8'd26} : s = 141;
	{8'd115,8'd27} : s = 142;
	{8'd115,8'd28} : s = 143;
	{8'd115,8'd29} : s = 144;
	{8'd115,8'd30} : s = 145;
	{8'd115,8'd31} : s = 146;
	{8'd115,8'd32} : s = 147;
	{8'd115,8'd33} : s = 148;
	{8'd115,8'd34} : s = 149;
	{8'd115,8'd35} : s = 150;
	{8'd115,8'd36} : s = 151;
	{8'd115,8'd37} : s = 152;
	{8'd115,8'd38} : s = 153;
	{8'd115,8'd39} : s = 154;
	{8'd115,8'd40} : s = 155;
	{8'd115,8'd41} : s = 156;
	{8'd115,8'd42} : s = 157;
	{8'd115,8'd43} : s = 158;
	{8'd115,8'd44} : s = 159;
	{8'd115,8'd45} : s = 160;
	{8'd115,8'd46} : s = 161;
	{8'd115,8'd47} : s = 162;
	{8'd115,8'd48} : s = 163;
	{8'd115,8'd49} : s = 164;
	{8'd115,8'd50} : s = 165;
	{8'd115,8'd51} : s = 166;
	{8'd115,8'd52} : s = 167;
	{8'd115,8'd53} : s = 168;
	{8'd115,8'd54} : s = 169;
	{8'd115,8'd55} : s = 170;
	{8'd115,8'd56} : s = 171;
	{8'd115,8'd57} : s = 172;
	{8'd115,8'd58} : s = 173;
	{8'd115,8'd59} : s = 174;
	{8'd115,8'd60} : s = 175;
	{8'd115,8'd61} : s = 176;
	{8'd115,8'd62} : s = 177;
	{8'd115,8'd63} : s = 178;
	{8'd115,8'd64} : s = 179;
	{8'd115,8'd65} : s = 180;
	{8'd115,8'd66} : s = 181;
	{8'd115,8'd67} : s = 182;
	{8'd115,8'd68} : s = 183;
	{8'd115,8'd69} : s = 184;
	{8'd115,8'd70} : s = 185;
	{8'd115,8'd71} : s = 186;
	{8'd115,8'd72} : s = 187;
	{8'd115,8'd73} : s = 188;
	{8'd115,8'd74} : s = 189;
	{8'd115,8'd75} : s = 190;
	{8'd115,8'd76} : s = 191;
	{8'd115,8'd77} : s = 192;
	{8'd115,8'd78} : s = 193;
	{8'd115,8'd79} : s = 194;
	{8'd115,8'd80} : s = 195;
	{8'd115,8'd81} : s = 196;
	{8'd115,8'd82} : s = 197;
	{8'd115,8'd83} : s = 198;
	{8'd115,8'd84} : s = 199;
	{8'd115,8'd85} : s = 200;
	{8'd115,8'd86} : s = 201;
	{8'd115,8'd87} : s = 202;
	{8'd115,8'd88} : s = 203;
	{8'd115,8'd89} : s = 204;
	{8'd115,8'd90} : s = 205;
	{8'd115,8'd91} : s = 206;
	{8'd115,8'd92} : s = 207;
	{8'd115,8'd93} : s = 208;
	{8'd115,8'd94} : s = 209;
	{8'd115,8'd95} : s = 210;
	{8'd115,8'd96} : s = 211;
	{8'd115,8'd97} : s = 212;
	{8'd115,8'd98} : s = 213;
	{8'd115,8'd99} : s = 214;
	{8'd115,8'd100} : s = 215;
	{8'd115,8'd101} : s = 216;
	{8'd115,8'd102} : s = 217;
	{8'd115,8'd103} : s = 218;
	{8'd115,8'd104} : s = 219;
	{8'd115,8'd105} : s = 220;
	{8'd115,8'd106} : s = 221;
	{8'd115,8'd107} : s = 222;
	{8'd115,8'd108} : s = 223;
	{8'd115,8'd109} : s = 224;
	{8'd115,8'd110} : s = 225;
	{8'd115,8'd111} : s = 226;
	{8'd115,8'd112} : s = 227;
	{8'd115,8'd113} : s = 228;
	{8'd115,8'd114} : s = 229;
	{8'd115,8'd115} : s = 230;
	{8'd115,8'd116} : s = 231;
	{8'd115,8'd117} : s = 232;
	{8'd115,8'd118} : s = 233;
	{8'd115,8'd119} : s = 234;
	{8'd115,8'd120} : s = 235;
	{8'd115,8'd121} : s = 236;
	{8'd115,8'd122} : s = 237;
	{8'd115,8'd123} : s = 238;
	{8'd115,8'd124} : s = 239;
	{8'd115,8'd125} : s = 240;
	{8'd115,8'd126} : s = 241;
	{8'd115,8'd127} : s = 242;
	{8'd115,8'd128} : s = 243;
	{8'd115,8'd129} : s = 244;
	{8'd115,8'd130} : s = 245;
	{8'd115,8'd131} : s = 246;
	{8'd115,8'd132} : s = 247;
	{8'd115,8'd133} : s = 248;
	{8'd115,8'd134} : s = 249;
	{8'd115,8'd135} : s = 250;
	{8'd115,8'd136} : s = 251;
	{8'd115,8'd137} : s = 252;
	{8'd115,8'd138} : s = 253;
	{8'd115,8'd139} : s = 254;
	{8'd115,8'd140} : s = 255;
	{8'd115,8'd141} : s = 256;
	{8'd115,8'd142} : s = 257;
	{8'd115,8'd143} : s = 258;
	{8'd115,8'd144} : s = 259;
	{8'd115,8'd145} : s = 260;
	{8'd115,8'd146} : s = 261;
	{8'd115,8'd147} : s = 262;
	{8'd115,8'd148} : s = 263;
	{8'd115,8'd149} : s = 264;
	{8'd115,8'd150} : s = 265;
	{8'd115,8'd151} : s = 266;
	{8'd115,8'd152} : s = 267;
	{8'd115,8'd153} : s = 268;
	{8'd115,8'd154} : s = 269;
	{8'd115,8'd155} : s = 270;
	{8'd115,8'd156} : s = 271;
	{8'd115,8'd157} : s = 272;
	{8'd115,8'd158} : s = 273;
	{8'd115,8'd159} : s = 274;
	{8'd115,8'd160} : s = 275;
	{8'd115,8'd161} : s = 276;
	{8'd115,8'd162} : s = 277;
	{8'd115,8'd163} : s = 278;
	{8'd115,8'd164} : s = 279;
	{8'd115,8'd165} : s = 280;
	{8'd115,8'd166} : s = 281;
	{8'd115,8'd167} : s = 282;
	{8'd115,8'd168} : s = 283;
	{8'd115,8'd169} : s = 284;
	{8'd115,8'd170} : s = 285;
	{8'd115,8'd171} : s = 286;
	{8'd115,8'd172} : s = 287;
	{8'd115,8'd173} : s = 288;
	{8'd115,8'd174} : s = 289;
	{8'd115,8'd175} : s = 290;
	{8'd115,8'd176} : s = 291;
	{8'd115,8'd177} : s = 292;
	{8'd115,8'd178} : s = 293;
	{8'd115,8'd179} : s = 294;
	{8'd115,8'd180} : s = 295;
	{8'd115,8'd181} : s = 296;
	{8'd115,8'd182} : s = 297;
	{8'd115,8'd183} : s = 298;
	{8'd115,8'd184} : s = 299;
	{8'd115,8'd185} : s = 300;
	{8'd115,8'd186} : s = 301;
	{8'd115,8'd187} : s = 302;
	{8'd115,8'd188} : s = 303;
	{8'd115,8'd189} : s = 304;
	{8'd115,8'd190} : s = 305;
	{8'd115,8'd191} : s = 306;
	{8'd115,8'd192} : s = 307;
	{8'd115,8'd193} : s = 308;
	{8'd115,8'd194} : s = 309;
	{8'd115,8'd195} : s = 310;
	{8'd115,8'd196} : s = 311;
	{8'd115,8'd197} : s = 312;
	{8'd115,8'd198} : s = 313;
	{8'd115,8'd199} : s = 314;
	{8'd115,8'd200} : s = 315;
	{8'd115,8'd201} : s = 316;
	{8'd115,8'd202} : s = 317;
	{8'd115,8'd203} : s = 318;
	{8'd115,8'd204} : s = 319;
	{8'd115,8'd205} : s = 320;
	{8'd115,8'd206} : s = 321;
	{8'd115,8'd207} : s = 322;
	{8'd115,8'd208} : s = 323;
	{8'd115,8'd209} : s = 324;
	{8'd115,8'd210} : s = 325;
	{8'd115,8'd211} : s = 326;
	{8'd115,8'd212} : s = 327;
	{8'd115,8'd213} : s = 328;
	{8'd115,8'd214} : s = 329;
	{8'd115,8'd215} : s = 330;
	{8'd115,8'd216} : s = 331;
	{8'd115,8'd217} : s = 332;
	{8'd115,8'd218} : s = 333;
	{8'd115,8'd219} : s = 334;
	{8'd115,8'd220} : s = 335;
	{8'd115,8'd221} : s = 336;
	{8'd115,8'd222} : s = 337;
	{8'd115,8'd223} : s = 338;
	{8'd115,8'd224} : s = 339;
	{8'd115,8'd225} : s = 340;
	{8'd115,8'd226} : s = 341;
	{8'd115,8'd227} : s = 342;
	{8'd115,8'd228} : s = 343;
	{8'd115,8'd229} : s = 344;
	{8'd115,8'd230} : s = 345;
	{8'd115,8'd231} : s = 346;
	{8'd115,8'd232} : s = 347;
	{8'd115,8'd233} : s = 348;
	{8'd115,8'd234} : s = 349;
	{8'd115,8'd235} : s = 350;
	{8'd115,8'd236} : s = 351;
	{8'd115,8'd237} : s = 352;
	{8'd115,8'd238} : s = 353;
	{8'd115,8'd239} : s = 354;
	{8'd115,8'd240} : s = 355;
	{8'd115,8'd241} : s = 356;
	{8'd115,8'd242} : s = 357;
	{8'd115,8'd243} : s = 358;
	{8'd115,8'd244} : s = 359;
	{8'd115,8'd245} : s = 360;
	{8'd115,8'd246} : s = 361;
	{8'd115,8'd247} : s = 362;
	{8'd115,8'd248} : s = 363;
	{8'd115,8'd249} : s = 364;
	{8'd115,8'd250} : s = 365;
	{8'd115,8'd251} : s = 366;
	{8'd115,8'd252} : s = 367;
	{8'd115,8'd253} : s = 368;
	{8'd115,8'd254} : s = 369;
	{8'd115,8'd255} : s = 370;
	{8'd116,8'd0} : s = 116;
	{8'd116,8'd1} : s = 117;
	{8'd116,8'd2} : s = 118;
	{8'd116,8'd3} : s = 119;
	{8'd116,8'd4} : s = 120;
	{8'd116,8'd5} : s = 121;
	{8'd116,8'd6} : s = 122;
	{8'd116,8'd7} : s = 123;
	{8'd116,8'd8} : s = 124;
	{8'd116,8'd9} : s = 125;
	{8'd116,8'd10} : s = 126;
	{8'd116,8'd11} : s = 127;
	{8'd116,8'd12} : s = 128;
	{8'd116,8'd13} : s = 129;
	{8'd116,8'd14} : s = 130;
	{8'd116,8'd15} : s = 131;
	{8'd116,8'd16} : s = 132;
	{8'd116,8'd17} : s = 133;
	{8'd116,8'd18} : s = 134;
	{8'd116,8'd19} : s = 135;
	{8'd116,8'd20} : s = 136;
	{8'd116,8'd21} : s = 137;
	{8'd116,8'd22} : s = 138;
	{8'd116,8'd23} : s = 139;
	{8'd116,8'd24} : s = 140;
	{8'd116,8'd25} : s = 141;
	{8'd116,8'd26} : s = 142;
	{8'd116,8'd27} : s = 143;
	{8'd116,8'd28} : s = 144;
	{8'd116,8'd29} : s = 145;
	{8'd116,8'd30} : s = 146;
	{8'd116,8'd31} : s = 147;
	{8'd116,8'd32} : s = 148;
	{8'd116,8'd33} : s = 149;
	{8'd116,8'd34} : s = 150;
	{8'd116,8'd35} : s = 151;
	{8'd116,8'd36} : s = 152;
	{8'd116,8'd37} : s = 153;
	{8'd116,8'd38} : s = 154;
	{8'd116,8'd39} : s = 155;
	{8'd116,8'd40} : s = 156;
	{8'd116,8'd41} : s = 157;
	{8'd116,8'd42} : s = 158;
	{8'd116,8'd43} : s = 159;
	{8'd116,8'd44} : s = 160;
	{8'd116,8'd45} : s = 161;
	{8'd116,8'd46} : s = 162;
	{8'd116,8'd47} : s = 163;
	{8'd116,8'd48} : s = 164;
	{8'd116,8'd49} : s = 165;
	{8'd116,8'd50} : s = 166;
	{8'd116,8'd51} : s = 167;
	{8'd116,8'd52} : s = 168;
	{8'd116,8'd53} : s = 169;
	{8'd116,8'd54} : s = 170;
	{8'd116,8'd55} : s = 171;
	{8'd116,8'd56} : s = 172;
	{8'd116,8'd57} : s = 173;
	{8'd116,8'd58} : s = 174;
	{8'd116,8'd59} : s = 175;
	{8'd116,8'd60} : s = 176;
	{8'd116,8'd61} : s = 177;
	{8'd116,8'd62} : s = 178;
	{8'd116,8'd63} : s = 179;
	{8'd116,8'd64} : s = 180;
	{8'd116,8'd65} : s = 181;
	{8'd116,8'd66} : s = 182;
	{8'd116,8'd67} : s = 183;
	{8'd116,8'd68} : s = 184;
	{8'd116,8'd69} : s = 185;
	{8'd116,8'd70} : s = 186;
	{8'd116,8'd71} : s = 187;
	{8'd116,8'd72} : s = 188;
	{8'd116,8'd73} : s = 189;
	{8'd116,8'd74} : s = 190;
	{8'd116,8'd75} : s = 191;
	{8'd116,8'd76} : s = 192;
	{8'd116,8'd77} : s = 193;
	{8'd116,8'd78} : s = 194;
	{8'd116,8'd79} : s = 195;
	{8'd116,8'd80} : s = 196;
	{8'd116,8'd81} : s = 197;
	{8'd116,8'd82} : s = 198;
	{8'd116,8'd83} : s = 199;
	{8'd116,8'd84} : s = 200;
	{8'd116,8'd85} : s = 201;
	{8'd116,8'd86} : s = 202;
	{8'd116,8'd87} : s = 203;
	{8'd116,8'd88} : s = 204;
	{8'd116,8'd89} : s = 205;
	{8'd116,8'd90} : s = 206;
	{8'd116,8'd91} : s = 207;
	{8'd116,8'd92} : s = 208;
	{8'd116,8'd93} : s = 209;
	{8'd116,8'd94} : s = 210;
	{8'd116,8'd95} : s = 211;
	{8'd116,8'd96} : s = 212;
	{8'd116,8'd97} : s = 213;
	{8'd116,8'd98} : s = 214;
	{8'd116,8'd99} : s = 215;
	{8'd116,8'd100} : s = 216;
	{8'd116,8'd101} : s = 217;
	{8'd116,8'd102} : s = 218;
	{8'd116,8'd103} : s = 219;
	{8'd116,8'd104} : s = 220;
	{8'd116,8'd105} : s = 221;
	{8'd116,8'd106} : s = 222;
	{8'd116,8'd107} : s = 223;
	{8'd116,8'd108} : s = 224;
	{8'd116,8'd109} : s = 225;
	{8'd116,8'd110} : s = 226;
	{8'd116,8'd111} : s = 227;
	{8'd116,8'd112} : s = 228;
	{8'd116,8'd113} : s = 229;
	{8'd116,8'd114} : s = 230;
	{8'd116,8'd115} : s = 231;
	{8'd116,8'd116} : s = 232;
	{8'd116,8'd117} : s = 233;
	{8'd116,8'd118} : s = 234;
	{8'd116,8'd119} : s = 235;
	{8'd116,8'd120} : s = 236;
	{8'd116,8'd121} : s = 237;
	{8'd116,8'd122} : s = 238;
	{8'd116,8'd123} : s = 239;
	{8'd116,8'd124} : s = 240;
	{8'd116,8'd125} : s = 241;
	{8'd116,8'd126} : s = 242;
	{8'd116,8'd127} : s = 243;
	{8'd116,8'd128} : s = 244;
	{8'd116,8'd129} : s = 245;
	{8'd116,8'd130} : s = 246;
	{8'd116,8'd131} : s = 247;
	{8'd116,8'd132} : s = 248;
	{8'd116,8'd133} : s = 249;
	{8'd116,8'd134} : s = 250;
	{8'd116,8'd135} : s = 251;
	{8'd116,8'd136} : s = 252;
	{8'd116,8'd137} : s = 253;
	{8'd116,8'd138} : s = 254;
	{8'd116,8'd139} : s = 255;
	{8'd116,8'd140} : s = 256;
	{8'd116,8'd141} : s = 257;
	{8'd116,8'd142} : s = 258;
	{8'd116,8'd143} : s = 259;
	{8'd116,8'd144} : s = 260;
	{8'd116,8'd145} : s = 261;
	{8'd116,8'd146} : s = 262;
	{8'd116,8'd147} : s = 263;
	{8'd116,8'd148} : s = 264;
	{8'd116,8'd149} : s = 265;
	{8'd116,8'd150} : s = 266;
	{8'd116,8'd151} : s = 267;
	{8'd116,8'd152} : s = 268;
	{8'd116,8'd153} : s = 269;
	{8'd116,8'd154} : s = 270;
	{8'd116,8'd155} : s = 271;
	{8'd116,8'd156} : s = 272;
	{8'd116,8'd157} : s = 273;
	{8'd116,8'd158} : s = 274;
	{8'd116,8'd159} : s = 275;
	{8'd116,8'd160} : s = 276;
	{8'd116,8'd161} : s = 277;
	{8'd116,8'd162} : s = 278;
	{8'd116,8'd163} : s = 279;
	{8'd116,8'd164} : s = 280;
	{8'd116,8'd165} : s = 281;
	{8'd116,8'd166} : s = 282;
	{8'd116,8'd167} : s = 283;
	{8'd116,8'd168} : s = 284;
	{8'd116,8'd169} : s = 285;
	{8'd116,8'd170} : s = 286;
	{8'd116,8'd171} : s = 287;
	{8'd116,8'd172} : s = 288;
	{8'd116,8'd173} : s = 289;
	{8'd116,8'd174} : s = 290;
	{8'd116,8'd175} : s = 291;
	{8'd116,8'd176} : s = 292;
	{8'd116,8'd177} : s = 293;
	{8'd116,8'd178} : s = 294;
	{8'd116,8'd179} : s = 295;
	{8'd116,8'd180} : s = 296;
	{8'd116,8'd181} : s = 297;
	{8'd116,8'd182} : s = 298;
	{8'd116,8'd183} : s = 299;
	{8'd116,8'd184} : s = 300;
	{8'd116,8'd185} : s = 301;
	{8'd116,8'd186} : s = 302;
	{8'd116,8'd187} : s = 303;
	{8'd116,8'd188} : s = 304;
	{8'd116,8'd189} : s = 305;
	{8'd116,8'd190} : s = 306;
	{8'd116,8'd191} : s = 307;
	{8'd116,8'd192} : s = 308;
	{8'd116,8'd193} : s = 309;
	{8'd116,8'd194} : s = 310;
	{8'd116,8'd195} : s = 311;
	{8'd116,8'd196} : s = 312;
	{8'd116,8'd197} : s = 313;
	{8'd116,8'd198} : s = 314;
	{8'd116,8'd199} : s = 315;
	{8'd116,8'd200} : s = 316;
	{8'd116,8'd201} : s = 317;
	{8'd116,8'd202} : s = 318;
	{8'd116,8'd203} : s = 319;
	{8'd116,8'd204} : s = 320;
	{8'd116,8'd205} : s = 321;
	{8'd116,8'd206} : s = 322;
	{8'd116,8'd207} : s = 323;
	{8'd116,8'd208} : s = 324;
	{8'd116,8'd209} : s = 325;
	{8'd116,8'd210} : s = 326;
	{8'd116,8'd211} : s = 327;
	{8'd116,8'd212} : s = 328;
	{8'd116,8'd213} : s = 329;
	{8'd116,8'd214} : s = 330;
	{8'd116,8'd215} : s = 331;
	{8'd116,8'd216} : s = 332;
	{8'd116,8'd217} : s = 333;
	{8'd116,8'd218} : s = 334;
	{8'd116,8'd219} : s = 335;
	{8'd116,8'd220} : s = 336;
	{8'd116,8'd221} : s = 337;
	{8'd116,8'd222} : s = 338;
	{8'd116,8'd223} : s = 339;
	{8'd116,8'd224} : s = 340;
	{8'd116,8'd225} : s = 341;
	{8'd116,8'd226} : s = 342;
	{8'd116,8'd227} : s = 343;
	{8'd116,8'd228} : s = 344;
	{8'd116,8'd229} : s = 345;
	{8'd116,8'd230} : s = 346;
	{8'd116,8'd231} : s = 347;
	{8'd116,8'd232} : s = 348;
	{8'd116,8'd233} : s = 349;
	{8'd116,8'd234} : s = 350;
	{8'd116,8'd235} : s = 351;
	{8'd116,8'd236} : s = 352;
	{8'd116,8'd237} : s = 353;
	{8'd116,8'd238} : s = 354;
	{8'd116,8'd239} : s = 355;
	{8'd116,8'd240} : s = 356;
	{8'd116,8'd241} : s = 357;
	{8'd116,8'd242} : s = 358;
	{8'd116,8'd243} : s = 359;
	{8'd116,8'd244} : s = 360;
	{8'd116,8'd245} : s = 361;
	{8'd116,8'd246} : s = 362;
	{8'd116,8'd247} : s = 363;
	{8'd116,8'd248} : s = 364;
	{8'd116,8'd249} : s = 365;
	{8'd116,8'd250} : s = 366;
	{8'd116,8'd251} : s = 367;
	{8'd116,8'd252} : s = 368;
	{8'd116,8'd253} : s = 369;
	{8'd116,8'd254} : s = 370;
	{8'd116,8'd255} : s = 371;
	{8'd117,8'd0} : s = 117;
	{8'd117,8'd1} : s = 118;
	{8'd117,8'd2} : s = 119;
	{8'd117,8'd3} : s = 120;
	{8'd117,8'd4} : s = 121;
	{8'd117,8'd5} : s = 122;
	{8'd117,8'd6} : s = 123;
	{8'd117,8'd7} : s = 124;
	{8'd117,8'd8} : s = 125;
	{8'd117,8'd9} : s = 126;
	{8'd117,8'd10} : s = 127;
	{8'd117,8'd11} : s = 128;
	{8'd117,8'd12} : s = 129;
	{8'd117,8'd13} : s = 130;
	{8'd117,8'd14} : s = 131;
	{8'd117,8'd15} : s = 132;
	{8'd117,8'd16} : s = 133;
	{8'd117,8'd17} : s = 134;
	{8'd117,8'd18} : s = 135;
	{8'd117,8'd19} : s = 136;
	{8'd117,8'd20} : s = 137;
	{8'd117,8'd21} : s = 138;
	{8'd117,8'd22} : s = 139;
	{8'd117,8'd23} : s = 140;
	{8'd117,8'd24} : s = 141;
	{8'd117,8'd25} : s = 142;
	{8'd117,8'd26} : s = 143;
	{8'd117,8'd27} : s = 144;
	{8'd117,8'd28} : s = 145;
	{8'd117,8'd29} : s = 146;
	{8'd117,8'd30} : s = 147;
	{8'd117,8'd31} : s = 148;
	{8'd117,8'd32} : s = 149;
	{8'd117,8'd33} : s = 150;
	{8'd117,8'd34} : s = 151;
	{8'd117,8'd35} : s = 152;
	{8'd117,8'd36} : s = 153;
	{8'd117,8'd37} : s = 154;
	{8'd117,8'd38} : s = 155;
	{8'd117,8'd39} : s = 156;
	{8'd117,8'd40} : s = 157;
	{8'd117,8'd41} : s = 158;
	{8'd117,8'd42} : s = 159;
	{8'd117,8'd43} : s = 160;
	{8'd117,8'd44} : s = 161;
	{8'd117,8'd45} : s = 162;
	{8'd117,8'd46} : s = 163;
	{8'd117,8'd47} : s = 164;
	{8'd117,8'd48} : s = 165;
	{8'd117,8'd49} : s = 166;
	{8'd117,8'd50} : s = 167;
	{8'd117,8'd51} : s = 168;
	{8'd117,8'd52} : s = 169;
	{8'd117,8'd53} : s = 170;
	{8'd117,8'd54} : s = 171;
	{8'd117,8'd55} : s = 172;
	{8'd117,8'd56} : s = 173;
	{8'd117,8'd57} : s = 174;
	{8'd117,8'd58} : s = 175;
	{8'd117,8'd59} : s = 176;
	{8'd117,8'd60} : s = 177;
	{8'd117,8'd61} : s = 178;
	{8'd117,8'd62} : s = 179;
	{8'd117,8'd63} : s = 180;
	{8'd117,8'd64} : s = 181;
	{8'd117,8'd65} : s = 182;
	{8'd117,8'd66} : s = 183;
	{8'd117,8'd67} : s = 184;
	{8'd117,8'd68} : s = 185;
	{8'd117,8'd69} : s = 186;
	{8'd117,8'd70} : s = 187;
	{8'd117,8'd71} : s = 188;
	{8'd117,8'd72} : s = 189;
	{8'd117,8'd73} : s = 190;
	{8'd117,8'd74} : s = 191;
	{8'd117,8'd75} : s = 192;
	{8'd117,8'd76} : s = 193;
	{8'd117,8'd77} : s = 194;
	{8'd117,8'd78} : s = 195;
	{8'd117,8'd79} : s = 196;
	{8'd117,8'd80} : s = 197;
	{8'd117,8'd81} : s = 198;
	{8'd117,8'd82} : s = 199;
	{8'd117,8'd83} : s = 200;
	{8'd117,8'd84} : s = 201;
	{8'd117,8'd85} : s = 202;
	{8'd117,8'd86} : s = 203;
	{8'd117,8'd87} : s = 204;
	{8'd117,8'd88} : s = 205;
	{8'd117,8'd89} : s = 206;
	{8'd117,8'd90} : s = 207;
	{8'd117,8'd91} : s = 208;
	{8'd117,8'd92} : s = 209;
	{8'd117,8'd93} : s = 210;
	{8'd117,8'd94} : s = 211;
	{8'd117,8'd95} : s = 212;
	{8'd117,8'd96} : s = 213;
	{8'd117,8'd97} : s = 214;
	{8'd117,8'd98} : s = 215;
	{8'd117,8'd99} : s = 216;
	{8'd117,8'd100} : s = 217;
	{8'd117,8'd101} : s = 218;
	{8'd117,8'd102} : s = 219;
	{8'd117,8'd103} : s = 220;
	{8'd117,8'd104} : s = 221;
	{8'd117,8'd105} : s = 222;
	{8'd117,8'd106} : s = 223;
	{8'd117,8'd107} : s = 224;
	{8'd117,8'd108} : s = 225;
	{8'd117,8'd109} : s = 226;
	{8'd117,8'd110} : s = 227;
	{8'd117,8'd111} : s = 228;
	{8'd117,8'd112} : s = 229;
	{8'd117,8'd113} : s = 230;
	{8'd117,8'd114} : s = 231;
	{8'd117,8'd115} : s = 232;
	{8'd117,8'd116} : s = 233;
	{8'd117,8'd117} : s = 234;
	{8'd117,8'd118} : s = 235;
	{8'd117,8'd119} : s = 236;
	{8'd117,8'd120} : s = 237;
	{8'd117,8'd121} : s = 238;
	{8'd117,8'd122} : s = 239;
	{8'd117,8'd123} : s = 240;
	{8'd117,8'd124} : s = 241;
	{8'd117,8'd125} : s = 242;
	{8'd117,8'd126} : s = 243;
	{8'd117,8'd127} : s = 244;
	{8'd117,8'd128} : s = 245;
	{8'd117,8'd129} : s = 246;
	{8'd117,8'd130} : s = 247;
	{8'd117,8'd131} : s = 248;
	{8'd117,8'd132} : s = 249;
	{8'd117,8'd133} : s = 250;
	{8'd117,8'd134} : s = 251;
	{8'd117,8'd135} : s = 252;
	{8'd117,8'd136} : s = 253;
	{8'd117,8'd137} : s = 254;
	{8'd117,8'd138} : s = 255;
	{8'd117,8'd139} : s = 256;
	{8'd117,8'd140} : s = 257;
	{8'd117,8'd141} : s = 258;
	{8'd117,8'd142} : s = 259;
	{8'd117,8'd143} : s = 260;
	{8'd117,8'd144} : s = 261;
	{8'd117,8'd145} : s = 262;
	{8'd117,8'd146} : s = 263;
	{8'd117,8'd147} : s = 264;
	{8'd117,8'd148} : s = 265;
	{8'd117,8'd149} : s = 266;
	{8'd117,8'd150} : s = 267;
	{8'd117,8'd151} : s = 268;
	{8'd117,8'd152} : s = 269;
	{8'd117,8'd153} : s = 270;
	{8'd117,8'd154} : s = 271;
	{8'd117,8'd155} : s = 272;
	{8'd117,8'd156} : s = 273;
	{8'd117,8'd157} : s = 274;
	{8'd117,8'd158} : s = 275;
	{8'd117,8'd159} : s = 276;
	{8'd117,8'd160} : s = 277;
	{8'd117,8'd161} : s = 278;
	{8'd117,8'd162} : s = 279;
	{8'd117,8'd163} : s = 280;
	{8'd117,8'd164} : s = 281;
	{8'd117,8'd165} : s = 282;
	{8'd117,8'd166} : s = 283;
	{8'd117,8'd167} : s = 284;
	{8'd117,8'd168} : s = 285;
	{8'd117,8'd169} : s = 286;
	{8'd117,8'd170} : s = 287;
	{8'd117,8'd171} : s = 288;
	{8'd117,8'd172} : s = 289;
	{8'd117,8'd173} : s = 290;
	{8'd117,8'd174} : s = 291;
	{8'd117,8'd175} : s = 292;
	{8'd117,8'd176} : s = 293;
	{8'd117,8'd177} : s = 294;
	{8'd117,8'd178} : s = 295;
	{8'd117,8'd179} : s = 296;
	{8'd117,8'd180} : s = 297;
	{8'd117,8'd181} : s = 298;
	{8'd117,8'd182} : s = 299;
	{8'd117,8'd183} : s = 300;
	{8'd117,8'd184} : s = 301;
	{8'd117,8'd185} : s = 302;
	{8'd117,8'd186} : s = 303;
	{8'd117,8'd187} : s = 304;
	{8'd117,8'd188} : s = 305;
	{8'd117,8'd189} : s = 306;
	{8'd117,8'd190} : s = 307;
	{8'd117,8'd191} : s = 308;
	{8'd117,8'd192} : s = 309;
	{8'd117,8'd193} : s = 310;
	{8'd117,8'd194} : s = 311;
	{8'd117,8'd195} : s = 312;
	{8'd117,8'd196} : s = 313;
	{8'd117,8'd197} : s = 314;
	{8'd117,8'd198} : s = 315;
	{8'd117,8'd199} : s = 316;
	{8'd117,8'd200} : s = 317;
	{8'd117,8'd201} : s = 318;
	{8'd117,8'd202} : s = 319;
	{8'd117,8'd203} : s = 320;
	{8'd117,8'd204} : s = 321;
	{8'd117,8'd205} : s = 322;
	{8'd117,8'd206} : s = 323;
	{8'd117,8'd207} : s = 324;
	{8'd117,8'd208} : s = 325;
	{8'd117,8'd209} : s = 326;
	{8'd117,8'd210} : s = 327;
	{8'd117,8'd211} : s = 328;
	{8'd117,8'd212} : s = 329;
	{8'd117,8'd213} : s = 330;
	{8'd117,8'd214} : s = 331;
	{8'd117,8'd215} : s = 332;
	{8'd117,8'd216} : s = 333;
	{8'd117,8'd217} : s = 334;
	{8'd117,8'd218} : s = 335;
	{8'd117,8'd219} : s = 336;
	{8'd117,8'd220} : s = 337;
	{8'd117,8'd221} : s = 338;
	{8'd117,8'd222} : s = 339;
	{8'd117,8'd223} : s = 340;
	{8'd117,8'd224} : s = 341;
	{8'd117,8'd225} : s = 342;
	{8'd117,8'd226} : s = 343;
	{8'd117,8'd227} : s = 344;
	{8'd117,8'd228} : s = 345;
	{8'd117,8'd229} : s = 346;
	{8'd117,8'd230} : s = 347;
	{8'd117,8'd231} : s = 348;
	{8'd117,8'd232} : s = 349;
	{8'd117,8'd233} : s = 350;
	{8'd117,8'd234} : s = 351;
	{8'd117,8'd235} : s = 352;
	{8'd117,8'd236} : s = 353;
	{8'd117,8'd237} : s = 354;
	{8'd117,8'd238} : s = 355;
	{8'd117,8'd239} : s = 356;
	{8'd117,8'd240} : s = 357;
	{8'd117,8'd241} : s = 358;
	{8'd117,8'd242} : s = 359;
	{8'd117,8'd243} : s = 360;
	{8'd117,8'd244} : s = 361;
	{8'd117,8'd245} : s = 362;
	{8'd117,8'd246} : s = 363;
	{8'd117,8'd247} : s = 364;
	{8'd117,8'd248} : s = 365;
	{8'd117,8'd249} : s = 366;
	{8'd117,8'd250} : s = 367;
	{8'd117,8'd251} : s = 368;
	{8'd117,8'd252} : s = 369;
	{8'd117,8'd253} : s = 370;
	{8'd117,8'd254} : s = 371;
	{8'd117,8'd255} : s = 372;
	{8'd118,8'd0} : s = 118;
	{8'd118,8'd1} : s = 119;
	{8'd118,8'd2} : s = 120;
	{8'd118,8'd3} : s = 121;
	{8'd118,8'd4} : s = 122;
	{8'd118,8'd5} : s = 123;
	{8'd118,8'd6} : s = 124;
	{8'd118,8'd7} : s = 125;
	{8'd118,8'd8} : s = 126;
	{8'd118,8'd9} : s = 127;
	{8'd118,8'd10} : s = 128;
	{8'd118,8'd11} : s = 129;
	{8'd118,8'd12} : s = 130;
	{8'd118,8'd13} : s = 131;
	{8'd118,8'd14} : s = 132;
	{8'd118,8'd15} : s = 133;
	{8'd118,8'd16} : s = 134;
	{8'd118,8'd17} : s = 135;
	{8'd118,8'd18} : s = 136;
	{8'd118,8'd19} : s = 137;
	{8'd118,8'd20} : s = 138;
	{8'd118,8'd21} : s = 139;
	{8'd118,8'd22} : s = 140;
	{8'd118,8'd23} : s = 141;
	{8'd118,8'd24} : s = 142;
	{8'd118,8'd25} : s = 143;
	{8'd118,8'd26} : s = 144;
	{8'd118,8'd27} : s = 145;
	{8'd118,8'd28} : s = 146;
	{8'd118,8'd29} : s = 147;
	{8'd118,8'd30} : s = 148;
	{8'd118,8'd31} : s = 149;
	{8'd118,8'd32} : s = 150;
	{8'd118,8'd33} : s = 151;
	{8'd118,8'd34} : s = 152;
	{8'd118,8'd35} : s = 153;
	{8'd118,8'd36} : s = 154;
	{8'd118,8'd37} : s = 155;
	{8'd118,8'd38} : s = 156;
	{8'd118,8'd39} : s = 157;
	{8'd118,8'd40} : s = 158;
	{8'd118,8'd41} : s = 159;
	{8'd118,8'd42} : s = 160;
	{8'd118,8'd43} : s = 161;
	{8'd118,8'd44} : s = 162;
	{8'd118,8'd45} : s = 163;
	{8'd118,8'd46} : s = 164;
	{8'd118,8'd47} : s = 165;
	{8'd118,8'd48} : s = 166;
	{8'd118,8'd49} : s = 167;
	{8'd118,8'd50} : s = 168;
	{8'd118,8'd51} : s = 169;
	{8'd118,8'd52} : s = 170;
	{8'd118,8'd53} : s = 171;
	{8'd118,8'd54} : s = 172;
	{8'd118,8'd55} : s = 173;
	{8'd118,8'd56} : s = 174;
	{8'd118,8'd57} : s = 175;
	{8'd118,8'd58} : s = 176;
	{8'd118,8'd59} : s = 177;
	{8'd118,8'd60} : s = 178;
	{8'd118,8'd61} : s = 179;
	{8'd118,8'd62} : s = 180;
	{8'd118,8'd63} : s = 181;
	{8'd118,8'd64} : s = 182;
	{8'd118,8'd65} : s = 183;
	{8'd118,8'd66} : s = 184;
	{8'd118,8'd67} : s = 185;
	{8'd118,8'd68} : s = 186;
	{8'd118,8'd69} : s = 187;
	{8'd118,8'd70} : s = 188;
	{8'd118,8'd71} : s = 189;
	{8'd118,8'd72} : s = 190;
	{8'd118,8'd73} : s = 191;
	{8'd118,8'd74} : s = 192;
	{8'd118,8'd75} : s = 193;
	{8'd118,8'd76} : s = 194;
	{8'd118,8'd77} : s = 195;
	{8'd118,8'd78} : s = 196;
	{8'd118,8'd79} : s = 197;
	{8'd118,8'd80} : s = 198;
	{8'd118,8'd81} : s = 199;
	{8'd118,8'd82} : s = 200;
	{8'd118,8'd83} : s = 201;
	{8'd118,8'd84} : s = 202;
	{8'd118,8'd85} : s = 203;
	{8'd118,8'd86} : s = 204;
	{8'd118,8'd87} : s = 205;
	{8'd118,8'd88} : s = 206;
	{8'd118,8'd89} : s = 207;
	{8'd118,8'd90} : s = 208;
	{8'd118,8'd91} : s = 209;
	{8'd118,8'd92} : s = 210;
	{8'd118,8'd93} : s = 211;
	{8'd118,8'd94} : s = 212;
	{8'd118,8'd95} : s = 213;
	{8'd118,8'd96} : s = 214;
	{8'd118,8'd97} : s = 215;
	{8'd118,8'd98} : s = 216;
	{8'd118,8'd99} : s = 217;
	{8'd118,8'd100} : s = 218;
	{8'd118,8'd101} : s = 219;
	{8'd118,8'd102} : s = 220;
	{8'd118,8'd103} : s = 221;
	{8'd118,8'd104} : s = 222;
	{8'd118,8'd105} : s = 223;
	{8'd118,8'd106} : s = 224;
	{8'd118,8'd107} : s = 225;
	{8'd118,8'd108} : s = 226;
	{8'd118,8'd109} : s = 227;
	{8'd118,8'd110} : s = 228;
	{8'd118,8'd111} : s = 229;
	{8'd118,8'd112} : s = 230;
	{8'd118,8'd113} : s = 231;
	{8'd118,8'd114} : s = 232;
	{8'd118,8'd115} : s = 233;
	{8'd118,8'd116} : s = 234;
	{8'd118,8'd117} : s = 235;
	{8'd118,8'd118} : s = 236;
	{8'd118,8'd119} : s = 237;
	{8'd118,8'd120} : s = 238;
	{8'd118,8'd121} : s = 239;
	{8'd118,8'd122} : s = 240;
	{8'd118,8'd123} : s = 241;
	{8'd118,8'd124} : s = 242;
	{8'd118,8'd125} : s = 243;
	{8'd118,8'd126} : s = 244;
	{8'd118,8'd127} : s = 245;
	{8'd118,8'd128} : s = 246;
	{8'd118,8'd129} : s = 247;
	{8'd118,8'd130} : s = 248;
	{8'd118,8'd131} : s = 249;
	{8'd118,8'd132} : s = 250;
	{8'd118,8'd133} : s = 251;
	{8'd118,8'd134} : s = 252;
	{8'd118,8'd135} : s = 253;
	{8'd118,8'd136} : s = 254;
	{8'd118,8'd137} : s = 255;
	{8'd118,8'd138} : s = 256;
	{8'd118,8'd139} : s = 257;
	{8'd118,8'd140} : s = 258;
	{8'd118,8'd141} : s = 259;
	{8'd118,8'd142} : s = 260;
	{8'd118,8'd143} : s = 261;
	{8'd118,8'd144} : s = 262;
	{8'd118,8'd145} : s = 263;
	{8'd118,8'd146} : s = 264;
	{8'd118,8'd147} : s = 265;
	{8'd118,8'd148} : s = 266;
	{8'd118,8'd149} : s = 267;
	{8'd118,8'd150} : s = 268;
	{8'd118,8'd151} : s = 269;
	{8'd118,8'd152} : s = 270;
	{8'd118,8'd153} : s = 271;
	{8'd118,8'd154} : s = 272;
	{8'd118,8'd155} : s = 273;
	{8'd118,8'd156} : s = 274;
	{8'd118,8'd157} : s = 275;
	{8'd118,8'd158} : s = 276;
	{8'd118,8'd159} : s = 277;
	{8'd118,8'd160} : s = 278;
	{8'd118,8'd161} : s = 279;
	{8'd118,8'd162} : s = 280;
	{8'd118,8'd163} : s = 281;
	{8'd118,8'd164} : s = 282;
	{8'd118,8'd165} : s = 283;
	{8'd118,8'd166} : s = 284;
	{8'd118,8'd167} : s = 285;
	{8'd118,8'd168} : s = 286;
	{8'd118,8'd169} : s = 287;
	{8'd118,8'd170} : s = 288;
	{8'd118,8'd171} : s = 289;
	{8'd118,8'd172} : s = 290;
	{8'd118,8'd173} : s = 291;
	{8'd118,8'd174} : s = 292;
	{8'd118,8'd175} : s = 293;
	{8'd118,8'd176} : s = 294;
	{8'd118,8'd177} : s = 295;
	{8'd118,8'd178} : s = 296;
	{8'd118,8'd179} : s = 297;
	{8'd118,8'd180} : s = 298;
	{8'd118,8'd181} : s = 299;
	{8'd118,8'd182} : s = 300;
	{8'd118,8'd183} : s = 301;
	{8'd118,8'd184} : s = 302;
	{8'd118,8'd185} : s = 303;
	{8'd118,8'd186} : s = 304;
	{8'd118,8'd187} : s = 305;
	{8'd118,8'd188} : s = 306;
	{8'd118,8'd189} : s = 307;
	{8'd118,8'd190} : s = 308;
	{8'd118,8'd191} : s = 309;
	{8'd118,8'd192} : s = 310;
	{8'd118,8'd193} : s = 311;
	{8'd118,8'd194} : s = 312;
	{8'd118,8'd195} : s = 313;
	{8'd118,8'd196} : s = 314;
	{8'd118,8'd197} : s = 315;
	{8'd118,8'd198} : s = 316;
	{8'd118,8'd199} : s = 317;
	{8'd118,8'd200} : s = 318;
	{8'd118,8'd201} : s = 319;
	{8'd118,8'd202} : s = 320;
	{8'd118,8'd203} : s = 321;
	{8'd118,8'd204} : s = 322;
	{8'd118,8'd205} : s = 323;
	{8'd118,8'd206} : s = 324;
	{8'd118,8'd207} : s = 325;
	{8'd118,8'd208} : s = 326;
	{8'd118,8'd209} : s = 327;
	{8'd118,8'd210} : s = 328;
	{8'd118,8'd211} : s = 329;
	{8'd118,8'd212} : s = 330;
	{8'd118,8'd213} : s = 331;
	{8'd118,8'd214} : s = 332;
	{8'd118,8'd215} : s = 333;
	{8'd118,8'd216} : s = 334;
	{8'd118,8'd217} : s = 335;
	{8'd118,8'd218} : s = 336;
	{8'd118,8'd219} : s = 337;
	{8'd118,8'd220} : s = 338;
	{8'd118,8'd221} : s = 339;
	{8'd118,8'd222} : s = 340;
	{8'd118,8'd223} : s = 341;
	{8'd118,8'd224} : s = 342;
	{8'd118,8'd225} : s = 343;
	{8'd118,8'd226} : s = 344;
	{8'd118,8'd227} : s = 345;
	{8'd118,8'd228} : s = 346;
	{8'd118,8'd229} : s = 347;
	{8'd118,8'd230} : s = 348;
	{8'd118,8'd231} : s = 349;
	{8'd118,8'd232} : s = 350;
	{8'd118,8'd233} : s = 351;
	{8'd118,8'd234} : s = 352;
	{8'd118,8'd235} : s = 353;
	{8'd118,8'd236} : s = 354;
	{8'd118,8'd237} : s = 355;
	{8'd118,8'd238} : s = 356;
	{8'd118,8'd239} : s = 357;
	{8'd118,8'd240} : s = 358;
	{8'd118,8'd241} : s = 359;
	{8'd118,8'd242} : s = 360;
	{8'd118,8'd243} : s = 361;
	{8'd118,8'd244} : s = 362;
	{8'd118,8'd245} : s = 363;
	{8'd118,8'd246} : s = 364;
	{8'd118,8'd247} : s = 365;
	{8'd118,8'd248} : s = 366;
	{8'd118,8'd249} : s = 367;
	{8'd118,8'd250} : s = 368;
	{8'd118,8'd251} : s = 369;
	{8'd118,8'd252} : s = 370;
	{8'd118,8'd253} : s = 371;
	{8'd118,8'd254} : s = 372;
	{8'd118,8'd255} : s = 373;
	{8'd119,8'd0} : s = 119;
	{8'd119,8'd1} : s = 120;
	{8'd119,8'd2} : s = 121;
	{8'd119,8'd3} : s = 122;
	{8'd119,8'd4} : s = 123;
	{8'd119,8'd5} : s = 124;
	{8'd119,8'd6} : s = 125;
	{8'd119,8'd7} : s = 126;
	{8'd119,8'd8} : s = 127;
	{8'd119,8'd9} : s = 128;
	{8'd119,8'd10} : s = 129;
	{8'd119,8'd11} : s = 130;
	{8'd119,8'd12} : s = 131;
	{8'd119,8'd13} : s = 132;
	{8'd119,8'd14} : s = 133;
	{8'd119,8'd15} : s = 134;
	{8'd119,8'd16} : s = 135;
	{8'd119,8'd17} : s = 136;
	{8'd119,8'd18} : s = 137;
	{8'd119,8'd19} : s = 138;
	{8'd119,8'd20} : s = 139;
	{8'd119,8'd21} : s = 140;
	{8'd119,8'd22} : s = 141;
	{8'd119,8'd23} : s = 142;
	{8'd119,8'd24} : s = 143;
	{8'd119,8'd25} : s = 144;
	{8'd119,8'd26} : s = 145;
	{8'd119,8'd27} : s = 146;
	{8'd119,8'd28} : s = 147;
	{8'd119,8'd29} : s = 148;
	{8'd119,8'd30} : s = 149;
	{8'd119,8'd31} : s = 150;
	{8'd119,8'd32} : s = 151;
	{8'd119,8'd33} : s = 152;
	{8'd119,8'd34} : s = 153;
	{8'd119,8'd35} : s = 154;
	{8'd119,8'd36} : s = 155;
	{8'd119,8'd37} : s = 156;
	{8'd119,8'd38} : s = 157;
	{8'd119,8'd39} : s = 158;
	{8'd119,8'd40} : s = 159;
	{8'd119,8'd41} : s = 160;
	{8'd119,8'd42} : s = 161;
	{8'd119,8'd43} : s = 162;
	{8'd119,8'd44} : s = 163;
	{8'd119,8'd45} : s = 164;
	{8'd119,8'd46} : s = 165;
	{8'd119,8'd47} : s = 166;
	{8'd119,8'd48} : s = 167;
	{8'd119,8'd49} : s = 168;
	{8'd119,8'd50} : s = 169;
	{8'd119,8'd51} : s = 170;
	{8'd119,8'd52} : s = 171;
	{8'd119,8'd53} : s = 172;
	{8'd119,8'd54} : s = 173;
	{8'd119,8'd55} : s = 174;
	{8'd119,8'd56} : s = 175;
	{8'd119,8'd57} : s = 176;
	{8'd119,8'd58} : s = 177;
	{8'd119,8'd59} : s = 178;
	{8'd119,8'd60} : s = 179;
	{8'd119,8'd61} : s = 180;
	{8'd119,8'd62} : s = 181;
	{8'd119,8'd63} : s = 182;
	{8'd119,8'd64} : s = 183;
	{8'd119,8'd65} : s = 184;
	{8'd119,8'd66} : s = 185;
	{8'd119,8'd67} : s = 186;
	{8'd119,8'd68} : s = 187;
	{8'd119,8'd69} : s = 188;
	{8'd119,8'd70} : s = 189;
	{8'd119,8'd71} : s = 190;
	{8'd119,8'd72} : s = 191;
	{8'd119,8'd73} : s = 192;
	{8'd119,8'd74} : s = 193;
	{8'd119,8'd75} : s = 194;
	{8'd119,8'd76} : s = 195;
	{8'd119,8'd77} : s = 196;
	{8'd119,8'd78} : s = 197;
	{8'd119,8'd79} : s = 198;
	{8'd119,8'd80} : s = 199;
	{8'd119,8'd81} : s = 200;
	{8'd119,8'd82} : s = 201;
	{8'd119,8'd83} : s = 202;
	{8'd119,8'd84} : s = 203;
	{8'd119,8'd85} : s = 204;
	{8'd119,8'd86} : s = 205;
	{8'd119,8'd87} : s = 206;
	{8'd119,8'd88} : s = 207;
	{8'd119,8'd89} : s = 208;
	{8'd119,8'd90} : s = 209;
	{8'd119,8'd91} : s = 210;
	{8'd119,8'd92} : s = 211;
	{8'd119,8'd93} : s = 212;
	{8'd119,8'd94} : s = 213;
	{8'd119,8'd95} : s = 214;
	{8'd119,8'd96} : s = 215;
	{8'd119,8'd97} : s = 216;
	{8'd119,8'd98} : s = 217;
	{8'd119,8'd99} : s = 218;
	{8'd119,8'd100} : s = 219;
	{8'd119,8'd101} : s = 220;
	{8'd119,8'd102} : s = 221;
	{8'd119,8'd103} : s = 222;
	{8'd119,8'd104} : s = 223;
	{8'd119,8'd105} : s = 224;
	{8'd119,8'd106} : s = 225;
	{8'd119,8'd107} : s = 226;
	{8'd119,8'd108} : s = 227;
	{8'd119,8'd109} : s = 228;
	{8'd119,8'd110} : s = 229;
	{8'd119,8'd111} : s = 230;
	{8'd119,8'd112} : s = 231;
	{8'd119,8'd113} : s = 232;
	{8'd119,8'd114} : s = 233;
	{8'd119,8'd115} : s = 234;
	{8'd119,8'd116} : s = 235;
	{8'd119,8'd117} : s = 236;
	{8'd119,8'd118} : s = 237;
	{8'd119,8'd119} : s = 238;
	{8'd119,8'd120} : s = 239;
	{8'd119,8'd121} : s = 240;
	{8'd119,8'd122} : s = 241;
	{8'd119,8'd123} : s = 242;
	{8'd119,8'd124} : s = 243;
	{8'd119,8'd125} : s = 244;
	{8'd119,8'd126} : s = 245;
	{8'd119,8'd127} : s = 246;
	{8'd119,8'd128} : s = 247;
	{8'd119,8'd129} : s = 248;
	{8'd119,8'd130} : s = 249;
	{8'd119,8'd131} : s = 250;
	{8'd119,8'd132} : s = 251;
	{8'd119,8'd133} : s = 252;
	{8'd119,8'd134} : s = 253;
	{8'd119,8'd135} : s = 254;
	{8'd119,8'd136} : s = 255;
	{8'd119,8'd137} : s = 256;
	{8'd119,8'd138} : s = 257;
	{8'd119,8'd139} : s = 258;
	{8'd119,8'd140} : s = 259;
	{8'd119,8'd141} : s = 260;
	{8'd119,8'd142} : s = 261;
	{8'd119,8'd143} : s = 262;
	{8'd119,8'd144} : s = 263;
	{8'd119,8'd145} : s = 264;
	{8'd119,8'd146} : s = 265;
	{8'd119,8'd147} : s = 266;
	{8'd119,8'd148} : s = 267;
	{8'd119,8'd149} : s = 268;
	{8'd119,8'd150} : s = 269;
	{8'd119,8'd151} : s = 270;
	{8'd119,8'd152} : s = 271;
	{8'd119,8'd153} : s = 272;
	{8'd119,8'd154} : s = 273;
	{8'd119,8'd155} : s = 274;
	{8'd119,8'd156} : s = 275;
	{8'd119,8'd157} : s = 276;
	{8'd119,8'd158} : s = 277;
	{8'd119,8'd159} : s = 278;
	{8'd119,8'd160} : s = 279;
	{8'd119,8'd161} : s = 280;
	{8'd119,8'd162} : s = 281;
	{8'd119,8'd163} : s = 282;
	{8'd119,8'd164} : s = 283;
	{8'd119,8'd165} : s = 284;
	{8'd119,8'd166} : s = 285;
	{8'd119,8'd167} : s = 286;
	{8'd119,8'd168} : s = 287;
	{8'd119,8'd169} : s = 288;
	{8'd119,8'd170} : s = 289;
	{8'd119,8'd171} : s = 290;
	{8'd119,8'd172} : s = 291;
	{8'd119,8'd173} : s = 292;
	{8'd119,8'd174} : s = 293;
	{8'd119,8'd175} : s = 294;
	{8'd119,8'd176} : s = 295;
	{8'd119,8'd177} : s = 296;
	{8'd119,8'd178} : s = 297;
	{8'd119,8'd179} : s = 298;
	{8'd119,8'd180} : s = 299;
	{8'd119,8'd181} : s = 300;
	{8'd119,8'd182} : s = 301;
	{8'd119,8'd183} : s = 302;
	{8'd119,8'd184} : s = 303;
	{8'd119,8'd185} : s = 304;
	{8'd119,8'd186} : s = 305;
	{8'd119,8'd187} : s = 306;
	{8'd119,8'd188} : s = 307;
	{8'd119,8'd189} : s = 308;
	{8'd119,8'd190} : s = 309;
	{8'd119,8'd191} : s = 310;
	{8'd119,8'd192} : s = 311;
	{8'd119,8'd193} : s = 312;
	{8'd119,8'd194} : s = 313;
	{8'd119,8'd195} : s = 314;
	{8'd119,8'd196} : s = 315;
	{8'd119,8'd197} : s = 316;
	{8'd119,8'd198} : s = 317;
	{8'd119,8'd199} : s = 318;
	{8'd119,8'd200} : s = 319;
	{8'd119,8'd201} : s = 320;
	{8'd119,8'd202} : s = 321;
	{8'd119,8'd203} : s = 322;
	{8'd119,8'd204} : s = 323;
	{8'd119,8'd205} : s = 324;
	{8'd119,8'd206} : s = 325;
	{8'd119,8'd207} : s = 326;
	{8'd119,8'd208} : s = 327;
	{8'd119,8'd209} : s = 328;
	{8'd119,8'd210} : s = 329;
	{8'd119,8'd211} : s = 330;
	{8'd119,8'd212} : s = 331;
	{8'd119,8'd213} : s = 332;
	{8'd119,8'd214} : s = 333;
	{8'd119,8'd215} : s = 334;
	{8'd119,8'd216} : s = 335;
	{8'd119,8'd217} : s = 336;
	{8'd119,8'd218} : s = 337;
	{8'd119,8'd219} : s = 338;
	{8'd119,8'd220} : s = 339;
	{8'd119,8'd221} : s = 340;
	{8'd119,8'd222} : s = 341;
	{8'd119,8'd223} : s = 342;
	{8'd119,8'd224} : s = 343;
	{8'd119,8'd225} : s = 344;
	{8'd119,8'd226} : s = 345;
	{8'd119,8'd227} : s = 346;
	{8'd119,8'd228} : s = 347;
	{8'd119,8'd229} : s = 348;
	{8'd119,8'd230} : s = 349;
	{8'd119,8'd231} : s = 350;
	{8'd119,8'd232} : s = 351;
	{8'd119,8'd233} : s = 352;
	{8'd119,8'd234} : s = 353;
	{8'd119,8'd235} : s = 354;
	{8'd119,8'd236} : s = 355;
	{8'd119,8'd237} : s = 356;
	{8'd119,8'd238} : s = 357;
	{8'd119,8'd239} : s = 358;
	{8'd119,8'd240} : s = 359;
	{8'd119,8'd241} : s = 360;
	{8'd119,8'd242} : s = 361;
	{8'd119,8'd243} : s = 362;
	{8'd119,8'd244} : s = 363;
	{8'd119,8'd245} : s = 364;
	{8'd119,8'd246} : s = 365;
	{8'd119,8'd247} : s = 366;
	{8'd119,8'd248} : s = 367;
	{8'd119,8'd249} : s = 368;
	{8'd119,8'd250} : s = 369;
	{8'd119,8'd251} : s = 370;
	{8'd119,8'd252} : s = 371;
	{8'd119,8'd253} : s = 372;
	{8'd119,8'd254} : s = 373;
	{8'd119,8'd255} : s = 374;
	{8'd120,8'd0} : s = 120;
	{8'd120,8'd1} : s = 121;
	{8'd120,8'd2} : s = 122;
	{8'd120,8'd3} : s = 123;
	{8'd120,8'd4} : s = 124;
	{8'd120,8'd5} : s = 125;
	{8'd120,8'd6} : s = 126;
	{8'd120,8'd7} : s = 127;
	{8'd120,8'd8} : s = 128;
	{8'd120,8'd9} : s = 129;
	{8'd120,8'd10} : s = 130;
	{8'd120,8'd11} : s = 131;
	{8'd120,8'd12} : s = 132;
	{8'd120,8'd13} : s = 133;
	{8'd120,8'd14} : s = 134;
	{8'd120,8'd15} : s = 135;
	{8'd120,8'd16} : s = 136;
	{8'd120,8'd17} : s = 137;
	{8'd120,8'd18} : s = 138;
	{8'd120,8'd19} : s = 139;
	{8'd120,8'd20} : s = 140;
	{8'd120,8'd21} : s = 141;
	{8'd120,8'd22} : s = 142;
	{8'd120,8'd23} : s = 143;
	{8'd120,8'd24} : s = 144;
	{8'd120,8'd25} : s = 145;
	{8'd120,8'd26} : s = 146;
	{8'd120,8'd27} : s = 147;
	{8'd120,8'd28} : s = 148;
	{8'd120,8'd29} : s = 149;
	{8'd120,8'd30} : s = 150;
	{8'd120,8'd31} : s = 151;
	{8'd120,8'd32} : s = 152;
	{8'd120,8'd33} : s = 153;
	{8'd120,8'd34} : s = 154;
	{8'd120,8'd35} : s = 155;
	{8'd120,8'd36} : s = 156;
	{8'd120,8'd37} : s = 157;
	{8'd120,8'd38} : s = 158;
	{8'd120,8'd39} : s = 159;
	{8'd120,8'd40} : s = 160;
	{8'd120,8'd41} : s = 161;
	{8'd120,8'd42} : s = 162;
	{8'd120,8'd43} : s = 163;
	{8'd120,8'd44} : s = 164;
	{8'd120,8'd45} : s = 165;
	{8'd120,8'd46} : s = 166;
	{8'd120,8'd47} : s = 167;
	{8'd120,8'd48} : s = 168;
	{8'd120,8'd49} : s = 169;
	{8'd120,8'd50} : s = 170;
	{8'd120,8'd51} : s = 171;
	{8'd120,8'd52} : s = 172;
	{8'd120,8'd53} : s = 173;
	{8'd120,8'd54} : s = 174;
	{8'd120,8'd55} : s = 175;
	{8'd120,8'd56} : s = 176;
	{8'd120,8'd57} : s = 177;
	{8'd120,8'd58} : s = 178;
	{8'd120,8'd59} : s = 179;
	{8'd120,8'd60} : s = 180;
	{8'd120,8'd61} : s = 181;
	{8'd120,8'd62} : s = 182;
	{8'd120,8'd63} : s = 183;
	{8'd120,8'd64} : s = 184;
	{8'd120,8'd65} : s = 185;
	{8'd120,8'd66} : s = 186;
	{8'd120,8'd67} : s = 187;
	{8'd120,8'd68} : s = 188;
	{8'd120,8'd69} : s = 189;
	{8'd120,8'd70} : s = 190;
	{8'd120,8'd71} : s = 191;
	{8'd120,8'd72} : s = 192;
	{8'd120,8'd73} : s = 193;
	{8'd120,8'd74} : s = 194;
	{8'd120,8'd75} : s = 195;
	{8'd120,8'd76} : s = 196;
	{8'd120,8'd77} : s = 197;
	{8'd120,8'd78} : s = 198;
	{8'd120,8'd79} : s = 199;
	{8'd120,8'd80} : s = 200;
	{8'd120,8'd81} : s = 201;
	{8'd120,8'd82} : s = 202;
	{8'd120,8'd83} : s = 203;
	{8'd120,8'd84} : s = 204;
	{8'd120,8'd85} : s = 205;
	{8'd120,8'd86} : s = 206;
	{8'd120,8'd87} : s = 207;
	{8'd120,8'd88} : s = 208;
	{8'd120,8'd89} : s = 209;
	{8'd120,8'd90} : s = 210;
	{8'd120,8'd91} : s = 211;
	{8'd120,8'd92} : s = 212;
	{8'd120,8'd93} : s = 213;
	{8'd120,8'd94} : s = 214;
	{8'd120,8'd95} : s = 215;
	{8'd120,8'd96} : s = 216;
	{8'd120,8'd97} : s = 217;
	{8'd120,8'd98} : s = 218;
	{8'd120,8'd99} : s = 219;
	{8'd120,8'd100} : s = 220;
	{8'd120,8'd101} : s = 221;
	{8'd120,8'd102} : s = 222;
	{8'd120,8'd103} : s = 223;
	{8'd120,8'd104} : s = 224;
	{8'd120,8'd105} : s = 225;
	{8'd120,8'd106} : s = 226;
	{8'd120,8'd107} : s = 227;
	{8'd120,8'd108} : s = 228;
	{8'd120,8'd109} : s = 229;
	{8'd120,8'd110} : s = 230;
	{8'd120,8'd111} : s = 231;
	{8'd120,8'd112} : s = 232;
	{8'd120,8'd113} : s = 233;
	{8'd120,8'd114} : s = 234;
	{8'd120,8'd115} : s = 235;
	{8'd120,8'd116} : s = 236;
	{8'd120,8'd117} : s = 237;
	{8'd120,8'd118} : s = 238;
	{8'd120,8'd119} : s = 239;
	{8'd120,8'd120} : s = 240;
	{8'd120,8'd121} : s = 241;
	{8'd120,8'd122} : s = 242;
	{8'd120,8'd123} : s = 243;
	{8'd120,8'd124} : s = 244;
	{8'd120,8'd125} : s = 245;
	{8'd120,8'd126} : s = 246;
	{8'd120,8'd127} : s = 247;
	{8'd120,8'd128} : s = 248;
	{8'd120,8'd129} : s = 249;
	{8'd120,8'd130} : s = 250;
	{8'd120,8'd131} : s = 251;
	{8'd120,8'd132} : s = 252;
	{8'd120,8'd133} : s = 253;
	{8'd120,8'd134} : s = 254;
	{8'd120,8'd135} : s = 255;
	{8'd120,8'd136} : s = 256;
	{8'd120,8'd137} : s = 257;
	{8'd120,8'd138} : s = 258;
	{8'd120,8'd139} : s = 259;
	{8'd120,8'd140} : s = 260;
	{8'd120,8'd141} : s = 261;
	{8'd120,8'd142} : s = 262;
	{8'd120,8'd143} : s = 263;
	{8'd120,8'd144} : s = 264;
	{8'd120,8'd145} : s = 265;
	{8'd120,8'd146} : s = 266;
	{8'd120,8'd147} : s = 267;
	{8'd120,8'd148} : s = 268;
	{8'd120,8'd149} : s = 269;
	{8'd120,8'd150} : s = 270;
	{8'd120,8'd151} : s = 271;
	{8'd120,8'd152} : s = 272;
	{8'd120,8'd153} : s = 273;
	{8'd120,8'd154} : s = 274;
	{8'd120,8'd155} : s = 275;
	{8'd120,8'd156} : s = 276;
	{8'd120,8'd157} : s = 277;
	{8'd120,8'd158} : s = 278;
	{8'd120,8'd159} : s = 279;
	{8'd120,8'd160} : s = 280;
	{8'd120,8'd161} : s = 281;
	{8'd120,8'd162} : s = 282;
	{8'd120,8'd163} : s = 283;
	{8'd120,8'd164} : s = 284;
	{8'd120,8'd165} : s = 285;
	{8'd120,8'd166} : s = 286;
	{8'd120,8'd167} : s = 287;
	{8'd120,8'd168} : s = 288;
	{8'd120,8'd169} : s = 289;
	{8'd120,8'd170} : s = 290;
	{8'd120,8'd171} : s = 291;
	{8'd120,8'd172} : s = 292;
	{8'd120,8'd173} : s = 293;
	{8'd120,8'd174} : s = 294;
	{8'd120,8'd175} : s = 295;
	{8'd120,8'd176} : s = 296;
	{8'd120,8'd177} : s = 297;
	{8'd120,8'd178} : s = 298;
	{8'd120,8'd179} : s = 299;
	{8'd120,8'd180} : s = 300;
	{8'd120,8'd181} : s = 301;
	{8'd120,8'd182} : s = 302;
	{8'd120,8'd183} : s = 303;
	{8'd120,8'd184} : s = 304;
	{8'd120,8'd185} : s = 305;
	{8'd120,8'd186} : s = 306;
	{8'd120,8'd187} : s = 307;
	{8'd120,8'd188} : s = 308;
	{8'd120,8'd189} : s = 309;
	{8'd120,8'd190} : s = 310;
	{8'd120,8'd191} : s = 311;
	{8'd120,8'd192} : s = 312;
	{8'd120,8'd193} : s = 313;
	{8'd120,8'd194} : s = 314;
	{8'd120,8'd195} : s = 315;
	{8'd120,8'd196} : s = 316;
	{8'd120,8'd197} : s = 317;
	{8'd120,8'd198} : s = 318;
	{8'd120,8'd199} : s = 319;
	{8'd120,8'd200} : s = 320;
	{8'd120,8'd201} : s = 321;
	{8'd120,8'd202} : s = 322;
	{8'd120,8'd203} : s = 323;
	{8'd120,8'd204} : s = 324;
	{8'd120,8'd205} : s = 325;
	{8'd120,8'd206} : s = 326;
	{8'd120,8'd207} : s = 327;
	{8'd120,8'd208} : s = 328;
	{8'd120,8'd209} : s = 329;
	{8'd120,8'd210} : s = 330;
	{8'd120,8'd211} : s = 331;
	{8'd120,8'd212} : s = 332;
	{8'd120,8'd213} : s = 333;
	{8'd120,8'd214} : s = 334;
	{8'd120,8'd215} : s = 335;
	{8'd120,8'd216} : s = 336;
	{8'd120,8'd217} : s = 337;
	{8'd120,8'd218} : s = 338;
	{8'd120,8'd219} : s = 339;
	{8'd120,8'd220} : s = 340;
	{8'd120,8'd221} : s = 341;
	{8'd120,8'd222} : s = 342;
	{8'd120,8'd223} : s = 343;
	{8'd120,8'd224} : s = 344;
	{8'd120,8'd225} : s = 345;
	{8'd120,8'd226} : s = 346;
	{8'd120,8'd227} : s = 347;
	{8'd120,8'd228} : s = 348;
	{8'd120,8'd229} : s = 349;
	{8'd120,8'd230} : s = 350;
	{8'd120,8'd231} : s = 351;
	{8'd120,8'd232} : s = 352;
	{8'd120,8'd233} : s = 353;
	{8'd120,8'd234} : s = 354;
	{8'd120,8'd235} : s = 355;
	{8'd120,8'd236} : s = 356;
	{8'd120,8'd237} : s = 357;
	{8'd120,8'd238} : s = 358;
	{8'd120,8'd239} : s = 359;
	{8'd120,8'd240} : s = 360;
	{8'd120,8'd241} : s = 361;
	{8'd120,8'd242} : s = 362;
	{8'd120,8'd243} : s = 363;
	{8'd120,8'd244} : s = 364;
	{8'd120,8'd245} : s = 365;
	{8'd120,8'd246} : s = 366;
	{8'd120,8'd247} : s = 367;
	{8'd120,8'd248} : s = 368;
	{8'd120,8'd249} : s = 369;
	{8'd120,8'd250} : s = 370;
	{8'd120,8'd251} : s = 371;
	{8'd120,8'd252} : s = 372;
	{8'd120,8'd253} : s = 373;
	{8'd120,8'd254} : s = 374;
	{8'd120,8'd255} : s = 375;
	{8'd121,8'd0} : s = 121;
	{8'd121,8'd1} : s = 122;
	{8'd121,8'd2} : s = 123;
	{8'd121,8'd3} : s = 124;
	{8'd121,8'd4} : s = 125;
	{8'd121,8'd5} : s = 126;
	{8'd121,8'd6} : s = 127;
	{8'd121,8'd7} : s = 128;
	{8'd121,8'd8} : s = 129;
	{8'd121,8'd9} : s = 130;
	{8'd121,8'd10} : s = 131;
	{8'd121,8'd11} : s = 132;
	{8'd121,8'd12} : s = 133;
	{8'd121,8'd13} : s = 134;
	{8'd121,8'd14} : s = 135;
	{8'd121,8'd15} : s = 136;
	{8'd121,8'd16} : s = 137;
	{8'd121,8'd17} : s = 138;
	{8'd121,8'd18} : s = 139;
	{8'd121,8'd19} : s = 140;
	{8'd121,8'd20} : s = 141;
	{8'd121,8'd21} : s = 142;
	{8'd121,8'd22} : s = 143;
	{8'd121,8'd23} : s = 144;
	{8'd121,8'd24} : s = 145;
	{8'd121,8'd25} : s = 146;
	{8'd121,8'd26} : s = 147;
	{8'd121,8'd27} : s = 148;
	{8'd121,8'd28} : s = 149;
	{8'd121,8'd29} : s = 150;
	{8'd121,8'd30} : s = 151;
	{8'd121,8'd31} : s = 152;
	{8'd121,8'd32} : s = 153;
	{8'd121,8'd33} : s = 154;
	{8'd121,8'd34} : s = 155;
	{8'd121,8'd35} : s = 156;
	{8'd121,8'd36} : s = 157;
	{8'd121,8'd37} : s = 158;
	{8'd121,8'd38} : s = 159;
	{8'd121,8'd39} : s = 160;
	{8'd121,8'd40} : s = 161;
	{8'd121,8'd41} : s = 162;
	{8'd121,8'd42} : s = 163;
	{8'd121,8'd43} : s = 164;
	{8'd121,8'd44} : s = 165;
	{8'd121,8'd45} : s = 166;
	{8'd121,8'd46} : s = 167;
	{8'd121,8'd47} : s = 168;
	{8'd121,8'd48} : s = 169;
	{8'd121,8'd49} : s = 170;
	{8'd121,8'd50} : s = 171;
	{8'd121,8'd51} : s = 172;
	{8'd121,8'd52} : s = 173;
	{8'd121,8'd53} : s = 174;
	{8'd121,8'd54} : s = 175;
	{8'd121,8'd55} : s = 176;
	{8'd121,8'd56} : s = 177;
	{8'd121,8'd57} : s = 178;
	{8'd121,8'd58} : s = 179;
	{8'd121,8'd59} : s = 180;
	{8'd121,8'd60} : s = 181;
	{8'd121,8'd61} : s = 182;
	{8'd121,8'd62} : s = 183;
	{8'd121,8'd63} : s = 184;
	{8'd121,8'd64} : s = 185;
	{8'd121,8'd65} : s = 186;
	{8'd121,8'd66} : s = 187;
	{8'd121,8'd67} : s = 188;
	{8'd121,8'd68} : s = 189;
	{8'd121,8'd69} : s = 190;
	{8'd121,8'd70} : s = 191;
	{8'd121,8'd71} : s = 192;
	{8'd121,8'd72} : s = 193;
	{8'd121,8'd73} : s = 194;
	{8'd121,8'd74} : s = 195;
	{8'd121,8'd75} : s = 196;
	{8'd121,8'd76} : s = 197;
	{8'd121,8'd77} : s = 198;
	{8'd121,8'd78} : s = 199;
	{8'd121,8'd79} : s = 200;
	{8'd121,8'd80} : s = 201;
	{8'd121,8'd81} : s = 202;
	{8'd121,8'd82} : s = 203;
	{8'd121,8'd83} : s = 204;
	{8'd121,8'd84} : s = 205;
	{8'd121,8'd85} : s = 206;
	{8'd121,8'd86} : s = 207;
	{8'd121,8'd87} : s = 208;
	{8'd121,8'd88} : s = 209;
	{8'd121,8'd89} : s = 210;
	{8'd121,8'd90} : s = 211;
	{8'd121,8'd91} : s = 212;
	{8'd121,8'd92} : s = 213;
	{8'd121,8'd93} : s = 214;
	{8'd121,8'd94} : s = 215;
	{8'd121,8'd95} : s = 216;
	{8'd121,8'd96} : s = 217;
	{8'd121,8'd97} : s = 218;
	{8'd121,8'd98} : s = 219;
	{8'd121,8'd99} : s = 220;
	{8'd121,8'd100} : s = 221;
	{8'd121,8'd101} : s = 222;
	{8'd121,8'd102} : s = 223;
	{8'd121,8'd103} : s = 224;
	{8'd121,8'd104} : s = 225;
	{8'd121,8'd105} : s = 226;
	{8'd121,8'd106} : s = 227;
	{8'd121,8'd107} : s = 228;
	{8'd121,8'd108} : s = 229;
	{8'd121,8'd109} : s = 230;
	{8'd121,8'd110} : s = 231;
	{8'd121,8'd111} : s = 232;
	{8'd121,8'd112} : s = 233;
	{8'd121,8'd113} : s = 234;
	{8'd121,8'd114} : s = 235;
	{8'd121,8'd115} : s = 236;
	{8'd121,8'd116} : s = 237;
	{8'd121,8'd117} : s = 238;
	{8'd121,8'd118} : s = 239;
	{8'd121,8'd119} : s = 240;
	{8'd121,8'd120} : s = 241;
	{8'd121,8'd121} : s = 242;
	{8'd121,8'd122} : s = 243;
	{8'd121,8'd123} : s = 244;
	{8'd121,8'd124} : s = 245;
	{8'd121,8'd125} : s = 246;
	{8'd121,8'd126} : s = 247;
	{8'd121,8'd127} : s = 248;
	{8'd121,8'd128} : s = 249;
	{8'd121,8'd129} : s = 250;
	{8'd121,8'd130} : s = 251;
	{8'd121,8'd131} : s = 252;
	{8'd121,8'd132} : s = 253;
	{8'd121,8'd133} : s = 254;
	{8'd121,8'd134} : s = 255;
	{8'd121,8'd135} : s = 256;
	{8'd121,8'd136} : s = 257;
	{8'd121,8'd137} : s = 258;
	{8'd121,8'd138} : s = 259;
	{8'd121,8'd139} : s = 260;
	{8'd121,8'd140} : s = 261;
	{8'd121,8'd141} : s = 262;
	{8'd121,8'd142} : s = 263;
	{8'd121,8'd143} : s = 264;
	{8'd121,8'd144} : s = 265;
	{8'd121,8'd145} : s = 266;
	{8'd121,8'd146} : s = 267;
	{8'd121,8'd147} : s = 268;
	{8'd121,8'd148} : s = 269;
	{8'd121,8'd149} : s = 270;
	{8'd121,8'd150} : s = 271;
	{8'd121,8'd151} : s = 272;
	{8'd121,8'd152} : s = 273;
	{8'd121,8'd153} : s = 274;
	{8'd121,8'd154} : s = 275;
	{8'd121,8'd155} : s = 276;
	{8'd121,8'd156} : s = 277;
	{8'd121,8'd157} : s = 278;
	{8'd121,8'd158} : s = 279;
	{8'd121,8'd159} : s = 280;
	{8'd121,8'd160} : s = 281;
	{8'd121,8'd161} : s = 282;
	{8'd121,8'd162} : s = 283;
	{8'd121,8'd163} : s = 284;
	{8'd121,8'd164} : s = 285;
	{8'd121,8'd165} : s = 286;
	{8'd121,8'd166} : s = 287;
	{8'd121,8'd167} : s = 288;
	{8'd121,8'd168} : s = 289;
	{8'd121,8'd169} : s = 290;
	{8'd121,8'd170} : s = 291;
	{8'd121,8'd171} : s = 292;
	{8'd121,8'd172} : s = 293;
	{8'd121,8'd173} : s = 294;
	{8'd121,8'd174} : s = 295;
	{8'd121,8'd175} : s = 296;
	{8'd121,8'd176} : s = 297;
	{8'd121,8'd177} : s = 298;
	{8'd121,8'd178} : s = 299;
	{8'd121,8'd179} : s = 300;
	{8'd121,8'd180} : s = 301;
	{8'd121,8'd181} : s = 302;
	{8'd121,8'd182} : s = 303;
	{8'd121,8'd183} : s = 304;
	{8'd121,8'd184} : s = 305;
	{8'd121,8'd185} : s = 306;
	{8'd121,8'd186} : s = 307;
	{8'd121,8'd187} : s = 308;
	{8'd121,8'd188} : s = 309;
	{8'd121,8'd189} : s = 310;
	{8'd121,8'd190} : s = 311;
	{8'd121,8'd191} : s = 312;
	{8'd121,8'd192} : s = 313;
	{8'd121,8'd193} : s = 314;
	{8'd121,8'd194} : s = 315;
	{8'd121,8'd195} : s = 316;
	{8'd121,8'd196} : s = 317;
	{8'd121,8'd197} : s = 318;
	{8'd121,8'd198} : s = 319;
	{8'd121,8'd199} : s = 320;
	{8'd121,8'd200} : s = 321;
	{8'd121,8'd201} : s = 322;
	{8'd121,8'd202} : s = 323;
	{8'd121,8'd203} : s = 324;
	{8'd121,8'd204} : s = 325;
	{8'd121,8'd205} : s = 326;
	{8'd121,8'd206} : s = 327;
	{8'd121,8'd207} : s = 328;
	{8'd121,8'd208} : s = 329;
	{8'd121,8'd209} : s = 330;
	{8'd121,8'd210} : s = 331;
	{8'd121,8'd211} : s = 332;
	{8'd121,8'd212} : s = 333;
	{8'd121,8'd213} : s = 334;
	{8'd121,8'd214} : s = 335;
	{8'd121,8'd215} : s = 336;
	{8'd121,8'd216} : s = 337;
	{8'd121,8'd217} : s = 338;
	{8'd121,8'd218} : s = 339;
	{8'd121,8'd219} : s = 340;
	{8'd121,8'd220} : s = 341;
	{8'd121,8'd221} : s = 342;
	{8'd121,8'd222} : s = 343;
	{8'd121,8'd223} : s = 344;
	{8'd121,8'd224} : s = 345;
	{8'd121,8'd225} : s = 346;
	{8'd121,8'd226} : s = 347;
	{8'd121,8'd227} : s = 348;
	{8'd121,8'd228} : s = 349;
	{8'd121,8'd229} : s = 350;
	{8'd121,8'd230} : s = 351;
	{8'd121,8'd231} : s = 352;
	{8'd121,8'd232} : s = 353;
	{8'd121,8'd233} : s = 354;
	{8'd121,8'd234} : s = 355;
	{8'd121,8'd235} : s = 356;
	{8'd121,8'd236} : s = 357;
	{8'd121,8'd237} : s = 358;
	{8'd121,8'd238} : s = 359;
	{8'd121,8'd239} : s = 360;
	{8'd121,8'd240} : s = 361;
	{8'd121,8'd241} : s = 362;
	{8'd121,8'd242} : s = 363;
	{8'd121,8'd243} : s = 364;
	{8'd121,8'd244} : s = 365;
	{8'd121,8'd245} : s = 366;
	{8'd121,8'd246} : s = 367;
	{8'd121,8'd247} : s = 368;
	{8'd121,8'd248} : s = 369;
	{8'd121,8'd249} : s = 370;
	{8'd121,8'd250} : s = 371;
	{8'd121,8'd251} : s = 372;
	{8'd121,8'd252} : s = 373;
	{8'd121,8'd253} : s = 374;
	{8'd121,8'd254} : s = 375;
	{8'd121,8'd255} : s = 376;
	{8'd122,8'd0} : s = 122;
	{8'd122,8'd1} : s = 123;
	{8'd122,8'd2} : s = 124;
	{8'd122,8'd3} : s = 125;
	{8'd122,8'd4} : s = 126;
	{8'd122,8'd5} : s = 127;
	{8'd122,8'd6} : s = 128;
	{8'd122,8'd7} : s = 129;
	{8'd122,8'd8} : s = 130;
	{8'd122,8'd9} : s = 131;
	{8'd122,8'd10} : s = 132;
	{8'd122,8'd11} : s = 133;
	{8'd122,8'd12} : s = 134;
	{8'd122,8'd13} : s = 135;
	{8'd122,8'd14} : s = 136;
	{8'd122,8'd15} : s = 137;
	{8'd122,8'd16} : s = 138;
	{8'd122,8'd17} : s = 139;
	{8'd122,8'd18} : s = 140;
	{8'd122,8'd19} : s = 141;
	{8'd122,8'd20} : s = 142;
	{8'd122,8'd21} : s = 143;
	{8'd122,8'd22} : s = 144;
	{8'd122,8'd23} : s = 145;
	{8'd122,8'd24} : s = 146;
	{8'd122,8'd25} : s = 147;
	{8'd122,8'd26} : s = 148;
	{8'd122,8'd27} : s = 149;
	{8'd122,8'd28} : s = 150;
	{8'd122,8'd29} : s = 151;
	{8'd122,8'd30} : s = 152;
	{8'd122,8'd31} : s = 153;
	{8'd122,8'd32} : s = 154;
	{8'd122,8'd33} : s = 155;
	{8'd122,8'd34} : s = 156;
	{8'd122,8'd35} : s = 157;
	{8'd122,8'd36} : s = 158;
	{8'd122,8'd37} : s = 159;
	{8'd122,8'd38} : s = 160;
	{8'd122,8'd39} : s = 161;
	{8'd122,8'd40} : s = 162;
	{8'd122,8'd41} : s = 163;
	{8'd122,8'd42} : s = 164;
	{8'd122,8'd43} : s = 165;
	{8'd122,8'd44} : s = 166;
	{8'd122,8'd45} : s = 167;
	{8'd122,8'd46} : s = 168;
	{8'd122,8'd47} : s = 169;
	{8'd122,8'd48} : s = 170;
	{8'd122,8'd49} : s = 171;
	{8'd122,8'd50} : s = 172;
	{8'd122,8'd51} : s = 173;
	{8'd122,8'd52} : s = 174;
	{8'd122,8'd53} : s = 175;
	{8'd122,8'd54} : s = 176;
	{8'd122,8'd55} : s = 177;
	{8'd122,8'd56} : s = 178;
	{8'd122,8'd57} : s = 179;
	{8'd122,8'd58} : s = 180;
	{8'd122,8'd59} : s = 181;
	{8'd122,8'd60} : s = 182;
	{8'd122,8'd61} : s = 183;
	{8'd122,8'd62} : s = 184;
	{8'd122,8'd63} : s = 185;
	{8'd122,8'd64} : s = 186;
	{8'd122,8'd65} : s = 187;
	{8'd122,8'd66} : s = 188;
	{8'd122,8'd67} : s = 189;
	{8'd122,8'd68} : s = 190;
	{8'd122,8'd69} : s = 191;
	{8'd122,8'd70} : s = 192;
	{8'd122,8'd71} : s = 193;
	{8'd122,8'd72} : s = 194;
	{8'd122,8'd73} : s = 195;
	{8'd122,8'd74} : s = 196;
	{8'd122,8'd75} : s = 197;
	{8'd122,8'd76} : s = 198;
	{8'd122,8'd77} : s = 199;
	{8'd122,8'd78} : s = 200;
	{8'd122,8'd79} : s = 201;
	{8'd122,8'd80} : s = 202;
	{8'd122,8'd81} : s = 203;
	{8'd122,8'd82} : s = 204;
	{8'd122,8'd83} : s = 205;
	{8'd122,8'd84} : s = 206;
	{8'd122,8'd85} : s = 207;
	{8'd122,8'd86} : s = 208;
	{8'd122,8'd87} : s = 209;
	{8'd122,8'd88} : s = 210;
	{8'd122,8'd89} : s = 211;
	{8'd122,8'd90} : s = 212;
	{8'd122,8'd91} : s = 213;
	{8'd122,8'd92} : s = 214;
	{8'd122,8'd93} : s = 215;
	{8'd122,8'd94} : s = 216;
	{8'd122,8'd95} : s = 217;
	{8'd122,8'd96} : s = 218;
	{8'd122,8'd97} : s = 219;
	{8'd122,8'd98} : s = 220;
	{8'd122,8'd99} : s = 221;
	{8'd122,8'd100} : s = 222;
	{8'd122,8'd101} : s = 223;
	{8'd122,8'd102} : s = 224;
	{8'd122,8'd103} : s = 225;
	{8'd122,8'd104} : s = 226;
	{8'd122,8'd105} : s = 227;
	{8'd122,8'd106} : s = 228;
	{8'd122,8'd107} : s = 229;
	{8'd122,8'd108} : s = 230;
	{8'd122,8'd109} : s = 231;
	{8'd122,8'd110} : s = 232;
	{8'd122,8'd111} : s = 233;
	{8'd122,8'd112} : s = 234;
	{8'd122,8'd113} : s = 235;
	{8'd122,8'd114} : s = 236;
	{8'd122,8'd115} : s = 237;
	{8'd122,8'd116} : s = 238;
	{8'd122,8'd117} : s = 239;
	{8'd122,8'd118} : s = 240;
	{8'd122,8'd119} : s = 241;
	{8'd122,8'd120} : s = 242;
	{8'd122,8'd121} : s = 243;
	{8'd122,8'd122} : s = 244;
	{8'd122,8'd123} : s = 245;
	{8'd122,8'd124} : s = 246;
	{8'd122,8'd125} : s = 247;
	{8'd122,8'd126} : s = 248;
	{8'd122,8'd127} : s = 249;
	{8'd122,8'd128} : s = 250;
	{8'd122,8'd129} : s = 251;
	{8'd122,8'd130} : s = 252;
	{8'd122,8'd131} : s = 253;
	{8'd122,8'd132} : s = 254;
	{8'd122,8'd133} : s = 255;
	{8'd122,8'd134} : s = 256;
	{8'd122,8'd135} : s = 257;
	{8'd122,8'd136} : s = 258;
	{8'd122,8'd137} : s = 259;
	{8'd122,8'd138} : s = 260;
	{8'd122,8'd139} : s = 261;
	{8'd122,8'd140} : s = 262;
	{8'd122,8'd141} : s = 263;
	{8'd122,8'd142} : s = 264;
	{8'd122,8'd143} : s = 265;
	{8'd122,8'd144} : s = 266;
	{8'd122,8'd145} : s = 267;
	{8'd122,8'd146} : s = 268;
	{8'd122,8'd147} : s = 269;
	{8'd122,8'd148} : s = 270;
	{8'd122,8'd149} : s = 271;
	{8'd122,8'd150} : s = 272;
	{8'd122,8'd151} : s = 273;
	{8'd122,8'd152} : s = 274;
	{8'd122,8'd153} : s = 275;
	{8'd122,8'd154} : s = 276;
	{8'd122,8'd155} : s = 277;
	{8'd122,8'd156} : s = 278;
	{8'd122,8'd157} : s = 279;
	{8'd122,8'd158} : s = 280;
	{8'd122,8'd159} : s = 281;
	{8'd122,8'd160} : s = 282;
	{8'd122,8'd161} : s = 283;
	{8'd122,8'd162} : s = 284;
	{8'd122,8'd163} : s = 285;
	{8'd122,8'd164} : s = 286;
	{8'd122,8'd165} : s = 287;
	{8'd122,8'd166} : s = 288;
	{8'd122,8'd167} : s = 289;
	{8'd122,8'd168} : s = 290;
	{8'd122,8'd169} : s = 291;
	{8'd122,8'd170} : s = 292;
	{8'd122,8'd171} : s = 293;
	{8'd122,8'd172} : s = 294;
	{8'd122,8'd173} : s = 295;
	{8'd122,8'd174} : s = 296;
	{8'd122,8'd175} : s = 297;
	{8'd122,8'd176} : s = 298;
	{8'd122,8'd177} : s = 299;
	{8'd122,8'd178} : s = 300;
	{8'd122,8'd179} : s = 301;
	{8'd122,8'd180} : s = 302;
	{8'd122,8'd181} : s = 303;
	{8'd122,8'd182} : s = 304;
	{8'd122,8'd183} : s = 305;
	{8'd122,8'd184} : s = 306;
	{8'd122,8'd185} : s = 307;
	{8'd122,8'd186} : s = 308;
	{8'd122,8'd187} : s = 309;
	{8'd122,8'd188} : s = 310;
	{8'd122,8'd189} : s = 311;
	{8'd122,8'd190} : s = 312;
	{8'd122,8'd191} : s = 313;
	{8'd122,8'd192} : s = 314;
	{8'd122,8'd193} : s = 315;
	{8'd122,8'd194} : s = 316;
	{8'd122,8'd195} : s = 317;
	{8'd122,8'd196} : s = 318;
	{8'd122,8'd197} : s = 319;
	{8'd122,8'd198} : s = 320;
	{8'd122,8'd199} : s = 321;
	{8'd122,8'd200} : s = 322;
	{8'd122,8'd201} : s = 323;
	{8'd122,8'd202} : s = 324;
	{8'd122,8'd203} : s = 325;
	{8'd122,8'd204} : s = 326;
	{8'd122,8'd205} : s = 327;
	{8'd122,8'd206} : s = 328;
	{8'd122,8'd207} : s = 329;
	{8'd122,8'd208} : s = 330;
	{8'd122,8'd209} : s = 331;
	{8'd122,8'd210} : s = 332;
	{8'd122,8'd211} : s = 333;
	{8'd122,8'd212} : s = 334;
	{8'd122,8'd213} : s = 335;
	{8'd122,8'd214} : s = 336;
	{8'd122,8'd215} : s = 337;
	{8'd122,8'd216} : s = 338;
	{8'd122,8'd217} : s = 339;
	{8'd122,8'd218} : s = 340;
	{8'd122,8'd219} : s = 341;
	{8'd122,8'd220} : s = 342;
	{8'd122,8'd221} : s = 343;
	{8'd122,8'd222} : s = 344;
	{8'd122,8'd223} : s = 345;
	{8'd122,8'd224} : s = 346;
	{8'd122,8'd225} : s = 347;
	{8'd122,8'd226} : s = 348;
	{8'd122,8'd227} : s = 349;
	{8'd122,8'd228} : s = 350;
	{8'd122,8'd229} : s = 351;
	{8'd122,8'd230} : s = 352;
	{8'd122,8'd231} : s = 353;
	{8'd122,8'd232} : s = 354;
	{8'd122,8'd233} : s = 355;
	{8'd122,8'd234} : s = 356;
	{8'd122,8'd235} : s = 357;
	{8'd122,8'd236} : s = 358;
	{8'd122,8'd237} : s = 359;
	{8'd122,8'd238} : s = 360;
	{8'd122,8'd239} : s = 361;
	{8'd122,8'd240} : s = 362;
	{8'd122,8'd241} : s = 363;
	{8'd122,8'd242} : s = 364;
	{8'd122,8'd243} : s = 365;
	{8'd122,8'd244} : s = 366;
	{8'd122,8'd245} : s = 367;
	{8'd122,8'd246} : s = 368;
	{8'd122,8'd247} : s = 369;
	{8'd122,8'd248} : s = 370;
	{8'd122,8'd249} : s = 371;
	{8'd122,8'd250} : s = 372;
	{8'd122,8'd251} : s = 373;
	{8'd122,8'd252} : s = 374;
	{8'd122,8'd253} : s = 375;
	{8'd122,8'd254} : s = 376;
	{8'd122,8'd255} : s = 377;
	{8'd123,8'd0} : s = 123;
	{8'd123,8'd1} : s = 124;
	{8'd123,8'd2} : s = 125;
	{8'd123,8'd3} : s = 126;
	{8'd123,8'd4} : s = 127;
	{8'd123,8'd5} : s = 128;
	{8'd123,8'd6} : s = 129;
	{8'd123,8'd7} : s = 130;
	{8'd123,8'd8} : s = 131;
	{8'd123,8'd9} : s = 132;
	{8'd123,8'd10} : s = 133;
	{8'd123,8'd11} : s = 134;
	{8'd123,8'd12} : s = 135;
	{8'd123,8'd13} : s = 136;
	{8'd123,8'd14} : s = 137;
	{8'd123,8'd15} : s = 138;
	{8'd123,8'd16} : s = 139;
	{8'd123,8'd17} : s = 140;
	{8'd123,8'd18} : s = 141;
	{8'd123,8'd19} : s = 142;
	{8'd123,8'd20} : s = 143;
	{8'd123,8'd21} : s = 144;
	{8'd123,8'd22} : s = 145;
	{8'd123,8'd23} : s = 146;
	{8'd123,8'd24} : s = 147;
	{8'd123,8'd25} : s = 148;
	{8'd123,8'd26} : s = 149;
	{8'd123,8'd27} : s = 150;
	{8'd123,8'd28} : s = 151;
	{8'd123,8'd29} : s = 152;
	{8'd123,8'd30} : s = 153;
	{8'd123,8'd31} : s = 154;
	{8'd123,8'd32} : s = 155;
	{8'd123,8'd33} : s = 156;
	{8'd123,8'd34} : s = 157;
	{8'd123,8'd35} : s = 158;
	{8'd123,8'd36} : s = 159;
	{8'd123,8'd37} : s = 160;
	{8'd123,8'd38} : s = 161;
	{8'd123,8'd39} : s = 162;
	{8'd123,8'd40} : s = 163;
	{8'd123,8'd41} : s = 164;
	{8'd123,8'd42} : s = 165;
	{8'd123,8'd43} : s = 166;
	{8'd123,8'd44} : s = 167;
	{8'd123,8'd45} : s = 168;
	{8'd123,8'd46} : s = 169;
	{8'd123,8'd47} : s = 170;
	{8'd123,8'd48} : s = 171;
	{8'd123,8'd49} : s = 172;
	{8'd123,8'd50} : s = 173;
	{8'd123,8'd51} : s = 174;
	{8'd123,8'd52} : s = 175;
	{8'd123,8'd53} : s = 176;
	{8'd123,8'd54} : s = 177;
	{8'd123,8'd55} : s = 178;
	{8'd123,8'd56} : s = 179;
	{8'd123,8'd57} : s = 180;
	{8'd123,8'd58} : s = 181;
	{8'd123,8'd59} : s = 182;
	{8'd123,8'd60} : s = 183;
	{8'd123,8'd61} : s = 184;
	{8'd123,8'd62} : s = 185;
	{8'd123,8'd63} : s = 186;
	{8'd123,8'd64} : s = 187;
	{8'd123,8'd65} : s = 188;
	{8'd123,8'd66} : s = 189;
	{8'd123,8'd67} : s = 190;
	{8'd123,8'd68} : s = 191;
	{8'd123,8'd69} : s = 192;
	{8'd123,8'd70} : s = 193;
	{8'd123,8'd71} : s = 194;
	{8'd123,8'd72} : s = 195;
	{8'd123,8'd73} : s = 196;
	{8'd123,8'd74} : s = 197;
	{8'd123,8'd75} : s = 198;
	{8'd123,8'd76} : s = 199;
	{8'd123,8'd77} : s = 200;
	{8'd123,8'd78} : s = 201;
	{8'd123,8'd79} : s = 202;
	{8'd123,8'd80} : s = 203;
	{8'd123,8'd81} : s = 204;
	{8'd123,8'd82} : s = 205;
	{8'd123,8'd83} : s = 206;
	{8'd123,8'd84} : s = 207;
	{8'd123,8'd85} : s = 208;
	{8'd123,8'd86} : s = 209;
	{8'd123,8'd87} : s = 210;
	{8'd123,8'd88} : s = 211;
	{8'd123,8'd89} : s = 212;
	{8'd123,8'd90} : s = 213;
	{8'd123,8'd91} : s = 214;
	{8'd123,8'd92} : s = 215;
	{8'd123,8'd93} : s = 216;
	{8'd123,8'd94} : s = 217;
	{8'd123,8'd95} : s = 218;
	{8'd123,8'd96} : s = 219;
	{8'd123,8'd97} : s = 220;
	{8'd123,8'd98} : s = 221;
	{8'd123,8'd99} : s = 222;
	{8'd123,8'd100} : s = 223;
	{8'd123,8'd101} : s = 224;
	{8'd123,8'd102} : s = 225;
	{8'd123,8'd103} : s = 226;
	{8'd123,8'd104} : s = 227;
	{8'd123,8'd105} : s = 228;
	{8'd123,8'd106} : s = 229;
	{8'd123,8'd107} : s = 230;
	{8'd123,8'd108} : s = 231;
	{8'd123,8'd109} : s = 232;
	{8'd123,8'd110} : s = 233;
	{8'd123,8'd111} : s = 234;
	{8'd123,8'd112} : s = 235;
	{8'd123,8'd113} : s = 236;
	{8'd123,8'd114} : s = 237;
	{8'd123,8'd115} : s = 238;
	{8'd123,8'd116} : s = 239;
	{8'd123,8'd117} : s = 240;
	{8'd123,8'd118} : s = 241;
	{8'd123,8'd119} : s = 242;
	{8'd123,8'd120} : s = 243;
	{8'd123,8'd121} : s = 244;
	{8'd123,8'd122} : s = 245;
	{8'd123,8'd123} : s = 246;
	{8'd123,8'd124} : s = 247;
	{8'd123,8'd125} : s = 248;
	{8'd123,8'd126} : s = 249;
	{8'd123,8'd127} : s = 250;
	{8'd123,8'd128} : s = 251;
	{8'd123,8'd129} : s = 252;
	{8'd123,8'd130} : s = 253;
	{8'd123,8'd131} : s = 254;
	{8'd123,8'd132} : s = 255;
	{8'd123,8'd133} : s = 256;
	{8'd123,8'd134} : s = 257;
	{8'd123,8'd135} : s = 258;
	{8'd123,8'd136} : s = 259;
	{8'd123,8'd137} : s = 260;
	{8'd123,8'd138} : s = 261;
	{8'd123,8'd139} : s = 262;
	{8'd123,8'd140} : s = 263;
	{8'd123,8'd141} : s = 264;
	{8'd123,8'd142} : s = 265;
	{8'd123,8'd143} : s = 266;
	{8'd123,8'd144} : s = 267;
	{8'd123,8'd145} : s = 268;
	{8'd123,8'd146} : s = 269;
	{8'd123,8'd147} : s = 270;
	{8'd123,8'd148} : s = 271;
	{8'd123,8'd149} : s = 272;
	{8'd123,8'd150} : s = 273;
	{8'd123,8'd151} : s = 274;
	{8'd123,8'd152} : s = 275;
	{8'd123,8'd153} : s = 276;
	{8'd123,8'd154} : s = 277;
	{8'd123,8'd155} : s = 278;
	{8'd123,8'd156} : s = 279;
	{8'd123,8'd157} : s = 280;
	{8'd123,8'd158} : s = 281;
	{8'd123,8'd159} : s = 282;
	{8'd123,8'd160} : s = 283;
	{8'd123,8'd161} : s = 284;
	{8'd123,8'd162} : s = 285;
	{8'd123,8'd163} : s = 286;
	{8'd123,8'd164} : s = 287;
	{8'd123,8'd165} : s = 288;
	{8'd123,8'd166} : s = 289;
	{8'd123,8'd167} : s = 290;
	{8'd123,8'd168} : s = 291;
	{8'd123,8'd169} : s = 292;
	{8'd123,8'd170} : s = 293;
	{8'd123,8'd171} : s = 294;
	{8'd123,8'd172} : s = 295;
	{8'd123,8'd173} : s = 296;
	{8'd123,8'd174} : s = 297;
	{8'd123,8'd175} : s = 298;
	{8'd123,8'd176} : s = 299;
	{8'd123,8'd177} : s = 300;
	{8'd123,8'd178} : s = 301;
	{8'd123,8'd179} : s = 302;
	{8'd123,8'd180} : s = 303;
	{8'd123,8'd181} : s = 304;
	{8'd123,8'd182} : s = 305;
	{8'd123,8'd183} : s = 306;
	{8'd123,8'd184} : s = 307;
	{8'd123,8'd185} : s = 308;
	{8'd123,8'd186} : s = 309;
	{8'd123,8'd187} : s = 310;
	{8'd123,8'd188} : s = 311;
	{8'd123,8'd189} : s = 312;
	{8'd123,8'd190} : s = 313;
	{8'd123,8'd191} : s = 314;
	{8'd123,8'd192} : s = 315;
	{8'd123,8'd193} : s = 316;
	{8'd123,8'd194} : s = 317;
	{8'd123,8'd195} : s = 318;
	{8'd123,8'd196} : s = 319;
	{8'd123,8'd197} : s = 320;
	{8'd123,8'd198} : s = 321;
	{8'd123,8'd199} : s = 322;
	{8'd123,8'd200} : s = 323;
	{8'd123,8'd201} : s = 324;
	{8'd123,8'd202} : s = 325;
	{8'd123,8'd203} : s = 326;
	{8'd123,8'd204} : s = 327;
	{8'd123,8'd205} : s = 328;
	{8'd123,8'd206} : s = 329;
	{8'd123,8'd207} : s = 330;
	{8'd123,8'd208} : s = 331;
	{8'd123,8'd209} : s = 332;
	{8'd123,8'd210} : s = 333;
	{8'd123,8'd211} : s = 334;
	{8'd123,8'd212} : s = 335;
	{8'd123,8'd213} : s = 336;
	{8'd123,8'd214} : s = 337;
	{8'd123,8'd215} : s = 338;
	{8'd123,8'd216} : s = 339;
	{8'd123,8'd217} : s = 340;
	{8'd123,8'd218} : s = 341;
	{8'd123,8'd219} : s = 342;
	{8'd123,8'd220} : s = 343;
	{8'd123,8'd221} : s = 344;
	{8'd123,8'd222} : s = 345;
	{8'd123,8'd223} : s = 346;
	{8'd123,8'd224} : s = 347;
	{8'd123,8'd225} : s = 348;
	{8'd123,8'd226} : s = 349;
	{8'd123,8'd227} : s = 350;
	{8'd123,8'd228} : s = 351;
	{8'd123,8'd229} : s = 352;
	{8'd123,8'd230} : s = 353;
	{8'd123,8'd231} : s = 354;
	{8'd123,8'd232} : s = 355;
	{8'd123,8'd233} : s = 356;
	{8'd123,8'd234} : s = 357;
	{8'd123,8'd235} : s = 358;
	{8'd123,8'd236} : s = 359;
	{8'd123,8'd237} : s = 360;
	{8'd123,8'd238} : s = 361;
	{8'd123,8'd239} : s = 362;
	{8'd123,8'd240} : s = 363;
	{8'd123,8'd241} : s = 364;
	{8'd123,8'd242} : s = 365;
	{8'd123,8'd243} : s = 366;
	{8'd123,8'd244} : s = 367;
	{8'd123,8'd245} : s = 368;
	{8'd123,8'd246} : s = 369;
	{8'd123,8'd247} : s = 370;
	{8'd123,8'd248} : s = 371;
	{8'd123,8'd249} : s = 372;
	{8'd123,8'd250} : s = 373;
	{8'd123,8'd251} : s = 374;
	{8'd123,8'd252} : s = 375;
	{8'd123,8'd253} : s = 376;
	{8'd123,8'd254} : s = 377;
	{8'd123,8'd255} : s = 378;
	{8'd124,8'd0} : s = 124;
	{8'd124,8'd1} : s = 125;
	{8'd124,8'd2} : s = 126;
	{8'd124,8'd3} : s = 127;
	{8'd124,8'd4} : s = 128;
	{8'd124,8'd5} : s = 129;
	{8'd124,8'd6} : s = 130;
	{8'd124,8'd7} : s = 131;
	{8'd124,8'd8} : s = 132;
	{8'd124,8'd9} : s = 133;
	{8'd124,8'd10} : s = 134;
	{8'd124,8'd11} : s = 135;
	{8'd124,8'd12} : s = 136;
	{8'd124,8'd13} : s = 137;
	{8'd124,8'd14} : s = 138;
	{8'd124,8'd15} : s = 139;
	{8'd124,8'd16} : s = 140;
	{8'd124,8'd17} : s = 141;
	{8'd124,8'd18} : s = 142;
	{8'd124,8'd19} : s = 143;
	{8'd124,8'd20} : s = 144;
	{8'd124,8'd21} : s = 145;
	{8'd124,8'd22} : s = 146;
	{8'd124,8'd23} : s = 147;
	{8'd124,8'd24} : s = 148;
	{8'd124,8'd25} : s = 149;
	{8'd124,8'd26} : s = 150;
	{8'd124,8'd27} : s = 151;
	{8'd124,8'd28} : s = 152;
	{8'd124,8'd29} : s = 153;
	{8'd124,8'd30} : s = 154;
	{8'd124,8'd31} : s = 155;
	{8'd124,8'd32} : s = 156;
	{8'd124,8'd33} : s = 157;
	{8'd124,8'd34} : s = 158;
	{8'd124,8'd35} : s = 159;
	{8'd124,8'd36} : s = 160;
	{8'd124,8'd37} : s = 161;
	{8'd124,8'd38} : s = 162;
	{8'd124,8'd39} : s = 163;
	{8'd124,8'd40} : s = 164;
	{8'd124,8'd41} : s = 165;
	{8'd124,8'd42} : s = 166;
	{8'd124,8'd43} : s = 167;
	{8'd124,8'd44} : s = 168;
	{8'd124,8'd45} : s = 169;
	{8'd124,8'd46} : s = 170;
	{8'd124,8'd47} : s = 171;
	{8'd124,8'd48} : s = 172;
	{8'd124,8'd49} : s = 173;
	{8'd124,8'd50} : s = 174;
	{8'd124,8'd51} : s = 175;
	{8'd124,8'd52} : s = 176;
	{8'd124,8'd53} : s = 177;
	{8'd124,8'd54} : s = 178;
	{8'd124,8'd55} : s = 179;
	{8'd124,8'd56} : s = 180;
	{8'd124,8'd57} : s = 181;
	{8'd124,8'd58} : s = 182;
	{8'd124,8'd59} : s = 183;
	{8'd124,8'd60} : s = 184;
	{8'd124,8'd61} : s = 185;
	{8'd124,8'd62} : s = 186;
	{8'd124,8'd63} : s = 187;
	{8'd124,8'd64} : s = 188;
	{8'd124,8'd65} : s = 189;
	{8'd124,8'd66} : s = 190;
	{8'd124,8'd67} : s = 191;
	{8'd124,8'd68} : s = 192;
	{8'd124,8'd69} : s = 193;
	{8'd124,8'd70} : s = 194;
	{8'd124,8'd71} : s = 195;
	{8'd124,8'd72} : s = 196;
	{8'd124,8'd73} : s = 197;
	{8'd124,8'd74} : s = 198;
	{8'd124,8'd75} : s = 199;
	{8'd124,8'd76} : s = 200;
	{8'd124,8'd77} : s = 201;
	{8'd124,8'd78} : s = 202;
	{8'd124,8'd79} : s = 203;
	{8'd124,8'd80} : s = 204;
	{8'd124,8'd81} : s = 205;
	{8'd124,8'd82} : s = 206;
	{8'd124,8'd83} : s = 207;
	{8'd124,8'd84} : s = 208;
	{8'd124,8'd85} : s = 209;
	{8'd124,8'd86} : s = 210;
	{8'd124,8'd87} : s = 211;
	{8'd124,8'd88} : s = 212;
	{8'd124,8'd89} : s = 213;
	{8'd124,8'd90} : s = 214;
	{8'd124,8'd91} : s = 215;
	{8'd124,8'd92} : s = 216;
	{8'd124,8'd93} : s = 217;
	{8'd124,8'd94} : s = 218;
	{8'd124,8'd95} : s = 219;
	{8'd124,8'd96} : s = 220;
	{8'd124,8'd97} : s = 221;
	{8'd124,8'd98} : s = 222;
	{8'd124,8'd99} : s = 223;
	{8'd124,8'd100} : s = 224;
	{8'd124,8'd101} : s = 225;
	{8'd124,8'd102} : s = 226;
	{8'd124,8'd103} : s = 227;
	{8'd124,8'd104} : s = 228;
	{8'd124,8'd105} : s = 229;
	{8'd124,8'd106} : s = 230;
	{8'd124,8'd107} : s = 231;
	{8'd124,8'd108} : s = 232;
	{8'd124,8'd109} : s = 233;
	{8'd124,8'd110} : s = 234;
	{8'd124,8'd111} : s = 235;
	{8'd124,8'd112} : s = 236;
	{8'd124,8'd113} : s = 237;
	{8'd124,8'd114} : s = 238;
	{8'd124,8'd115} : s = 239;
	{8'd124,8'd116} : s = 240;
	{8'd124,8'd117} : s = 241;
	{8'd124,8'd118} : s = 242;
	{8'd124,8'd119} : s = 243;
	{8'd124,8'd120} : s = 244;
	{8'd124,8'd121} : s = 245;
	{8'd124,8'd122} : s = 246;
	{8'd124,8'd123} : s = 247;
	{8'd124,8'd124} : s = 248;
	{8'd124,8'd125} : s = 249;
	{8'd124,8'd126} : s = 250;
	{8'd124,8'd127} : s = 251;
	{8'd124,8'd128} : s = 252;
	{8'd124,8'd129} : s = 253;
	{8'd124,8'd130} : s = 254;
	{8'd124,8'd131} : s = 255;
	{8'd124,8'd132} : s = 256;
	{8'd124,8'd133} : s = 257;
	{8'd124,8'd134} : s = 258;
	{8'd124,8'd135} : s = 259;
	{8'd124,8'd136} : s = 260;
	{8'd124,8'd137} : s = 261;
	{8'd124,8'd138} : s = 262;
	{8'd124,8'd139} : s = 263;
	{8'd124,8'd140} : s = 264;
	{8'd124,8'd141} : s = 265;
	{8'd124,8'd142} : s = 266;
	{8'd124,8'd143} : s = 267;
	{8'd124,8'd144} : s = 268;
	{8'd124,8'd145} : s = 269;
	{8'd124,8'd146} : s = 270;
	{8'd124,8'd147} : s = 271;
	{8'd124,8'd148} : s = 272;
	{8'd124,8'd149} : s = 273;
	{8'd124,8'd150} : s = 274;
	{8'd124,8'd151} : s = 275;
	{8'd124,8'd152} : s = 276;
	{8'd124,8'd153} : s = 277;
	{8'd124,8'd154} : s = 278;
	{8'd124,8'd155} : s = 279;
	{8'd124,8'd156} : s = 280;
	{8'd124,8'd157} : s = 281;
	{8'd124,8'd158} : s = 282;
	{8'd124,8'd159} : s = 283;
	{8'd124,8'd160} : s = 284;
	{8'd124,8'd161} : s = 285;
	{8'd124,8'd162} : s = 286;
	{8'd124,8'd163} : s = 287;
	{8'd124,8'd164} : s = 288;
	{8'd124,8'd165} : s = 289;
	{8'd124,8'd166} : s = 290;
	{8'd124,8'd167} : s = 291;
	{8'd124,8'd168} : s = 292;
	{8'd124,8'd169} : s = 293;
	{8'd124,8'd170} : s = 294;
	{8'd124,8'd171} : s = 295;
	{8'd124,8'd172} : s = 296;
	{8'd124,8'd173} : s = 297;
	{8'd124,8'd174} : s = 298;
	{8'd124,8'd175} : s = 299;
	{8'd124,8'd176} : s = 300;
	{8'd124,8'd177} : s = 301;
	{8'd124,8'd178} : s = 302;
	{8'd124,8'd179} : s = 303;
	{8'd124,8'd180} : s = 304;
	{8'd124,8'd181} : s = 305;
	{8'd124,8'd182} : s = 306;
	{8'd124,8'd183} : s = 307;
	{8'd124,8'd184} : s = 308;
	{8'd124,8'd185} : s = 309;
	{8'd124,8'd186} : s = 310;
	{8'd124,8'd187} : s = 311;
	{8'd124,8'd188} : s = 312;
	{8'd124,8'd189} : s = 313;
	{8'd124,8'd190} : s = 314;
	{8'd124,8'd191} : s = 315;
	{8'd124,8'd192} : s = 316;
	{8'd124,8'd193} : s = 317;
	{8'd124,8'd194} : s = 318;
	{8'd124,8'd195} : s = 319;
	{8'd124,8'd196} : s = 320;
	{8'd124,8'd197} : s = 321;
	{8'd124,8'd198} : s = 322;
	{8'd124,8'd199} : s = 323;
	{8'd124,8'd200} : s = 324;
	{8'd124,8'd201} : s = 325;
	{8'd124,8'd202} : s = 326;
	{8'd124,8'd203} : s = 327;
	{8'd124,8'd204} : s = 328;
	{8'd124,8'd205} : s = 329;
	{8'd124,8'd206} : s = 330;
	{8'd124,8'd207} : s = 331;
	{8'd124,8'd208} : s = 332;
	{8'd124,8'd209} : s = 333;
	{8'd124,8'd210} : s = 334;
	{8'd124,8'd211} : s = 335;
	{8'd124,8'd212} : s = 336;
	{8'd124,8'd213} : s = 337;
	{8'd124,8'd214} : s = 338;
	{8'd124,8'd215} : s = 339;
	{8'd124,8'd216} : s = 340;
	{8'd124,8'd217} : s = 341;
	{8'd124,8'd218} : s = 342;
	{8'd124,8'd219} : s = 343;
	{8'd124,8'd220} : s = 344;
	{8'd124,8'd221} : s = 345;
	{8'd124,8'd222} : s = 346;
	{8'd124,8'd223} : s = 347;
	{8'd124,8'd224} : s = 348;
	{8'd124,8'd225} : s = 349;
	{8'd124,8'd226} : s = 350;
	{8'd124,8'd227} : s = 351;
	{8'd124,8'd228} : s = 352;
	{8'd124,8'd229} : s = 353;
	{8'd124,8'd230} : s = 354;
	{8'd124,8'd231} : s = 355;
	{8'd124,8'd232} : s = 356;
	{8'd124,8'd233} : s = 357;
	{8'd124,8'd234} : s = 358;
	{8'd124,8'd235} : s = 359;
	{8'd124,8'd236} : s = 360;
	{8'd124,8'd237} : s = 361;
	{8'd124,8'd238} : s = 362;
	{8'd124,8'd239} : s = 363;
	{8'd124,8'd240} : s = 364;
	{8'd124,8'd241} : s = 365;
	{8'd124,8'd242} : s = 366;
	{8'd124,8'd243} : s = 367;
	{8'd124,8'd244} : s = 368;
	{8'd124,8'd245} : s = 369;
	{8'd124,8'd246} : s = 370;
	{8'd124,8'd247} : s = 371;
	{8'd124,8'd248} : s = 372;
	{8'd124,8'd249} : s = 373;
	{8'd124,8'd250} : s = 374;
	{8'd124,8'd251} : s = 375;
	{8'd124,8'd252} : s = 376;
	{8'd124,8'd253} : s = 377;
	{8'd124,8'd254} : s = 378;
	{8'd124,8'd255} : s = 379;
	{8'd125,8'd0} : s = 125;
	{8'd125,8'd1} : s = 126;
	{8'd125,8'd2} : s = 127;
	{8'd125,8'd3} : s = 128;
	{8'd125,8'd4} : s = 129;
	{8'd125,8'd5} : s = 130;
	{8'd125,8'd6} : s = 131;
	{8'd125,8'd7} : s = 132;
	{8'd125,8'd8} : s = 133;
	{8'd125,8'd9} : s = 134;
	{8'd125,8'd10} : s = 135;
	{8'd125,8'd11} : s = 136;
	{8'd125,8'd12} : s = 137;
	{8'd125,8'd13} : s = 138;
	{8'd125,8'd14} : s = 139;
	{8'd125,8'd15} : s = 140;
	{8'd125,8'd16} : s = 141;
	{8'd125,8'd17} : s = 142;
	{8'd125,8'd18} : s = 143;
	{8'd125,8'd19} : s = 144;
	{8'd125,8'd20} : s = 145;
	{8'd125,8'd21} : s = 146;
	{8'd125,8'd22} : s = 147;
	{8'd125,8'd23} : s = 148;
	{8'd125,8'd24} : s = 149;
	{8'd125,8'd25} : s = 150;
	{8'd125,8'd26} : s = 151;
	{8'd125,8'd27} : s = 152;
	{8'd125,8'd28} : s = 153;
	{8'd125,8'd29} : s = 154;
	{8'd125,8'd30} : s = 155;
	{8'd125,8'd31} : s = 156;
	{8'd125,8'd32} : s = 157;
	{8'd125,8'd33} : s = 158;
	{8'd125,8'd34} : s = 159;
	{8'd125,8'd35} : s = 160;
	{8'd125,8'd36} : s = 161;
	{8'd125,8'd37} : s = 162;
	{8'd125,8'd38} : s = 163;
	{8'd125,8'd39} : s = 164;
	{8'd125,8'd40} : s = 165;
	{8'd125,8'd41} : s = 166;
	{8'd125,8'd42} : s = 167;
	{8'd125,8'd43} : s = 168;
	{8'd125,8'd44} : s = 169;
	{8'd125,8'd45} : s = 170;
	{8'd125,8'd46} : s = 171;
	{8'd125,8'd47} : s = 172;
	{8'd125,8'd48} : s = 173;
	{8'd125,8'd49} : s = 174;
	{8'd125,8'd50} : s = 175;
	{8'd125,8'd51} : s = 176;
	{8'd125,8'd52} : s = 177;
	{8'd125,8'd53} : s = 178;
	{8'd125,8'd54} : s = 179;
	{8'd125,8'd55} : s = 180;
	{8'd125,8'd56} : s = 181;
	{8'd125,8'd57} : s = 182;
	{8'd125,8'd58} : s = 183;
	{8'd125,8'd59} : s = 184;
	{8'd125,8'd60} : s = 185;
	{8'd125,8'd61} : s = 186;
	{8'd125,8'd62} : s = 187;
	{8'd125,8'd63} : s = 188;
	{8'd125,8'd64} : s = 189;
	{8'd125,8'd65} : s = 190;
	{8'd125,8'd66} : s = 191;
	{8'd125,8'd67} : s = 192;
	{8'd125,8'd68} : s = 193;
	{8'd125,8'd69} : s = 194;
	{8'd125,8'd70} : s = 195;
	{8'd125,8'd71} : s = 196;
	{8'd125,8'd72} : s = 197;
	{8'd125,8'd73} : s = 198;
	{8'd125,8'd74} : s = 199;
	{8'd125,8'd75} : s = 200;
	{8'd125,8'd76} : s = 201;
	{8'd125,8'd77} : s = 202;
	{8'd125,8'd78} : s = 203;
	{8'd125,8'd79} : s = 204;
	{8'd125,8'd80} : s = 205;
	{8'd125,8'd81} : s = 206;
	{8'd125,8'd82} : s = 207;
	{8'd125,8'd83} : s = 208;
	{8'd125,8'd84} : s = 209;
	{8'd125,8'd85} : s = 210;
	{8'd125,8'd86} : s = 211;
	{8'd125,8'd87} : s = 212;
	{8'd125,8'd88} : s = 213;
	{8'd125,8'd89} : s = 214;
	{8'd125,8'd90} : s = 215;
	{8'd125,8'd91} : s = 216;
	{8'd125,8'd92} : s = 217;
	{8'd125,8'd93} : s = 218;
	{8'd125,8'd94} : s = 219;
	{8'd125,8'd95} : s = 220;
	{8'd125,8'd96} : s = 221;
	{8'd125,8'd97} : s = 222;
	{8'd125,8'd98} : s = 223;
	{8'd125,8'd99} : s = 224;
	{8'd125,8'd100} : s = 225;
	{8'd125,8'd101} : s = 226;
	{8'd125,8'd102} : s = 227;
	{8'd125,8'd103} : s = 228;
	{8'd125,8'd104} : s = 229;
	{8'd125,8'd105} : s = 230;
	{8'd125,8'd106} : s = 231;
	{8'd125,8'd107} : s = 232;
	{8'd125,8'd108} : s = 233;
	{8'd125,8'd109} : s = 234;
	{8'd125,8'd110} : s = 235;
	{8'd125,8'd111} : s = 236;
	{8'd125,8'd112} : s = 237;
	{8'd125,8'd113} : s = 238;
	{8'd125,8'd114} : s = 239;
	{8'd125,8'd115} : s = 240;
	{8'd125,8'd116} : s = 241;
	{8'd125,8'd117} : s = 242;
	{8'd125,8'd118} : s = 243;
	{8'd125,8'd119} : s = 244;
	{8'd125,8'd120} : s = 245;
	{8'd125,8'd121} : s = 246;
	{8'd125,8'd122} : s = 247;
	{8'd125,8'd123} : s = 248;
	{8'd125,8'd124} : s = 249;
	{8'd125,8'd125} : s = 250;
	{8'd125,8'd126} : s = 251;
	{8'd125,8'd127} : s = 252;
	{8'd125,8'd128} : s = 253;
	{8'd125,8'd129} : s = 254;
	{8'd125,8'd130} : s = 255;
	{8'd125,8'd131} : s = 256;
	{8'd125,8'd132} : s = 257;
	{8'd125,8'd133} : s = 258;
	{8'd125,8'd134} : s = 259;
	{8'd125,8'd135} : s = 260;
	{8'd125,8'd136} : s = 261;
	{8'd125,8'd137} : s = 262;
	{8'd125,8'd138} : s = 263;
	{8'd125,8'd139} : s = 264;
	{8'd125,8'd140} : s = 265;
	{8'd125,8'd141} : s = 266;
	{8'd125,8'd142} : s = 267;
	{8'd125,8'd143} : s = 268;
	{8'd125,8'd144} : s = 269;
	{8'd125,8'd145} : s = 270;
	{8'd125,8'd146} : s = 271;
	{8'd125,8'd147} : s = 272;
	{8'd125,8'd148} : s = 273;
	{8'd125,8'd149} : s = 274;
	{8'd125,8'd150} : s = 275;
	{8'd125,8'd151} : s = 276;
	{8'd125,8'd152} : s = 277;
	{8'd125,8'd153} : s = 278;
	{8'd125,8'd154} : s = 279;
	{8'd125,8'd155} : s = 280;
	{8'd125,8'd156} : s = 281;
	{8'd125,8'd157} : s = 282;
	{8'd125,8'd158} : s = 283;
	{8'd125,8'd159} : s = 284;
	{8'd125,8'd160} : s = 285;
	{8'd125,8'd161} : s = 286;
	{8'd125,8'd162} : s = 287;
	{8'd125,8'd163} : s = 288;
	{8'd125,8'd164} : s = 289;
	{8'd125,8'd165} : s = 290;
	{8'd125,8'd166} : s = 291;
	{8'd125,8'd167} : s = 292;
	{8'd125,8'd168} : s = 293;
	{8'd125,8'd169} : s = 294;
	{8'd125,8'd170} : s = 295;
	{8'd125,8'd171} : s = 296;
	{8'd125,8'd172} : s = 297;
	{8'd125,8'd173} : s = 298;
	{8'd125,8'd174} : s = 299;
	{8'd125,8'd175} : s = 300;
	{8'd125,8'd176} : s = 301;
	{8'd125,8'd177} : s = 302;
	{8'd125,8'd178} : s = 303;
	{8'd125,8'd179} : s = 304;
	{8'd125,8'd180} : s = 305;
	{8'd125,8'd181} : s = 306;
	{8'd125,8'd182} : s = 307;
	{8'd125,8'd183} : s = 308;
	{8'd125,8'd184} : s = 309;
	{8'd125,8'd185} : s = 310;
	{8'd125,8'd186} : s = 311;
	{8'd125,8'd187} : s = 312;
	{8'd125,8'd188} : s = 313;
	{8'd125,8'd189} : s = 314;
	{8'd125,8'd190} : s = 315;
	{8'd125,8'd191} : s = 316;
	{8'd125,8'd192} : s = 317;
	{8'd125,8'd193} : s = 318;
	{8'd125,8'd194} : s = 319;
	{8'd125,8'd195} : s = 320;
	{8'd125,8'd196} : s = 321;
	{8'd125,8'd197} : s = 322;
	{8'd125,8'd198} : s = 323;
	{8'd125,8'd199} : s = 324;
	{8'd125,8'd200} : s = 325;
	{8'd125,8'd201} : s = 326;
	{8'd125,8'd202} : s = 327;
	{8'd125,8'd203} : s = 328;
	{8'd125,8'd204} : s = 329;
	{8'd125,8'd205} : s = 330;
	{8'd125,8'd206} : s = 331;
	{8'd125,8'd207} : s = 332;
	{8'd125,8'd208} : s = 333;
	{8'd125,8'd209} : s = 334;
	{8'd125,8'd210} : s = 335;
	{8'd125,8'd211} : s = 336;
	{8'd125,8'd212} : s = 337;
	{8'd125,8'd213} : s = 338;
	{8'd125,8'd214} : s = 339;
	{8'd125,8'd215} : s = 340;
	{8'd125,8'd216} : s = 341;
	{8'd125,8'd217} : s = 342;
	{8'd125,8'd218} : s = 343;
	{8'd125,8'd219} : s = 344;
	{8'd125,8'd220} : s = 345;
	{8'd125,8'd221} : s = 346;
	{8'd125,8'd222} : s = 347;
	{8'd125,8'd223} : s = 348;
	{8'd125,8'd224} : s = 349;
	{8'd125,8'd225} : s = 350;
	{8'd125,8'd226} : s = 351;
	{8'd125,8'd227} : s = 352;
	{8'd125,8'd228} : s = 353;
	{8'd125,8'd229} : s = 354;
	{8'd125,8'd230} : s = 355;
	{8'd125,8'd231} : s = 356;
	{8'd125,8'd232} : s = 357;
	{8'd125,8'd233} : s = 358;
	{8'd125,8'd234} : s = 359;
	{8'd125,8'd235} : s = 360;
	{8'd125,8'd236} : s = 361;
	{8'd125,8'd237} : s = 362;
	{8'd125,8'd238} : s = 363;
	{8'd125,8'd239} : s = 364;
	{8'd125,8'd240} : s = 365;
	{8'd125,8'd241} : s = 366;
	{8'd125,8'd242} : s = 367;
	{8'd125,8'd243} : s = 368;
	{8'd125,8'd244} : s = 369;
	{8'd125,8'd245} : s = 370;
	{8'd125,8'd246} : s = 371;
	{8'd125,8'd247} : s = 372;
	{8'd125,8'd248} : s = 373;
	{8'd125,8'd249} : s = 374;
	{8'd125,8'd250} : s = 375;
	{8'd125,8'd251} : s = 376;
	{8'd125,8'd252} : s = 377;
	{8'd125,8'd253} : s = 378;
	{8'd125,8'd254} : s = 379;
	{8'd125,8'd255} : s = 380;
	{8'd126,8'd0} : s = 126;
	{8'd126,8'd1} : s = 127;
	{8'd126,8'd2} : s = 128;
	{8'd126,8'd3} : s = 129;
	{8'd126,8'd4} : s = 130;
	{8'd126,8'd5} : s = 131;
	{8'd126,8'd6} : s = 132;
	{8'd126,8'd7} : s = 133;
	{8'd126,8'd8} : s = 134;
	{8'd126,8'd9} : s = 135;
	{8'd126,8'd10} : s = 136;
	{8'd126,8'd11} : s = 137;
	{8'd126,8'd12} : s = 138;
	{8'd126,8'd13} : s = 139;
	{8'd126,8'd14} : s = 140;
	{8'd126,8'd15} : s = 141;
	{8'd126,8'd16} : s = 142;
	{8'd126,8'd17} : s = 143;
	{8'd126,8'd18} : s = 144;
	{8'd126,8'd19} : s = 145;
	{8'd126,8'd20} : s = 146;
	{8'd126,8'd21} : s = 147;
	{8'd126,8'd22} : s = 148;
	{8'd126,8'd23} : s = 149;
	{8'd126,8'd24} : s = 150;
	{8'd126,8'd25} : s = 151;
	{8'd126,8'd26} : s = 152;
	{8'd126,8'd27} : s = 153;
	{8'd126,8'd28} : s = 154;
	{8'd126,8'd29} : s = 155;
	{8'd126,8'd30} : s = 156;
	{8'd126,8'd31} : s = 157;
	{8'd126,8'd32} : s = 158;
	{8'd126,8'd33} : s = 159;
	{8'd126,8'd34} : s = 160;
	{8'd126,8'd35} : s = 161;
	{8'd126,8'd36} : s = 162;
	{8'd126,8'd37} : s = 163;
	{8'd126,8'd38} : s = 164;
	{8'd126,8'd39} : s = 165;
	{8'd126,8'd40} : s = 166;
	{8'd126,8'd41} : s = 167;
	{8'd126,8'd42} : s = 168;
	{8'd126,8'd43} : s = 169;
	{8'd126,8'd44} : s = 170;
	{8'd126,8'd45} : s = 171;
	{8'd126,8'd46} : s = 172;
	{8'd126,8'd47} : s = 173;
	{8'd126,8'd48} : s = 174;
	{8'd126,8'd49} : s = 175;
	{8'd126,8'd50} : s = 176;
	{8'd126,8'd51} : s = 177;
	{8'd126,8'd52} : s = 178;
	{8'd126,8'd53} : s = 179;
	{8'd126,8'd54} : s = 180;
	{8'd126,8'd55} : s = 181;
	{8'd126,8'd56} : s = 182;
	{8'd126,8'd57} : s = 183;
	{8'd126,8'd58} : s = 184;
	{8'd126,8'd59} : s = 185;
	{8'd126,8'd60} : s = 186;
	{8'd126,8'd61} : s = 187;
	{8'd126,8'd62} : s = 188;
	{8'd126,8'd63} : s = 189;
	{8'd126,8'd64} : s = 190;
	{8'd126,8'd65} : s = 191;
	{8'd126,8'd66} : s = 192;
	{8'd126,8'd67} : s = 193;
	{8'd126,8'd68} : s = 194;
	{8'd126,8'd69} : s = 195;
	{8'd126,8'd70} : s = 196;
	{8'd126,8'd71} : s = 197;
	{8'd126,8'd72} : s = 198;
	{8'd126,8'd73} : s = 199;
	{8'd126,8'd74} : s = 200;
	{8'd126,8'd75} : s = 201;
	{8'd126,8'd76} : s = 202;
	{8'd126,8'd77} : s = 203;
	{8'd126,8'd78} : s = 204;
	{8'd126,8'd79} : s = 205;
	{8'd126,8'd80} : s = 206;
	{8'd126,8'd81} : s = 207;
	{8'd126,8'd82} : s = 208;
	{8'd126,8'd83} : s = 209;
	{8'd126,8'd84} : s = 210;
	{8'd126,8'd85} : s = 211;
	{8'd126,8'd86} : s = 212;
	{8'd126,8'd87} : s = 213;
	{8'd126,8'd88} : s = 214;
	{8'd126,8'd89} : s = 215;
	{8'd126,8'd90} : s = 216;
	{8'd126,8'd91} : s = 217;
	{8'd126,8'd92} : s = 218;
	{8'd126,8'd93} : s = 219;
	{8'd126,8'd94} : s = 220;
	{8'd126,8'd95} : s = 221;
	{8'd126,8'd96} : s = 222;
	{8'd126,8'd97} : s = 223;
	{8'd126,8'd98} : s = 224;
	{8'd126,8'd99} : s = 225;
	{8'd126,8'd100} : s = 226;
	{8'd126,8'd101} : s = 227;
	{8'd126,8'd102} : s = 228;
	{8'd126,8'd103} : s = 229;
	{8'd126,8'd104} : s = 230;
	{8'd126,8'd105} : s = 231;
	{8'd126,8'd106} : s = 232;
	{8'd126,8'd107} : s = 233;
	{8'd126,8'd108} : s = 234;
	{8'd126,8'd109} : s = 235;
	{8'd126,8'd110} : s = 236;
	{8'd126,8'd111} : s = 237;
	{8'd126,8'd112} : s = 238;
	{8'd126,8'd113} : s = 239;
	{8'd126,8'd114} : s = 240;
	{8'd126,8'd115} : s = 241;
	{8'd126,8'd116} : s = 242;
	{8'd126,8'd117} : s = 243;
	{8'd126,8'd118} : s = 244;
	{8'd126,8'd119} : s = 245;
	{8'd126,8'd120} : s = 246;
	{8'd126,8'd121} : s = 247;
	{8'd126,8'd122} : s = 248;
	{8'd126,8'd123} : s = 249;
	{8'd126,8'd124} : s = 250;
	{8'd126,8'd125} : s = 251;
	{8'd126,8'd126} : s = 252;
	{8'd126,8'd127} : s = 253;
	{8'd126,8'd128} : s = 254;
	{8'd126,8'd129} : s = 255;
	{8'd126,8'd130} : s = 256;
	{8'd126,8'd131} : s = 257;
	{8'd126,8'd132} : s = 258;
	{8'd126,8'd133} : s = 259;
	{8'd126,8'd134} : s = 260;
	{8'd126,8'd135} : s = 261;
	{8'd126,8'd136} : s = 262;
	{8'd126,8'd137} : s = 263;
	{8'd126,8'd138} : s = 264;
	{8'd126,8'd139} : s = 265;
	{8'd126,8'd140} : s = 266;
	{8'd126,8'd141} : s = 267;
	{8'd126,8'd142} : s = 268;
	{8'd126,8'd143} : s = 269;
	{8'd126,8'd144} : s = 270;
	{8'd126,8'd145} : s = 271;
	{8'd126,8'd146} : s = 272;
	{8'd126,8'd147} : s = 273;
	{8'd126,8'd148} : s = 274;
	{8'd126,8'd149} : s = 275;
	{8'd126,8'd150} : s = 276;
	{8'd126,8'd151} : s = 277;
	{8'd126,8'd152} : s = 278;
	{8'd126,8'd153} : s = 279;
	{8'd126,8'd154} : s = 280;
	{8'd126,8'd155} : s = 281;
	{8'd126,8'd156} : s = 282;
	{8'd126,8'd157} : s = 283;
	{8'd126,8'd158} : s = 284;
	{8'd126,8'd159} : s = 285;
	{8'd126,8'd160} : s = 286;
	{8'd126,8'd161} : s = 287;
	{8'd126,8'd162} : s = 288;
	{8'd126,8'd163} : s = 289;
	{8'd126,8'd164} : s = 290;
	{8'd126,8'd165} : s = 291;
	{8'd126,8'd166} : s = 292;
	{8'd126,8'd167} : s = 293;
	{8'd126,8'd168} : s = 294;
	{8'd126,8'd169} : s = 295;
	{8'd126,8'd170} : s = 296;
	{8'd126,8'd171} : s = 297;
	{8'd126,8'd172} : s = 298;
	{8'd126,8'd173} : s = 299;
	{8'd126,8'd174} : s = 300;
	{8'd126,8'd175} : s = 301;
	{8'd126,8'd176} : s = 302;
	{8'd126,8'd177} : s = 303;
	{8'd126,8'd178} : s = 304;
	{8'd126,8'd179} : s = 305;
	{8'd126,8'd180} : s = 306;
	{8'd126,8'd181} : s = 307;
	{8'd126,8'd182} : s = 308;
	{8'd126,8'd183} : s = 309;
	{8'd126,8'd184} : s = 310;
	{8'd126,8'd185} : s = 311;
	{8'd126,8'd186} : s = 312;
	{8'd126,8'd187} : s = 313;
	{8'd126,8'd188} : s = 314;
	{8'd126,8'd189} : s = 315;
	{8'd126,8'd190} : s = 316;
	{8'd126,8'd191} : s = 317;
	{8'd126,8'd192} : s = 318;
	{8'd126,8'd193} : s = 319;
	{8'd126,8'd194} : s = 320;
	{8'd126,8'd195} : s = 321;
	{8'd126,8'd196} : s = 322;
	{8'd126,8'd197} : s = 323;
	{8'd126,8'd198} : s = 324;
	{8'd126,8'd199} : s = 325;
	{8'd126,8'd200} : s = 326;
	{8'd126,8'd201} : s = 327;
	{8'd126,8'd202} : s = 328;
	{8'd126,8'd203} : s = 329;
	{8'd126,8'd204} : s = 330;
	{8'd126,8'd205} : s = 331;
	{8'd126,8'd206} : s = 332;
	{8'd126,8'd207} : s = 333;
	{8'd126,8'd208} : s = 334;
	{8'd126,8'd209} : s = 335;
	{8'd126,8'd210} : s = 336;
	{8'd126,8'd211} : s = 337;
	{8'd126,8'd212} : s = 338;
	{8'd126,8'd213} : s = 339;
	{8'd126,8'd214} : s = 340;
	{8'd126,8'd215} : s = 341;
	{8'd126,8'd216} : s = 342;
	{8'd126,8'd217} : s = 343;
	{8'd126,8'd218} : s = 344;
	{8'd126,8'd219} : s = 345;
	{8'd126,8'd220} : s = 346;
	{8'd126,8'd221} : s = 347;
	{8'd126,8'd222} : s = 348;
	{8'd126,8'd223} : s = 349;
	{8'd126,8'd224} : s = 350;
	{8'd126,8'd225} : s = 351;
	{8'd126,8'd226} : s = 352;
	{8'd126,8'd227} : s = 353;
	{8'd126,8'd228} : s = 354;
	{8'd126,8'd229} : s = 355;
	{8'd126,8'd230} : s = 356;
	{8'd126,8'd231} : s = 357;
	{8'd126,8'd232} : s = 358;
	{8'd126,8'd233} : s = 359;
	{8'd126,8'd234} : s = 360;
	{8'd126,8'd235} : s = 361;
	{8'd126,8'd236} : s = 362;
	{8'd126,8'd237} : s = 363;
	{8'd126,8'd238} : s = 364;
	{8'd126,8'd239} : s = 365;
	{8'd126,8'd240} : s = 366;
	{8'd126,8'd241} : s = 367;
	{8'd126,8'd242} : s = 368;
	{8'd126,8'd243} : s = 369;
	{8'd126,8'd244} : s = 370;
	{8'd126,8'd245} : s = 371;
	{8'd126,8'd246} : s = 372;
	{8'd126,8'd247} : s = 373;
	{8'd126,8'd248} : s = 374;
	{8'd126,8'd249} : s = 375;
	{8'd126,8'd250} : s = 376;
	{8'd126,8'd251} : s = 377;
	{8'd126,8'd252} : s = 378;
	{8'd126,8'd253} : s = 379;
	{8'd126,8'd254} : s = 380;
	{8'd126,8'd255} : s = 381;
	{8'd127,8'd0} : s = 127;
	{8'd127,8'd1} : s = 128;
	{8'd127,8'd2} : s = 129;
	{8'd127,8'd3} : s = 130;
	{8'd127,8'd4} : s = 131;
	{8'd127,8'd5} : s = 132;
	{8'd127,8'd6} : s = 133;
	{8'd127,8'd7} : s = 134;
	{8'd127,8'd8} : s = 135;
	{8'd127,8'd9} : s = 136;
	{8'd127,8'd10} : s = 137;
	{8'd127,8'd11} : s = 138;
	{8'd127,8'd12} : s = 139;
	{8'd127,8'd13} : s = 140;
	{8'd127,8'd14} : s = 141;
	{8'd127,8'd15} : s = 142;
	{8'd127,8'd16} : s = 143;
	{8'd127,8'd17} : s = 144;
	{8'd127,8'd18} : s = 145;
	{8'd127,8'd19} : s = 146;
	{8'd127,8'd20} : s = 147;
	{8'd127,8'd21} : s = 148;
	{8'd127,8'd22} : s = 149;
	{8'd127,8'd23} : s = 150;
	{8'd127,8'd24} : s = 151;
	{8'd127,8'd25} : s = 152;
	{8'd127,8'd26} : s = 153;
	{8'd127,8'd27} : s = 154;
	{8'd127,8'd28} : s = 155;
	{8'd127,8'd29} : s = 156;
	{8'd127,8'd30} : s = 157;
	{8'd127,8'd31} : s = 158;
	{8'd127,8'd32} : s = 159;
	{8'd127,8'd33} : s = 160;
	{8'd127,8'd34} : s = 161;
	{8'd127,8'd35} : s = 162;
	{8'd127,8'd36} : s = 163;
	{8'd127,8'd37} : s = 164;
	{8'd127,8'd38} : s = 165;
	{8'd127,8'd39} : s = 166;
	{8'd127,8'd40} : s = 167;
	{8'd127,8'd41} : s = 168;
	{8'd127,8'd42} : s = 169;
	{8'd127,8'd43} : s = 170;
	{8'd127,8'd44} : s = 171;
	{8'd127,8'd45} : s = 172;
	{8'd127,8'd46} : s = 173;
	{8'd127,8'd47} : s = 174;
	{8'd127,8'd48} : s = 175;
	{8'd127,8'd49} : s = 176;
	{8'd127,8'd50} : s = 177;
	{8'd127,8'd51} : s = 178;
	{8'd127,8'd52} : s = 179;
	{8'd127,8'd53} : s = 180;
	{8'd127,8'd54} : s = 181;
	{8'd127,8'd55} : s = 182;
	{8'd127,8'd56} : s = 183;
	{8'd127,8'd57} : s = 184;
	{8'd127,8'd58} : s = 185;
	{8'd127,8'd59} : s = 186;
	{8'd127,8'd60} : s = 187;
	{8'd127,8'd61} : s = 188;
	{8'd127,8'd62} : s = 189;
	{8'd127,8'd63} : s = 190;
	{8'd127,8'd64} : s = 191;
	{8'd127,8'd65} : s = 192;
	{8'd127,8'd66} : s = 193;
	{8'd127,8'd67} : s = 194;
	{8'd127,8'd68} : s = 195;
	{8'd127,8'd69} : s = 196;
	{8'd127,8'd70} : s = 197;
	{8'd127,8'd71} : s = 198;
	{8'd127,8'd72} : s = 199;
	{8'd127,8'd73} : s = 200;
	{8'd127,8'd74} : s = 201;
	{8'd127,8'd75} : s = 202;
	{8'd127,8'd76} : s = 203;
	{8'd127,8'd77} : s = 204;
	{8'd127,8'd78} : s = 205;
	{8'd127,8'd79} : s = 206;
	{8'd127,8'd80} : s = 207;
	{8'd127,8'd81} : s = 208;
	{8'd127,8'd82} : s = 209;
	{8'd127,8'd83} : s = 210;
	{8'd127,8'd84} : s = 211;
	{8'd127,8'd85} : s = 212;
	{8'd127,8'd86} : s = 213;
	{8'd127,8'd87} : s = 214;
	{8'd127,8'd88} : s = 215;
	{8'd127,8'd89} : s = 216;
	{8'd127,8'd90} : s = 217;
	{8'd127,8'd91} : s = 218;
	{8'd127,8'd92} : s = 219;
	{8'd127,8'd93} : s = 220;
	{8'd127,8'd94} : s = 221;
	{8'd127,8'd95} : s = 222;
	{8'd127,8'd96} : s = 223;
	{8'd127,8'd97} : s = 224;
	{8'd127,8'd98} : s = 225;
	{8'd127,8'd99} : s = 226;
	{8'd127,8'd100} : s = 227;
	{8'd127,8'd101} : s = 228;
	{8'd127,8'd102} : s = 229;
	{8'd127,8'd103} : s = 230;
	{8'd127,8'd104} : s = 231;
	{8'd127,8'd105} : s = 232;
	{8'd127,8'd106} : s = 233;
	{8'd127,8'd107} : s = 234;
	{8'd127,8'd108} : s = 235;
	{8'd127,8'd109} : s = 236;
	{8'd127,8'd110} : s = 237;
	{8'd127,8'd111} : s = 238;
	{8'd127,8'd112} : s = 239;
	{8'd127,8'd113} : s = 240;
	{8'd127,8'd114} : s = 241;
	{8'd127,8'd115} : s = 242;
	{8'd127,8'd116} : s = 243;
	{8'd127,8'd117} : s = 244;
	{8'd127,8'd118} : s = 245;
	{8'd127,8'd119} : s = 246;
	{8'd127,8'd120} : s = 247;
	{8'd127,8'd121} : s = 248;
	{8'd127,8'd122} : s = 249;
	{8'd127,8'd123} : s = 250;
	{8'd127,8'd124} : s = 251;
	{8'd127,8'd125} : s = 252;
	{8'd127,8'd126} : s = 253;
	{8'd127,8'd127} : s = 254;
	{8'd127,8'd128} : s = 255;
	{8'd127,8'd129} : s = 256;
	{8'd127,8'd130} : s = 257;
	{8'd127,8'd131} : s = 258;
	{8'd127,8'd132} : s = 259;
	{8'd127,8'd133} : s = 260;
	{8'd127,8'd134} : s = 261;
	{8'd127,8'd135} : s = 262;
	{8'd127,8'd136} : s = 263;
	{8'd127,8'd137} : s = 264;
	{8'd127,8'd138} : s = 265;
	{8'd127,8'd139} : s = 266;
	{8'd127,8'd140} : s = 267;
	{8'd127,8'd141} : s = 268;
	{8'd127,8'd142} : s = 269;
	{8'd127,8'd143} : s = 270;
	{8'd127,8'd144} : s = 271;
	{8'd127,8'd145} : s = 272;
	{8'd127,8'd146} : s = 273;
	{8'd127,8'd147} : s = 274;
	{8'd127,8'd148} : s = 275;
	{8'd127,8'd149} : s = 276;
	{8'd127,8'd150} : s = 277;
	{8'd127,8'd151} : s = 278;
	{8'd127,8'd152} : s = 279;
	{8'd127,8'd153} : s = 280;
	{8'd127,8'd154} : s = 281;
	{8'd127,8'd155} : s = 282;
	{8'd127,8'd156} : s = 283;
	{8'd127,8'd157} : s = 284;
	{8'd127,8'd158} : s = 285;
	{8'd127,8'd159} : s = 286;
	{8'd127,8'd160} : s = 287;
	{8'd127,8'd161} : s = 288;
	{8'd127,8'd162} : s = 289;
	{8'd127,8'd163} : s = 290;
	{8'd127,8'd164} : s = 291;
	{8'd127,8'd165} : s = 292;
	{8'd127,8'd166} : s = 293;
	{8'd127,8'd167} : s = 294;
	{8'd127,8'd168} : s = 295;
	{8'd127,8'd169} : s = 296;
	{8'd127,8'd170} : s = 297;
	{8'd127,8'd171} : s = 298;
	{8'd127,8'd172} : s = 299;
	{8'd127,8'd173} : s = 300;
	{8'd127,8'd174} : s = 301;
	{8'd127,8'd175} : s = 302;
	{8'd127,8'd176} : s = 303;
	{8'd127,8'd177} : s = 304;
	{8'd127,8'd178} : s = 305;
	{8'd127,8'd179} : s = 306;
	{8'd127,8'd180} : s = 307;
	{8'd127,8'd181} : s = 308;
	{8'd127,8'd182} : s = 309;
	{8'd127,8'd183} : s = 310;
	{8'd127,8'd184} : s = 311;
	{8'd127,8'd185} : s = 312;
	{8'd127,8'd186} : s = 313;
	{8'd127,8'd187} : s = 314;
	{8'd127,8'd188} : s = 315;
	{8'd127,8'd189} : s = 316;
	{8'd127,8'd190} : s = 317;
	{8'd127,8'd191} : s = 318;
	{8'd127,8'd192} : s = 319;
	{8'd127,8'd193} : s = 320;
	{8'd127,8'd194} : s = 321;
	{8'd127,8'd195} : s = 322;
	{8'd127,8'd196} : s = 323;
	{8'd127,8'd197} : s = 324;
	{8'd127,8'd198} : s = 325;
	{8'd127,8'd199} : s = 326;
	{8'd127,8'd200} : s = 327;
	{8'd127,8'd201} : s = 328;
	{8'd127,8'd202} : s = 329;
	{8'd127,8'd203} : s = 330;
	{8'd127,8'd204} : s = 331;
	{8'd127,8'd205} : s = 332;
	{8'd127,8'd206} : s = 333;
	{8'd127,8'd207} : s = 334;
	{8'd127,8'd208} : s = 335;
	{8'd127,8'd209} : s = 336;
	{8'd127,8'd210} : s = 337;
	{8'd127,8'd211} : s = 338;
	{8'd127,8'd212} : s = 339;
	{8'd127,8'd213} : s = 340;
	{8'd127,8'd214} : s = 341;
	{8'd127,8'd215} : s = 342;
	{8'd127,8'd216} : s = 343;
	{8'd127,8'd217} : s = 344;
	{8'd127,8'd218} : s = 345;
	{8'd127,8'd219} : s = 346;
	{8'd127,8'd220} : s = 347;
	{8'd127,8'd221} : s = 348;
	{8'd127,8'd222} : s = 349;
	{8'd127,8'd223} : s = 350;
	{8'd127,8'd224} : s = 351;
	{8'd127,8'd225} : s = 352;
	{8'd127,8'd226} : s = 353;
	{8'd127,8'd227} : s = 354;
	{8'd127,8'd228} : s = 355;
	{8'd127,8'd229} : s = 356;
	{8'd127,8'd230} : s = 357;
	{8'd127,8'd231} : s = 358;
	{8'd127,8'd232} : s = 359;
	{8'd127,8'd233} : s = 360;
	{8'd127,8'd234} : s = 361;
	{8'd127,8'd235} : s = 362;
	{8'd127,8'd236} : s = 363;
	{8'd127,8'd237} : s = 364;
	{8'd127,8'd238} : s = 365;
	{8'd127,8'd239} : s = 366;
	{8'd127,8'd240} : s = 367;
	{8'd127,8'd241} : s = 368;
	{8'd127,8'd242} : s = 369;
	{8'd127,8'd243} : s = 370;
	{8'd127,8'd244} : s = 371;
	{8'd127,8'd245} : s = 372;
	{8'd127,8'd246} : s = 373;
	{8'd127,8'd247} : s = 374;
	{8'd127,8'd248} : s = 375;
	{8'd127,8'd249} : s = 376;
	{8'd127,8'd250} : s = 377;
	{8'd127,8'd251} : s = 378;
	{8'd127,8'd252} : s = 379;
	{8'd127,8'd253} : s = 380;
	{8'd127,8'd254} : s = 381;
	{8'd127,8'd255} : s = 382;
	{8'd128,8'd0} : s = 128;
	{8'd128,8'd1} : s = 129;
	{8'd128,8'd2} : s = 130;
	{8'd128,8'd3} : s = 131;
	{8'd128,8'd4} : s = 132;
	{8'd128,8'd5} : s = 133;
	{8'd128,8'd6} : s = 134;
	{8'd128,8'd7} : s = 135;
	{8'd128,8'd8} : s = 136;
	{8'd128,8'd9} : s = 137;
	{8'd128,8'd10} : s = 138;
	{8'd128,8'd11} : s = 139;
	{8'd128,8'd12} : s = 140;
	{8'd128,8'd13} : s = 141;
	{8'd128,8'd14} : s = 142;
	{8'd128,8'd15} : s = 143;
	{8'd128,8'd16} : s = 144;
	{8'd128,8'd17} : s = 145;
	{8'd128,8'd18} : s = 146;
	{8'd128,8'd19} : s = 147;
	{8'd128,8'd20} : s = 148;
	{8'd128,8'd21} : s = 149;
	{8'd128,8'd22} : s = 150;
	{8'd128,8'd23} : s = 151;
	{8'd128,8'd24} : s = 152;
	{8'd128,8'd25} : s = 153;
	{8'd128,8'd26} : s = 154;
	{8'd128,8'd27} : s = 155;
	{8'd128,8'd28} : s = 156;
	{8'd128,8'd29} : s = 157;
	{8'd128,8'd30} : s = 158;
	{8'd128,8'd31} : s = 159;
	{8'd128,8'd32} : s = 160;
	{8'd128,8'd33} : s = 161;
	{8'd128,8'd34} : s = 162;
	{8'd128,8'd35} : s = 163;
	{8'd128,8'd36} : s = 164;
	{8'd128,8'd37} : s = 165;
	{8'd128,8'd38} : s = 166;
	{8'd128,8'd39} : s = 167;
	{8'd128,8'd40} : s = 168;
	{8'd128,8'd41} : s = 169;
	{8'd128,8'd42} : s = 170;
	{8'd128,8'd43} : s = 171;
	{8'd128,8'd44} : s = 172;
	{8'd128,8'd45} : s = 173;
	{8'd128,8'd46} : s = 174;
	{8'd128,8'd47} : s = 175;
	{8'd128,8'd48} : s = 176;
	{8'd128,8'd49} : s = 177;
	{8'd128,8'd50} : s = 178;
	{8'd128,8'd51} : s = 179;
	{8'd128,8'd52} : s = 180;
	{8'd128,8'd53} : s = 181;
	{8'd128,8'd54} : s = 182;
	{8'd128,8'd55} : s = 183;
	{8'd128,8'd56} : s = 184;
	{8'd128,8'd57} : s = 185;
	{8'd128,8'd58} : s = 186;
	{8'd128,8'd59} : s = 187;
	{8'd128,8'd60} : s = 188;
	{8'd128,8'd61} : s = 189;
	{8'd128,8'd62} : s = 190;
	{8'd128,8'd63} : s = 191;
	{8'd128,8'd64} : s = 192;
	{8'd128,8'd65} : s = 193;
	{8'd128,8'd66} : s = 194;
	{8'd128,8'd67} : s = 195;
	{8'd128,8'd68} : s = 196;
	{8'd128,8'd69} : s = 197;
	{8'd128,8'd70} : s = 198;
	{8'd128,8'd71} : s = 199;
	{8'd128,8'd72} : s = 200;
	{8'd128,8'd73} : s = 201;
	{8'd128,8'd74} : s = 202;
	{8'd128,8'd75} : s = 203;
	{8'd128,8'd76} : s = 204;
	{8'd128,8'd77} : s = 205;
	{8'd128,8'd78} : s = 206;
	{8'd128,8'd79} : s = 207;
	{8'd128,8'd80} : s = 208;
	{8'd128,8'd81} : s = 209;
	{8'd128,8'd82} : s = 210;
	{8'd128,8'd83} : s = 211;
	{8'd128,8'd84} : s = 212;
	{8'd128,8'd85} : s = 213;
	{8'd128,8'd86} : s = 214;
	{8'd128,8'd87} : s = 215;
	{8'd128,8'd88} : s = 216;
	{8'd128,8'd89} : s = 217;
	{8'd128,8'd90} : s = 218;
	{8'd128,8'd91} : s = 219;
	{8'd128,8'd92} : s = 220;
	{8'd128,8'd93} : s = 221;
	{8'd128,8'd94} : s = 222;
	{8'd128,8'd95} : s = 223;
	{8'd128,8'd96} : s = 224;
	{8'd128,8'd97} : s = 225;
	{8'd128,8'd98} : s = 226;
	{8'd128,8'd99} : s = 227;
	{8'd128,8'd100} : s = 228;
	{8'd128,8'd101} : s = 229;
	{8'd128,8'd102} : s = 230;
	{8'd128,8'd103} : s = 231;
	{8'd128,8'd104} : s = 232;
	{8'd128,8'd105} : s = 233;
	{8'd128,8'd106} : s = 234;
	{8'd128,8'd107} : s = 235;
	{8'd128,8'd108} : s = 236;
	{8'd128,8'd109} : s = 237;
	{8'd128,8'd110} : s = 238;
	{8'd128,8'd111} : s = 239;
	{8'd128,8'd112} : s = 240;
	{8'd128,8'd113} : s = 241;
	{8'd128,8'd114} : s = 242;
	{8'd128,8'd115} : s = 243;
	{8'd128,8'd116} : s = 244;
	{8'd128,8'd117} : s = 245;
	{8'd128,8'd118} : s = 246;
	{8'd128,8'd119} : s = 247;
	{8'd128,8'd120} : s = 248;
	{8'd128,8'd121} : s = 249;
	{8'd128,8'd122} : s = 250;
	{8'd128,8'd123} : s = 251;
	{8'd128,8'd124} : s = 252;
	{8'd128,8'd125} : s = 253;
	{8'd128,8'd126} : s = 254;
	{8'd128,8'd127} : s = 255;
	{8'd128,8'd128} : s = 256;
	{8'd128,8'd129} : s = 257;
	{8'd128,8'd130} : s = 258;
	{8'd128,8'd131} : s = 259;
	{8'd128,8'd132} : s = 260;
	{8'd128,8'd133} : s = 261;
	{8'd128,8'd134} : s = 262;
	{8'd128,8'd135} : s = 263;
	{8'd128,8'd136} : s = 264;
	{8'd128,8'd137} : s = 265;
	{8'd128,8'd138} : s = 266;
	{8'd128,8'd139} : s = 267;
	{8'd128,8'd140} : s = 268;
	{8'd128,8'd141} : s = 269;
	{8'd128,8'd142} : s = 270;
	{8'd128,8'd143} : s = 271;
	{8'd128,8'd144} : s = 272;
	{8'd128,8'd145} : s = 273;
	{8'd128,8'd146} : s = 274;
	{8'd128,8'd147} : s = 275;
	{8'd128,8'd148} : s = 276;
	{8'd128,8'd149} : s = 277;
	{8'd128,8'd150} : s = 278;
	{8'd128,8'd151} : s = 279;
	{8'd128,8'd152} : s = 280;
	{8'd128,8'd153} : s = 281;
	{8'd128,8'd154} : s = 282;
	{8'd128,8'd155} : s = 283;
	{8'd128,8'd156} : s = 284;
	{8'd128,8'd157} : s = 285;
	{8'd128,8'd158} : s = 286;
	{8'd128,8'd159} : s = 287;
	{8'd128,8'd160} : s = 288;
	{8'd128,8'd161} : s = 289;
	{8'd128,8'd162} : s = 290;
	{8'd128,8'd163} : s = 291;
	{8'd128,8'd164} : s = 292;
	{8'd128,8'd165} : s = 293;
	{8'd128,8'd166} : s = 294;
	{8'd128,8'd167} : s = 295;
	{8'd128,8'd168} : s = 296;
	{8'd128,8'd169} : s = 297;
	{8'd128,8'd170} : s = 298;
	{8'd128,8'd171} : s = 299;
	{8'd128,8'd172} : s = 300;
	{8'd128,8'd173} : s = 301;
	{8'd128,8'd174} : s = 302;
	{8'd128,8'd175} : s = 303;
	{8'd128,8'd176} : s = 304;
	{8'd128,8'd177} : s = 305;
	{8'd128,8'd178} : s = 306;
	{8'd128,8'd179} : s = 307;
	{8'd128,8'd180} : s = 308;
	{8'd128,8'd181} : s = 309;
	{8'd128,8'd182} : s = 310;
	{8'd128,8'd183} : s = 311;
	{8'd128,8'd184} : s = 312;
	{8'd128,8'd185} : s = 313;
	{8'd128,8'd186} : s = 314;
	{8'd128,8'd187} : s = 315;
	{8'd128,8'd188} : s = 316;
	{8'd128,8'd189} : s = 317;
	{8'd128,8'd190} : s = 318;
	{8'd128,8'd191} : s = 319;
	{8'd128,8'd192} : s = 320;
	{8'd128,8'd193} : s = 321;
	{8'd128,8'd194} : s = 322;
	{8'd128,8'd195} : s = 323;
	{8'd128,8'd196} : s = 324;
	{8'd128,8'd197} : s = 325;
	{8'd128,8'd198} : s = 326;
	{8'd128,8'd199} : s = 327;
	{8'd128,8'd200} : s = 328;
	{8'd128,8'd201} : s = 329;
	{8'd128,8'd202} : s = 330;
	{8'd128,8'd203} : s = 331;
	{8'd128,8'd204} : s = 332;
	{8'd128,8'd205} : s = 333;
	{8'd128,8'd206} : s = 334;
	{8'd128,8'd207} : s = 335;
	{8'd128,8'd208} : s = 336;
	{8'd128,8'd209} : s = 337;
	{8'd128,8'd210} : s = 338;
	{8'd128,8'd211} : s = 339;
	{8'd128,8'd212} : s = 340;
	{8'd128,8'd213} : s = 341;
	{8'd128,8'd214} : s = 342;
	{8'd128,8'd215} : s = 343;
	{8'd128,8'd216} : s = 344;
	{8'd128,8'd217} : s = 345;
	{8'd128,8'd218} : s = 346;
	{8'd128,8'd219} : s = 347;
	{8'd128,8'd220} : s = 348;
	{8'd128,8'd221} : s = 349;
	{8'd128,8'd222} : s = 350;
	{8'd128,8'd223} : s = 351;
	{8'd128,8'd224} : s = 352;
	{8'd128,8'd225} : s = 353;
	{8'd128,8'd226} : s = 354;
	{8'd128,8'd227} : s = 355;
	{8'd128,8'd228} : s = 356;
	{8'd128,8'd229} : s = 357;
	{8'd128,8'd230} : s = 358;
	{8'd128,8'd231} : s = 359;
	{8'd128,8'd232} : s = 360;
	{8'd128,8'd233} : s = 361;
	{8'd128,8'd234} : s = 362;
	{8'd128,8'd235} : s = 363;
	{8'd128,8'd236} : s = 364;
	{8'd128,8'd237} : s = 365;
	{8'd128,8'd238} : s = 366;
	{8'd128,8'd239} : s = 367;
	{8'd128,8'd240} : s = 368;
	{8'd128,8'd241} : s = 369;
	{8'd128,8'd242} : s = 370;
	{8'd128,8'd243} : s = 371;
	{8'd128,8'd244} : s = 372;
	{8'd128,8'd245} : s = 373;
	{8'd128,8'd246} : s = 374;
	{8'd128,8'd247} : s = 375;
	{8'd128,8'd248} : s = 376;
	{8'd128,8'd249} : s = 377;
	{8'd128,8'd250} : s = 378;
	{8'd128,8'd251} : s = 379;
	{8'd128,8'd252} : s = 380;
	{8'd128,8'd253} : s = 381;
	{8'd128,8'd254} : s = 382;
	{8'd128,8'd255} : s = 383;
	{8'd129,8'd0} : s = 129;
	{8'd129,8'd1} : s = 130;
	{8'd129,8'd2} : s = 131;
	{8'd129,8'd3} : s = 132;
	{8'd129,8'd4} : s = 133;
	{8'd129,8'd5} : s = 134;
	{8'd129,8'd6} : s = 135;
	{8'd129,8'd7} : s = 136;
	{8'd129,8'd8} : s = 137;
	{8'd129,8'd9} : s = 138;
	{8'd129,8'd10} : s = 139;
	{8'd129,8'd11} : s = 140;
	{8'd129,8'd12} : s = 141;
	{8'd129,8'd13} : s = 142;
	{8'd129,8'd14} : s = 143;
	{8'd129,8'd15} : s = 144;
	{8'd129,8'd16} : s = 145;
	{8'd129,8'd17} : s = 146;
	{8'd129,8'd18} : s = 147;
	{8'd129,8'd19} : s = 148;
	{8'd129,8'd20} : s = 149;
	{8'd129,8'd21} : s = 150;
	{8'd129,8'd22} : s = 151;
	{8'd129,8'd23} : s = 152;
	{8'd129,8'd24} : s = 153;
	{8'd129,8'd25} : s = 154;
	{8'd129,8'd26} : s = 155;
	{8'd129,8'd27} : s = 156;
	{8'd129,8'd28} : s = 157;
	{8'd129,8'd29} : s = 158;
	{8'd129,8'd30} : s = 159;
	{8'd129,8'd31} : s = 160;
	{8'd129,8'd32} : s = 161;
	{8'd129,8'd33} : s = 162;
	{8'd129,8'd34} : s = 163;
	{8'd129,8'd35} : s = 164;
	{8'd129,8'd36} : s = 165;
	{8'd129,8'd37} : s = 166;
	{8'd129,8'd38} : s = 167;
	{8'd129,8'd39} : s = 168;
	{8'd129,8'd40} : s = 169;
	{8'd129,8'd41} : s = 170;
	{8'd129,8'd42} : s = 171;
	{8'd129,8'd43} : s = 172;
	{8'd129,8'd44} : s = 173;
	{8'd129,8'd45} : s = 174;
	{8'd129,8'd46} : s = 175;
	{8'd129,8'd47} : s = 176;
	{8'd129,8'd48} : s = 177;
	{8'd129,8'd49} : s = 178;
	{8'd129,8'd50} : s = 179;
	{8'd129,8'd51} : s = 180;
	{8'd129,8'd52} : s = 181;
	{8'd129,8'd53} : s = 182;
	{8'd129,8'd54} : s = 183;
	{8'd129,8'd55} : s = 184;
	{8'd129,8'd56} : s = 185;
	{8'd129,8'd57} : s = 186;
	{8'd129,8'd58} : s = 187;
	{8'd129,8'd59} : s = 188;
	{8'd129,8'd60} : s = 189;
	{8'd129,8'd61} : s = 190;
	{8'd129,8'd62} : s = 191;
	{8'd129,8'd63} : s = 192;
	{8'd129,8'd64} : s = 193;
	{8'd129,8'd65} : s = 194;
	{8'd129,8'd66} : s = 195;
	{8'd129,8'd67} : s = 196;
	{8'd129,8'd68} : s = 197;
	{8'd129,8'd69} : s = 198;
	{8'd129,8'd70} : s = 199;
	{8'd129,8'd71} : s = 200;
	{8'd129,8'd72} : s = 201;
	{8'd129,8'd73} : s = 202;
	{8'd129,8'd74} : s = 203;
	{8'd129,8'd75} : s = 204;
	{8'd129,8'd76} : s = 205;
	{8'd129,8'd77} : s = 206;
	{8'd129,8'd78} : s = 207;
	{8'd129,8'd79} : s = 208;
	{8'd129,8'd80} : s = 209;
	{8'd129,8'd81} : s = 210;
	{8'd129,8'd82} : s = 211;
	{8'd129,8'd83} : s = 212;
	{8'd129,8'd84} : s = 213;
	{8'd129,8'd85} : s = 214;
	{8'd129,8'd86} : s = 215;
	{8'd129,8'd87} : s = 216;
	{8'd129,8'd88} : s = 217;
	{8'd129,8'd89} : s = 218;
	{8'd129,8'd90} : s = 219;
	{8'd129,8'd91} : s = 220;
	{8'd129,8'd92} : s = 221;
	{8'd129,8'd93} : s = 222;
	{8'd129,8'd94} : s = 223;
	{8'd129,8'd95} : s = 224;
	{8'd129,8'd96} : s = 225;
	{8'd129,8'd97} : s = 226;
	{8'd129,8'd98} : s = 227;
	{8'd129,8'd99} : s = 228;
	{8'd129,8'd100} : s = 229;
	{8'd129,8'd101} : s = 230;
	{8'd129,8'd102} : s = 231;
	{8'd129,8'd103} : s = 232;
	{8'd129,8'd104} : s = 233;
	{8'd129,8'd105} : s = 234;
	{8'd129,8'd106} : s = 235;
	{8'd129,8'd107} : s = 236;
	{8'd129,8'd108} : s = 237;
	{8'd129,8'd109} : s = 238;
	{8'd129,8'd110} : s = 239;
	{8'd129,8'd111} : s = 240;
	{8'd129,8'd112} : s = 241;
	{8'd129,8'd113} : s = 242;
	{8'd129,8'd114} : s = 243;
	{8'd129,8'd115} : s = 244;
	{8'd129,8'd116} : s = 245;
	{8'd129,8'd117} : s = 246;
	{8'd129,8'd118} : s = 247;
	{8'd129,8'd119} : s = 248;
	{8'd129,8'd120} : s = 249;
	{8'd129,8'd121} : s = 250;
	{8'd129,8'd122} : s = 251;
	{8'd129,8'd123} : s = 252;
	{8'd129,8'd124} : s = 253;
	{8'd129,8'd125} : s = 254;
	{8'd129,8'd126} : s = 255;
	{8'd129,8'd127} : s = 256;
	{8'd129,8'd128} : s = 257;
	{8'd129,8'd129} : s = 258;
	{8'd129,8'd130} : s = 259;
	{8'd129,8'd131} : s = 260;
	{8'd129,8'd132} : s = 261;
	{8'd129,8'd133} : s = 262;
	{8'd129,8'd134} : s = 263;
	{8'd129,8'd135} : s = 264;
	{8'd129,8'd136} : s = 265;
	{8'd129,8'd137} : s = 266;
	{8'd129,8'd138} : s = 267;
	{8'd129,8'd139} : s = 268;
	{8'd129,8'd140} : s = 269;
	{8'd129,8'd141} : s = 270;
	{8'd129,8'd142} : s = 271;
	{8'd129,8'd143} : s = 272;
	{8'd129,8'd144} : s = 273;
	{8'd129,8'd145} : s = 274;
	{8'd129,8'd146} : s = 275;
	{8'd129,8'd147} : s = 276;
	{8'd129,8'd148} : s = 277;
	{8'd129,8'd149} : s = 278;
	{8'd129,8'd150} : s = 279;
	{8'd129,8'd151} : s = 280;
	{8'd129,8'd152} : s = 281;
	{8'd129,8'd153} : s = 282;
	{8'd129,8'd154} : s = 283;
	{8'd129,8'd155} : s = 284;
	{8'd129,8'd156} : s = 285;
	{8'd129,8'd157} : s = 286;
	{8'd129,8'd158} : s = 287;
	{8'd129,8'd159} : s = 288;
	{8'd129,8'd160} : s = 289;
	{8'd129,8'd161} : s = 290;
	{8'd129,8'd162} : s = 291;
	{8'd129,8'd163} : s = 292;
	{8'd129,8'd164} : s = 293;
	{8'd129,8'd165} : s = 294;
	{8'd129,8'd166} : s = 295;
	{8'd129,8'd167} : s = 296;
	{8'd129,8'd168} : s = 297;
	{8'd129,8'd169} : s = 298;
	{8'd129,8'd170} : s = 299;
	{8'd129,8'd171} : s = 300;
	{8'd129,8'd172} : s = 301;
	{8'd129,8'd173} : s = 302;
	{8'd129,8'd174} : s = 303;
	{8'd129,8'd175} : s = 304;
	{8'd129,8'd176} : s = 305;
	{8'd129,8'd177} : s = 306;
	{8'd129,8'd178} : s = 307;
	{8'd129,8'd179} : s = 308;
	{8'd129,8'd180} : s = 309;
	{8'd129,8'd181} : s = 310;
	{8'd129,8'd182} : s = 311;
	{8'd129,8'd183} : s = 312;
	{8'd129,8'd184} : s = 313;
	{8'd129,8'd185} : s = 314;
	{8'd129,8'd186} : s = 315;
	{8'd129,8'd187} : s = 316;
	{8'd129,8'd188} : s = 317;
	{8'd129,8'd189} : s = 318;
	{8'd129,8'd190} : s = 319;
	{8'd129,8'd191} : s = 320;
	{8'd129,8'd192} : s = 321;
	{8'd129,8'd193} : s = 322;
	{8'd129,8'd194} : s = 323;
	{8'd129,8'd195} : s = 324;
	{8'd129,8'd196} : s = 325;
	{8'd129,8'd197} : s = 326;
	{8'd129,8'd198} : s = 327;
	{8'd129,8'd199} : s = 328;
	{8'd129,8'd200} : s = 329;
	{8'd129,8'd201} : s = 330;
	{8'd129,8'd202} : s = 331;
	{8'd129,8'd203} : s = 332;
	{8'd129,8'd204} : s = 333;
	{8'd129,8'd205} : s = 334;
	{8'd129,8'd206} : s = 335;
	{8'd129,8'd207} : s = 336;
	{8'd129,8'd208} : s = 337;
	{8'd129,8'd209} : s = 338;
	{8'd129,8'd210} : s = 339;
	{8'd129,8'd211} : s = 340;
	{8'd129,8'd212} : s = 341;
	{8'd129,8'd213} : s = 342;
	{8'd129,8'd214} : s = 343;
	{8'd129,8'd215} : s = 344;
	{8'd129,8'd216} : s = 345;
	{8'd129,8'd217} : s = 346;
	{8'd129,8'd218} : s = 347;
	{8'd129,8'd219} : s = 348;
	{8'd129,8'd220} : s = 349;
	{8'd129,8'd221} : s = 350;
	{8'd129,8'd222} : s = 351;
	{8'd129,8'd223} : s = 352;
	{8'd129,8'd224} : s = 353;
	{8'd129,8'd225} : s = 354;
	{8'd129,8'd226} : s = 355;
	{8'd129,8'd227} : s = 356;
	{8'd129,8'd228} : s = 357;
	{8'd129,8'd229} : s = 358;
	{8'd129,8'd230} : s = 359;
	{8'd129,8'd231} : s = 360;
	{8'd129,8'd232} : s = 361;
	{8'd129,8'd233} : s = 362;
	{8'd129,8'd234} : s = 363;
	{8'd129,8'd235} : s = 364;
	{8'd129,8'd236} : s = 365;
	{8'd129,8'd237} : s = 366;
	{8'd129,8'd238} : s = 367;
	{8'd129,8'd239} : s = 368;
	{8'd129,8'd240} : s = 369;
	{8'd129,8'd241} : s = 370;
	{8'd129,8'd242} : s = 371;
	{8'd129,8'd243} : s = 372;
	{8'd129,8'd244} : s = 373;
	{8'd129,8'd245} : s = 374;
	{8'd129,8'd246} : s = 375;
	{8'd129,8'd247} : s = 376;
	{8'd129,8'd248} : s = 377;
	{8'd129,8'd249} : s = 378;
	{8'd129,8'd250} : s = 379;
	{8'd129,8'd251} : s = 380;
	{8'd129,8'd252} : s = 381;
	{8'd129,8'd253} : s = 382;
	{8'd129,8'd254} : s = 383;
	{8'd129,8'd255} : s = 384;
	{8'd130,8'd0} : s = 130;
	{8'd130,8'd1} : s = 131;
	{8'd130,8'd2} : s = 132;
	{8'd130,8'd3} : s = 133;
	{8'd130,8'd4} : s = 134;
	{8'd130,8'd5} : s = 135;
	{8'd130,8'd6} : s = 136;
	{8'd130,8'd7} : s = 137;
	{8'd130,8'd8} : s = 138;
	{8'd130,8'd9} : s = 139;
	{8'd130,8'd10} : s = 140;
	{8'd130,8'd11} : s = 141;
	{8'd130,8'd12} : s = 142;
	{8'd130,8'd13} : s = 143;
	{8'd130,8'd14} : s = 144;
	{8'd130,8'd15} : s = 145;
	{8'd130,8'd16} : s = 146;
	{8'd130,8'd17} : s = 147;
	{8'd130,8'd18} : s = 148;
	{8'd130,8'd19} : s = 149;
	{8'd130,8'd20} : s = 150;
	{8'd130,8'd21} : s = 151;
	{8'd130,8'd22} : s = 152;
	{8'd130,8'd23} : s = 153;
	{8'd130,8'd24} : s = 154;
	{8'd130,8'd25} : s = 155;
	{8'd130,8'd26} : s = 156;
	{8'd130,8'd27} : s = 157;
	{8'd130,8'd28} : s = 158;
	{8'd130,8'd29} : s = 159;
	{8'd130,8'd30} : s = 160;
	{8'd130,8'd31} : s = 161;
	{8'd130,8'd32} : s = 162;
	{8'd130,8'd33} : s = 163;
	{8'd130,8'd34} : s = 164;
	{8'd130,8'd35} : s = 165;
	{8'd130,8'd36} : s = 166;
	{8'd130,8'd37} : s = 167;
	{8'd130,8'd38} : s = 168;
	{8'd130,8'd39} : s = 169;
	{8'd130,8'd40} : s = 170;
	{8'd130,8'd41} : s = 171;
	{8'd130,8'd42} : s = 172;
	{8'd130,8'd43} : s = 173;
	{8'd130,8'd44} : s = 174;
	{8'd130,8'd45} : s = 175;
	{8'd130,8'd46} : s = 176;
	{8'd130,8'd47} : s = 177;
	{8'd130,8'd48} : s = 178;
	{8'd130,8'd49} : s = 179;
	{8'd130,8'd50} : s = 180;
	{8'd130,8'd51} : s = 181;
	{8'd130,8'd52} : s = 182;
	{8'd130,8'd53} : s = 183;
	{8'd130,8'd54} : s = 184;
	{8'd130,8'd55} : s = 185;
	{8'd130,8'd56} : s = 186;
	{8'd130,8'd57} : s = 187;
	{8'd130,8'd58} : s = 188;
	{8'd130,8'd59} : s = 189;
	{8'd130,8'd60} : s = 190;
	{8'd130,8'd61} : s = 191;
	{8'd130,8'd62} : s = 192;
	{8'd130,8'd63} : s = 193;
	{8'd130,8'd64} : s = 194;
	{8'd130,8'd65} : s = 195;
	{8'd130,8'd66} : s = 196;
	{8'd130,8'd67} : s = 197;
	{8'd130,8'd68} : s = 198;
	{8'd130,8'd69} : s = 199;
	{8'd130,8'd70} : s = 200;
	{8'd130,8'd71} : s = 201;
	{8'd130,8'd72} : s = 202;
	{8'd130,8'd73} : s = 203;
	{8'd130,8'd74} : s = 204;
	{8'd130,8'd75} : s = 205;
	{8'd130,8'd76} : s = 206;
	{8'd130,8'd77} : s = 207;
	{8'd130,8'd78} : s = 208;
	{8'd130,8'd79} : s = 209;
	{8'd130,8'd80} : s = 210;
	{8'd130,8'd81} : s = 211;
	{8'd130,8'd82} : s = 212;
	{8'd130,8'd83} : s = 213;
	{8'd130,8'd84} : s = 214;
	{8'd130,8'd85} : s = 215;
	{8'd130,8'd86} : s = 216;
	{8'd130,8'd87} : s = 217;
	{8'd130,8'd88} : s = 218;
	{8'd130,8'd89} : s = 219;
	{8'd130,8'd90} : s = 220;
	{8'd130,8'd91} : s = 221;
	{8'd130,8'd92} : s = 222;
	{8'd130,8'd93} : s = 223;
	{8'd130,8'd94} : s = 224;
	{8'd130,8'd95} : s = 225;
	{8'd130,8'd96} : s = 226;
	{8'd130,8'd97} : s = 227;
	{8'd130,8'd98} : s = 228;
	{8'd130,8'd99} : s = 229;
	{8'd130,8'd100} : s = 230;
	{8'd130,8'd101} : s = 231;
	{8'd130,8'd102} : s = 232;
	{8'd130,8'd103} : s = 233;
	{8'd130,8'd104} : s = 234;
	{8'd130,8'd105} : s = 235;
	{8'd130,8'd106} : s = 236;
	{8'd130,8'd107} : s = 237;
	{8'd130,8'd108} : s = 238;
	{8'd130,8'd109} : s = 239;
	{8'd130,8'd110} : s = 240;
	{8'd130,8'd111} : s = 241;
	{8'd130,8'd112} : s = 242;
	{8'd130,8'd113} : s = 243;
	{8'd130,8'd114} : s = 244;
	{8'd130,8'd115} : s = 245;
	{8'd130,8'd116} : s = 246;
	{8'd130,8'd117} : s = 247;
	{8'd130,8'd118} : s = 248;
	{8'd130,8'd119} : s = 249;
	{8'd130,8'd120} : s = 250;
	{8'd130,8'd121} : s = 251;
	{8'd130,8'd122} : s = 252;
	{8'd130,8'd123} : s = 253;
	{8'd130,8'd124} : s = 254;
	{8'd130,8'd125} : s = 255;
	{8'd130,8'd126} : s = 256;
	{8'd130,8'd127} : s = 257;
	{8'd130,8'd128} : s = 258;
	{8'd130,8'd129} : s = 259;
	{8'd130,8'd130} : s = 260;
	{8'd130,8'd131} : s = 261;
	{8'd130,8'd132} : s = 262;
	{8'd130,8'd133} : s = 263;
	{8'd130,8'd134} : s = 264;
	{8'd130,8'd135} : s = 265;
	{8'd130,8'd136} : s = 266;
	{8'd130,8'd137} : s = 267;
	{8'd130,8'd138} : s = 268;
	{8'd130,8'd139} : s = 269;
	{8'd130,8'd140} : s = 270;
	{8'd130,8'd141} : s = 271;
	{8'd130,8'd142} : s = 272;
	{8'd130,8'd143} : s = 273;
	{8'd130,8'd144} : s = 274;
	{8'd130,8'd145} : s = 275;
	{8'd130,8'd146} : s = 276;
	{8'd130,8'd147} : s = 277;
	{8'd130,8'd148} : s = 278;
	{8'd130,8'd149} : s = 279;
	{8'd130,8'd150} : s = 280;
	{8'd130,8'd151} : s = 281;
	{8'd130,8'd152} : s = 282;
	{8'd130,8'd153} : s = 283;
	{8'd130,8'd154} : s = 284;
	{8'd130,8'd155} : s = 285;
	{8'd130,8'd156} : s = 286;
	{8'd130,8'd157} : s = 287;
	{8'd130,8'd158} : s = 288;
	{8'd130,8'd159} : s = 289;
	{8'd130,8'd160} : s = 290;
	{8'd130,8'd161} : s = 291;
	{8'd130,8'd162} : s = 292;
	{8'd130,8'd163} : s = 293;
	{8'd130,8'd164} : s = 294;
	{8'd130,8'd165} : s = 295;
	{8'd130,8'd166} : s = 296;
	{8'd130,8'd167} : s = 297;
	{8'd130,8'd168} : s = 298;
	{8'd130,8'd169} : s = 299;
	{8'd130,8'd170} : s = 300;
	{8'd130,8'd171} : s = 301;
	{8'd130,8'd172} : s = 302;
	{8'd130,8'd173} : s = 303;
	{8'd130,8'd174} : s = 304;
	{8'd130,8'd175} : s = 305;
	{8'd130,8'd176} : s = 306;
	{8'd130,8'd177} : s = 307;
	{8'd130,8'd178} : s = 308;
	{8'd130,8'd179} : s = 309;
	{8'd130,8'd180} : s = 310;
	{8'd130,8'd181} : s = 311;
	{8'd130,8'd182} : s = 312;
	{8'd130,8'd183} : s = 313;
	{8'd130,8'd184} : s = 314;
	{8'd130,8'd185} : s = 315;
	{8'd130,8'd186} : s = 316;
	{8'd130,8'd187} : s = 317;
	{8'd130,8'd188} : s = 318;
	{8'd130,8'd189} : s = 319;
	{8'd130,8'd190} : s = 320;
	{8'd130,8'd191} : s = 321;
	{8'd130,8'd192} : s = 322;
	{8'd130,8'd193} : s = 323;
	{8'd130,8'd194} : s = 324;
	{8'd130,8'd195} : s = 325;
	{8'd130,8'd196} : s = 326;
	{8'd130,8'd197} : s = 327;
	{8'd130,8'd198} : s = 328;
	{8'd130,8'd199} : s = 329;
	{8'd130,8'd200} : s = 330;
	{8'd130,8'd201} : s = 331;
	{8'd130,8'd202} : s = 332;
	{8'd130,8'd203} : s = 333;
	{8'd130,8'd204} : s = 334;
	{8'd130,8'd205} : s = 335;
	{8'd130,8'd206} : s = 336;
	{8'd130,8'd207} : s = 337;
	{8'd130,8'd208} : s = 338;
	{8'd130,8'd209} : s = 339;
	{8'd130,8'd210} : s = 340;
	{8'd130,8'd211} : s = 341;
	{8'd130,8'd212} : s = 342;
	{8'd130,8'd213} : s = 343;
	{8'd130,8'd214} : s = 344;
	{8'd130,8'd215} : s = 345;
	{8'd130,8'd216} : s = 346;
	{8'd130,8'd217} : s = 347;
	{8'd130,8'd218} : s = 348;
	{8'd130,8'd219} : s = 349;
	{8'd130,8'd220} : s = 350;
	{8'd130,8'd221} : s = 351;
	{8'd130,8'd222} : s = 352;
	{8'd130,8'd223} : s = 353;
	{8'd130,8'd224} : s = 354;
	{8'd130,8'd225} : s = 355;
	{8'd130,8'd226} : s = 356;
	{8'd130,8'd227} : s = 357;
	{8'd130,8'd228} : s = 358;
	{8'd130,8'd229} : s = 359;
	{8'd130,8'd230} : s = 360;
	{8'd130,8'd231} : s = 361;
	{8'd130,8'd232} : s = 362;
	{8'd130,8'd233} : s = 363;
	{8'd130,8'd234} : s = 364;
	{8'd130,8'd235} : s = 365;
	{8'd130,8'd236} : s = 366;
	{8'd130,8'd237} : s = 367;
	{8'd130,8'd238} : s = 368;
	{8'd130,8'd239} : s = 369;
	{8'd130,8'd240} : s = 370;
	{8'd130,8'd241} : s = 371;
	{8'd130,8'd242} : s = 372;
	{8'd130,8'd243} : s = 373;
	{8'd130,8'd244} : s = 374;
	{8'd130,8'd245} : s = 375;
	{8'd130,8'd246} : s = 376;
	{8'd130,8'd247} : s = 377;
	{8'd130,8'd248} : s = 378;
	{8'd130,8'd249} : s = 379;
	{8'd130,8'd250} : s = 380;
	{8'd130,8'd251} : s = 381;
	{8'd130,8'd252} : s = 382;
	{8'd130,8'd253} : s = 383;
	{8'd130,8'd254} : s = 384;
	{8'd130,8'd255} : s = 385;
	{8'd131,8'd0} : s = 131;
	{8'd131,8'd1} : s = 132;
	{8'd131,8'd2} : s = 133;
	{8'd131,8'd3} : s = 134;
	{8'd131,8'd4} : s = 135;
	{8'd131,8'd5} : s = 136;
	{8'd131,8'd6} : s = 137;
	{8'd131,8'd7} : s = 138;
	{8'd131,8'd8} : s = 139;
	{8'd131,8'd9} : s = 140;
	{8'd131,8'd10} : s = 141;
	{8'd131,8'd11} : s = 142;
	{8'd131,8'd12} : s = 143;
	{8'd131,8'd13} : s = 144;
	{8'd131,8'd14} : s = 145;
	{8'd131,8'd15} : s = 146;
	{8'd131,8'd16} : s = 147;
	{8'd131,8'd17} : s = 148;
	{8'd131,8'd18} : s = 149;
	{8'd131,8'd19} : s = 150;
	{8'd131,8'd20} : s = 151;
	{8'd131,8'd21} : s = 152;
	{8'd131,8'd22} : s = 153;
	{8'd131,8'd23} : s = 154;
	{8'd131,8'd24} : s = 155;
	{8'd131,8'd25} : s = 156;
	{8'd131,8'd26} : s = 157;
	{8'd131,8'd27} : s = 158;
	{8'd131,8'd28} : s = 159;
	{8'd131,8'd29} : s = 160;
	{8'd131,8'd30} : s = 161;
	{8'd131,8'd31} : s = 162;
	{8'd131,8'd32} : s = 163;
	{8'd131,8'd33} : s = 164;
	{8'd131,8'd34} : s = 165;
	{8'd131,8'd35} : s = 166;
	{8'd131,8'd36} : s = 167;
	{8'd131,8'd37} : s = 168;
	{8'd131,8'd38} : s = 169;
	{8'd131,8'd39} : s = 170;
	{8'd131,8'd40} : s = 171;
	{8'd131,8'd41} : s = 172;
	{8'd131,8'd42} : s = 173;
	{8'd131,8'd43} : s = 174;
	{8'd131,8'd44} : s = 175;
	{8'd131,8'd45} : s = 176;
	{8'd131,8'd46} : s = 177;
	{8'd131,8'd47} : s = 178;
	{8'd131,8'd48} : s = 179;
	{8'd131,8'd49} : s = 180;
	{8'd131,8'd50} : s = 181;
	{8'd131,8'd51} : s = 182;
	{8'd131,8'd52} : s = 183;
	{8'd131,8'd53} : s = 184;
	{8'd131,8'd54} : s = 185;
	{8'd131,8'd55} : s = 186;
	{8'd131,8'd56} : s = 187;
	{8'd131,8'd57} : s = 188;
	{8'd131,8'd58} : s = 189;
	{8'd131,8'd59} : s = 190;
	{8'd131,8'd60} : s = 191;
	{8'd131,8'd61} : s = 192;
	{8'd131,8'd62} : s = 193;
	{8'd131,8'd63} : s = 194;
	{8'd131,8'd64} : s = 195;
	{8'd131,8'd65} : s = 196;
	{8'd131,8'd66} : s = 197;
	{8'd131,8'd67} : s = 198;
	{8'd131,8'd68} : s = 199;
	{8'd131,8'd69} : s = 200;
	{8'd131,8'd70} : s = 201;
	{8'd131,8'd71} : s = 202;
	{8'd131,8'd72} : s = 203;
	{8'd131,8'd73} : s = 204;
	{8'd131,8'd74} : s = 205;
	{8'd131,8'd75} : s = 206;
	{8'd131,8'd76} : s = 207;
	{8'd131,8'd77} : s = 208;
	{8'd131,8'd78} : s = 209;
	{8'd131,8'd79} : s = 210;
	{8'd131,8'd80} : s = 211;
	{8'd131,8'd81} : s = 212;
	{8'd131,8'd82} : s = 213;
	{8'd131,8'd83} : s = 214;
	{8'd131,8'd84} : s = 215;
	{8'd131,8'd85} : s = 216;
	{8'd131,8'd86} : s = 217;
	{8'd131,8'd87} : s = 218;
	{8'd131,8'd88} : s = 219;
	{8'd131,8'd89} : s = 220;
	{8'd131,8'd90} : s = 221;
	{8'd131,8'd91} : s = 222;
	{8'd131,8'd92} : s = 223;
	{8'd131,8'd93} : s = 224;
	{8'd131,8'd94} : s = 225;
	{8'd131,8'd95} : s = 226;
	{8'd131,8'd96} : s = 227;
	{8'd131,8'd97} : s = 228;
	{8'd131,8'd98} : s = 229;
	{8'd131,8'd99} : s = 230;
	{8'd131,8'd100} : s = 231;
	{8'd131,8'd101} : s = 232;
	{8'd131,8'd102} : s = 233;
	{8'd131,8'd103} : s = 234;
	{8'd131,8'd104} : s = 235;
	{8'd131,8'd105} : s = 236;
	{8'd131,8'd106} : s = 237;
	{8'd131,8'd107} : s = 238;
	{8'd131,8'd108} : s = 239;
	{8'd131,8'd109} : s = 240;
	{8'd131,8'd110} : s = 241;
	{8'd131,8'd111} : s = 242;
	{8'd131,8'd112} : s = 243;
	{8'd131,8'd113} : s = 244;
	{8'd131,8'd114} : s = 245;
	{8'd131,8'd115} : s = 246;
	{8'd131,8'd116} : s = 247;
	{8'd131,8'd117} : s = 248;
	{8'd131,8'd118} : s = 249;
	{8'd131,8'd119} : s = 250;
	{8'd131,8'd120} : s = 251;
	{8'd131,8'd121} : s = 252;
	{8'd131,8'd122} : s = 253;
	{8'd131,8'd123} : s = 254;
	{8'd131,8'd124} : s = 255;
	{8'd131,8'd125} : s = 256;
	{8'd131,8'd126} : s = 257;
	{8'd131,8'd127} : s = 258;
	{8'd131,8'd128} : s = 259;
	{8'd131,8'd129} : s = 260;
	{8'd131,8'd130} : s = 261;
	{8'd131,8'd131} : s = 262;
	{8'd131,8'd132} : s = 263;
	{8'd131,8'd133} : s = 264;
	{8'd131,8'd134} : s = 265;
	{8'd131,8'd135} : s = 266;
	{8'd131,8'd136} : s = 267;
	{8'd131,8'd137} : s = 268;
	{8'd131,8'd138} : s = 269;
	{8'd131,8'd139} : s = 270;
	{8'd131,8'd140} : s = 271;
	{8'd131,8'd141} : s = 272;
	{8'd131,8'd142} : s = 273;
	{8'd131,8'd143} : s = 274;
	{8'd131,8'd144} : s = 275;
	{8'd131,8'd145} : s = 276;
	{8'd131,8'd146} : s = 277;
	{8'd131,8'd147} : s = 278;
	{8'd131,8'd148} : s = 279;
	{8'd131,8'd149} : s = 280;
	{8'd131,8'd150} : s = 281;
	{8'd131,8'd151} : s = 282;
	{8'd131,8'd152} : s = 283;
	{8'd131,8'd153} : s = 284;
	{8'd131,8'd154} : s = 285;
	{8'd131,8'd155} : s = 286;
	{8'd131,8'd156} : s = 287;
	{8'd131,8'd157} : s = 288;
	{8'd131,8'd158} : s = 289;
	{8'd131,8'd159} : s = 290;
	{8'd131,8'd160} : s = 291;
	{8'd131,8'd161} : s = 292;
	{8'd131,8'd162} : s = 293;
	{8'd131,8'd163} : s = 294;
	{8'd131,8'd164} : s = 295;
	{8'd131,8'd165} : s = 296;
	{8'd131,8'd166} : s = 297;
	{8'd131,8'd167} : s = 298;
	{8'd131,8'd168} : s = 299;
	{8'd131,8'd169} : s = 300;
	{8'd131,8'd170} : s = 301;
	{8'd131,8'd171} : s = 302;
	{8'd131,8'd172} : s = 303;
	{8'd131,8'd173} : s = 304;
	{8'd131,8'd174} : s = 305;
	{8'd131,8'd175} : s = 306;
	{8'd131,8'd176} : s = 307;
	{8'd131,8'd177} : s = 308;
	{8'd131,8'd178} : s = 309;
	{8'd131,8'd179} : s = 310;
	{8'd131,8'd180} : s = 311;
	{8'd131,8'd181} : s = 312;
	{8'd131,8'd182} : s = 313;
	{8'd131,8'd183} : s = 314;
	{8'd131,8'd184} : s = 315;
	{8'd131,8'd185} : s = 316;
	{8'd131,8'd186} : s = 317;
	{8'd131,8'd187} : s = 318;
	{8'd131,8'd188} : s = 319;
	{8'd131,8'd189} : s = 320;
	{8'd131,8'd190} : s = 321;
	{8'd131,8'd191} : s = 322;
	{8'd131,8'd192} : s = 323;
	{8'd131,8'd193} : s = 324;
	{8'd131,8'd194} : s = 325;
	{8'd131,8'd195} : s = 326;
	{8'd131,8'd196} : s = 327;
	{8'd131,8'd197} : s = 328;
	{8'd131,8'd198} : s = 329;
	{8'd131,8'd199} : s = 330;
	{8'd131,8'd200} : s = 331;
	{8'd131,8'd201} : s = 332;
	{8'd131,8'd202} : s = 333;
	{8'd131,8'd203} : s = 334;
	{8'd131,8'd204} : s = 335;
	{8'd131,8'd205} : s = 336;
	{8'd131,8'd206} : s = 337;
	{8'd131,8'd207} : s = 338;
	{8'd131,8'd208} : s = 339;
	{8'd131,8'd209} : s = 340;
	{8'd131,8'd210} : s = 341;
	{8'd131,8'd211} : s = 342;
	{8'd131,8'd212} : s = 343;
	{8'd131,8'd213} : s = 344;
	{8'd131,8'd214} : s = 345;
	{8'd131,8'd215} : s = 346;
	{8'd131,8'd216} : s = 347;
	{8'd131,8'd217} : s = 348;
	{8'd131,8'd218} : s = 349;
	{8'd131,8'd219} : s = 350;
	{8'd131,8'd220} : s = 351;
	{8'd131,8'd221} : s = 352;
	{8'd131,8'd222} : s = 353;
	{8'd131,8'd223} : s = 354;
	{8'd131,8'd224} : s = 355;
	{8'd131,8'd225} : s = 356;
	{8'd131,8'd226} : s = 357;
	{8'd131,8'd227} : s = 358;
	{8'd131,8'd228} : s = 359;
	{8'd131,8'd229} : s = 360;
	{8'd131,8'd230} : s = 361;
	{8'd131,8'd231} : s = 362;
	{8'd131,8'd232} : s = 363;
	{8'd131,8'd233} : s = 364;
	{8'd131,8'd234} : s = 365;
	{8'd131,8'd235} : s = 366;
	{8'd131,8'd236} : s = 367;
	{8'd131,8'd237} : s = 368;
	{8'd131,8'd238} : s = 369;
	{8'd131,8'd239} : s = 370;
	{8'd131,8'd240} : s = 371;
	{8'd131,8'd241} : s = 372;
	{8'd131,8'd242} : s = 373;
	{8'd131,8'd243} : s = 374;
	{8'd131,8'd244} : s = 375;
	{8'd131,8'd245} : s = 376;
	{8'd131,8'd246} : s = 377;
	{8'd131,8'd247} : s = 378;
	{8'd131,8'd248} : s = 379;
	{8'd131,8'd249} : s = 380;
	{8'd131,8'd250} : s = 381;
	{8'd131,8'd251} : s = 382;
	{8'd131,8'd252} : s = 383;
	{8'd131,8'd253} : s = 384;
	{8'd131,8'd254} : s = 385;
	{8'd131,8'd255} : s = 386;
	{8'd132,8'd0} : s = 132;
	{8'd132,8'd1} : s = 133;
	{8'd132,8'd2} : s = 134;
	{8'd132,8'd3} : s = 135;
	{8'd132,8'd4} : s = 136;
	{8'd132,8'd5} : s = 137;
	{8'd132,8'd6} : s = 138;
	{8'd132,8'd7} : s = 139;
	{8'd132,8'd8} : s = 140;
	{8'd132,8'd9} : s = 141;
	{8'd132,8'd10} : s = 142;
	{8'd132,8'd11} : s = 143;
	{8'd132,8'd12} : s = 144;
	{8'd132,8'd13} : s = 145;
	{8'd132,8'd14} : s = 146;
	{8'd132,8'd15} : s = 147;
	{8'd132,8'd16} : s = 148;
	{8'd132,8'd17} : s = 149;
	{8'd132,8'd18} : s = 150;
	{8'd132,8'd19} : s = 151;
	{8'd132,8'd20} : s = 152;
	{8'd132,8'd21} : s = 153;
	{8'd132,8'd22} : s = 154;
	{8'd132,8'd23} : s = 155;
	{8'd132,8'd24} : s = 156;
	{8'd132,8'd25} : s = 157;
	{8'd132,8'd26} : s = 158;
	{8'd132,8'd27} : s = 159;
	{8'd132,8'd28} : s = 160;
	{8'd132,8'd29} : s = 161;
	{8'd132,8'd30} : s = 162;
	{8'd132,8'd31} : s = 163;
	{8'd132,8'd32} : s = 164;
	{8'd132,8'd33} : s = 165;
	{8'd132,8'd34} : s = 166;
	{8'd132,8'd35} : s = 167;
	{8'd132,8'd36} : s = 168;
	{8'd132,8'd37} : s = 169;
	{8'd132,8'd38} : s = 170;
	{8'd132,8'd39} : s = 171;
	{8'd132,8'd40} : s = 172;
	{8'd132,8'd41} : s = 173;
	{8'd132,8'd42} : s = 174;
	{8'd132,8'd43} : s = 175;
	{8'd132,8'd44} : s = 176;
	{8'd132,8'd45} : s = 177;
	{8'd132,8'd46} : s = 178;
	{8'd132,8'd47} : s = 179;
	{8'd132,8'd48} : s = 180;
	{8'd132,8'd49} : s = 181;
	{8'd132,8'd50} : s = 182;
	{8'd132,8'd51} : s = 183;
	{8'd132,8'd52} : s = 184;
	{8'd132,8'd53} : s = 185;
	{8'd132,8'd54} : s = 186;
	{8'd132,8'd55} : s = 187;
	{8'd132,8'd56} : s = 188;
	{8'd132,8'd57} : s = 189;
	{8'd132,8'd58} : s = 190;
	{8'd132,8'd59} : s = 191;
	{8'd132,8'd60} : s = 192;
	{8'd132,8'd61} : s = 193;
	{8'd132,8'd62} : s = 194;
	{8'd132,8'd63} : s = 195;
	{8'd132,8'd64} : s = 196;
	{8'd132,8'd65} : s = 197;
	{8'd132,8'd66} : s = 198;
	{8'd132,8'd67} : s = 199;
	{8'd132,8'd68} : s = 200;
	{8'd132,8'd69} : s = 201;
	{8'd132,8'd70} : s = 202;
	{8'd132,8'd71} : s = 203;
	{8'd132,8'd72} : s = 204;
	{8'd132,8'd73} : s = 205;
	{8'd132,8'd74} : s = 206;
	{8'd132,8'd75} : s = 207;
	{8'd132,8'd76} : s = 208;
	{8'd132,8'd77} : s = 209;
	{8'd132,8'd78} : s = 210;
	{8'd132,8'd79} : s = 211;
	{8'd132,8'd80} : s = 212;
	{8'd132,8'd81} : s = 213;
	{8'd132,8'd82} : s = 214;
	{8'd132,8'd83} : s = 215;
	{8'd132,8'd84} : s = 216;
	{8'd132,8'd85} : s = 217;
	{8'd132,8'd86} : s = 218;
	{8'd132,8'd87} : s = 219;
	{8'd132,8'd88} : s = 220;
	{8'd132,8'd89} : s = 221;
	{8'd132,8'd90} : s = 222;
	{8'd132,8'd91} : s = 223;
	{8'd132,8'd92} : s = 224;
	{8'd132,8'd93} : s = 225;
	{8'd132,8'd94} : s = 226;
	{8'd132,8'd95} : s = 227;
	{8'd132,8'd96} : s = 228;
	{8'd132,8'd97} : s = 229;
	{8'd132,8'd98} : s = 230;
	{8'd132,8'd99} : s = 231;
	{8'd132,8'd100} : s = 232;
	{8'd132,8'd101} : s = 233;
	{8'd132,8'd102} : s = 234;
	{8'd132,8'd103} : s = 235;
	{8'd132,8'd104} : s = 236;
	{8'd132,8'd105} : s = 237;
	{8'd132,8'd106} : s = 238;
	{8'd132,8'd107} : s = 239;
	{8'd132,8'd108} : s = 240;
	{8'd132,8'd109} : s = 241;
	{8'd132,8'd110} : s = 242;
	{8'd132,8'd111} : s = 243;
	{8'd132,8'd112} : s = 244;
	{8'd132,8'd113} : s = 245;
	{8'd132,8'd114} : s = 246;
	{8'd132,8'd115} : s = 247;
	{8'd132,8'd116} : s = 248;
	{8'd132,8'd117} : s = 249;
	{8'd132,8'd118} : s = 250;
	{8'd132,8'd119} : s = 251;
	{8'd132,8'd120} : s = 252;
	{8'd132,8'd121} : s = 253;
	{8'd132,8'd122} : s = 254;
	{8'd132,8'd123} : s = 255;
	{8'd132,8'd124} : s = 256;
	{8'd132,8'd125} : s = 257;
	{8'd132,8'd126} : s = 258;
	{8'd132,8'd127} : s = 259;
	{8'd132,8'd128} : s = 260;
	{8'd132,8'd129} : s = 261;
	{8'd132,8'd130} : s = 262;
	{8'd132,8'd131} : s = 263;
	{8'd132,8'd132} : s = 264;
	{8'd132,8'd133} : s = 265;
	{8'd132,8'd134} : s = 266;
	{8'd132,8'd135} : s = 267;
	{8'd132,8'd136} : s = 268;
	{8'd132,8'd137} : s = 269;
	{8'd132,8'd138} : s = 270;
	{8'd132,8'd139} : s = 271;
	{8'd132,8'd140} : s = 272;
	{8'd132,8'd141} : s = 273;
	{8'd132,8'd142} : s = 274;
	{8'd132,8'd143} : s = 275;
	{8'd132,8'd144} : s = 276;
	{8'd132,8'd145} : s = 277;
	{8'd132,8'd146} : s = 278;
	{8'd132,8'd147} : s = 279;
	{8'd132,8'd148} : s = 280;
	{8'd132,8'd149} : s = 281;
	{8'd132,8'd150} : s = 282;
	{8'd132,8'd151} : s = 283;
	{8'd132,8'd152} : s = 284;
	{8'd132,8'd153} : s = 285;
	{8'd132,8'd154} : s = 286;
	{8'd132,8'd155} : s = 287;
	{8'd132,8'd156} : s = 288;
	{8'd132,8'd157} : s = 289;
	{8'd132,8'd158} : s = 290;
	{8'd132,8'd159} : s = 291;
	{8'd132,8'd160} : s = 292;
	{8'd132,8'd161} : s = 293;
	{8'd132,8'd162} : s = 294;
	{8'd132,8'd163} : s = 295;
	{8'd132,8'd164} : s = 296;
	{8'd132,8'd165} : s = 297;
	{8'd132,8'd166} : s = 298;
	{8'd132,8'd167} : s = 299;
	{8'd132,8'd168} : s = 300;
	{8'd132,8'd169} : s = 301;
	{8'd132,8'd170} : s = 302;
	{8'd132,8'd171} : s = 303;
	{8'd132,8'd172} : s = 304;
	{8'd132,8'd173} : s = 305;
	{8'd132,8'd174} : s = 306;
	{8'd132,8'd175} : s = 307;
	{8'd132,8'd176} : s = 308;
	{8'd132,8'd177} : s = 309;
	{8'd132,8'd178} : s = 310;
	{8'd132,8'd179} : s = 311;
	{8'd132,8'd180} : s = 312;
	{8'd132,8'd181} : s = 313;
	{8'd132,8'd182} : s = 314;
	{8'd132,8'd183} : s = 315;
	{8'd132,8'd184} : s = 316;
	{8'd132,8'd185} : s = 317;
	{8'd132,8'd186} : s = 318;
	{8'd132,8'd187} : s = 319;
	{8'd132,8'd188} : s = 320;
	{8'd132,8'd189} : s = 321;
	{8'd132,8'd190} : s = 322;
	{8'd132,8'd191} : s = 323;
	{8'd132,8'd192} : s = 324;
	{8'd132,8'd193} : s = 325;
	{8'd132,8'd194} : s = 326;
	{8'd132,8'd195} : s = 327;
	{8'd132,8'd196} : s = 328;
	{8'd132,8'd197} : s = 329;
	{8'd132,8'd198} : s = 330;
	{8'd132,8'd199} : s = 331;
	{8'd132,8'd200} : s = 332;
	{8'd132,8'd201} : s = 333;
	{8'd132,8'd202} : s = 334;
	{8'd132,8'd203} : s = 335;
	{8'd132,8'd204} : s = 336;
	{8'd132,8'd205} : s = 337;
	{8'd132,8'd206} : s = 338;
	{8'd132,8'd207} : s = 339;
	{8'd132,8'd208} : s = 340;
	{8'd132,8'd209} : s = 341;
	{8'd132,8'd210} : s = 342;
	{8'd132,8'd211} : s = 343;
	{8'd132,8'd212} : s = 344;
	{8'd132,8'd213} : s = 345;
	{8'd132,8'd214} : s = 346;
	{8'd132,8'd215} : s = 347;
	{8'd132,8'd216} : s = 348;
	{8'd132,8'd217} : s = 349;
	{8'd132,8'd218} : s = 350;
	{8'd132,8'd219} : s = 351;
	{8'd132,8'd220} : s = 352;
	{8'd132,8'd221} : s = 353;
	{8'd132,8'd222} : s = 354;
	{8'd132,8'd223} : s = 355;
	{8'd132,8'd224} : s = 356;
	{8'd132,8'd225} : s = 357;
	{8'd132,8'd226} : s = 358;
	{8'd132,8'd227} : s = 359;
	{8'd132,8'd228} : s = 360;
	{8'd132,8'd229} : s = 361;
	{8'd132,8'd230} : s = 362;
	{8'd132,8'd231} : s = 363;
	{8'd132,8'd232} : s = 364;
	{8'd132,8'd233} : s = 365;
	{8'd132,8'd234} : s = 366;
	{8'd132,8'd235} : s = 367;
	{8'd132,8'd236} : s = 368;
	{8'd132,8'd237} : s = 369;
	{8'd132,8'd238} : s = 370;
	{8'd132,8'd239} : s = 371;
	{8'd132,8'd240} : s = 372;
	{8'd132,8'd241} : s = 373;
	{8'd132,8'd242} : s = 374;
	{8'd132,8'd243} : s = 375;
	{8'd132,8'd244} : s = 376;
	{8'd132,8'd245} : s = 377;
	{8'd132,8'd246} : s = 378;
	{8'd132,8'd247} : s = 379;
	{8'd132,8'd248} : s = 380;
	{8'd132,8'd249} : s = 381;
	{8'd132,8'd250} : s = 382;
	{8'd132,8'd251} : s = 383;
	{8'd132,8'd252} : s = 384;
	{8'd132,8'd253} : s = 385;
	{8'd132,8'd254} : s = 386;
	{8'd132,8'd255} : s = 387;
	{8'd133,8'd0} : s = 133;
	{8'd133,8'd1} : s = 134;
	{8'd133,8'd2} : s = 135;
	{8'd133,8'd3} : s = 136;
	{8'd133,8'd4} : s = 137;
	{8'd133,8'd5} : s = 138;
	{8'd133,8'd6} : s = 139;
	{8'd133,8'd7} : s = 140;
	{8'd133,8'd8} : s = 141;
	{8'd133,8'd9} : s = 142;
	{8'd133,8'd10} : s = 143;
	{8'd133,8'd11} : s = 144;
	{8'd133,8'd12} : s = 145;
	{8'd133,8'd13} : s = 146;
	{8'd133,8'd14} : s = 147;
	{8'd133,8'd15} : s = 148;
	{8'd133,8'd16} : s = 149;
	{8'd133,8'd17} : s = 150;
	{8'd133,8'd18} : s = 151;
	{8'd133,8'd19} : s = 152;
	{8'd133,8'd20} : s = 153;
	{8'd133,8'd21} : s = 154;
	{8'd133,8'd22} : s = 155;
	{8'd133,8'd23} : s = 156;
	{8'd133,8'd24} : s = 157;
	{8'd133,8'd25} : s = 158;
	{8'd133,8'd26} : s = 159;
	{8'd133,8'd27} : s = 160;
	{8'd133,8'd28} : s = 161;
	{8'd133,8'd29} : s = 162;
	{8'd133,8'd30} : s = 163;
	{8'd133,8'd31} : s = 164;
	{8'd133,8'd32} : s = 165;
	{8'd133,8'd33} : s = 166;
	{8'd133,8'd34} : s = 167;
	{8'd133,8'd35} : s = 168;
	{8'd133,8'd36} : s = 169;
	{8'd133,8'd37} : s = 170;
	{8'd133,8'd38} : s = 171;
	{8'd133,8'd39} : s = 172;
	{8'd133,8'd40} : s = 173;
	{8'd133,8'd41} : s = 174;
	{8'd133,8'd42} : s = 175;
	{8'd133,8'd43} : s = 176;
	{8'd133,8'd44} : s = 177;
	{8'd133,8'd45} : s = 178;
	{8'd133,8'd46} : s = 179;
	{8'd133,8'd47} : s = 180;
	{8'd133,8'd48} : s = 181;
	{8'd133,8'd49} : s = 182;
	{8'd133,8'd50} : s = 183;
	{8'd133,8'd51} : s = 184;
	{8'd133,8'd52} : s = 185;
	{8'd133,8'd53} : s = 186;
	{8'd133,8'd54} : s = 187;
	{8'd133,8'd55} : s = 188;
	{8'd133,8'd56} : s = 189;
	{8'd133,8'd57} : s = 190;
	{8'd133,8'd58} : s = 191;
	{8'd133,8'd59} : s = 192;
	{8'd133,8'd60} : s = 193;
	{8'd133,8'd61} : s = 194;
	{8'd133,8'd62} : s = 195;
	{8'd133,8'd63} : s = 196;
	{8'd133,8'd64} : s = 197;
	{8'd133,8'd65} : s = 198;
	{8'd133,8'd66} : s = 199;
	{8'd133,8'd67} : s = 200;
	{8'd133,8'd68} : s = 201;
	{8'd133,8'd69} : s = 202;
	{8'd133,8'd70} : s = 203;
	{8'd133,8'd71} : s = 204;
	{8'd133,8'd72} : s = 205;
	{8'd133,8'd73} : s = 206;
	{8'd133,8'd74} : s = 207;
	{8'd133,8'd75} : s = 208;
	{8'd133,8'd76} : s = 209;
	{8'd133,8'd77} : s = 210;
	{8'd133,8'd78} : s = 211;
	{8'd133,8'd79} : s = 212;
	{8'd133,8'd80} : s = 213;
	{8'd133,8'd81} : s = 214;
	{8'd133,8'd82} : s = 215;
	{8'd133,8'd83} : s = 216;
	{8'd133,8'd84} : s = 217;
	{8'd133,8'd85} : s = 218;
	{8'd133,8'd86} : s = 219;
	{8'd133,8'd87} : s = 220;
	{8'd133,8'd88} : s = 221;
	{8'd133,8'd89} : s = 222;
	{8'd133,8'd90} : s = 223;
	{8'd133,8'd91} : s = 224;
	{8'd133,8'd92} : s = 225;
	{8'd133,8'd93} : s = 226;
	{8'd133,8'd94} : s = 227;
	{8'd133,8'd95} : s = 228;
	{8'd133,8'd96} : s = 229;
	{8'd133,8'd97} : s = 230;
	{8'd133,8'd98} : s = 231;
	{8'd133,8'd99} : s = 232;
	{8'd133,8'd100} : s = 233;
	{8'd133,8'd101} : s = 234;
	{8'd133,8'd102} : s = 235;
	{8'd133,8'd103} : s = 236;
	{8'd133,8'd104} : s = 237;
	{8'd133,8'd105} : s = 238;
	{8'd133,8'd106} : s = 239;
	{8'd133,8'd107} : s = 240;
	{8'd133,8'd108} : s = 241;
	{8'd133,8'd109} : s = 242;
	{8'd133,8'd110} : s = 243;
	{8'd133,8'd111} : s = 244;
	{8'd133,8'd112} : s = 245;
	{8'd133,8'd113} : s = 246;
	{8'd133,8'd114} : s = 247;
	{8'd133,8'd115} : s = 248;
	{8'd133,8'd116} : s = 249;
	{8'd133,8'd117} : s = 250;
	{8'd133,8'd118} : s = 251;
	{8'd133,8'd119} : s = 252;
	{8'd133,8'd120} : s = 253;
	{8'd133,8'd121} : s = 254;
	{8'd133,8'd122} : s = 255;
	{8'd133,8'd123} : s = 256;
	{8'd133,8'd124} : s = 257;
	{8'd133,8'd125} : s = 258;
	{8'd133,8'd126} : s = 259;
	{8'd133,8'd127} : s = 260;
	{8'd133,8'd128} : s = 261;
	{8'd133,8'd129} : s = 262;
	{8'd133,8'd130} : s = 263;
	{8'd133,8'd131} : s = 264;
	{8'd133,8'd132} : s = 265;
	{8'd133,8'd133} : s = 266;
	{8'd133,8'd134} : s = 267;
	{8'd133,8'd135} : s = 268;
	{8'd133,8'd136} : s = 269;
	{8'd133,8'd137} : s = 270;
	{8'd133,8'd138} : s = 271;
	{8'd133,8'd139} : s = 272;
	{8'd133,8'd140} : s = 273;
	{8'd133,8'd141} : s = 274;
	{8'd133,8'd142} : s = 275;
	{8'd133,8'd143} : s = 276;
	{8'd133,8'd144} : s = 277;
	{8'd133,8'd145} : s = 278;
	{8'd133,8'd146} : s = 279;
	{8'd133,8'd147} : s = 280;
	{8'd133,8'd148} : s = 281;
	{8'd133,8'd149} : s = 282;
	{8'd133,8'd150} : s = 283;
	{8'd133,8'd151} : s = 284;
	{8'd133,8'd152} : s = 285;
	{8'd133,8'd153} : s = 286;
	{8'd133,8'd154} : s = 287;
	{8'd133,8'd155} : s = 288;
	{8'd133,8'd156} : s = 289;
	{8'd133,8'd157} : s = 290;
	{8'd133,8'd158} : s = 291;
	{8'd133,8'd159} : s = 292;
	{8'd133,8'd160} : s = 293;
	{8'd133,8'd161} : s = 294;
	{8'd133,8'd162} : s = 295;
	{8'd133,8'd163} : s = 296;
	{8'd133,8'd164} : s = 297;
	{8'd133,8'd165} : s = 298;
	{8'd133,8'd166} : s = 299;
	{8'd133,8'd167} : s = 300;
	{8'd133,8'd168} : s = 301;
	{8'd133,8'd169} : s = 302;
	{8'd133,8'd170} : s = 303;
	{8'd133,8'd171} : s = 304;
	{8'd133,8'd172} : s = 305;
	{8'd133,8'd173} : s = 306;
	{8'd133,8'd174} : s = 307;
	{8'd133,8'd175} : s = 308;
	{8'd133,8'd176} : s = 309;
	{8'd133,8'd177} : s = 310;
	{8'd133,8'd178} : s = 311;
	{8'd133,8'd179} : s = 312;
	{8'd133,8'd180} : s = 313;
	{8'd133,8'd181} : s = 314;
	{8'd133,8'd182} : s = 315;
	{8'd133,8'd183} : s = 316;
	{8'd133,8'd184} : s = 317;
	{8'd133,8'd185} : s = 318;
	{8'd133,8'd186} : s = 319;
	{8'd133,8'd187} : s = 320;
	{8'd133,8'd188} : s = 321;
	{8'd133,8'd189} : s = 322;
	{8'd133,8'd190} : s = 323;
	{8'd133,8'd191} : s = 324;
	{8'd133,8'd192} : s = 325;
	{8'd133,8'd193} : s = 326;
	{8'd133,8'd194} : s = 327;
	{8'd133,8'd195} : s = 328;
	{8'd133,8'd196} : s = 329;
	{8'd133,8'd197} : s = 330;
	{8'd133,8'd198} : s = 331;
	{8'd133,8'd199} : s = 332;
	{8'd133,8'd200} : s = 333;
	{8'd133,8'd201} : s = 334;
	{8'd133,8'd202} : s = 335;
	{8'd133,8'd203} : s = 336;
	{8'd133,8'd204} : s = 337;
	{8'd133,8'd205} : s = 338;
	{8'd133,8'd206} : s = 339;
	{8'd133,8'd207} : s = 340;
	{8'd133,8'd208} : s = 341;
	{8'd133,8'd209} : s = 342;
	{8'd133,8'd210} : s = 343;
	{8'd133,8'd211} : s = 344;
	{8'd133,8'd212} : s = 345;
	{8'd133,8'd213} : s = 346;
	{8'd133,8'd214} : s = 347;
	{8'd133,8'd215} : s = 348;
	{8'd133,8'd216} : s = 349;
	{8'd133,8'd217} : s = 350;
	{8'd133,8'd218} : s = 351;
	{8'd133,8'd219} : s = 352;
	{8'd133,8'd220} : s = 353;
	{8'd133,8'd221} : s = 354;
	{8'd133,8'd222} : s = 355;
	{8'd133,8'd223} : s = 356;
	{8'd133,8'd224} : s = 357;
	{8'd133,8'd225} : s = 358;
	{8'd133,8'd226} : s = 359;
	{8'd133,8'd227} : s = 360;
	{8'd133,8'd228} : s = 361;
	{8'd133,8'd229} : s = 362;
	{8'd133,8'd230} : s = 363;
	{8'd133,8'd231} : s = 364;
	{8'd133,8'd232} : s = 365;
	{8'd133,8'd233} : s = 366;
	{8'd133,8'd234} : s = 367;
	{8'd133,8'd235} : s = 368;
	{8'd133,8'd236} : s = 369;
	{8'd133,8'd237} : s = 370;
	{8'd133,8'd238} : s = 371;
	{8'd133,8'd239} : s = 372;
	{8'd133,8'd240} : s = 373;
	{8'd133,8'd241} : s = 374;
	{8'd133,8'd242} : s = 375;
	{8'd133,8'd243} : s = 376;
	{8'd133,8'd244} : s = 377;
	{8'd133,8'd245} : s = 378;
	{8'd133,8'd246} : s = 379;
	{8'd133,8'd247} : s = 380;
	{8'd133,8'd248} : s = 381;
	{8'd133,8'd249} : s = 382;
	{8'd133,8'd250} : s = 383;
	{8'd133,8'd251} : s = 384;
	{8'd133,8'd252} : s = 385;
	{8'd133,8'd253} : s = 386;
	{8'd133,8'd254} : s = 387;
	{8'd133,8'd255} : s = 388;
	{8'd134,8'd0} : s = 134;
	{8'd134,8'd1} : s = 135;
	{8'd134,8'd2} : s = 136;
	{8'd134,8'd3} : s = 137;
	{8'd134,8'd4} : s = 138;
	{8'd134,8'd5} : s = 139;
	{8'd134,8'd6} : s = 140;
	{8'd134,8'd7} : s = 141;
	{8'd134,8'd8} : s = 142;
	{8'd134,8'd9} : s = 143;
	{8'd134,8'd10} : s = 144;
	{8'd134,8'd11} : s = 145;
	{8'd134,8'd12} : s = 146;
	{8'd134,8'd13} : s = 147;
	{8'd134,8'd14} : s = 148;
	{8'd134,8'd15} : s = 149;
	{8'd134,8'd16} : s = 150;
	{8'd134,8'd17} : s = 151;
	{8'd134,8'd18} : s = 152;
	{8'd134,8'd19} : s = 153;
	{8'd134,8'd20} : s = 154;
	{8'd134,8'd21} : s = 155;
	{8'd134,8'd22} : s = 156;
	{8'd134,8'd23} : s = 157;
	{8'd134,8'd24} : s = 158;
	{8'd134,8'd25} : s = 159;
	{8'd134,8'd26} : s = 160;
	{8'd134,8'd27} : s = 161;
	{8'd134,8'd28} : s = 162;
	{8'd134,8'd29} : s = 163;
	{8'd134,8'd30} : s = 164;
	{8'd134,8'd31} : s = 165;
	{8'd134,8'd32} : s = 166;
	{8'd134,8'd33} : s = 167;
	{8'd134,8'd34} : s = 168;
	{8'd134,8'd35} : s = 169;
	{8'd134,8'd36} : s = 170;
	{8'd134,8'd37} : s = 171;
	{8'd134,8'd38} : s = 172;
	{8'd134,8'd39} : s = 173;
	{8'd134,8'd40} : s = 174;
	{8'd134,8'd41} : s = 175;
	{8'd134,8'd42} : s = 176;
	{8'd134,8'd43} : s = 177;
	{8'd134,8'd44} : s = 178;
	{8'd134,8'd45} : s = 179;
	{8'd134,8'd46} : s = 180;
	{8'd134,8'd47} : s = 181;
	{8'd134,8'd48} : s = 182;
	{8'd134,8'd49} : s = 183;
	{8'd134,8'd50} : s = 184;
	{8'd134,8'd51} : s = 185;
	{8'd134,8'd52} : s = 186;
	{8'd134,8'd53} : s = 187;
	{8'd134,8'd54} : s = 188;
	{8'd134,8'd55} : s = 189;
	{8'd134,8'd56} : s = 190;
	{8'd134,8'd57} : s = 191;
	{8'd134,8'd58} : s = 192;
	{8'd134,8'd59} : s = 193;
	{8'd134,8'd60} : s = 194;
	{8'd134,8'd61} : s = 195;
	{8'd134,8'd62} : s = 196;
	{8'd134,8'd63} : s = 197;
	{8'd134,8'd64} : s = 198;
	{8'd134,8'd65} : s = 199;
	{8'd134,8'd66} : s = 200;
	{8'd134,8'd67} : s = 201;
	{8'd134,8'd68} : s = 202;
	{8'd134,8'd69} : s = 203;
	{8'd134,8'd70} : s = 204;
	{8'd134,8'd71} : s = 205;
	{8'd134,8'd72} : s = 206;
	{8'd134,8'd73} : s = 207;
	{8'd134,8'd74} : s = 208;
	{8'd134,8'd75} : s = 209;
	{8'd134,8'd76} : s = 210;
	{8'd134,8'd77} : s = 211;
	{8'd134,8'd78} : s = 212;
	{8'd134,8'd79} : s = 213;
	{8'd134,8'd80} : s = 214;
	{8'd134,8'd81} : s = 215;
	{8'd134,8'd82} : s = 216;
	{8'd134,8'd83} : s = 217;
	{8'd134,8'd84} : s = 218;
	{8'd134,8'd85} : s = 219;
	{8'd134,8'd86} : s = 220;
	{8'd134,8'd87} : s = 221;
	{8'd134,8'd88} : s = 222;
	{8'd134,8'd89} : s = 223;
	{8'd134,8'd90} : s = 224;
	{8'd134,8'd91} : s = 225;
	{8'd134,8'd92} : s = 226;
	{8'd134,8'd93} : s = 227;
	{8'd134,8'd94} : s = 228;
	{8'd134,8'd95} : s = 229;
	{8'd134,8'd96} : s = 230;
	{8'd134,8'd97} : s = 231;
	{8'd134,8'd98} : s = 232;
	{8'd134,8'd99} : s = 233;
	{8'd134,8'd100} : s = 234;
	{8'd134,8'd101} : s = 235;
	{8'd134,8'd102} : s = 236;
	{8'd134,8'd103} : s = 237;
	{8'd134,8'd104} : s = 238;
	{8'd134,8'd105} : s = 239;
	{8'd134,8'd106} : s = 240;
	{8'd134,8'd107} : s = 241;
	{8'd134,8'd108} : s = 242;
	{8'd134,8'd109} : s = 243;
	{8'd134,8'd110} : s = 244;
	{8'd134,8'd111} : s = 245;
	{8'd134,8'd112} : s = 246;
	{8'd134,8'd113} : s = 247;
	{8'd134,8'd114} : s = 248;
	{8'd134,8'd115} : s = 249;
	{8'd134,8'd116} : s = 250;
	{8'd134,8'd117} : s = 251;
	{8'd134,8'd118} : s = 252;
	{8'd134,8'd119} : s = 253;
	{8'd134,8'd120} : s = 254;
	{8'd134,8'd121} : s = 255;
	{8'd134,8'd122} : s = 256;
	{8'd134,8'd123} : s = 257;
	{8'd134,8'd124} : s = 258;
	{8'd134,8'd125} : s = 259;
	{8'd134,8'd126} : s = 260;
	{8'd134,8'd127} : s = 261;
	{8'd134,8'd128} : s = 262;
	{8'd134,8'd129} : s = 263;
	{8'd134,8'd130} : s = 264;
	{8'd134,8'd131} : s = 265;
	{8'd134,8'd132} : s = 266;
	{8'd134,8'd133} : s = 267;
	{8'd134,8'd134} : s = 268;
	{8'd134,8'd135} : s = 269;
	{8'd134,8'd136} : s = 270;
	{8'd134,8'd137} : s = 271;
	{8'd134,8'd138} : s = 272;
	{8'd134,8'd139} : s = 273;
	{8'd134,8'd140} : s = 274;
	{8'd134,8'd141} : s = 275;
	{8'd134,8'd142} : s = 276;
	{8'd134,8'd143} : s = 277;
	{8'd134,8'd144} : s = 278;
	{8'd134,8'd145} : s = 279;
	{8'd134,8'd146} : s = 280;
	{8'd134,8'd147} : s = 281;
	{8'd134,8'd148} : s = 282;
	{8'd134,8'd149} : s = 283;
	{8'd134,8'd150} : s = 284;
	{8'd134,8'd151} : s = 285;
	{8'd134,8'd152} : s = 286;
	{8'd134,8'd153} : s = 287;
	{8'd134,8'd154} : s = 288;
	{8'd134,8'd155} : s = 289;
	{8'd134,8'd156} : s = 290;
	{8'd134,8'd157} : s = 291;
	{8'd134,8'd158} : s = 292;
	{8'd134,8'd159} : s = 293;
	{8'd134,8'd160} : s = 294;
	{8'd134,8'd161} : s = 295;
	{8'd134,8'd162} : s = 296;
	{8'd134,8'd163} : s = 297;
	{8'd134,8'd164} : s = 298;
	{8'd134,8'd165} : s = 299;
	{8'd134,8'd166} : s = 300;
	{8'd134,8'd167} : s = 301;
	{8'd134,8'd168} : s = 302;
	{8'd134,8'd169} : s = 303;
	{8'd134,8'd170} : s = 304;
	{8'd134,8'd171} : s = 305;
	{8'd134,8'd172} : s = 306;
	{8'd134,8'd173} : s = 307;
	{8'd134,8'd174} : s = 308;
	{8'd134,8'd175} : s = 309;
	{8'd134,8'd176} : s = 310;
	{8'd134,8'd177} : s = 311;
	{8'd134,8'd178} : s = 312;
	{8'd134,8'd179} : s = 313;
	{8'd134,8'd180} : s = 314;
	{8'd134,8'd181} : s = 315;
	{8'd134,8'd182} : s = 316;
	{8'd134,8'd183} : s = 317;
	{8'd134,8'd184} : s = 318;
	{8'd134,8'd185} : s = 319;
	{8'd134,8'd186} : s = 320;
	{8'd134,8'd187} : s = 321;
	{8'd134,8'd188} : s = 322;
	{8'd134,8'd189} : s = 323;
	{8'd134,8'd190} : s = 324;
	{8'd134,8'd191} : s = 325;
	{8'd134,8'd192} : s = 326;
	{8'd134,8'd193} : s = 327;
	{8'd134,8'd194} : s = 328;
	{8'd134,8'd195} : s = 329;
	{8'd134,8'd196} : s = 330;
	{8'd134,8'd197} : s = 331;
	{8'd134,8'd198} : s = 332;
	{8'd134,8'd199} : s = 333;
	{8'd134,8'd200} : s = 334;
	{8'd134,8'd201} : s = 335;
	{8'd134,8'd202} : s = 336;
	{8'd134,8'd203} : s = 337;
	{8'd134,8'd204} : s = 338;
	{8'd134,8'd205} : s = 339;
	{8'd134,8'd206} : s = 340;
	{8'd134,8'd207} : s = 341;
	{8'd134,8'd208} : s = 342;
	{8'd134,8'd209} : s = 343;
	{8'd134,8'd210} : s = 344;
	{8'd134,8'd211} : s = 345;
	{8'd134,8'd212} : s = 346;
	{8'd134,8'd213} : s = 347;
	{8'd134,8'd214} : s = 348;
	{8'd134,8'd215} : s = 349;
	{8'd134,8'd216} : s = 350;
	{8'd134,8'd217} : s = 351;
	{8'd134,8'd218} : s = 352;
	{8'd134,8'd219} : s = 353;
	{8'd134,8'd220} : s = 354;
	{8'd134,8'd221} : s = 355;
	{8'd134,8'd222} : s = 356;
	{8'd134,8'd223} : s = 357;
	{8'd134,8'd224} : s = 358;
	{8'd134,8'd225} : s = 359;
	{8'd134,8'd226} : s = 360;
	{8'd134,8'd227} : s = 361;
	{8'd134,8'd228} : s = 362;
	{8'd134,8'd229} : s = 363;
	{8'd134,8'd230} : s = 364;
	{8'd134,8'd231} : s = 365;
	{8'd134,8'd232} : s = 366;
	{8'd134,8'd233} : s = 367;
	{8'd134,8'd234} : s = 368;
	{8'd134,8'd235} : s = 369;
	{8'd134,8'd236} : s = 370;
	{8'd134,8'd237} : s = 371;
	{8'd134,8'd238} : s = 372;
	{8'd134,8'd239} : s = 373;
	{8'd134,8'd240} : s = 374;
	{8'd134,8'd241} : s = 375;
	{8'd134,8'd242} : s = 376;
	{8'd134,8'd243} : s = 377;
	{8'd134,8'd244} : s = 378;
	{8'd134,8'd245} : s = 379;
	{8'd134,8'd246} : s = 380;
	{8'd134,8'd247} : s = 381;
	{8'd134,8'd248} : s = 382;
	{8'd134,8'd249} : s = 383;
	{8'd134,8'd250} : s = 384;
	{8'd134,8'd251} : s = 385;
	{8'd134,8'd252} : s = 386;
	{8'd134,8'd253} : s = 387;
	{8'd134,8'd254} : s = 388;
	{8'd134,8'd255} : s = 389;
	{8'd135,8'd0} : s = 135;
	{8'd135,8'd1} : s = 136;
	{8'd135,8'd2} : s = 137;
	{8'd135,8'd3} : s = 138;
	{8'd135,8'd4} : s = 139;
	{8'd135,8'd5} : s = 140;
	{8'd135,8'd6} : s = 141;
	{8'd135,8'd7} : s = 142;
	{8'd135,8'd8} : s = 143;
	{8'd135,8'd9} : s = 144;
	{8'd135,8'd10} : s = 145;
	{8'd135,8'd11} : s = 146;
	{8'd135,8'd12} : s = 147;
	{8'd135,8'd13} : s = 148;
	{8'd135,8'd14} : s = 149;
	{8'd135,8'd15} : s = 150;
	{8'd135,8'd16} : s = 151;
	{8'd135,8'd17} : s = 152;
	{8'd135,8'd18} : s = 153;
	{8'd135,8'd19} : s = 154;
	{8'd135,8'd20} : s = 155;
	{8'd135,8'd21} : s = 156;
	{8'd135,8'd22} : s = 157;
	{8'd135,8'd23} : s = 158;
	{8'd135,8'd24} : s = 159;
	{8'd135,8'd25} : s = 160;
	{8'd135,8'd26} : s = 161;
	{8'd135,8'd27} : s = 162;
	{8'd135,8'd28} : s = 163;
	{8'd135,8'd29} : s = 164;
	{8'd135,8'd30} : s = 165;
	{8'd135,8'd31} : s = 166;
	{8'd135,8'd32} : s = 167;
	{8'd135,8'd33} : s = 168;
	{8'd135,8'd34} : s = 169;
	{8'd135,8'd35} : s = 170;
	{8'd135,8'd36} : s = 171;
	{8'd135,8'd37} : s = 172;
	{8'd135,8'd38} : s = 173;
	{8'd135,8'd39} : s = 174;
	{8'd135,8'd40} : s = 175;
	{8'd135,8'd41} : s = 176;
	{8'd135,8'd42} : s = 177;
	{8'd135,8'd43} : s = 178;
	{8'd135,8'd44} : s = 179;
	{8'd135,8'd45} : s = 180;
	{8'd135,8'd46} : s = 181;
	{8'd135,8'd47} : s = 182;
	{8'd135,8'd48} : s = 183;
	{8'd135,8'd49} : s = 184;
	{8'd135,8'd50} : s = 185;
	{8'd135,8'd51} : s = 186;
	{8'd135,8'd52} : s = 187;
	{8'd135,8'd53} : s = 188;
	{8'd135,8'd54} : s = 189;
	{8'd135,8'd55} : s = 190;
	{8'd135,8'd56} : s = 191;
	{8'd135,8'd57} : s = 192;
	{8'd135,8'd58} : s = 193;
	{8'd135,8'd59} : s = 194;
	{8'd135,8'd60} : s = 195;
	{8'd135,8'd61} : s = 196;
	{8'd135,8'd62} : s = 197;
	{8'd135,8'd63} : s = 198;
	{8'd135,8'd64} : s = 199;
	{8'd135,8'd65} : s = 200;
	{8'd135,8'd66} : s = 201;
	{8'd135,8'd67} : s = 202;
	{8'd135,8'd68} : s = 203;
	{8'd135,8'd69} : s = 204;
	{8'd135,8'd70} : s = 205;
	{8'd135,8'd71} : s = 206;
	{8'd135,8'd72} : s = 207;
	{8'd135,8'd73} : s = 208;
	{8'd135,8'd74} : s = 209;
	{8'd135,8'd75} : s = 210;
	{8'd135,8'd76} : s = 211;
	{8'd135,8'd77} : s = 212;
	{8'd135,8'd78} : s = 213;
	{8'd135,8'd79} : s = 214;
	{8'd135,8'd80} : s = 215;
	{8'd135,8'd81} : s = 216;
	{8'd135,8'd82} : s = 217;
	{8'd135,8'd83} : s = 218;
	{8'd135,8'd84} : s = 219;
	{8'd135,8'd85} : s = 220;
	{8'd135,8'd86} : s = 221;
	{8'd135,8'd87} : s = 222;
	{8'd135,8'd88} : s = 223;
	{8'd135,8'd89} : s = 224;
	{8'd135,8'd90} : s = 225;
	{8'd135,8'd91} : s = 226;
	{8'd135,8'd92} : s = 227;
	{8'd135,8'd93} : s = 228;
	{8'd135,8'd94} : s = 229;
	{8'd135,8'd95} : s = 230;
	{8'd135,8'd96} : s = 231;
	{8'd135,8'd97} : s = 232;
	{8'd135,8'd98} : s = 233;
	{8'd135,8'd99} : s = 234;
	{8'd135,8'd100} : s = 235;
	{8'd135,8'd101} : s = 236;
	{8'd135,8'd102} : s = 237;
	{8'd135,8'd103} : s = 238;
	{8'd135,8'd104} : s = 239;
	{8'd135,8'd105} : s = 240;
	{8'd135,8'd106} : s = 241;
	{8'd135,8'd107} : s = 242;
	{8'd135,8'd108} : s = 243;
	{8'd135,8'd109} : s = 244;
	{8'd135,8'd110} : s = 245;
	{8'd135,8'd111} : s = 246;
	{8'd135,8'd112} : s = 247;
	{8'd135,8'd113} : s = 248;
	{8'd135,8'd114} : s = 249;
	{8'd135,8'd115} : s = 250;
	{8'd135,8'd116} : s = 251;
	{8'd135,8'd117} : s = 252;
	{8'd135,8'd118} : s = 253;
	{8'd135,8'd119} : s = 254;
	{8'd135,8'd120} : s = 255;
	{8'd135,8'd121} : s = 256;
	{8'd135,8'd122} : s = 257;
	{8'd135,8'd123} : s = 258;
	{8'd135,8'd124} : s = 259;
	{8'd135,8'd125} : s = 260;
	{8'd135,8'd126} : s = 261;
	{8'd135,8'd127} : s = 262;
	{8'd135,8'd128} : s = 263;
	{8'd135,8'd129} : s = 264;
	{8'd135,8'd130} : s = 265;
	{8'd135,8'd131} : s = 266;
	{8'd135,8'd132} : s = 267;
	{8'd135,8'd133} : s = 268;
	{8'd135,8'd134} : s = 269;
	{8'd135,8'd135} : s = 270;
	{8'd135,8'd136} : s = 271;
	{8'd135,8'd137} : s = 272;
	{8'd135,8'd138} : s = 273;
	{8'd135,8'd139} : s = 274;
	{8'd135,8'd140} : s = 275;
	{8'd135,8'd141} : s = 276;
	{8'd135,8'd142} : s = 277;
	{8'd135,8'd143} : s = 278;
	{8'd135,8'd144} : s = 279;
	{8'd135,8'd145} : s = 280;
	{8'd135,8'd146} : s = 281;
	{8'd135,8'd147} : s = 282;
	{8'd135,8'd148} : s = 283;
	{8'd135,8'd149} : s = 284;
	{8'd135,8'd150} : s = 285;
	{8'd135,8'd151} : s = 286;
	{8'd135,8'd152} : s = 287;
	{8'd135,8'd153} : s = 288;
	{8'd135,8'd154} : s = 289;
	{8'd135,8'd155} : s = 290;
	{8'd135,8'd156} : s = 291;
	{8'd135,8'd157} : s = 292;
	{8'd135,8'd158} : s = 293;
	{8'd135,8'd159} : s = 294;
	{8'd135,8'd160} : s = 295;
	{8'd135,8'd161} : s = 296;
	{8'd135,8'd162} : s = 297;
	{8'd135,8'd163} : s = 298;
	{8'd135,8'd164} : s = 299;
	{8'd135,8'd165} : s = 300;
	{8'd135,8'd166} : s = 301;
	{8'd135,8'd167} : s = 302;
	{8'd135,8'd168} : s = 303;
	{8'd135,8'd169} : s = 304;
	{8'd135,8'd170} : s = 305;
	{8'd135,8'd171} : s = 306;
	{8'd135,8'd172} : s = 307;
	{8'd135,8'd173} : s = 308;
	{8'd135,8'd174} : s = 309;
	{8'd135,8'd175} : s = 310;
	{8'd135,8'd176} : s = 311;
	{8'd135,8'd177} : s = 312;
	{8'd135,8'd178} : s = 313;
	{8'd135,8'd179} : s = 314;
	{8'd135,8'd180} : s = 315;
	{8'd135,8'd181} : s = 316;
	{8'd135,8'd182} : s = 317;
	{8'd135,8'd183} : s = 318;
	{8'd135,8'd184} : s = 319;
	{8'd135,8'd185} : s = 320;
	{8'd135,8'd186} : s = 321;
	{8'd135,8'd187} : s = 322;
	{8'd135,8'd188} : s = 323;
	{8'd135,8'd189} : s = 324;
	{8'd135,8'd190} : s = 325;
	{8'd135,8'd191} : s = 326;
	{8'd135,8'd192} : s = 327;
	{8'd135,8'd193} : s = 328;
	{8'd135,8'd194} : s = 329;
	{8'd135,8'd195} : s = 330;
	{8'd135,8'd196} : s = 331;
	{8'd135,8'd197} : s = 332;
	{8'd135,8'd198} : s = 333;
	{8'd135,8'd199} : s = 334;
	{8'd135,8'd200} : s = 335;
	{8'd135,8'd201} : s = 336;
	{8'd135,8'd202} : s = 337;
	{8'd135,8'd203} : s = 338;
	{8'd135,8'd204} : s = 339;
	{8'd135,8'd205} : s = 340;
	{8'd135,8'd206} : s = 341;
	{8'd135,8'd207} : s = 342;
	{8'd135,8'd208} : s = 343;
	{8'd135,8'd209} : s = 344;
	{8'd135,8'd210} : s = 345;
	{8'd135,8'd211} : s = 346;
	{8'd135,8'd212} : s = 347;
	{8'd135,8'd213} : s = 348;
	{8'd135,8'd214} : s = 349;
	{8'd135,8'd215} : s = 350;
	{8'd135,8'd216} : s = 351;
	{8'd135,8'd217} : s = 352;
	{8'd135,8'd218} : s = 353;
	{8'd135,8'd219} : s = 354;
	{8'd135,8'd220} : s = 355;
	{8'd135,8'd221} : s = 356;
	{8'd135,8'd222} : s = 357;
	{8'd135,8'd223} : s = 358;
	{8'd135,8'd224} : s = 359;
	{8'd135,8'd225} : s = 360;
	{8'd135,8'd226} : s = 361;
	{8'd135,8'd227} : s = 362;
	{8'd135,8'd228} : s = 363;
	{8'd135,8'd229} : s = 364;
	{8'd135,8'd230} : s = 365;
	{8'd135,8'd231} : s = 366;
	{8'd135,8'd232} : s = 367;
	{8'd135,8'd233} : s = 368;
	{8'd135,8'd234} : s = 369;
	{8'd135,8'd235} : s = 370;
	{8'd135,8'd236} : s = 371;
	{8'd135,8'd237} : s = 372;
	{8'd135,8'd238} : s = 373;
	{8'd135,8'd239} : s = 374;
	{8'd135,8'd240} : s = 375;
	{8'd135,8'd241} : s = 376;
	{8'd135,8'd242} : s = 377;
	{8'd135,8'd243} : s = 378;
	{8'd135,8'd244} : s = 379;
	{8'd135,8'd245} : s = 380;
	{8'd135,8'd246} : s = 381;
	{8'd135,8'd247} : s = 382;
	{8'd135,8'd248} : s = 383;
	{8'd135,8'd249} : s = 384;
	{8'd135,8'd250} : s = 385;
	{8'd135,8'd251} : s = 386;
	{8'd135,8'd252} : s = 387;
	{8'd135,8'd253} : s = 388;
	{8'd135,8'd254} : s = 389;
	{8'd135,8'd255} : s = 390;
	{8'd136,8'd0} : s = 136;
	{8'd136,8'd1} : s = 137;
	{8'd136,8'd2} : s = 138;
	{8'd136,8'd3} : s = 139;
	{8'd136,8'd4} : s = 140;
	{8'd136,8'd5} : s = 141;
	{8'd136,8'd6} : s = 142;
	{8'd136,8'd7} : s = 143;
	{8'd136,8'd8} : s = 144;
	{8'd136,8'd9} : s = 145;
	{8'd136,8'd10} : s = 146;
	{8'd136,8'd11} : s = 147;
	{8'd136,8'd12} : s = 148;
	{8'd136,8'd13} : s = 149;
	{8'd136,8'd14} : s = 150;
	{8'd136,8'd15} : s = 151;
	{8'd136,8'd16} : s = 152;
	{8'd136,8'd17} : s = 153;
	{8'd136,8'd18} : s = 154;
	{8'd136,8'd19} : s = 155;
	{8'd136,8'd20} : s = 156;
	{8'd136,8'd21} : s = 157;
	{8'd136,8'd22} : s = 158;
	{8'd136,8'd23} : s = 159;
	{8'd136,8'd24} : s = 160;
	{8'd136,8'd25} : s = 161;
	{8'd136,8'd26} : s = 162;
	{8'd136,8'd27} : s = 163;
	{8'd136,8'd28} : s = 164;
	{8'd136,8'd29} : s = 165;
	{8'd136,8'd30} : s = 166;
	{8'd136,8'd31} : s = 167;
	{8'd136,8'd32} : s = 168;
	{8'd136,8'd33} : s = 169;
	{8'd136,8'd34} : s = 170;
	{8'd136,8'd35} : s = 171;
	{8'd136,8'd36} : s = 172;
	{8'd136,8'd37} : s = 173;
	{8'd136,8'd38} : s = 174;
	{8'd136,8'd39} : s = 175;
	{8'd136,8'd40} : s = 176;
	{8'd136,8'd41} : s = 177;
	{8'd136,8'd42} : s = 178;
	{8'd136,8'd43} : s = 179;
	{8'd136,8'd44} : s = 180;
	{8'd136,8'd45} : s = 181;
	{8'd136,8'd46} : s = 182;
	{8'd136,8'd47} : s = 183;
	{8'd136,8'd48} : s = 184;
	{8'd136,8'd49} : s = 185;
	{8'd136,8'd50} : s = 186;
	{8'd136,8'd51} : s = 187;
	{8'd136,8'd52} : s = 188;
	{8'd136,8'd53} : s = 189;
	{8'd136,8'd54} : s = 190;
	{8'd136,8'd55} : s = 191;
	{8'd136,8'd56} : s = 192;
	{8'd136,8'd57} : s = 193;
	{8'd136,8'd58} : s = 194;
	{8'd136,8'd59} : s = 195;
	{8'd136,8'd60} : s = 196;
	{8'd136,8'd61} : s = 197;
	{8'd136,8'd62} : s = 198;
	{8'd136,8'd63} : s = 199;
	{8'd136,8'd64} : s = 200;
	{8'd136,8'd65} : s = 201;
	{8'd136,8'd66} : s = 202;
	{8'd136,8'd67} : s = 203;
	{8'd136,8'd68} : s = 204;
	{8'd136,8'd69} : s = 205;
	{8'd136,8'd70} : s = 206;
	{8'd136,8'd71} : s = 207;
	{8'd136,8'd72} : s = 208;
	{8'd136,8'd73} : s = 209;
	{8'd136,8'd74} : s = 210;
	{8'd136,8'd75} : s = 211;
	{8'd136,8'd76} : s = 212;
	{8'd136,8'd77} : s = 213;
	{8'd136,8'd78} : s = 214;
	{8'd136,8'd79} : s = 215;
	{8'd136,8'd80} : s = 216;
	{8'd136,8'd81} : s = 217;
	{8'd136,8'd82} : s = 218;
	{8'd136,8'd83} : s = 219;
	{8'd136,8'd84} : s = 220;
	{8'd136,8'd85} : s = 221;
	{8'd136,8'd86} : s = 222;
	{8'd136,8'd87} : s = 223;
	{8'd136,8'd88} : s = 224;
	{8'd136,8'd89} : s = 225;
	{8'd136,8'd90} : s = 226;
	{8'd136,8'd91} : s = 227;
	{8'd136,8'd92} : s = 228;
	{8'd136,8'd93} : s = 229;
	{8'd136,8'd94} : s = 230;
	{8'd136,8'd95} : s = 231;
	{8'd136,8'd96} : s = 232;
	{8'd136,8'd97} : s = 233;
	{8'd136,8'd98} : s = 234;
	{8'd136,8'd99} : s = 235;
	{8'd136,8'd100} : s = 236;
	{8'd136,8'd101} : s = 237;
	{8'd136,8'd102} : s = 238;
	{8'd136,8'd103} : s = 239;
	{8'd136,8'd104} : s = 240;
	{8'd136,8'd105} : s = 241;
	{8'd136,8'd106} : s = 242;
	{8'd136,8'd107} : s = 243;
	{8'd136,8'd108} : s = 244;
	{8'd136,8'd109} : s = 245;
	{8'd136,8'd110} : s = 246;
	{8'd136,8'd111} : s = 247;
	{8'd136,8'd112} : s = 248;
	{8'd136,8'd113} : s = 249;
	{8'd136,8'd114} : s = 250;
	{8'd136,8'd115} : s = 251;
	{8'd136,8'd116} : s = 252;
	{8'd136,8'd117} : s = 253;
	{8'd136,8'd118} : s = 254;
	{8'd136,8'd119} : s = 255;
	{8'd136,8'd120} : s = 256;
	{8'd136,8'd121} : s = 257;
	{8'd136,8'd122} : s = 258;
	{8'd136,8'd123} : s = 259;
	{8'd136,8'd124} : s = 260;
	{8'd136,8'd125} : s = 261;
	{8'd136,8'd126} : s = 262;
	{8'd136,8'd127} : s = 263;
	{8'd136,8'd128} : s = 264;
	{8'd136,8'd129} : s = 265;
	{8'd136,8'd130} : s = 266;
	{8'd136,8'd131} : s = 267;
	{8'd136,8'd132} : s = 268;
	{8'd136,8'd133} : s = 269;
	{8'd136,8'd134} : s = 270;
	{8'd136,8'd135} : s = 271;
	{8'd136,8'd136} : s = 272;
	{8'd136,8'd137} : s = 273;
	{8'd136,8'd138} : s = 274;
	{8'd136,8'd139} : s = 275;
	{8'd136,8'd140} : s = 276;
	{8'd136,8'd141} : s = 277;
	{8'd136,8'd142} : s = 278;
	{8'd136,8'd143} : s = 279;
	{8'd136,8'd144} : s = 280;
	{8'd136,8'd145} : s = 281;
	{8'd136,8'd146} : s = 282;
	{8'd136,8'd147} : s = 283;
	{8'd136,8'd148} : s = 284;
	{8'd136,8'd149} : s = 285;
	{8'd136,8'd150} : s = 286;
	{8'd136,8'd151} : s = 287;
	{8'd136,8'd152} : s = 288;
	{8'd136,8'd153} : s = 289;
	{8'd136,8'd154} : s = 290;
	{8'd136,8'd155} : s = 291;
	{8'd136,8'd156} : s = 292;
	{8'd136,8'd157} : s = 293;
	{8'd136,8'd158} : s = 294;
	{8'd136,8'd159} : s = 295;
	{8'd136,8'd160} : s = 296;
	{8'd136,8'd161} : s = 297;
	{8'd136,8'd162} : s = 298;
	{8'd136,8'd163} : s = 299;
	{8'd136,8'd164} : s = 300;
	{8'd136,8'd165} : s = 301;
	{8'd136,8'd166} : s = 302;
	{8'd136,8'd167} : s = 303;
	{8'd136,8'd168} : s = 304;
	{8'd136,8'd169} : s = 305;
	{8'd136,8'd170} : s = 306;
	{8'd136,8'd171} : s = 307;
	{8'd136,8'd172} : s = 308;
	{8'd136,8'd173} : s = 309;
	{8'd136,8'd174} : s = 310;
	{8'd136,8'd175} : s = 311;
	{8'd136,8'd176} : s = 312;
	{8'd136,8'd177} : s = 313;
	{8'd136,8'd178} : s = 314;
	{8'd136,8'd179} : s = 315;
	{8'd136,8'd180} : s = 316;
	{8'd136,8'd181} : s = 317;
	{8'd136,8'd182} : s = 318;
	{8'd136,8'd183} : s = 319;
	{8'd136,8'd184} : s = 320;
	{8'd136,8'd185} : s = 321;
	{8'd136,8'd186} : s = 322;
	{8'd136,8'd187} : s = 323;
	{8'd136,8'd188} : s = 324;
	{8'd136,8'd189} : s = 325;
	{8'd136,8'd190} : s = 326;
	{8'd136,8'd191} : s = 327;
	{8'd136,8'd192} : s = 328;
	{8'd136,8'd193} : s = 329;
	{8'd136,8'd194} : s = 330;
	{8'd136,8'd195} : s = 331;
	{8'd136,8'd196} : s = 332;
	{8'd136,8'd197} : s = 333;
	{8'd136,8'd198} : s = 334;
	{8'd136,8'd199} : s = 335;
	{8'd136,8'd200} : s = 336;
	{8'd136,8'd201} : s = 337;
	{8'd136,8'd202} : s = 338;
	{8'd136,8'd203} : s = 339;
	{8'd136,8'd204} : s = 340;
	{8'd136,8'd205} : s = 341;
	{8'd136,8'd206} : s = 342;
	{8'd136,8'd207} : s = 343;
	{8'd136,8'd208} : s = 344;
	{8'd136,8'd209} : s = 345;
	{8'd136,8'd210} : s = 346;
	{8'd136,8'd211} : s = 347;
	{8'd136,8'd212} : s = 348;
	{8'd136,8'd213} : s = 349;
	{8'd136,8'd214} : s = 350;
	{8'd136,8'd215} : s = 351;
	{8'd136,8'd216} : s = 352;
	{8'd136,8'd217} : s = 353;
	{8'd136,8'd218} : s = 354;
	{8'd136,8'd219} : s = 355;
	{8'd136,8'd220} : s = 356;
	{8'd136,8'd221} : s = 357;
	{8'd136,8'd222} : s = 358;
	{8'd136,8'd223} : s = 359;
	{8'd136,8'd224} : s = 360;
	{8'd136,8'd225} : s = 361;
	{8'd136,8'd226} : s = 362;
	{8'd136,8'd227} : s = 363;
	{8'd136,8'd228} : s = 364;
	{8'd136,8'd229} : s = 365;
	{8'd136,8'd230} : s = 366;
	{8'd136,8'd231} : s = 367;
	{8'd136,8'd232} : s = 368;
	{8'd136,8'd233} : s = 369;
	{8'd136,8'd234} : s = 370;
	{8'd136,8'd235} : s = 371;
	{8'd136,8'd236} : s = 372;
	{8'd136,8'd237} : s = 373;
	{8'd136,8'd238} : s = 374;
	{8'd136,8'd239} : s = 375;
	{8'd136,8'd240} : s = 376;
	{8'd136,8'd241} : s = 377;
	{8'd136,8'd242} : s = 378;
	{8'd136,8'd243} : s = 379;
	{8'd136,8'd244} : s = 380;
	{8'd136,8'd245} : s = 381;
	{8'd136,8'd246} : s = 382;
	{8'd136,8'd247} : s = 383;
	{8'd136,8'd248} : s = 384;
	{8'd136,8'd249} : s = 385;
	{8'd136,8'd250} : s = 386;
	{8'd136,8'd251} : s = 387;
	{8'd136,8'd252} : s = 388;
	{8'd136,8'd253} : s = 389;
	{8'd136,8'd254} : s = 390;
	{8'd136,8'd255} : s = 391;
	{8'd137,8'd0} : s = 137;
	{8'd137,8'd1} : s = 138;
	{8'd137,8'd2} : s = 139;
	{8'd137,8'd3} : s = 140;
	{8'd137,8'd4} : s = 141;
	{8'd137,8'd5} : s = 142;
	{8'd137,8'd6} : s = 143;
	{8'd137,8'd7} : s = 144;
	{8'd137,8'd8} : s = 145;
	{8'd137,8'd9} : s = 146;
	{8'd137,8'd10} : s = 147;
	{8'd137,8'd11} : s = 148;
	{8'd137,8'd12} : s = 149;
	{8'd137,8'd13} : s = 150;
	{8'd137,8'd14} : s = 151;
	{8'd137,8'd15} : s = 152;
	{8'd137,8'd16} : s = 153;
	{8'd137,8'd17} : s = 154;
	{8'd137,8'd18} : s = 155;
	{8'd137,8'd19} : s = 156;
	{8'd137,8'd20} : s = 157;
	{8'd137,8'd21} : s = 158;
	{8'd137,8'd22} : s = 159;
	{8'd137,8'd23} : s = 160;
	{8'd137,8'd24} : s = 161;
	{8'd137,8'd25} : s = 162;
	{8'd137,8'd26} : s = 163;
	{8'd137,8'd27} : s = 164;
	{8'd137,8'd28} : s = 165;
	{8'd137,8'd29} : s = 166;
	{8'd137,8'd30} : s = 167;
	{8'd137,8'd31} : s = 168;
	{8'd137,8'd32} : s = 169;
	{8'd137,8'd33} : s = 170;
	{8'd137,8'd34} : s = 171;
	{8'd137,8'd35} : s = 172;
	{8'd137,8'd36} : s = 173;
	{8'd137,8'd37} : s = 174;
	{8'd137,8'd38} : s = 175;
	{8'd137,8'd39} : s = 176;
	{8'd137,8'd40} : s = 177;
	{8'd137,8'd41} : s = 178;
	{8'd137,8'd42} : s = 179;
	{8'd137,8'd43} : s = 180;
	{8'd137,8'd44} : s = 181;
	{8'd137,8'd45} : s = 182;
	{8'd137,8'd46} : s = 183;
	{8'd137,8'd47} : s = 184;
	{8'd137,8'd48} : s = 185;
	{8'd137,8'd49} : s = 186;
	{8'd137,8'd50} : s = 187;
	{8'd137,8'd51} : s = 188;
	{8'd137,8'd52} : s = 189;
	{8'd137,8'd53} : s = 190;
	{8'd137,8'd54} : s = 191;
	{8'd137,8'd55} : s = 192;
	{8'd137,8'd56} : s = 193;
	{8'd137,8'd57} : s = 194;
	{8'd137,8'd58} : s = 195;
	{8'd137,8'd59} : s = 196;
	{8'd137,8'd60} : s = 197;
	{8'd137,8'd61} : s = 198;
	{8'd137,8'd62} : s = 199;
	{8'd137,8'd63} : s = 200;
	{8'd137,8'd64} : s = 201;
	{8'd137,8'd65} : s = 202;
	{8'd137,8'd66} : s = 203;
	{8'd137,8'd67} : s = 204;
	{8'd137,8'd68} : s = 205;
	{8'd137,8'd69} : s = 206;
	{8'd137,8'd70} : s = 207;
	{8'd137,8'd71} : s = 208;
	{8'd137,8'd72} : s = 209;
	{8'd137,8'd73} : s = 210;
	{8'd137,8'd74} : s = 211;
	{8'd137,8'd75} : s = 212;
	{8'd137,8'd76} : s = 213;
	{8'd137,8'd77} : s = 214;
	{8'd137,8'd78} : s = 215;
	{8'd137,8'd79} : s = 216;
	{8'd137,8'd80} : s = 217;
	{8'd137,8'd81} : s = 218;
	{8'd137,8'd82} : s = 219;
	{8'd137,8'd83} : s = 220;
	{8'd137,8'd84} : s = 221;
	{8'd137,8'd85} : s = 222;
	{8'd137,8'd86} : s = 223;
	{8'd137,8'd87} : s = 224;
	{8'd137,8'd88} : s = 225;
	{8'd137,8'd89} : s = 226;
	{8'd137,8'd90} : s = 227;
	{8'd137,8'd91} : s = 228;
	{8'd137,8'd92} : s = 229;
	{8'd137,8'd93} : s = 230;
	{8'd137,8'd94} : s = 231;
	{8'd137,8'd95} : s = 232;
	{8'd137,8'd96} : s = 233;
	{8'd137,8'd97} : s = 234;
	{8'd137,8'd98} : s = 235;
	{8'd137,8'd99} : s = 236;
	{8'd137,8'd100} : s = 237;
	{8'd137,8'd101} : s = 238;
	{8'd137,8'd102} : s = 239;
	{8'd137,8'd103} : s = 240;
	{8'd137,8'd104} : s = 241;
	{8'd137,8'd105} : s = 242;
	{8'd137,8'd106} : s = 243;
	{8'd137,8'd107} : s = 244;
	{8'd137,8'd108} : s = 245;
	{8'd137,8'd109} : s = 246;
	{8'd137,8'd110} : s = 247;
	{8'd137,8'd111} : s = 248;
	{8'd137,8'd112} : s = 249;
	{8'd137,8'd113} : s = 250;
	{8'd137,8'd114} : s = 251;
	{8'd137,8'd115} : s = 252;
	{8'd137,8'd116} : s = 253;
	{8'd137,8'd117} : s = 254;
	{8'd137,8'd118} : s = 255;
	{8'd137,8'd119} : s = 256;
	{8'd137,8'd120} : s = 257;
	{8'd137,8'd121} : s = 258;
	{8'd137,8'd122} : s = 259;
	{8'd137,8'd123} : s = 260;
	{8'd137,8'd124} : s = 261;
	{8'd137,8'd125} : s = 262;
	{8'd137,8'd126} : s = 263;
	{8'd137,8'd127} : s = 264;
	{8'd137,8'd128} : s = 265;
	{8'd137,8'd129} : s = 266;
	{8'd137,8'd130} : s = 267;
	{8'd137,8'd131} : s = 268;
	{8'd137,8'd132} : s = 269;
	{8'd137,8'd133} : s = 270;
	{8'd137,8'd134} : s = 271;
	{8'd137,8'd135} : s = 272;
	{8'd137,8'd136} : s = 273;
	{8'd137,8'd137} : s = 274;
	{8'd137,8'd138} : s = 275;
	{8'd137,8'd139} : s = 276;
	{8'd137,8'd140} : s = 277;
	{8'd137,8'd141} : s = 278;
	{8'd137,8'd142} : s = 279;
	{8'd137,8'd143} : s = 280;
	{8'd137,8'd144} : s = 281;
	{8'd137,8'd145} : s = 282;
	{8'd137,8'd146} : s = 283;
	{8'd137,8'd147} : s = 284;
	{8'd137,8'd148} : s = 285;
	{8'd137,8'd149} : s = 286;
	{8'd137,8'd150} : s = 287;
	{8'd137,8'd151} : s = 288;
	{8'd137,8'd152} : s = 289;
	{8'd137,8'd153} : s = 290;
	{8'd137,8'd154} : s = 291;
	{8'd137,8'd155} : s = 292;
	{8'd137,8'd156} : s = 293;
	{8'd137,8'd157} : s = 294;
	{8'd137,8'd158} : s = 295;
	{8'd137,8'd159} : s = 296;
	{8'd137,8'd160} : s = 297;
	{8'd137,8'd161} : s = 298;
	{8'd137,8'd162} : s = 299;
	{8'd137,8'd163} : s = 300;
	{8'd137,8'd164} : s = 301;
	{8'd137,8'd165} : s = 302;
	{8'd137,8'd166} : s = 303;
	{8'd137,8'd167} : s = 304;
	{8'd137,8'd168} : s = 305;
	{8'd137,8'd169} : s = 306;
	{8'd137,8'd170} : s = 307;
	{8'd137,8'd171} : s = 308;
	{8'd137,8'd172} : s = 309;
	{8'd137,8'd173} : s = 310;
	{8'd137,8'd174} : s = 311;
	{8'd137,8'd175} : s = 312;
	{8'd137,8'd176} : s = 313;
	{8'd137,8'd177} : s = 314;
	{8'd137,8'd178} : s = 315;
	{8'd137,8'd179} : s = 316;
	{8'd137,8'd180} : s = 317;
	{8'd137,8'd181} : s = 318;
	{8'd137,8'd182} : s = 319;
	{8'd137,8'd183} : s = 320;
	{8'd137,8'd184} : s = 321;
	{8'd137,8'd185} : s = 322;
	{8'd137,8'd186} : s = 323;
	{8'd137,8'd187} : s = 324;
	{8'd137,8'd188} : s = 325;
	{8'd137,8'd189} : s = 326;
	{8'd137,8'd190} : s = 327;
	{8'd137,8'd191} : s = 328;
	{8'd137,8'd192} : s = 329;
	{8'd137,8'd193} : s = 330;
	{8'd137,8'd194} : s = 331;
	{8'd137,8'd195} : s = 332;
	{8'd137,8'd196} : s = 333;
	{8'd137,8'd197} : s = 334;
	{8'd137,8'd198} : s = 335;
	{8'd137,8'd199} : s = 336;
	{8'd137,8'd200} : s = 337;
	{8'd137,8'd201} : s = 338;
	{8'd137,8'd202} : s = 339;
	{8'd137,8'd203} : s = 340;
	{8'd137,8'd204} : s = 341;
	{8'd137,8'd205} : s = 342;
	{8'd137,8'd206} : s = 343;
	{8'd137,8'd207} : s = 344;
	{8'd137,8'd208} : s = 345;
	{8'd137,8'd209} : s = 346;
	{8'd137,8'd210} : s = 347;
	{8'd137,8'd211} : s = 348;
	{8'd137,8'd212} : s = 349;
	{8'd137,8'd213} : s = 350;
	{8'd137,8'd214} : s = 351;
	{8'd137,8'd215} : s = 352;
	{8'd137,8'd216} : s = 353;
	{8'd137,8'd217} : s = 354;
	{8'd137,8'd218} : s = 355;
	{8'd137,8'd219} : s = 356;
	{8'd137,8'd220} : s = 357;
	{8'd137,8'd221} : s = 358;
	{8'd137,8'd222} : s = 359;
	{8'd137,8'd223} : s = 360;
	{8'd137,8'd224} : s = 361;
	{8'd137,8'd225} : s = 362;
	{8'd137,8'd226} : s = 363;
	{8'd137,8'd227} : s = 364;
	{8'd137,8'd228} : s = 365;
	{8'd137,8'd229} : s = 366;
	{8'd137,8'd230} : s = 367;
	{8'd137,8'd231} : s = 368;
	{8'd137,8'd232} : s = 369;
	{8'd137,8'd233} : s = 370;
	{8'd137,8'd234} : s = 371;
	{8'd137,8'd235} : s = 372;
	{8'd137,8'd236} : s = 373;
	{8'd137,8'd237} : s = 374;
	{8'd137,8'd238} : s = 375;
	{8'd137,8'd239} : s = 376;
	{8'd137,8'd240} : s = 377;
	{8'd137,8'd241} : s = 378;
	{8'd137,8'd242} : s = 379;
	{8'd137,8'd243} : s = 380;
	{8'd137,8'd244} : s = 381;
	{8'd137,8'd245} : s = 382;
	{8'd137,8'd246} : s = 383;
	{8'd137,8'd247} : s = 384;
	{8'd137,8'd248} : s = 385;
	{8'd137,8'd249} : s = 386;
	{8'd137,8'd250} : s = 387;
	{8'd137,8'd251} : s = 388;
	{8'd137,8'd252} : s = 389;
	{8'd137,8'd253} : s = 390;
	{8'd137,8'd254} : s = 391;
	{8'd137,8'd255} : s = 392;
	{8'd138,8'd0} : s = 138;
	{8'd138,8'd1} : s = 139;
	{8'd138,8'd2} : s = 140;
	{8'd138,8'd3} : s = 141;
	{8'd138,8'd4} : s = 142;
	{8'd138,8'd5} : s = 143;
	{8'd138,8'd6} : s = 144;
	{8'd138,8'd7} : s = 145;
	{8'd138,8'd8} : s = 146;
	{8'd138,8'd9} : s = 147;
	{8'd138,8'd10} : s = 148;
	{8'd138,8'd11} : s = 149;
	{8'd138,8'd12} : s = 150;
	{8'd138,8'd13} : s = 151;
	{8'd138,8'd14} : s = 152;
	{8'd138,8'd15} : s = 153;
	{8'd138,8'd16} : s = 154;
	{8'd138,8'd17} : s = 155;
	{8'd138,8'd18} : s = 156;
	{8'd138,8'd19} : s = 157;
	{8'd138,8'd20} : s = 158;
	{8'd138,8'd21} : s = 159;
	{8'd138,8'd22} : s = 160;
	{8'd138,8'd23} : s = 161;
	{8'd138,8'd24} : s = 162;
	{8'd138,8'd25} : s = 163;
	{8'd138,8'd26} : s = 164;
	{8'd138,8'd27} : s = 165;
	{8'd138,8'd28} : s = 166;
	{8'd138,8'd29} : s = 167;
	{8'd138,8'd30} : s = 168;
	{8'd138,8'd31} : s = 169;
	{8'd138,8'd32} : s = 170;
	{8'd138,8'd33} : s = 171;
	{8'd138,8'd34} : s = 172;
	{8'd138,8'd35} : s = 173;
	{8'd138,8'd36} : s = 174;
	{8'd138,8'd37} : s = 175;
	{8'd138,8'd38} : s = 176;
	{8'd138,8'd39} : s = 177;
	{8'd138,8'd40} : s = 178;
	{8'd138,8'd41} : s = 179;
	{8'd138,8'd42} : s = 180;
	{8'd138,8'd43} : s = 181;
	{8'd138,8'd44} : s = 182;
	{8'd138,8'd45} : s = 183;
	{8'd138,8'd46} : s = 184;
	{8'd138,8'd47} : s = 185;
	{8'd138,8'd48} : s = 186;
	{8'd138,8'd49} : s = 187;
	{8'd138,8'd50} : s = 188;
	{8'd138,8'd51} : s = 189;
	{8'd138,8'd52} : s = 190;
	{8'd138,8'd53} : s = 191;
	{8'd138,8'd54} : s = 192;
	{8'd138,8'd55} : s = 193;
	{8'd138,8'd56} : s = 194;
	{8'd138,8'd57} : s = 195;
	{8'd138,8'd58} : s = 196;
	{8'd138,8'd59} : s = 197;
	{8'd138,8'd60} : s = 198;
	{8'd138,8'd61} : s = 199;
	{8'd138,8'd62} : s = 200;
	{8'd138,8'd63} : s = 201;
	{8'd138,8'd64} : s = 202;
	{8'd138,8'd65} : s = 203;
	{8'd138,8'd66} : s = 204;
	{8'd138,8'd67} : s = 205;
	{8'd138,8'd68} : s = 206;
	{8'd138,8'd69} : s = 207;
	{8'd138,8'd70} : s = 208;
	{8'd138,8'd71} : s = 209;
	{8'd138,8'd72} : s = 210;
	{8'd138,8'd73} : s = 211;
	{8'd138,8'd74} : s = 212;
	{8'd138,8'd75} : s = 213;
	{8'd138,8'd76} : s = 214;
	{8'd138,8'd77} : s = 215;
	{8'd138,8'd78} : s = 216;
	{8'd138,8'd79} : s = 217;
	{8'd138,8'd80} : s = 218;
	{8'd138,8'd81} : s = 219;
	{8'd138,8'd82} : s = 220;
	{8'd138,8'd83} : s = 221;
	{8'd138,8'd84} : s = 222;
	{8'd138,8'd85} : s = 223;
	{8'd138,8'd86} : s = 224;
	{8'd138,8'd87} : s = 225;
	{8'd138,8'd88} : s = 226;
	{8'd138,8'd89} : s = 227;
	{8'd138,8'd90} : s = 228;
	{8'd138,8'd91} : s = 229;
	{8'd138,8'd92} : s = 230;
	{8'd138,8'd93} : s = 231;
	{8'd138,8'd94} : s = 232;
	{8'd138,8'd95} : s = 233;
	{8'd138,8'd96} : s = 234;
	{8'd138,8'd97} : s = 235;
	{8'd138,8'd98} : s = 236;
	{8'd138,8'd99} : s = 237;
	{8'd138,8'd100} : s = 238;
	{8'd138,8'd101} : s = 239;
	{8'd138,8'd102} : s = 240;
	{8'd138,8'd103} : s = 241;
	{8'd138,8'd104} : s = 242;
	{8'd138,8'd105} : s = 243;
	{8'd138,8'd106} : s = 244;
	{8'd138,8'd107} : s = 245;
	{8'd138,8'd108} : s = 246;
	{8'd138,8'd109} : s = 247;
	{8'd138,8'd110} : s = 248;
	{8'd138,8'd111} : s = 249;
	{8'd138,8'd112} : s = 250;
	{8'd138,8'd113} : s = 251;
	{8'd138,8'd114} : s = 252;
	{8'd138,8'd115} : s = 253;
	{8'd138,8'd116} : s = 254;
	{8'd138,8'd117} : s = 255;
	{8'd138,8'd118} : s = 256;
	{8'd138,8'd119} : s = 257;
	{8'd138,8'd120} : s = 258;
	{8'd138,8'd121} : s = 259;
	{8'd138,8'd122} : s = 260;
	{8'd138,8'd123} : s = 261;
	{8'd138,8'd124} : s = 262;
	{8'd138,8'd125} : s = 263;
	{8'd138,8'd126} : s = 264;
	{8'd138,8'd127} : s = 265;
	{8'd138,8'd128} : s = 266;
	{8'd138,8'd129} : s = 267;
	{8'd138,8'd130} : s = 268;
	{8'd138,8'd131} : s = 269;
	{8'd138,8'd132} : s = 270;
	{8'd138,8'd133} : s = 271;
	{8'd138,8'd134} : s = 272;
	{8'd138,8'd135} : s = 273;
	{8'd138,8'd136} : s = 274;
	{8'd138,8'd137} : s = 275;
	{8'd138,8'd138} : s = 276;
	{8'd138,8'd139} : s = 277;
	{8'd138,8'd140} : s = 278;
	{8'd138,8'd141} : s = 279;
	{8'd138,8'd142} : s = 280;
	{8'd138,8'd143} : s = 281;
	{8'd138,8'd144} : s = 282;
	{8'd138,8'd145} : s = 283;
	{8'd138,8'd146} : s = 284;
	{8'd138,8'd147} : s = 285;
	{8'd138,8'd148} : s = 286;
	{8'd138,8'd149} : s = 287;
	{8'd138,8'd150} : s = 288;
	{8'd138,8'd151} : s = 289;
	{8'd138,8'd152} : s = 290;
	{8'd138,8'd153} : s = 291;
	{8'd138,8'd154} : s = 292;
	{8'd138,8'd155} : s = 293;
	{8'd138,8'd156} : s = 294;
	{8'd138,8'd157} : s = 295;
	{8'd138,8'd158} : s = 296;
	{8'd138,8'd159} : s = 297;
	{8'd138,8'd160} : s = 298;
	{8'd138,8'd161} : s = 299;
	{8'd138,8'd162} : s = 300;
	{8'd138,8'd163} : s = 301;
	{8'd138,8'd164} : s = 302;
	{8'd138,8'd165} : s = 303;
	{8'd138,8'd166} : s = 304;
	{8'd138,8'd167} : s = 305;
	{8'd138,8'd168} : s = 306;
	{8'd138,8'd169} : s = 307;
	{8'd138,8'd170} : s = 308;
	{8'd138,8'd171} : s = 309;
	{8'd138,8'd172} : s = 310;
	{8'd138,8'd173} : s = 311;
	{8'd138,8'd174} : s = 312;
	{8'd138,8'd175} : s = 313;
	{8'd138,8'd176} : s = 314;
	{8'd138,8'd177} : s = 315;
	{8'd138,8'd178} : s = 316;
	{8'd138,8'd179} : s = 317;
	{8'd138,8'd180} : s = 318;
	{8'd138,8'd181} : s = 319;
	{8'd138,8'd182} : s = 320;
	{8'd138,8'd183} : s = 321;
	{8'd138,8'd184} : s = 322;
	{8'd138,8'd185} : s = 323;
	{8'd138,8'd186} : s = 324;
	{8'd138,8'd187} : s = 325;
	{8'd138,8'd188} : s = 326;
	{8'd138,8'd189} : s = 327;
	{8'd138,8'd190} : s = 328;
	{8'd138,8'd191} : s = 329;
	{8'd138,8'd192} : s = 330;
	{8'd138,8'd193} : s = 331;
	{8'd138,8'd194} : s = 332;
	{8'd138,8'd195} : s = 333;
	{8'd138,8'd196} : s = 334;
	{8'd138,8'd197} : s = 335;
	{8'd138,8'd198} : s = 336;
	{8'd138,8'd199} : s = 337;
	{8'd138,8'd200} : s = 338;
	{8'd138,8'd201} : s = 339;
	{8'd138,8'd202} : s = 340;
	{8'd138,8'd203} : s = 341;
	{8'd138,8'd204} : s = 342;
	{8'd138,8'd205} : s = 343;
	{8'd138,8'd206} : s = 344;
	{8'd138,8'd207} : s = 345;
	{8'd138,8'd208} : s = 346;
	{8'd138,8'd209} : s = 347;
	{8'd138,8'd210} : s = 348;
	{8'd138,8'd211} : s = 349;
	{8'd138,8'd212} : s = 350;
	{8'd138,8'd213} : s = 351;
	{8'd138,8'd214} : s = 352;
	{8'd138,8'd215} : s = 353;
	{8'd138,8'd216} : s = 354;
	{8'd138,8'd217} : s = 355;
	{8'd138,8'd218} : s = 356;
	{8'd138,8'd219} : s = 357;
	{8'd138,8'd220} : s = 358;
	{8'd138,8'd221} : s = 359;
	{8'd138,8'd222} : s = 360;
	{8'd138,8'd223} : s = 361;
	{8'd138,8'd224} : s = 362;
	{8'd138,8'd225} : s = 363;
	{8'd138,8'd226} : s = 364;
	{8'd138,8'd227} : s = 365;
	{8'd138,8'd228} : s = 366;
	{8'd138,8'd229} : s = 367;
	{8'd138,8'd230} : s = 368;
	{8'd138,8'd231} : s = 369;
	{8'd138,8'd232} : s = 370;
	{8'd138,8'd233} : s = 371;
	{8'd138,8'd234} : s = 372;
	{8'd138,8'd235} : s = 373;
	{8'd138,8'd236} : s = 374;
	{8'd138,8'd237} : s = 375;
	{8'd138,8'd238} : s = 376;
	{8'd138,8'd239} : s = 377;
	{8'd138,8'd240} : s = 378;
	{8'd138,8'd241} : s = 379;
	{8'd138,8'd242} : s = 380;
	{8'd138,8'd243} : s = 381;
	{8'd138,8'd244} : s = 382;
	{8'd138,8'd245} : s = 383;
	{8'd138,8'd246} : s = 384;
	{8'd138,8'd247} : s = 385;
	{8'd138,8'd248} : s = 386;
	{8'd138,8'd249} : s = 387;
	{8'd138,8'd250} : s = 388;
	{8'd138,8'd251} : s = 389;
	{8'd138,8'd252} : s = 390;
	{8'd138,8'd253} : s = 391;
	{8'd138,8'd254} : s = 392;
	{8'd138,8'd255} : s = 393;
	{8'd139,8'd0} : s = 139;
	{8'd139,8'd1} : s = 140;
	{8'd139,8'd2} : s = 141;
	{8'd139,8'd3} : s = 142;
	{8'd139,8'd4} : s = 143;
	{8'd139,8'd5} : s = 144;
	{8'd139,8'd6} : s = 145;
	{8'd139,8'd7} : s = 146;
	{8'd139,8'd8} : s = 147;
	{8'd139,8'd9} : s = 148;
	{8'd139,8'd10} : s = 149;
	{8'd139,8'd11} : s = 150;
	{8'd139,8'd12} : s = 151;
	{8'd139,8'd13} : s = 152;
	{8'd139,8'd14} : s = 153;
	{8'd139,8'd15} : s = 154;
	{8'd139,8'd16} : s = 155;
	{8'd139,8'd17} : s = 156;
	{8'd139,8'd18} : s = 157;
	{8'd139,8'd19} : s = 158;
	{8'd139,8'd20} : s = 159;
	{8'd139,8'd21} : s = 160;
	{8'd139,8'd22} : s = 161;
	{8'd139,8'd23} : s = 162;
	{8'd139,8'd24} : s = 163;
	{8'd139,8'd25} : s = 164;
	{8'd139,8'd26} : s = 165;
	{8'd139,8'd27} : s = 166;
	{8'd139,8'd28} : s = 167;
	{8'd139,8'd29} : s = 168;
	{8'd139,8'd30} : s = 169;
	{8'd139,8'd31} : s = 170;
	{8'd139,8'd32} : s = 171;
	{8'd139,8'd33} : s = 172;
	{8'd139,8'd34} : s = 173;
	{8'd139,8'd35} : s = 174;
	{8'd139,8'd36} : s = 175;
	{8'd139,8'd37} : s = 176;
	{8'd139,8'd38} : s = 177;
	{8'd139,8'd39} : s = 178;
	{8'd139,8'd40} : s = 179;
	{8'd139,8'd41} : s = 180;
	{8'd139,8'd42} : s = 181;
	{8'd139,8'd43} : s = 182;
	{8'd139,8'd44} : s = 183;
	{8'd139,8'd45} : s = 184;
	{8'd139,8'd46} : s = 185;
	{8'd139,8'd47} : s = 186;
	{8'd139,8'd48} : s = 187;
	{8'd139,8'd49} : s = 188;
	{8'd139,8'd50} : s = 189;
	{8'd139,8'd51} : s = 190;
	{8'd139,8'd52} : s = 191;
	{8'd139,8'd53} : s = 192;
	{8'd139,8'd54} : s = 193;
	{8'd139,8'd55} : s = 194;
	{8'd139,8'd56} : s = 195;
	{8'd139,8'd57} : s = 196;
	{8'd139,8'd58} : s = 197;
	{8'd139,8'd59} : s = 198;
	{8'd139,8'd60} : s = 199;
	{8'd139,8'd61} : s = 200;
	{8'd139,8'd62} : s = 201;
	{8'd139,8'd63} : s = 202;
	{8'd139,8'd64} : s = 203;
	{8'd139,8'd65} : s = 204;
	{8'd139,8'd66} : s = 205;
	{8'd139,8'd67} : s = 206;
	{8'd139,8'd68} : s = 207;
	{8'd139,8'd69} : s = 208;
	{8'd139,8'd70} : s = 209;
	{8'd139,8'd71} : s = 210;
	{8'd139,8'd72} : s = 211;
	{8'd139,8'd73} : s = 212;
	{8'd139,8'd74} : s = 213;
	{8'd139,8'd75} : s = 214;
	{8'd139,8'd76} : s = 215;
	{8'd139,8'd77} : s = 216;
	{8'd139,8'd78} : s = 217;
	{8'd139,8'd79} : s = 218;
	{8'd139,8'd80} : s = 219;
	{8'd139,8'd81} : s = 220;
	{8'd139,8'd82} : s = 221;
	{8'd139,8'd83} : s = 222;
	{8'd139,8'd84} : s = 223;
	{8'd139,8'd85} : s = 224;
	{8'd139,8'd86} : s = 225;
	{8'd139,8'd87} : s = 226;
	{8'd139,8'd88} : s = 227;
	{8'd139,8'd89} : s = 228;
	{8'd139,8'd90} : s = 229;
	{8'd139,8'd91} : s = 230;
	{8'd139,8'd92} : s = 231;
	{8'd139,8'd93} : s = 232;
	{8'd139,8'd94} : s = 233;
	{8'd139,8'd95} : s = 234;
	{8'd139,8'd96} : s = 235;
	{8'd139,8'd97} : s = 236;
	{8'd139,8'd98} : s = 237;
	{8'd139,8'd99} : s = 238;
	{8'd139,8'd100} : s = 239;
	{8'd139,8'd101} : s = 240;
	{8'd139,8'd102} : s = 241;
	{8'd139,8'd103} : s = 242;
	{8'd139,8'd104} : s = 243;
	{8'd139,8'd105} : s = 244;
	{8'd139,8'd106} : s = 245;
	{8'd139,8'd107} : s = 246;
	{8'd139,8'd108} : s = 247;
	{8'd139,8'd109} : s = 248;
	{8'd139,8'd110} : s = 249;
	{8'd139,8'd111} : s = 250;
	{8'd139,8'd112} : s = 251;
	{8'd139,8'd113} : s = 252;
	{8'd139,8'd114} : s = 253;
	{8'd139,8'd115} : s = 254;
	{8'd139,8'd116} : s = 255;
	{8'd139,8'd117} : s = 256;
	{8'd139,8'd118} : s = 257;
	{8'd139,8'd119} : s = 258;
	{8'd139,8'd120} : s = 259;
	{8'd139,8'd121} : s = 260;
	{8'd139,8'd122} : s = 261;
	{8'd139,8'd123} : s = 262;
	{8'd139,8'd124} : s = 263;
	{8'd139,8'd125} : s = 264;
	{8'd139,8'd126} : s = 265;
	{8'd139,8'd127} : s = 266;
	{8'd139,8'd128} : s = 267;
	{8'd139,8'd129} : s = 268;
	{8'd139,8'd130} : s = 269;
	{8'd139,8'd131} : s = 270;
	{8'd139,8'd132} : s = 271;
	{8'd139,8'd133} : s = 272;
	{8'd139,8'd134} : s = 273;
	{8'd139,8'd135} : s = 274;
	{8'd139,8'd136} : s = 275;
	{8'd139,8'd137} : s = 276;
	{8'd139,8'd138} : s = 277;
	{8'd139,8'd139} : s = 278;
	{8'd139,8'd140} : s = 279;
	{8'd139,8'd141} : s = 280;
	{8'd139,8'd142} : s = 281;
	{8'd139,8'd143} : s = 282;
	{8'd139,8'd144} : s = 283;
	{8'd139,8'd145} : s = 284;
	{8'd139,8'd146} : s = 285;
	{8'd139,8'd147} : s = 286;
	{8'd139,8'd148} : s = 287;
	{8'd139,8'd149} : s = 288;
	{8'd139,8'd150} : s = 289;
	{8'd139,8'd151} : s = 290;
	{8'd139,8'd152} : s = 291;
	{8'd139,8'd153} : s = 292;
	{8'd139,8'd154} : s = 293;
	{8'd139,8'd155} : s = 294;
	{8'd139,8'd156} : s = 295;
	{8'd139,8'd157} : s = 296;
	{8'd139,8'd158} : s = 297;
	{8'd139,8'd159} : s = 298;
	{8'd139,8'd160} : s = 299;
	{8'd139,8'd161} : s = 300;
	{8'd139,8'd162} : s = 301;
	{8'd139,8'd163} : s = 302;
	{8'd139,8'd164} : s = 303;
	{8'd139,8'd165} : s = 304;
	{8'd139,8'd166} : s = 305;
	{8'd139,8'd167} : s = 306;
	{8'd139,8'd168} : s = 307;
	{8'd139,8'd169} : s = 308;
	{8'd139,8'd170} : s = 309;
	{8'd139,8'd171} : s = 310;
	{8'd139,8'd172} : s = 311;
	{8'd139,8'd173} : s = 312;
	{8'd139,8'd174} : s = 313;
	{8'd139,8'd175} : s = 314;
	{8'd139,8'd176} : s = 315;
	{8'd139,8'd177} : s = 316;
	{8'd139,8'd178} : s = 317;
	{8'd139,8'd179} : s = 318;
	{8'd139,8'd180} : s = 319;
	{8'd139,8'd181} : s = 320;
	{8'd139,8'd182} : s = 321;
	{8'd139,8'd183} : s = 322;
	{8'd139,8'd184} : s = 323;
	{8'd139,8'd185} : s = 324;
	{8'd139,8'd186} : s = 325;
	{8'd139,8'd187} : s = 326;
	{8'd139,8'd188} : s = 327;
	{8'd139,8'd189} : s = 328;
	{8'd139,8'd190} : s = 329;
	{8'd139,8'd191} : s = 330;
	{8'd139,8'd192} : s = 331;
	{8'd139,8'd193} : s = 332;
	{8'd139,8'd194} : s = 333;
	{8'd139,8'd195} : s = 334;
	{8'd139,8'd196} : s = 335;
	{8'd139,8'd197} : s = 336;
	{8'd139,8'd198} : s = 337;
	{8'd139,8'd199} : s = 338;
	{8'd139,8'd200} : s = 339;
	{8'd139,8'd201} : s = 340;
	{8'd139,8'd202} : s = 341;
	{8'd139,8'd203} : s = 342;
	{8'd139,8'd204} : s = 343;
	{8'd139,8'd205} : s = 344;
	{8'd139,8'd206} : s = 345;
	{8'd139,8'd207} : s = 346;
	{8'd139,8'd208} : s = 347;
	{8'd139,8'd209} : s = 348;
	{8'd139,8'd210} : s = 349;
	{8'd139,8'd211} : s = 350;
	{8'd139,8'd212} : s = 351;
	{8'd139,8'd213} : s = 352;
	{8'd139,8'd214} : s = 353;
	{8'd139,8'd215} : s = 354;
	{8'd139,8'd216} : s = 355;
	{8'd139,8'd217} : s = 356;
	{8'd139,8'd218} : s = 357;
	{8'd139,8'd219} : s = 358;
	{8'd139,8'd220} : s = 359;
	{8'd139,8'd221} : s = 360;
	{8'd139,8'd222} : s = 361;
	{8'd139,8'd223} : s = 362;
	{8'd139,8'd224} : s = 363;
	{8'd139,8'd225} : s = 364;
	{8'd139,8'd226} : s = 365;
	{8'd139,8'd227} : s = 366;
	{8'd139,8'd228} : s = 367;
	{8'd139,8'd229} : s = 368;
	{8'd139,8'd230} : s = 369;
	{8'd139,8'd231} : s = 370;
	{8'd139,8'd232} : s = 371;
	{8'd139,8'd233} : s = 372;
	{8'd139,8'd234} : s = 373;
	{8'd139,8'd235} : s = 374;
	{8'd139,8'd236} : s = 375;
	{8'd139,8'd237} : s = 376;
	{8'd139,8'd238} : s = 377;
	{8'd139,8'd239} : s = 378;
	{8'd139,8'd240} : s = 379;
	{8'd139,8'd241} : s = 380;
	{8'd139,8'd242} : s = 381;
	{8'd139,8'd243} : s = 382;
	{8'd139,8'd244} : s = 383;
	{8'd139,8'd245} : s = 384;
	{8'd139,8'd246} : s = 385;
	{8'd139,8'd247} : s = 386;
	{8'd139,8'd248} : s = 387;
	{8'd139,8'd249} : s = 388;
	{8'd139,8'd250} : s = 389;
	{8'd139,8'd251} : s = 390;
	{8'd139,8'd252} : s = 391;
	{8'd139,8'd253} : s = 392;
	{8'd139,8'd254} : s = 393;
	{8'd139,8'd255} : s = 394;
	{8'd140,8'd0} : s = 140;
	{8'd140,8'd1} : s = 141;
	{8'd140,8'd2} : s = 142;
	{8'd140,8'd3} : s = 143;
	{8'd140,8'd4} : s = 144;
	{8'd140,8'd5} : s = 145;
	{8'd140,8'd6} : s = 146;
	{8'd140,8'd7} : s = 147;
	{8'd140,8'd8} : s = 148;
	{8'd140,8'd9} : s = 149;
	{8'd140,8'd10} : s = 150;
	{8'd140,8'd11} : s = 151;
	{8'd140,8'd12} : s = 152;
	{8'd140,8'd13} : s = 153;
	{8'd140,8'd14} : s = 154;
	{8'd140,8'd15} : s = 155;
	{8'd140,8'd16} : s = 156;
	{8'd140,8'd17} : s = 157;
	{8'd140,8'd18} : s = 158;
	{8'd140,8'd19} : s = 159;
	{8'd140,8'd20} : s = 160;
	{8'd140,8'd21} : s = 161;
	{8'd140,8'd22} : s = 162;
	{8'd140,8'd23} : s = 163;
	{8'd140,8'd24} : s = 164;
	{8'd140,8'd25} : s = 165;
	{8'd140,8'd26} : s = 166;
	{8'd140,8'd27} : s = 167;
	{8'd140,8'd28} : s = 168;
	{8'd140,8'd29} : s = 169;
	{8'd140,8'd30} : s = 170;
	{8'd140,8'd31} : s = 171;
	{8'd140,8'd32} : s = 172;
	{8'd140,8'd33} : s = 173;
	{8'd140,8'd34} : s = 174;
	{8'd140,8'd35} : s = 175;
	{8'd140,8'd36} : s = 176;
	{8'd140,8'd37} : s = 177;
	{8'd140,8'd38} : s = 178;
	{8'd140,8'd39} : s = 179;
	{8'd140,8'd40} : s = 180;
	{8'd140,8'd41} : s = 181;
	{8'd140,8'd42} : s = 182;
	{8'd140,8'd43} : s = 183;
	{8'd140,8'd44} : s = 184;
	{8'd140,8'd45} : s = 185;
	{8'd140,8'd46} : s = 186;
	{8'd140,8'd47} : s = 187;
	{8'd140,8'd48} : s = 188;
	{8'd140,8'd49} : s = 189;
	{8'd140,8'd50} : s = 190;
	{8'd140,8'd51} : s = 191;
	{8'd140,8'd52} : s = 192;
	{8'd140,8'd53} : s = 193;
	{8'd140,8'd54} : s = 194;
	{8'd140,8'd55} : s = 195;
	{8'd140,8'd56} : s = 196;
	{8'd140,8'd57} : s = 197;
	{8'd140,8'd58} : s = 198;
	{8'd140,8'd59} : s = 199;
	{8'd140,8'd60} : s = 200;
	{8'd140,8'd61} : s = 201;
	{8'd140,8'd62} : s = 202;
	{8'd140,8'd63} : s = 203;
	{8'd140,8'd64} : s = 204;
	{8'd140,8'd65} : s = 205;
	{8'd140,8'd66} : s = 206;
	{8'd140,8'd67} : s = 207;
	{8'd140,8'd68} : s = 208;
	{8'd140,8'd69} : s = 209;
	{8'd140,8'd70} : s = 210;
	{8'd140,8'd71} : s = 211;
	{8'd140,8'd72} : s = 212;
	{8'd140,8'd73} : s = 213;
	{8'd140,8'd74} : s = 214;
	{8'd140,8'd75} : s = 215;
	{8'd140,8'd76} : s = 216;
	{8'd140,8'd77} : s = 217;
	{8'd140,8'd78} : s = 218;
	{8'd140,8'd79} : s = 219;
	{8'd140,8'd80} : s = 220;
	{8'd140,8'd81} : s = 221;
	{8'd140,8'd82} : s = 222;
	{8'd140,8'd83} : s = 223;
	{8'd140,8'd84} : s = 224;
	{8'd140,8'd85} : s = 225;
	{8'd140,8'd86} : s = 226;
	{8'd140,8'd87} : s = 227;
	{8'd140,8'd88} : s = 228;
	{8'd140,8'd89} : s = 229;
	{8'd140,8'd90} : s = 230;
	{8'd140,8'd91} : s = 231;
	{8'd140,8'd92} : s = 232;
	{8'd140,8'd93} : s = 233;
	{8'd140,8'd94} : s = 234;
	{8'd140,8'd95} : s = 235;
	{8'd140,8'd96} : s = 236;
	{8'd140,8'd97} : s = 237;
	{8'd140,8'd98} : s = 238;
	{8'd140,8'd99} : s = 239;
	{8'd140,8'd100} : s = 240;
	{8'd140,8'd101} : s = 241;
	{8'd140,8'd102} : s = 242;
	{8'd140,8'd103} : s = 243;
	{8'd140,8'd104} : s = 244;
	{8'd140,8'd105} : s = 245;
	{8'd140,8'd106} : s = 246;
	{8'd140,8'd107} : s = 247;
	{8'd140,8'd108} : s = 248;
	{8'd140,8'd109} : s = 249;
	{8'd140,8'd110} : s = 250;
	{8'd140,8'd111} : s = 251;
	{8'd140,8'd112} : s = 252;
	{8'd140,8'd113} : s = 253;
	{8'd140,8'd114} : s = 254;
	{8'd140,8'd115} : s = 255;
	{8'd140,8'd116} : s = 256;
	{8'd140,8'd117} : s = 257;
	{8'd140,8'd118} : s = 258;
	{8'd140,8'd119} : s = 259;
	{8'd140,8'd120} : s = 260;
	{8'd140,8'd121} : s = 261;
	{8'd140,8'd122} : s = 262;
	{8'd140,8'd123} : s = 263;
	{8'd140,8'd124} : s = 264;
	{8'd140,8'd125} : s = 265;
	{8'd140,8'd126} : s = 266;
	{8'd140,8'd127} : s = 267;
	{8'd140,8'd128} : s = 268;
	{8'd140,8'd129} : s = 269;
	{8'd140,8'd130} : s = 270;
	{8'd140,8'd131} : s = 271;
	{8'd140,8'd132} : s = 272;
	{8'd140,8'd133} : s = 273;
	{8'd140,8'd134} : s = 274;
	{8'd140,8'd135} : s = 275;
	{8'd140,8'd136} : s = 276;
	{8'd140,8'd137} : s = 277;
	{8'd140,8'd138} : s = 278;
	{8'd140,8'd139} : s = 279;
	{8'd140,8'd140} : s = 280;
	{8'd140,8'd141} : s = 281;
	{8'd140,8'd142} : s = 282;
	{8'd140,8'd143} : s = 283;
	{8'd140,8'd144} : s = 284;
	{8'd140,8'd145} : s = 285;
	{8'd140,8'd146} : s = 286;
	{8'd140,8'd147} : s = 287;
	{8'd140,8'd148} : s = 288;
	{8'd140,8'd149} : s = 289;
	{8'd140,8'd150} : s = 290;
	{8'd140,8'd151} : s = 291;
	{8'd140,8'd152} : s = 292;
	{8'd140,8'd153} : s = 293;
	{8'd140,8'd154} : s = 294;
	{8'd140,8'd155} : s = 295;
	{8'd140,8'd156} : s = 296;
	{8'd140,8'd157} : s = 297;
	{8'd140,8'd158} : s = 298;
	{8'd140,8'd159} : s = 299;
	{8'd140,8'd160} : s = 300;
	{8'd140,8'd161} : s = 301;
	{8'd140,8'd162} : s = 302;
	{8'd140,8'd163} : s = 303;
	{8'd140,8'd164} : s = 304;
	{8'd140,8'd165} : s = 305;
	{8'd140,8'd166} : s = 306;
	{8'd140,8'd167} : s = 307;
	{8'd140,8'd168} : s = 308;
	{8'd140,8'd169} : s = 309;
	{8'd140,8'd170} : s = 310;
	{8'd140,8'd171} : s = 311;
	{8'd140,8'd172} : s = 312;
	{8'd140,8'd173} : s = 313;
	{8'd140,8'd174} : s = 314;
	{8'd140,8'd175} : s = 315;
	{8'd140,8'd176} : s = 316;
	{8'd140,8'd177} : s = 317;
	{8'd140,8'd178} : s = 318;
	{8'd140,8'd179} : s = 319;
	{8'd140,8'd180} : s = 320;
	{8'd140,8'd181} : s = 321;
	{8'd140,8'd182} : s = 322;
	{8'd140,8'd183} : s = 323;
	{8'd140,8'd184} : s = 324;
	{8'd140,8'd185} : s = 325;
	{8'd140,8'd186} : s = 326;
	{8'd140,8'd187} : s = 327;
	{8'd140,8'd188} : s = 328;
	{8'd140,8'd189} : s = 329;
	{8'd140,8'd190} : s = 330;
	{8'd140,8'd191} : s = 331;
	{8'd140,8'd192} : s = 332;
	{8'd140,8'd193} : s = 333;
	{8'd140,8'd194} : s = 334;
	{8'd140,8'd195} : s = 335;
	{8'd140,8'd196} : s = 336;
	{8'd140,8'd197} : s = 337;
	{8'd140,8'd198} : s = 338;
	{8'd140,8'd199} : s = 339;
	{8'd140,8'd200} : s = 340;
	{8'd140,8'd201} : s = 341;
	{8'd140,8'd202} : s = 342;
	{8'd140,8'd203} : s = 343;
	{8'd140,8'd204} : s = 344;
	{8'd140,8'd205} : s = 345;
	{8'd140,8'd206} : s = 346;
	{8'd140,8'd207} : s = 347;
	{8'd140,8'd208} : s = 348;
	{8'd140,8'd209} : s = 349;
	{8'd140,8'd210} : s = 350;
	{8'd140,8'd211} : s = 351;
	{8'd140,8'd212} : s = 352;
	{8'd140,8'd213} : s = 353;
	{8'd140,8'd214} : s = 354;
	{8'd140,8'd215} : s = 355;
	{8'd140,8'd216} : s = 356;
	{8'd140,8'd217} : s = 357;
	{8'd140,8'd218} : s = 358;
	{8'd140,8'd219} : s = 359;
	{8'd140,8'd220} : s = 360;
	{8'd140,8'd221} : s = 361;
	{8'd140,8'd222} : s = 362;
	{8'd140,8'd223} : s = 363;
	{8'd140,8'd224} : s = 364;
	{8'd140,8'd225} : s = 365;
	{8'd140,8'd226} : s = 366;
	{8'd140,8'd227} : s = 367;
	{8'd140,8'd228} : s = 368;
	{8'd140,8'd229} : s = 369;
	{8'd140,8'd230} : s = 370;
	{8'd140,8'd231} : s = 371;
	{8'd140,8'd232} : s = 372;
	{8'd140,8'd233} : s = 373;
	{8'd140,8'd234} : s = 374;
	{8'd140,8'd235} : s = 375;
	{8'd140,8'd236} : s = 376;
	{8'd140,8'd237} : s = 377;
	{8'd140,8'd238} : s = 378;
	{8'd140,8'd239} : s = 379;
	{8'd140,8'd240} : s = 380;
	{8'd140,8'd241} : s = 381;
	{8'd140,8'd242} : s = 382;
	{8'd140,8'd243} : s = 383;
	{8'd140,8'd244} : s = 384;
	{8'd140,8'd245} : s = 385;
	{8'd140,8'd246} : s = 386;
	{8'd140,8'd247} : s = 387;
	{8'd140,8'd248} : s = 388;
	{8'd140,8'd249} : s = 389;
	{8'd140,8'd250} : s = 390;
	{8'd140,8'd251} : s = 391;
	{8'd140,8'd252} : s = 392;
	{8'd140,8'd253} : s = 393;
	{8'd140,8'd254} : s = 394;
	{8'd140,8'd255} : s = 395;
	{8'd141,8'd0} : s = 141;
	{8'd141,8'd1} : s = 142;
	{8'd141,8'd2} : s = 143;
	{8'd141,8'd3} : s = 144;
	{8'd141,8'd4} : s = 145;
	{8'd141,8'd5} : s = 146;
	{8'd141,8'd6} : s = 147;
	{8'd141,8'd7} : s = 148;
	{8'd141,8'd8} : s = 149;
	{8'd141,8'd9} : s = 150;
	{8'd141,8'd10} : s = 151;
	{8'd141,8'd11} : s = 152;
	{8'd141,8'd12} : s = 153;
	{8'd141,8'd13} : s = 154;
	{8'd141,8'd14} : s = 155;
	{8'd141,8'd15} : s = 156;
	{8'd141,8'd16} : s = 157;
	{8'd141,8'd17} : s = 158;
	{8'd141,8'd18} : s = 159;
	{8'd141,8'd19} : s = 160;
	{8'd141,8'd20} : s = 161;
	{8'd141,8'd21} : s = 162;
	{8'd141,8'd22} : s = 163;
	{8'd141,8'd23} : s = 164;
	{8'd141,8'd24} : s = 165;
	{8'd141,8'd25} : s = 166;
	{8'd141,8'd26} : s = 167;
	{8'd141,8'd27} : s = 168;
	{8'd141,8'd28} : s = 169;
	{8'd141,8'd29} : s = 170;
	{8'd141,8'd30} : s = 171;
	{8'd141,8'd31} : s = 172;
	{8'd141,8'd32} : s = 173;
	{8'd141,8'd33} : s = 174;
	{8'd141,8'd34} : s = 175;
	{8'd141,8'd35} : s = 176;
	{8'd141,8'd36} : s = 177;
	{8'd141,8'd37} : s = 178;
	{8'd141,8'd38} : s = 179;
	{8'd141,8'd39} : s = 180;
	{8'd141,8'd40} : s = 181;
	{8'd141,8'd41} : s = 182;
	{8'd141,8'd42} : s = 183;
	{8'd141,8'd43} : s = 184;
	{8'd141,8'd44} : s = 185;
	{8'd141,8'd45} : s = 186;
	{8'd141,8'd46} : s = 187;
	{8'd141,8'd47} : s = 188;
	{8'd141,8'd48} : s = 189;
	{8'd141,8'd49} : s = 190;
	{8'd141,8'd50} : s = 191;
	{8'd141,8'd51} : s = 192;
	{8'd141,8'd52} : s = 193;
	{8'd141,8'd53} : s = 194;
	{8'd141,8'd54} : s = 195;
	{8'd141,8'd55} : s = 196;
	{8'd141,8'd56} : s = 197;
	{8'd141,8'd57} : s = 198;
	{8'd141,8'd58} : s = 199;
	{8'd141,8'd59} : s = 200;
	{8'd141,8'd60} : s = 201;
	{8'd141,8'd61} : s = 202;
	{8'd141,8'd62} : s = 203;
	{8'd141,8'd63} : s = 204;
	{8'd141,8'd64} : s = 205;
	{8'd141,8'd65} : s = 206;
	{8'd141,8'd66} : s = 207;
	{8'd141,8'd67} : s = 208;
	{8'd141,8'd68} : s = 209;
	{8'd141,8'd69} : s = 210;
	{8'd141,8'd70} : s = 211;
	{8'd141,8'd71} : s = 212;
	{8'd141,8'd72} : s = 213;
	{8'd141,8'd73} : s = 214;
	{8'd141,8'd74} : s = 215;
	{8'd141,8'd75} : s = 216;
	{8'd141,8'd76} : s = 217;
	{8'd141,8'd77} : s = 218;
	{8'd141,8'd78} : s = 219;
	{8'd141,8'd79} : s = 220;
	{8'd141,8'd80} : s = 221;
	{8'd141,8'd81} : s = 222;
	{8'd141,8'd82} : s = 223;
	{8'd141,8'd83} : s = 224;
	{8'd141,8'd84} : s = 225;
	{8'd141,8'd85} : s = 226;
	{8'd141,8'd86} : s = 227;
	{8'd141,8'd87} : s = 228;
	{8'd141,8'd88} : s = 229;
	{8'd141,8'd89} : s = 230;
	{8'd141,8'd90} : s = 231;
	{8'd141,8'd91} : s = 232;
	{8'd141,8'd92} : s = 233;
	{8'd141,8'd93} : s = 234;
	{8'd141,8'd94} : s = 235;
	{8'd141,8'd95} : s = 236;
	{8'd141,8'd96} : s = 237;
	{8'd141,8'd97} : s = 238;
	{8'd141,8'd98} : s = 239;
	{8'd141,8'd99} : s = 240;
	{8'd141,8'd100} : s = 241;
	{8'd141,8'd101} : s = 242;
	{8'd141,8'd102} : s = 243;
	{8'd141,8'd103} : s = 244;
	{8'd141,8'd104} : s = 245;
	{8'd141,8'd105} : s = 246;
	{8'd141,8'd106} : s = 247;
	{8'd141,8'd107} : s = 248;
	{8'd141,8'd108} : s = 249;
	{8'd141,8'd109} : s = 250;
	{8'd141,8'd110} : s = 251;
	{8'd141,8'd111} : s = 252;
	{8'd141,8'd112} : s = 253;
	{8'd141,8'd113} : s = 254;
	{8'd141,8'd114} : s = 255;
	{8'd141,8'd115} : s = 256;
	{8'd141,8'd116} : s = 257;
	{8'd141,8'd117} : s = 258;
	{8'd141,8'd118} : s = 259;
	{8'd141,8'd119} : s = 260;
	{8'd141,8'd120} : s = 261;
	{8'd141,8'd121} : s = 262;
	{8'd141,8'd122} : s = 263;
	{8'd141,8'd123} : s = 264;
	{8'd141,8'd124} : s = 265;
	{8'd141,8'd125} : s = 266;
	{8'd141,8'd126} : s = 267;
	{8'd141,8'd127} : s = 268;
	{8'd141,8'd128} : s = 269;
	{8'd141,8'd129} : s = 270;
	{8'd141,8'd130} : s = 271;
	{8'd141,8'd131} : s = 272;
	{8'd141,8'd132} : s = 273;
	{8'd141,8'd133} : s = 274;
	{8'd141,8'd134} : s = 275;
	{8'd141,8'd135} : s = 276;
	{8'd141,8'd136} : s = 277;
	{8'd141,8'd137} : s = 278;
	{8'd141,8'd138} : s = 279;
	{8'd141,8'd139} : s = 280;
	{8'd141,8'd140} : s = 281;
	{8'd141,8'd141} : s = 282;
	{8'd141,8'd142} : s = 283;
	{8'd141,8'd143} : s = 284;
	{8'd141,8'd144} : s = 285;
	{8'd141,8'd145} : s = 286;
	{8'd141,8'd146} : s = 287;
	{8'd141,8'd147} : s = 288;
	{8'd141,8'd148} : s = 289;
	{8'd141,8'd149} : s = 290;
	{8'd141,8'd150} : s = 291;
	{8'd141,8'd151} : s = 292;
	{8'd141,8'd152} : s = 293;
	{8'd141,8'd153} : s = 294;
	{8'd141,8'd154} : s = 295;
	{8'd141,8'd155} : s = 296;
	{8'd141,8'd156} : s = 297;
	{8'd141,8'd157} : s = 298;
	{8'd141,8'd158} : s = 299;
	{8'd141,8'd159} : s = 300;
	{8'd141,8'd160} : s = 301;
	{8'd141,8'd161} : s = 302;
	{8'd141,8'd162} : s = 303;
	{8'd141,8'd163} : s = 304;
	{8'd141,8'd164} : s = 305;
	{8'd141,8'd165} : s = 306;
	{8'd141,8'd166} : s = 307;
	{8'd141,8'd167} : s = 308;
	{8'd141,8'd168} : s = 309;
	{8'd141,8'd169} : s = 310;
	{8'd141,8'd170} : s = 311;
	{8'd141,8'd171} : s = 312;
	{8'd141,8'd172} : s = 313;
	{8'd141,8'd173} : s = 314;
	{8'd141,8'd174} : s = 315;
	{8'd141,8'd175} : s = 316;
	{8'd141,8'd176} : s = 317;
	{8'd141,8'd177} : s = 318;
	{8'd141,8'd178} : s = 319;
	{8'd141,8'd179} : s = 320;
	{8'd141,8'd180} : s = 321;
	{8'd141,8'd181} : s = 322;
	{8'd141,8'd182} : s = 323;
	{8'd141,8'd183} : s = 324;
	{8'd141,8'd184} : s = 325;
	{8'd141,8'd185} : s = 326;
	{8'd141,8'd186} : s = 327;
	{8'd141,8'd187} : s = 328;
	{8'd141,8'd188} : s = 329;
	{8'd141,8'd189} : s = 330;
	{8'd141,8'd190} : s = 331;
	{8'd141,8'd191} : s = 332;
	{8'd141,8'd192} : s = 333;
	{8'd141,8'd193} : s = 334;
	{8'd141,8'd194} : s = 335;
	{8'd141,8'd195} : s = 336;
	{8'd141,8'd196} : s = 337;
	{8'd141,8'd197} : s = 338;
	{8'd141,8'd198} : s = 339;
	{8'd141,8'd199} : s = 340;
	{8'd141,8'd200} : s = 341;
	{8'd141,8'd201} : s = 342;
	{8'd141,8'd202} : s = 343;
	{8'd141,8'd203} : s = 344;
	{8'd141,8'd204} : s = 345;
	{8'd141,8'd205} : s = 346;
	{8'd141,8'd206} : s = 347;
	{8'd141,8'd207} : s = 348;
	{8'd141,8'd208} : s = 349;
	{8'd141,8'd209} : s = 350;
	{8'd141,8'd210} : s = 351;
	{8'd141,8'd211} : s = 352;
	{8'd141,8'd212} : s = 353;
	{8'd141,8'd213} : s = 354;
	{8'd141,8'd214} : s = 355;
	{8'd141,8'd215} : s = 356;
	{8'd141,8'd216} : s = 357;
	{8'd141,8'd217} : s = 358;
	{8'd141,8'd218} : s = 359;
	{8'd141,8'd219} : s = 360;
	{8'd141,8'd220} : s = 361;
	{8'd141,8'd221} : s = 362;
	{8'd141,8'd222} : s = 363;
	{8'd141,8'd223} : s = 364;
	{8'd141,8'd224} : s = 365;
	{8'd141,8'd225} : s = 366;
	{8'd141,8'd226} : s = 367;
	{8'd141,8'd227} : s = 368;
	{8'd141,8'd228} : s = 369;
	{8'd141,8'd229} : s = 370;
	{8'd141,8'd230} : s = 371;
	{8'd141,8'd231} : s = 372;
	{8'd141,8'd232} : s = 373;
	{8'd141,8'd233} : s = 374;
	{8'd141,8'd234} : s = 375;
	{8'd141,8'd235} : s = 376;
	{8'd141,8'd236} : s = 377;
	{8'd141,8'd237} : s = 378;
	{8'd141,8'd238} : s = 379;
	{8'd141,8'd239} : s = 380;
	{8'd141,8'd240} : s = 381;
	{8'd141,8'd241} : s = 382;
	{8'd141,8'd242} : s = 383;
	{8'd141,8'd243} : s = 384;
	{8'd141,8'd244} : s = 385;
	{8'd141,8'd245} : s = 386;
	{8'd141,8'd246} : s = 387;
	{8'd141,8'd247} : s = 388;
	{8'd141,8'd248} : s = 389;
	{8'd141,8'd249} : s = 390;
	{8'd141,8'd250} : s = 391;
	{8'd141,8'd251} : s = 392;
	{8'd141,8'd252} : s = 393;
	{8'd141,8'd253} : s = 394;
	{8'd141,8'd254} : s = 395;
	{8'd141,8'd255} : s = 396;
	{8'd142,8'd0} : s = 142;
	{8'd142,8'd1} : s = 143;
	{8'd142,8'd2} : s = 144;
	{8'd142,8'd3} : s = 145;
	{8'd142,8'd4} : s = 146;
	{8'd142,8'd5} : s = 147;
	{8'd142,8'd6} : s = 148;
	{8'd142,8'd7} : s = 149;
	{8'd142,8'd8} : s = 150;
	{8'd142,8'd9} : s = 151;
	{8'd142,8'd10} : s = 152;
	{8'd142,8'd11} : s = 153;
	{8'd142,8'd12} : s = 154;
	{8'd142,8'd13} : s = 155;
	{8'd142,8'd14} : s = 156;
	{8'd142,8'd15} : s = 157;
	{8'd142,8'd16} : s = 158;
	{8'd142,8'd17} : s = 159;
	{8'd142,8'd18} : s = 160;
	{8'd142,8'd19} : s = 161;
	{8'd142,8'd20} : s = 162;
	{8'd142,8'd21} : s = 163;
	{8'd142,8'd22} : s = 164;
	{8'd142,8'd23} : s = 165;
	{8'd142,8'd24} : s = 166;
	{8'd142,8'd25} : s = 167;
	{8'd142,8'd26} : s = 168;
	{8'd142,8'd27} : s = 169;
	{8'd142,8'd28} : s = 170;
	{8'd142,8'd29} : s = 171;
	{8'd142,8'd30} : s = 172;
	{8'd142,8'd31} : s = 173;
	{8'd142,8'd32} : s = 174;
	{8'd142,8'd33} : s = 175;
	{8'd142,8'd34} : s = 176;
	{8'd142,8'd35} : s = 177;
	{8'd142,8'd36} : s = 178;
	{8'd142,8'd37} : s = 179;
	{8'd142,8'd38} : s = 180;
	{8'd142,8'd39} : s = 181;
	{8'd142,8'd40} : s = 182;
	{8'd142,8'd41} : s = 183;
	{8'd142,8'd42} : s = 184;
	{8'd142,8'd43} : s = 185;
	{8'd142,8'd44} : s = 186;
	{8'd142,8'd45} : s = 187;
	{8'd142,8'd46} : s = 188;
	{8'd142,8'd47} : s = 189;
	{8'd142,8'd48} : s = 190;
	{8'd142,8'd49} : s = 191;
	{8'd142,8'd50} : s = 192;
	{8'd142,8'd51} : s = 193;
	{8'd142,8'd52} : s = 194;
	{8'd142,8'd53} : s = 195;
	{8'd142,8'd54} : s = 196;
	{8'd142,8'd55} : s = 197;
	{8'd142,8'd56} : s = 198;
	{8'd142,8'd57} : s = 199;
	{8'd142,8'd58} : s = 200;
	{8'd142,8'd59} : s = 201;
	{8'd142,8'd60} : s = 202;
	{8'd142,8'd61} : s = 203;
	{8'd142,8'd62} : s = 204;
	{8'd142,8'd63} : s = 205;
	{8'd142,8'd64} : s = 206;
	{8'd142,8'd65} : s = 207;
	{8'd142,8'd66} : s = 208;
	{8'd142,8'd67} : s = 209;
	{8'd142,8'd68} : s = 210;
	{8'd142,8'd69} : s = 211;
	{8'd142,8'd70} : s = 212;
	{8'd142,8'd71} : s = 213;
	{8'd142,8'd72} : s = 214;
	{8'd142,8'd73} : s = 215;
	{8'd142,8'd74} : s = 216;
	{8'd142,8'd75} : s = 217;
	{8'd142,8'd76} : s = 218;
	{8'd142,8'd77} : s = 219;
	{8'd142,8'd78} : s = 220;
	{8'd142,8'd79} : s = 221;
	{8'd142,8'd80} : s = 222;
	{8'd142,8'd81} : s = 223;
	{8'd142,8'd82} : s = 224;
	{8'd142,8'd83} : s = 225;
	{8'd142,8'd84} : s = 226;
	{8'd142,8'd85} : s = 227;
	{8'd142,8'd86} : s = 228;
	{8'd142,8'd87} : s = 229;
	{8'd142,8'd88} : s = 230;
	{8'd142,8'd89} : s = 231;
	{8'd142,8'd90} : s = 232;
	{8'd142,8'd91} : s = 233;
	{8'd142,8'd92} : s = 234;
	{8'd142,8'd93} : s = 235;
	{8'd142,8'd94} : s = 236;
	{8'd142,8'd95} : s = 237;
	{8'd142,8'd96} : s = 238;
	{8'd142,8'd97} : s = 239;
	{8'd142,8'd98} : s = 240;
	{8'd142,8'd99} : s = 241;
	{8'd142,8'd100} : s = 242;
	{8'd142,8'd101} : s = 243;
	{8'd142,8'd102} : s = 244;
	{8'd142,8'd103} : s = 245;
	{8'd142,8'd104} : s = 246;
	{8'd142,8'd105} : s = 247;
	{8'd142,8'd106} : s = 248;
	{8'd142,8'd107} : s = 249;
	{8'd142,8'd108} : s = 250;
	{8'd142,8'd109} : s = 251;
	{8'd142,8'd110} : s = 252;
	{8'd142,8'd111} : s = 253;
	{8'd142,8'd112} : s = 254;
	{8'd142,8'd113} : s = 255;
	{8'd142,8'd114} : s = 256;
	{8'd142,8'd115} : s = 257;
	{8'd142,8'd116} : s = 258;
	{8'd142,8'd117} : s = 259;
	{8'd142,8'd118} : s = 260;
	{8'd142,8'd119} : s = 261;
	{8'd142,8'd120} : s = 262;
	{8'd142,8'd121} : s = 263;
	{8'd142,8'd122} : s = 264;
	{8'd142,8'd123} : s = 265;
	{8'd142,8'd124} : s = 266;
	{8'd142,8'd125} : s = 267;
	{8'd142,8'd126} : s = 268;
	{8'd142,8'd127} : s = 269;
	{8'd142,8'd128} : s = 270;
	{8'd142,8'd129} : s = 271;
	{8'd142,8'd130} : s = 272;
	{8'd142,8'd131} : s = 273;
	{8'd142,8'd132} : s = 274;
	{8'd142,8'd133} : s = 275;
	{8'd142,8'd134} : s = 276;
	{8'd142,8'd135} : s = 277;
	{8'd142,8'd136} : s = 278;
	{8'd142,8'd137} : s = 279;
	{8'd142,8'd138} : s = 280;
	{8'd142,8'd139} : s = 281;
	{8'd142,8'd140} : s = 282;
	{8'd142,8'd141} : s = 283;
	{8'd142,8'd142} : s = 284;
	{8'd142,8'd143} : s = 285;
	{8'd142,8'd144} : s = 286;
	{8'd142,8'd145} : s = 287;
	{8'd142,8'd146} : s = 288;
	{8'd142,8'd147} : s = 289;
	{8'd142,8'd148} : s = 290;
	{8'd142,8'd149} : s = 291;
	{8'd142,8'd150} : s = 292;
	{8'd142,8'd151} : s = 293;
	{8'd142,8'd152} : s = 294;
	{8'd142,8'd153} : s = 295;
	{8'd142,8'd154} : s = 296;
	{8'd142,8'd155} : s = 297;
	{8'd142,8'd156} : s = 298;
	{8'd142,8'd157} : s = 299;
	{8'd142,8'd158} : s = 300;
	{8'd142,8'd159} : s = 301;
	{8'd142,8'd160} : s = 302;
	{8'd142,8'd161} : s = 303;
	{8'd142,8'd162} : s = 304;
	{8'd142,8'd163} : s = 305;
	{8'd142,8'd164} : s = 306;
	{8'd142,8'd165} : s = 307;
	{8'd142,8'd166} : s = 308;
	{8'd142,8'd167} : s = 309;
	{8'd142,8'd168} : s = 310;
	{8'd142,8'd169} : s = 311;
	{8'd142,8'd170} : s = 312;
	{8'd142,8'd171} : s = 313;
	{8'd142,8'd172} : s = 314;
	{8'd142,8'd173} : s = 315;
	{8'd142,8'd174} : s = 316;
	{8'd142,8'd175} : s = 317;
	{8'd142,8'd176} : s = 318;
	{8'd142,8'd177} : s = 319;
	{8'd142,8'd178} : s = 320;
	{8'd142,8'd179} : s = 321;
	{8'd142,8'd180} : s = 322;
	{8'd142,8'd181} : s = 323;
	{8'd142,8'd182} : s = 324;
	{8'd142,8'd183} : s = 325;
	{8'd142,8'd184} : s = 326;
	{8'd142,8'd185} : s = 327;
	{8'd142,8'd186} : s = 328;
	{8'd142,8'd187} : s = 329;
	{8'd142,8'd188} : s = 330;
	{8'd142,8'd189} : s = 331;
	{8'd142,8'd190} : s = 332;
	{8'd142,8'd191} : s = 333;
	{8'd142,8'd192} : s = 334;
	{8'd142,8'd193} : s = 335;
	{8'd142,8'd194} : s = 336;
	{8'd142,8'd195} : s = 337;
	{8'd142,8'd196} : s = 338;
	{8'd142,8'd197} : s = 339;
	{8'd142,8'd198} : s = 340;
	{8'd142,8'd199} : s = 341;
	{8'd142,8'd200} : s = 342;
	{8'd142,8'd201} : s = 343;
	{8'd142,8'd202} : s = 344;
	{8'd142,8'd203} : s = 345;
	{8'd142,8'd204} : s = 346;
	{8'd142,8'd205} : s = 347;
	{8'd142,8'd206} : s = 348;
	{8'd142,8'd207} : s = 349;
	{8'd142,8'd208} : s = 350;
	{8'd142,8'd209} : s = 351;
	{8'd142,8'd210} : s = 352;
	{8'd142,8'd211} : s = 353;
	{8'd142,8'd212} : s = 354;
	{8'd142,8'd213} : s = 355;
	{8'd142,8'd214} : s = 356;
	{8'd142,8'd215} : s = 357;
	{8'd142,8'd216} : s = 358;
	{8'd142,8'd217} : s = 359;
	{8'd142,8'd218} : s = 360;
	{8'd142,8'd219} : s = 361;
	{8'd142,8'd220} : s = 362;
	{8'd142,8'd221} : s = 363;
	{8'd142,8'd222} : s = 364;
	{8'd142,8'd223} : s = 365;
	{8'd142,8'd224} : s = 366;
	{8'd142,8'd225} : s = 367;
	{8'd142,8'd226} : s = 368;
	{8'd142,8'd227} : s = 369;
	{8'd142,8'd228} : s = 370;
	{8'd142,8'd229} : s = 371;
	{8'd142,8'd230} : s = 372;
	{8'd142,8'd231} : s = 373;
	{8'd142,8'd232} : s = 374;
	{8'd142,8'd233} : s = 375;
	{8'd142,8'd234} : s = 376;
	{8'd142,8'd235} : s = 377;
	{8'd142,8'd236} : s = 378;
	{8'd142,8'd237} : s = 379;
	{8'd142,8'd238} : s = 380;
	{8'd142,8'd239} : s = 381;
	{8'd142,8'd240} : s = 382;
	{8'd142,8'd241} : s = 383;
	{8'd142,8'd242} : s = 384;
	{8'd142,8'd243} : s = 385;
	{8'd142,8'd244} : s = 386;
	{8'd142,8'd245} : s = 387;
	{8'd142,8'd246} : s = 388;
	{8'd142,8'd247} : s = 389;
	{8'd142,8'd248} : s = 390;
	{8'd142,8'd249} : s = 391;
	{8'd142,8'd250} : s = 392;
	{8'd142,8'd251} : s = 393;
	{8'd142,8'd252} : s = 394;
	{8'd142,8'd253} : s = 395;
	{8'd142,8'd254} : s = 396;
	{8'd142,8'd255} : s = 397;
	{8'd143,8'd0} : s = 143;
	{8'd143,8'd1} : s = 144;
	{8'd143,8'd2} : s = 145;
	{8'd143,8'd3} : s = 146;
	{8'd143,8'd4} : s = 147;
	{8'd143,8'd5} : s = 148;
	{8'd143,8'd6} : s = 149;
	{8'd143,8'd7} : s = 150;
	{8'd143,8'd8} : s = 151;
	{8'd143,8'd9} : s = 152;
	{8'd143,8'd10} : s = 153;
	{8'd143,8'd11} : s = 154;
	{8'd143,8'd12} : s = 155;
	{8'd143,8'd13} : s = 156;
	{8'd143,8'd14} : s = 157;
	{8'd143,8'd15} : s = 158;
	{8'd143,8'd16} : s = 159;
	{8'd143,8'd17} : s = 160;
	{8'd143,8'd18} : s = 161;
	{8'd143,8'd19} : s = 162;
	{8'd143,8'd20} : s = 163;
	{8'd143,8'd21} : s = 164;
	{8'd143,8'd22} : s = 165;
	{8'd143,8'd23} : s = 166;
	{8'd143,8'd24} : s = 167;
	{8'd143,8'd25} : s = 168;
	{8'd143,8'd26} : s = 169;
	{8'd143,8'd27} : s = 170;
	{8'd143,8'd28} : s = 171;
	{8'd143,8'd29} : s = 172;
	{8'd143,8'd30} : s = 173;
	{8'd143,8'd31} : s = 174;
	{8'd143,8'd32} : s = 175;
	{8'd143,8'd33} : s = 176;
	{8'd143,8'd34} : s = 177;
	{8'd143,8'd35} : s = 178;
	{8'd143,8'd36} : s = 179;
	{8'd143,8'd37} : s = 180;
	{8'd143,8'd38} : s = 181;
	{8'd143,8'd39} : s = 182;
	{8'd143,8'd40} : s = 183;
	{8'd143,8'd41} : s = 184;
	{8'd143,8'd42} : s = 185;
	{8'd143,8'd43} : s = 186;
	{8'd143,8'd44} : s = 187;
	{8'd143,8'd45} : s = 188;
	{8'd143,8'd46} : s = 189;
	{8'd143,8'd47} : s = 190;
	{8'd143,8'd48} : s = 191;
	{8'd143,8'd49} : s = 192;
	{8'd143,8'd50} : s = 193;
	{8'd143,8'd51} : s = 194;
	{8'd143,8'd52} : s = 195;
	{8'd143,8'd53} : s = 196;
	{8'd143,8'd54} : s = 197;
	{8'd143,8'd55} : s = 198;
	{8'd143,8'd56} : s = 199;
	{8'd143,8'd57} : s = 200;
	{8'd143,8'd58} : s = 201;
	{8'd143,8'd59} : s = 202;
	{8'd143,8'd60} : s = 203;
	{8'd143,8'd61} : s = 204;
	{8'd143,8'd62} : s = 205;
	{8'd143,8'd63} : s = 206;
	{8'd143,8'd64} : s = 207;
	{8'd143,8'd65} : s = 208;
	{8'd143,8'd66} : s = 209;
	{8'd143,8'd67} : s = 210;
	{8'd143,8'd68} : s = 211;
	{8'd143,8'd69} : s = 212;
	{8'd143,8'd70} : s = 213;
	{8'd143,8'd71} : s = 214;
	{8'd143,8'd72} : s = 215;
	{8'd143,8'd73} : s = 216;
	{8'd143,8'd74} : s = 217;
	{8'd143,8'd75} : s = 218;
	{8'd143,8'd76} : s = 219;
	{8'd143,8'd77} : s = 220;
	{8'd143,8'd78} : s = 221;
	{8'd143,8'd79} : s = 222;
	{8'd143,8'd80} : s = 223;
	{8'd143,8'd81} : s = 224;
	{8'd143,8'd82} : s = 225;
	{8'd143,8'd83} : s = 226;
	{8'd143,8'd84} : s = 227;
	{8'd143,8'd85} : s = 228;
	{8'd143,8'd86} : s = 229;
	{8'd143,8'd87} : s = 230;
	{8'd143,8'd88} : s = 231;
	{8'd143,8'd89} : s = 232;
	{8'd143,8'd90} : s = 233;
	{8'd143,8'd91} : s = 234;
	{8'd143,8'd92} : s = 235;
	{8'd143,8'd93} : s = 236;
	{8'd143,8'd94} : s = 237;
	{8'd143,8'd95} : s = 238;
	{8'd143,8'd96} : s = 239;
	{8'd143,8'd97} : s = 240;
	{8'd143,8'd98} : s = 241;
	{8'd143,8'd99} : s = 242;
	{8'd143,8'd100} : s = 243;
	{8'd143,8'd101} : s = 244;
	{8'd143,8'd102} : s = 245;
	{8'd143,8'd103} : s = 246;
	{8'd143,8'd104} : s = 247;
	{8'd143,8'd105} : s = 248;
	{8'd143,8'd106} : s = 249;
	{8'd143,8'd107} : s = 250;
	{8'd143,8'd108} : s = 251;
	{8'd143,8'd109} : s = 252;
	{8'd143,8'd110} : s = 253;
	{8'd143,8'd111} : s = 254;
	{8'd143,8'd112} : s = 255;
	{8'd143,8'd113} : s = 256;
	{8'd143,8'd114} : s = 257;
	{8'd143,8'd115} : s = 258;
	{8'd143,8'd116} : s = 259;
	{8'd143,8'd117} : s = 260;
	{8'd143,8'd118} : s = 261;
	{8'd143,8'd119} : s = 262;
	{8'd143,8'd120} : s = 263;
	{8'd143,8'd121} : s = 264;
	{8'd143,8'd122} : s = 265;
	{8'd143,8'd123} : s = 266;
	{8'd143,8'd124} : s = 267;
	{8'd143,8'd125} : s = 268;
	{8'd143,8'd126} : s = 269;
	{8'd143,8'd127} : s = 270;
	{8'd143,8'd128} : s = 271;
	{8'd143,8'd129} : s = 272;
	{8'd143,8'd130} : s = 273;
	{8'd143,8'd131} : s = 274;
	{8'd143,8'd132} : s = 275;
	{8'd143,8'd133} : s = 276;
	{8'd143,8'd134} : s = 277;
	{8'd143,8'd135} : s = 278;
	{8'd143,8'd136} : s = 279;
	{8'd143,8'd137} : s = 280;
	{8'd143,8'd138} : s = 281;
	{8'd143,8'd139} : s = 282;
	{8'd143,8'd140} : s = 283;
	{8'd143,8'd141} : s = 284;
	{8'd143,8'd142} : s = 285;
	{8'd143,8'd143} : s = 286;
	{8'd143,8'd144} : s = 287;
	{8'd143,8'd145} : s = 288;
	{8'd143,8'd146} : s = 289;
	{8'd143,8'd147} : s = 290;
	{8'd143,8'd148} : s = 291;
	{8'd143,8'd149} : s = 292;
	{8'd143,8'd150} : s = 293;
	{8'd143,8'd151} : s = 294;
	{8'd143,8'd152} : s = 295;
	{8'd143,8'd153} : s = 296;
	{8'd143,8'd154} : s = 297;
	{8'd143,8'd155} : s = 298;
	{8'd143,8'd156} : s = 299;
	{8'd143,8'd157} : s = 300;
	{8'd143,8'd158} : s = 301;
	{8'd143,8'd159} : s = 302;
	{8'd143,8'd160} : s = 303;
	{8'd143,8'd161} : s = 304;
	{8'd143,8'd162} : s = 305;
	{8'd143,8'd163} : s = 306;
	{8'd143,8'd164} : s = 307;
	{8'd143,8'd165} : s = 308;
	{8'd143,8'd166} : s = 309;
	{8'd143,8'd167} : s = 310;
	{8'd143,8'd168} : s = 311;
	{8'd143,8'd169} : s = 312;
	{8'd143,8'd170} : s = 313;
	{8'd143,8'd171} : s = 314;
	{8'd143,8'd172} : s = 315;
	{8'd143,8'd173} : s = 316;
	{8'd143,8'd174} : s = 317;
	{8'd143,8'd175} : s = 318;
	{8'd143,8'd176} : s = 319;
	{8'd143,8'd177} : s = 320;
	{8'd143,8'd178} : s = 321;
	{8'd143,8'd179} : s = 322;
	{8'd143,8'd180} : s = 323;
	{8'd143,8'd181} : s = 324;
	{8'd143,8'd182} : s = 325;
	{8'd143,8'd183} : s = 326;
	{8'd143,8'd184} : s = 327;
	{8'd143,8'd185} : s = 328;
	{8'd143,8'd186} : s = 329;
	{8'd143,8'd187} : s = 330;
	{8'd143,8'd188} : s = 331;
	{8'd143,8'd189} : s = 332;
	{8'd143,8'd190} : s = 333;
	{8'd143,8'd191} : s = 334;
	{8'd143,8'd192} : s = 335;
	{8'd143,8'd193} : s = 336;
	{8'd143,8'd194} : s = 337;
	{8'd143,8'd195} : s = 338;
	{8'd143,8'd196} : s = 339;
	{8'd143,8'd197} : s = 340;
	{8'd143,8'd198} : s = 341;
	{8'd143,8'd199} : s = 342;
	{8'd143,8'd200} : s = 343;
	{8'd143,8'd201} : s = 344;
	{8'd143,8'd202} : s = 345;
	{8'd143,8'd203} : s = 346;
	{8'd143,8'd204} : s = 347;
	{8'd143,8'd205} : s = 348;
	{8'd143,8'd206} : s = 349;
	{8'd143,8'd207} : s = 350;
	{8'd143,8'd208} : s = 351;
	{8'd143,8'd209} : s = 352;
	{8'd143,8'd210} : s = 353;
	{8'd143,8'd211} : s = 354;
	{8'd143,8'd212} : s = 355;
	{8'd143,8'd213} : s = 356;
	{8'd143,8'd214} : s = 357;
	{8'd143,8'd215} : s = 358;
	{8'd143,8'd216} : s = 359;
	{8'd143,8'd217} : s = 360;
	{8'd143,8'd218} : s = 361;
	{8'd143,8'd219} : s = 362;
	{8'd143,8'd220} : s = 363;
	{8'd143,8'd221} : s = 364;
	{8'd143,8'd222} : s = 365;
	{8'd143,8'd223} : s = 366;
	{8'd143,8'd224} : s = 367;
	{8'd143,8'd225} : s = 368;
	{8'd143,8'd226} : s = 369;
	{8'd143,8'd227} : s = 370;
	{8'd143,8'd228} : s = 371;
	{8'd143,8'd229} : s = 372;
	{8'd143,8'd230} : s = 373;
	{8'd143,8'd231} : s = 374;
	{8'd143,8'd232} : s = 375;
	{8'd143,8'd233} : s = 376;
	{8'd143,8'd234} : s = 377;
	{8'd143,8'd235} : s = 378;
	{8'd143,8'd236} : s = 379;
	{8'd143,8'd237} : s = 380;
	{8'd143,8'd238} : s = 381;
	{8'd143,8'd239} : s = 382;
	{8'd143,8'd240} : s = 383;
	{8'd143,8'd241} : s = 384;
	{8'd143,8'd242} : s = 385;
	{8'd143,8'd243} : s = 386;
	{8'd143,8'd244} : s = 387;
	{8'd143,8'd245} : s = 388;
	{8'd143,8'd246} : s = 389;
	{8'd143,8'd247} : s = 390;
	{8'd143,8'd248} : s = 391;
	{8'd143,8'd249} : s = 392;
	{8'd143,8'd250} : s = 393;
	{8'd143,8'd251} : s = 394;
	{8'd143,8'd252} : s = 395;
	{8'd143,8'd253} : s = 396;
	{8'd143,8'd254} : s = 397;
	{8'd143,8'd255} : s = 398;
	{8'd144,8'd0} : s = 144;
	{8'd144,8'd1} : s = 145;
	{8'd144,8'd2} : s = 146;
	{8'd144,8'd3} : s = 147;
	{8'd144,8'd4} : s = 148;
	{8'd144,8'd5} : s = 149;
	{8'd144,8'd6} : s = 150;
	{8'd144,8'd7} : s = 151;
	{8'd144,8'd8} : s = 152;
	{8'd144,8'd9} : s = 153;
	{8'd144,8'd10} : s = 154;
	{8'd144,8'd11} : s = 155;
	{8'd144,8'd12} : s = 156;
	{8'd144,8'd13} : s = 157;
	{8'd144,8'd14} : s = 158;
	{8'd144,8'd15} : s = 159;
	{8'd144,8'd16} : s = 160;
	{8'd144,8'd17} : s = 161;
	{8'd144,8'd18} : s = 162;
	{8'd144,8'd19} : s = 163;
	{8'd144,8'd20} : s = 164;
	{8'd144,8'd21} : s = 165;
	{8'd144,8'd22} : s = 166;
	{8'd144,8'd23} : s = 167;
	{8'd144,8'd24} : s = 168;
	{8'd144,8'd25} : s = 169;
	{8'd144,8'd26} : s = 170;
	{8'd144,8'd27} : s = 171;
	{8'd144,8'd28} : s = 172;
	{8'd144,8'd29} : s = 173;
	{8'd144,8'd30} : s = 174;
	{8'd144,8'd31} : s = 175;
	{8'd144,8'd32} : s = 176;
	{8'd144,8'd33} : s = 177;
	{8'd144,8'd34} : s = 178;
	{8'd144,8'd35} : s = 179;
	{8'd144,8'd36} : s = 180;
	{8'd144,8'd37} : s = 181;
	{8'd144,8'd38} : s = 182;
	{8'd144,8'd39} : s = 183;
	{8'd144,8'd40} : s = 184;
	{8'd144,8'd41} : s = 185;
	{8'd144,8'd42} : s = 186;
	{8'd144,8'd43} : s = 187;
	{8'd144,8'd44} : s = 188;
	{8'd144,8'd45} : s = 189;
	{8'd144,8'd46} : s = 190;
	{8'd144,8'd47} : s = 191;
	{8'd144,8'd48} : s = 192;
	{8'd144,8'd49} : s = 193;
	{8'd144,8'd50} : s = 194;
	{8'd144,8'd51} : s = 195;
	{8'd144,8'd52} : s = 196;
	{8'd144,8'd53} : s = 197;
	{8'd144,8'd54} : s = 198;
	{8'd144,8'd55} : s = 199;
	{8'd144,8'd56} : s = 200;
	{8'd144,8'd57} : s = 201;
	{8'd144,8'd58} : s = 202;
	{8'd144,8'd59} : s = 203;
	{8'd144,8'd60} : s = 204;
	{8'd144,8'd61} : s = 205;
	{8'd144,8'd62} : s = 206;
	{8'd144,8'd63} : s = 207;
	{8'd144,8'd64} : s = 208;
	{8'd144,8'd65} : s = 209;
	{8'd144,8'd66} : s = 210;
	{8'd144,8'd67} : s = 211;
	{8'd144,8'd68} : s = 212;
	{8'd144,8'd69} : s = 213;
	{8'd144,8'd70} : s = 214;
	{8'd144,8'd71} : s = 215;
	{8'd144,8'd72} : s = 216;
	{8'd144,8'd73} : s = 217;
	{8'd144,8'd74} : s = 218;
	{8'd144,8'd75} : s = 219;
	{8'd144,8'd76} : s = 220;
	{8'd144,8'd77} : s = 221;
	{8'd144,8'd78} : s = 222;
	{8'd144,8'd79} : s = 223;
	{8'd144,8'd80} : s = 224;
	{8'd144,8'd81} : s = 225;
	{8'd144,8'd82} : s = 226;
	{8'd144,8'd83} : s = 227;
	{8'd144,8'd84} : s = 228;
	{8'd144,8'd85} : s = 229;
	{8'd144,8'd86} : s = 230;
	{8'd144,8'd87} : s = 231;
	{8'd144,8'd88} : s = 232;
	{8'd144,8'd89} : s = 233;
	{8'd144,8'd90} : s = 234;
	{8'd144,8'd91} : s = 235;
	{8'd144,8'd92} : s = 236;
	{8'd144,8'd93} : s = 237;
	{8'd144,8'd94} : s = 238;
	{8'd144,8'd95} : s = 239;
	{8'd144,8'd96} : s = 240;
	{8'd144,8'd97} : s = 241;
	{8'd144,8'd98} : s = 242;
	{8'd144,8'd99} : s = 243;
	{8'd144,8'd100} : s = 244;
	{8'd144,8'd101} : s = 245;
	{8'd144,8'd102} : s = 246;
	{8'd144,8'd103} : s = 247;
	{8'd144,8'd104} : s = 248;
	{8'd144,8'd105} : s = 249;
	{8'd144,8'd106} : s = 250;
	{8'd144,8'd107} : s = 251;
	{8'd144,8'd108} : s = 252;
	{8'd144,8'd109} : s = 253;
	{8'd144,8'd110} : s = 254;
	{8'd144,8'd111} : s = 255;
	{8'd144,8'd112} : s = 256;
	{8'd144,8'd113} : s = 257;
	{8'd144,8'd114} : s = 258;
	{8'd144,8'd115} : s = 259;
	{8'd144,8'd116} : s = 260;
	{8'd144,8'd117} : s = 261;
	{8'd144,8'd118} : s = 262;
	{8'd144,8'd119} : s = 263;
	{8'd144,8'd120} : s = 264;
	{8'd144,8'd121} : s = 265;
	{8'd144,8'd122} : s = 266;
	{8'd144,8'd123} : s = 267;
	{8'd144,8'd124} : s = 268;
	{8'd144,8'd125} : s = 269;
	{8'd144,8'd126} : s = 270;
	{8'd144,8'd127} : s = 271;
	{8'd144,8'd128} : s = 272;
	{8'd144,8'd129} : s = 273;
	{8'd144,8'd130} : s = 274;
	{8'd144,8'd131} : s = 275;
	{8'd144,8'd132} : s = 276;
	{8'd144,8'd133} : s = 277;
	{8'd144,8'd134} : s = 278;
	{8'd144,8'd135} : s = 279;
	{8'd144,8'd136} : s = 280;
	{8'd144,8'd137} : s = 281;
	{8'd144,8'd138} : s = 282;
	{8'd144,8'd139} : s = 283;
	{8'd144,8'd140} : s = 284;
	{8'd144,8'd141} : s = 285;
	{8'd144,8'd142} : s = 286;
	{8'd144,8'd143} : s = 287;
	{8'd144,8'd144} : s = 288;
	{8'd144,8'd145} : s = 289;
	{8'd144,8'd146} : s = 290;
	{8'd144,8'd147} : s = 291;
	{8'd144,8'd148} : s = 292;
	{8'd144,8'd149} : s = 293;
	{8'd144,8'd150} : s = 294;
	{8'd144,8'd151} : s = 295;
	{8'd144,8'd152} : s = 296;
	{8'd144,8'd153} : s = 297;
	{8'd144,8'd154} : s = 298;
	{8'd144,8'd155} : s = 299;
	{8'd144,8'd156} : s = 300;
	{8'd144,8'd157} : s = 301;
	{8'd144,8'd158} : s = 302;
	{8'd144,8'd159} : s = 303;
	{8'd144,8'd160} : s = 304;
	{8'd144,8'd161} : s = 305;
	{8'd144,8'd162} : s = 306;
	{8'd144,8'd163} : s = 307;
	{8'd144,8'd164} : s = 308;
	{8'd144,8'd165} : s = 309;
	{8'd144,8'd166} : s = 310;
	{8'd144,8'd167} : s = 311;
	{8'd144,8'd168} : s = 312;
	{8'd144,8'd169} : s = 313;
	{8'd144,8'd170} : s = 314;
	{8'd144,8'd171} : s = 315;
	{8'd144,8'd172} : s = 316;
	{8'd144,8'd173} : s = 317;
	{8'd144,8'd174} : s = 318;
	{8'd144,8'd175} : s = 319;
	{8'd144,8'd176} : s = 320;
	{8'd144,8'd177} : s = 321;
	{8'd144,8'd178} : s = 322;
	{8'd144,8'd179} : s = 323;
	{8'd144,8'd180} : s = 324;
	{8'd144,8'd181} : s = 325;
	{8'd144,8'd182} : s = 326;
	{8'd144,8'd183} : s = 327;
	{8'd144,8'd184} : s = 328;
	{8'd144,8'd185} : s = 329;
	{8'd144,8'd186} : s = 330;
	{8'd144,8'd187} : s = 331;
	{8'd144,8'd188} : s = 332;
	{8'd144,8'd189} : s = 333;
	{8'd144,8'd190} : s = 334;
	{8'd144,8'd191} : s = 335;
	{8'd144,8'd192} : s = 336;
	{8'd144,8'd193} : s = 337;
	{8'd144,8'd194} : s = 338;
	{8'd144,8'd195} : s = 339;
	{8'd144,8'd196} : s = 340;
	{8'd144,8'd197} : s = 341;
	{8'd144,8'd198} : s = 342;
	{8'd144,8'd199} : s = 343;
	{8'd144,8'd200} : s = 344;
	{8'd144,8'd201} : s = 345;
	{8'd144,8'd202} : s = 346;
	{8'd144,8'd203} : s = 347;
	{8'd144,8'd204} : s = 348;
	{8'd144,8'd205} : s = 349;
	{8'd144,8'd206} : s = 350;
	{8'd144,8'd207} : s = 351;
	{8'd144,8'd208} : s = 352;
	{8'd144,8'd209} : s = 353;
	{8'd144,8'd210} : s = 354;
	{8'd144,8'd211} : s = 355;
	{8'd144,8'd212} : s = 356;
	{8'd144,8'd213} : s = 357;
	{8'd144,8'd214} : s = 358;
	{8'd144,8'd215} : s = 359;
	{8'd144,8'd216} : s = 360;
	{8'd144,8'd217} : s = 361;
	{8'd144,8'd218} : s = 362;
	{8'd144,8'd219} : s = 363;
	{8'd144,8'd220} : s = 364;
	{8'd144,8'd221} : s = 365;
	{8'd144,8'd222} : s = 366;
	{8'd144,8'd223} : s = 367;
	{8'd144,8'd224} : s = 368;
	{8'd144,8'd225} : s = 369;
	{8'd144,8'd226} : s = 370;
	{8'd144,8'd227} : s = 371;
	{8'd144,8'd228} : s = 372;
	{8'd144,8'd229} : s = 373;
	{8'd144,8'd230} : s = 374;
	{8'd144,8'd231} : s = 375;
	{8'd144,8'd232} : s = 376;
	{8'd144,8'd233} : s = 377;
	{8'd144,8'd234} : s = 378;
	{8'd144,8'd235} : s = 379;
	{8'd144,8'd236} : s = 380;
	{8'd144,8'd237} : s = 381;
	{8'd144,8'd238} : s = 382;
	{8'd144,8'd239} : s = 383;
	{8'd144,8'd240} : s = 384;
	{8'd144,8'd241} : s = 385;
	{8'd144,8'd242} : s = 386;
	{8'd144,8'd243} : s = 387;
	{8'd144,8'd244} : s = 388;
	{8'd144,8'd245} : s = 389;
	{8'd144,8'd246} : s = 390;
	{8'd144,8'd247} : s = 391;
	{8'd144,8'd248} : s = 392;
	{8'd144,8'd249} : s = 393;
	{8'd144,8'd250} : s = 394;
	{8'd144,8'd251} : s = 395;
	{8'd144,8'd252} : s = 396;
	{8'd144,8'd253} : s = 397;
	{8'd144,8'd254} : s = 398;
	{8'd144,8'd255} : s = 399;
	{8'd145,8'd0} : s = 145;
	{8'd145,8'd1} : s = 146;
	{8'd145,8'd2} : s = 147;
	{8'd145,8'd3} : s = 148;
	{8'd145,8'd4} : s = 149;
	{8'd145,8'd5} : s = 150;
	{8'd145,8'd6} : s = 151;
	{8'd145,8'd7} : s = 152;
	{8'd145,8'd8} : s = 153;
	{8'd145,8'd9} : s = 154;
	{8'd145,8'd10} : s = 155;
	{8'd145,8'd11} : s = 156;
	{8'd145,8'd12} : s = 157;
	{8'd145,8'd13} : s = 158;
	{8'd145,8'd14} : s = 159;
	{8'd145,8'd15} : s = 160;
	{8'd145,8'd16} : s = 161;
	{8'd145,8'd17} : s = 162;
	{8'd145,8'd18} : s = 163;
	{8'd145,8'd19} : s = 164;
	{8'd145,8'd20} : s = 165;
	{8'd145,8'd21} : s = 166;
	{8'd145,8'd22} : s = 167;
	{8'd145,8'd23} : s = 168;
	{8'd145,8'd24} : s = 169;
	{8'd145,8'd25} : s = 170;
	{8'd145,8'd26} : s = 171;
	{8'd145,8'd27} : s = 172;
	{8'd145,8'd28} : s = 173;
	{8'd145,8'd29} : s = 174;
	{8'd145,8'd30} : s = 175;
	{8'd145,8'd31} : s = 176;
	{8'd145,8'd32} : s = 177;
	{8'd145,8'd33} : s = 178;
	{8'd145,8'd34} : s = 179;
	{8'd145,8'd35} : s = 180;
	{8'd145,8'd36} : s = 181;
	{8'd145,8'd37} : s = 182;
	{8'd145,8'd38} : s = 183;
	{8'd145,8'd39} : s = 184;
	{8'd145,8'd40} : s = 185;
	{8'd145,8'd41} : s = 186;
	{8'd145,8'd42} : s = 187;
	{8'd145,8'd43} : s = 188;
	{8'd145,8'd44} : s = 189;
	{8'd145,8'd45} : s = 190;
	{8'd145,8'd46} : s = 191;
	{8'd145,8'd47} : s = 192;
	{8'd145,8'd48} : s = 193;
	{8'd145,8'd49} : s = 194;
	{8'd145,8'd50} : s = 195;
	{8'd145,8'd51} : s = 196;
	{8'd145,8'd52} : s = 197;
	{8'd145,8'd53} : s = 198;
	{8'd145,8'd54} : s = 199;
	{8'd145,8'd55} : s = 200;
	{8'd145,8'd56} : s = 201;
	{8'd145,8'd57} : s = 202;
	{8'd145,8'd58} : s = 203;
	{8'd145,8'd59} : s = 204;
	{8'd145,8'd60} : s = 205;
	{8'd145,8'd61} : s = 206;
	{8'd145,8'd62} : s = 207;
	{8'd145,8'd63} : s = 208;
	{8'd145,8'd64} : s = 209;
	{8'd145,8'd65} : s = 210;
	{8'd145,8'd66} : s = 211;
	{8'd145,8'd67} : s = 212;
	{8'd145,8'd68} : s = 213;
	{8'd145,8'd69} : s = 214;
	{8'd145,8'd70} : s = 215;
	{8'd145,8'd71} : s = 216;
	{8'd145,8'd72} : s = 217;
	{8'd145,8'd73} : s = 218;
	{8'd145,8'd74} : s = 219;
	{8'd145,8'd75} : s = 220;
	{8'd145,8'd76} : s = 221;
	{8'd145,8'd77} : s = 222;
	{8'd145,8'd78} : s = 223;
	{8'd145,8'd79} : s = 224;
	{8'd145,8'd80} : s = 225;
	{8'd145,8'd81} : s = 226;
	{8'd145,8'd82} : s = 227;
	{8'd145,8'd83} : s = 228;
	{8'd145,8'd84} : s = 229;
	{8'd145,8'd85} : s = 230;
	{8'd145,8'd86} : s = 231;
	{8'd145,8'd87} : s = 232;
	{8'd145,8'd88} : s = 233;
	{8'd145,8'd89} : s = 234;
	{8'd145,8'd90} : s = 235;
	{8'd145,8'd91} : s = 236;
	{8'd145,8'd92} : s = 237;
	{8'd145,8'd93} : s = 238;
	{8'd145,8'd94} : s = 239;
	{8'd145,8'd95} : s = 240;
	{8'd145,8'd96} : s = 241;
	{8'd145,8'd97} : s = 242;
	{8'd145,8'd98} : s = 243;
	{8'd145,8'd99} : s = 244;
	{8'd145,8'd100} : s = 245;
	{8'd145,8'd101} : s = 246;
	{8'd145,8'd102} : s = 247;
	{8'd145,8'd103} : s = 248;
	{8'd145,8'd104} : s = 249;
	{8'd145,8'd105} : s = 250;
	{8'd145,8'd106} : s = 251;
	{8'd145,8'd107} : s = 252;
	{8'd145,8'd108} : s = 253;
	{8'd145,8'd109} : s = 254;
	{8'd145,8'd110} : s = 255;
	{8'd145,8'd111} : s = 256;
	{8'd145,8'd112} : s = 257;
	{8'd145,8'd113} : s = 258;
	{8'd145,8'd114} : s = 259;
	{8'd145,8'd115} : s = 260;
	{8'd145,8'd116} : s = 261;
	{8'd145,8'd117} : s = 262;
	{8'd145,8'd118} : s = 263;
	{8'd145,8'd119} : s = 264;
	{8'd145,8'd120} : s = 265;
	{8'd145,8'd121} : s = 266;
	{8'd145,8'd122} : s = 267;
	{8'd145,8'd123} : s = 268;
	{8'd145,8'd124} : s = 269;
	{8'd145,8'd125} : s = 270;
	{8'd145,8'd126} : s = 271;
	{8'd145,8'd127} : s = 272;
	{8'd145,8'd128} : s = 273;
	{8'd145,8'd129} : s = 274;
	{8'd145,8'd130} : s = 275;
	{8'd145,8'd131} : s = 276;
	{8'd145,8'd132} : s = 277;
	{8'd145,8'd133} : s = 278;
	{8'd145,8'd134} : s = 279;
	{8'd145,8'd135} : s = 280;
	{8'd145,8'd136} : s = 281;
	{8'd145,8'd137} : s = 282;
	{8'd145,8'd138} : s = 283;
	{8'd145,8'd139} : s = 284;
	{8'd145,8'd140} : s = 285;
	{8'd145,8'd141} : s = 286;
	{8'd145,8'd142} : s = 287;
	{8'd145,8'd143} : s = 288;
	{8'd145,8'd144} : s = 289;
	{8'd145,8'd145} : s = 290;
	{8'd145,8'd146} : s = 291;
	{8'd145,8'd147} : s = 292;
	{8'd145,8'd148} : s = 293;
	{8'd145,8'd149} : s = 294;
	{8'd145,8'd150} : s = 295;
	{8'd145,8'd151} : s = 296;
	{8'd145,8'd152} : s = 297;
	{8'd145,8'd153} : s = 298;
	{8'd145,8'd154} : s = 299;
	{8'd145,8'd155} : s = 300;
	{8'd145,8'd156} : s = 301;
	{8'd145,8'd157} : s = 302;
	{8'd145,8'd158} : s = 303;
	{8'd145,8'd159} : s = 304;
	{8'd145,8'd160} : s = 305;
	{8'd145,8'd161} : s = 306;
	{8'd145,8'd162} : s = 307;
	{8'd145,8'd163} : s = 308;
	{8'd145,8'd164} : s = 309;
	{8'd145,8'd165} : s = 310;
	{8'd145,8'd166} : s = 311;
	{8'd145,8'd167} : s = 312;
	{8'd145,8'd168} : s = 313;
	{8'd145,8'd169} : s = 314;
	{8'd145,8'd170} : s = 315;
	{8'd145,8'd171} : s = 316;
	{8'd145,8'd172} : s = 317;
	{8'd145,8'd173} : s = 318;
	{8'd145,8'd174} : s = 319;
	{8'd145,8'd175} : s = 320;
	{8'd145,8'd176} : s = 321;
	{8'd145,8'd177} : s = 322;
	{8'd145,8'd178} : s = 323;
	{8'd145,8'd179} : s = 324;
	{8'd145,8'd180} : s = 325;
	{8'd145,8'd181} : s = 326;
	{8'd145,8'd182} : s = 327;
	{8'd145,8'd183} : s = 328;
	{8'd145,8'd184} : s = 329;
	{8'd145,8'd185} : s = 330;
	{8'd145,8'd186} : s = 331;
	{8'd145,8'd187} : s = 332;
	{8'd145,8'd188} : s = 333;
	{8'd145,8'd189} : s = 334;
	{8'd145,8'd190} : s = 335;
	{8'd145,8'd191} : s = 336;
	{8'd145,8'd192} : s = 337;
	{8'd145,8'd193} : s = 338;
	{8'd145,8'd194} : s = 339;
	{8'd145,8'd195} : s = 340;
	{8'd145,8'd196} : s = 341;
	{8'd145,8'd197} : s = 342;
	{8'd145,8'd198} : s = 343;
	{8'd145,8'd199} : s = 344;
	{8'd145,8'd200} : s = 345;
	{8'd145,8'd201} : s = 346;
	{8'd145,8'd202} : s = 347;
	{8'd145,8'd203} : s = 348;
	{8'd145,8'd204} : s = 349;
	{8'd145,8'd205} : s = 350;
	{8'd145,8'd206} : s = 351;
	{8'd145,8'd207} : s = 352;
	{8'd145,8'd208} : s = 353;
	{8'd145,8'd209} : s = 354;
	{8'd145,8'd210} : s = 355;
	{8'd145,8'd211} : s = 356;
	{8'd145,8'd212} : s = 357;
	{8'd145,8'd213} : s = 358;
	{8'd145,8'd214} : s = 359;
	{8'd145,8'd215} : s = 360;
	{8'd145,8'd216} : s = 361;
	{8'd145,8'd217} : s = 362;
	{8'd145,8'd218} : s = 363;
	{8'd145,8'd219} : s = 364;
	{8'd145,8'd220} : s = 365;
	{8'd145,8'd221} : s = 366;
	{8'd145,8'd222} : s = 367;
	{8'd145,8'd223} : s = 368;
	{8'd145,8'd224} : s = 369;
	{8'd145,8'd225} : s = 370;
	{8'd145,8'd226} : s = 371;
	{8'd145,8'd227} : s = 372;
	{8'd145,8'd228} : s = 373;
	{8'd145,8'd229} : s = 374;
	{8'd145,8'd230} : s = 375;
	{8'd145,8'd231} : s = 376;
	{8'd145,8'd232} : s = 377;
	{8'd145,8'd233} : s = 378;
	{8'd145,8'd234} : s = 379;
	{8'd145,8'd235} : s = 380;
	{8'd145,8'd236} : s = 381;
	{8'd145,8'd237} : s = 382;
	{8'd145,8'd238} : s = 383;
	{8'd145,8'd239} : s = 384;
	{8'd145,8'd240} : s = 385;
	{8'd145,8'd241} : s = 386;
	{8'd145,8'd242} : s = 387;
	{8'd145,8'd243} : s = 388;
	{8'd145,8'd244} : s = 389;
	{8'd145,8'd245} : s = 390;
	{8'd145,8'd246} : s = 391;
	{8'd145,8'd247} : s = 392;
	{8'd145,8'd248} : s = 393;
	{8'd145,8'd249} : s = 394;
	{8'd145,8'd250} : s = 395;
	{8'd145,8'd251} : s = 396;
	{8'd145,8'd252} : s = 397;
	{8'd145,8'd253} : s = 398;
	{8'd145,8'd254} : s = 399;
	{8'd145,8'd255} : s = 400;
	{8'd146,8'd0} : s = 146;
	{8'd146,8'd1} : s = 147;
	{8'd146,8'd2} : s = 148;
	{8'd146,8'd3} : s = 149;
	{8'd146,8'd4} : s = 150;
	{8'd146,8'd5} : s = 151;
	{8'd146,8'd6} : s = 152;
	{8'd146,8'd7} : s = 153;
	{8'd146,8'd8} : s = 154;
	{8'd146,8'd9} : s = 155;
	{8'd146,8'd10} : s = 156;
	{8'd146,8'd11} : s = 157;
	{8'd146,8'd12} : s = 158;
	{8'd146,8'd13} : s = 159;
	{8'd146,8'd14} : s = 160;
	{8'd146,8'd15} : s = 161;
	{8'd146,8'd16} : s = 162;
	{8'd146,8'd17} : s = 163;
	{8'd146,8'd18} : s = 164;
	{8'd146,8'd19} : s = 165;
	{8'd146,8'd20} : s = 166;
	{8'd146,8'd21} : s = 167;
	{8'd146,8'd22} : s = 168;
	{8'd146,8'd23} : s = 169;
	{8'd146,8'd24} : s = 170;
	{8'd146,8'd25} : s = 171;
	{8'd146,8'd26} : s = 172;
	{8'd146,8'd27} : s = 173;
	{8'd146,8'd28} : s = 174;
	{8'd146,8'd29} : s = 175;
	{8'd146,8'd30} : s = 176;
	{8'd146,8'd31} : s = 177;
	{8'd146,8'd32} : s = 178;
	{8'd146,8'd33} : s = 179;
	{8'd146,8'd34} : s = 180;
	{8'd146,8'd35} : s = 181;
	{8'd146,8'd36} : s = 182;
	{8'd146,8'd37} : s = 183;
	{8'd146,8'd38} : s = 184;
	{8'd146,8'd39} : s = 185;
	{8'd146,8'd40} : s = 186;
	{8'd146,8'd41} : s = 187;
	{8'd146,8'd42} : s = 188;
	{8'd146,8'd43} : s = 189;
	{8'd146,8'd44} : s = 190;
	{8'd146,8'd45} : s = 191;
	{8'd146,8'd46} : s = 192;
	{8'd146,8'd47} : s = 193;
	{8'd146,8'd48} : s = 194;
	{8'd146,8'd49} : s = 195;
	{8'd146,8'd50} : s = 196;
	{8'd146,8'd51} : s = 197;
	{8'd146,8'd52} : s = 198;
	{8'd146,8'd53} : s = 199;
	{8'd146,8'd54} : s = 200;
	{8'd146,8'd55} : s = 201;
	{8'd146,8'd56} : s = 202;
	{8'd146,8'd57} : s = 203;
	{8'd146,8'd58} : s = 204;
	{8'd146,8'd59} : s = 205;
	{8'd146,8'd60} : s = 206;
	{8'd146,8'd61} : s = 207;
	{8'd146,8'd62} : s = 208;
	{8'd146,8'd63} : s = 209;
	{8'd146,8'd64} : s = 210;
	{8'd146,8'd65} : s = 211;
	{8'd146,8'd66} : s = 212;
	{8'd146,8'd67} : s = 213;
	{8'd146,8'd68} : s = 214;
	{8'd146,8'd69} : s = 215;
	{8'd146,8'd70} : s = 216;
	{8'd146,8'd71} : s = 217;
	{8'd146,8'd72} : s = 218;
	{8'd146,8'd73} : s = 219;
	{8'd146,8'd74} : s = 220;
	{8'd146,8'd75} : s = 221;
	{8'd146,8'd76} : s = 222;
	{8'd146,8'd77} : s = 223;
	{8'd146,8'd78} : s = 224;
	{8'd146,8'd79} : s = 225;
	{8'd146,8'd80} : s = 226;
	{8'd146,8'd81} : s = 227;
	{8'd146,8'd82} : s = 228;
	{8'd146,8'd83} : s = 229;
	{8'd146,8'd84} : s = 230;
	{8'd146,8'd85} : s = 231;
	{8'd146,8'd86} : s = 232;
	{8'd146,8'd87} : s = 233;
	{8'd146,8'd88} : s = 234;
	{8'd146,8'd89} : s = 235;
	{8'd146,8'd90} : s = 236;
	{8'd146,8'd91} : s = 237;
	{8'd146,8'd92} : s = 238;
	{8'd146,8'd93} : s = 239;
	{8'd146,8'd94} : s = 240;
	{8'd146,8'd95} : s = 241;
	{8'd146,8'd96} : s = 242;
	{8'd146,8'd97} : s = 243;
	{8'd146,8'd98} : s = 244;
	{8'd146,8'd99} : s = 245;
	{8'd146,8'd100} : s = 246;
	{8'd146,8'd101} : s = 247;
	{8'd146,8'd102} : s = 248;
	{8'd146,8'd103} : s = 249;
	{8'd146,8'd104} : s = 250;
	{8'd146,8'd105} : s = 251;
	{8'd146,8'd106} : s = 252;
	{8'd146,8'd107} : s = 253;
	{8'd146,8'd108} : s = 254;
	{8'd146,8'd109} : s = 255;
	{8'd146,8'd110} : s = 256;
	{8'd146,8'd111} : s = 257;
	{8'd146,8'd112} : s = 258;
	{8'd146,8'd113} : s = 259;
	{8'd146,8'd114} : s = 260;
	{8'd146,8'd115} : s = 261;
	{8'd146,8'd116} : s = 262;
	{8'd146,8'd117} : s = 263;
	{8'd146,8'd118} : s = 264;
	{8'd146,8'd119} : s = 265;
	{8'd146,8'd120} : s = 266;
	{8'd146,8'd121} : s = 267;
	{8'd146,8'd122} : s = 268;
	{8'd146,8'd123} : s = 269;
	{8'd146,8'd124} : s = 270;
	{8'd146,8'd125} : s = 271;
	{8'd146,8'd126} : s = 272;
	{8'd146,8'd127} : s = 273;
	{8'd146,8'd128} : s = 274;
	{8'd146,8'd129} : s = 275;
	{8'd146,8'd130} : s = 276;
	{8'd146,8'd131} : s = 277;
	{8'd146,8'd132} : s = 278;
	{8'd146,8'd133} : s = 279;
	{8'd146,8'd134} : s = 280;
	{8'd146,8'd135} : s = 281;
	{8'd146,8'd136} : s = 282;
	{8'd146,8'd137} : s = 283;
	{8'd146,8'd138} : s = 284;
	{8'd146,8'd139} : s = 285;
	{8'd146,8'd140} : s = 286;
	{8'd146,8'd141} : s = 287;
	{8'd146,8'd142} : s = 288;
	{8'd146,8'd143} : s = 289;
	{8'd146,8'd144} : s = 290;
	{8'd146,8'd145} : s = 291;
	{8'd146,8'd146} : s = 292;
	{8'd146,8'd147} : s = 293;
	{8'd146,8'd148} : s = 294;
	{8'd146,8'd149} : s = 295;
	{8'd146,8'd150} : s = 296;
	{8'd146,8'd151} : s = 297;
	{8'd146,8'd152} : s = 298;
	{8'd146,8'd153} : s = 299;
	{8'd146,8'd154} : s = 300;
	{8'd146,8'd155} : s = 301;
	{8'd146,8'd156} : s = 302;
	{8'd146,8'd157} : s = 303;
	{8'd146,8'd158} : s = 304;
	{8'd146,8'd159} : s = 305;
	{8'd146,8'd160} : s = 306;
	{8'd146,8'd161} : s = 307;
	{8'd146,8'd162} : s = 308;
	{8'd146,8'd163} : s = 309;
	{8'd146,8'd164} : s = 310;
	{8'd146,8'd165} : s = 311;
	{8'd146,8'd166} : s = 312;
	{8'd146,8'd167} : s = 313;
	{8'd146,8'd168} : s = 314;
	{8'd146,8'd169} : s = 315;
	{8'd146,8'd170} : s = 316;
	{8'd146,8'd171} : s = 317;
	{8'd146,8'd172} : s = 318;
	{8'd146,8'd173} : s = 319;
	{8'd146,8'd174} : s = 320;
	{8'd146,8'd175} : s = 321;
	{8'd146,8'd176} : s = 322;
	{8'd146,8'd177} : s = 323;
	{8'd146,8'd178} : s = 324;
	{8'd146,8'd179} : s = 325;
	{8'd146,8'd180} : s = 326;
	{8'd146,8'd181} : s = 327;
	{8'd146,8'd182} : s = 328;
	{8'd146,8'd183} : s = 329;
	{8'd146,8'd184} : s = 330;
	{8'd146,8'd185} : s = 331;
	{8'd146,8'd186} : s = 332;
	{8'd146,8'd187} : s = 333;
	{8'd146,8'd188} : s = 334;
	{8'd146,8'd189} : s = 335;
	{8'd146,8'd190} : s = 336;
	{8'd146,8'd191} : s = 337;
	{8'd146,8'd192} : s = 338;
	{8'd146,8'd193} : s = 339;
	{8'd146,8'd194} : s = 340;
	{8'd146,8'd195} : s = 341;
	{8'd146,8'd196} : s = 342;
	{8'd146,8'd197} : s = 343;
	{8'd146,8'd198} : s = 344;
	{8'd146,8'd199} : s = 345;
	{8'd146,8'd200} : s = 346;
	{8'd146,8'd201} : s = 347;
	{8'd146,8'd202} : s = 348;
	{8'd146,8'd203} : s = 349;
	{8'd146,8'd204} : s = 350;
	{8'd146,8'd205} : s = 351;
	{8'd146,8'd206} : s = 352;
	{8'd146,8'd207} : s = 353;
	{8'd146,8'd208} : s = 354;
	{8'd146,8'd209} : s = 355;
	{8'd146,8'd210} : s = 356;
	{8'd146,8'd211} : s = 357;
	{8'd146,8'd212} : s = 358;
	{8'd146,8'd213} : s = 359;
	{8'd146,8'd214} : s = 360;
	{8'd146,8'd215} : s = 361;
	{8'd146,8'd216} : s = 362;
	{8'd146,8'd217} : s = 363;
	{8'd146,8'd218} : s = 364;
	{8'd146,8'd219} : s = 365;
	{8'd146,8'd220} : s = 366;
	{8'd146,8'd221} : s = 367;
	{8'd146,8'd222} : s = 368;
	{8'd146,8'd223} : s = 369;
	{8'd146,8'd224} : s = 370;
	{8'd146,8'd225} : s = 371;
	{8'd146,8'd226} : s = 372;
	{8'd146,8'd227} : s = 373;
	{8'd146,8'd228} : s = 374;
	{8'd146,8'd229} : s = 375;
	{8'd146,8'd230} : s = 376;
	{8'd146,8'd231} : s = 377;
	{8'd146,8'd232} : s = 378;
	{8'd146,8'd233} : s = 379;
	{8'd146,8'd234} : s = 380;
	{8'd146,8'd235} : s = 381;
	{8'd146,8'd236} : s = 382;
	{8'd146,8'd237} : s = 383;
	{8'd146,8'd238} : s = 384;
	{8'd146,8'd239} : s = 385;
	{8'd146,8'd240} : s = 386;
	{8'd146,8'd241} : s = 387;
	{8'd146,8'd242} : s = 388;
	{8'd146,8'd243} : s = 389;
	{8'd146,8'd244} : s = 390;
	{8'd146,8'd245} : s = 391;
	{8'd146,8'd246} : s = 392;
	{8'd146,8'd247} : s = 393;
	{8'd146,8'd248} : s = 394;
	{8'd146,8'd249} : s = 395;
	{8'd146,8'd250} : s = 396;
	{8'd146,8'd251} : s = 397;
	{8'd146,8'd252} : s = 398;
	{8'd146,8'd253} : s = 399;
	{8'd146,8'd254} : s = 400;
	{8'd146,8'd255} : s = 401;
	{8'd147,8'd0} : s = 147;
	{8'd147,8'd1} : s = 148;
	{8'd147,8'd2} : s = 149;
	{8'd147,8'd3} : s = 150;
	{8'd147,8'd4} : s = 151;
	{8'd147,8'd5} : s = 152;
	{8'd147,8'd6} : s = 153;
	{8'd147,8'd7} : s = 154;
	{8'd147,8'd8} : s = 155;
	{8'd147,8'd9} : s = 156;
	{8'd147,8'd10} : s = 157;
	{8'd147,8'd11} : s = 158;
	{8'd147,8'd12} : s = 159;
	{8'd147,8'd13} : s = 160;
	{8'd147,8'd14} : s = 161;
	{8'd147,8'd15} : s = 162;
	{8'd147,8'd16} : s = 163;
	{8'd147,8'd17} : s = 164;
	{8'd147,8'd18} : s = 165;
	{8'd147,8'd19} : s = 166;
	{8'd147,8'd20} : s = 167;
	{8'd147,8'd21} : s = 168;
	{8'd147,8'd22} : s = 169;
	{8'd147,8'd23} : s = 170;
	{8'd147,8'd24} : s = 171;
	{8'd147,8'd25} : s = 172;
	{8'd147,8'd26} : s = 173;
	{8'd147,8'd27} : s = 174;
	{8'd147,8'd28} : s = 175;
	{8'd147,8'd29} : s = 176;
	{8'd147,8'd30} : s = 177;
	{8'd147,8'd31} : s = 178;
	{8'd147,8'd32} : s = 179;
	{8'd147,8'd33} : s = 180;
	{8'd147,8'd34} : s = 181;
	{8'd147,8'd35} : s = 182;
	{8'd147,8'd36} : s = 183;
	{8'd147,8'd37} : s = 184;
	{8'd147,8'd38} : s = 185;
	{8'd147,8'd39} : s = 186;
	{8'd147,8'd40} : s = 187;
	{8'd147,8'd41} : s = 188;
	{8'd147,8'd42} : s = 189;
	{8'd147,8'd43} : s = 190;
	{8'd147,8'd44} : s = 191;
	{8'd147,8'd45} : s = 192;
	{8'd147,8'd46} : s = 193;
	{8'd147,8'd47} : s = 194;
	{8'd147,8'd48} : s = 195;
	{8'd147,8'd49} : s = 196;
	{8'd147,8'd50} : s = 197;
	{8'd147,8'd51} : s = 198;
	{8'd147,8'd52} : s = 199;
	{8'd147,8'd53} : s = 200;
	{8'd147,8'd54} : s = 201;
	{8'd147,8'd55} : s = 202;
	{8'd147,8'd56} : s = 203;
	{8'd147,8'd57} : s = 204;
	{8'd147,8'd58} : s = 205;
	{8'd147,8'd59} : s = 206;
	{8'd147,8'd60} : s = 207;
	{8'd147,8'd61} : s = 208;
	{8'd147,8'd62} : s = 209;
	{8'd147,8'd63} : s = 210;
	{8'd147,8'd64} : s = 211;
	{8'd147,8'd65} : s = 212;
	{8'd147,8'd66} : s = 213;
	{8'd147,8'd67} : s = 214;
	{8'd147,8'd68} : s = 215;
	{8'd147,8'd69} : s = 216;
	{8'd147,8'd70} : s = 217;
	{8'd147,8'd71} : s = 218;
	{8'd147,8'd72} : s = 219;
	{8'd147,8'd73} : s = 220;
	{8'd147,8'd74} : s = 221;
	{8'd147,8'd75} : s = 222;
	{8'd147,8'd76} : s = 223;
	{8'd147,8'd77} : s = 224;
	{8'd147,8'd78} : s = 225;
	{8'd147,8'd79} : s = 226;
	{8'd147,8'd80} : s = 227;
	{8'd147,8'd81} : s = 228;
	{8'd147,8'd82} : s = 229;
	{8'd147,8'd83} : s = 230;
	{8'd147,8'd84} : s = 231;
	{8'd147,8'd85} : s = 232;
	{8'd147,8'd86} : s = 233;
	{8'd147,8'd87} : s = 234;
	{8'd147,8'd88} : s = 235;
	{8'd147,8'd89} : s = 236;
	{8'd147,8'd90} : s = 237;
	{8'd147,8'd91} : s = 238;
	{8'd147,8'd92} : s = 239;
	{8'd147,8'd93} : s = 240;
	{8'd147,8'd94} : s = 241;
	{8'd147,8'd95} : s = 242;
	{8'd147,8'd96} : s = 243;
	{8'd147,8'd97} : s = 244;
	{8'd147,8'd98} : s = 245;
	{8'd147,8'd99} : s = 246;
	{8'd147,8'd100} : s = 247;
	{8'd147,8'd101} : s = 248;
	{8'd147,8'd102} : s = 249;
	{8'd147,8'd103} : s = 250;
	{8'd147,8'd104} : s = 251;
	{8'd147,8'd105} : s = 252;
	{8'd147,8'd106} : s = 253;
	{8'd147,8'd107} : s = 254;
	{8'd147,8'd108} : s = 255;
	{8'd147,8'd109} : s = 256;
	{8'd147,8'd110} : s = 257;
	{8'd147,8'd111} : s = 258;
	{8'd147,8'd112} : s = 259;
	{8'd147,8'd113} : s = 260;
	{8'd147,8'd114} : s = 261;
	{8'd147,8'd115} : s = 262;
	{8'd147,8'd116} : s = 263;
	{8'd147,8'd117} : s = 264;
	{8'd147,8'd118} : s = 265;
	{8'd147,8'd119} : s = 266;
	{8'd147,8'd120} : s = 267;
	{8'd147,8'd121} : s = 268;
	{8'd147,8'd122} : s = 269;
	{8'd147,8'd123} : s = 270;
	{8'd147,8'd124} : s = 271;
	{8'd147,8'd125} : s = 272;
	{8'd147,8'd126} : s = 273;
	{8'd147,8'd127} : s = 274;
	{8'd147,8'd128} : s = 275;
	{8'd147,8'd129} : s = 276;
	{8'd147,8'd130} : s = 277;
	{8'd147,8'd131} : s = 278;
	{8'd147,8'd132} : s = 279;
	{8'd147,8'd133} : s = 280;
	{8'd147,8'd134} : s = 281;
	{8'd147,8'd135} : s = 282;
	{8'd147,8'd136} : s = 283;
	{8'd147,8'd137} : s = 284;
	{8'd147,8'd138} : s = 285;
	{8'd147,8'd139} : s = 286;
	{8'd147,8'd140} : s = 287;
	{8'd147,8'd141} : s = 288;
	{8'd147,8'd142} : s = 289;
	{8'd147,8'd143} : s = 290;
	{8'd147,8'd144} : s = 291;
	{8'd147,8'd145} : s = 292;
	{8'd147,8'd146} : s = 293;
	{8'd147,8'd147} : s = 294;
	{8'd147,8'd148} : s = 295;
	{8'd147,8'd149} : s = 296;
	{8'd147,8'd150} : s = 297;
	{8'd147,8'd151} : s = 298;
	{8'd147,8'd152} : s = 299;
	{8'd147,8'd153} : s = 300;
	{8'd147,8'd154} : s = 301;
	{8'd147,8'd155} : s = 302;
	{8'd147,8'd156} : s = 303;
	{8'd147,8'd157} : s = 304;
	{8'd147,8'd158} : s = 305;
	{8'd147,8'd159} : s = 306;
	{8'd147,8'd160} : s = 307;
	{8'd147,8'd161} : s = 308;
	{8'd147,8'd162} : s = 309;
	{8'd147,8'd163} : s = 310;
	{8'd147,8'd164} : s = 311;
	{8'd147,8'd165} : s = 312;
	{8'd147,8'd166} : s = 313;
	{8'd147,8'd167} : s = 314;
	{8'd147,8'd168} : s = 315;
	{8'd147,8'd169} : s = 316;
	{8'd147,8'd170} : s = 317;
	{8'd147,8'd171} : s = 318;
	{8'd147,8'd172} : s = 319;
	{8'd147,8'd173} : s = 320;
	{8'd147,8'd174} : s = 321;
	{8'd147,8'd175} : s = 322;
	{8'd147,8'd176} : s = 323;
	{8'd147,8'd177} : s = 324;
	{8'd147,8'd178} : s = 325;
	{8'd147,8'd179} : s = 326;
	{8'd147,8'd180} : s = 327;
	{8'd147,8'd181} : s = 328;
	{8'd147,8'd182} : s = 329;
	{8'd147,8'd183} : s = 330;
	{8'd147,8'd184} : s = 331;
	{8'd147,8'd185} : s = 332;
	{8'd147,8'd186} : s = 333;
	{8'd147,8'd187} : s = 334;
	{8'd147,8'd188} : s = 335;
	{8'd147,8'd189} : s = 336;
	{8'd147,8'd190} : s = 337;
	{8'd147,8'd191} : s = 338;
	{8'd147,8'd192} : s = 339;
	{8'd147,8'd193} : s = 340;
	{8'd147,8'd194} : s = 341;
	{8'd147,8'd195} : s = 342;
	{8'd147,8'd196} : s = 343;
	{8'd147,8'd197} : s = 344;
	{8'd147,8'd198} : s = 345;
	{8'd147,8'd199} : s = 346;
	{8'd147,8'd200} : s = 347;
	{8'd147,8'd201} : s = 348;
	{8'd147,8'd202} : s = 349;
	{8'd147,8'd203} : s = 350;
	{8'd147,8'd204} : s = 351;
	{8'd147,8'd205} : s = 352;
	{8'd147,8'd206} : s = 353;
	{8'd147,8'd207} : s = 354;
	{8'd147,8'd208} : s = 355;
	{8'd147,8'd209} : s = 356;
	{8'd147,8'd210} : s = 357;
	{8'd147,8'd211} : s = 358;
	{8'd147,8'd212} : s = 359;
	{8'd147,8'd213} : s = 360;
	{8'd147,8'd214} : s = 361;
	{8'd147,8'd215} : s = 362;
	{8'd147,8'd216} : s = 363;
	{8'd147,8'd217} : s = 364;
	{8'd147,8'd218} : s = 365;
	{8'd147,8'd219} : s = 366;
	{8'd147,8'd220} : s = 367;
	{8'd147,8'd221} : s = 368;
	{8'd147,8'd222} : s = 369;
	{8'd147,8'd223} : s = 370;
	{8'd147,8'd224} : s = 371;
	{8'd147,8'd225} : s = 372;
	{8'd147,8'd226} : s = 373;
	{8'd147,8'd227} : s = 374;
	{8'd147,8'd228} : s = 375;
	{8'd147,8'd229} : s = 376;
	{8'd147,8'd230} : s = 377;
	{8'd147,8'd231} : s = 378;
	{8'd147,8'd232} : s = 379;
	{8'd147,8'd233} : s = 380;
	{8'd147,8'd234} : s = 381;
	{8'd147,8'd235} : s = 382;
	{8'd147,8'd236} : s = 383;
	{8'd147,8'd237} : s = 384;
	{8'd147,8'd238} : s = 385;
	{8'd147,8'd239} : s = 386;
	{8'd147,8'd240} : s = 387;
	{8'd147,8'd241} : s = 388;
	{8'd147,8'd242} : s = 389;
	{8'd147,8'd243} : s = 390;
	{8'd147,8'd244} : s = 391;
	{8'd147,8'd245} : s = 392;
	{8'd147,8'd246} : s = 393;
	{8'd147,8'd247} : s = 394;
	{8'd147,8'd248} : s = 395;
	{8'd147,8'd249} : s = 396;
	{8'd147,8'd250} : s = 397;
	{8'd147,8'd251} : s = 398;
	{8'd147,8'd252} : s = 399;
	{8'd147,8'd253} : s = 400;
	{8'd147,8'd254} : s = 401;
	{8'd147,8'd255} : s = 402;
	{8'd148,8'd0} : s = 148;
	{8'd148,8'd1} : s = 149;
	{8'd148,8'd2} : s = 150;
	{8'd148,8'd3} : s = 151;
	{8'd148,8'd4} : s = 152;
	{8'd148,8'd5} : s = 153;
	{8'd148,8'd6} : s = 154;
	{8'd148,8'd7} : s = 155;
	{8'd148,8'd8} : s = 156;
	{8'd148,8'd9} : s = 157;
	{8'd148,8'd10} : s = 158;
	{8'd148,8'd11} : s = 159;
	{8'd148,8'd12} : s = 160;
	{8'd148,8'd13} : s = 161;
	{8'd148,8'd14} : s = 162;
	{8'd148,8'd15} : s = 163;
	{8'd148,8'd16} : s = 164;
	{8'd148,8'd17} : s = 165;
	{8'd148,8'd18} : s = 166;
	{8'd148,8'd19} : s = 167;
	{8'd148,8'd20} : s = 168;
	{8'd148,8'd21} : s = 169;
	{8'd148,8'd22} : s = 170;
	{8'd148,8'd23} : s = 171;
	{8'd148,8'd24} : s = 172;
	{8'd148,8'd25} : s = 173;
	{8'd148,8'd26} : s = 174;
	{8'd148,8'd27} : s = 175;
	{8'd148,8'd28} : s = 176;
	{8'd148,8'd29} : s = 177;
	{8'd148,8'd30} : s = 178;
	{8'd148,8'd31} : s = 179;
	{8'd148,8'd32} : s = 180;
	{8'd148,8'd33} : s = 181;
	{8'd148,8'd34} : s = 182;
	{8'd148,8'd35} : s = 183;
	{8'd148,8'd36} : s = 184;
	{8'd148,8'd37} : s = 185;
	{8'd148,8'd38} : s = 186;
	{8'd148,8'd39} : s = 187;
	{8'd148,8'd40} : s = 188;
	{8'd148,8'd41} : s = 189;
	{8'd148,8'd42} : s = 190;
	{8'd148,8'd43} : s = 191;
	{8'd148,8'd44} : s = 192;
	{8'd148,8'd45} : s = 193;
	{8'd148,8'd46} : s = 194;
	{8'd148,8'd47} : s = 195;
	{8'd148,8'd48} : s = 196;
	{8'd148,8'd49} : s = 197;
	{8'd148,8'd50} : s = 198;
	{8'd148,8'd51} : s = 199;
	{8'd148,8'd52} : s = 200;
	{8'd148,8'd53} : s = 201;
	{8'd148,8'd54} : s = 202;
	{8'd148,8'd55} : s = 203;
	{8'd148,8'd56} : s = 204;
	{8'd148,8'd57} : s = 205;
	{8'd148,8'd58} : s = 206;
	{8'd148,8'd59} : s = 207;
	{8'd148,8'd60} : s = 208;
	{8'd148,8'd61} : s = 209;
	{8'd148,8'd62} : s = 210;
	{8'd148,8'd63} : s = 211;
	{8'd148,8'd64} : s = 212;
	{8'd148,8'd65} : s = 213;
	{8'd148,8'd66} : s = 214;
	{8'd148,8'd67} : s = 215;
	{8'd148,8'd68} : s = 216;
	{8'd148,8'd69} : s = 217;
	{8'd148,8'd70} : s = 218;
	{8'd148,8'd71} : s = 219;
	{8'd148,8'd72} : s = 220;
	{8'd148,8'd73} : s = 221;
	{8'd148,8'd74} : s = 222;
	{8'd148,8'd75} : s = 223;
	{8'd148,8'd76} : s = 224;
	{8'd148,8'd77} : s = 225;
	{8'd148,8'd78} : s = 226;
	{8'd148,8'd79} : s = 227;
	{8'd148,8'd80} : s = 228;
	{8'd148,8'd81} : s = 229;
	{8'd148,8'd82} : s = 230;
	{8'd148,8'd83} : s = 231;
	{8'd148,8'd84} : s = 232;
	{8'd148,8'd85} : s = 233;
	{8'd148,8'd86} : s = 234;
	{8'd148,8'd87} : s = 235;
	{8'd148,8'd88} : s = 236;
	{8'd148,8'd89} : s = 237;
	{8'd148,8'd90} : s = 238;
	{8'd148,8'd91} : s = 239;
	{8'd148,8'd92} : s = 240;
	{8'd148,8'd93} : s = 241;
	{8'd148,8'd94} : s = 242;
	{8'd148,8'd95} : s = 243;
	{8'd148,8'd96} : s = 244;
	{8'd148,8'd97} : s = 245;
	{8'd148,8'd98} : s = 246;
	{8'd148,8'd99} : s = 247;
	{8'd148,8'd100} : s = 248;
	{8'd148,8'd101} : s = 249;
	{8'd148,8'd102} : s = 250;
	{8'd148,8'd103} : s = 251;
	{8'd148,8'd104} : s = 252;
	{8'd148,8'd105} : s = 253;
	{8'd148,8'd106} : s = 254;
	{8'd148,8'd107} : s = 255;
	{8'd148,8'd108} : s = 256;
	{8'd148,8'd109} : s = 257;
	{8'd148,8'd110} : s = 258;
	{8'd148,8'd111} : s = 259;
	{8'd148,8'd112} : s = 260;
	{8'd148,8'd113} : s = 261;
	{8'd148,8'd114} : s = 262;
	{8'd148,8'd115} : s = 263;
	{8'd148,8'd116} : s = 264;
	{8'd148,8'd117} : s = 265;
	{8'd148,8'd118} : s = 266;
	{8'd148,8'd119} : s = 267;
	{8'd148,8'd120} : s = 268;
	{8'd148,8'd121} : s = 269;
	{8'd148,8'd122} : s = 270;
	{8'd148,8'd123} : s = 271;
	{8'd148,8'd124} : s = 272;
	{8'd148,8'd125} : s = 273;
	{8'd148,8'd126} : s = 274;
	{8'd148,8'd127} : s = 275;
	{8'd148,8'd128} : s = 276;
	{8'd148,8'd129} : s = 277;
	{8'd148,8'd130} : s = 278;
	{8'd148,8'd131} : s = 279;
	{8'd148,8'd132} : s = 280;
	{8'd148,8'd133} : s = 281;
	{8'd148,8'd134} : s = 282;
	{8'd148,8'd135} : s = 283;
	{8'd148,8'd136} : s = 284;
	{8'd148,8'd137} : s = 285;
	{8'd148,8'd138} : s = 286;
	{8'd148,8'd139} : s = 287;
	{8'd148,8'd140} : s = 288;
	{8'd148,8'd141} : s = 289;
	{8'd148,8'd142} : s = 290;
	{8'd148,8'd143} : s = 291;
	{8'd148,8'd144} : s = 292;
	{8'd148,8'd145} : s = 293;
	{8'd148,8'd146} : s = 294;
	{8'd148,8'd147} : s = 295;
	{8'd148,8'd148} : s = 296;
	{8'd148,8'd149} : s = 297;
	{8'd148,8'd150} : s = 298;
	{8'd148,8'd151} : s = 299;
	{8'd148,8'd152} : s = 300;
	{8'd148,8'd153} : s = 301;
	{8'd148,8'd154} : s = 302;
	{8'd148,8'd155} : s = 303;
	{8'd148,8'd156} : s = 304;
	{8'd148,8'd157} : s = 305;
	{8'd148,8'd158} : s = 306;
	{8'd148,8'd159} : s = 307;
	{8'd148,8'd160} : s = 308;
	{8'd148,8'd161} : s = 309;
	{8'd148,8'd162} : s = 310;
	{8'd148,8'd163} : s = 311;
	{8'd148,8'd164} : s = 312;
	{8'd148,8'd165} : s = 313;
	{8'd148,8'd166} : s = 314;
	{8'd148,8'd167} : s = 315;
	{8'd148,8'd168} : s = 316;
	{8'd148,8'd169} : s = 317;
	{8'd148,8'd170} : s = 318;
	{8'd148,8'd171} : s = 319;
	{8'd148,8'd172} : s = 320;
	{8'd148,8'd173} : s = 321;
	{8'd148,8'd174} : s = 322;
	{8'd148,8'd175} : s = 323;
	{8'd148,8'd176} : s = 324;
	{8'd148,8'd177} : s = 325;
	{8'd148,8'd178} : s = 326;
	{8'd148,8'd179} : s = 327;
	{8'd148,8'd180} : s = 328;
	{8'd148,8'd181} : s = 329;
	{8'd148,8'd182} : s = 330;
	{8'd148,8'd183} : s = 331;
	{8'd148,8'd184} : s = 332;
	{8'd148,8'd185} : s = 333;
	{8'd148,8'd186} : s = 334;
	{8'd148,8'd187} : s = 335;
	{8'd148,8'd188} : s = 336;
	{8'd148,8'd189} : s = 337;
	{8'd148,8'd190} : s = 338;
	{8'd148,8'd191} : s = 339;
	{8'd148,8'd192} : s = 340;
	{8'd148,8'd193} : s = 341;
	{8'd148,8'd194} : s = 342;
	{8'd148,8'd195} : s = 343;
	{8'd148,8'd196} : s = 344;
	{8'd148,8'd197} : s = 345;
	{8'd148,8'd198} : s = 346;
	{8'd148,8'd199} : s = 347;
	{8'd148,8'd200} : s = 348;
	{8'd148,8'd201} : s = 349;
	{8'd148,8'd202} : s = 350;
	{8'd148,8'd203} : s = 351;
	{8'd148,8'd204} : s = 352;
	{8'd148,8'd205} : s = 353;
	{8'd148,8'd206} : s = 354;
	{8'd148,8'd207} : s = 355;
	{8'd148,8'd208} : s = 356;
	{8'd148,8'd209} : s = 357;
	{8'd148,8'd210} : s = 358;
	{8'd148,8'd211} : s = 359;
	{8'd148,8'd212} : s = 360;
	{8'd148,8'd213} : s = 361;
	{8'd148,8'd214} : s = 362;
	{8'd148,8'd215} : s = 363;
	{8'd148,8'd216} : s = 364;
	{8'd148,8'd217} : s = 365;
	{8'd148,8'd218} : s = 366;
	{8'd148,8'd219} : s = 367;
	{8'd148,8'd220} : s = 368;
	{8'd148,8'd221} : s = 369;
	{8'd148,8'd222} : s = 370;
	{8'd148,8'd223} : s = 371;
	{8'd148,8'd224} : s = 372;
	{8'd148,8'd225} : s = 373;
	{8'd148,8'd226} : s = 374;
	{8'd148,8'd227} : s = 375;
	{8'd148,8'd228} : s = 376;
	{8'd148,8'd229} : s = 377;
	{8'd148,8'd230} : s = 378;
	{8'd148,8'd231} : s = 379;
	{8'd148,8'd232} : s = 380;
	{8'd148,8'd233} : s = 381;
	{8'd148,8'd234} : s = 382;
	{8'd148,8'd235} : s = 383;
	{8'd148,8'd236} : s = 384;
	{8'd148,8'd237} : s = 385;
	{8'd148,8'd238} : s = 386;
	{8'd148,8'd239} : s = 387;
	{8'd148,8'd240} : s = 388;
	{8'd148,8'd241} : s = 389;
	{8'd148,8'd242} : s = 390;
	{8'd148,8'd243} : s = 391;
	{8'd148,8'd244} : s = 392;
	{8'd148,8'd245} : s = 393;
	{8'd148,8'd246} : s = 394;
	{8'd148,8'd247} : s = 395;
	{8'd148,8'd248} : s = 396;
	{8'd148,8'd249} : s = 397;
	{8'd148,8'd250} : s = 398;
	{8'd148,8'd251} : s = 399;
	{8'd148,8'd252} : s = 400;
	{8'd148,8'd253} : s = 401;
	{8'd148,8'd254} : s = 402;
	{8'd148,8'd255} : s = 403;
	{8'd149,8'd0} : s = 149;
	{8'd149,8'd1} : s = 150;
	{8'd149,8'd2} : s = 151;
	{8'd149,8'd3} : s = 152;
	{8'd149,8'd4} : s = 153;
	{8'd149,8'd5} : s = 154;
	{8'd149,8'd6} : s = 155;
	{8'd149,8'd7} : s = 156;
	{8'd149,8'd8} : s = 157;
	{8'd149,8'd9} : s = 158;
	{8'd149,8'd10} : s = 159;
	{8'd149,8'd11} : s = 160;
	{8'd149,8'd12} : s = 161;
	{8'd149,8'd13} : s = 162;
	{8'd149,8'd14} : s = 163;
	{8'd149,8'd15} : s = 164;
	{8'd149,8'd16} : s = 165;
	{8'd149,8'd17} : s = 166;
	{8'd149,8'd18} : s = 167;
	{8'd149,8'd19} : s = 168;
	{8'd149,8'd20} : s = 169;
	{8'd149,8'd21} : s = 170;
	{8'd149,8'd22} : s = 171;
	{8'd149,8'd23} : s = 172;
	{8'd149,8'd24} : s = 173;
	{8'd149,8'd25} : s = 174;
	{8'd149,8'd26} : s = 175;
	{8'd149,8'd27} : s = 176;
	{8'd149,8'd28} : s = 177;
	{8'd149,8'd29} : s = 178;
	{8'd149,8'd30} : s = 179;
	{8'd149,8'd31} : s = 180;
	{8'd149,8'd32} : s = 181;
	{8'd149,8'd33} : s = 182;
	{8'd149,8'd34} : s = 183;
	{8'd149,8'd35} : s = 184;
	{8'd149,8'd36} : s = 185;
	{8'd149,8'd37} : s = 186;
	{8'd149,8'd38} : s = 187;
	{8'd149,8'd39} : s = 188;
	{8'd149,8'd40} : s = 189;
	{8'd149,8'd41} : s = 190;
	{8'd149,8'd42} : s = 191;
	{8'd149,8'd43} : s = 192;
	{8'd149,8'd44} : s = 193;
	{8'd149,8'd45} : s = 194;
	{8'd149,8'd46} : s = 195;
	{8'd149,8'd47} : s = 196;
	{8'd149,8'd48} : s = 197;
	{8'd149,8'd49} : s = 198;
	{8'd149,8'd50} : s = 199;
	{8'd149,8'd51} : s = 200;
	{8'd149,8'd52} : s = 201;
	{8'd149,8'd53} : s = 202;
	{8'd149,8'd54} : s = 203;
	{8'd149,8'd55} : s = 204;
	{8'd149,8'd56} : s = 205;
	{8'd149,8'd57} : s = 206;
	{8'd149,8'd58} : s = 207;
	{8'd149,8'd59} : s = 208;
	{8'd149,8'd60} : s = 209;
	{8'd149,8'd61} : s = 210;
	{8'd149,8'd62} : s = 211;
	{8'd149,8'd63} : s = 212;
	{8'd149,8'd64} : s = 213;
	{8'd149,8'd65} : s = 214;
	{8'd149,8'd66} : s = 215;
	{8'd149,8'd67} : s = 216;
	{8'd149,8'd68} : s = 217;
	{8'd149,8'd69} : s = 218;
	{8'd149,8'd70} : s = 219;
	{8'd149,8'd71} : s = 220;
	{8'd149,8'd72} : s = 221;
	{8'd149,8'd73} : s = 222;
	{8'd149,8'd74} : s = 223;
	{8'd149,8'd75} : s = 224;
	{8'd149,8'd76} : s = 225;
	{8'd149,8'd77} : s = 226;
	{8'd149,8'd78} : s = 227;
	{8'd149,8'd79} : s = 228;
	{8'd149,8'd80} : s = 229;
	{8'd149,8'd81} : s = 230;
	{8'd149,8'd82} : s = 231;
	{8'd149,8'd83} : s = 232;
	{8'd149,8'd84} : s = 233;
	{8'd149,8'd85} : s = 234;
	{8'd149,8'd86} : s = 235;
	{8'd149,8'd87} : s = 236;
	{8'd149,8'd88} : s = 237;
	{8'd149,8'd89} : s = 238;
	{8'd149,8'd90} : s = 239;
	{8'd149,8'd91} : s = 240;
	{8'd149,8'd92} : s = 241;
	{8'd149,8'd93} : s = 242;
	{8'd149,8'd94} : s = 243;
	{8'd149,8'd95} : s = 244;
	{8'd149,8'd96} : s = 245;
	{8'd149,8'd97} : s = 246;
	{8'd149,8'd98} : s = 247;
	{8'd149,8'd99} : s = 248;
	{8'd149,8'd100} : s = 249;
	{8'd149,8'd101} : s = 250;
	{8'd149,8'd102} : s = 251;
	{8'd149,8'd103} : s = 252;
	{8'd149,8'd104} : s = 253;
	{8'd149,8'd105} : s = 254;
	{8'd149,8'd106} : s = 255;
	{8'd149,8'd107} : s = 256;
	{8'd149,8'd108} : s = 257;
	{8'd149,8'd109} : s = 258;
	{8'd149,8'd110} : s = 259;
	{8'd149,8'd111} : s = 260;
	{8'd149,8'd112} : s = 261;
	{8'd149,8'd113} : s = 262;
	{8'd149,8'd114} : s = 263;
	{8'd149,8'd115} : s = 264;
	{8'd149,8'd116} : s = 265;
	{8'd149,8'd117} : s = 266;
	{8'd149,8'd118} : s = 267;
	{8'd149,8'd119} : s = 268;
	{8'd149,8'd120} : s = 269;
	{8'd149,8'd121} : s = 270;
	{8'd149,8'd122} : s = 271;
	{8'd149,8'd123} : s = 272;
	{8'd149,8'd124} : s = 273;
	{8'd149,8'd125} : s = 274;
	{8'd149,8'd126} : s = 275;
	{8'd149,8'd127} : s = 276;
	{8'd149,8'd128} : s = 277;
	{8'd149,8'd129} : s = 278;
	{8'd149,8'd130} : s = 279;
	{8'd149,8'd131} : s = 280;
	{8'd149,8'd132} : s = 281;
	{8'd149,8'd133} : s = 282;
	{8'd149,8'd134} : s = 283;
	{8'd149,8'd135} : s = 284;
	{8'd149,8'd136} : s = 285;
	{8'd149,8'd137} : s = 286;
	{8'd149,8'd138} : s = 287;
	{8'd149,8'd139} : s = 288;
	{8'd149,8'd140} : s = 289;
	{8'd149,8'd141} : s = 290;
	{8'd149,8'd142} : s = 291;
	{8'd149,8'd143} : s = 292;
	{8'd149,8'd144} : s = 293;
	{8'd149,8'd145} : s = 294;
	{8'd149,8'd146} : s = 295;
	{8'd149,8'd147} : s = 296;
	{8'd149,8'd148} : s = 297;
	{8'd149,8'd149} : s = 298;
	{8'd149,8'd150} : s = 299;
	{8'd149,8'd151} : s = 300;
	{8'd149,8'd152} : s = 301;
	{8'd149,8'd153} : s = 302;
	{8'd149,8'd154} : s = 303;
	{8'd149,8'd155} : s = 304;
	{8'd149,8'd156} : s = 305;
	{8'd149,8'd157} : s = 306;
	{8'd149,8'd158} : s = 307;
	{8'd149,8'd159} : s = 308;
	{8'd149,8'd160} : s = 309;
	{8'd149,8'd161} : s = 310;
	{8'd149,8'd162} : s = 311;
	{8'd149,8'd163} : s = 312;
	{8'd149,8'd164} : s = 313;
	{8'd149,8'd165} : s = 314;
	{8'd149,8'd166} : s = 315;
	{8'd149,8'd167} : s = 316;
	{8'd149,8'd168} : s = 317;
	{8'd149,8'd169} : s = 318;
	{8'd149,8'd170} : s = 319;
	{8'd149,8'd171} : s = 320;
	{8'd149,8'd172} : s = 321;
	{8'd149,8'd173} : s = 322;
	{8'd149,8'd174} : s = 323;
	{8'd149,8'd175} : s = 324;
	{8'd149,8'd176} : s = 325;
	{8'd149,8'd177} : s = 326;
	{8'd149,8'd178} : s = 327;
	{8'd149,8'd179} : s = 328;
	{8'd149,8'd180} : s = 329;
	{8'd149,8'd181} : s = 330;
	{8'd149,8'd182} : s = 331;
	{8'd149,8'd183} : s = 332;
	{8'd149,8'd184} : s = 333;
	{8'd149,8'd185} : s = 334;
	{8'd149,8'd186} : s = 335;
	{8'd149,8'd187} : s = 336;
	{8'd149,8'd188} : s = 337;
	{8'd149,8'd189} : s = 338;
	{8'd149,8'd190} : s = 339;
	{8'd149,8'd191} : s = 340;
	{8'd149,8'd192} : s = 341;
	{8'd149,8'd193} : s = 342;
	{8'd149,8'd194} : s = 343;
	{8'd149,8'd195} : s = 344;
	{8'd149,8'd196} : s = 345;
	{8'd149,8'd197} : s = 346;
	{8'd149,8'd198} : s = 347;
	{8'd149,8'd199} : s = 348;
	{8'd149,8'd200} : s = 349;
	{8'd149,8'd201} : s = 350;
	{8'd149,8'd202} : s = 351;
	{8'd149,8'd203} : s = 352;
	{8'd149,8'd204} : s = 353;
	{8'd149,8'd205} : s = 354;
	{8'd149,8'd206} : s = 355;
	{8'd149,8'd207} : s = 356;
	{8'd149,8'd208} : s = 357;
	{8'd149,8'd209} : s = 358;
	{8'd149,8'd210} : s = 359;
	{8'd149,8'd211} : s = 360;
	{8'd149,8'd212} : s = 361;
	{8'd149,8'd213} : s = 362;
	{8'd149,8'd214} : s = 363;
	{8'd149,8'd215} : s = 364;
	{8'd149,8'd216} : s = 365;
	{8'd149,8'd217} : s = 366;
	{8'd149,8'd218} : s = 367;
	{8'd149,8'd219} : s = 368;
	{8'd149,8'd220} : s = 369;
	{8'd149,8'd221} : s = 370;
	{8'd149,8'd222} : s = 371;
	{8'd149,8'd223} : s = 372;
	{8'd149,8'd224} : s = 373;
	{8'd149,8'd225} : s = 374;
	{8'd149,8'd226} : s = 375;
	{8'd149,8'd227} : s = 376;
	{8'd149,8'd228} : s = 377;
	{8'd149,8'd229} : s = 378;
	{8'd149,8'd230} : s = 379;
	{8'd149,8'd231} : s = 380;
	{8'd149,8'd232} : s = 381;
	{8'd149,8'd233} : s = 382;
	{8'd149,8'd234} : s = 383;
	{8'd149,8'd235} : s = 384;
	{8'd149,8'd236} : s = 385;
	{8'd149,8'd237} : s = 386;
	{8'd149,8'd238} : s = 387;
	{8'd149,8'd239} : s = 388;
	{8'd149,8'd240} : s = 389;
	{8'd149,8'd241} : s = 390;
	{8'd149,8'd242} : s = 391;
	{8'd149,8'd243} : s = 392;
	{8'd149,8'd244} : s = 393;
	{8'd149,8'd245} : s = 394;
	{8'd149,8'd246} : s = 395;
	{8'd149,8'd247} : s = 396;
	{8'd149,8'd248} : s = 397;
	{8'd149,8'd249} : s = 398;
	{8'd149,8'd250} : s = 399;
	{8'd149,8'd251} : s = 400;
	{8'd149,8'd252} : s = 401;
	{8'd149,8'd253} : s = 402;
	{8'd149,8'd254} : s = 403;
	{8'd149,8'd255} : s = 404;
	{8'd150,8'd0} : s = 150;
	{8'd150,8'd1} : s = 151;
	{8'd150,8'd2} : s = 152;
	{8'd150,8'd3} : s = 153;
	{8'd150,8'd4} : s = 154;
	{8'd150,8'd5} : s = 155;
	{8'd150,8'd6} : s = 156;
	{8'd150,8'd7} : s = 157;
	{8'd150,8'd8} : s = 158;
	{8'd150,8'd9} : s = 159;
	{8'd150,8'd10} : s = 160;
	{8'd150,8'd11} : s = 161;
	{8'd150,8'd12} : s = 162;
	{8'd150,8'd13} : s = 163;
	{8'd150,8'd14} : s = 164;
	{8'd150,8'd15} : s = 165;
	{8'd150,8'd16} : s = 166;
	{8'd150,8'd17} : s = 167;
	{8'd150,8'd18} : s = 168;
	{8'd150,8'd19} : s = 169;
	{8'd150,8'd20} : s = 170;
	{8'd150,8'd21} : s = 171;
	{8'd150,8'd22} : s = 172;
	{8'd150,8'd23} : s = 173;
	{8'd150,8'd24} : s = 174;
	{8'd150,8'd25} : s = 175;
	{8'd150,8'd26} : s = 176;
	{8'd150,8'd27} : s = 177;
	{8'd150,8'd28} : s = 178;
	{8'd150,8'd29} : s = 179;
	{8'd150,8'd30} : s = 180;
	{8'd150,8'd31} : s = 181;
	{8'd150,8'd32} : s = 182;
	{8'd150,8'd33} : s = 183;
	{8'd150,8'd34} : s = 184;
	{8'd150,8'd35} : s = 185;
	{8'd150,8'd36} : s = 186;
	{8'd150,8'd37} : s = 187;
	{8'd150,8'd38} : s = 188;
	{8'd150,8'd39} : s = 189;
	{8'd150,8'd40} : s = 190;
	{8'd150,8'd41} : s = 191;
	{8'd150,8'd42} : s = 192;
	{8'd150,8'd43} : s = 193;
	{8'd150,8'd44} : s = 194;
	{8'd150,8'd45} : s = 195;
	{8'd150,8'd46} : s = 196;
	{8'd150,8'd47} : s = 197;
	{8'd150,8'd48} : s = 198;
	{8'd150,8'd49} : s = 199;
	{8'd150,8'd50} : s = 200;
	{8'd150,8'd51} : s = 201;
	{8'd150,8'd52} : s = 202;
	{8'd150,8'd53} : s = 203;
	{8'd150,8'd54} : s = 204;
	{8'd150,8'd55} : s = 205;
	{8'd150,8'd56} : s = 206;
	{8'd150,8'd57} : s = 207;
	{8'd150,8'd58} : s = 208;
	{8'd150,8'd59} : s = 209;
	{8'd150,8'd60} : s = 210;
	{8'd150,8'd61} : s = 211;
	{8'd150,8'd62} : s = 212;
	{8'd150,8'd63} : s = 213;
	{8'd150,8'd64} : s = 214;
	{8'd150,8'd65} : s = 215;
	{8'd150,8'd66} : s = 216;
	{8'd150,8'd67} : s = 217;
	{8'd150,8'd68} : s = 218;
	{8'd150,8'd69} : s = 219;
	{8'd150,8'd70} : s = 220;
	{8'd150,8'd71} : s = 221;
	{8'd150,8'd72} : s = 222;
	{8'd150,8'd73} : s = 223;
	{8'd150,8'd74} : s = 224;
	{8'd150,8'd75} : s = 225;
	{8'd150,8'd76} : s = 226;
	{8'd150,8'd77} : s = 227;
	{8'd150,8'd78} : s = 228;
	{8'd150,8'd79} : s = 229;
	{8'd150,8'd80} : s = 230;
	{8'd150,8'd81} : s = 231;
	{8'd150,8'd82} : s = 232;
	{8'd150,8'd83} : s = 233;
	{8'd150,8'd84} : s = 234;
	{8'd150,8'd85} : s = 235;
	{8'd150,8'd86} : s = 236;
	{8'd150,8'd87} : s = 237;
	{8'd150,8'd88} : s = 238;
	{8'd150,8'd89} : s = 239;
	{8'd150,8'd90} : s = 240;
	{8'd150,8'd91} : s = 241;
	{8'd150,8'd92} : s = 242;
	{8'd150,8'd93} : s = 243;
	{8'd150,8'd94} : s = 244;
	{8'd150,8'd95} : s = 245;
	{8'd150,8'd96} : s = 246;
	{8'd150,8'd97} : s = 247;
	{8'd150,8'd98} : s = 248;
	{8'd150,8'd99} : s = 249;
	{8'd150,8'd100} : s = 250;
	{8'd150,8'd101} : s = 251;
	{8'd150,8'd102} : s = 252;
	{8'd150,8'd103} : s = 253;
	{8'd150,8'd104} : s = 254;
	{8'd150,8'd105} : s = 255;
	{8'd150,8'd106} : s = 256;
	{8'd150,8'd107} : s = 257;
	{8'd150,8'd108} : s = 258;
	{8'd150,8'd109} : s = 259;
	{8'd150,8'd110} : s = 260;
	{8'd150,8'd111} : s = 261;
	{8'd150,8'd112} : s = 262;
	{8'd150,8'd113} : s = 263;
	{8'd150,8'd114} : s = 264;
	{8'd150,8'd115} : s = 265;
	{8'd150,8'd116} : s = 266;
	{8'd150,8'd117} : s = 267;
	{8'd150,8'd118} : s = 268;
	{8'd150,8'd119} : s = 269;
	{8'd150,8'd120} : s = 270;
	{8'd150,8'd121} : s = 271;
	{8'd150,8'd122} : s = 272;
	{8'd150,8'd123} : s = 273;
	{8'd150,8'd124} : s = 274;
	{8'd150,8'd125} : s = 275;
	{8'd150,8'd126} : s = 276;
	{8'd150,8'd127} : s = 277;
	{8'd150,8'd128} : s = 278;
	{8'd150,8'd129} : s = 279;
	{8'd150,8'd130} : s = 280;
	{8'd150,8'd131} : s = 281;
	{8'd150,8'd132} : s = 282;
	{8'd150,8'd133} : s = 283;
	{8'd150,8'd134} : s = 284;
	{8'd150,8'd135} : s = 285;
	{8'd150,8'd136} : s = 286;
	{8'd150,8'd137} : s = 287;
	{8'd150,8'd138} : s = 288;
	{8'd150,8'd139} : s = 289;
	{8'd150,8'd140} : s = 290;
	{8'd150,8'd141} : s = 291;
	{8'd150,8'd142} : s = 292;
	{8'd150,8'd143} : s = 293;
	{8'd150,8'd144} : s = 294;
	{8'd150,8'd145} : s = 295;
	{8'd150,8'd146} : s = 296;
	{8'd150,8'd147} : s = 297;
	{8'd150,8'd148} : s = 298;
	{8'd150,8'd149} : s = 299;
	{8'd150,8'd150} : s = 300;
	{8'd150,8'd151} : s = 301;
	{8'd150,8'd152} : s = 302;
	{8'd150,8'd153} : s = 303;
	{8'd150,8'd154} : s = 304;
	{8'd150,8'd155} : s = 305;
	{8'd150,8'd156} : s = 306;
	{8'd150,8'd157} : s = 307;
	{8'd150,8'd158} : s = 308;
	{8'd150,8'd159} : s = 309;
	{8'd150,8'd160} : s = 310;
	{8'd150,8'd161} : s = 311;
	{8'd150,8'd162} : s = 312;
	{8'd150,8'd163} : s = 313;
	{8'd150,8'd164} : s = 314;
	{8'd150,8'd165} : s = 315;
	{8'd150,8'd166} : s = 316;
	{8'd150,8'd167} : s = 317;
	{8'd150,8'd168} : s = 318;
	{8'd150,8'd169} : s = 319;
	{8'd150,8'd170} : s = 320;
	{8'd150,8'd171} : s = 321;
	{8'd150,8'd172} : s = 322;
	{8'd150,8'd173} : s = 323;
	{8'd150,8'd174} : s = 324;
	{8'd150,8'd175} : s = 325;
	{8'd150,8'd176} : s = 326;
	{8'd150,8'd177} : s = 327;
	{8'd150,8'd178} : s = 328;
	{8'd150,8'd179} : s = 329;
	{8'd150,8'd180} : s = 330;
	{8'd150,8'd181} : s = 331;
	{8'd150,8'd182} : s = 332;
	{8'd150,8'd183} : s = 333;
	{8'd150,8'd184} : s = 334;
	{8'd150,8'd185} : s = 335;
	{8'd150,8'd186} : s = 336;
	{8'd150,8'd187} : s = 337;
	{8'd150,8'd188} : s = 338;
	{8'd150,8'd189} : s = 339;
	{8'd150,8'd190} : s = 340;
	{8'd150,8'd191} : s = 341;
	{8'd150,8'd192} : s = 342;
	{8'd150,8'd193} : s = 343;
	{8'd150,8'd194} : s = 344;
	{8'd150,8'd195} : s = 345;
	{8'd150,8'd196} : s = 346;
	{8'd150,8'd197} : s = 347;
	{8'd150,8'd198} : s = 348;
	{8'd150,8'd199} : s = 349;
	{8'd150,8'd200} : s = 350;
	{8'd150,8'd201} : s = 351;
	{8'd150,8'd202} : s = 352;
	{8'd150,8'd203} : s = 353;
	{8'd150,8'd204} : s = 354;
	{8'd150,8'd205} : s = 355;
	{8'd150,8'd206} : s = 356;
	{8'd150,8'd207} : s = 357;
	{8'd150,8'd208} : s = 358;
	{8'd150,8'd209} : s = 359;
	{8'd150,8'd210} : s = 360;
	{8'd150,8'd211} : s = 361;
	{8'd150,8'd212} : s = 362;
	{8'd150,8'd213} : s = 363;
	{8'd150,8'd214} : s = 364;
	{8'd150,8'd215} : s = 365;
	{8'd150,8'd216} : s = 366;
	{8'd150,8'd217} : s = 367;
	{8'd150,8'd218} : s = 368;
	{8'd150,8'd219} : s = 369;
	{8'd150,8'd220} : s = 370;
	{8'd150,8'd221} : s = 371;
	{8'd150,8'd222} : s = 372;
	{8'd150,8'd223} : s = 373;
	{8'd150,8'd224} : s = 374;
	{8'd150,8'd225} : s = 375;
	{8'd150,8'd226} : s = 376;
	{8'd150,8'd227} : s = 377;
	{8'd150,8'd228} : s = 378;
	{8'd150,8'd229} : s = 379;
	{8'd150,8'd230} : s = 380;
	{8'd150,8'd231} : s = 381;
	{8'd150,8'd232} : s = 382;
	{8'd150,8'd233} : s = 383;
	{8'd150,8'd234} : s = 384;
	{8'd150,8'd235} : s = 385;
	{8'd150,8'd236} : s = 386;
	{8'd150,8'd237} : s = 387;
	{8'd150,8'd238} : s = 388;
	{8'd150,8'd239} : s = 389;
	{8'd150,8'd240} : s = 390;
	{8'd150,8'd241} : s = 391;
	{8'd150,8'd242} : s = 392;
	{8'd150,8'd243} : s = 393;
	{8'd150,8'd244} : s = 394;
	{8'd150,8'd245} : s = 395;
	{8'd150,8'd246} : s = 396;
	{8'd150,8'd247} : s = 397;
	{8'd150,8'd248} : s = 398;
	{8'd150,8'd249} : s = 399;
	{8'd150,8'd250} : s = 400;
	{8'd150,8'd251} : s = 401;
	{8'd150,8'd252} : s = 402;
	{8'd150,8'd253} : s = 403;
	{8'd150,8'd254} : s = 404;
	{8'd150,8'd255} : s = 405;
	{8'd151,8'd0} : s = 151;
	{8'd151,8'd1} : s = 152;
	{8'd151,8'd2} : s = 153;
	{8'd151,8'd3} : s = 154;
	{8'd151,8'd4} : s = 155;
	{8'd151,8'd5} : s = 156;
	{8'd151,8'd6} : s = 157;
	{8'd151,8'd7} : s = 158;
	{8'd151,8'd8} : s = 159;
	{8'd151,8'd9} : s = 160;
	{8'd151,8'd10} : s = 161;
	{8'd151,8'd11} : s = 162;
	{8'd151,8'd12} : s = 163;
	{8'd151,8'd13} : s = 164;
	{8'd151,8'd14} : s = 165;
	{8'd151,8'd15} : s = 166;
	{8'd151,8'd16} : s = 167;
	{8'd151,8'd17} : s = 168;
	{8'd151,8'd18} : s = 169;
	{8'd151,8'd19} : s = 170;
	{8'd151,8'd20} : s = 171;
	{8'd151,8'd21} : s = 172;
	{8'd151,8'd22} : s = 173;
	{8'd151,8'd23} : s = 174;
	{8'd151,8'd24} : s = 175;
	{8'd151,8'd25} : s = 176;
	{8'd151,8'd26} : s = 177;
	{8'd151,8'd27} : s = 178;
	{8'd151,8'd28} : s = 179;
	{8'd151,8'd29} : s = 180;
	{8'd151,8'd30} : s = 181;
	{8'd151,8'd31} : s = 182;
	{8'd151,8'd32} : s = 183;
	{8'd151,8'd33} : s = 184;
	{8'd151,8'd34} : s = 185;
	{8'd151,8'd35} : s = 186;
	{8'd151,8'd36} : s = 187;
	{8'd151,8'd37} : s = 188;
	{8'd151,8'd38} : s = 189;
	{8'd151,8'd39} : s = 190;
	{8'd151,8'd40} : s = 191;
	{8'd151,8'd41} : s = 192;
	{8'd151,8'd42} : s = 193;
	{8'd151,8'd43} : s = 194;
	{8'd151,8'd44} : s = 195;
	{8'd151,8'd45} : s = 196;
	{8'd151,8'd46} : s = 197;
	{8'd151,8'd47} : s = 198;
	{8'd151,8'd48} : s = 199;
	{8'd151,8'd49} : s = 200;
	{8'd151,8'd50} : s = 201;
	{8'd151,8'd51} : s = 202;
	{8'd151,8'd52} : s = 203;
	{8'd151,8'd53} : s = 204;
	{8'd151,8'd54} : s = 205;
	{8'd151,8'd55} : s = 206;
	{8'd151,8'd56} : s = 207;
	{8'd151,8'd57} : s = 208;
	{8'd151,8'd58} : s = 209;
	{8'd151,8'd59} : s = 210;
	{8'd151,8'd60} : s = 211;
	{8'd151,8'd61} : s = 212;
	{8'd151,8'd62} : s = 213;
	{8'd151,8'd63} : s = 214;
	{8'd151,8'd64} : s = 215;
	{8'd151,8'd65} : s = 216;
	{8'd151,8'd66} : s = 217;
	{8'd151,8'd67} : s = 218;
	{8'd151,8'd68} : s = 219;
	{8'd151,8'd69} : s = 220;
	{8'd151,8'd70} : s = 221;
	{8'd151,8'd71} : s = 222;
	{8'd151,8'd72} : s = 223;
	{8'd151,8'd73} : s = 224;
	{8'd151,8'd74} : s = 225;
	{8'd151,8'd75} : s = 226;
	{8'd151,8'd76} : s = 227;
	{8'd151,8'd77} : s = 228;
	{8'd151,8'd78} : s = 229;
	{8'd151,8'd79} : s = 230;
	{8'd151,8'd80} : s = 231;
	{8'd151,8'd81} : s = 232;
	{8'd151,8'd82} : s = 233;
	{8'd151,8'd83} : s = 234;
	{8'd151,8'd84} : s = 235;
	{8'd151,8'd85} : s = 236;
	{8'd151,8'd86} : s = 237;
	{8'd151,8'd87} : s = 238;
	{8'd151,8'd88} : s = 239;
	{8'd151,8'd89} : s = 240;
	{8'd151,8'd90} : s = 241;
	{8'd151,8'd91} : s = 242;
	{8'd151,8'd92} : s = 243;
	{8'd151,8'd93} : s = 244;
	{8'd151,8'd94} : s = 245;
	{8'd151,8'd95} : s = 246;
	{8'd151,8'd96} : s = 247;
	{8'd151,8'd97} : s = 248;
	{8'd151,8'd98} : s = 249;
	{8'd151,8'd99} : s = 250;
	{8'd151,8'd100} : s = 251;
	{8'd151,8'd101} : s = 252;
	{8'd151,8'd102} : s = 253;
	{8'd151,8'd103} : s = 254;
	{8'd151,8'd104} : s = 255;
	{8'd151,8'd105} : s = 256;
	{8'd151,8'd106} : s = 257;
	{8'd151,8'd107} : s = 258;
	{8'd151,8'd108} : s = 259;
	{8'd151,8'd109} : s = 260;
	{8'd151,8'd110} : s = 261;
	{8'd151,8'd111} : s = 262;
	{8'd151,8'd112} : s = 263;
	{8'd151,8'd113} : s = 264;
	{8'd151,8'd114} : s = 265;
	{8'd151,8'd115} : s = 266;
	{8'd151,8'd116} : s = 267;
	{8'd151,8'd117} : s = 268;
	{8'd151,8'd118} : s = 269;
	{8'd151,8'd119} : s = 270;
	{8'd151,8'd120} : s = 271;
	{8'd151,8'd121} : s = 272;
	{8'd151,8'd122} : s = 273;
	{8'd151,8'd123} : s = 274;
	{8'd151,8'd124} : s = 275;
	{8'd151,8'd125} : s = 276;
	{8'd151,8'd126} : s = 277;
	{8'd151,8'd127} : s = 278;
	{8'd151,8'd128} : s = 279;
	{8'd151,8'd129} : s = 280;
	{8'd151,8'd130} : s = 281;
	{8'd151,8'd131} : s = 282;
	{8'd151,8'd132} : s = 283;
	{8'd151,8'd133} : s = 284;
	{8'd151,8'd134} : s = 285;
	{8'd151,8'd135} : s = 286;
	{8'd151,8'd136} : s = 287;
	{8'd151,8'd137} : s = 288;
	{8'd151,8'd138} : s = 289;
	{8'd151,8'd139} : s = 290;
	{8'd151,8'd140} : s = 291;
	{8'd151,8'd141} : s = 292;
	{8'd151,8'd142} : s = 293;
	{8'd151,8'd143} : s = 294;
	{8'd151,8'd144} : s = 295;
	{8'd151,8'd145} : s = 296;
	{8'd151,8'd146} : s = 297;
	{8'd151,8'd147} : s = 298;
	{8'd151,8'd148} : s = 299;
	{8'd151,8'd149} : s = 300;
	{8'd151,8'd150} : s = 301;
	{8'd151,8'd151} : s = 302;
	{8'd151,8'd152} : s = 303;
	{8'd151,8'd153} : s = 304;
	{8'd151,8'd154} : s = 305;
	{8'd151,8'd155} : s = 306;
	{8'd151,8'd156} : s = 307;
	{8'd151,8'd157} : s = 308;
	{8'd151,8'd158} : s = 309;
	{8'd151,8'd159} : s = 310;
	{8'd151,8'd160} : s = 311;
	{8'd151,8'd161} : s = 312;
	{8'd151,8'd162} : s = 313;
	{8'd151,8'd163} : s = 314;
	{8'd151,8'd164} : s = 315;
	{8'd151,8'd165} : s = 316;
	{8'd151,8'd166} : s = 317;
	{8'd151,8'd167} : s = 318;
	{8'd151,8'd168} : s = 319;
	{8'd151,8'd169} : s = 320;
	{8'd151,8'd170} : s = 321;
	{8'd151,8'd171} : s = 322;
	{8'd151,8'd172} : s = 323;
	{8'd151,8'd173} : s = 324;
	{8'd151,8'd174} : s = 325;
	{8'd151,8'd175} : s = 326;
	{8'd151,8'd176} : s = 327;
	{8'd151,8'd177} : s = 328;
	{8'd151,8'd178} : s = 329;
	{8'd151,8'd179} : s = 330;
	{8'd151,8'd180} : s = 331;
	{8'd151,8'd181} : s = 332;
	{8'd151,8'd182} : s = 333;
	{8'd151,8'd183} : s = 334;
	{8'd151,8'd184} : s = 335;
	{8'd151,8'd185} : s = 336;
	{8'd151,8'd186} : s = 337;
	{8'd151,8'd187} : s = 338;
	{8'd151,8'd188} : s = 339;
	{8'd151,8'd189} : s = 340;
	{8'd151,8'd190} : s = 341;
	{8'd151,8'd191} : s = 342;
	{8'd151,8'd192} : s = 343;
	{8'd151,8'd193} : s = 344;
	{8'd151,8'd194} : s = 345;
	{8'd151,8'd195} : s = 346;
	{8'd151,8'd196} : s = 347;
	{8'd151,8'd197} : s = 348;
	{8'd151,8'd198} : s = 349;
	{8'd151,8'd199} : s = 350;
	{8'd151,8'd200} : s = 351;
	{8'd151,8'd201} : s = 352;
	{8'd151,8'd202} : s = 353;
	{8'd151,8'd203} : s = 354;
	{8'd151,8'd204} : s = 355;
	{8'd151,8'd205} : s = 356;
	{8'd151,8'd206} : s = 357;
	{8'd151,8'd207} : s = 358;
	{8'd151,8'd208} : s = 359;
	{8'd151,8'd209} : s = 360;
	{8'd151,8'd210} : s = 361;
	{8'd151,8'd211} : s = 362;
	{8'd151,8'd212} : s = 363;
	{8'd151,8'd213} : s = 364;
	{8'd151,8'd214} : s = 365;
	{8'd151,8'd215} : s = 366;
	{8'd151,8'd216} : s = 367;
	{8'd151,8'd217} : s = 368;
	{8'd151,8'd218} : s = 369;
	{8'd151,8'd219} : s = 370;
	{8'd151,8'd220} : s = 371;
	{8'd151,8'd221} : s = 372;
	{8'd151,8'd222} : s = 373;
	{8'd151,8'd223} : s = 374;
	{8'd151,8'd224} : s = 375;
	{8'd151,8'd225} : s = 376;
	{8'd151,8'd226} : s = 377;
	{8'd151,8'd227} : s = 378;
	{8'd151,8'd228} : s = 379;
	{8'd151,8'd229} : s = 380;
	{8'd151,8'd230} : s = 381;
	{8'd151,8'd231} : s = 382;
	{8'd151,8'd232} : s = 383;
	{8'd151,8'd233} : s = 384;
	{8'd151,8'd234} : s = 385;
	{8'd151,8'd235} : s = 386;
	{8'd151,8'd236} : s = 387;
	{8'd151,8'd237} : s = 388;
	{8'd151,8'd238} : s = 389;
	{8'd151,8'd239} : s = 390;
	{8'd151,8'd240} : s = 391;
	{8'd151,8'd241} : s = 392;
	{8'd151,8'd242} : s = 393;
	{8'd151,8'd243} : s = 394;
	{8'd151,8'd244} : s = 395;
	{8'd151,8'd245} : s = 396;
	{8'd151,8'd246} : s = 397;
	{8'd151,8'd247} : s = 398;
	{8'd151,8'd248} : s = 399;
	{8'd151,8'd249} : s = 400;
	{8'd151,8'd250} : s = 401;
	{8'd151,8'd251} : s = 402;
	{8'd151,8'd252} : s = 403;
	{8'd151,8'd253} : s = 404;
	{8'd151,8'd254} : s = 405;
	{8'd151,8'd255} : s = 406;
	{8'd152,8'd0} : s = 152;
	{8'd152,8'd1} : s = 153;
	{8'd152,8'd2} : s = 154;
	{8'd152,8'd3} : s = 155;
	{8'd152,8'd4} : s = 156;
	{8'd152,8'd5} : s = 157;
	{8'd152,8'd6} : s = 158;
	{8'd152,8'd7} : s = 159;
	{8'd152,8'd8} : s = 160;
	{8'd152,8'd9} : s = 161;
	{8'd152,8'd10} : s = 162;
	{8'd152,8'd11} : s = 163;
	{8'd152,8'd12} : s = 164;
	{8'd152,8'd13} : s = 165;
	{8'd152,8'd14} : s = 166;
	{8'd152,8'd15} : s = 167;
	{8'd152,8'd16} : s = 168;
	{8'd152,8'd17} : s = 169;
	{8'd152,8'd18} : s = 170;
	{8'd152,8'd19} : s = 171;
	{8'd152,8'd20} : s = 172;
	{8'd152,8'd21} : s = 173;
	{8'd152,8'd22} : s = 174;
	{8'd152,8'd23} : s = 175;
	{8'd152,8'd24} : s = 176;
	{8'd152,8'd25} : s = 177;
	{8'd152,8'd26} : s = 178;
	{8'd152,8'd27} : s = 179;
	{8'd152,8'd28} : s = 180;
	{8'd152,8'd29} : s = 181;
	{8'd152,8'd30} : s = 182;
	{8'd152,8'd31} : s = 183;
	{8'd152,8'd32} : s = 184;
	{8'd152,8'd33} : s = 185;
	{8'd152,8'd34} : s = 186;
	{8'd152,8'd35} : s = 187;
	{8'd152,8'd36} : s = 188;
	{8'd152,8'd37} : s = 189;
	{8'd152,8'd38} : s = 190;
	{8'd152,8'd39} : s = 191;
	{8'd152,8'd40} : s = 192;
	{8'd152,8'd41} : s = 193;
	{8'd152,8'd42} : s = 194;
	{8'd152,8'd43} : s = 195;
	{8'd152,8'd44} : s = 196;
	{8'd152,8'd45} : s = 197;
	{8'd152,8'd46} : s = 198;
	{8'd152,8'd47} : s = 199;
	{8'd152,8'd48} : s = 200;
	{8'd152,8'd49} : s = 201;
	{8'd152,8'd50} : s = 202;
	{8'd152,8'd51} : s = 203;
	{8'd152,8'd52} : s = 204;
	{8'd152,8'd53} : s = 205;
	{8'd152,8'd54} : s = 206;
	{8'd152,8'd55} : s = 207;
	{8'd152,8'd56} : s = 208;
	{8'd152,8'd57} : s = 209;
	{8'd152,8'd58} : s = 210;
	{8'd152,8'd59} : s = 211;
	{8'd152,8'd60} : s = 212;
	{8'd152,8'd61} : s = 213;
	{8'd152,8'd62} : s = 214;
	{8'd152,8'd63} : s = 215;
	{8'd152,8'd64} : s = 216;
	{8'd152,8'd65} : s = 217;
	{8'd152,8'd66} : s = 218;
	{8'd152,8'd67} : s = 219;
	{8'd152,8'd68} : s = 220;
	{8'd152,8'd69} : s = 221;
	{8'd152,8'd70} : s = 222;
	{8'd152,8'd71} : s = 223;
	{8'd152,8'd72} : s = 224;
	{8'd152,8'd73} : s = 225;
	{8'd152,8'd74} : s = 226;
	{8'd152,8'd75} : s = 227;
	{8'd152,8'd76} : s = 228;
	{8'd152,8'd77} : s = 229;
	{8'd152,8'd78} : s = 230;
	{8'd152,8'd79} : s = 231;
	{8'd152,8'd80} : s = 232;
	{8'd152,8'd81} : s = 233;
	{8'd152,8'd82} : s = 234;
	{8'd152,8'd83} : s = 235;
	{8'd152,8'd84} : s = 236;
	{8'd152,8'd85} : s = 237;
	{8'd152,8'd86} : s = 238;
	{8'd152,8'd87} : s = 239;
	{8'd152,8'd88} : s = 240;
	{8'd152,8'd89} : s = 241;
	{8'd152,8'd90} : s = 242;
	{8'd152,8'd91} : s = 243;
	{8'd152,8'd92} : s = 244;
	{8'd152,8'd93} : s = 245;
	{8'd152,8'd94} : s = 246;
	{8'd152,8'd95} : s = 247;
	{8'd152,8'd96} : s = 248;
	{8'd152,8'd97} : s = 249;
	{8'd152,8'd98} : s = 250;
	{8'd152,8'd99} : s = 251;
	{8'd152,8'd100} : s = 252;
	{8'd152,8'd101} : s = 253;
	{8'd152,8'd102} : s = 254;
	{8'd152,8'd103} : s = 255;
	{8'd152,8'd104} : s = 256;
	{8'd152,8'd105} : s = 257;
	{8'd152,8'd106} : s = 258;
	{8'd152,8'd107} : s = 259;
	{8'd152,8'd108} : s = 260;
	{8'd152,8'd109} : s = 261;
	{8'd152,8'd110} : s = 262;
	{8'd152,8'd111} : s = 263;
	{8'd152,8'd112} : s = 264;
	{8'd152,8'd113} : s = 265;
	{8'd152,8'd114} : s = 266;
	{8'd152,8'd115} : s = 267;
	{8'd152,8'd116} : s = 268;
	{8'd152,8'd117} : s = 269;
	{8'd152,8'd118} : s = 270;
	{8'd152,8'd119} : s = 271;
	{8'd152,8'd120} : s = 272;
	{8'd152,8'd121} : s = 273;
	{8'd152,8'd122} : s = 274;
	{8'd152,8'd123} : s = 275;
	{8'd152,8'd124} : s = 276;
	{8'd152,8'd125} : s = 277;
	{8'd152,8'd126} : s = 278;
	{8'd152,8'd127} : s = 279;
	{8'd152,8'd128} : s = 280;
	{8'd152,8'd129} : s = 281;
	{8'd152,8'd130} : s = 282;
	{8'd152,8'd131} : s = 283;
	{8'd152,8'd132} : s = 284;
	{8'd152,8'd133} : s = 285;
	{8'd152,8'd134} : s = 286;
	{8'd152,8'd135} : s = 287;
	{8'd152,8'd136} : s = 288;
	{8'd152,8'd137} : s = 289;
	{8'd152,8'd138} : s = 290;
	{8'd152,8'd139} : s = 291;
	{8'd152,8'd140} : s = 292;
	{8'd152,8'd141} : s = 293;
	{8'd152,8'd142} : s = 294;
	{8'd152,8'd143} : s = 295;
	{8'd152,8'd144} : s = 296;
	{8'd152,8'd145} : s = 297;
	{8'd152,8'd146} : s = 298;
	{8'd152,8'd147} : s = 299;
	{8'd152,8'd148} : s = 300;
	{8'd152,8'd149} : s = 301;
	{8'd152,8'd150} : s = 302;
	{8'd152,8'd151} : s = 303;
	{8'd152,8'd152} : s = 304;
	{8'd152,8'd153} : s = 305;
	{8'd152,8'd154} : s = 306;
	{8'd152,8'd155} : s = 307;
	{8'd152,8'd156} : s = 308;
	{8'd152,8'd157} : s = 309;
	{8'd152,8'd158} : s = 310;
	{8'd152,8'd159} : s = 311;
	{8'd152,8'd160} : s = 312;
	{8'd152,8'd161} : s = 313;
	{8'd152,8'd162} : s = 314;
	{8'd152,8'd163} : s = 315;
	{8'd152,8'd164} : s = 316;
	{8'd152,8'd165} : s = 317;
	{8'd152,8'd166} : s = 318;
	{8'd152,8'd167} : s = 319;
	{8'd152,8'd168} : s = 320;
	{8'd152,8'd169} : s = 321;
	{8'd152,8'd170} : s = 322;
	{8'd152,8'd171} : s = 323;
	{8'd152,8'd172} : s = 324;
	{8'd152,8'd173} : s = 325;
	{8'd152,8'd174} : s = 326;
	{8'd152,8'd175} : s = 327;
	{8'd152,8'd176} : s = 328;
	{8'd152,8'd177} : s = 329;
	{8'd152,8'd178} : s = 330;
	{8'd152,8'd179} : s = 331;
	{8'd152,8'd180} : s = 332;
	{8'd152,8'd181} : s = 333;
	{8'd152,8'd182} : s = 334;
	{8'd152,8'd183} : s = 335;
	{8'd152,8'd184} : s = 336;
	{8'd152,8'd185} : s = 337;
	{8'd152,8'd186} : s = 338;
	{8'd152,8'd187} : s = 339;
	{8'd152,8'd188} : s = 340;
	{8'd152,8'd189} : s = 341;
	{8'd152,8'd190} : s = 342;
	{8'd152,8'd191} : s = 343;
	{8'd152,8'd192} : s = 344;
	{8'd152,8'd193} : s = 345;
	{8'd152,8'd194} : s = 346;
	{8'd152,8'd195} : s = 347;
	{8'd152,8'd196} : s = 348;
	{8'd152,8'd197} : s = 349;
	{8'd152,8'd198} : s = 350;
	{8'd152,8'd199} : s = 351;
	{8'd152,8'd200} : s = 352;
	{8'd152,8'd201} : s = 353;
	{8'd152,8'd202} : s = 354;
	{8'd152,8'd203} : s = 355;
	{8'd152,8'd204} : s = 356;
	{8'd152,8'd205} : s = 357;
	{8'd152,8'd206} : s = 358;
	{8'd152,8'd207} : s = 359;
	{8'd152,8'd208} : s = 360;
	{8'd152,8'd209} : s = 361;
	{8'd152,8'd210} : s = 362;
	{8'd152,8'd211} : s = 363;
	{8'd152,8'd212} : s = 364;
	{8'd152,8'd213} : s = 365;
	{8'd152,8'd214} : s = 366;
	{8'd152,8'd215} : s = 367;
	{8'd152,8'd216} : s = 368;
	{8'd152,8'd217} : s = 369;
	{8'd152,8'd218} : s = 370;
	{8'd152,8'd219} : s = 371;
	{8'd152,8'd220} : s = 372;
	{8'd152,8'd221} : s = 373;
	{8'd152,8'd222} : s = 374;
	{8'd152,8'd223} : s = 375;
	{8'd152,8'd224} : s = 376;
	{8'd152,8'd225} : s = 377;
	{8'd152,8'd226} : s = 378;
	{8'd152,8'd227} : s = 379;
	{8'd152,8'd228} : s = 380;
	{8'd152,8'd229} : s = 381;
	{8'd152,8'd230} : s = 382;
	{8'd152,8'd231} : s = 383;
	{8'd152,8'd232} : s = 384;
	{8'd152,8'd233} : s = 385;
	{8'd152,8'd234} : s = 386;
	{8'd152,8'd235} : s = 387;
	{8'd152,8'd236} : s = 388;
	{8'd152,8'd237} : s = 389;
	{8'd152,8'd238} : s = 390;
	{8'd152,8'd239} : s = 391;
	{8'd152,8'd240} : s = 392;
	{8'd152,8'd241} : s = 393;
	{8'd152,8'd242} : s = 394;
	{8'd152,8'd243} : s = 395;
	{8'd152,8'd244} : s = 396;
	{8'd152,8'd245} : s = 397;
	{8'd152,8'd246} : s = 398;
	{8'd152,8'd247} : s = 399;
	{8'd152,8'd248} : s = 400;
	{8'd152,8'd249} : s = 401;
	{8'd152,8'd250} : s = 402;
	{8'd152,8'd251} : s = 403;
	{8'd152,8'd252} : s = 404;
	{8'd152,8'd253} : s = 405;
	{8'd152,8'd254} : s = 406;
	{8'd152,8'd255} : s = 407;
	{8'd153,8'd0} : s = 153;
	{8'd153,8'd1} : s = 154;
	{8'd153,8'd2} : s = 155;
	{8'd153,8'd3} : s = 156;
	{8'd153,8'd4} : s = 157;
	{8'd153,8'd5} : s = 158;
	{8'd153,8'd6} : s = 159;
	{8'd153,8'd7} : s = 160;
	{8'd153,8'd8} : s = 161;
	{8'd153,8'd9} : s = 162;
	{8'd153,8'd10} : s = 163;
	{8'd153,8'd11} : s = 164;
	{8'd153,8'd12} : s = 165;
	{8'd153,8'd13} : s = 166;
	{8'd153,8'd14} : s = 167;
	{8'd153,8'd15} : s = 168;
	{8'd153,8'd16} : s = 169;
	{8'd153,8'd17} : s = 170;
	{8'd153,8'd18} : s = 171;
	{8'd153,8'd19} : s = 172;
	{8'd153,8'd20} : s = 173;
	{8'd153,8'd21} : s = 174;
	{8'd153,8'd22} : s = 175;
	{8'd153,8'd23} : s = 176;
	{8'd153,8'd24} : s = 177;
	{8'd153,8'd25} : s = 178;
	{8'd153,8'd26} : s = 179;
	{8'd153,8'd27} : s = 180;
	{8'd153,8'd28} : s = 181;
	{8'd153,8'd29} : s = 182;
	{8'd153,8'd30} : s = 183;
	{8'd153,8'd31} : s = 184;
	{8'd153,8'd32} : s = 185;
	{8'd153,8'd33} : s = 186;
	{8'd153,8'd34} : s = 187;
	{8'd153,8'd35} : s = 188;
	{8'd153,8'd36} : s = 189;
	{8'd153,8'd37} : s = 190;
	{8'd153,8'd38} : s = 191;
	{8'd153,8'd39} : s = 192;
	{8'd153,8'd40} : s = 193;
	{8'd153,8'd41} : s = 194;
	{8'd153,8'd42} : s = 195;
	{8'd153,8'd43} : s = 196;
	{8'd153,8'd44} : s = 197;
	{8'd153,8'd45} : s = 198;
	{8'd153,8'd46} : s = 199;
	{8'd153,8'd47} : s = 200;
	{8'd153,8'd48} : s = 201;
	{8'd153,8'd49} : s = 202;
	{8'd153,8'd50} : s = 203;
	{8'd153,8'd51} : s = 204;
	{8'd153,8'd52} : s = 205;
	{8'd153,8'd53} : s = 206;
	{8'd153,8'd54} : s = 207;
	{8'd153,8'd55} : s = 208;
	{8'd153,8'd56} : s = 209;
	{8'd153,8'd57} : s = 210;
	{8'd153,8'd58} : s = 211;
	{8'd153,8'd59} : s = 212;
	{8'd153,8'd60} : s = 213;
	{8'd153,8'd61} : s = 214;
	{8'd153,8'd62} : s = 215;
	{8'd153,8'd63} : s = 216;
	{8'd153,8'd64} : s = 217;
	{8'd153,8'd65} : s = 218;
	{8'd153,8'd66} : s = 219;
	{8'd153,8'd67} : s = 220;
	{8'd153,8'd68} : s = 221;
	{8'd153,8'd69} : s = 222;
	{8'd153,8'd70} : s = 223;
	{8'd153,8'd71} : s = 224;
	{8'd153,8'd72} : s = 225;
	{8'd153,8'd73} : s = 226;
	{8'd153,8'd74} : s = 227;
	{8'd153,8'd75} : s = 228;
	{8'd153,8'd76} : s = 229;
	{8'd153,8'd77} : s = 230;
	{8'd153,8'd78} : s = 231;
	{8'd153,8'd79} : s = 232;
	{8'd153,8'd80} : s = 233;
	{8'd153,8'd81} : s = 234;
	{8'd153,8'd82} : s = 235;
	{8'd153,8'd83} : s = 236;
	{8'd153,8'd84} : s = 237;
	{8'd153,8'd85} : s = 238;
	{8'd153,8'd86} : s = 239;
	{8'd153,8'd87} : s = 240;
	{8'd153,8'd88} : s = 241;
	{8'd153,8'd89} : s = 242;
	{8'd153,8'd90} : s = 243;
	{8'd153,8'd91} : s = 244;
	{8'd153,8'd92} : s = 245;
	{8'd153,8'd93} : s = 246;
	{8'd153,8'd94} : s = 247;
	{8'd153,8'd95} : s = 248;
	{8'd153,8'd96} : s = 249;
	{8'd153,8'd97} : s = 250;
	{8'd153,8'd98} : s = 251;
	{8'd153,8'd99} : s = 252;
	{8'd153,8'd100} : s = 253;
	{8'd153,8'd101} : s = 254;
	{8'd153,8'd102} : s = 255;
	{8'd153,8'd103} : s = 256;
	{8'd153,8'd104} : s = 257;
	{8'd153,8'd105} : s = 258;
	{8'd153,8'd106} : s = 259;
	{8'd153,8'd107} : s = 260;
	{8'd153,8'd108} : s = 261;
	{8'd153,8'd109} : s = 262;
	{8'd153,8'd110} : s = 263;
	{8'd153,8'd111} : s = 264;
	{8'd153,8'd112} : s = 265;
	{8'd153,8'd113} : s = 266;
	{8'd153,8'd114} : s = 267;
	{8'd153,8'd115} : s = 268;
	{8'd153,8'd116} : s = 269;
	{8'd153,8'd117} : s = 270;
	{8'd153,8'd118} : s = 271;
	{8'd153,8'd119} : s = 272;
	{8'd153,8'd120} : s = 273;
	{8'd153,8'd121} : s = 274;
	{8'd153,8'd122} : s = 275;
	{8'd153,8'd123} : s = 276;
	{8'd153,8'd124} : s = 277;
	{8'd153,8'd125} : s = 278;
	{8'd153,8'd126} : s = 279;
	{8'd153,8'd127} : s = 280;
	{8'd153,8'd128} : s = 281;
	{8'd153,8'd129} : s = 282;
	{8'd153,8'd130} : s = 283;
	{8'd153,8'd131} : s = 284;
	{8'd153,8'd132} : s = 285;
	{8'd153,8'd133} : s = 286;
	{8'd153,8'd134} : s = 287;
	{8'd153,8'd135} : s = 288;
	{8'd153,8'd136} : s = 289;
	{8'd153,8'd137} : s = 290;
	{8'd153,8'd138} : s = 291;
	{8'd153,8'd139} : s = 292;
	{8'd153,8'd140} : s = 293;
	{8'd153,8'd141} : s = 294;
	{8'd153,8'd142} : s = 295;
	{8'd153,8'd143} : s = 296;
	{8'd153,8'd144} : s = 297;
	{8'd153,8'd145} : s = 298;
	{8'd153,8'd146} : s = 299;
	{8'd153,8'd147} : s = 300;
	{8'd153,8'd148} : s = 301;
	{8'd153,8'd149} : s = 302;
	{8'd153,8'd150} : s = 303;
	{8'd153,8'd151} : s = 304;
	{8'd153,8'd152} : s = 305;
	{8'd153,8'd153} : s = 306;
	{8'd153,8'd154} : s = 307;
	{8'd153,8'd155} : s = 308;
	{8'd153,8'd156} : s = 309;
	{8'd153,8'd157} : s = 310;
	{8'd153,8'd158} : s = 311;
	{8'd153,8'd159} : s = 312;
	{8'd153,8'd160} : s = 313;
	{8'd153,8'd161} : s = 314;
	{8'd153,8'd162} : s = 315;
	{8'd153,8'd163} : s = 316;
	{8'd153,8'd164} : s = 317;
	{8'd153,8'd165} : s = 318;
	{8'd153,8'd166} : s = 319;
	{8'd153,8'd167} : s = 320;
	{8'd153,8'd168} : s = 321;
	{8'd153,8'd169} : s = 322;
	{8'd153,8'd170} : s = 323;
	{8'd153,8'd171} : s = 324;
	{8'd153,8'd172} : s = 325;
	{8'd153,8'd173} : s = 326;
	{8'd153,8'd174} : s = 327;
	{8'd153,8'd175} : s = 328;
	{8'd153,8'd176} : s = 329;
	{8'd153,8'd177} : s = 330;
	{8'd153,8'd178} : s = 331;
	{8'd153,8'd179} : s = 332;
	{8'd153,8'd180} : s = 333;
	{8'd153,8'd181} : s = 334;
	{8'd153,8'd182} : s = 335;
	{8'd153,8'd183} : s = 336;
	{8'd153,8'd184} : s = 337;
	{8'd153,8'd185} : s = 338;
	{8'd153,8'd186} : s = 339;
	{8'd153,8'd187} : s = 340;
	{8'd153,8'd188} : s = 341;
	{8'd153,8'd189} : s = 342;
	{8'd153,8'd190} : s = 343;
	{8'd153,8'd191} : s = 344;
	{8'd153,8'd192} : s = 345;
	{8'd153,8'd193} : s = 346;
	{8'd153,8'd194} : s = 347;
	{8'd153,8'd195} : s = 348;
	{8'd153,8'd196} : s = 349;
	{8'd153,8'd197} : s = 350;
	{8'd153,8'd198} : s = 351;
	{8'd153,8'd199} : s = 352;
	{8'd153,8'd200} : s = 353;
	{8'd153,8'd201} : s = 354;
	{8'd153,8'd202} : s = 355;
	{8'd153,8'd203} : s = 356;
	{8'd153,8'd204} : s = 357;
	{8'd153,8'd205} : s = 358;
	{8'd153,8'd206} : s = 359;
	{8'd153,8'd207} : s = 360;
	{8'd153,8'd208} : s = 361;
	{8'd153,8'd209} : s = 362;
	{8'd153,8'd210} : s = 363;
	{8'd153,8'd211} : s = 364;
	{8'd153,8'd212} : s = 365;
	{8'd153,8'd213} : s = 366;
	{8'd153,8'd214} : s = 367;
	{8'd153,8'd215} : s = 368;
	{8'd153,8'd216} : s = 369;
	{8'd153,8'd217} : s = 370;
	{8'd153,8'd218} : s = 371;
	{8'd153,8'd219} : s = 372;
	{8'd153,8'd220} : s = 373;
	{8'd153,8'd221} : s = 374;
	{8'd153,8'd222} : s = 375;
	{8'd153,8'd223} : s = 376;
	{8'd153,8'd224} : s = 377;
	{8'd153,8'd225} : s = 378;
	{8'd153,8'd226} : s = 379;
	{8'd153,8'd227} : s = 380;
	{8'd153,8'd228} : s = 381;
	{8'd153,8'd229} : s = 382;
	{8'd153,8'd230} : s = 383;
	{8'd153,8'd231} : s = 384;
	{8'd153,8'd232} : s = 385;
	{8'd153,8'd233} : s = 386;
	{8'd153,8'd234} : s = 387;
	{8'd153,8'd235} : s = 388;
	{8'd153,8'd236} : s = 389;
	{8'd153,8'd237} : s = 390;
	{8'd153,8'd238} : s = 391;
	{8'd153,8'd239} : s = 392;
	{8'd153,8'd240} : s = 393;
	{8'd153,8'd241} : s = 394;
	{8'd153,8'd242} : s = 395;
	{8'd153,8'd243} : s = 396;
	{8'd153,8'd244} : s = 397;
	{8'd153,8'd245} : s = 398;
	{8'd153,8'd246} : s = 399;
	{8'd153,8'd247} : s = 400;
	{8'd153,8'd248} : s = 401;
	{8'd153,8'd249} : s = 402;
	{8'd153,8'd250} : s = 403;
	{8'd153,8'd251} : s = 404;
	{8'd153,8'd252} : s = 405;
	{8'd153,8'd253} : s = 406;
	{8'd153,8'd254} : s = 407;
	{8'd153,8'd255} : s = 408;
	{8'd154,8'd0} : s = 154;
	{8'd154,8'd1} : s = 155;
	{8'd154,8'd2} : s = 156;
	{8'd154,8'd3} : s = 157;
	{8'd154,8'd4} : s = 158;
	{8'd154,8'd5} : s = 159;
	{8'd154,8'd6} : s = 160;
	{8'd154,8'd7} : s = 161;
	{8'd154,8'd8} : s = 162;
	{8'd154,8'd9} : s = 163;
	{8'd154,8'd10} : s = 164;
	{8'd154,8'd11} : s = 165;
	{8'd154,8'd12} : s = 166;
	{8'd154,8'd13} : s = 167;
	{8'd154,8'd14} : s = 168;
	{8'd154,8'd15} : s = 169;
	{8'd154,8'd16} : s = 170;
	{8'd154,8'd17} : s = 171;
	{8'd154,8'd18} : s = 172;
	{8'd154,8'd19} : s = 173;
	{8'd154,8'd20} : s = 174;
	{8'd154,8'd21} : s = 175;
	{8'd154,8'd22} : s = 176;
	{8'd154,8'd23} : s = 177;
	{8'd154,8'd24} : s = 178;
	{8'd154,8'd25} : s = 179;
	{8'd154,8'd26} : s = 180;
	{8'd154,8'd27} : s = 181;
	{8'd154,8'd28} : s = 182;
	{8'd154,8'd29} : s = 183;
	{8'd154,8'd30} : s = 184;
	{8'd154,8'd31} : s = 185;
	{8'd154,8'd32} : s = 186;
	{8'd154,8'd33} : s = 187;
	{8'd154,8'd34} : s = 188;
	{8'd154,8'd35} : s = 189;
	{8'd154,8'd36} : s = 190;
	{8'd154,8'd37} : s = 191;
	{8'd154,8'd38} : s = 192;
	{8'd154,8'd39} : s = 193;
	{8'd154,8'd40} : s = 194;
	{8'd154,8'd41} : s = 195;
	{8'd154,8'd42} : s = 196;
	{8'd154,8'd43} : s = 197;
	{8'd154,8'd44} : s = 198;
	{8'd154,8'd45} : s = 199;
	{8'd154,8'd46} : s = 200;
	{8'd154,8'd47} : s = 201;
	{8'd154,8'd48} : s = 202;
	{8'd154,8'd49} : s = 203;
	{8'd154,8'd50} : s = 204;
	{8'd154,8'd51} : s = 205;
	{8'd154,8'd52} : s = 206;
	{8'd154,8'd53} : s = 207;
	{8'd154,8'd54} : s = 208;
	{8'd154,8'd55} : s = 209;
	{8'd154,8'd56} : s = 210;
	{8'd154,8'd57} : s = 211;
	{8'd154,8'd58} : s = 212;
	{8'd154,8'd59} : s = 213;
	{8'd154,8'd60} : s = 214;
	{8'd154,8'd61} : s = 215;
	{8'd154,8'd62} : s = 216;
	{8'd154,8'd63} : s = 217;
	{8'd154,8'd64} : s = 218;
	{8'd154,8'd65} : s = 219;
	{8'd154,8'd66} : s = 220;
	{8'd154,8'd67} : s = 221;
	{8'd154,8'd68} : s = 222;
	{8'd154,8'd69} : s = 223;
	{8'd154,8'd70} : s = 224;
	{8'd154,8'd71} : s = 225;
	{8'd154,8'd72} : s = 226;
	{8'd154,8'd73} : s = 227;
	{8'd154,8'd74} : s = 228;
	{8'd154,8'd75} : s = 229;
	{8'd154,8'd76} : s = 230;
	{8'd154,8'd77} : s = 231;
	{8'd154,8'd78} : s = 232;
	{8'd154,8'd79} : s = 233;
	{8'd154,8'd80} : s = 234;
	{8'd154,8'd81} : s = 235;
	{8'd154,8'd82} : s = 236;
	{8'd154,8'd83} : s = 237;
	{8'd154,8'd84} : s = 238;
	{8'd154,8'd85} : s = 239;
	{8'd154,8'd86} : s = 240;
	{8'd154,8'd87} : s = 241;
	{8'd154,8'd88} : s = 242;
	{8'd154,8'd89} : s = 243;
	{8'd154,8'd90} : s = 244;
	{8'd154,8'd91} : s = 245;
	{8'd154,8'd92} : s = 246;
	{8'd154,8'd93} : s = 247;
	{8'd154,8'd94} : s = 248;
	{8'd154,8'd95} : s = 249;
	{8'd154,8'd96} : s = 250;
	{8'd154,8'd97} : s = 251;
	{8'd154,8'd98} : s = 252;
	{8'd154,8'd99} : s = 253;
	{8'd154,8'd100} : s = 254;
	{8'd154,8'd101} : s = 255;
	{8'd154,8'd102} : s = 256;
	{8'd154,8'd103} : s = 257;
	{8'd154,8'd104} : s = 258;
	{8'd154,8'd105} : s = 259;
	{8'd154,8'd106} : s = 260;
	{8'd154,8'd107} : s = 261;
	{8'd154,8'd108} : s = 262;
	{8'd154,8'd109} : s = 263;
	{8'd154,8'd110} : s = 264;
	{8'd154,8'd111} : s = 265;
	{8'd154,8'd112} : s = 266;
	{8'd154,8'd113} : s = 267;
	{8'd154,8'd114} : s = 268;
	{8'd154,8'd115} : s = 269;
	{8'd154,8'd116} : s = 270;
	{8'd154,8'd117} : s = 271;
	{8'd154,8'd118} : s = 272;
	{8'd154,8'd119} : s = 273;
	{8'd154,8'd120} : s = 274;
	{8'd154,8'd121} : s = 275;
	{8'd154,8'd122} : s = 276;
	{8'd154,8'd123} : s = 277;
	{8'd154,8'd124} : s = 278;
	{8'd154,8'd125} : s = 279;
	{8'd154,8'd126} : s = 280;
	{8'd154,8'd127} : s = 281;
	{8'd154,8'd128} : s = 282;
	{8'd154,8'd129} : s = 283;
	{8'd154,8'd130} : s = 284;
	{8'd154,8'd131} : s = 285;
	{8'd154,8'd132} : s = 286;
	{8'd154,8'd133} : s = 287;
	{8'd154,8'd134} : s = 288;
	{8'd154,8'd135} : s = 289;
	{8'd154,8'd136} : s = 290;
	{8'd154,8'd137} : s = 291;
	{8'd154,8'd138} : s = 292;
	{8'd154,8'd139} : s = 293;
	{8'd154,8'd140} : s = 294;
	{8'd154,8'd141} : s = 295;
	{8'd154,8'd142} : s = 296;
	{8'd154,8'd143} : s = 297;
	{8'd154,8'd144} : s = 298;
	{8'd154,8'd145} : s = 299;
	{8'd154,8'd146} : s = 300;
	{8'd154,8'd147} : s = 301;
	{8'd154,8'd148} : s = 302;
	{8'd154,8'd149} : s = 303;
	{8'd154,8'd150} : s = 304;
	{8'd154,8'd151} : s = 305;
	{8'd154,8'd152} : s = 306;
	{8'd154,8'd153} : s = 307;
	{8'd154,8'd154} : s = 308;
	{8'd154,8'd155} : s = 309;
	{8'd154,8'd156} : s = 310;
	{8'd154,8'd157} : s = 311;
	{8'd154,8'd158} : s = 312;
	{8'd154,8'd159} : s = 313;
	{8'd154,8'd160} : s = 314;
	{8'd154,8'd161} : s = 315;
	{8'd154,8'd162} : s = 316;
	{8'd154,8'd163} : s = 317;
	{8'd154,8'd164} : s = 318;
	{8'd154,8'd165} : s = 319;
	{8'd154,8'd166} : s = 320;
	{8'd154,8'd167} : s = 321;
	{8'd154,8'd168} : s = 322;
	{8'd154,8'd169} : s = 323;
	{8'd154,8'd170} : s = 324;
	{8'd154,8'd171} : s = 325;
	{8'd154,8'd172} : s = 326;
	{8'd154,8'd173} : s = 327;
	{8'd154,8'd174} : s = 328;
	{8'd154,8'd175} : s = 329;
	{8'd154,8'd176} : s = 330;
	{8'd154,8'd177} : s = 331;
	{8'd154,8'd178} : s = 332;
	{8'd154,8'd179} : s = 333;
	{8'd154,8'd180} : s = 334;
	{8'd154,8'd181} : s = 335;
	{8'd154,8'd182} : s = 336;
	{8'd154,8'd183} : s = 337;
	{8'd154,8'd184} : s = 338;
	{8'd154,8'd185} : s = 339;
	{8'd154,8'd186} : s = 340;
	{8'd154,8'd187} : s = 341;
	{8'd154,8'd188} : s = 342;
	{8'd154,8'd189} : s = 343;
	{8'd154,8'd190} : s = 344;
	{8'd154,8'd191} : s = 345;
	{8'd154,8'd192} : s = 346;
	{8'd154,8'd193} : s = 347;
	{8'd154,8'd194} : s = 348;
	{8'd154,8'd195} : s = 349;
	{8'd154,8'd196} : s = 350;
	{8'd154,8'd197} : s = 351;
	{8'd154,8'd198} : s = 352;
	{8'd154,8'd199} : s = 353;
	{8'd154,8'd200} : s = 354;
	{8'd154,8'd201} : s = 355;
	{8'd154,8'd202} : s = 356;
	{8'd154,8'd203} : s = 357;
	{8'd154,8'd204} : s = 358;
	{8'd154,8'd205} : s = 359;
	{8'd154,8'd206} : s = 360;
	{8'd154,8'd207} : s = 361;
	{8'd154,8'd208} : s = 362;
	{8'd154,8'd209} : s = 363;
	{8'd154,8'd210} : s = 364;
	{8'd154,8'd211} : s = 365;
	{8'd154,8'd212} : s = 366;
	{8'd154,8'd213} : s = 367;
	{8'd154,8'd214} : s = 368;
	{8'd154,8'd215} : s = 369;
	{8'd154,8'd216} : s = 370;
	{8'd154,8'd217} : s = 371;
	{8'd154,8'd218} : s = 372;
	{8'd154,8'd219} : s = 373;
	{8'd154,8'd220} : s = 374;
	{8'd154,8'd221} : s = 375;
	{8'd154,8'd222} : s = 376;
	{8'd154,8'd223} : s = 377;
	{8'd154,8'd224} : s = 378;
	{8'd154,8'd225} : s = 379;
	{8'd154,8'd226} : s = 380;
	{8'd154,8'd227} : s = 381;
	{8'd154,8'd228} : s = 382;
	{8'd154,8'd229} : s = 383;
	{8'd154,8'd230} : s = 384;
	{8'd154,8'd231} : s = 385;
	{8'd154,8'd232} : s = 386;
	{8'd154,8'd233} : s = 387;
	{8'd154,8'd234} : s = 388;
	{8'd154,8'd235} : s = 389;
	{8'd154,8'd236} : s = 390;
	{8'd154,8'd237} : s = 391;
	{8'd154,8'd238} : s = 392;
	{8'd154,8'd239} : s = 393;
	{8'd154,8'd240} : s = 394;
	{8'd154,8'd241} : s = 395;
	{8'd154,8'd242} : s = 396;
	{8'd154,8'd243} : s = 397;
	{8'd154,8'd244} : s = 398;
	{8'd154,8'd245} : s = 399;
	{8'd154,8'd246} : s = 400;
	{8'd154,8'd247} : s = 401;
	{8'd154,8'd248} : s = 402;
	{8'd154,8'd249} : s = 403;
	{8'd154,8'd250} : s = 404;
	{8'd154,8'd251} : s = 405;
	{8'd154,8'd252} : s = 406;
	{8'd154,8'd253} : s = 407;
	{8'd154,8'd254} : s = 408;
	{8'd154,8'd255} : s = 409;
	{8'd155,8'd0} : s = 155;
	{8'd155,8'd1} : s = 156;
	{8'd155,8'd2} : s = 157;
	{8'd155,8'd3} : s = 158;
	{8'd155,8'd4} : s = 159;
	{8'd155,8'd5} : s = 160;
	{8'd155,8'd6} : s = 161;
	{8'd155,8'd7} : s = 162;
	{8'd155,8'd8} : s = 163;
	{8'd155,8'd9} : s = 164;
	{8'd155,8'd10} : s = 165;
	{8'd155,8'd11} : s = 166;
	{8'd155,8'd12} : s = 167;
	{8'd155,8'd13} : s = 168;
	{8'd155,8'd14} : s = 169;
	{8'd155,8'd15} : s = 170;
	{8'd155,8'd16} : s = 171;
	{8'd155,8'd17} : s = 172;
	{8'd155,8'd18} : s = 173;
	{8'd155,8'd19} : s = 174;
	{8'd155,8'd20} : s = 175;
	{8'd155,8'd21} : s = 176;
	{8'd155,8'd22} : s = 177;
	{8'd155,8'd23} : s = 178;
	{8'd155,8'd24} : s = 179;
	{8'd155,8'd25} : s = 180;
	{8'd155,8'd26} : s = 181;
	{8'd155,8'd27} : s = 182;
	{8'd155,8'd28} : s = 183;
	{8'd155,8'd29} : s = 184;
	{8'd155,8'd30} : s = 185;
	{8'd155,8'd31} : s = 186;
	{8'd155,8'd32} : s = 187;
	{8'd155,8'd33} : s = 188;
	{8'd155,8'd34} : s = 189;
	{8'd155,8'd35} : s = 190;
	{8'd155,8'd36} : s = 191;
	{8'd155,8'd37} : s = 192;
	{8'd155,8'd38} : s = 193;
	{8'd155,8'd39} : s = 194;
	{8'd155,8'd40} : s = 195;
	{8'd155,8'd41} : s = 196;
	{8'd155,8'd42} : s = 197;
	{8'd155,8'd43} : s = 198;
	{8'd155,8'd44} : s = 199;
	{8'd155,8'd45} : s = 200;
	{8'd155,8'd46} : s = 201;
	{8'd155,8'd47} : s = 202;
	{8'd155,8'd48} : s = 203;
	{8'd155,8'd49} : s = 204;
	{8'd155,8'd50} : s = 205;
	{8'd155,8'd51} : s = 206;
	{8'd155,8'd52} : s = 207;
	{8'd155,8'd53} : s = 208;
	{8'd155,8'd54} : s = 209;
	{8'd155,8'd55} : s = 210;
	{8'd155,8'd56} : s = 211;
	{8'd155,8'd57} : s = 212;
	{8'd155,8'd58} : s = 213;
	{8'd155,8'd59} : s = 214;
	{8'd155,8'd60} : s = 215;
	{8'd155,8'd61} : s = 216;
	{8'd155,8'd62} : s = 217;
	{8'd155,8'd63} : s = 218;
	{8'd155,8'd64} : s = 219;
	{8'd155,8'd65} : s = 220;
	{8'd155,8'd66} : s = 221;
	{8'd155,8'd67} : s = 222;
	{8'd155,8'd68} : s = 223;
	{8'd155,8'd69} : s = 224;
	{8'd155,8'd70} : s = 225;
	{8'd155,8'd71} : s = 226;
	{8'd155,8'd72} : s = 227;
	{8'd155,8'd73} : s = 228;
	{8'd155,8'd74} : s = 229;
	{8'd155,8'd75} : s = 230;
	{8'd155,8'd76} : s = 231;
	{8'd155,8'd77} : s = 232;
	{8'd155,8'd78} : s = 233;
	{8'd155,8'd79} : s = 234;
	{8'd155,8'd80} : s = 235;
	{8'd155,8'd81} : s = 236;
	{8'd155,8'd82} : s = 237;
	{8'd155,8'd83} : s = 238;
	{8'd155,8'd84} : s = 239;
	{8'd155,8'd85} : s = 240;
	{8'd155,8'd86} : s = 241;
	{8'd155,8'd87} : s = 242;
	{8'd155,8'd88} : s = 243;
	{8'd155,8'd89} : s = 244;
	{8'd155,8'd90} : s = 245;
	{8'd155,8'd91} : s = 246;
	{8'd155,8'd92} : s = 247;
	{8'd155,8'd93} : s = 248;
	{8'd155,8'd94} : s = 249;
	{8'd155,8'd95} : s = 250;
	{8'd155,8'd96} : s = 251;
	{8'd155,8'd97} : s = 252;
	{8'd155,8'd98} : s = 253;
	{8'd155,8'd99} : s = 254;
	{8'd155,8'd100} : s = 255;
	{8'd155,8'd101} : s = 256;
	{8'd155,8'd102} : s = 257;
	{8'd155,8'd103} : s = 258;
	{8'd155,8'd104} : s = 259;
	{8'd155,8'd105} : s = 260;
	{8'd155,8'd106} : s = 261;
	{8'd155,8'd107} : s = 262;
	{8'd155,8'd108} : s = 263;
	{8'd155,8'd109} : s = 264;
	{8'd155,8'd110} : s = 265;
	{8'd155,8'd111} : s = 266;
	{8'd155,8'd112} : s = 267;
	{8'd155,8'd113} : s = 268;
	{8'd155,8'd114} : s = 269;
	{8'd155,8'd115} : s = 270;
	{8'd155,8'd116} : s = 271;
	{8'd155,8'd117} : s = 272;
	{8'd155,8'd118} : s = 273;
	{8'd155,8'd119} : s = 274;
	{8'd155,8'd120} : s = 275;
	{8'd155,8'd121} : s = 276;
	{8'd155,8'd122} : s = 277;
	{8'd155,8'd123} : s = 278;
	{8'd155,8'd124} : s = 279;
	{8'd155,8'd125} : s = 280;
	{8'd155,8'd126} : s = 281;
	{8'd155,8'd127} : s = 282;
	{8'd155,8'd128} : s = 283;
	{8'd155,8'd129} : s = 284;
	{8'd155,8'd130} : s = 285;
	{8'd155,8'd131} : s = 286;
	{8'd155,8'd132} : s = 287;
	{8'd155,8'd133} : s = 288;
	{8'd155,8'd134} : s = 289;
	{8'd155,8'd135} : s = 290;
	{8'd155,8'd136} : s = 291;
	{8'd155,8'd137} : s = 292;
	{8'd155,8'd138} : s = 293;
	{8'd155,8'd139} : s = 294;
	{8'd155,8'd140} : s = 295;
	{8'd155,8'd141} : s = 296;
	{8'd155,8'd142} : s = 297;
	{8'd155,8'd143} : s = 298;
	{8'd155,8'd144} : s = 299;
	{8'd155,8'd145} : s = 300;
	{8'd155,8'd146} : s = 301;
	{8'd155,8'd147} : s = 302;
	{8'd155,8'd148} : s = 303;
	{8'd155,8'd149} : s = 304;
	{8'd155,8'd150} : s = 305;
	{8'd155,8'd151} : s = 306;
	{8'd155,8'd152} : s = 307;
	{8'd155,8'd153} : s = 308;
	{8'd155,8'd154} : s = 309;
	{8'd155,8'd155} : s = 310;
	{8'd155,8'd156} : s = 311;
	{8'd155,8'd157} : s = 312;
	{8'd155,8'd158} : s = 313;
	{8'd155,8'd159} : s = 314;
	{8'd155,8'd160} : s = 315;
	{8'd155,8'd161} : s = 316;
	{8'd155,8'd162} : s = 317;
	{8'd155,8'd163} : s = 318;
	{8'd155,8'd164} : s = 319;
	{8'd155,8'd165} : s = 320;
	{8'd155,8'd166} : s = 321;
	{8'd155,8'd167} : s = 322;
	{8'd155,8'd168} : s = 323;
	{8'd155,8'd169} : s = 324;
	{8'd155,8'd170} : s = 325;
	{8'd155,8'd171} : s = 326;
	{8'd155,8'd172} : s = 327;
	{8'd155,8'd173} : s = 328;
	{8'd155,8'd174} : s = 329;
	{8'd155,8'd175} : s = 330;
	{8'd155,8'd176} : s = 331;
	{8'd155,8'd177} : s = 332;
	{8'd155,8'd178} : s = 333;
	{8'd155,8'd179} : s = 334;
	{8'd155,8'd180} : s = 335;
	{8'd155,8'd181} : s = 336;
	{8'd155,8'd182} : s = 337;
	{8'd155,8'd183} : s = 338;
	{8'd155,8'd184} : s = 339;
	{8'd155,8'd185} : s = 340;
	{8'd155,8'd186} : s = 341;
	{8'd155,8'd187} : s = 342;
	{8'd155,8'd188} : s = 343;
	{8'd155,8'd189} : s = 344;
	{8'd155,8'd190} : s = 345;
	{8'd155,8'd191} : s = 346;
	{8'd155,8'd192} : s = 347;
	{8'd155,8'd193} : s = 348;
	{8'd155,8'd194} : s = 349;
	{8'd155,8'd195} : s = 350;
	{8'd155,8'd196} : s = 351;
	{8'd155,8'd197} : s = 352;
	{8'd155,8'd198} : s = 353;
	{8'd155,8'd199} : s = 354;
	{8'd155,8'd200} : s = 355;
	{8'd155,8'd201} : s = 356;
	{8'd155,8'd202} : s = 357;
	{8'd155,8'd203} : s = 358;
	{8'd155,8'd204} : s = 359;
	{8'd155,8'd205} : s = 360;
	{8'd155,8'd206} : s = 361;
	{8'd155,8'd207} : s = 362;
	{8'd155,8'd208} : s = 363;
	{8'd155,8'd209} : s = 364;
	{8'd155,8'd210} : s = 365;
	{8'd155,8'd211} : s = 366;
	{8'd155,8'd212} : s = 367;
	{8'd155,8'd213} : s = 368;
	{8'd155,8'd214} : s = 369;
	{8'd155,8'd215} : s = 370;
	{8'd155,8'd216} : s = 371;
	{8'd155,8'd217} : s = 372;
	{8'd155,8'd218} : s = 373;
	{8'd155,8'd219} : s = 374;
	{8'd155,8'd220} : s = 375;
	{8'd155,8'd221} : s = 376;
	{8'd155,8'd222} : s = 377;
	{8'd155,8'd223} : s = 378;
	{8'd155,8'd224} : s = 379;
	{8'd155,8'd225} : s = 380;
	{8'd155,8'd226} : s = 381;
	{8'd155,8'd227} : s = 382;
	{8'd155,8'd228} : s = 383;
	{8'd155,8'd229} : s = 384;
	{8'd155,8'd230} : s = 385;
	{8'd155,8'd231} : s = 386;
	{8'd155,8'd232} : s = 387;
	{8'd155,8'd233} : s = 388;
	{8'd155,8'd234} : s = 389;
	{8'd155,8'd235} : s = 390;
	{8'd155,8'd236} : s = 391;
	{8'd155,8'd237} : s = 392;
	{8'd155,8'd238} : s = 393;
	{8'd155,8'd239} : s = 394;
	{8'd155,8'd240} : s = 395;
	{8'd155,8'd241} : s = 396;
	{8'd155,8'd242} : s = 397;
	{8'd155,8'd243} : s = 398;
	{8'd155,8'd244} : s = 399;
	{8'd155,8'd245} : s = 400;
	{8'd155,8'd246} : s = 401;
	{8'd155,8'd247} : s = 402;
	{8'd155,8'd248} : s = 403;
	{8'd155,8'd249} : s = 404;
	{8'd155,8'd250} : s = 405;
	{8'd155,8'd251} : s = 406;
	{8'd155,8'd252} : s = 407;
	{8'd155,8'd253} : s = 408;
	{8'd155,8'd254} : s = 409;
	{8'd155,8'd255} : s = 410;
	{8'd156,8'd0} : s = 156;
	{8'd156,8'd1} : s = 157;
	{8'd156,8'd2} : s = 158;
	{8'd156,8'd3} : s = 159;
	{8'd156,8'd4} : s = 160;
	{8'd156,8'd5} : s = 161;
	{8'd156,8'd6} : s = 162;
	{8'd156,8'd7} : s = 163;
	{8'd156,8'd8} : s = 164;
	{8'd156,8'd9} : s = 165;
	{8'd156,8'd10} : s = 166;
	{8'd156,8'd11} : s = 167;
	{8'd156,8'd12} : s = 168;
	{8'd156,8'd13} : s = 169;
	{8'd156,8'd14} : s = 170;
	{8'd156,8'd15} : s = 171;
	{8'd156,8'd16} : s = 172;
	{8'd156,8'd17} : s = 173;
	{8'd156,8'd18} : s = 174;
	{8'd156,8'd19} : s = 175;
	{8'd156,8'd20} : s = 176;
	{8'd156,8'd21} : s = 177;
	{8'd156,8'd22} : s = 178;
	{8'd156,8'd23} : s = 179;
	{8'd156,8'd24} : s = 180;
	{8'd156,8'd25} : s = 181;
	{8'd156,8'd26} : s = 182;
	{8'd156,8'd27} : s = 183;
	{8'd156,8'd28} : s = 184;
	{8'd156,8'd29} : s = 185;
	{8'd156,8'd30} : s = 186;
	{8'd156,8'd31} : s = 187;
	{8'd156,8'd32} : s = 188;
	{8'd156,8'd33} : s = 189;
	{8'd156,8'd34} : s = 190;
	{8'd156,8'd35} : s = 191;
	{8'd156,8'd36} : s = 192;
	{8'd156,8'd37} : s = 193;
	{8'd156,8'd38} : s = 194;
	{8'd156,8'd39} : s = 195;
	{8'd156,8'd40} : s = 196;
	{8'd156,8'd41} : s = 197;
	{8'd156,8'd42} : s = 198;
	{8'd156,8'd43} : s = 199;
	{8'd156,8'd44} : s = 200;
	{8'd156,8'd45} : s = 201;
	{8'd156,8'd46} : s = 202;
	{8'd156,8'd47} : s = 203;
	{8'd156,8'd48} : s = 204;
	{8'd156,8'd49} : s = 205;
	{8'd156,8'd50} : s = 206;
	{8'd156,8'd51} : s = 207;
	{8'd156,8'd52} : s = 208;
	{8'd156,8'd53} : s = 209;
	{8'd156,8'd54} : s = 210;
	{8'd156,8'd55} : s = 211;
	{8'd156,8'd56} : s = 212;
	{8'd156,8'd57} : s = 213;
	{8'd156,8'd58} : s = 214;
	{8'd156,8'd59} : s = 215;
	{8'd156,8'd60} : s = 216;
	{8'd156,8'd61} : s = 217;
	{8'd156,8'd62} : s = 218;
	{8'd156,8'd63} : s = 219;
	{8'd156,8'd64} : s = 220;
	{8'd156,8'd65} : s = 221;
	{8'd156,8'd66} : s = 222;
	{8'd156,8'd67} : s = 223;
	{8'd156,8'd68} : s = 224;
	{8'd156,8'd69} : s = 225;
	{8'd156,8'd70} : s = 226;
	{8'd156,8'd71} : s = 227;
	{8'd156,8'd72} : s = 228;
	{8'd156,8'd73} : s = 229;
	{8'd156,8'd74} : s = 230;
	{8'd156,8'd75} : s = 231;
	{8'd156,8'd76} : s = 232;
	{8'd156,8'd77} : s = 233;
	{8'd156,8'd78} : s = 234;
	{8'd156,8'd79} : s = 235;
	{8'd156,8'd80} : s = 236;
	{8'd156,8'd81} : s = 237;
	{8'd156,8'd82} : s = 238;
	{8'd156,8'd83} : s = 239;
	{8'd156,8'd84} : s = 240;
	{8'd156,8'd85} : s = 241;
	{8'd156,8'd86} : s = 242;
	{8'd156,8'd87} : s = 243;
	{8'd156,8'd88} : s = 244;
	{8'd156,8'd89} : s = 245;
	{8'd156,8'd90} : s = 246;
	{8'd156,8'd91} : s = 247;
	{8'd156,8'd92} : s = 248;
	{8'd156,8'd93} : s = 249;
	{8'd156,8'd94} : s = 250;
	{8'd156,8'd95} : s = 251;
	{8'd156,8'd96} : s = 252;
	{8'd156,8'd97} : s = 253;
	{8'd156,8'd98} : s = 254;
	{8'd156,8'd99} : s = 255;
	{8'd156,8'd100} : s = 256;
	{8'd156,8'd101} : s = 257;
	{8'd156,8'd102} : s = 258;
	{8'd156,8'd103} : s = 259;
	{8'd156,8'd104} : s = 260;
	{8'd156,8'd105} : s = 261;
	{8'd156,8'd106} : s = 262;
	{8'd156,8'd107} : s = 263;
	{8'd156,8'd108} : s = 264;
	{8'd156,8'd109} : s = 265;
	{8'd156,8'd110} : s = 266;
	{8'd156,8'd111} : s = 267;
	{8'd156,8'd112} : s = 268;
	{8'd156,8'd113} : s = 269;
	{8'd156,8'd114} : s = 270;
	{8'd156,8'd115} : s = 271;
	{8'd156,8'd116} : s = 272;
	{8'd156,8'd117} : s = 273;
	{8'd156,8'd118} : s = 274;
	{8'd156,8'd119} : s = 275;
	{8'd156,8'd120} : s = 276;
	{8'd156,8'd121} : s = 277;
	{8'd156,8'd122} : s = 278;
	{8'd156,8'd123} : s = 279;
	{8'd156,8'd124} : s = 280;
	{8'd156,8'd125} : s = 281;
	{8'd156,8'd126} : s = 282;
	{8'd156,8'd127} : s = 283;
	{8'd156,8'd128} : s = 284;
	{8'd156,8'd129} : s = 285;
	{8'd156,8'd130} : s = 286;
	{8'd156,8'd131} : s = 287;
	{8'd156,8'd132} : s = 288;
	{8'd156,8'd133} : s = 289;
	{8'd156,8'd134} : s = 290;
	{8'd156,8'd135} : s = 291;
	{8'd156,8'd136} : s = 292;
	{8'd156,8'd137} : s = 293;
	{8'd156,8'd138} : s = 294;
	{8'd156,8'd139} : s = 295;
	{8'd156,8'd140} : s = 296;
	{8'd156,8'd141} : s = 297;
	{8'd156,8'd142} : s = 298;
	{8'd156,8'd143} : s = 299;
	{8'd156,8'd144} : s = 300;
	{8'd156,8'd145} : s = 301;
	{8'd156,8'd146} : s = 302;
	{8'd156,8'd147} : s = 303;
	{8'd156,8'd148} : s = 304;
	{8'd156,8'd149} : s = 305;
	{8'd156,8'd150} : s = 306;
	{8'd156,8'd151} : s = 307;
	{8'd156,8'd152} : s = 308;
	{8'd156,8'd153} : s = 309;
	{8'd156,8'd154} : s = 310;
	{8'd156,8'd155} : s = 311;
	{8'd156,8'd156} : s = 312;
	{8'd156,8'd157} : s = 313;
	{8'd156,8'd158} : s = 314;
	{8'd156,8'd159} : s = 315;
	{8'd156,8'd160} : s = 316;
	{8'd156,8'd161} : s = 317;
	{8'd156,8'd162} : s = 318;
	{8'd156,8'd163} : s = 319;
	{8'd156,8'd164} : s = 320;
	{8'd156,8'd165} : s = 321;
	{8'd156,8'd166} : s = 322;
	{8'd156,8'd167} : s = 323;
	{8'd156,8'd168} : s = 324;
	{8'd156,8'd169} : s = 325;
	{8'd156,8'd170} : s = 326;
	{8'd156,8'd171} : s = 327;
	{8'd156,8'd172} : s = 328;
	{8'd156,8'd173} : s = 329;
	{8'd156,8'd174} : s = 330;
	{8'd156,8'd175} : s = 331;
	{8'd156,8'd176} : s = 332;
	{8'd156,8'd177} : s = 333;
	{8'd156,8'd178} : s = 334;
	{8'd156,8'd179} : s = 335;
	{8'd156,8'd180} : s = 336;
	{8'd156,8'd181} : s = 337;
	{8'd156,8'd182} : s = 338;
	{8'd156,8'd183} : s = 339;
	{8'd156,8'd184} : s = 340;
	{8'd156,8'd185} : s = 341;
	{8'd156,8'd186} : s = 342;
	{8'd156,8'd187} : s = 343;
	{8'd156,8'd188} : s = 344;
	{8'd156,8'd189} : s = 345;
	{8'd156,8'd190} : s = 346;
	{8'd156,8'd191} : s = 347;
	{8'd156,8'd192} : s = 348;
	{8'd156,8'd193} : s = 349;
	{8'd156,8'd194} : s = 350;
	{8'd156,8'd195} : s = 351;
	{8'd156,8'd196} : s = 352;
	{8'd156,8'd197} : s = 353;
	{8'd156,8'd198} : s = 354;
	{8'd156,8'd199} : s = 355;
	{8'd156,8'd200} : s = 356;
	{8'd156,8'd201} : s = 357;
	{8'd156,8'd202} : s = 358;
	{8'd156,8'd203} : s = 359;
	{8'd156,8'd204} : s = 360;
	{8'd156,8'd205} : s = 361;
	{8'd156,8'd206} : s = 362;
	{8'd156,8'd207} : s = 363;
	{8'd156,8'd208} : s = 364;
	{8'd156,8'd209} : s = 365;
	{8'd156,8'd210} : s = 366;
	{8'd156,8'd211} : s = 367;
	{8'd156,8'd212} : s = 368;
	{8'd156,8'd213} : s = 369;
	{8'd156,8'd214} : s = 370;
	{8'd156,8'd215} : s = 371;
	{8'd156,8'd216} : s = 372;
	{8'd156,8'd217} : s = 373;
	{8'd156,8'd218} : s = 374;
	{8'd156,8'd219} : s = 375;
	{8'd156,8'd220} : s = 376;
	{8'd156,8'd221} : s = 377;
	{8'd156,8'd222} : s = 378;
	{8'd156,8'd223} : s = 379;
	{8'd156,8'd224} : s = 380;
	{8'd156,8'd225} : s = 381;
	{8'd156,8'd226} : s = 382;
	{8'd156,8'd227} : s = 383;
	{8'd156,8'd228} : s = 384;
	{8'd156,8'd229} : s = 385;
	{8'd156,8'd230} : s = 386;
	{8'd156,8'd231} : s = 387;
	{8'd156,8'd232} : s = 388;
	{8'd156,8'd233} : s = 389;
	{8'd156,8'd234} : s = 390;
	{8'd156,8'd235} : s = 391;
	{8'd156,8'd236} : s = 392;
	{8'd156,8'd237} : s = 393;
	{8'd156,8'd238} : s = 394;
	{8'd156,8'd239} : s = 395;
	{8'd156,8'd240} : s = 396;
	{8'd156,8'd241} : s = 397;
	{8'd156,8'd242} : s = 398;
	{8'd156,8'd243} : s = 399;
	{8'd156,8'd244} : s = 400;
	{8'd156,8'd245} : s = 401;
	{8'd156,8'd246} : s = 402;
	{8'd156,8'd247} : s = 403;
	{8'd156,8'd248} : s = 404;
	{8'd156,8'd249} : s = 405;
	{8'd156,8'd250} : s = 406;
	{8'd156,8'd251} : s = 407;
	{8'd156,8'd252} : s = 408;
	{8'd156,8'd253} : s = 409;
	{8'd156,8'd254} : s = 410;
	{8'd156,8'd255} : s = 411;
	{8'd157,8'd0} : s = 157;
	{8'd157,8'd1} : s = 158;
	{8'd157,8'd2} : s = 159;
	{8'd157,8'd3} : s = 160;
	{8'd157,8'd4} : s = 161;
	{8'd157,8'd5} : s = 162;
	{8'd157,8'd6} : s = 163;
	{8'd157,8'd7} : s = 164;
	{8'd157,8'd8} : s = 165;
	{8'd157,8'd9} : s = 166;
	{8'd157,8'd10} : s = 167;
	{8'd157,8'd11} : s = 168;
	{8'd157,8'd12} : s = 169;
	{8'd157,8'd13} : s = 170;
	{8'd157,8'd14} : s = 171;
	{8'd157,8'd15} : s = 172;
	{8'd157,8'd16} : s = 173;
	{8'd157,8'd17} : s = 174;
	{8'd157,8'd18} : s = 175;
	{8'd157,8'd19} : s = 176;
	{8'd157,8'd20} : s = 177;
	{8'd157,8'd21} : s = 178;
	{8'd157,8'd22} : s = 179;
	{8'd157,8'd23} : s = 180;
	{8'd157,8'd24} : s = 181;
	{8'd157,8'd25} : s = 182;
	{8'd157,8'd26} : s = 183;
	{8'd157,8'd27} : s = 184;
	{8'd157,8'd28} : s = 185;
	{8'd157,8'd29} : s = 186;
	{8'd157,8'd30} : s = 187;
	{8'd157,8'd31} : s = 188;
	{8'd157,8'd32} : s = 189;
	{8'd157,8'd33} : s = 190;
	{8'd157,8'd34} : s = 191;
	{8'd157,8'd35} : s = 192;
	{8'd157,8'd36} : s = 193;
	{8'd157,8'd37} : s = 194;
	{8'd157,8'd38} : s = 195;
	{8'd157,8'd39} : s = 196;
	{8'd157,8'd40} : s = 197;
	{8'd157,8'd41} : s = 198;
	{8'd157,8'd42} : s = 199;
	{8'd157,8'd43} : s = 200;
	{8'd157,8'd44} : s = 201;
	{8'd157,8'd45} : s = 202;
	{8'd157,8'd46} : s = 203;
	{8'd157,8'd47} : s = 204;
	{8'd157,8'd48} : s = 205;
	{8'd157,8'd49} : s = 206;
	{8'd157,8'd50} : s = 207;
	{8'd157,8'd51} : s = 208;
	{8'd157,8'd52} : s = 209;
	{8'd157,8'd53} : s = 210;
	{8'd157,8'd54} : s = 211;
	{8'd157,8'd55} : s = 212;
	{8'd157,8'd56} : s = 213;
	{8'd157,8'd57} : s = 214;
	{8'd157,8'd58} : s = 215;
	{8'd157,8'd59} : s = 216;
	{8'd157,8'd60} : s = 217;
	{8'd157,8'd61} : s = 218;
	{8'd157,8'd62} : s = 219;
	{8'd157,8'd63} : s = 220;
	{8'd157,8'd64} : s = 221;
	{8'd157,8'd65} : s = 222;
	{8'd157,8'd66} : s = 223;
	{8'd157,8'd67} : s = 224;
	{8'd157,8'd68} : s = 225;
	{8'd157,8'd69} : s = 226;
	{8'd157,8'd70} : s = 227;
	{8'd157,8'd71} : s = 228;
	{8'd157,8'd72} : s = 229;
	{8'd157,8'd73} : s = 230;
	{8'd157,8'd74} : s = 231;
	{8'd157,8'd75} : s = 232;
	{8'd157,8'd76} : s = 233;
	{8'd157,8'd77} : s = 234;
	{8'd157,8'd78} : s = 235;
	{8'd157,8'd79} : s = 236;
	{8'd157,8'd80} : s = 237;
	{8'd157,8'd81} : s = 238;
	{8'd157,8'd82} : s = 239;
	{8'd157,8'd83} : s = 240;
	{8'd157,8'd84} : s = 241;
	{8'd157,8'd85} : s = 242;
	{8'd157,8'd86} : s = 243;
	{8'd157,8'd87} : s = 244;
	{8'd157,8'd88} : s = 245;
	{8'd157,8'd89} : s = 246;
	{8'd157,8'd90} : s = 247;
	{8'd157,8'd91} : s = 248;
	{8'd157,8'd92} : s = 249;
	{8'd157,8'd93} : s = 250;
	{8'd157,8'd94} : s = 251;
	{8'd157,8'd95} : s = 252;
	{8'd157,8'd96} : s = 253;
	{8'd157,8'd97} : s = 254;
	{8'd157,8'd98} : s = 255;
	{8'd157,8'd99} : s = 256;
	{8'd157,8'd100} : s = 257;
	{8'd157,8'd101} : s = 258;
	{8'd157,8'd102} : s = 259;
	{8'd157,8'd103} : s = 260;
	{8'd157,8'd104} : s = 261;
	{8'd157,8'd105} : s = 262;
	{8'd157,8'd106} : s = 263;
	{8'd157,8'd107} : s = 264;
	{8'd157,8'd108} : s = 265;
	{8'd157,8'd109} : s = 266;
	{8'd157,8'd110} : s = 267;
	{8'd157,8'd111} : s = 268;
	{8'd157,8'd112} : s = 269;
	{8'd157,8'd113} : s = 270;
	{8'd157,8'd114} : s = 271;
	{8'd157,8'd115} : s = 272;
	{8'd157,8'd116} : s = 273;
	{8'd157,8'd117} : s = 274;
	{8'd157,8'd118} : s = 275;
	{8'd157,8'd119} : s = 276;
	{8'd157,8'd120} : s = 277;
	{8'd157,8'd121} : s = 278;
	{8'd157,8'd122} : s = 279;
	{8'd157,8'd123} : s = 280;
	{8'd157,8'd124} : s = 281;
	{8'd157,8'd125} : s = 282;
	{8'd157,8'd126} : s = 283;
	{8'd157,8'd127} : s = 284;
	{8'd157,8'd128} : s = 285;
	{8'd157,8'd129} : s = 286;
	{8'd157,8'd130} : s = 287;
	{8'd157,8'd131} : s = 288;
	{8'd157,8'd132} : s = 289;
	{8'd157,8'd133} : s = 290;
	{8'd157,8'd134} : s = 291;
	{8'd157,8'd135} : s = 292;
	{8'd157,8'd136} : s = 293;
	{8'd157,8'd137} : s = 294;
	{8'd157,8'd138} : s = 295;
	{8'd157,8'd139} : s = 296;
	{8'd157,8'd140} : s = 297;
	{8'd157,8'd141} : s = 298;
	{8'd157,8'd142} : s = 299;
	{8'd157,8'd143} : s = 300;
	{8'd157,8'd144} : s = 301;
	{8'd157,8'd145} : s = 302;
	{8'd157,8'd146} : s = 303;
	{8'd157,8'd147} : s = 304;
	{8'd157,8'd148} : s = 305;
	{8'd157,8'd149} : s = 306;
	{8'd157,8'd150} : s = 307;
	{8'd157,8'd151} : s = 308;
	{8'd157,8'd152} : s = 309;
	{8'd157,8'd153} : s = 310;
	{8'd157,8'd154} : s = 311;
	{8'd157,8'd155} : s = 312;
	{8'd157,8'd156} : s = 313;
	{8'd157,8'd157} : s = 314;
	{8'd157,8'd158} : s = 315;
	{8'd157,8'd159} : s = 316;
	{8'd157,8'd160} : s = 317;
	{8'd157,8'd161} : s = 318;
	{8'd157,8'd162} : s = 319;
	{8'd157,8'd163} : s = 320;
	{8'd157,8'd164} : s = 321;
	{8'd157,8'd165} : s = 322;
	{8'd157,8'd166} : s = 323;
	{8'd157,8'd167} : s = 324;
	{8'd157,8'd168} : s = 325;
	{8'd157,8'd169} : s = 326;
	{8'd157,8'd170} : s = 327;
	{8'd157,8'd171} : s = 328;
	{8'd157,8'd172} : s = 329;
	{8'd157,8'd173} : s = 330;
	{8'd157,8'd174} : s = 331;
	{8'd157,8'd175} : s = 332;
	{8'd157,8'd176} : s = 333;
	{8'd157,8'd177} : s = 334;
	{8'd157,8'd178} : s = 335;
	{8'd157,8'd179} : s = 336;
	{8'd157,8'd180} : s = 337;
	{8'd157,8'd181} : s = 338;
	{8'd157,8'd182} : s = 339;
	{8'd157,8'd183} : s = 340;
	{8'd157,8'd184} : s = 341;
	{8'd157,8'd185} : s = 342;
	{8'd157,8'd186} : s = 343;
	{8'd157,8'd187} : s = 344;
	{8'd157,8'd188} : s = 345;
	{8'd157,8'd189} : s = 346;
	{8'd157,8'd190} : s = 347;
	{8'd157,8'd191} : s = 348;
	{8'd157,8'd192} : s = 349;
	{8'd157,8'd193} : s = 350;
	{8'd157,8'd194} : s = 351;
	{8'd157,8'd195} : s = 352;
	{8'd157,8'd196} : s = 353;
	{8'd157,8'd197} : s = 354;
	{8'd157,8'd198} : s = 355;
	{8'd157,8'd199} : s = 356;
	{8'd157,8'd200} : s = 357;
	{8'd157,8'd201} : s = 358;
	{8'd157,8'd202} : s = 359;
	{8'd157,8'd203} : s = 360;
	{8'd157,8'd204} : s = 361;
	{8'd157,8'd205} : s = 362;
	{8'd157,8'd206} : s = 363;
	{8'd157,8'd207} : s = 364;
	{8'd157,8'd208} : s = 365;
	{8'd157,8'd209} : s = 366;
	{8'd157,8'd210} : s = 367;
	{8'd157,8'd211} : s = 368;
	{8'd157,8'd212} : s = 369;
	{8'd157,8'd213} : s = 370;
	{8'd157,8'd214} : s = 371;
	{8'd157,8'd215} : s = 372;
	{8'd157,8'd216} : s = 373;
	{8'd157,8'd217} : s = 374;
	{8'd157,8'd218} : s = 375;
	{8'd157,8'd219} : s = 376;
	{8'd157,8'd220} : s = 377;
	{8'd157,8'd221} : s = 378;
	{8'd157,8'd222} : s = 379;
	{8'd157,8'd223} : s = 380;
	{8'd157,8'd224} : s = 381;
	{8'd157,8'd225} : s = 382;
	{8'd157,8'd226} : s = 383;
	{8'd157,8'd227} : s = 384;
	{8'd157,8'd228} : s = 385;
	{8'd157,8'd229} : s = 386;
	{8'd157,8'd230} : s = 387;
	{8'd157,8'd231} : s = 388;
	{8'd157,8'd232} : s = 389;
	{8'd157,8'd233} : s = 390;
	{8'd157,8'd234} : s = 391;
	{8'd157,8'd235} : s = 392;
	{8'd157,8'd236} : s = 393;
	{8'd157,8'd237} : s = 394;
	{8'd157,8'd238} : s = 395;
	{8'd157,8'd239} : s = 396;
	{8'd157,8'd240} : s = 397;
	{8'd157,8'd241} : s = 398;
	{8'd157,8'd242} : s = 399;
	{8'd157,8'd243} : s = 400;
	{8'd157,8'd244} : s = 401;
	{8'd157,8'd245} : s = 402;
	{8'd157,8'd246} : s = 403;
	{8'd157,8'd247} : s = 404;
	{8'd157,8'd248} : s = 405;
	{8'd157,8'd249} : s = 406;
	{8'd157,8'd250} : s = 407;
	{8'd157,8'd251} : s = 408;
	{8'd157,8'd252} : s = 409;
	{8'd157,8'd253} : s = 410;
	{8'd157,8'd254} : s = 411;
	{8'd157,8'd255} : s = 412;
	{8'd158,8'd0} : s = 158;
	{8'd158,8'd1} : s = 159;
	{8'd158,8'd2} : s = 160;
	{8'd158,8'd3} : s = 161;
	{8'd158,8'd4} : s = 162;
	{8'd158,8'd5} : s = 163;
	{8'd158,8'd6} : s = 164;
	{8'd158,8'd7} : s = 165;
	{8'd158,8'd8} : s = 166;
	{8'd158,8'd9} : s = 167;
	{8'd158,8'd10} : s = 168;
	{8'd158,8'd11} : s = 169;
	{8'd158,8'd12} : s = 170;
	{8'd158,8'd13} : s = 171;
	{8'd158,8'd14} : s = 172;
	{8'd158,8'd15} : s = 173;
	{8'd158,8'd16} : s = 174;
	{8'd158,8'd17} : s = 175;
	{8'd158,8'd18} : s = 176;
	{8'd158,8'd19} : s = 177;
	{8'd158,8'd20} : s = 178;
	{8'd158,8'd21} : s = 179;
	{8'd158,8'd22} : s = 180;
	{8'd158,8'd23} : s = 181;
	{8'd158,8'd24} : s = 182;
	{8'd158,8'd25} : s = 183;
	{8'd158,8'd26} : s = 184;
	{8'd158,8'd27} : s = 185;
	{8'd158,8'd28} : s = 186;
	{8'd158,8'd29} : s = 187;
	{8'd158,8'd30} : s = 188;
	{8'd158,8'd31} : s = 189;
	{8'd158,8'd32} : s = 190;
	{8'd158,8'd33} : s = 191;
	{8'd158,8'd34} : s = 192;
	{8'd158,8'd35} : s = 193;
	{8'd158,8'd36} : s = 194;
	{8'd158,8'd37} : s = 195;
	{8'd158,8'd38} : s = 196;
	{8'd158,8'd39} : s = 197;
	{8'd158,8'd40} : s = 198;
	{8'd158,8'd41} : s = 199;
	{8'd158,8'd42} : s = 200;
	{8'd158,8'd43} : s = 201;
	{8'd158,8'd44} : s = 202;
	{8'd158,8'd45} : s = 203;
	{8'd158,8'd46} : s = 204;
	{8'd158,8'd47} : s = 205;
	{8'd158,8'd48} : s = 206;
	{8'd158,8'd49} : s = 207;
	{8'd158,8'd50} : s = 208;
	{8'd158,8'd51} : s = 209;
	{8'd158,8'd52} : s = 210;
	{8'd158,8'd53} : s = 211;
	{8'd158,8'd54} : s = 212;
	{8'd158,8'd55} : s = 213;
	{8'd158,8'd56} : s = 214;
	{8'd158,8'd57} : s = 215;
	{8'd158,8'd58} : s = 216;
	{8'd158,8'd59} : s = 217;
	{8'd158,8'd60} : s = 218;
	{8'd158,8'd61} : s = 219;
	{8'd158,8'd62} : s = 220;
	{8'd158,8'd63} : s = 221;
	{8'd158,8'd64} : s = 222;
	{8'd158,8'd65} : s = 223;
	{8'd158,8'd66} : s = 224;
	{8'd158,8'd67} : s = 225;
	{8'd158,8'd68} : s = 226;
	{8'd158,8'd69} : s = 227;
	{8'd158,8'd70} : s = 228;
	{8'd158,8'd71} : s = 229;
	{8'd158,8'd72} : s = 230;
	{8'd158,8'd73} : s = 231;
	{8'd158,8'd74} : s = 232;
	{8'd158,8'd75} : s = 233;
	{8'd158,8'd76} : s = 234;
	{8'd158,8'd77} : s = 235;
	{8'd158,8'd78} : s = 236;
	{8'd158,8'd79} : s = 237;
	{8'd158,8'd80} : s = 238;
	{8'd158,8'd81} : s = 239;
	{8'd158,8'd82} : s = 240;
	{8'd158,8'd83} : s = 241;
	{8'd158,8'd84} : s = 242;
	{8'd158,8'd85} : s = 243;
	{8'd158,8'd86} : s = 244;
	{8'd158,8'd87} : s = 245;
	{8'd158,8'd88} : s = 246;
	{8'd158,8'd89} : s = 247;
	{8'd158,8'd90} : s = 248;
	{8'd158,8'd91} : s = 249;
	{8'd158,8'd92} : s = 250;
	{8'd158,8'd93} : s = 251;
	{8'd158,8'd94} : s = 252;
	{8'd158,8'd95} : s = 253;
	{8'd158,8'd96} : s = 254;
	{8'd158,8'd97} : s = 255;
	{8'd158,8'd98} : s = 256;
	{8'd158,8'd99} : s = 257;
	{8'd158,8'd100} : s = 258;
	{8'd158,8'd101} : s = 259;
	{8'd158,8'd102} : s = 260;
	{8'd158,8'd103} : s = 261;
	{8'd158,8'd104} : s = 262;
	{8'd158,8'd105} : s = 263;
	{8'd158,8'd106} : s = 264;
	{8'd158,8'd107} : s = 265;
	{8'd158,8'd108} : s = 266;
	{8'd158,8'd109} : s = 267;
	{8'd158,8'd110} : s = 268;
	{8'd158,8'd111} : s = 269;
	{8'd158,8'd112} : s = 270;
	{8'd158,8'd113} : s = 271;
	{8'd158,8'd114} : s = 272;
	{8'd158,8'd115} : s = 273;
	{8'd158,8'd116} : s = 274;
	{8'd158,8'd117} : s = 275;
	{8'd158,8'd118} : s = 276;
	{8'd158,8'd119} : s = 277;
	{8'd158,8'd120} : s = 278;
	{8'd158,8'd121} : s = 279;
	{8'd158,8'd122} : s = 280;
	{8'd158,8'd123} : s = 281;
	{8'd158,8'd124} : s = 282;
	{8'd158,8'd125} : s = 283;
	{8'd158,8'd126} : s = 284;
	{8'd158,8'd127} : s = 285;
	{8'd158,8'd128} : s = 286;
	{8'd158,8'd129} : s = 287;
	{8'd158,8'd130} : s = 288;
	{8'd158,8'd131} : s = 289;
	{8'd158,8'd132} : s = 290;
	{8'd158,8'd133} : s = 291;
	{8'd158,8'd134} : s = 292;
	{8'd158,8'd135} : s = 293;
	{8'd158,8'd136} : s = 294;
	{8'd158,8'd137} : s = 295;
	{8'd158,8'd138} : s = 296;
	{8'd158,8'd139} : s = 297;
	{8'd158,8'd140} : s = 298;
	{8'd158,8'd141} : s = 299;
	{8'd158,8'd142} : s = 300;
	{8'd158,8'd143} : s = 301;
	{8'd158,8'd144} : s = 302;
	{8'd158,8'd145} : s = 303;
	{8'd158,8'd146} : s = 304;
	{8'd158,8'd147} : s = 305;
	{8'd158,8'd148} : s = 306;
	{8'd158,8'd149} : s = 307;
	{8'd158,8'd150} : s = 308;
	{8'd158,8'd151} : s = 309;
	{8'd158,8'd152} : s = 310;
	{8'd158,8'd153} : s = 311;
	{8'd158,8'd154} : s = 312;
	{8'd158,8'd155} : s = 313;
	{8'd158,8'd156} : s = 314;
	{8'd158,8'd157} : s = 315;
	{8'd158,8'd158} : s = 316;
	{8'd158,8'd159} : s = 317;
	{8'd158,8'd160} : s = 318;
	{8'd158,8'd161} : s = 319;
	{8'd158,8'd162} : s = 320;
	{8'd158,8'd163} : s = 321;
	{8'd158,8'd164} : s = 322;
	{8'd158,8'd165} : s = 323;
	{8'd158,8'd166} : s = 324;
	{8'd158,8'd167} : s = 325;
	{8'd158,8'd168} : s = 326;
	{8'd158,8'd169} : s = 327;
	{8'd158,8'd170} : s = 328;
	{8'd158,8'd171} : s = 329;
	{8'd158,8'd172} : s = 330;
	{8'd158,8'd173} : s = 331;
	{8'd158,8'd174} : s = 332;
	{8'd158,8'd175} : s = 333;
	{8'd158,8'd176} : s = 334;
	{8'd158,8'd177} : s = 335;
	{8'd158,8'd178} : s = 336;
	{8'd158,8'd179} : s = 337;
	{8'd158,8'd180} : s = 338;
	{8'd158,8'd181} : s = 339;
	{8'd158,8'd182} : s = 340;
	{8'd158,8'd183} : s = 341;
	{8'd158,8'd184} : s = 342;
	{8'd158,8'd185} : s = 343;
	{8'd158,8'd186} : s = 344;
	{8'd158,8'd187} : s = 345;
	{8'd158,8'd188} : s = 346;
	{8'd158,8'd189} : s = 347;
	{8'd158,8'd190} : s = 348;
	{8'd158,8'd191} : s = 349;
	{8'd158,8'd192} : s = 350;
	{8'd158,8'd193} : s = 351;
	{8'd158,8'd194} : s = 352;
	{8'd158,8'd195} : s = 353;
	{8'd158,8'd196} : s = 354;
	{8'd158,8'd197} : s = 355;
	{8'd158,8'd198} : s = 356;
	{8'd158,8'd199} : s = 357;
	{8'd158,8'd200} : s = 358;
	{8'd158,8'd201} : s = 359;
	{8'd158,8'd202} : s = 360;
	{8'd158,8'd203} : s = 361;
	{8'd158,8'd204} : s = 362;
	{8'd158,8'd205} : s = 363;
	{8'd158,8'd206} : s = 364;
	{8'd158,8'd207} : s = 365;
	{8'd158,8'd208} : s = 366;
	{8'd158,8'd209} : s = 367;
	{8'd158,8'd210} : s = 368;
	{8'd158,8'd211} : s = 369;
	{8'd158,8'd212} : s = 370;
	{8'd158,8'd213} : s = 371;
	{8'd158,8'd214} : s = 372;
	{8'd158,8'd215} : s = 373;
	{8'd158,8'd216} : s = 374;
	{8'd158,8'd217} : s = 375;
	{8'd158,8'd218} : s = 376;
	{8'd158,8'd219} : s = 377;
	{8'd158,8'd220} : s = 378;
	{8'd158,8'd221} : s = 379;
	{8'd158,8'd222} : s = 380;
	{8'd158,8'd223} : s = 381;
	{8'd158,8'd224} : s = 382;
	{8'd158,8'd225} : s = 383;
	{8'd158,8'd226} : s = 384;
	{8'd158,8'd227} : s = 385;
	{8'd158,8'd228} : s = 386;
	{8'd158,8'd229} : s = 387;
	{8'd158,8'd230} : s = 388;
	{8'd158,8'd231} : s = 389;
	{8'd158,8'd232} : s = 390;
	{8'd158,8'd233} : s = 391;
	{8'd158,8'd234} : s = 392;
	{8'd158,8'd235} : s = 393;
	{8'd158,8'd236} : s = 394;
	{8'd158,8'd237} : s = 395;
	{8'd158,8'd238} : s = 396;
	{8'd158,8'd239} : s = 397;
	{8'd158,8'd240} : s = 398;
	{8'd158,8'd241} : s = 399;
	{8'd158,8'd242} : s = 400;
	{8'd158,8'd243} : s = 401;
	{8'd158,8'd244} : s = 402;
	{8'd158,8'd245} : s = 403;
	{8'd158,8'd246} : s = 404;
	{8'd158,8'd247} : s = 405;
	{8'd158,8'd248} : s = 406;
	{8'd158,8'd249} : s = 407;
	{8'd158,8'd250} : s = 408;
	{8'd158,8'd251} : s = 409;
	{8'd158,8'd252} : s = 410;
	{8'd158,8'd253} : s = 411;
	{8'd158,8'd254} : s = 412;
	{8'd158,8'd255} : s = 413;
	{8'd159,8'd0} : s = 159;
	{8'd159,8'd1} : s = 160;
	{8'd159,8'd2} : s = 161;
	{8'd159,8'd3} : s = 162;
	{8'd159,8'd4} : s = 163;
	{8'd159,8'd5} : s = 164;
	{8'd159,8'd6} : s = 165;
	{8'd159,8'd7} : s = 166;
	{8'd159,8'd8} : s = 167;
	{8'd159,8'd9} : s = 168;
	{8'd159,8'd10} : s = 169;
	{8'd159,8'd11} : s = 170;
	{8'd159,8'd12} : s = 171;
	{8'd159,8'd13} : s = 172;
	{8'd159,8'd14} : s = 173;
	{8'd159,8'd15} : s = 174;
	{8'd159,8'd16} : s = 175;
	{8'd159,8'd17} : s = 176;
	{8'd159,8'd18} : s = 177;
	{8'd159,8'd19} : s = 178;
	{8'd159,8'd20} : s = 179;
	{8'd159,8'd21} : s = 180;
	{8'd159,8'd22} : s = 181;
	{8'd159,8'd23} : s = 182;
	{8'd159,8'd24} : s = 183;
	{8'd159,8'd25} : s = 184;
	{8'd159,8'd26} : s = 185;
	{8'd159,8'd27} : s = 186;
	{8'd159,8'd28} : s = 187;
	{8'd159,8'd29} : s = 188;
	{8'd159,8'd30} : s = 189;
	{8'd159,8'd31} : s = 190;
	{8'd159,8'd32} : s = 191;
	{8'd159,8'd33} : s = 192;
	{8'd159,8'd34} : s = 193;
	{8'd159,8'd35} : s = 194;
	{8'd159,8'd36} : s = 195;
	{8'd159,8'd37} : s = 196;
	{8'd159,8'd38} : s = 197;
	{8'd159,8'd39} : s = 198;
	{8'd159,8'd40} : s = 199;
	{8'd159,8'd41} : s = 200;
	{8'd159,8'd42} : s = 201;
	{8'd159,8'd43} : s = 202;
	{8'd159,8'd44} : s = 203;
	{8'd159,8'd45} : s = 204;
	{8'd159,8'd46} : s = 205;
	{8'd159,8'd47} : s = 206;
	{8'd159,8'd48} : s = 207;
	{8'd159,8'd49} : s = 208;
	{8'd159,8'd50} : s = 209;
	{8'd159,8'd51} : s = 210;
	{8'd159,8'd52} : s = 211;
	{8'd159,8'd53} : s = 212;
	{8'd159,8'd54} : s = 213;
	{8'd159,8'd55} : s = 214;
	{8'd159,8'd56} : s = 215;
	{8'd159,8'd57} : s = 216;
	{8'd159,8'd58} : s = 217;
	{8'd159,8'd59} : s = 218;
	{8'd159,8'd60} : s = 219;
	{8'd159,8'd61} : s = 220;
	{8'd159,8'd62} : s = 221;
	{8'd159,8'd63} : s = 222;
	{8'd159,8'd64} : s = 223;
	{8'd159,8'd65} : s = 224;
	{8'd159,8'd66} : s = 225;
	{8'd159,8'd67} : s = 226;
	{8'd159,8'd68} : s = 227;
	{8'd159,8'd69} : s = 228;
	{8'd159,8'd70} : s = 229;
	{8'd159,8'd71} : s = 230;
	{8'd159,8'd72} : s = 231;
	{8'd159,8'd73} : s = 232;
	{8'd159,8'd74} : s = 233;
	{8'd159,8'd75} : s = 234;
	{8'd159,8'd76} : s = 235;
	{8'd159,8'd77} : s = 236;
	{8'd159,8'd78} : s = 237;
	{8'd159,8'd79} : s = 238;
	{8'd159,8'd80} : s = 239;
	{8'd159,8'd81} : s = 240;
	{8'd159,8'd82} : s = 241;
	{8'd159,8'd83} : s = 242;
	{8'd159,8'd84} : s = 243;
	{8'd159,8'd85} : s = 244;
	{8'd159,8'd86} : s = 245;
	{8'd159,8'd87} : s = 246;
	{8'd159,8'd88} : s = 247;
	{8'd159,8'd89} : s = 248;
	{8'd159,8'd90} : s = 249;
	{8'd159,8'd91} : s = 250;
	{8'd159,8'd92} : s = 251;
	{8'd159,8'd93} : s = 252;
	{8'd159,8'd94} : s = 253;
	{8'd159,8'd95} : s = 254;
	{8'd159,8'd96} : s = 255;
	{8'd159,8'd97} : s = 256;
	{8'd159,8'd98} : s = 257;
	{8'd159,8'd99} : s = 258;
	{8'd159,8'd100} : s = 259;
	{8'd159,8'd101} : s = 260;
	{8'd159,8'd102} : s = 261;
	{8'd159,8'd103} : s = 262;
	{8'd159,8'd104} : s = 263;
	{8'd159,8'd105} : s = 264;
	{8'd159,8'd106} : s = 265;
	{8'd159,8'd107} : s = 266;
	{8'd159,8'd108} : s = 267;
	{8'd159,8'd109} : s = 268;
	{8'd159,8'd110} : s = 269;
	{8'd159,8'd111} : s = 270;
	{8'd159,8'd112} : s = 271;
	{8'd159,8'd113} : s = 272;
	{8'd159,8'd114} : s = 273;
	{8'd159,8'd115} : s = 274;
	{8'd159,8'd116} : s = 275;
	{8'd159,8'd117} : s = 276;
	{8'd159,8'd118} : s = 277;
	{8'd159,8'd119} : s = 278;
	{8'd159,8'd120} : s = 279;
	{8'd159,8'd121} : s = 280;
	{8'd159,8'd122} : s = 281;
	{8'd159,8'd123} : s = 282;
	{8'd159,8'd124} : s = 283;
	{8'd159,8'd125} : s = 284;
	{8'd159,8'd126} : s = 285;
	{8'd159,8'd127} : s = 286;
	{8'd159,8'd128} : s = 287;
	{8'd159,8'd129} : s = 288;
	{8'd159,8'd130} : s = 289;
	{8'd159,8'd131} : s = 290;
	{8'd159,8'd132} : s = 291;
	{8'd159,8'd133} : s = 292;
	{8'd159,8'd134} : s = 293;
	{8'd159,8'd135} : s = 294;
	{8'd159,8'd136} : s = 295;
	{8'd159,8'd137} : s = 296;
	{8'd159,8'd138} : s = 297;
	{8'd159,8'd139} : s = 298;
	{8'd159,8'd140} : s = 299;
	{8'd159,8'd141} : s = 300;
	{8'd159,8'd142} : s = 301;
	{8'd159,8'd143} : s = 302;
	{8'd159,8'd144} : s = 303;
	{8'd159,8'd145} : s = 304;
	{8'd159,8'd146} : s = 305;
	{8'd159,8'd147} : s = 306;
	{8'd159,8'd148} : s = 307;
	{8'd159,8'd149} : s = 308;
	{8'd159,8'd150} : s = 309;
	{8'd159,8'd151} : s = 310;
	{8'd159,8'd152} : s = 311;
	{8'd159,8'd153} : s = 312;
	{8'd159,8'd154} : s = 313;
	{8'd159,8'd155} : s = 314;
	{8'd159,8'd156} : s = 315;
	{8'd159,8'd157} : s = 316;
	{8'd159,8'd158} : s = 317;
	{8'd159,8'd159} : s = 318;
	{8'd159,8'd160} : s = 319;
	{8'd159,8'd161} : s = 320;
	{8'd159,8'd162} : s = 321;
	{8'd159,8'd163} : s = 322;
	{8'd159,8'd164} : s = 323;
	{8'd159,8'd165} : s = 324;
	{8'd159,8'd166} : s = 325;
	{8'd159,8'd167} : s = 326;
	{8'd159,8'd168} : s = 327;
	{8'd159,8'd169} : s = 328;
	{8'd159,8'd170} : s = 329;
	{8'd159,8'd171} : s = 330;
	{8'd159,8'd172} : s = 331;
	{8'd159,8'd173} : s = 332;
	{8'd159,8'd174} : s = 333;
	{8'd159,8'd175} : s = 334;
	{8'd159,8'd176} : s = 335;
	{8'd159,8'd177} : s = 336;
	{8'd159,8'd178} : s = 337;
	{8'd159,8'd179} : s = 338;
	{8'd159,8'd180} : s = 339;
	{8'd159,8'd181} : s = 340;
	{8'd159,8'd182} : s = 341;
	{8'd159,8'd183} : s = 342;
	{8'd159,8'd184} : s = 343;
	{8'd159,8'd185} : s = 344;
	{8'd159,8'd186} : s = 345;
	{8'd159,8'd187} : s = 346;
	{8'd159,8'd188} : s = 347;
	{8'd159,8'd189} : s = 348;
	{8'd159,8'd190} : s = 349;
	{8'd159,8'd191} : s = 350;
	{8'd159,8'd192} : s = 351;
	{8'd159,8'd193} : s = 352;
	{8'd159,8'd194} : s = 353;
	{8'd159,8'd195} : s = 354;
	{8'd159,8'd196} : s = 355;
	{8'd159,8'd197} : s = 356;
	{8'd159,8'd198} : s = 357;
	{8'd159,8'd199} : s = 358;
	{8'd159,8'd200} : s = 359;
	{8'd159,8'd201} : s = 360;
	{8'd159,8'd202} : s = 361;
	{8'd159,8'd203} : s = 362;
	{8'd159,8'd204} : s = 363;
	{8'd159,8'd205} : s = 364;
	{8'd159,8'd206} : s = 365;
	{8'd159,8'd207} : s = 366;
	{8'd159,8'd208} : s = 367;
	{8'd159,8'd209} : s = 368;
	{8'd159,8'd210} : s = 369;
	{8'd159,8'd211} : s = 370;
	{8'd159,8'd212} : s = 371;
	{8'd159,8'd213} : s = 372;
	{8'd159,8'd214} : s = 373;
	{8'd159,8'd215} : s = 374;
	{8'd159,8'd216} : s = 375;
	{8'd159,8'd217} : s = 376;
	{8'd159,8'd218} : s = 377;
	{8'd159,8'd219} : s = 378;
	{8'd159,8'd220} : s = 379;
	{8'd159,8'd221} : s = 380;
	{8'd159,8'd222} : s = 381;
	{8'd159,8'd223} : s = 382;
	{8'd159,8'd224} : s = 383;
	{8'd159,8'd225} : s = 384;
	{8'd159,8'd226} : s = 385;
	{8'd159,8'd227} : s = 386;
	{8'd159,8'd228} : s = 387;
	{8'd159,8'd229} : s = 388;
	{8'd159,8'd230} : s = 389;
	{8'd159,8'd231} : s = 390;
	{8'd159,8'd232} : s = 391;
	{8'd159,8'd233} : s = 392;
	{8'd159,8'd234} : s = 393;
	{8'd159,8'd235} : s = 394;
	{8'd159,8'd236} : s = 395;
	{8'd159,8'd237} : s = 396;
	{8'd159,8'd238} : s = 397;
	{8'd159,8'd239} : s = 398;
	{8'd159,8'd240} : s = 399;
	{8'd159,8'd241} : s = 400;
	{8'd159,8'd242} : s = 401;
	{8'd159,8'd243} : s = 402;
	{8'd159,8'd244} : s = 403;
	{8'd159,8'd245} : s = 404;
	{8'd159,8'd246} : s = 405;
	{8'd159,8'd247} : s = 406;
	{8'd159,8'd248} : s = 407;
	{8'd159,8'd249} : s = 408;
	{8'd159,8'd250} : s = 409;
	{8'd159,8'd251} : s = 410;
	{8'd159,8'd252} : s = 411;
	{8'd159,8'd253} : s = 412;
	{8'd159,8'd254} : s = 413;
	{8'd159,8'd255} : s = 414;
	{8'd160,8'd0} : s = 160;
	{8'd160,8'd1} : s = 161;
	{8'd160,8'd2} : s = 162;
	{8'd160,8'd3} : s = 163;
	{8'd160,8'd4} : s = 164;
	{8'd160,8'd5} : s = 165;
	{8'd160,8'd6} : s = 166;
	{8'd160,8'd7} : s = 167;
	{8'd160,8'd8} : s = 168;
	{8'd160,8'd9} : s = 169;
	{8'd160,8'd10} : s = 170;
	{8'd160,8'd11} : s = 171;
	{8'd160,8'd12} : s = 172;
	{8'd160,8'd13} : s = 173;
	{8'd160,8'd14} : s = 174;
	{8'd160,8'd15} : s = 175;
	{8'd160,8'd16} : s = 176;
	{8'd160,8'd17} : s = 177;
	{8'd160,8'd18} : s = 178;
	{8'd160,8'd19} : s = 179;
	{8'd160,8'd20} : s = 180;
	{8'd160,8'd21} : s = 181;
	{8'd160,8'd22} : s = 182;
	{8'd160,8'd23} : s = 183;
	{8'd160,8'd24} : s = 184;
	{8'd160,8'd25} : s = 185;
	{8'd160,8'd26} : s = 186;
	{8'd160,8'd27} : s = 187;
	{8'd160,8'd28} : s = 188;
	{8'd160,8'd29} : s = 189;
	{8'd160,8'd30} : s = 190;
	{8'd160,8'd31} : s = 191;
	{8'd160,8'd32} : s = 192;
	{8'd160,8'd33} : s = 193;
	{8'd160,8'd34} : s = 194;
	{8'd160,8'd35} : s = 195;
	{8'd160,8'd36} : s = 196;
	{8'd160,8'd37} : s = 197;
	{8'd160,8'd38} : s = 198;
	{8'd160,8'd39} : s = 199;
	{8'd160,8'd40} : s = 200;
	{8'd160,8'd41} : s = 201;
	{8'd160,8'd42} : s = 202;
	{8'd160,8'd43} : s = 203;
	{8'd160,8'd44} : s = 204;
	{8'd160,8'd45} : s = 205;
	{8'd160,8'd46} : s = 206;
	{8'd160,8'd47} : s = 207;
	{8'd160,8'd48} : s = 208;
	{8'd160,8'd49} : s = 209;
	{8'd160,8'd50} : s = 210;
	{8'd160,8'd51} : s = 211;
	{8'd160,8'd52} : s = 212;
	{8'd160,8'd53} : s = 213;
	{8'd160,8'd54} : s = 214;
	{8'd160,8'd55} : s = 215;
	{8'd160,8'd56} : s = 216;
	{8'd160,8'd57} : s = 217;
	{8'd160,8'd58} : s = 218;
	{8'd160,8'd59} : s = 219;
	{8'd160,8'd60} : s = 220;
	{8'd160,8'd61} : s = 221;
	{8'd160,8'd62} : s = 222;
	{8'd160,8'd63} : s = 223;
	{8'd160,8'd64} : s = 224;
	{8'd160,8'd65} : s = 225;
	{8'd160,8'd66} : s = 226;
	{8'd160,8'd67} : s = 227;
	{8'd160,8'd68} : s = 228;
	{8'd160,8'd69} : s = 229;
	{8'd160,8'd70} : s = 230;
	{8'd160,8'd71} : s = 231;
	{8'd160,8'd72} : s = 232;
	{8'd160,8'd73} : s = 233;
	{8'd160,8'd74} : s = 234;
	{8'd160,8'd75} : s = 235;
	{8'd160,8'd76} : s = 236;
	{8'd160,8'd77} : s = 237;
	{8'd160,8'd78} : s = 238;
	{8'd160,8'd79} : s = 239;
	{8'd160,8'd80} : s = 240;
	{8'd160,8'd81} : s = 241;
	{8'd160,8'd82} : s = 242;
	{8'd160,8'd83} : s = 243;
	{8'd160,8'd84} : s = 244;
	{8'd160,8'd85} : s = 245;
	{8'd160,8'd86} : s = 246;
	{8'd160,8'd87} : s = 247;
	{8'd160,8'd88} : s = 248;
	{8'd160,8'd89} : s = 249;
	{8'd160,8'd90} : s = 250;
	{8'd160,8'd91} : s = 251;
	{8'd160,8'd92} : s = 252;
	{8'd160,8'd93} : s = 253;
	{8'd160,8'd94} : s = 254;
	{8'd160,8'd95} : s = 255;
	{8'd160,8'd96} : s = 256;
	{8'd160,8'd97} : s = 257;
	{8'd160,8'd98} : s = 258;
	{8'd160,8'd99} : s = 259;
	{8'd160,8'd100} : s = 260;
	{8'd160,8'd101} : s = 261;
	{8'd160,8'd102} : s = 262;
	{8'd160,8'd103} : s = 263;
	{8'd160,8'd104} : s = 264;
	{8'd160,8'd105} : s = 265;
	{8'd160,8'd106} : s = 266;
	{8'd160,8'd107} : s = 267;
	{8'd160,8'd108} : s = 268;
	{8'd160,8'd109} : s = 269;
	{8'd160,8'd110} : s = 270;
	{8'd160,8'd111} : s = 271;
	{8'd160,8'd112} : s = 272;
	{8'd160,8'd113} : s = 273;
	{8'd160,8'd114} : s = 274;
	{8'd160,8'd115} : s = 275;
	{8'd160,8'd116} : s = 276;
	{8'd160,8'd117} : s = 277;
	{8'd160,8'd118} : s = 278;
	{8'd160,8'd119} : s = 279;
	{8'd160,8'd120} : s = 280;
	{8'd160,8'd121} : s = 281;
	{8'd160,8'd122} : s = 282;
	{8'd160,8'd123} : s = 283;
	{8'd160,8'd124} : s = 284;
	{8'd160,8'd125} : s = 285;
	{8'd160,8'd126} : s = 286;
	{8'd160,8'd127} : s = 287;
	{8'd160,8'd128} : s = 288;
	{8'd160,8'd129} : s = 289;
	{8'd160,8'd130} : s = 290;
	{8'd160,8'd131} : s = 291;
	{8'd160,8'd132} : s = 292;
	{8'd160,8'd133} : s = 293;
	{8'd160,8'd134} : s = 294;
	{8'd160,8'd135} : s = 295;
	{8'd160,8'd136} : s = 296;
	{8'd160,8'd137} : s = 297;
	{8'd160,8'd138} : s = 298;
	{8'd160,8'd139} : s = 299;
	{8'd160,8'd140} : s = 300;
	{8'd160,8'd141} : s = 301;
	{8'd160,8'd142} : s = 302;
	{8'd160,8'd143} : s = 303;
	{8'd160,8'd144} : s = 304;
	{8'd160,8'd145} : s = 305;
	{8'd160,8'd146} : s = 306;
	{8'd160,8'd147} : s = 307;
	{8'd160,8'd148} : s = 308;
	{8'd160,8'd149} : s = 309;
	{8'd160,8'd150} : s = 310;
	{8'd160,8'd151} : s = 311;
	{8'd160,8'd152} : s = 312;
	{8'd160,8'd153} : s = 313;
	{8'd160,8'd154} : s = 314;
	{8'd160,8'd155} : s = 315;
	{8'd160,8'd156} : s = 316;
	{8'd160,8'd157} : s = 317;
	{8'd160,8'd158} : s = 318;
	{8'd160,8'd159} : s = 319;
	{8'd160,8'd160} : s = 320;
	{8'd160,8'd161} : s = 321;
	{8'd160,8'd162} : s = 322;
	{8'd160,8'd163} : s = 323;
	{8'd160,8'd164} : s = 324;
	{8'd160,8'd165} : s = 325;
	{8'd160,8'd166} : s = 326;
	{8'd160,8'd167} : s = 327;
	{8'd160,8'd168} : s = 328;
	{8'd160,8'd169} : s = 329;
	{8'd160,8'd170} : s = 330;
	{8'd160,8'd171} : s = 331;
	{8'd160,8'd172} : s = 332;
	{8'd160,8'd173} : s = 333;
	{8'd160,8'd174} : s = 334;
	{8'd160,8'd175} : s = 335;
	{8'd160,8'd176} : s = 336;
	{8'd160,8'd177} : s = 337;
	{8'd160,8'd178} : s = 338;
	{8'd160,8'd179} : s = 339;
	{8'd160,8'd180} : s = 340;
	{8'd160,8'd181} : s = 341;
	{8'd160,8'd182} : s = 342;
	{8'd160,8'd183} : s = 343;
	{8'd160,8'd184} : s = 344;
	{8'd160,8'd185} : s = 345;
	{8'd160,8'd186} : s = 346;
	{8'd160,8'd187} : s = 347;
	{8'd160,8'd188} : s = 348;
	{8'd160,8'd189} : s = 349;
	{8'd160,8'd190} : s = 350;
	{8'd160,8'd191} : s = 351;
	{8'd160,8'd192} : s = 352;
	{8'd160,8'd193} : s = 353;
	{8'd160,8'd194} : s = 354;
	{8'd160,8'd195} : s = 355;
	{8'd160,8'd196} : s = 356;
	{8'd160,8'd197} : s = 357;
	{8'd160,8'd198} : s = 358;
	{8'd160,8'd199} : s = 359;
	{8'd160,8'd200} : s = 360;
	{8'd160,8'd201} : s = 361;
	{8'd160,8'd202} : s = 362;
	{8'd160,8'd203} : s = 363;
	{8'd160,8'd204} : s = 364;
	{8'd160,8'd205} : s = 365;
	{8'd160,8'd206} : s = 366;
	{8'd160,8'd207} : s = 367;
	{8'd160,8'd208} : s = 368;
	{8'd160,8'd209} : s = 369;
	{8'd160,8'd210} : s = 370;
	{8'd160,8'd211} : s = 371;
	{8'd160,8'd212} : s = 372;
	{8'd160,8'd213} : s = 373;
	{8'd160,8'd214} : s = 374;
	{8'd160,8'd215} : s = 375;
	{8'd160,8'd216} : s = 376;
	{8'd160,8'd217} : s = 377;
	{8'd160,8'd218} : s = 378;
	{8'd160,8'd219} : s = 379;
	{8'd160,8'd220} : s = 380;
	{8'd160,8'd221} : s = 381;
	{8'd160,8'd222} : s = 382;
	{8'd160,8'd223} : s = 383;
	{8'd160,8'd224} : s = 384;
	{8'd160,8'd225} : s = 385;
	{8'd160,8'd226} : s = 386;
	{8'd160,8'd227} : s = 387;
	{8'd160,8'd228} : s = 388;
	{8'd160,8'd229} : s = 389;
	{8'd160,8'd230} : s = 390;
	{8'd160,8'd231} : s = 391;
	{8'd160,8'd232} : s = 392;
	{8'd160,8'd233} : s = 393;
	{8'd160,8'd234} : s = 394;
	{8'd160,8'd235} : s = 395;
	{8'd160,8'd236} : s = 396;
	{8'd160,8'd237} : s = 397;
	{8'd160,8'd238} : s = 398;
	{8'd160,8'd239} : s = 399;
	{8'd160,8'd240} : s = 400;
	{8'd160,8'd241} : s = 401;
	{8'd160,8'd242} : s = 402;
	{8'd160,8'd243} : s = 403;
	{8'd160,8'd244} : s = 404;
	{8'd160,8'd245} : s = 405;
	{8'd160,8'd246} : s = 406;
	{8'd160,8'd247} : s = 407;
	{8'd160,8'd248} : s = 408;
	{8'd160,8'd249} : s = 409;
	{8'd160,8'd250} : s = 410;
	{8'd160,8'd251} : s = 411;
	{8'd160,8'd252} : s = 412;
	{8'd160,8'd253} : s = 413;
	{8'd160,8'd254} : s = 414;
	{8'd160,8'd255} : s = 415;
	{8'd161,8'd0} : s = 161;
	{8'd161,8'd1} : s = 162;
	{8'd161,8'd2} : s = 163;
	{8'd161,8'd3} : s = 164;
	{8'd161,8'd4} : s = 165;
	{8'd161,8'd5} : s = 166;
	{8'd161,8'd6} : s = 167;
	{8'd161,8'd7} : s = 168;
	{8'd161,8'd8} : s = 169;
	{8'd161,8'd9} : s = 170;
	{8'd161,8'd10} : s = 171;
	{8'd161,8'd11} : s = 172;
	{8'd161,8'd12} : s = 173;
	{8'd161,8'd13} : s = 174;
	{8'd161,8'd14} : s = 175;
	{8'd161,8'd15} : s = 176;
	{8'd161,8'd16} : s = 177;
	{8'd161,8'd17} : s = 178;
	{8'd161,8'd18} : s = 179;
	{8'd161,8'd19} : s = 180;
	{8'd161,8'd20} : s = 181;
	{8'd161,8'd21} : s = 182;
	{8'd161,8'd22} : s = 183;
	{8'd161,8'd23} : s = 184;
	{8'd161,8'd24} : s = 185;
	{8'd161,8'd25} : s = 186;
	{8'd161,8'd26} : s = 187;
	{8'd161,8'd27} : s = 188;
	{8'd161,8'd28} : s = 189;
	{8'd161,8'd29} : s = 190;
	{8'd161,8'd30} : s = 191;
	{8'd161,8'd31} : s = 192;
	{8'd161,8'd32} : s = 193;
	{8'd161,8'd33} : s = 194;
	{8'd161,8'd34} : s = 195;
	{8'd161,8'd35} : s = 196;
	{8'd161,8'd36} : s = 197;
	{8'd161,8'd37} : s = 198;
	{8'd161,8'd38} : s = 199;
	{8'd161,8'd39} : s = 200;
	{8'd161,8'd40} : s = 201;
	{8'd161,8'd41} : s = 202;
	{8'd161,8'd42} : s = 203;
	{8'd161,8'd43} : s = 204;
	{8'd161,8'd44} : s = 205;
	{8'd161,8'd45} : s = 206;
	{8'd161,8'd46} : s = 207;
	{8'd161,8'd47} : s = 208;
	{8'd161,8'd48} : s = 209;
	{8'd161,8'd49} : s = 210;
	{8'd161,8'd50} : s = 211;
	{8'd161,8'd51} : s = 212;
	{8'd161,8'd52} : s = 213;
	{8'd161,8'd53} : s = 214;
	{8'd161,8'd54} : s = 215;
	{8'd161,8'd55} : s = 216;
	{8'd161,8'd56} : s = 217;
	{8'd161,8'd57} : s = 218;
	{8'd161,8'd58} : s = 219;
	{8'd161,8'd59} : s = 220;
	{8'd161,8'd60} : s = 221;
	{8'd161,8'd61} : s = 222;
	{8'd161,8'd62} : s = 223;
	{8'd161,8'd63} : s = 224;
	{8'd161,8'd64} : s = 225;
	{8'd161,8'd65} : s = 226;
	{8'd161,8'd66} : s = 227;
	{8'd161,8'd67} : s = 228;
	{8'd161,8'd68} : s = 229;
	{8'd161,8'd69} : s = 230;
	{8'd161,8'd70} : s = 231;
	{8'd161,8'd71} : s = 232;
	{8'd161,8'd72} : s = 233;
	{8'd161,8'd73} : s = 234;
	{8'd161,8'd74} : s = 235;
	{8'd161,8'd75} : s = 236;
	{8'd161,8'd76} : s = 237;
	{8'd161,8'd77} : s = 238;
	{8'd161,8'd78} : s = 239;
	{8'd161,8'd79} : s = 240;
	{8'd161,8'd80} : s = 241;
	{8'd161,8'd81} : s = 242;
	{8'd161,8'd82} : s = 243;
	{8'd161,8'd83} : s = 244;
	{8'd161,8'd84} : s = 245;
	{8'd161,8'd85} : s = 246;
	{8'd161,8'd86} : s = 247;
	{8'd161,8'd87} : s = 248;
	{8'd161,8'd88} : s = 249;
	{8'd161,8'd89} : s = 250;
	{8'd161,8'd90} : s = 251;
	{8'd161,8'd91} : s = 252;
	{8'd161,8'd92} : s = 253;
	{8'd161,8'd93} : s = 254;
	{8'd161,8'd94} : s = 255;
	{8'd161,8'd95} : s = 256;
	{8'd161,8'd96} : s = 257;
	{8'd161,8'd97} : s = 258;
	{8'd161,8'd98} : s = 259;
	{8'd161,8'd99} : s = 260;
	{8'd161,8'd100} : s = 261;
	{8'd161,8'd101} : s = 262;
	{8'd161,8'd102} : s = 263;
	{8'd161,8'd103} : s = 264;
	{8'd161,8'd104} : s = 265;
	{8'd161,8'd105} : s = 266;
	{8'd161,8'd106} : s = 267;
	{8'd161,8'd107} : s = 268;
	{8'd161,8'd108} : s = 269;
	{8'd161,8'd109} : s = 270;
	{8'd161,8'd110} : s = 271;
	{8'd161,8'd111} : s = 272;
	{8'd161,8'd112} : s = 273;
	{8'd161,8'd113} : s = 274;
	{8'd161,8'd114} : s = 275;
	{8'd161,8'd115} : s = 276;
	{8'd161,8'd116} : s = 277;
	{8'd161,8'd117} : s = 278;
	{8'd161,8'd118} : s = 279;
	{8'd161,8'd119} : s = 280;
	{8'd161,8'd120} : s = 281;
	{8'd161,8'd121} : s = 282;
	{8'd161,8'd122} : s = 283;
	{8'd161,8'd123} : s = 284;
	{8'd161,8'd124} : s = 285;
	{8'd161,8'd125} : s = 286;
	{8'd161,8'd126} : s = 287;
	{8'd161,8'd127} : s = 288;
	{8'd161,8'd128} : s = 289;
	{8'd161,8'd129} : s = 290;
	{8'd161,8'd130} : s = 291;
	{8'd161,8'd131} : s = 292;
	{8'd161,8'd132} : s = 293;
	{8'd161,8'd133} : s = 294;
	{8'd161,8'd134} : s = 295;
	{8'd161,8'd135} : s = 296;
	{8'd161,8'd136} : s = 297;
	{8'd161,8'd137} : s = 298;
	{8'd161,8'd138} : s = 299;
	{8'd161,8'd139} : s = 300;
	{8'd161,8'd140} : s = 301;
	{8'd161,8'd141} : s = 302;
	{8'd161,8'd142} : s = 303;
	{8'd161,8'd143} : s = 304;
	{8'd161,8'd144} : s = 305;
	{8'd161,8'd145} : s = 306;
	{8'd161,8'd146} : s = 307;
	{8'd161,8'd147} : s = 308;
	{8'd161,8'd148} : s = 309;
	{8'd161,8'd149} : s = 310;
	{8'd161,8'd150} : s = 311;
	{8'd161,8'd151} : s = 312;
	{8'd161,8'd152} : s = 313;
	{8'd161,8'd153} : s = 314;
	{8'd161,8'd154} : s = 315;
	{8'd161,8'd155} : s = 316;
	{8'd161,8'd156} : s = 317;
	{8'd161,8'd157} : s = 318;
	{8'd161,8'd158} : s = 319;
	{8'd161,8'd159} : s = 320;
	{8'd161,8'd160} : s = 321;
	{8'd161,8'd161} : s = 322;
	{8'd161,8'd162} : s = 323;
	{8'd161,8'd163} : s = 324;
	{8'd161,8'd164} : s = 325;
	{8'd161,8'd165} : s = 326;
	{8'd161,8'd166} : s = 327;
	{8'd161,8'd167} : s = 328;
	{8'd161,8'd168} : s = 329;
	{8'd161,8'd169} : s = 330;
	{8'd161,8'd170} : s = 331;
	{8'd161,8'd171} : s = 332;
	{8'd161,8'd172} : s = 333;
	{8'd161,8'd173} : s = 334;
	{8'd161,8'd174} : s = 335;
	{8'd161,8'd175} : s = 336;
	{8'd161,8'd176} : s = 337;
	{8'd161,8'd177} : s = 338;
	{8'd161,8'd178} : s = 339;
	{8'd161,8'd179} : s = 340;
	{8'd161,8'd180} : s = 341;
	{8'd161,8'd181} : s = 342;
	{8'd161,8'd182} : s = 343;
	{8'd161,8'd183} : s = 344;
	{8'd161,8'd184} : s = 345;
	{8'd161,8'd185} : s = 346;
	{8'd161,8'd186} : s = 347;
	{8'd161,8'd187} : s = 348;
	{8'd161,8'd188} : s = 349;
	{8'd161,8'd189} : s = 350;
	{8'd161,8'd190} : s = 351;
	{8'd161,8'd191} : s = 352;
	{8'd161,8'd192} : s = 353;
	{8'd161,8'd193} : s = 354;
	{8'd161,8'd194} : s = 355;
	{8'd161,8'd195} : s = 356;
	{8'd161,8'd196} : s = 357;
	{8'd161,8'd197} : s = 358;
	{8'd161,8'd198} : s = 359;
	{8'd161,8'd199} : s = 360;
	{8'd161,8'd200} : s = 361;
	{8'd161,8'd201} : s = 362;
	{8'd161,8'd202} : s = 363;
	{8'd161,8'd203} : s = 364;
	{8'd161,8'd204} : s = 365;
	{8'd161,8'd205} : s = 366;
	{8'd161,8'd206} : s = 367;
	{8'd161,8'd207} : s = 368;
	{8'd161,8'd208} : s = 369;
	{8'd161,8'd209} : s = 370;
	{8'd161,8'd210} : s = 371;
	{8'd161,8'd211} : s = 372;
	{8'd161,8'd212} : s = 373;
	{8'd161,8'd213} : s = 374;
	{8'd161,8'd214} : s = 375;
	{8'd161,8'd215} : s = 376;
	{8'd161,8'd216} : s = 377;
	{8'd161,8'd217} : s = 378;
	{8'd161,8'd218} : s = 379;
	{8'd161,8'd219} : s = 380;
	{8'd161,8'd220} : s = 381;
	{8'd161,8'd221} : s = 382;
	{8'd161,8'd222} : s = 383;
	{8'd161,8'd223} : s = 384;
	{8'd161,8'd224} : s = 385;
	{8'd161,8'd225} : s = 386;
	{8'd161,8'd226} : s = 387;
	{8'd161,8'd227} : s = 388;
	{8'd161,8'd228} : s = 389;
	{8'd161,8'd229} : s = 390;
	{8'd161,8'd230} : s = 391;
	{8'd161,8'd231} : s = 392;
	{8'd161,8'd232} : s = 393;
	{8'd161,8'd233} : s = 394;
	{8'd161,8'd234} : s = 395;
	{8'd161,8'd235} : s = 396;
	{8'd161,8'd236} : s = 397;
	{8'd161,8'd237} : s = 398;
	{8'd161,8'd238} : s = 399;
	{8'd161,8'd239} : s = 400;
	{8'd161,8'd240} : s = 401;
	{8'd161,8'd241} : s = 402;
	{8'd161,8'd242} : s = 403;
	{8'd161,8'd243} : s = 404;
	{8'd161,8'd244} : s = 405;
	{8'd161,8'd245} : s = 406;
	{8'd161,8'd246} : s = 407;
	{8'd161,8'd247} : s = 408;
	{8'd161,8'd248} : s = 409;
	{8'd161,8'd249} : s = 410;
	{8'd161,8'd250} : s = 411;
	{8'd161,8'd251} : s = 412;
	{8'd161,8'd252} : s = 413;
	{8'd161,8'd253} : s = 414;
	{8'd161,8'd254} : s = 415;
	{8'd161,8'd255} : s = 416;
	{8'd162,8'd0} : s = 162;
	{8'd162,8'd1} : s = 163;
	{8'd162,8'd2} : s = 164;
	{8'd162,8'd3} : s = 165;
	{8'd162,8'd4} : s = 166;
	{8'd162,8'd5} : s = 167;
	{8'd162,8'd6} : s = 168;
	{8'd162,8'd7} : s = 169;
	{8'd162,8'd8} : s = 170;
	{8'd162,8'd9} : s = 171;
	{8'd162,8'd10} : s = 172;
	{8'd162,8'd11} : s = 173;
	{8'd162,8'd12} : s = 174;
	{8'd162,8'd13} : s = 175;
	{8'd162,8'd14} : s = 176;
	{8'd162,8'd15} : s = 177;
	{8'd162,8'd16} : s = 178;
	{8'd162,8'd17} : s = 179;
	{8'd162,8'd18} : s = 180;
	{8'd162,8'd19} : s = 181;
	{8'd162,8'd20} : s = 182;
	{8'd162,8'd21} : s = 183;
	{8'd162,8'd22} : s = 184;
	{8'd162,8'd23} : s = 185;
	{8'd162,8'd24} : s = 186;
	{8'd162,8'd25} : s = 187;
	{8'd162,8'd26} : s = 188;
	{8'd162,8'd27} : s = 189;
	{8'd162,8'd28} : s = 190;
	{8'd162,8'd29} : s = 191;
	{8'd162,8'd30} : s = 192;
	{8'd162,8'd31} : s = 193;
	{8'd162,8'd32} : s = 194;
	{8'd162,8'd33} : s = 195;
	{8'd162,8'd34} : s = 196;
	{8'd162,8'd35} : s = 197;
	{8'd162,8'd36} : s = 198;
	{8'd162,8'd37} : s = 199;
	{8'd162,8'd38} : s = 200;
	{8'd162,8'd39} : s = 201;
	{8'd162,8'd40} : s = 202;
	{8'd162,8'd41} : s = 203;
	{8'd162,8'd42} : s = 204;
	{8'd162,8'd43} : s = 205;
	{8'd162,8'd44} : s = 206;
	{8'd162,8'd45} : s = 207;
	{8'd162,8'd46} : s = 208;
	{8'd162,8'd47} : s = 209;
	{8'd162,8'd48} : s = 210;
	{8'd162,8'd49} : s = 211;
	{8'd162,8'd50} : s = 212;
	{8'd162,8'd51} : s = 213;
	{8'd162,8'd52} : s = 214;
	{8'd162,8'd53} : s = 215;
	{8'd162,8'd54} : s = 216;
	{8'd162,8'd55} : s = 217;
	{8'd162,8'd56} : s = 218;
	{8'd162,8'd57} : s = 219;
	{8'd162,8'd58} : s = 220;
	{8'd162,8'd59} : s = 221;
	{8'd162,8'd60} : s = 222;
	{8'd162,8'd61} : s = 223;
	{8'd162,8'd62} : s = 224;
	{8'd162,8'd63} : s = 225;
	{8'd162,8'd64} : s = 226;
	{8'd162,8'd65} : s = 227;
	{8'd162,8'd66} : s = 228;
	{8'd162,8'd67} : s = 229;
	{8'd162,8'd68} : s = 230;
	{8'd162,8'd69} : s = 231;
	{8'd162,8'd70} : s = 232;
	{8'd162,8'd71} : s = 233;
	{8'd162,8'd72} : s = 234;
	{8'd162,8'd73} : s = 235;
	{8'd162,8'd74} : s = 236;
	{8'd162,8'd75} : s = 237;
	{8'd162,8'd76} : s = 238;
	{8'd162,8'd77} : s = 239;
	{8'd162,8'd78} : s = 240;
	{8'd162,8'd79} : s = 241;
	{8'd162,8'd80} : s = 242;
	{8'd162,8'd81} : s = 243;
	{8'd162,8'd82} : s = 244;
	{8'd162,8'd83} : s = 245;
	{8'd162,8'd84} : s = 246;
	{8'd162,8'd85} : s = 247;
	{8'd162,8'd86} : s = 248;
	{8'd162,8'd87} : s = 249;
	{8'd162,8'd88} : s = 250;
	{8'd162,8'd89} : s = 251;
	{8'd162,8'd90} : s = 252;
	{8'd162,8'd91} : s = 253;
	{8'd162,8'd92} : s = 254;
	{8'd162,8'd93} : s = 255;
	{8'd162,8'd94} : s = 256;
	{8'd162,8'd95} : s = 257;
	{8'd162,8'd96} : s = 258;
	{8'd162,8'd97} : s = 259;
	{8'd162,8'd98} : s = 260;
	{8'd162,8'd99} : s = 261;
	{8'd162,8'd100} : s = 262;
	{8'd162,8'd101} : s = 263;
	{8'd162,8'd102} : s = 264;
	{8'd162,8'd103} : s = 265;
	{8'd162,8'd104} : s = 266;
	{8'd162,8'd105} : s = 267;
	{8'd162,8'd106} : s = 268;
	{8'd162,8'd107} : s = 269;
	{8'd162,8'd108} : s = 270;
	{8'd162,8'd109} : s = 271;
	{8'd162,8'd110} : s = 272;
	{8'd162,8'd111} : s = 273;
	{8'd162,8'd112} : s = 274;
	{8'd162,8'd113} : s = 275;
	{8'd162,8'd114} : s = 276;
	{8'd162,8'd115} : s = 277;
	{8'd162,8'd116} : s = 278;
	{8'd162,8'd117} : s = 279;
	{8'd162,8'd118} : s = 280;
	{8'd162,8'd119} : s = 281;
	{8'd162,8'd120} : s = 282;
	{8'd162,8'd121} : s = 283;
	{8'd162,8'd122} : s = 284;
	{8'd162,8'd123} : s = 285;
	{8'd162,8'd124} : s = 286;
	{8'd162,8'd125} : s = 287;
	{8'd162,8'd126} : s = 288;
	{8'd162,8'd127} : s = 289;
	{8'd162,8'd128} : s = 290;
	{8'd162,8'd129} : s = 291;
	{8'd162,8'd130} : s = 292;
	{8'd162,8'd131} : s = 293;
	{8'd162,8'd132} : s = 294;
	{8'd162,8'd133} : s = 295;
	{8'd162,8'd134} : s = 296;
	{8'd162,8'd135} : s = 297;
	{8'd162,8'd136} : s = 298;
	{8'd162,8'd137} : s = 299;
	{8'd162,8'd138} : s = 300;
	{8'd162,8'd139} : s = 301;
	{8'd162,8'd140} : s = 302;
	{8'd162,8'd141} : s = 303;
	{8'd162,8'd142} : s = 304;
	{8'd162,8'd143} : s = 305;
	{8'd162,8'd144} : s = 306;
	{8'd162,8'd145} : s = 307;
	{8'd162,8'd146} : s = 308;
	{8'd162,8'd147} : s = 309;
	{8'd162,8'd148} : s = 310;
	{8'd162,8'd149} : s = 311;
	{8'd162,8'd150} : s = 312;
	{8'd162,8'd151} : s = 313;
	{8'd162,8'd152} : s = 314;
	{8'd162,8'd153} : s = 315;
	{8'd162,8'd154} : s = 316;
	{8'd162,8'd155} : s = 317;
	{8'd162,8'd156} : s = 318;
	{8'd162,8'd157} : s = 319;
	{8'd162,8'd158} : s = 320;
	{8'd162,8'd159} : s = 321;
	{8'd162,8'd160} : s = 322;
	{8'd162,8'd161} : s = 323;
	{8'd162,8'd162} : s = 324;
	{8'd162,8'd163} : s = 325;
	{8'd162,8'd164} : s = 326;
	{8'd162,8'd165} : s = 327;
	{8'd162,8'd166} : s = 328;
	{8'd162,8'd167} : s = 329;
	{8'd162,8'd168} : s = 330;
	{8'd162,8'd169} : s = 331;
	{8'd162,8'd170} : s = 332;
	{8'd162,8'd171} : s = 333;
	{8'd162,8'd172} : s = 334;
	{8'd162,8'd173} : s = 335;
	{8'd162,8'd174} : s = 336;
	{8'd162,8'd175} : s = 337;
	{8'd162,8'd176} : s = 338;
	{8'd162,8'd177} : s = 339;
	{8'd162,8'd178} : s = 340;
	{8'd162,8'd179} : s = 341;
	{8'd162,8'd180} : s = 342;
	{8'd162,8'd181} : s = 343;
	{8'd162,8'd182} : s = 344;
	{8'd162,8'd183} : s = 345;
	{8'd162,8'd184} : s = 346;
	{8'd162,8'd185} : s = 347;
	{8'd162,8'd186} : s = 348;
	{8'd162,8'd187} : s = 349;
	{8'd162,8'd188} : s = 350;
	{8'd162,8'd189} : s = 351;
	{8'd162,8'd190} : s = 352;
	{8'd162,8'd191} : s = 353;
	{8'd162,8'd192} : s = 354;
	{8'd162,8'd193} : s = 355;
	{8'd162,8'd194} : s = 356;
	{8'd162,8'd195} : s = 357;
	{8'd162,8'd196} : s = 358;
	{8'd162,8'd197} : s = 359;
	{8'd162,8'd198} : s = 360;
	{8'd162,8'd199} : s = 361;
	{8'd162,8'd200} : s = 362;
	{8'd162,8'd201} : s = 363;
	{8'd162,8'd202} : s = 364;
	{8'd162,8'd203} : s = 365;
	{8'd162,8'd204} : s = 366;
	{8'd162,8'd205} : s = 367;
	{8'd162,8'd206} : s = 368;
	{8'd162,8'd207} : s = 369;
	{8'd162,8'd208} : s = 370;
	{8'd162,8'd209} : s = 371;
	{8'd162,8'd210} : s = 372;
	{8'd162,8'd211} : s = 373;
	{8'd162,8'd212} : s = 374;
	{8'd162,8'd213} : s = 375;
	{8'd162,8'd214} : s = 376;
	{8'd162,8'd215} : s = 377;
	{8'd162,8'd216} : s = 378;
	{8'd162,8'd217} : s = 379;
	{8'd162,8'd218} : s = 380;
	{8'd162,8'd219} : s = 381;
	{8'd162,8'd220} : s = 382;
	{8'd162,8'd221} : s = 383;
	{8'd162,8'd222} : s = 384;
	{8'd162,8'd223} : s = 385;
	{8'd162,8'd224} : s = 386;
	{8'd162,8'd225} : s = 387;
	{8'd162,8'd226} : s = 388;
	{8'd162,8'd227} : s = 389;
	{8'd162,8'd228} : s = 390;
	{8'd162,8'd229} : s = 391;
	{8'd162,8'd230} : s = 392;
	{8'd162,8'd231} : s = 393;
	{8'd162,8'd232} : s = 394;
	{8'd162,8'd233} : s = 395;
	{8'd162,8'd234} : s = 396;
	{8'd162,8'd235} : s = 397;
	{8'd162,8'd236} : s = 398;
	{8'd162,8'd237} : s = 399;
	{8'd162,8'd238} : s = 400;
	{8'd162,8'd239} : s = 401;
	{8'd162,8'd240} : s = 402;
	{8'd162,8'd241} : s = 403;
	{8'd162,8'd242} : s = 404;
	{8'd162,8'd243} : s = 405;
	{8'd162,8'd244} : s = 406;
	{8'd162,8'd245} : s = 407;
	{8'd162,8'd246} : s = 408;
	{8'd162,8'd247} : s = 409;
	{8'd162,8'd248} : s = 410;
	{8'd162,8'd249} : s = 411;
	{8'd162,8'd250} : s = 412;
	{8'd162,8'd251} : s = 413;
	{8'd162,8'd252} : s = 414;
	{8'd162,8'd253} : s = 415;
	{8'd162,8'd254} : s = 416;
	{8'd162,8'd255} : s = 417;
	{8'd163,8'd0} : s = 163;
	{8'd163,8'd1} : s = 164;
	{8'd163,8'd2} : s = 165;
	{8'd163,8'd3} : s = 166;
	{8'd163,8'd4} : s = 167;
	{8'd163,8'd5} : s = 168;
	{8'd163,8'd6} : s = 169;
	{8'd163,8'd7} : s = 170;
	{8'd163,8'd8} : s = 171;
	{8'd163,8'd9} : s = 172;
	{8'd163,8'd10} : s = 173;
	{8'd163,8'd11} : s = 174;
	{8'd163,8'd12} : s = 175;
	{8'd163,8'd13} : s = 176;
	{8'd163,8'd14} : s = 177;
	{8'd163,8'd15} : s = 178;
	{8'd163,8'd16} : s = 179;
	{8'd163,8'd17} : s = 180;
	{8'd163,8'd18} : s = 181;
	{8'd163,8'd19} : s = 182;
	{8'd163,8'd20} : s = 183;
	{8'd163,8'd21} : s = 184;
	{8'd163,8'd22} : s = 185;
	{8'd163,8'd23} : s = 186;
	{8'd163,8'd24} : s = 187;
	{8'd163,8'd25} : s = 188;
	{8'd163,8'd26} : s = 189;
	{8'd163,8'd27} : s = 190;
	{8'd163,8'd28} : s = 191;
	{8'd163,8'd29} : s = 192;
	{8'd163,8'd30} : s = 193;
	{8'd163,8'd31} : s = 194;
	{8'd163,8'd32} : s = 195;
	{8'd163,8'd33} : s = 196;
	{8'd163,8'd34} : s = 197;
	{8'd163,8'd35} : s = 198;
	{8'd163,8'd36} : s = 199;
	{8'd163,8'd37} : s = 200;
	{8'd163,8'd38} : s = 201;
	{8'd163,8'd39} : s = 202;
	{8'd163,8'd40} : s = 203;
	{8'd163,8'd41} : s = 204;
	{8'd163,8'd42} : s = 205;
	{8'd163,8'd43} : s = 206;
	{8'd163,8'd44} : s = 207;
	{8'd163,8'd45} : s = 208;
	{8'd163,8'd46} : s = 209;
	{8'd163,8'd47} : s = 210;
	{8'd163,8'd48} : s = 211;
	{8'd163,8'd49} : s = 212;
	{8'd163,8'd50} : s = 213;
	{8'd163,8'd51} : s = 214;
	{8'd163,8'd52} : s = 215;
	{8'd163,8'd53} : s = 216;
	{8'd163,8'd54} : s = 217;
	{8'd163,8'd55} : s = 218;
	{8'd163,8'd56} : s = 219;
	{8'd163,8'd57} : s = 220;
	{8'd163,8'd58} : s = 221;
	{8'd163,8'd59} : s = 222;
	{8'd163,8'd60} : s = 223;
	{8'd163,8'd61} : s = 224;
	{8'd163,8'd62} : s = 225;
	{8'd163,8'd63} : s = 226;
	{8'd163,8'd64} : s = 227;
	{8'd163,8'd65} : s = 228;
	{8'd163,8'd66} : s = 229;
	{8'd163,8'd67} : s = 230;
	{8'd163,8'd68} : s = 231;
	{8'd163,8'd69} : s = 232;
	{8'd163,8'd70} : s = 233;
	{8'd163,8'd71} : s = 234;
	{8'd163,8'd72} : s = 235;
	{8'd163,8'd73} : s = 236;
	{8'd163,8'd74} : s = 237;
	{8'd163,8'd75} : s = 238;
	{8'd163,8'd76} : s = 239;
	{8'd163,8'd77} : s = 240;
	{8'd163,8'd78} : s = 241;
	{8'd163,8'd79} : s = 242;
	{8'd163,8'd80} : s = 243;
	{8'd163,8'd81} : s = 244;
	{8'd163,8'd82} : s = 245;
	{8'd163,8'd83} : s = 246;
	{8'd163,8'd84} : s = 247;
	{8'd163,8'd85} : s = 248;
	{8'd163,8'd86} : s = 249;
	{8'd163,8'd87} : s = 250;
	{8'd163,8'd88} : s = 251;
	{8'd163,8'd89} : s = 252;
	{8'd163,8'd90} : s = 253;
	{8'd163,8'd91} : s = 254;
	{8'd163,8'd92} : s = 255;
	{8'd163,8'd93} : s = 256;
	{8'd163,8'd94} : s = 257;
	{8'd163,8'd95} : s = 258;
	{8'd163,8'd96} : s = 259;
	{8'd163,8'd97} : s = 260;
	{8'd163,8'd98} : s = 261;
	{8'd163,8'd99} : s = 262;
	{8'd163,8'd100} : s = 263;
	{8'd163,8'd101} : s = 264;
	{8'd163,8'd102} : s = 265;
	{8'd163,8'd103} : s = 266;
	{8'd163,8'd104} : s = 267;
	{8'd163,8'd105} : s = 268;
	{8'd163,8'd106} : s = 269;
	{8'd163,8'd107} : s = 270;
	{8'd163,8'd108} : s = 271;
	{8'd163,8'd109} : s = 272;
	{8'd163,8'd110} : s = 273;
	{8'd163,8'd111} : s = 274;
	{8'd163,8'd112} : s = 275;
	{8'd163,8'd113} : s = 276;
	{8'd163,8'd114} : s = 277;
	{8'd163,8'd115} : s = 278;
	{8'd163,8'd116} : s = 279;
	{8'd163,8'd117} : s = 280;
	{8'd163,8'd118} : s = 281;
	{8'd163,8'd119} : s = 282;
	{8'd163,8'd120} : s = 283;
	{8'd163,8'd121} : s = 284;
	{8'd163,8'd122} : s = 285;
	{8'd163,8'd123} : s = 286;
	{8'd163,8'd124} : s = 287;
	{8'd163,8'd125} : s = 288;
	{8'd163,8'd126} : s = 289;
	{8'd163,8'd127} : s = 290;
	{8'd163,8'd128} : s = 291;
	{8'd163,8'd129} : s = 292;
	{8'd163,8'd130} : s = 293;
	{8'd163,8'd131} : s = 294;
	{8'd163,8'd132} : s = 295;
	{8'd163,8'd133} : s = 296;
	{8'd163,8'd134} : s = 297;
	{8'd163,8'd135} : s = 298;
	{8'd163,8'd136} : s = 299;
	{8'd163,8'd137} : s = 300;
	{8'd163,8'd138} : s = 301;
	{8'd163,8'd139} : s = 302;
	{8'd163,8'd140} : s = 303;
	{8'd163,8'd141} : s = 304;
	{8'd163,8'd142} : s = 305;
	{8'd163,8'd143} : s = 306;
	{8'd163,8'd144} : s = 307;
	{8'd163,8'd145} : s = 308;
	{8'd163,8'd146} : s = 309;
	{8'd163,8'd147} : s = 310;
	{8'd163,8'd148} : s = 311;
	{8'd163,8'd149} : s = 312;
	{8'd163,8'd150} : s = 313;
	{8'd163,8'd151} : s = 314;
	{8'd163,8'd152} : s = 315;
	{8'd163,8'd153} : s = 316;
	{8'd163,8'd154} : s = 317;
	{8'd163,8'd155} : s = 318;
	{8'd163,8'd156} : s = 319;
	{8'd163,8'd157} : s = 320;
	{8'd163,8'd158} : s = 321;
	{8'd163,8'd159} : s = 322;
	{8'd163,8'd160} : s = 323;
	{8'd163,8'd161} : s = 324;
	{8'd163,8'd162} : s = 325;
	{8'd163,8'd163} : s = 326;
	{8'd163,8'd164} : s = 327;
	{8'd163,8'd165} : s = 328;
	{8'd163,8'd166} : s = 329;
	{8'd163,8'd167} : s = 330;
	{8'd163,8'd168} : s = 331;
	{8'd163,8'd169} : s = 332;
	{8'd163,8'd170} : s = 333;
	{8'd163,8'd171} : s = 334;
	{8'd163,8'd172} : s = 335;
	{8'd163,8'd173} : s = 336;
	{8'd163,8'd174} : s = 337;
	{8'd163,8'd175} : s = 338;
	{8'd163,8'd176} : s = 339;
	{8'd163,8'd177} : s = 340;
	{8'd163,8'd178} : s = 341;
	{8'd163,8'd179} : s = 342;
	{8'd163,8'd180} : s = 343;
	{8'd163,8'd181} : s = 344;
	{8'd163,8'd182} : s = 345;
	{8'd163,8'd183} : s = 346;
	{8'd163,8'd184} : s = 347;
	{8'd163,8'd185} : s = 348;
	{8'd163,8'd186} : s = 349;
	{8'd163,8'd187} : s = 350;
	{8'd163,8'd188} : s = 351;
	{8'd163,8'd189} : s = 352;
	{8'd163,8'd190} : s = 353;
	{8'd163,8'd191} : s = 354;
	{8'd163,8'd192} : s = 355;
	{8'd163,8'd193} : s = 356;
	{8'd163,8'd194} : s = 357;
	{8'd163,8'd195} : s = 358;
	{8'd163,8'd196} : s = 359;
	{8'd163,8'd197} : s = 360;
	{8'd163,8'd198} : s = 361;
	{8'd163,8'd199} : s = 362;
	{8'd163,8'd200} : s = 363;
	{8'd163,8'd201} : s = 364;
	{8'd163,8'd202} : s = 365;
	{8'd163,8'd203} : s = 366;
	{8'd163,8'd204} : s = 367;
	{8'd163,8'd205} : s = 368;
	{8'd163,8'd206} : s = 369;
	{8'd163,8'd207} : s = 370;
	{8'd163,8'd208} : s = 371;
	{8'd163,8'd209} : s = 372;
	{8'd163,8'd210} : s = 373;
	{8'd163,8'd211} : s = 374;
	{8'd163,8'd212} : s = 375;
	{8'd163,8'd213} : s = 376;
	{8'd163,8'd214} : s = 377;
	{8'd163,8'd215} : s = 378;
	{8'd163,8'd216} : s = 379;
	{8'd163,8'd217} : s = 380;
	{8'd163,8'd218} : s = 381;
	{8'd163,8'd219} : s = 382;
	{8'd163,8'd220} : s = 383;
	{8'd163,8'd221} : s = 384;
	{8'd163,8'd222} : s = 385;
	{8'd163,8'd223} : s = 386;
	{8'd163,8'd224} : s = 387;
	{8'd163,8'd225} : s = 388;
	{8'd163,8'd226} : s = 389;
	{8'd163,8'd227} : s = 390;
	{8'd163,8'd228} : s = 391;
	{8'd163,8'd229} : s = 392;
	{8'd163,8'd230} : s = 393;
	{8'd163,8'd231} : s = 394;
	{8'd163,8'd232} : s = 395;
	{8'd163,8'd233} : s = 396;
	{8'd163,8'd234} : s = 397;
	{8'd163,8'd235} : s = 398;
	{8'd163,8'd236} : s = 399;
	{8'd163,8'd237} : s = 400;
	{8'd163,8'd238} : s = 401;
	{8'd163,8'd239} : s = 402;
	{8'd163,8'd240} : s = 403;
	{8'd163,8'd241} : s = 404;
	{8'd163,8'd242} : s = 405;
	{8'd163,8'd243} : s = 406;
	{8'd163,8'd244} : s = 407;
	{8'd163,8'd245} : s = 408;
	{8'd163,8'd246} : s = 409;
	{8'd163,8'd247} : s = 410;
	{8'd163,8'd248} : s = 411;
	{8'd163,8'd249} : s = 412;
	{8'd163,8'd250} : s = 413;
	{8'd163,8'd251} : s = 414;
	{8'd163,8'd252} : s = 415;
	{8'd163,8'd253} : s = 416;
	{8'd163,8'd254} : s = 417;
	{8'd163,8'd255} : s = 418;
	{8'd164,8'd0} : s = 164;
	{8'd164,8'd1} : s = 165;
	{8'd164,8'd2} : s = 166;
	{8'd164,8'd3} : s = 167;
	{8'd164,8'd4} : s = 168;
	{8'd164,8'd5} : s = 169;
	{8'd164,8'd6} : s = 170;
	{8'd164,8'd7} : s = 171;
	{8'd164,8'd8} : s = 172;
	{8'd164,8'd9} : s = 173;
	{8'd164,8'd10} : s = 174;
	{8'd164,8'd11} : s = 175;
	{8'd164,8'd12} : s = 176;
	{8'd164,8'd13} : s = 177;
	{8'd164,8'd14} : s = 178;
	{8'd164,8'd15} : s = 179;
	{8'd164,8'd16} : s = 180;
	{8'd164,8'd17} : s = 181;
	{8'd164,8'd18} : s = 182;
	{8'd164,8'd19} : s = 183;
	{8'd164,8'd20} : s = 184;
	{8'd164,8'd21} : s = 185;
	{8'd164,8'd22} : s = 186;
	{8'd164,8'd23} : s = 187;
	{8'd164,8'd24} : s = 188;
	{8'd164,8'd25} : s = 189;
	{8'd164,8'd26} : s = 190;
	{8'd164,8'd27} : s = 191;
	{8'd164,8'd28} : s = 192;
	{8'd164,8'd29} : s = 193;
	{8'd164,8'd30} : s = 194;
	{8'd164,8'd31} : s = 195;
	{8'd164,8'd32} : s = 196;
	{8'd164,8'd33} : s = 197;
	{8'd164,8'd34} : s = 198;
	{8'd164,8'd35} : s = 199;
	{8'd164,8'd36} : s = 200;
	{8'd164,8'd37} : s = 201;
	{8'd164,8'd38} : s = 202;
	{8'd164,8'd39} : s = 203;
	{8'd164,8'd40} : s = 204;
	{8'd164,8'd41} : s = 205;
	{8'd164,8'd42} : s = 206;
	{8'd164,8'd43} : s = 207;
	{8'd164,8'd44} : s = 208;
	{8'd164,8'd45} : s = 209;
	{8'd164,8'd46} : s = 210;
	{8'd164,8'd47} : s = 211;
	{8'd164,8'd48} : s = 212;
	{8'd164,8'd49} : s = 213;
	{8'd164,8'd50} : s = 214;
	{8'd164,8'd51} : s = 215;
	{8'd164,8'd52} : s = 216;
	{8'd164,8'd53} : s = 217;
	{8'd164,8'd54} : s = 218;
	{8'd164,8'd55} : s = 219;
	{8'd164,8'd56} : s = 220;
	{8'd164,8'd57} : s = 221;
	{8'd164,8'd58} : s = 222;
	{8'd164,8'd59} : s = 223;
	{8'd164,8'd60} : s = 224;
	{8'd164,8'd61} : s = 225;
	{8'd164,8'd62} : s = 226;
	{8'd164,8'd63} : s = 227;
	{8'd164,8'd64} : s = 228;
	{8'd164,8'd65} : s = 229;
	{8'd164,8'd66} : s = 230;
	{8'd164,8'd67} : s = 231;
	{8'd164,8'd68} : s = 232;
	{8'd164,8'd69} : s = 233;
	{8'd164,8'd70} : s = 234;
	{8'd164,8'd71} : s = 235;
	{8'd164,8'd72} : s = 236;
	{8'd164,8'd73} : s = 237;
	{8'd164,8'd74} : s = 238;
	{8'd164,8'd75} : s = 239;
	{8'd164,8'd76} : s = 240;
	{8'd164,8'd77} : s = 241;
	{8'd164,8'd78} : s = 242;
	{8'd164,8'd79} : s = 243;
	{8'd164,8'd80} : s = 244;
	{8'd164,8'd81} : s = 245;
	{8'd164,8'd82} : s = 246;
	{8'd164,8'd83} : s = 247;
	{8'd164,8'd84} : s = 248;
	{8'd164,8'd85} : s = 249;
	{8'd164,8'd86} : s = 250;
	{8'd164,8'd87} : s = 251;
	{8'd164,8'd88} : s = 252;
	{8'd164,8'd89} : s = 253;
	{8'd164,8'd90} : s = 254;
	{8'd164,8'd91} : s = 255;
	{8'd164,8'd92} : s = 256;
	{8'd164,8'd93} : s = 257;
	{8'd164,8'd94} : s = 258;
	{8'd164,8'd95} : s = 259;
	{8'd164,8'd96} : s = 260;
	{8'd164,8'd97} : s = 261;
	{8'd164,8'd98} : s = 262;
	{8'd164,8'd99} : s = 263;
	{8'd164,8'd100} : s = 264;
	{8'd164,8'd101} : s = 265;
	{8'd164,8'd102} : s = 266;
	{8'd164,8'd103} : s = 267;
	{8'd164,8'd104} : s = 268;
	{8'd164,8'd105} : s = 269;
	{8'd164,8'd106} : s = 270;
	{8'd164,8'd107} : s = 271;
	{8'd164,8'd108} : s = 272;
	{8'd164,8'd109} : s = 273;
	{8'd164,8'd110} : s = 274;
	{8'd164,8'd111} : s = 275;
	{8'd164,8'd112} : s = 276;
	{8'd164,8'd113} : s = 277;
	{8'd164,8'd114} : s = 278;
	{8'd164,8'd115} : s = 279;
	{8'd164,8'd116} : s = 280;
	{8'd164,8'd117} : s = 281;
	{8'd164,8'd118} : s = 282;
	{8'd164,8'd119} : s = 283;
	{8'd164,8'd120} : s = 284;
	{8'd164,8'd121} : s = 285;
	{8'd164,8'd122} : s = 286;
	{8'd164,8'd123} : s = 287;
	{8'd164,8'd124} : s = 288;
	{8'd164,8'd125} : s = 289;
	{8'd164,8'd126} : s = 290;
	{8'd164,8'd127} : s = 291;
	{8'd164,8'd128} : s = 292;
	{8'd164,8'd129} : s = 293;
	{8'd164,8'd130} : s = 294;
	{8'd164,8'd131} : s = 295;
	{8'd164,8'd132} : s = 296;
	{8'd164,8'd133} : s = 297;
	{8'd164,8'd134} : s = 298;
	{8'd164,8'd135} : s = 299;
	{8'd164,8'd136} : s = 300;
	{8'd164,8'd137} : s = 301;
	{8'd164,8'd138} : s = 302;
	{8'd164,8'd139} : s = 303;
	{8'd164,8'd140} : s = 304;
	{8'd164,8'd141} : s = 305;
	{8'd164,8'd142} : s = 306;
	{8'd164,8'd143} : s = 307;
	{8'd164,8'd144} : s = 308;
	{8'd164,8'd145} : s = 309;
	{8'd164,8'd146} : s = 310;
	{8'd164,8'd147} : s = 311;
	{8'd164,8'd148} : s = 312;
	{8'd164,8'd149} : s = 313;
	{8'd164,8'd150} : s = 314;
	{8'd164,8'd151} : s = 315;
	{8'd164,8'd152} : s = 316;
	{8'd164,8'd153} : s = 317;
	{8'd164,8'd154} : s = 318;
	{8'd164,8'd155} : s = 319;
	{8'd164,8'd156} : s = 320;
	{8'd164,8'd157} : s = 321;
	{8'd164,8'd158} : s = 322;
	{8'd164,8'd159} : s = 323;
	{8'd164,8'd160} : s = 324;
	{8'd164,8'd161} : s = 325;
	{8'd164,8'd162} : s = 326;
	{8'd164,8'd163} : s = 327;
	{8'd164,8'd164} : s = 328;
	{8'd164,8'd165} : s = 329;
	{8'd164,8'd166} : s = 330;
	{8'd164,8'd167} : s = 331;
	{8'd164,8'd168} : s = 332;
	{8'd164,8'd169} : s = 333;
	{8'd164,8'd170} : s = 334;
	{8'd164,8'd171} : s = 335;
	{8'd164,8'd172} : s = 336;
	{8'd164,8'd173} : s = 337;
	{8'd164,8'd174} : s = 338;
	{8'd164,8'd175} : s = 339;
	{8'd164,8'd176} : s = 340;
	{8'd164,8'd177} : s = 341;
	{8'd164,8'd178} : s = 342;
	{8'd164,8'd179} : s = 343;
	{8'd164,8'd180} : s = 344;
	{8'd164,8'd181} : s = 345;
	{8'd164,8'd182} : s = 346;
	{8'd164,8'd183} : s = 347;
	{8'd164,8'd184} : s = 348;
	{8'd164,8'd185} : s = 349;
	{8'd164,8'd186} : s = 350;
	{8'd164,8'd187} : s = 351;
	{8'd164,8'd188} : s = 352;
	{8'd164,8'd189} : s = 353;
	{8'd164,8'd190} : s = 354;
	{8'd164,8'd191} : s = 355;
	{8'd164,8'd192} : s = 356;
	{8'd164,8'd193} : s = 357;
	{8'd164,8'd194} : s = 358;
	{8'd164,8'd195} : s = 359;
	{8'd164,8'd196} : s = 360;
	{8'd164,8'd197} : s = 361;
	{8'd164,8'd198} : s = 362;
	{8'd164,8'd199} : s = 363;
	{8'd164,8'd200} : s = 364;
	{8'd164,8'd201} : s = 365;
	{8'd164,8'd202} : s = 366;
	{8'd164,8'd203} : s = 367;
	{8'd164,8'd204} : s = 368;
	{8'd164,8'd205} : s = 369;
	{8'd164,8'd206} : s = 370;
	{8'd164,8'd207} : s = 371;
	{8'd164,8'd208} : s = 372;
	{8'd164,8'd209} : s = 373;
	{8'd164,8'd210} : s = 374;
	{8'd164,8'd211} : s = 375;
	{8'd164,8'd212} : s = 376;
	{8'd164,8'd213} : s = 377;
	{8'd164,8'd214} : s = 378;
	{8'd164,8'd215} : s = 379;
	{8'd164,8'd216} : s = 380;
	{8'd164,8'd217} : s = 381;
	{8'd164,8'd218} : s = 382;
	{8'd164,8'd219} : s = 383;
	{8'd164,8'd220} : s = 384;
	{8'd164,8'd221} : s = 385;
	{8'd164,8'd222} : s = 386;
	{8'd164,8'd223} : s = 387;
	{8'd164,8'd224} : s = 388;
	{8'd164,8'd225} : s = 389;
	{8'd164,8'd226} : s = 390;
	{8'd164,8'd227} : s = 391;
	{8'd164,8'd228} : s = 392;
	{8'd164,8'd229} : s = 393;
	{8'd164,8'd230} : s = 394;
	{8'd164,8'd231} : s = 395;
	{8'd164,8'd232} : s = 396;
	{8'd164,8'd233} : s = 397;
	{8'd164,8'd234} : s = 398;
	{8'd164,8'd235} : s = 399;
	{8'd164,8'd236} : s = 400;
	{8'd164,8'd237} : s = 401;
	{8'd164,8'd238} : s = 402;
	{8'd164,8'd239} : s = 403;
	{8'd164,8'd240} : s = 404;
	{8'd164,8'd241} : s = 405;
	{8'd164,8'd242} : s = 406;
	{8'd164,8'd243} : s = 407;
	{8'd164,8'd244} : s = 408;
	{8'd164,8'd245} : s = 409;
	{8'd164,8'd246} : s = 410;
	{8'd164,8'd247} : s = 411;
	{8'd164,8'd248} : s = 412;
	{8'd164,8'd249} : s = 413;
	{8'd164,8'd250} : s = 414;
	{8'd164,8'd251} : s = 415;
	{8'd164,8'd252} : s = 416;
	{8'd164,8'd253} : s = 417;
	{8'd164,8'd254} : s = 418;
	{8'd164,8'd255} : s = 419;
	{8'd165,8'd0} : s = 165;
	{8'd165,8'd1} : s = 166;
	{8'd165,8'd2} : s = 167;
	{8'd165,8'd3} : s = 168;
	{8'd165,8'd4} : s = 169;
	{8'd165,8'd5} : s = 170;
	{8'd165,8'd6} : s = 171;
	{8'd165,8'd7} : s = 172;
	{8'd165,8'd8} : s = 173;
	{8'd165,8'd9} : s = 174;
	{8'd165,8'd10} : s = 175;
	{8'd165,8'd11} : s = 176;
	{8'd165,8'd12} : s = 177;
	{8'd165,8'd13} : s = 178;
	{8'd165,8'd14} : s = 179;
	{8'd165,8'd15} : s = 180;
	{8'd165,8'd16} : s = 181;
	{8'd165,8'd17} : s = 182;
	{8'd165,8'd18} : s = 183;
	{8'd165,8'd19} : s = 184;
	{8'd165,8'd20} : s = 185;
	{8'd165,8'd21} : s = 186;
	{8'd165,8'd22} : s = 187;
	{8'd165,8'd23} : s = 188;
	{8'd165,8'd24} : s = 189;
	{8'd165,8'd25} : s = 190;
	{8'd165,8'd26} : s = 191;
	{8'd165,8'd27} : s = 192;
	{8'd165,8'd28} : s = 193;
	{8'd165,8'd29} : s = 194;
	{8'd165,8'd30} : s = 195;
	{8'd165,8'd31} : s = 196;
	{8'd165,8'd32} : s = 197;
	{8'd165,8'd33} : s = 198;
	{8'd165,8'd34} : s = 199;
	{8'd165,8'd35} : s = 200;
	{8'd165,8'd36} : s = 201;
	{8'd165,8'd37} : s = 202;
	{8'd165,8'd38} : s = 203;
	{8'd165,8'd39} : s = 204;
	{8'd165,8'd40} : s = 205;
	{8'd165,8'd41} : s = 206;
	{8'd165,8'd42} : s = 207;
	{8'd165,8'd43} : s = 208;
	{8'd165,8'd44} : s = 209;
	{8'd165,8'd45} : s = 210;
	{8'd165,8'd46} : s = 211;
	{8'd165,8'd47} : s = 212;
	{8'd165,8'd48} : s = 213;
	{8'd165,8'd49} : s = 214;
	{8'd165,8'd50} : s = 215;
	{8'd165,8'd51} : s = 216;
	{8'd165,8'd52} : s = 217;
	{8'd165,8'd53} : s = 218;
	{8'd165,8'd54} : s = 219;
	{8'd165,8'd55} : s = 220;
	{8'd165,8'd56} : s = 221;
	{8'd165,8'd57} : s = 222;
	{8'd165,8'd58} : s = 223;
	{8'd165,8'd59} : s = 224;
	{8'd165,8'd60} : s = 225;
	{8'd165,8'd61} : s = 226;
	{8'd165,8'd62} : s = 227;
	{8'd165,8'd63} : s = 228;
	{8'd165,8'd64} : s = 229;
	{8'd165,8'd65} : s = 230;
	{8'd165,8'd66} : s = 231;
	{8'd165,8'd67} : s = 232;
	{8'd165,8'd68} : s = 233;
	{8'd165,8'd69} : s = 234;
	{8'd165,8'd70} : s = 235;
	{8'd165,8'd71} : s = 236;
	{8'd165,8'd72} : s = 237;
	{8'd165,8'd73} : s = 238;
	{8'd165,8'd74} : s = 239;
	{8'd165,8'd75} : s = 240;
	{8'd165,8'd76} : s = 241;
	{8'd165,8'd77} : s = 242;
	{8'd165,8'd78} : s = 243;
	{8'd165,8'd79} : s = 244;
	{8'd165,8'd80} : s = 245;
	{8'd165,8'd81} : s = 246;
	{8'd165,8'd82} : s = 247;
	{8'd165,8'd83} : s = 248;
	{8'd165,8'd84} : s = 249;
	{8'd165,8'd85} : s = 250;
	{8'd165,8'd86} : s = 251;
	{8'd165,8'd87} : s = 252;
	{8'd165,8'd88} : s = 253;
	{8'd165,8'd89} : s = 254;
	{8'd165,8'd90} : s = 255;
	{8'd165,8'd91} : s = 256;
	{8'd165,8'd92} : s = 257;
	{8'd165,8'd93} : s = 258;
	{8'd165,8'd94} : s = 259;
	{8'd165,8'd95} : s = 260;
	{8'd165,8'd96} : s = 261;
	{8'd165,8'd97} : s = 262;
	{8'd165,8'd98} : s = 263;
	{8'd165,8'd99} : s = 264;
	{8'd165,8'd100} : s = 265;
	{8'd165,8'd101} : s = 266;
	{8'd165,8'd102} : s = 267;
	{8'd165,8'd103} : s = 268;
	{8'd165,8'd104} : s = 269;
	{8'd165,8'd105} : s = 270;
	{8'd165,8'd106} : s = 271;
	{8'd165,8'd107} : s = 272;
	{8'd165,8'd108} : s = 273;
	{8'd165,8'd109} : s = 274;
	{8'd165,8'd110} : s = 275;
	{8'd165,8'd111} : s = 276;
	{8'd165,8'd112} : s = 277;
	{8'd165,8'd113} : s = 278;
	{8'd165,8'd114} : s = 279;
	{8'd165,8'd115} : s = 280;
	{8'd165,8'd116} : s = 281;
	{8'd165,8'd117} : s = 282;
	{8'd165,8'd118} : s = 283;
	{8'd165,8'd119} : s = 284;
	{8'd165,8'd120} : s = 285;
	{8'd165,8'd121} : s = 286;
	{8'd165,8'd122} : s = 287;
	{8'd165,8'd123} : s = 288;
	{8'd165,8'd124} : s = 289;
	{8'd165,8'd125} : s = 290;
	{8'd165,8'd126} : s = 291;
	{8'd165,8'd127} : s = 292;
	{8'd165,8'd128} : s = 293;
	{8'd165,8'd129} : s = 294;
	{8'd165,8'd130} : s = 295;
	{8'd165,8'd131} : s = 296;
	{8'd165,8'd132} : s = 297;
	{8'd165,8'd133} : s = 298;
	{8'd165,8'd134} : s = 299;
	{8'd165,8'd135} : s = 300;
	{8'd165,8'd136} : s = 301;
	{8'd165,8'd137} : s = 302;
	{8'd165,8'd138} : s = 303;
	{8'd165,8'd139} : s = 304;
	{8'd165,8'd140} : s = 305;
	{8'd165,8'd141} : s = 306;
	{8'd165,8'd142} : s = 307;
	{8'd165,8'd143} : s = 308;
	{8'd165,8'd144} : s = 309;
	{8'd165,8'd145} : s = 310;
	{8'd165,8'd146} : s = 311;
	{8'd165,8'd147} : s = 312;
	{8'd165,8'd148} : s = 313;
	{8'd165,8'd149} : s = 314;
	{8'd165,8'd150} : s = 315;
	{8'd165,8'd151} : s = 316;
	{8'd165,8'd152} : s = 317;
	{8'd165,8'd153} : s = 318;
	{8'd165,8'd154} : s = 319;
	{8'd165,8'd155} : s = 320;
	{8'd165,8'd156} : s = 321;
	{8'd165,8'd157} : s = 322;
	{8'd165,8'd158} : s = 323;
	{8'd165,8'd159} : s = 324;
	{8'd165,8'd160} : s = 325;
	{8'd165,8'd161} : s = 326;
	{8'd165,8'd162} : s = 327;
	{8'd165,8'd163} : s = 328;
	{8'd165,8'd164} : s = 329;
	{8'd165,8'd165} : s = 330;
	{8'd165,8'd166} : s = 331;
	{8'd165,8'd167} : s = 332;
	{8'd165,8'd168} : s = 333;
	{8'd165,8'd169} : s = 334;
	{8'd165,8'd170} : s = 335;
	{8'd165,8'd171} : s = 336;
	{8'd165,8'd172} : s = 337;
	{8'd165,8'd173} : s = 338;
	{8'd165,8'd174} : s = 339;
	{8'd165,8'd175} : s = 340;
	{8'd165,8'd176} : s = 341;
	{8'd165,8'd177} : s = 342;
	{8'd165,8'd178} : s = 343;
	{8'd165,8'd179} : s = 344;
	{8'd165,8'd180} : s = 345;
	{8'd165,8'd181} : s = 346;
	{8'd165,8'd182} : s = 347;
	{8'd165,8'd183} : s = 348;
	{8'd165,8'd184} : s = 349;
	{8'd165,8'd185} : s = 350;
	{8'd165,8'd186} : s = 351;
	{8'd165,8'd187} : s = 352;
	{8'd165,8'd188} : s = 353;
	{8'd165,8'd189} : s = 354;
	{8'd165,8'd190} : s = 355;
	{8'd165,8'd191} : s = 356;
	{8'd165,8'd192} : s = 357;
	{8'd165,8'd193} : s = 358;
	{8'd165,8'd194} : s = 359;
	{8'd165,8'd195} : s = 360;
	{8'd165,8'd196} : s = 361;
	{8'd165,8'd197} : s = 362;
	{8'd165,8'd198} : s = 363;
	{8'd165,8'd199} : s = 364;
	{8'd165,8'd200} : s = 365;
	{8'd165,8'd201} : s = 366;
	{8'd165,8'd202} : s = 367;
	{8'd165,8'd203} : s = 368;
	{8'd165,8'd204} : s = 369;
	{8'd165,8'd205} : s = 370;
	{8'd165,8'd206} : s = 371;
	{8'd165,8'd207} : s = 372;
	{8'd165,8'd208} : s = 373;
	{8'd165,8'd209} : s = 374;
	{8'd165,8'd210} : s = 375;
	{8'd165,8'd211} : s = 376;
	{8'd165,8'd212} : s = 377;
	{8'd165,8'd213} : s = 378;
	{8'd165,8'd214} : s = 379;
	{8'd165,8'd215} : s = 380;
	{8'd165,8'd216} : s = 381;
	{8'd165,8'd217} : s = 382;
	{8'd165,8'd218} : s = 383;
	{8'd165,8'd219} : s = 384;
	{8'd165,8'd220} : s = 385;
	{8'd165,8'd221} : s = 386;
	{8'd165,8'd222} : s = 387;
	{8'd165,8'd223} : s = 388;
	{8'd165,8'd224} : s = 389;
	{8'd165,8'd225} : s = 390;
	{8'd165,8'd226} : s = 391;
	{8'd165,8'd227} : s = 392;
	{8'd165,8'd228} : s = 393;
	{8'd165,8'd229} : s = 394;
	{8'd165,8'd230} : s = 395;
	{8'd165,8'd231} : s = 396;
	{8'd165,8'd232} : s = 397;
	{8'd165,8'd233} : s = 398;
	{8'd165,8'd234} : s = 399;
	{8'd165,8'd235} : s = 400;
	{8'd165,8'd236} : s = 401;
	{8'd165,8'd237} : s = 402;
	{8'd165,8'd238} : s = 403;
	{8'd165,8'd239} : s = 404;
	{8'd165,8'd240} : s = 405;
	{8'd165,8'd241} : s = 406;
	{8'd165,8'd242} : s = 407;
	{8'd165,8'd243} : s = 408;
	{8'd165,8'd244} : s = 409;
	{8'd165,8'd245} : s = 410;
	{8'd165,8'd246} : s = 411;
	{8'd165,8'd247} : s = 412;
	{8'd165,8'd248} : s = 413;
	{8'd165,8'd249} : s = 414;
	{8'd165,8'd250} : s = 415;
	{8'd165,8'd251} : s = 416;
	{8'd165,8'd252} : s = 417;
	{8'd165,8'd253} : s = 418;
	{8'd165,8'd254} : s = 419;
	{8'd165,8'd255} : s = 420;
	{8'd166,8'd0} : s = 166;
	{8'd166,8'd1} : s = 167;
	{8'd166,8'd2} : s = 168;
	{8'd166,8'd3} : s = 169;
	{8'd166,8'd4} : s = 170;
	{8'd166,8'd5} : s = 171;
	{8'd166,8'd6} : s = 172;
	{8'd166,8'd7} : s = 173;
	{8'd166,8'd8} : s = 174;
	{8'd166,8'd9} : s = 175;
	{8'd166,8'd10} : s = 176;
	{8'd166,8'd11} : s = 177;
	{8'd166,8'd12} : s = 178;
	{8'd166,8'd13} : s = 179;
	{8'd166,8'd14} : s = 180;
	{8'd166,8'd15} : s = 181;
	{8'd166,8'd16} : s = 182;
	{8'd166,8'd17} : s = 183;
	{8'd166,8'd18} : s = 184;
	{8'd166,8'd19} : s = 185;
	{8'd166,8'd20} : s = 186;
	{8'd166,8'd21} : s = 187;
	{8'd166,8'd22} : s = 188;
	{8'd166,8'd23} : s = 189;
	{8'd166,8'd24} : s = 190;
	{8'd166,8'd25} : s = 191;
	{8'd166,8'd26} : s = 192;
	{8'd166,8'd27} : s = 193;
	{8'd166,8'd28} : s = 194;
	{8'd166,8'd29} : s = 195;
	{8'd166,8'd30} : s = 196;
	{8'd166,8'd31} : s = 197;
	{8'd166,8'd32} : s = 198;
	{8'd166,8'd33} : s = 199;
	{8'd166,8'd34} : s = 200;
	{8'd166,8'd35} : s = 201;
	{8'd166,8'd36} : s = 202;
	{8'd166,8'd37} : s = 203;
	{8'd166,8'd38} : s = 204;
	{8'd166,8'd39} : s = 205;
	{8'd166,8'd40} : s = 206;
	{8'd166,8'd41} : s = 207;
	{8'd166,8'd42} : s = 208;
	{8'd166,8'd43} : s = 209;
	{8'd166,8'd44} : s = 210;
	{8'd166,8'd45} : s = 211;
	{8'd166,8'd46} : s = 212;
	{8'd166,8'd47} : s = 213;
	{8'd166,8'd48} : s = 214;
	{8'd166,8'd49} : s = 215;
	{8'd166,8'd50} : s = 216;
	{8'd166,8'd51} : s = 217;
	{8'd166,8'd52} : s = 218;
	{8'd166,8'd53} : s = 219;
	{8'd166,8'd54} : s = 220;
	{8'd166,8'd55} : s = 221;
	{8'd166,8'd56} : s = 222;
	{8'd166,8'd57} : s = 223;
	{8'd166,8'd58} : s = 224;
	{8'd166,8'd59} : s = 225;
	{8'd166,8'd60} : s = 226;
	{8'd166,8'd61} : s = 227;
	{8'd166,8'd62} : s = 228;
	{8'd166,8'd63} : s = 229;
	{8'd166,8'd64} : s = 230;
	{8'd166,8'd65} : s = 231;
	{8'd166,8'd66} : s = 232;
	{8'd166,8'd67} : s = 233;
	{8'd166,8'd68} : s = 234;
	{8'd166,8'd69} : s = 235;
	{8'd166,8'd70} : s = 236;
	{8'd166,8'd71} : s = 237;
	{8'd166,8'd72} : s = 238;
	{8'd166,8'd73} : s = 239;
	{8'd166,8'd74} : s = 240;
	{8'd166,8'd75} : s = 241;
	{8'd166,8'd76} : s = 242;
	{8'd166,8'd77} : s = 243;
	{8'd166,8'd78} : s = 244;
	{8'd166,8'd79} : s = 245;
	{8'd166,8'd80} : s = 246;
	{8'd166,8'd81} : s = 247;
	{8'd166,8'd82} : s = 248;
	{8'd166,8'd83} : s = 249;
	{8'd166,8'd84} : s = 250;
	{8'd166,8'd85} : s = 251;
	{8'd166,8'd86} : s = 252;
	{8'd166,8'd87} : s = 253;
	{8'd166,8'd88} : s = 254;
	{8'd166,8'd89} : s = 255;
	{8'd166,8'd90} : s = 256;
	{8'd166,8'd91} : s = 257;
	{8'd166,8'd92} : s = 258;
	{8'd166,8'd93} : s = 259;
	{8'd166,8'd94} : s = 260;
	{8'd166,8'd95} : s = 261;
	{8'd166,8'd96} : s = 262;
	{8'd166,8'd97} : s = 263;
	{8'd166,8'd98} : s = 264;
	{8'd166,8'd99} : s = 265;
	{8'd166,8'd100} : s = 266;
	{8'd166,8'd101} : s = 267;
	{8'd166,8'd102} : s = 268;
	{8'd166,8'd103} : s = 269;
	{8'd166,8'd104} : s = 270;
	{8'd166,8'd105} : s = 271;
	{8'd166,8'd106} : s = 272;
	{8'd166,8'd107} : s = 273;
	{8'd166,8'd108} : s = 274;
	{8'd166,8'd109} : s = 275;
	{8'd166,8'd110} : s = 276;
	{8'd166,8'd111} : s = 277;
	{8'd166,8'd112} : s = 278;
	{8'd166,8'd113} : s = 279;
	{8'd166,8'd114} : s = 280;
	{8'd166,8'd115} : s = 281;
	{8'd166,8'd116} : s = 282;
	{8'd166,8'd117} : s = 283;
	{8'd166,8'd118} : s = 284;
	{8'd166,8'd119} : s = 285;
	{8'd166,8'd120} : s = 286;
	{8'd166,8'd121} : s = 287;
	{8'd166,8'd122} : s = 288;
	{8'd166,8'd123} : s = 289;
	{8'd166,8'd124} : s = 290;
	{8'd166,8'd125} : s = 291;
	{8'd166,8'd126} : s = 292;
	{8'd166,8'd127} : s = 293;
	{8'd166,8'd128} : s = 294;
	{8'd166,8'd129} : s = 295;
	{8'd166,8'd130} : s = 296;
	{8'd166,8'd131} : s = 297;
	{8'd166,8'd132} : s = 298;
	{8'd166,8'd133} : s = 299;
	{8'd166,8'd134} : s = 300;
	{8'd166,8'd135} : s = 301;
	{8'd166,8'd136} : s = 302;
	{8'd166,8'd137} : s = 303;
	{8'd166,8'd138} : s = 304;
	{8'd166,8'd139} : s = 305;
	{8'd166,8'd140} : s = 306;
	{8'd166,8'd141} : s = 307;
	{8'd166,8'd142} : s = 308;
	{8'd166,8'd143} : s = 309;
	{8'd166,8'd144} : s = 310;
	{8'd166,8'd145} : s = 311;
	{8'd166,8'd146} : s = 312;
	{8'd166,8'd147} : s = 313;
	{8'd166,8'd148} : s = 314;
	{8'd166,8'd149} : s = 315;
	{8'd166,8'd150} : s = 316;
	{8'd166,8'd151} : s = 317;
	{8'd166,8'd152} : s = 318;
	{8'd166,8'd153} : s = 319;
	{8'd166,8'd154} : s = 320;
	{8'd166,8'd155} : s = 321;
	{8'd166,8'd156} : s = 322;
	{8'd166,8'd157} : s = 323;
	{8'd166,8'd158} : s = 324;
	{8'd166,8'd159} : s = 325;
	{8'd166,8'd160} : s = 326;
	{8'd166,8'd161} : s = 327;
	{8'd166,8'd162} : s = 328;
	{8'd166,8'd163} : s = 329;
	{8'd166,8'd164} : s = 330;
	{8'd166,8'd165} : s = 331;
	{8'd166,8'd166} : s = 332;
	{8'd166,8'd167} : s = 333;
	{8'd166,8'd168} : s = 334;
	{8'd166,8'd169} : s = 335;
	{8'd166,8'd170} : s = 336;
	{8'd166,8'd171} : s = 337;
	{8'd166,8'd172} : s = 338;
	{8'd166,8'd173} : s = 339;
	{8'd166,8'd174} : s = 340;
	{8'd166,8'd175} : s = 341;
	{8'd166,8'd176} : s = 342;
	{8'd166,8'd177} : s = 343;
	{8'd166,8'd178} : s = 344;
	{8'd166,8'd179} : s = 345;
	{8'd166,8'd180} : s = 346;
	{8'd166,8'd181} : s = 347;
	{8'd166,8'd182} : s = 348;
	{8'd166,8'd183} : s = 349;
	{8'd166,8'd184} : s = 350;
	{8'd166,8'd185} : s = 351;
	{8'd166,8'd186} : s = 352;
	{8'd166,8'd187} : s = 353;
	{8'd166,8'd188} : s = 354;
	{8'd166,8'd189} : s = 355;
	{8'd166,8'd190} : s = 356;
	{8'd166,8'd191} : s = 357;
	{8'd166,8'd192} : s = 358;
	{8'd166,8'd193} : s = 359;
	{8'd166,8'd194} : s = 360;
	{8'd166,8'd195} : s = 361;
	{8'd166,8'd196} : s = 362;
	{8'd166,8'd197} : s = 363;
	{8'd166,8'd198} : s = 364;
	{8'd166,8'd199} : s = 365;
	{8'd166,8'd200} : s = 366;
	{8'd166,8'd201} : s = 367;
	{8'd166,8'd202} : s = 368;
	{8'd166,8'd203} : s = 369;
	{8'd166,8'd204} : s = 370;
	{8'd166,8'd205} : s = 371;
	{8'd166,8'd206} : s = 372;
	{8'd166,8'd207} : s = 373;
	{8'd166,8'd208} : s = 374;
	{8'd166,8'd209} : s = 375;
	{8'd166,8'd210} : s = 376;
	{8'd166,8'd211} : s = 377;
	{8'd166,8'd212} : s = 378;
	{8'd166,8'd213} : s = 379;
	{8'd166,8'd214} : s = 380;
	{8'd166,8'd215} : s = 381;
	{8'd166,8'd216} : s = 382;
	{8'd166,8'd217} : s = 383;
	{8'd166,8'd218} : s = 384;
	{8'd166,8'd219} : s = 385;
	{8'd166,8'd220} : s = 386;
	{8'd166,8'd221} : s = 387;
	{8'd166,8'd222} : s = 388;
	{8'd166,8'd223} : s = 389;
	{8'd166,8'd224} : s = 390;
	{8'd166,8'd225} : s = 391;
	{8'd166,8'd226} : s = 392;
	{8'd166,8'd227} : s = 393;
	{8'd166,8'd228} : s = 394;
	{8'd166,8'd229} : s = 395;
	{8'd166,8'd230} : s = 396;
	{8'd166,8'd231} : s = 397;
	{8'd166,8'd232} : s = 398;
	{8'd166,8'd233} : s = 399;
	{8'd166,8'd234} : s = 400;
	{8'd166,8'd235} : s = 401;
	{8'd166,8'd236} : s = 402;
	{8'd166,8'd237} : s = 403;
	{8'd166,8'd238} : s = 404;
	{8'd166,8'd239} : s = 405;
	{8'd166,8'd240} : s = 406;
	{8'd166,8'd241} : s = 407;
	{8'd166,8'd242} : s = 408;
	{8'd166,8'd243} : s = 409;
	{8'd166,8'd244} : s = 410;
	{8'd166,8'd245} : s = 411;
	{8'd166,8'd246} : s = 412;
	{8'd166,8'd247} : s = 413;
	{8'd166,8'd248} : s = 414;
	{8'd166,8'd249} : s = 415;
	{8'd166,8'd250} : s = 416;
	{8'd166,8'd251} : s = 417;
	{8'd166,8'd252} : s = 418;
	{8'd166,8'd253} : s = 419;
	{8'd166,8'd254} : s = 420;
	{8'd166,8'd255} : s = 421;
	{8'd167,8'd0} : s = 167;
	{8'd167,8'd1} : s = 168;
	{8'd167,8'd2} : s = 169;
	{8'd167,8'd3} : s = 170;
	{8'd167,8'd4} : s = 171;
	{8'd167,8'd5} : s = 172;
	{8'd167,8'd6} : s = 173;
	{8'd167,8'd7} : s = 174;
	{8'd167,8'd8} : s = 175;
	{8'd167,8'd9} : s = 176;
	{8'd167,8'd10} : s = 177;
	{8'd167,8'd11} : s = 178;
	{8'd167,8'd12} : s = 179;
	{8'd167,8'd13} : s = 180;
	{8'd167,8'd14} : s = 181;
	{8'd167,8'd15} : s = 182;
	{8'd167,8'd16} : s = 183;
	{8'd167,8'd17} : s = 184;
	{8'd167,8'd18} : s = 185;
	{8'd167,8'd19} : s = 186;
	{8'd167,8'd20} : s = 187;
	{8'd167,8'd21} : s = 188;
	{8'd167,8'd22} : s = 189;
	{8'd167,8'd23} : s = 190;
	{8'd167,8'd24} : s = 191;
	{8'd167,8'd25} : s = 192;
	{8'd167,8'd26} : s = 193;
	{8'd167,8'd27} : s = 194;
	{8'd167,8'd28} : s = 195;
	{8'd167,8'd29} : s = 196;
	{8'd167,8'd30} : s = 197;
	{8'd167,8'd31} : s = 198;
	{8'd167,8'd32} : s = 199;
	{8'd167,8'd33} : s = 200;
	{8'd167,8'd34} : s = 201;
	{8'd167,8'd35} : s = 202;
	{8'd167,8'd36} : s = 203;
	{8'd167,8'd37} : s = 204;
	{8'd167,8'd38} : s = 205;
	{8'd167,8'd39} : s = 206;
	{8'd167,8'd40} : s = 207;
	{8'd167,8'd41} : s = 208;
	{8'd167,8'd42} : s = 209;
	{8'd167,8'd43} : s = 210;
	{8'd167,8'd44} : s = 211;
	{8'd167,8'd45} : s = 212;
	{8'd167,8'd46} : s = 213;
	{8'd167,8'd47} : s = 214;
	{8'd167,8'd48} : s = 215;
	{8'd167,8'd49} : s = 216;
	{8'd167,8'd50} : s = 217;
	{8'd167,8'd51} : s = 218;
	{8'd167,8'd52} : s = 219;
	{8'd167,8'd53} : s = 220;
	{8'd167,8'd54} : s = 221;
	{8'd167,8'd55} : s = 222;
	{8'd167,8'd56} : s = 223;
	{8'd167,8'd57} : s = 224;
	{8'd167,8'd58} : s = 225;
	{8'd167,8'd59} : s = 226;
	{8'd167,8'd60} : s = 227;
	{8'd167,8'd61} : s = 228;
	{8'd167,8'd62} : s = 229;
	{8'd167,8'd63} : s = 230;
	{8'd167,8'd64} : s = 231;
	{8'd167,8'd65} : s = 232;
	{8'd167,8'd66} : s = 233;
	{8'd167,8'd67} : s = 234;
	{8'd167,8'd68} : s = 235;
	{8'd167,8'd69} : s = 236;
	{8'd167,8'd70} : s = 237;
	{8'd167,8'd71} : s = 238;
	{8'd167,8'd72} : s = 239;
	{8'd167,8'd73} : s = 240;
	{8'd167,8'd74} : s = 241;
	{8'd167,8'd75} : s = 242;
	{8'd167,8'd76} : s = 243;
	{8'd167,8'd77} : s = 244;
	{8'd167,8'd78} : s = 245;
	{8'd167,8'd79} : s = 246;
	{8'd167,8'd80} : s = 247;
	{8'd167,8'd81} : s = 248;
	{8'd167,8'd82} : s = 249;
	{8'd167,8'd83} : s = 250;
	{8'd167,8'd84} : s = 251;
	{8'd167,8'd85} : s = 252;
	{8'd167,8'd86} : s = 253;
	{8'd167,8'd87} : s = 254;
	{8'd167,8'd88} : s = 255;
	{8'd167,8'd89} : s = 256;
	{8'd167,8'd90} : s = 257;
	{8'd167,8'd91} : s = 258;
	{8'd167,8'd92} : s = 259;
	{8'd167,8'd93} : s = 260;
	{8'd167,8'd94} : s = 261;
	{8'd167,8'd95} : s = 262;
	{8'd167,8'd96} : s = 263;
	{8'd167,8'd97} : s = 264;
	{8'd167,8'd98} : s = 265;
	{8'd167,8'd99} : s = 266;
	{8'd167,8'd100} : s = 267;
	{8'd167,8'd101} : s = 268;
	{8'd167,8'd102} : s = 269;
	{8'd167,8'd103} : s = 270;
	{8'd167,8'd104} : s = 271;
	{8'd167,8'd105} : s = 272;
	{8'd167,8'd106} : s = 273;
	{8'd167,8'd107} : s = 274;
	{8'd167,8'd108} : s = 275;
	{8'd167,8'd109} : s = 276;
	{8'd167,8'd110} : s = 277;
	{8'd167,8'd111} : s = 278;
	{8'd167,8'd112} : s = 279;
	{8'd167,8'd113} : s = 280;
	{8'd167,8'd114} : s = 281;
	{8'd167,8'd115} : s = 282;
	{8'd167,8'd116} : s = 283;
	{8'd167,8'd117} : s = 284;
	{8'd167,8'd118} : s = 285;
	{8'd167,8'd119} : s = 286;
	{8'd167,8'd120} : s = 287;
	{8'd167,8'd121} : s = 288;
	{8'd167,8'd122} : s = 289;
	{8'd167,8'd123} : s = 290;
	{8'd167,8'd124} : s = 291;
	{8'd167,8'd125} : s = 292;
	{8'd167,8'd126} : s = 293;
	{8'd167,8'd127} : s = 294;
	{8'd167,8'd128} : s = 295;
	{8'd167,8'd129} : s = 296;
	{8'd167,8'd130} : s = 297;
	{8'd167,8'd131} : s = 298;
	{8'd167,8'd132} : s = 299;
	{8'd167,8'd133} : s = 300;
	{8'd167,8'd134} : s = 301;
	{8'd167,8'd135} : s = 302;
	{8'd167,8'd136} : s = 303;
	{8'd167,8'd137} : s = 304;
	{8'd167,8'd138} : s = 305;
	{8'd167,8'd139} : s = 306;
	{8'd167,8'd140} : s = 307;
	{8'd167,8'd141} : s = 308;
	{8'd167,8'd142} : s = 309;
	{8'd167,8'd143} : s = 310;
	{8'd167,8'd144} : s = 311;
	{8'd167,8'd145} : s = 312;
	{8'd167,8'd146} : s = 313;
	{8'd167,8'd147} : s = 314;
	{8'd167,8'd148} : s = 315;
	{8'd167,8'd149} : s = 316;
	{8'd167,8'd150} : s = 317;
	{8'd167,8'd151} : s = 318;
	{8'd167,8'd152} : s = 319;
	{8'd167,8'd153} : s = 320;
	{8'd167,8'd154} : s = 321;
	{8'd167,8'd155} : s = 322;
	{8'd167,8'd156} : s = 323;
	{8'd167,8'd157} : s = 324;
	{8'd167,8'd158} : s = 325;
	{8'd167,8'd159} : s = 326;
	{8'd167,8'd160} : s = 327;
	{8'd167,8'd161} : s = 328;
	{8'd167,8'd162} : s = 329;
	{8'd167,8'd163} : s = 330;
	{8'd167,8'd164} : s = 331;
	{8'd167,8'd165} : s = 332;
	{8'd167,8'd166} : s = 333;
	{8'd167,8'd167} : s = 334;
	{8'd167,8'd168} : s = 335;
	{8'd167,8'd169} : s = 336;
	{8'd167,8'd170} : s = 337;
	{8'd167,8'd171} : s = 338;
	{8'd167,8'd172} : s = 339;
	{8'd167,8'd173} : s = 340;
	{8'd167,8'd174} : s = 341;
	{8'd167,8'd175} : s = 342;
	{8'd167,8'd176} : s = 343;
	{8'd167,8'd177} : s = 344;
	{8'd167,8'd178} : s = 345;
	{8'd167,8'd179} : s = 346;
	{8'd167,8'd180} : s = 347;
	{8'd167,8'd181} : s = 348;
	{8'd167,8'd182} : s = 349;
	{8'd167,8'd183} : s = 350;
	{8'd167,8'd184} : s = 351;
	{8'd167,8'd185} : s = 352;
	{8'd167,8'd186} : s = 353;
	{8'd167,8'd187} : s = 354;
	{8'd167,8'd188} : s = 355;
	{8'd167,8'd189} : s = 356;
	{8'd167,8'd190} : s = 357;
	{8'd167,8'd191} : s = 358;
	{8'd167,8'd192} : s = 359;
	{8'd167,8'd193} : s = 360;
	{8'd167,8'd194} : s = 361;
	{8'd167,8'd195} : s = 362;
	{8'd167,8'd196} : s = 363;
	{8'd167,8'd197} : s = 364;
	{8'd167,8'd198} : s = 365;
	{8'd167,8'd199} : s = 366;
	{8'd167,8'd200} : s = 367;
	{8'd167,8'd201} : s = 368;
	{8'd167,8'd202} : s = 369;
	{8'd167,8'd203} : s = 370;
	{8'd167,8'd204} : s = 371;
	{8'd167,8'd205} : s = 372;
	{8'd167,8'd206} : s = 373;
	{8'd167,8'd207} : s = 374;
	{8'd167,8'd208} : s = 375;
	{8'd167,8'd209} : s = 376;
	{8'd167,8'd210} : s = 377;
	{8'd167,8'd211} : s = 378;
	{8'd167,8'd212} : s = 379;
	{8'd167,8'd213} : s = 380;
	{8'd167,8'd214} : s = 381;
	{8'd167,8'd215} : s = 382;
	{8'd167,8'd216} : s = 383;
	{8'd167,8'd217} : s = 384;
	{8'd167,8'd218} : s = 385;
	{8'd167,8'd219} : s = 386;
	{8'd167,8'd220} : s = 387;
	{8'd167,8'd221} : s = 388;
	{8'd167,8'd222} : s = 389;
	{8'd167,8'd223} : s = 390;
	{8'd167,8'd224} : s = 391;
	{8'd167,8'd225} : s = 392;
	{8'd167,8'd226} : s = 393;
	{8'd167,8'd227} : s = 394;
	{8'd167,8'd228} : s = 395;
	{8'd167,8'd229} : s = 396;
	{8'd167,8'd230} : s = 397;
	{8'd167,8'd231} : s = 398;
	{8'd167,8'd232} : s = 399;
	{8'd167,8'd233} : s = 400;
	{8'd167,8'd234} : s = 401;
	{8'd167,8'd235} : s = 402;
	{8'd167,8'd236} : s = 403;
	{8'd167,8'd237} : s = 404;
	{8'd167,8'd238} : s = 405;
	{8'd167,8'd239} : s = 406;
	{8'd167,8'd240} : s = 407;
	{8'd167,8'd241} : s = 408;
	{8'd167,8'd242} : s = 409;
	{8'd167,8'd243} : s = 410;
	{8'd167,8'd244} : s = 411;
	{8'd167,8'd245} : s = 412;
	{8'd167,8'd246} : s = 413;
	{8'd167,8'd247} : s = 414;
	{8'd167,8'd248} : s = 415;
	{8'd167,8'd249} : s = 416;
	{8'd167,8'd250} : s = 417;
	{8'd167,8'd251} : s = 418;
	{8'd167,8'd252} : s = 419;
	{8'd167,8'd253} : s = 420;
	{8'd167,8'd254} : s = 421;
	{8'd167,8'd255} : s = 422;
	{8'd168,8'd0} : s = 168;
	{8'd168,8'd1} : s = 169;
	{8'd168,8'd2} : s = 170;
	{8'd168,8'd3} : s = 171;
	{8'd168,8'd4} : s = 172;
	{8'd168,8'd5} : s = 173;
	{8'd168,8'd6} : s = 174;
	{8'd168,8'd7} : s = 175;
	{8'd168,8'd8} : s = 176;
	{8'd168,8'd9} : s = 177;
	{8'd168,8'd10} : s = 178;
	{8'd168,8'd11} : s = 179;
	{8'd168,8'd12} : s = 180;
	{8'd168,8'd13} : s = 181;
	{8'd168,8'd14} : s = 182;
	{8'd168,8'd15} : s = 183;
	{8'd168,8'd16} : s = 184;
	{8'd168,8'd17} : s = 185;
	{8'd168,8'd18} : s = 186;
	{8'd168,8'd19} : s = 187;
	{8'd168,8'd20} : s = 188;
	{8'd168,8'd21} : s = 189;
	{8'd168,8'd22} : s = 190;
	{8'd168,8'd23} : s = 191;
	{8'd168,8'd24} : s = 192;
	{8'd168,8'd25} : s = 193;
	{8'd168,8'd26} : s = 194;
	{8'd168,8'd27} : s = 195;
	{8'd168,8'd28} : s = 196;
	{8'd168,8'd29} : s = 197;
	{8'd168,8'd30} : s = 198;
	{8'd168,8'd31} : s = 199;
	{8'd168,8'd32} : s = 200;
	{8'd168,8'd33} : s = 201;
	{8'd168,8'd34} : s = 202;
	{8'd168,8'd35} : s = 203;
	{8'd168,8'd36} : s = 204;
	{8'd168,8'd37} : s = 205;
	{8'd168,8'd38} : s = 206;
	{8'd168,8'd39} : s = 207;
	{8'd168,8'd40} : s = 208;
	{8'd168,8'd41} : s = 209;
	{8'd168,8'd42} : s = 210;
	{8'd168,8'd43} : s = 211;
	{8'd168,8'd44} : s = 212;
	{8'd168,8'd45} : s = 213;
	{8'd168,8'd46} : s = 214;
	{8'd168,8'd47} : s = 215;
	{8'd168,8'd48} : s = 216;
	{8'd168,8'd49} : s = 217;
	{8'd168,8'd50} : s = 218;
	{8'd168,8'd51} : s = 219;
	{8'd168,8'd52} : s = 220;
	{8'd168,8'd53} : s = 221;
	{8'd168,8'd54} : s = 222;
	{8'd168,8'd55} : s = 223;
	{8'd168,8'd56} : s = 224;
	{8'd168,8'd57} : s = 225;
	{8'd168,8'd58} : s = 226;
	{8'd168,8'd59} : s = 227;
	{8'd168,8'd60} : s = 228;
	{8'd168,8'd61} : s = 229;
	{8'd168,8'd62} : s = 230;
	{8'd168,8'd63} : s = 231;
	{8'd168,8'd64} : s = 232;
	{8'd168,8'd65} : s = 233;
	{8'd168,8'd66} : s = 234;
	{8'd168,8'd67} : s = 235;
	{8'd168,8'd68} : s = 236;
	{8'd168,8'd69} : s = 237;
	{8'd168,8'd70} : s = 238;
	{8'd168,8'd71} : s = 239;
	{8'd168,8'd72} : s = 240;
	{8'd168,8'd73} : s = 241;
	{8'd168,8'd74} : s = 242;
	{8'd168,8'd75} : s = 243;
	{8'd168,8'd76} : s = 244;
	{8'd168,8'd77} : s = 245;
	{8'd168,8'd78} : s = 246;
	{8'd168,8'd79} : s = 247;
	{8'd168,8'd80} : s = 248;
	{8'd168,8'd81} : s = 249;
	{8'd168,8'd82} : s = 250;
	{8'd168,8'd83} : s = 251;
	{8'd168,8'd84} : s = 252;
	{8'd168,8'd85} : s = 253;
	{8'd168,8'd86} : s = 254;
	{8'd168,8'd87} : s = 255;
	{8'd168,8'd88} : s = 256;
	{8'd168,8'd89} : s = 257;
	{8'd168,8'd90} : s = 258;
	{8'd168,8'd91} : s = 259;
	{8'd168,8'd92} : s = 260;
	{8'd168,8'd93} : s = 261;
	{8'd168,8'd94} : s = 262;
	{8'd168,8'd95} : s = 263;
	{8'd168,8'd96} : s = 264;
	{8'd168,8'd97} : s = 265;
	{8'd168,8'd98} : s = 266;
	{8'd168,8'd99} : s = 267;
	{8'd168,8'd100} : s = 268;
	{8'd168,8'd101} : s = 269;
	{8'd168,8'd102} : s = 270;
	{8'd168,8'd103} : s = 271;
	{8'd168,8'd104} : s = 272;
	{8'd168,8'd105} : s = 273;
	{8'd168,8'd106} : s = 274;
	{8'd168,8'd107} : s = 275;
	{8'd168,8'd108} : s = 276;
	{8'd168,8'd109} : s = 277;
	{8'd168,8'd110} : s = 278;
	{8'd168,8'd111} : s = 279;
	{8'd168,8'd112} : s = 280;
	{8'd168,8'd113} : s = 281;
	{8'd168,8'd114} : s = 282;
	{8'd168,8'd115} : s = 283;
	{8'd168,8'd116} : s = 284;
	{8'd168,8'd117} : s = 285;
	{8'd168,8'd118} : s = 286;
	{8'd168,8'd119} : s = 287;
	{8'd168,8'd120} : s = 288;
	{8'd168,8'd121} : s = 289;
	{8'd168,8'd122} : s = 290;
	{8'd168,8'd123} : s = 291;
	{8'd168,8'd124} : s = 292;
	{8'd168,8'd125} : s = 293;
	{8'd168,8'd126} : s = 294;
	{8'd168,8'd127} : s = 295;
	{8'd168,8'd128} : s = 296;
	{8'd168,8'd129} : s = 297;
	{8'd168,8'd130} : s = 298;
	{8'd168,8'd131} : s = 299;
	{8'd168,8'd132} : s = 300;
	{8'd168,8'd133} : s = 301;
	{8'd168,8'd134} : s = 302;
	{8'd168,8'd135} : s = 303;
	{8'd168,8'd136} : s = 304;
	{8'd168,8'd137} : s = 305;
	{8'd168,8'd138} : s = 306;
	{8'd168,8'd139} : s = 307;
	{8'd168,8'd140} : s = 308;
	{8'd168,8'd141} : s = 309;
	{8'd168,8'd142} : s = 310;
	{8'd168,8'd143} : s = 311;
	{8'd168,8'd144} : s = 312;
	{8'd168,8'd145} : s = 313;
	{8'd168,8'd146} : s = 314;
	{8'd168,8'd147} : s = 315;
	{8'd168,8'd148} : s = 316;
	{8'd168,8'd149} : s = 317;
	{8'd168,8'd150} : s = 318;
	{8'd168,8'd151} : s = 319;
	{8'd168,8'd152} : s = 320;
	{8'd168,8'd153} : s = 321;
	{8'd168,8'd154} : s = 322;
	{8'd168,8'd155} : s = 323;
	{8'd168,8'd156} : s = 324;
	{8'd168,8'd157} : s = 325;
	{8'd168,8'd158} : s = 326;
	{8'd168,8'd159} : s = 327;
	{8'd168,8'd160} : s = 328;
	{8'd168,8'd161} : s = 329;
	{8'd168,8'd162} : s = 330;
	{8'd168,8'd163} : s = 331;
	{8'd168,8'd164} : s = 332;
	{8'd168,8'd165} : s = 333;
	{8'd168,8'd166} : s = 334;
	{8'd168,8'd167} : s = 335;
	{8'd168,8'd168} : s = 336;
	{8'd168,8'd169} : s = 337;
	{8'd168,8'd170} : s = 338;
	{8'd168,8'd171} : s = 339;
	{8'd168,8'd172} : s = 340;
	{8'd168,8'd173} : s = 341;
	{8'd168,8'd174} : s = 342;
	{8'd168,8'd175} : s = 343;
	{8'd168,8'd176} : s = 344;
	{8'd168,8'd177} : s = 345;
	{8'd168,8'd178} : s = 346;
	{8'd168,8'd179} : s = 347;
	{8'd168,8'd180} : s = 348;
	{8'd168,8'd181} : s = 349;
	{8'd168,8'd182} : s = 350;
	{8'd168,8'd183} : s = 351;
	{8'd168,8'd184} : s = 352;
	{8'd168,8'd185} : s = 353;
	{8'd168,8'd186} : s = 354;
	{8'd168,8'd187} : s = 355;
	{8'd168,8'd188} : s = 356;
	{8'd168,8'd189} : s = 357;
	{8'd168,8'd190} : s = 358;
	{8'd168,8'd191} : s = 359;
	{8'd168,8'd192} : s = 360;
	{8'd168,8'd193} : s = 361;
	{8'd168,8'd194} : s = 362;
	{8'd168,8'd195} : s = 363;
	{8'd168,8'd196} : s = 364;
	{8'd168,8'd197} : s = 365;
	{8'd168,8'd198} : s = 366;
	{8'd168,8'd199} : s = 367;
	{8'd168,8'd200} : s = 368;
	{8'd168,8'd201} : s = 369;
	{8'd168,8'd202} : s = 370;
	{8'd168,8'd203} : s = 371;
	{8'd168,8'd204} : s = 372;
	{8'd168,8'd205} : s = 373;
	{8'd168,8'd206} : s = 374;
	{8'd168,8'd207} : s = 375;
	{8'd168,8'd208} : s = 376;
	{8'd168,8'd209} : s = 377;
	{8'd168,8'd210} : s = 378;
	{8'd168,8'd211} : s = 379;
	{8'd168,8'd212} : s = 380;
	{8'd168,8'd213} : s = 381;
	{8'd168,8'd214} : s = 382;
	{8'd168,8'd215} : s = 383;
	{8'd168,8'd216} : s = 384;
	{8'd168,8'd217} : s = 385;
	{8'd168,8'd218} : s = 386;
	{8'd168,8'd219} : s = 387;
	{8'd168,8'd220} : s = 388;
	{8'd168,8'd221} : s = 389;
	{8'd168,8'd222} : s = 390;
	{8'd168,8'd223} : s = 391;
	{8'd168,8'd224} : s = 392;
	{8'd168,8'd225} : s = 393;
	{8'd168,8'd226} : s = 394;
	{8'd168,8'd227} : s = 395;
	{8'd168,8'd228} : s = 396;
	{8'd168,8'd229} : s = 397;
	{8'd168,8'd230} : s = 398;
	{8'd168,8'd231} : s = 399;
	{8'd168,8'd232} : s = 400;
	{8'd168,8'd233} : s = 401;
	{8'd168,8'd234} : s = 402;
	{8'd168,8'd235} : s = 403;
	{8'd168,8'd236} : s = 404;
	{8'd168,8'd237} : s = 405;
	{8'd168,8'd238} : s = 406;
	{8'd168,8'd239} : s = 407;
	{8'd168,8'd240} : s = 408;
	{8'd168,8'd241} : s = 409;
	{8'd168,8'd242} : s = 410;
	{8'd168,8'd243} : s = 411;
	{8'd168,8'd244} : s = 412;
	{8'd168,8'd245} : s = 413;
	{8'd168,8'd246} : s = 414;
	{8'd168,8'd247} : s = 415;
	{8'd168,8'd248} : s = 416;
	{8'd168,8'd249} : s = 417;
	{8'd168,8'd250} : s = 418;
	{8'd168,8'd251} : s = 419;
	{8'd168,8'd252} : s = 420;
	{8'd168,8'd253} : s = 421;
	{8'd168,8'd254} : s = 422;
	{8'd168,8'd255} : s = 423;
	{8'd169,8'd0} : s = 169;
	{8'd169,8'd1} : s = 170;
	{8'd169,8'd2} : s = 171;
	{8'd169,8'd3} : s = 172;
	{8'd169,8'd4} : s = 173;
	{8'd169,8'd5} : s = 174;
	{8'd169,8'd6} : s = 175;
	{8'd169,8'd7} : s = 176;
	{8'd169,8'd8} : s = 177;
	{8'd169,8'd9} : s = 178;
	{8'd169,8'd10} : s = 179;
	{8'd169,8'd11} : s = 180;
	{8'd169,8'd12} : s = 181;
	{8'd169,8'd13} : s = 182;
	{8'd169,8'd14} : s = 183;
	{8'd169,8'd15} : s = 184;
	{8'd169,8'd16} : s = 185;
	{8'd169,8'd17} : s = 186;
	{8'd169,8'd18} : s = 187;
	{8'd169,8'd19} : s = 188;
	{8'd169,8'd20} : s = 189;
	{8'd169,8'd21} : s = 190;
	{8'd169,8'd22} : s = 191;
	{8'd169,8'd23} : s = 192;
	{8'd169,8'd24} : s = 193;
	{8'd169,8'd25} : s = 194;
	{8'd169,8'd26} : s = 195;
	{8'd169,8'd27} : s = 196;
	{8'd169,8'd28} : s = 197;
	{8'd169,8'd29} : s = 198;
	{8'd169,8'd30} : s = 199;
	{8'd169,8'd31} : s = 200;
	{8'd169,8'd32} : s = 201;
	{8'd169,8'd33} : s = 202;
	{8'd169,8'd34} : s = 203;
	{8'd169,8'd35} : s = 204;
	{8'd169,8'd36} : s = 205;
	{8'd169,8'd37} : s = 206;
	{8'd169,8'd38} : s = 207;
	{8'd169,8'd39} : s = 208;
	{8'd169,8'd40} : s = 209;
	{8'd169,8'd41} : s = 210;
	{8'd169,8'd42} : s = 211;
	{8'd169,8'd43} : s = 212;
	{8'd169,8'd44} : s = 213;
	{8'd169,8'd45} : s = 214;
	{8'd169,8'd46} : s = 215;
	{8'd169,8'd47} : s = 216;
	{8'd169,8'd48} : s = 217;
	{8'd169,8'd49} : s = 218;
	{8'd169,8'd50} : s = 219;
	{8'd169,8'd51} : s = 220;
	{8'd169,8'd52} : s = 221;
	{8'd169,8'd53} : s = 222;
	{8'd169,8'd54} : s = 223;
	{8'd169,8'd55} : s = 224;
	{8'd169,8'd56} : s = 225;
	{8'd169,8'd57} : s = 226;
	{8'd169,8'd58} : s = 227;
	{8'd169,8'd59} : s = 228;
	{8'd169,8'd60} : s = 229;
	{8'd169,8'd61} : s = 230;
	{8'd169,8'd62} : s = 231;
	{8'd169,8'd63} : s = 232;
	{8'd169,8'd64} : s = 233;
	{8'd169,8'd65} : s = 234;
	{8'd169,8'd66} : s = 235;
	{8'd169,8'd67} : s = 236;
	{8'd169,8'd68} : s = 237;
	{8'd169,8'd69} : s = 238;
	{8'd169,8'd70} : s = 239;
	{8'd169,8'd71} : s = 240;
	{8'd169,8'd72} : s = 241;
	{8'd169,8'd73} : s = 242;
	{8'd169,8'd74} : s = 243;
	{8'd169,8'd75} : s = 244;
	{8'd169,8'd76} : s = 245;
	{8'd169,8'd77} : s = 246;
	{8'd169,8'd78} : s = 247;
	{8'd169,8'd79} : s = 248;
	{8'd169,8'd80} : s = 249;
	{8'd169,8'd81} : s = 250;
	{8'd169,8'd82} : s = 251;
	{8'd169,8'd83} : s = 252;
	{8'd169,8'd84} : s = 253;
	{8'd169,8'd85} : s = 254;
	{8'd169,8'd86} : s = 255;
	{8'd169,8'd87} : s = 256;
	{8'd169,8'd88} : s = 257;
	{8'd169,8'd89} : s = 258;
	{8'd169,8'd90} : s = 259;
	{8'd169,8'd91} : s = 260;
	{8'd169,8'd92} : s = 261;
	{8'd169,8'd93} : s = 262;
	{8'd169,8'd94} : s = 263;
	{8'd169,8'd95} : s = 264;
	{8'd169,8'd96} : s = 265;
	{8'd169,8'd97} : s = 266;
	{8'd169,8'd98} : s = 267;
	{8'd169,8'd99} : s = 268;
	{8'd169,8'd100} : s = 269;
	{8'd169,8'd101} : s = 270;
	{8'd169,8'd102} : s = 271;
	{8'd169,8'd103} : s = 272;
	{8'd169,8'd104} : s = 273;
	{8'd169,8'd105} : s = 274;
	{8'd169,8'd106} : s = 275;
	{8'd169,8'd107} : s = 276;
	{8'd169,8'd108} : s = 277;
	{8'd169,8'd109} : s = 278;
	{8'd169,8'd110} : s = 279;
	{8'd169,8'd111} : s = 280;
	{8'd169,8'd112} : s = 281;
	{8'd169,8'd113} : s = 282;
	{8'd169,8'd114} : s = 283;
	{8'd169,8'd115} : s = 284;
	{8'd169,8'd116} : s = 285;
	{8'd169,8'd117} : s = 286;
	{8'd169,8'd118} : s = 287;
	{8'd169,8'd119} : s = 288;
	{8'd169,8'd120} : s = 289;
	{8'd169,8'd121} : s = 290;
	{8'd169,8'd122} : s = 291;
	{8'd169,8'd123} : s = 292;
	{8'd169,8'd124} : s = 293;
	{8'd169,8'd125} : s = 294;
	{8'd169,8'd126} : s = 295;
	{8'd169,8'd127} : s = 296;
	{8'd169,8'd128} : s = 297;
	{8'd169,8'd129} : s = 298;
	{8'd169,8'd130} : s = 299;
	{8'd169,8'd131} : s = 300;
	{8'd169,8'd132} : s = 301;
	{8'd169,8'd133} : s = 302;
	{8'd169,8'd134} : s = 303;
	{8'd169,8'd135} : s = 304;
	{8'd169,8'd136} : s = 305;
	{8'd169,8'd137} : s = 306;
	{8'd169,8'd138} : s = 307;
	{8'd169,8'd139} : s = 308;
	{8'd169,8'd140} : s = 309;
	{8'd169,8'd141} : s = 310;
	{8'd169,8'd142} : s = 311;
	{8'd169,8'd143} : s = 312;
	{8'd169,8'd144} : s = 313;
	{8'd169,8'd145} : s = 314;
	{8'd169,8'd146} : s = 315;
	{8'd169,8'd147} : s = 316;
	{8'd169,8'd148} : s = 317;
	{8'd169,8'd149} : s = 318;
	{8'd169,8'd150} : s = 319;
	{8'd169,8'd151} : s = 320;
	{8'd169,8'd152} : s = 321;
	{8'd169,8'd153} : s = 322;
	{8'd169,8'd154} : s = 323;
	{8'd169,8'd155} : s = 324;
	{8'd169,8'd156} : s = 325;
	{8'd169,8'd157} : s = 326;
	{8'd169,8'd158} : s = 327;
	{8'd169,8'd159} : s = 328;
	{8'd169,8'd160} : s = 329;
	{8'd169,8'd161} : s = 330;
	{8'd169,8'd162} : s = 331;
	{8'd169,8'd163} : s = 332;
	{8'd169,8'd164} : s = 333;
	{8'd169,8'd165} : s = 334;
	{8'd169,8'd166} : s = 335;
	{8'd169,8'd167} : s = 336;
	{8'd169,8'd168} : s = 337;
	{8'd169,8'd169} : s = 338;
	{8'd169,8'd170} : s = 339;
	{8'd169,8'd171} : s = 340;
	{8'd169,8'd172} : s = 341;
	{8'd169,8'd173} : s = 342;
	{8'd169,8'd174} : s = 343;
	{8'd169,8'd175} : s = 344;
	{8'd169,8'd176} : s = 345;
	{8'd169,8'd177} : s = 346;
	{8'd169,8'd178} : s = 347;
	{8'd169,8'd179} : s = 348;
	{8'd169,8'd180} : s = 349;
	{8'd169,8'd181} : s = 350;
	{8'd169,8'd182} : s = 351;
	{8'd169,8'd183} : s = 352;
	{8'd169,8'd184} : s = 353;
	{8'd169,8'd185} : s = 354;
	{8'd169,8'd186} : s = 355;
	{8'd169,8'd187} : s = 356;
	{8'd169,8'd188} : s = 357;
	{8'd169,8'd189} : s = 358;
	{8'd169,8'd190} : s = 359;
	{8'd169,8'd191} : s = 360;
	{8'd169,8'd192} : s = 361;
	{8'd169,8'd193} : s = 362;
	{8'd169,8'd194} : s = 363;
	{8'd169,8'd195} : s = 364;
	{8'd169,8'd196} : s = 365;
	{8'd169,8'd197} : s = 366;
	{8'd169,8'd198} : s = 367;
	{8'd169,8'd199} : s = 368;
	{8'd169,8'd200} : s = 369;
	{8'd169,8'd201} : s = 370;
	{8'd169,8'd202} : s = 371;
	{8'd169,8'd203} : s = 372;
	{8'd169,8'd204} : s = 373;
	{8'd169,8'd205} : s = 374;
	{8'd169,8'd206} : s = 375;
	{8'd169,8'd207} : s = 376;
	{8'd169,8'd208} : s = 377;
	{8'd169,8'd209} : s = 378;
	{8'd169,8'd210} : s = 379;
	{8'd169,8'd211} : s = 380;
	{8'd169,8'd212} : s = 381;
	{8'd169,8'd213} : s = 382;
	{8'd169,8'd214} : s = 383;
	{8'd169,8'd215} : s = 384;
	{8'd169,8'd216} : s = 385;
	{8'd169,8'd217} : s = 386;
	{8'd169,8'd218} : s = 387;
	{8'd169,8'd219} : s = 388;
	{8'd169,8'd220} : s = 389;
	{8'd169,8'd221} : s = 390;
	{8'd169,8'd222} : s = 391;
	{8'd169,8'd223} : s = 392;
	{8'd169,8'd224} : s = 393;
	{8'd169,8'd225} : s = 394;
	{8'd169,8'd226} : s = 395;
	{8'd169,8'd227} : s = 396;
	{8'd169,8'd228} : s = 397;
	{8'd169,8'd229} : s = 398;
	{8'd169,8'd230} : s = 399;
	{8'd169,8'd231} : s = 400;
	{8'd169,8'd232} : s = 401;
	{8'd169,8'd233} : s = 402;
	{8'd169,8'd234} : s = 403;
	{8'd169,8'd235} : s = 404;
	{8'd169,8'd236} : s = 405;
	{8'd169,8'd237} : s = 406;
	{8'd169,8'd238} : s = 407;
	{8'd169,8'd239} : s = 408;
	{8'd169,8'd240} : s = 409;
	{8'd169,8'd241} : s = 410;
	{8'd169,8'd242} : s = 411;
	{8'd169,8'd243} : s = 412;
	{8'd169,8'd244} : s = 413;
	{8'd169,8'd245} : s = 414;
	{8'd169,8'd246} : s = 415;
	{8'd169,8'd247} : s = 416;
	{8'd169,8'd248} : s = 417;
	{8'd169,8'd249} : s = 418;
	{8'd169,8'd250} : s = 419;
	{8'd169,8'd251} : s = 420;
	{8'd169,8'd252} : s = 421;
	{8'd169,8'd253} : s = 422;
	{8'd169,8'd254} : s = 423;
	{8'd169,8'd255} : s = 424;
	{8'd170,8'd0} : s = 170;
	{8'd170,8'd1} : s = 171;
	{8'd170,8'd2} : s = 172;
	{8'd170,8'd3} : s = 173;
	{8'd170,8'd4} : s = 174;
	{8'd170,8'd5} : s = 175;
	{8'd170,8'd6} : s = 176;
	{8'd170,8'd7} : s = 177;
	{8'd170,8'd8} : s = 178;
	{8'd170,8'd9} : s = 179;
	{8'd170,8'd10} : s = 180;
	{8'd170,8'd11} : s = 181;
	{8'd170,8'd12} : s = 182;
	{8'd170,8'd13} : s = 183;
	{8'd170,8'd14} : s = 184;
	{8'd170,8'd15} : s = 185;
	{8'd170,8'd16} : s = 186;
	{8'd170,8'd17} : s = 187;
	{8'd170,8'd18} : s = 188;
	{8'd170,8'd19} : s = 189;
	{8'd170,8'd20} : s = 190;
	{8'd170,8'd21} : s = 191;
	{8'd170,8'd22} : s = 192;
	{8'd170,8'd23} : s = 193;
	{8'd170,8'd24} : s = 194;
	{8'd170,8'd25} : s = 195;
	{8'd170,8'd26} : s = 196;
	{8'd170,8'd27} : s = 197;
	{8'd170,8'd28} : s = 198;
	{8'd170,8'd29} : s = 199;
	{8'd170,8'd30} : s = 200;
	{8'd170,8'd31} : s = 201;
	{8'd170,8'd32} : s = 202;
	{8'd170,8'd33} : s = 203;
	{8'd170,8'd34} : s = 204;
	{8'd170,8'd35} : s = 205;
	{8'd170,8'd36} : s = 206;
	{8'd170,8'd37} : s = 207;
	{8'd170,8'd38} : s = 208;
	{8'd170,8'd39} : s = 209;
	{8'd170,8'd40} : s = 210;
	{8'd170,8'd41} : s = 211;
	{8'd170,8'd42} : s = 212;
	{8'd170,8'd43} : s = 213;
	{8'd170,8'd44} : s = 214;
	{8'd170,8'd45} : s = 215;
	{8'd170,8'd46} : s = 216;
	{8'd170,8'd47} : s = 217;
	{8'd170,8'd48} : s = 218;
	{8'd170,8'd49} : s = 219;
	{8'd170,8'd50} : s = 220;
	{8'd170,8'd51} : s = 221;
	{8'd170,8'd52} : s = 222;
	{8'd170,8'd53} : s = 223;
	{8'd170,8'd54} : s = 224;
	{8'd170,8'd55} : s = 225;
	{8'd170,8'd56} : s = 226;
	{8'd170,8'd57} : s = 227;
	{8'd170,8'd58} : s = 228;
	{8'd170,8'd59} : s = 229;
	{8'd170,8'd60} : s = 230;
	{8'd170,8'd61} : s = 231;
	{8'd170,8'd62} : s = 232;
	{8'd170,8'd63} : s = 233;
	{8'd170,8'd64} : s = 234;
	{8'd170,8'd65} : s = 235;
	{8'd170,8'd66} : s = 236;
	{8'd170,8'd67} : s = 237;
	{8'd170,8'd68} : s = 238;
	{8'd170,8'd69} : s = 239;
	{8'd170,8'd70} : s = 240;
	{8'd170,8'd71} : s = 241;
	{8'd170,8'd72} : s = 242;
	{8'd170,8'd73} : s = 243;
	{8'd170,8'd74} : s = 244;
	{8'd170,8'd75} : s = 245;
	{8'd170,8'd76} : s = 246;
	{8'd170,8'd77} : s = 247;
	{8'd170,8'd78} : s = 248;
	{8'd170,8'd79} : s = 249;
	{8'd170,8'd80} : s = 250;
	{8'd170,8'd81} : s = 251;
	{8'd170,8'd82} : s = 252;
	{8'd170,8'd83} : s = 253;
	{8'd170,8'd84} : s = 254;
	{8'd170,8'd85} : s = 255;
	{8'd170,8'd86} : s = 256;
	{8'd170,8'd87} : s = 257;
	{8'd170,8'd88} : s = 258;
	{8'd170,8'd89} : s = 259;
	{8'd170,8'd90} : s = 260;
	{8'd170,8'd91} : s = 261;
	{8'd170,8'd92} : s = 262;
	{8'd170,8'd93} : s = 263;
	{8'd170,8'd94} : s = 264;
	{8'd170,8'd95} : s = 265;
	{8'd170,8'd96} : s = 266;
	{8'd170,8'd97} : s = 267;
	{8'd170,8'd98} : s = 268;
	{8'd170,8'd99} : s = 269;
	{8'd170,8'd100} : s = 270;
	{8'd170,8'd101} : s = 271;
	{8'd170,8'd102} : s = 272;
	{8'd170,8'd103} : s = 273;
	{8'd170,8'd104} : s = 274;
	{8'd170,8'd105} : s = 275;
	{8'd170,8'd106} : s = 276;
	{8'd170,8'd107} : s = 277;
	{8'd170,8'd108} : s = 278;
	{8'd170,8'd109} : s = 279;
	{8'd170,8'd110} : s = 280;
	{8'd170,8'd111} : s = 281;
	{8'd170,8'd112} : s = 282;
	{8'd170,8'd113} : s = 283;
	{8'd170,8'd114} : s = 284;
	{8'd170,8'd115} : s = 285;
	{8'd170,8'd116} : s = 286;
	{8'd170,8'd117} : s = 287;
	{8'd170,8'd118} : s = 288;
	{8'd170,8'd119} : s = 289;
	{8'd170,8'd120} : s = 290;
	{8'd170,8'd121} : s = 291;
	{8'd170,8'd122} : s = 292;
	{8'd170,8'd123} : s = 293;
	{8'd170,8'd124} : s = 294;
	{8'd170,8'd125} : s = 295;
	{8'd170,8'd126} : s = 296;
	{8'd170,8'd127} : s = 297;
	{8'd170,8'd128} : s = 298;
	{8'd170,8'd129} : s = 299;
	{8'd170,8'd130} : s = 300;
	{8'd170,8'd131} : s = 301;
	{8'd170,8'd132} : s = 302;
	{8'd170,8'd133} : s = 303;
	{8'd170,8'd134} : s = 304;
	{8'd170,8'd135} : s = 305;
	{8'd170,8'd136} : s = 306;
	{8'd170,8'd137} : s = 307;
	{8'd170,8'd138} : s = 308;
	{8'd170,8'd139} : s = 309;
	{8'd170,8'd140} : s = 310;
	{8'd170,8'd141} : s = 311;
	{8'd170,8'd142} : s = 312;
	{8'd170,8'd143} : s = 313;
	{8'd170,8'd144} : s = 314;
	{8'd170,8'd145} : s = 315;
	{8'd170,8'd146} : s = 316;
	{8'd170,8'd147} : s = 317;
	{8'd170,8'd148} : s = 318;
	{8'd170,8'd149} : s = 319;
	{8'd170,8'd150} : s = 320;
	{8'd170,8'd151} : s = 321;
	{8'd170,8'd152} : s = 322;
	{8'd170,8'd153} : s = 323;
	{8'd170,8'd154} : s = 324;
	{8'd170,8'd155} : s = 325;
	{8'd170,8'd156} : s = 326;
	{8'd170,8'd157} : s = 327;
	{8'd170,8'd158} : s = 328;
	{8'd170,8'd159} : s = 329;
	{8'd170,8'd160} : s = 330;
	{8'd170,8'd161} : s = 331;
	{8'd170,8'd162} : s = 332;
	{8'd170,8'd163} : s = 333;
	{8'd170,8'd164} : s = 334;
	{8'd170,8'd165} : s = 335;
	{8'd170,8'd166} : s = 336;
	{8'd170,8'd167} : s = 337;
	{8'd170,8'd168} : s = 338;
	{8'd170,8'd169} : s = 339;
	{8'd170,8'd170} : s = 340;
	{8'd170,8'd171} : s = 341;
	{8'd170,8'd172} : s = 342;
	{8'd170,8'd173} : s = 343;
	{8'd170,8'd174} : s = 344;
	{8'd170,8'd175} : s = 345;
	{8'd170,8'd176} : s = 346;
	{8'd170,8'd177} : s = 347;
	{8'd170,8'd178} : s = 348;
	{8'd170,8'd179} : s = 349;
	{8'd170,8'd180} : s = 350;
	{8'd170,8'd181} : s = 351;
	{8'd170,8'd182} : s = 352;
	{8'd170,8'd183} : s = 353;
	{8'd170,8'd184} : s = 354;
	{8'd170,8'd185} : s = 355;
	{8'd170,8'd186} : s = 356;
	{8'd170,8'd187} : s = 357;
	{8'd170,8'd188} : s = 358;
	{8'd170,8'd189} : s = 359;
	{8'd170,8'd190} : s = 360;
	{8'd170,8'd191} : s = 361;
	{8'd170,8'd192} : s = 362;
	{8'd170,8'd193} : s = 363;
	{8'd170,8'd194} : s = 364;
	{8'd170,8'd195} : s = 365;
	{8'd170,8'd196} : s = 366;
	{8'd170,8'd197} : s = 367;
	{8'd170,8'd198} : s = 368;
	{8'd170,8'd199} : s = 369;
	{8'd170,8'd200} : s = 370;
	{8'd170,8'd201} : s = 371;
	{8'd170,8'd202} : s = 372;
	{8'd170,8'd203} : s = 373;
	{8'd170,8'd204} : s = 374;
	{8'd170,8'd205} : s = 375;
	{8'd170,8'd206} : s = 376;
	{8'd170,8'd207} : s = 377;
	{8'd170,8'd208} : s = 378;
	{8'd170,8'd209} : s = 379;
	{8'd170,8'd210} : s = 380;
	{8'd170,8'd211} : s = 381;
	{8'd170,8'd212} : s = 382;
	{8'd170,8'd213} : s = 383;
	{8'd170,8'd214} : s = 384;
	{8'd170,8'd215} : s = 385;
	{8'd170,8'd216} : s = 386;
	{8'd170,8'd217} : s = 387;
	{8'd170,8'd218} : s = 388;
	{8'd170,8'd219} : s = 389;
	{8'd170,8'd220} : s = 390;
	{8'd170,8'd221} : s = 391;
	{8'd170,8'd222} : s = 392;
	{8'd170,8'd223} : s = 393;
	{8'd170,8'd224} : s = 394;
	{8'd170,8'd225} : s = 395;
	{8'd170,8'd226} : s = 396;
	{8'd170,8'd227} : s = 397;
	{8'd170,8'd228} : s = 398;
	{8'd170,8'd229} : s = 399;
	{8'd170,8'd230} : s = 400;
	{8'd170,8'd231} : s = 401;
	{8'd170,8'd232} : s = 402;
	{8'd170,8'd233} : s = 403;
	{8'd170,8'd234} : s = 404;
	{8'd170,8'd235} : s = 405;
	{8'd170,8'd236} : s = 406;
	{8'd170,8'd237} : s = 407;
	{8'd170,8'd238} : s = 408;
	{8'd170,8'd239} : s = 409;
	{8'd170,8'd240} : s = 410;
	{8'd170,8'd241} : s = 411;
	{8'd170,8'd242} : s = 412;
	{8'd170,8'd243} : s = 413;
	{8'd170,8'd244} : s = 414;
	{8'd170,8'd245} : s = 415;
	{8'd170,8'd246} : s = 416;
	{8'd170,8'd247} : s = 417;
	{8'd170,8'd248} : s = 418;
	{8'd170,8'd249} : s = 419;
	{8'd170,8'd250} : s = 420;
	{8'd170,8'd251} : s = 421;
	{8'd170,8'd252} : s = 422;
	{8'd170,8'd253} : s = 423;
	{8'd170,8'd254} : s = 424;
	{8'd170,8'd255} : s = 425;
	{8'd171,8'd0} : s = 171;
	{8'd171,8'd1} : s = 172;
	{8'd171,8'd2} : s = 173;
	{8'd171,8'd3} : s = 174;
	{8'd171,8'd4} : s = 175;
	{8'd171,8'd5} : s = 176;
	{8'd171,8'd6} : s = 177;
	{8'd171,8'd7} : s = 178;
	{8'd171,8'd8} : s = 179;
	{8'd171,8'd9} : s = 180;
	{8'd171,8'd10} : s = 181;
	{8'd171,8'd11} : s = 182;
	{8'd171,8'd12} : s = 183;
	{8'd171,8'd13} : s = 184;
	{8'd171,8'd14} : s = 185;
	{8'd171,8'd15} : s = 186;
	{8'd171,8'd16} : s = 187;
	{8'd171,8'd17} : s = 188;
	{8'd171,8'd18} : s = 189;
	{8'd171,8'd19} : s = 190;
	{8'd171,8'd20} : s = 191;
	{8'd171,8'd21} : s = 192;
	{8'd171,8'd22} : s = 193;
	{8'd171,8'd23} : s = 194;
	{8'd171,8'd24} : s = 195;
	{8'd171,8'd25} : s = 196;
	{8'd171,8'd26} : s = 197;
	{8'd171,8'd27} : s = 198;
	{8'd171,8'd28} : s = 199;
	{8'd171,8'd29} : s = 200;
	{8'd171,8'd30} : s = 201;
	{8'd171,8'd31} : s = 202;
	{8'd171,8'd32} : s = 203;
	{8'd171,8'd33} : s = 204;
	{8'd171,8'd34} : s = 205;
	{8'd171,8'd35} : s = 206;
	{8'd171,8'd36} : s = 207;
	{8'd171,8'd37} : s = 208;
	{8'd171,8'd38} : s = 209;
	{8'd171,8'd39} : s = 210;
	{8'd171,8'd40} : s = 211;
	{8'd171,8'd41} : s = 212;
	{8'd171,8'd42} : s = 213;
	{8'd171,8'd43} : s = 214;
	{8'd171,8'd44} : s = 215;
	{8'd171,8'd45} : s = 216;
	{8'd171,8'd46} : s = 217;
	{8'd171,8'd47} : s = 218;
	{8'd171,8'd48} : s = 219;
	{8'd171,8'd49} : s = 220;
	{8'd171,8'd50} : s = 221;
	{8'd171,8'd51} : s = 222;
	{8'd171,8'd52} : s = 223;
	{8'd171,8'd53} : s = 224;
	{8'd171,8'd54} : s = 225;
	{8'd171,8'd55} : s = 226;
	{8'd171,8'd56} : s = 227;
	{8'd171,8'd57} : s = 228;
	{8'd171,8'd58} : s = 229;
	{8'd171,8'd59} : s = 230;
	{8'd171,8'd60} : s = 231;
	{8'd171,8'd61} : s = 232;
	{8'd171,8'd62} : s = 233;
	{8'd171,8'd63} : s = 234;
	{8'd171,8'd64} : s = 235;
	{8'd171,8'd65} : s = 236;
	{8'd171,8'd66} : s = 237;
	{8'd171,8'd67} : s = 238;
	{8'd171,8'd68} : s = 239;
	{8'd171,8'd69} : s = 240;
	{8'd171,8'd70} : s = 241;
	{8'd171,8'd71} : s = 242;
	{8'd171,8'd72} : s = 243;
	{8'd171,8'd73} : s = 244;
	{8'd171,8'd74} : s = 245;
	{8'd171,8'd75} : s = 246;
	{8'd171,8'd76} : s = 247;
	{8'd171,8'd77} : s = 248;
	{8'd171,8'd78} : s = 249;
	{8'd171,8'd79} : s = 250;
	{8'd171,8'd80} : s = 251;
	{8'd171,8'd81} : s = 252;
	{8'd171,8'd82} : s = 253;
	{8'd171,8'd83} : s = 254;
	{8'd171,8'd84} : s = 255;
	{8'd171,8'd85} : s = 256;
	{8'd171,8'd86} : s = 257;
	{8'd171,8'd87} : s = 258;
	{8'd171,8'd88} : s = 259;
	{8'd171,8'd89} : s = 260;
	{8'd171,8'd90} : s = 261;
	{8'd171,8'd91} : s = 262;
	{8'd171,8'd92} : s = 263;
	{8'd171,8'd93} : s = 264;
	{8'd171,8'd94} : s = 265;
	{8'd171,8'd95} : s = 266;
	{8'd171,8'd96} : s = 267;
	{8'd171,8'd97} : s = 268;
	{8'd171,8'd98} : s = 269;
	{8'd171,8'd99} : s = 270;
	{8'd171,8'd100} : s = 271;
	{8'd171,8'd101} : s = 272;
	{8'd171,8'd102} : s = 273;
	{8'd171,8'd103} : s = 274;
	{8'd171,8'd104} : s = 275;
	{8'd171,8'd105} : s = 276;
	{8'd171,8'd106} : s = 277;
	{8'd171,8'd107} : s = 278;
	{8'd171,8'd108} : s = 279;
	{8'd171,8'd109} : s = 280;
	{8'd171,8'd110} : s = 281;
	{8'd171,8'd111} : s = 282;
	{8'd171,8'd112} : s = 283;
	{8'd171,8'd113} : s = 284;
	{8'd171,8'd114} : s = 285;
	{8'd171,8'd115} : s = 286;
	{8'd171,8'd116} : s = 287;
	{8'd171,8'd117} : s = 288;
	{8'd171,8'd118} : s = 289;
	{8'd171,8'd119} : s = 290;
	{8'd171,8'd120} : s = 291;
	{8'd171,8'd121} : s = 292;
	{8'd171,8'd122} : s = 293;
	{8'd171,8'd123} : s = 294;
	{8'd171,8'd124} : s = 295;
	{8'd171,8'd125} : s = 296;
	{8'd171,8'd126} : s = 297;
	{8'd171,8'd127} : s = 298;
	{8'd171,8'd128} : s = 299;
	{8'd171,8'd129} : s = 300;
	{8'd171,8'd130} : s = 301;
	{8'd171,8'd131} : s = 302;
	{8'd171,8'd132} : s = 303;
	{8'd171,8'd133} : s = 304;
	{8'd171,8'd134} : s = 305;
	{8'd171,8'd135} : s = 306;
	{8'd171,8'd136} : s = 307;
	{8'd171,8'd137} : s = 308;
	{8'd171,8'd138} : s = 309;
	{8'd171,8'd139} : s = 310;
	{8'd171,8'd140} : s = 311;
	{8'd171,8'd141} : s = 312;
	{8'd171,8'd142} : s = 313;
	{8'd171,8'd143} : s = 314;
	{8'd171,8'd144} : s = 315;
	{8'd171,8'd145} : s = 316;
	{8'd171,8'd146} : s = 317;
	{8'd171,8'd147} : s = 318;
	{8'd171,8'd148} : s = 319;
	{8'd171,8'd149} : s = 320;
	{8'd171,8'd150} : s = 321;
	{8'd171,8'd151} : s = 322;
	{8'd171,8'd152} : s = 323;
	{8'd171,8'd153} : s = 324;
	{8'd171,8'd154} : s = 325;
	{8'd171,8'd155} : s = 326;
	{8'd171,8'd156} : s = 327;
	{8'd171,8'd157} : s = 328;
	{8'd171,8'd158} : s = 329;
	{8'd171,8'd159} : s = 330;
	{8'd171,8'd160} : s = 331;
	{8'd171,8'd161} : s = 332;
	{8'd171,8'd162} : s = 333;
	{8'd171,8'd163} : s = 334;
	{8'd171,8'd164} : s = 335;
	{8'd171,8'd165} : s = 336;
	{8'd171,8'd166} : s = 337;
	{8'd171,8'd167} : s = 338;
	{8'd171,8'd168} : s = 339;
	{8'd171,8'd169} : s = 340;
	{8'd171,8'd170} : s = 341;
	{8'd171,8'd171} : s = 342;
	{8'd171,8'd172} : s = 343;
	{8'd171,8'd173} : s = 344;
	{8'd171,8'd174} : s = 345;
	{8'd171,8'd175} : s = 346;
	{8'd171,8'd176} : s = 347;
	{8'd171,8'd177} : s = 348;
	{8'd171,8'd178} : s = 349;
	{8'd171,8'd179} : s = 350;
	{8'd171,8'd180} : s = 351;
	{8'd171,8'd181} : s = 352;
	{8'd171,8'd182} : s = 353;
	{8'd171,8'd183} : s = 354;
	{8'd171,8'd184} : s = 355;
	{8'd171,8'd185} : s = 356;
	{8'd171,8'd186} : s = 357;
	{8'd171,8'd187} : s = 358;
	{8'd171,8'd188} : s = 359;
	{8'd171,8'd189} : s = 360;
	{8'd171,8'd190} : s = 361;
	{8'd171,8'd191} : s = 362;
	{8'd171,8'd192} : s = 363;
	{8'd171,8'd193} : s = 364;
	{8'd171,8'd194} : s = 365;
	{8'd171,8'd195} : s = 366;
	{8'd171,8'd196} : s = 367;
	{8'd171,8'd197} : s = 368;
	{8'd171,8'd198} : s = 369;
	{8'd171,8'd199} : s = 370;
	{8'd171,8'd200} : s = 371;
	{8'd171,8'd201} : s = 372;
	{8'd171,8'd202} : s = 373;
	{8'd171,8'd203} : s = 374;
	{8'd171,8'd204} : s = 375;
	{8'd171,8'd205} : s = 376;
	{8'd171,8'd206} : s = 377;
	{8'd171,8'd207} : s = 378;
	{8'd171,8'd208} : s = 379;
	{8'd171,8'd209} : s = 380;
	{8'd171,8'd210} : s = 381;
	{8'd171,8'd211} : s = 382;
	{8'd171,8'd212} : s = 383;
	{8'd171,8'd213} : s = 384;
	{8'd171,8'd214} : s = 385;
	{8'd171,8'd215} : s = 386;
	{8'd171,8'd216} : s = 387;
	{8'd171,8'd217} : s = 388;
	{8'd171,8'd218} : s = 389;
	{8'd171,8'd219} : s = 390;
	{8'd171,8'd220} : s = 391;
	{8'd171,8'd221} : s = 392;
	{8'd171,8'd222} : s = 393;
	{8'd171,8'd223} : s = 394;
	{8'd171,8'd224} : s = 395;
	{8'd171,8'd225} : s = 396;
	{8'd171,8'd226} : s = 397;
	{8'd171,8'd227} : s = 398;
	{8'd171,8'd228} : s = 399;
	{8'd171,8'd229} : s = 400;
	{8'd171,8'd230} : s = 401;
	{8'd171,8'd231} : s = 402;
	{8'd171,8'd232} : s = 403;
	{8'd171,8'd233} : s = 404;
	{8'd171,8'd234} : s = 405;
	{8'd171,8'd235} : s = 406;
	{8'd171,8'd236} : s = 407;
	{8'd171,8'd237} : s = 408;
	{8'd171,8'd238} : s = 409;
	{8'd171,8'd239} : s = 410;
	{8'd171,8'd240} : s = 411;
	{8'd171,8'd241} : s = 412;
	{8'd171,8'd242} : s = 413;
	{8'd171,8'd243} : s = 414;
	{8'd171,8'd244} : s = 415;
	{8'd171,8'd245} : s = 416;
	{8'd171,8'd246} : s = 417;
	{8'd171,8'd247} : s = 418;
	{8'd171,8'd248} : s = 419;
	{8'd171,8'd249} : s = 420;
	{8'd171,8'd250} : s = 421;
	{8'd171,8'd251} : s = 422;
	{8'd171,8'd252} : s = 423;
	{8'd171,8'd253} : s = 424;
	{8'd171,8'd254} : s = 425;
	{8'd171,8'd255} : s = 426;
	{8'd172,8'd0} : s = 172;
	{8'd172,8'd1} : s = 173;
	{8'd172,8'd2} : s = 174;
	{8'd172,8'd3} : s = 175;
	{8'd172,8'd4} : s = 176;
	{8'd172,8'd5} : s = 177;
	{8'd172,8'd6} : s = 178;
	{8'd172,8'd7} : s = 179;
	{8'd172,8'd8} : s = 180;
	{8'd172,8'd9} : s = 181;
	{8'd172,8'd10} : s = 182;
	{8'd172,8'd11} : s = 183;
	{8'd172,8'd12} : s = 184;
	{8'd172,8'd13} : s = 185;
	{8'd172,8'd14} : s = 186;
	{8'd172,8'd15} : s = 187;
	{8'd172,8'd16} : s = 188;
	{8'd172,8'd17} : s = 189;
	{8'd172,8'd18} : s = 190;
	{8'd172,8'd19} : s = 191;
	{8'd172,8'd20} : s = 192;
	{8'd172,8'd21} : s = 193;
	{8'd172,8'd22} : s = 194;
	{8'd172,8'd23} : s = 195;
	{8'd172,8'd24} : s = 196;
	{8'd172,8'd25} : s = 197;
	{8'd172,8'd26} : s = 198;
	{8'd172,8'd27} : s = 199;
	{8'd172,8'd28} : s = 200;
	{8'd172,8'd29} : s = 201;
	{8'd172,8'd30} : s = 202;
	{8'd172,8'd31} : s = 203;
	{8'd172,8'd32} : s = 204;
	{8'd172,8'd33} : s = 205;
	{8'd172,8'd34} : s = 206;
	{8'd172,8'd35} : s = 207;
	{8'd172,8'd36} : s = 208;
	{8'd172,8'd37} : s = 209;
	{8'd172,8'd38} : s = 210;
	{8'd172,8'd39} : s = 211;
	{8'd172,8'd40} : s = 212;
	{8'd172,8'd41} : s = 213;
	{8'd172,8'd42} : s = 214;
	{8'd172,8'd43} : s = 215;
	{8'd172,8'd44} : s = 216;
	{8'd172,8'd45} : s = 217;
	{8'd172,8'd46} : s = 218;
	{8'd172,8'd47} : s = 219;
	{8'd172,8'd48} : s = 220;
	{8'd172,8'd49} : s = 221;
	{8'd172,8'd50} : s = 222;
	{8'd172,8'd51} : s = 223;
	{8'd172,8'd52} : s = 224;
	{8'd172,8'd53} : s = 225;
	{8'd172,8'd54} : s = 226;
	{8'd172,8'd55} : s = 227;
	{8'd172,8'd56} : s = 228;
	{8'd172,8'd57} : s = 229;
	{8'd172,8'd58} : s = 230;
	{8'd172,8'd59} : s = 231;
	{8'd172,8'd60} : s = 232;
	{8'd172,8'd61} : s = 233;
	{8'd172,8'd62} : s = 234;
	{8'd172,8'd63} : s = 235;
	{8'd172,8'd64} : s = 236;
	{8'd172,8'd65} : s = 237;
	{8'd172,8'd66} : s = 238;
	{8'd172,8'd67} : s = 239;
	{8'd172,8'd68} : s = 240;
	{8'd172,8'd69} : s = 241;
	{8'd172,8'd70} : s = 242;
	{8'd172,8'd71} : s = 243;
	{8'd172,8'd72} : s = 244;
	{8'd172,8'd73} : s = 245;
	{8'd172,8'd74} : s = 246;
	{8'd172,8'd75} : s = 247;
	{8'd172,8'd76} : s = 248;
	{8'd172,8'd77} : s = 249;
	{8'd172,8'd78} : s = 250;
	{8'd172,8'd79} : s = 251;
	{8'd172,8'd80} : s = 252;
	{8'd172,8'd81} : s = 253;
	{8'd172,8'd82} : s = 254;
	{8'd172,8'd83} : s = 255;
	{8'd172,8'd84} : s = 256;
	{8'd172,8'd85} : s = 257;
	{8'd172,8'd86} : s = 258;
	{8'd172,8'd87} : s = 259;
	{8'd172,8'd88} : s = 260;
	{8'd172,8'd89} : s = 261;
	{8'd172,8'd90} : s = 262;
	{8'd172,8'd91} : s = 263;
	{8'd172,8'd92} : s = 264;
	{8'd172,8'd93} : s = 265;
	{8'd172,8'd94} : s = 266;
	{8'd172,8'd95} : s = 267;
	{8'd172,8'd96} : s = 268;
	{8'd172,8'd97} : s = 269;
	{8'd172,8'd98} : s = 270;
	{8'd172,8'd99} : s = 271;
	{8'd172,8'd100} : s = 272;
	{8'd172,8'd101} : s = 273;
	{8'd172,8'd102} : s = 274;
	{8'd172,8'd103} : s = 275;
	{8'd172,8'd104} : s = 276;
	{8'd172,8'd105} : s = 277;
	{8'd172,8'd106} : s = 278;
	{8'd172,8'd107} : s = 279;
	{8'd172,8'd108} : s = 280;
	{8'd172,8'd109} : s = 281;
	{8'd172,8'd110} : s = 282;
	{8'd172,8'd111} : s = 283;
	{8'd172,8'd112} : s = 284;
	{8'd172,8'd113} : s = 285;
	{8'd172,8'd114} : s = 286;
	{8'd172,8'd115} : s = 287;
	{8'd172,8'd116} : s = 288;
	{8'd172,8'd117} : s = 289;
	{8'd172,8'd118} : s = 290;
	{8'd172,8'd119} : s = 291;
	{8'd172,8'd120} : s = 292;
	{8'd172,8'd121} : s = 293;
	{8'd172,8'd122} : s = 294;
	{8'd172,8'd123} : s = 295;
	{8'd172,8'd124} : s = 296;
	{8'd172,8'd125} : s = 297;
	{8'd172,8'd126} : s = 298;
	{8'd172,8'd127} : s = 299;
	{8'd172,8'd128} : s = 300;
	{8'd172,8'd129} : s = 301;
	{8'd172,8'd130} : s = 302;
	{8'd172,8'd131} : s = 303;
	{8'd172,8'd132} : s = 304;
	{8'd172,8'd133} : s = 305;
	{8'd172,8'd134} : s = 306;
	{8'd172,8'd135} : s = 307;
	{8'd172,8'd136} : s = 308;
	{8'd172,8'd137} : s = 309;
	{8'd172,8'd138} : s = 310;
	{8'd172,8'd139} : s = 311;
	{8'd172,8'd140} : s = 312;
	{8'd172,8'd141} : s = 313;
	{8'd172,8'd142} : s = 314;
	{8'd172,8'd143} : s = 315;
	{8'd172,8'd144} : s = 316;
	{8'd172,8'd145} : s = 317;
	{8'd172,8'd146} : s = 318;
	{8'd172,8'd147} : s = 319;
	{8'd172,8'd148} : s = 320;
	{8'd172,8'd149} : s = 321;
	{8'd172,8'd150} : s = 322;
	{8'd172,8'd151} : s = 323;
	{8'd172,8'd152} : s = 324;
	{8'd172,8'd153} : s = 325;
	{8'd172,8'd154} : s = 326;
	{8'd172,8'd155} : s = 327;
	{8'd172,8'd156} : s = 328;
	{8'd172,8'd157} : s = 329;
	{8'd172,8'd158} : s = 330;
	{8'd172,8'd159} : s = 331;
	{8'd172,8'd160} : s = 332;
	{8'd172,8'd161} : s = 333;
	{8'd172,8'd162} : s = 334;
	{8'd172,8'd163} : s = 335;
	{8'd172,8'd164} : s = 336;
	{8'd172,8'd165} : s = 337;
	{8'd172,8'd166} : s = 338;
	{8'd172,8'd167} : s = 339;
	{8'd172,8'd168} : s = 340;
	{8'd172,8'd169} : s = 341;
	{8'd172,8'd170} : s = 342;
	{8'd172,8'd171} : s = 343;
	{8'd172,8'd172} : s = 344;
	{8'd172,8'd173} : s = 345;
	{8'd172,8'd174} : s = 346;
	{8'd172,8'd175} : s = 347;
	{8'd172,8'd176} : s = 348;
	{8'd172,8'd177} : s = 349;
	{8'd172,8'd178} : s = 350;
	{8'd172,8'd179} : s = 351;
	{8'd172,8'd180} : s = 352;
	{8'd172,8'd181} : s = 353;
	{8'd172,8'd182} : s = 354;
	{8'd172,8'd183} : s = 355;
	{8'd172,8'd184} : s = 356;
	{8'd172,8'd185} : s = 357;
	{8'd172,8'd186} : s = 358;
	{8'd172,8'd187} : s = 359;
	{8'd172,8'd188} : s = 360;
	{8'd172,8'd189} : s = 361;
	{8'd172,8'd190} : s = 362;
	{8'd172,8'd191} : s = 363;
	{8'd172,8'd192} : s = 364;
	{8'd172,8'd193} : s = 365;
	{8'd172,8'd194} : s = 366;
	{8'd172,8'd195} : s = 367;
	{8'd172,8'd196} : s = 368;
	{8'd172,8'd197} : s = 369;
	{8'd172,8'd198} : s = 370;
	{8'd172,8'd199} : s = 371;
	{8'd172,8'd200} : s = 372;
	{8'd172,8'd201} : s = 373;
	{8'd172,8'd202} : s = 374;
	{8'd172,8'd203} : s = 375;
	{8'd172,8'd204} : s = 376;
	{8'd172,8'd205} : s = 377;
	{8'd172,8'd206} : s = 378;
	{8'd172,8'd207} : s = 379;
	{8'd172,8'd208} : s = 380;
	{8'd172,8'd209} : s = 381;
	{8'd172,8'd210} : s = 382;
	{8'd172,8'd211} : s = 383;
	{8'd172,8'd212} : s = 384;
	{8'd172,8'd213} : s = 385;
	{8'd172,8'd214} : s = 386;
	{8'd172,8'd215} : s = 387;
	{8'd172,8'd216} : s = 388;
	{8'd172,8'd217} : s = 389;
	{8'd172,8'd218} : s = 390;
	{8'd172,8'd219} : s = 391;
	{8'd172,8'd220} : s = 392;
	{8'd172,8'd221} : s = 393;
	{8'd172,8'd222} : s = 394;
	{8'd172,8'd223} : s = 395;
	{8'd172,8'd224} : s = 396;
	{8'd172,8'd225} : s = 397;
	{8'd172,8'd226} : s = 398;
	{8'd172,8'd227} : s = 399;
	{8'd172,8'd228} : s = 400;
	{8'd172,8'd229} : s = 401;
	{8'd172,8'd230} : s = 402;
	{8'd172,8'd231} : s = 403;
	{8'd172,8'd232} : s = 404;
	{8'd172,8'd233} : s = 405;
	{8'd172,8'd234} : s = 406;
	{8'd172,8'd235} : s = 407;
	{8'd172,8'd236} : s = 408;
	{8'd172,8'd237} : s = 409;
	{8'd172,8'd238} : s = 410;
	{8'd172,8'd239} : s = 411;
	{8'd172,8'd240} : s = 412;
	{8'd172,8'd241} : s = 413;
	{8'd172,8'd242} : s = 414;
	{8'd172,8'd243} : s = 415;
	{8'd172,8'd244} : s = 416;
	{8'd172,8'd245} : s = 417;
	{8'd172,8'd246} : s = 418;
	{8'd172,8'd247} : s = 419;
	{8'd172,8'd248} : s = 420;
	{8'd172,8'd249} : s = 421;
	{8'd172,8'd250} : s = 422;
	{8'd172,8'd251} : s = 423;
	{8'd172,8'd252} : s = 424;
	{8'd172,8'd253} : s = 425;
	{8'd172,8'd254} : s = 426;
	{8'd172,8'd255} : s = 427;
	{8'd173,8'd0} : s = 173;
	{8'd173,8'd1} : s = 174;
	{8'd173,8'd2} : s = 175;
	{8'd173,8'd3} : s = 176;
	{8'd173,8'd4} : s = 177;
	{8'd173,8'd5} : s = 178;
	{8'd173,8'd6} : s = 179;
	{8'd173,8'd7} : s = 180;
	{8'd173,8'd8} : s = 181;
	{8'd173,8'd9} : s = 182;
	{8'd173,8'd10} : s = 183;
	{8'd173,8'd11} : s = 184;
	{8'd173,8'd12} : s = 185;
	{8'd173,8'd13} : s = 186;
	{8'd173,8'd14} : s = 187;
	{8'd173,8'd15} : s = 188;
	{8'd173,8'd16} : s = 189;
	{8'd173,8'd17} : s = 190;
	{8'd173,8'd18} : s = 191;
	{8'd173,8'd19} : s = 192;
	{8'd173,8'd20} : s = 193;
	{8'd173,8'd21} : s = 194;
	{8'd173,8'd22} : s = 195;
	{8'd173,8'd23} : s = 196;
	{8'd173,8'd24} : s = 197;
	{8'd173,8'd25} : s = 198;
	{8'd173,8'd26} : s = 199;
	{8'd173,8'd27} : s = 200;
	{8'd173,8'd28} : s = 201;
	{8'd173,8'd29} : s = 202;
	{8'd173,8'd30} : s = 203;
	{8'd173,8'd31} : s = 204;
	{8'd173,8'd32} : s = 205;
	{8'd173,8'd33} : s = 206;
	{8'd173,8'd34} : s = 207;
	{8'd173,8'd35} : s = 208;
	{8'd173,8'd36} : s = 209;
	{8'd173,8'd37} : s = 210;
	{8'd173,8'd38} : s = 211;
	{8'd173,8'd39} : s = 212;
	{8'd173,8'd40} : s = 213;
	{8'd173,8'd41} : s = 214;
	{8'd173,8'd42} : s = 215;
	{8'd173,8'd43} : s = 216;
	{8'd173,8'd44} : s = 217;
	{8'd173,8'd45} : s = 218;
	{8'd173,8'd46} : s = 219;
	{8'd173,8'd47} : s = 220;
	{8'd173,8'd48} : s = 221;
	{8'd173,8'd49} : s = 222;
	{8'd173,8'd50} : s = 223;
	{8'd173,8'd51} : s = 224;
	{8'd173,8'd52} : s = 225;
	{8'd173,8'd53} : s = 226;
	{8'd173,8'd54} : s = 227;
	{8'd173,8'd55} : s = 228;
	{8'd173,8'd56} : s = 229;
	{8'd173,8'd57} : s = 230;
	{8'd173,8'd58} : s = 231;
	{8'd173,8'd59} : s = 232;
	{8'd173,8'd60} : s = 233;
	{8'd173,8'd61} : s = 234;
	{8'd173,8'd62} : s = 235;
	{8'd173,8'd63} : s = 236;
	{8'd173,8'd64} : s = 237;
	{8'd173,8'd65} : s = 238;
	{8'd173,8'd66} : s = 239;
	{8'd173,8'd67} : s = 240;
	{8'd173,8'd68} : s = 241;
	{8'd173,8'd69} : s = 242;
	{8'd173,8'd70} : s = 243;
	{8'd173,8'd71} : s = 244;
	{8'd173,8'd72} : s = 245;
	{8'd173,8'd73} : s = 246;
	{8'd173,8'd74} : s = 247;
	{8'd173,8'd75} : s = 248;
	{8'd173,8'd76} : s = 249;
	{8'd173,8'd77} : s = 250;
	{8'd173,8'd78} : s = 251;
	{8'd173,8'd79} : s = 252;
	{8'd173,8'd80} : s = 253;
	{8'd173,8'd81} : s = 254;
	{8'd173,8'd82} : s = 255;
	{8'd173,8'd83} : s = 256;
	{8'd173,8'd84} : s = 257;
	{8'd173,8'd85} : s = 258;
	{8'd173,8'd86} : s = 259;
	{8'd173,8'd87} : s = 260;
	{8'd173,8'd88} : s = 261;
	{8'd173,8'd89} : s = 262;
	{8'd173,8'd90} : s = 263;
	{8'd173,8'd91} : s = 264;
	{8'd173,8'd92} : s = 265;
	{8'd173,8'd93} : s = 266;
	{8'd173,8'd94} : s = 267;
	{8'd173,8'd95} : s = 268;
	{8'd173,8'd96} : s = 269;
	{8'd173,8'd97} : s = 270;
	{8'd173,8'd98} : s = 271;
	{8'd173,8'd99} : s = 272;
	{8'd173,8'd100} : s = 273;
	{8'd173,8'd101} : s = 274;
	{8'd173,8'd102} : s = 275;
	{8'd173,8'd103} : s = 276;
	{8'd173,8'd104} : s = 277;
	{8'd173,8'd105} : s = 278;
	{8'd173,8'd106} : s = 279;
	{8'd173,8'd107} : s = 280;
	{8'd173,8'd108} : s = 281;
	{8'd173,8'd109} : s = 282;
	{8'd173,8'd110} : s = 283;
	{8'd173,8'd111} : s = 284;
	{8'd173,8'd112} : s = 285;
	{8'd173,8'd113} : s = 286;
	{8'd173,8'd114} : s = 287;
	{8'd173,8'd115} : s = 288;
	{8'd173,8'd116} : s = 289;
	{8'd173,8'd117} : s = 290;
	{8'd173,8'd118} : s = 291;
	{8'd173,8'd119} : s = 292;
	{8'd173,8'd120} : s = 293;
	{8'd173,8'd121} : s = 294;
	{8'd173,8'd122} : s = 295;
	{8'd173,8'd123} : s = 296;
	{8'd173,8'd124} : s = 297;
	{8'd173,8'd125} : s = 298;
	{8'd173,8'd126} : s = 299;
	{8'd173,8'd127} : s = 300;
	{8'd173,8'd128} : s = 301;
	{8'd173,8'd129} : s = 302;
	{8'd173,8'd130} : s = 303;
	{8'd173,8'd131} : s = 304;
	{8'd173,8'd132} : s = 305;
	{8'd173,8'd133} : s = 306;
	{8'd173,8'd134} : s = 307;
	{8'd173,8'd135} : s = 308;
	{8'd173,8'd136} : s = 309;
	{8'd173,8'd137} : s = 310;
	{8'd173,8'd138} : s = 311;
	{8'd173,8'd139} : s = 312;
	{8'd173,8'd140} : s = 313;
	{8'd173,8'd141} : s = 314;
	{8'd173,8'd142} : s = 315;
	{8'd173,8'd143} : s = 316;
	{8'd173,8'd144} : s = 317;
	{8'd173,8'd145} : s = 318;
	{8'd173,8'd146} : s = 319;
	{8'd173,8'd147} : s = 320;
	{8'd173,8'd148} : s = 321;
	{8'd173,8'd149} : s = 322;
	{8'd173,8'd150} : s = 323;
	{8'd173,8'd151} : s = 324;
	{8'd173,8'd152} : s = 325;
	{8'd173,8'd153} : s = 326;
	{8'd173,8'd154} : s = 327;
	{8'd173,8'd155} : s = 328;
	{8'd173,8'd156} : s = 329;
	{8'd173,8'd157} : s = 330;
	{8'd173,8'd158} : s = 331;
	{8'd173,8'd159} : s = 332;
	{8'd173,8'd160} : s = 333;
	{8'd173,8'd161} : s = 334;
	{8'd173,8'd162} : s = 335;
	{8'd173,8'd163} : s = 336;
	{8'd173,8'd164} : s = 337;
	{8'd173,8'd165} : s = 338;
	{8'd173,8'd166} : s = 339;
	{8'd173,8'd167} : s = 340;
	{8'd173,8'd168} : s = 341;
	{8'd173,8'd169} : s = 342;
	{8'd173,8'd170} : s = 343;
	{8'd173,8'd171} : s = 344;
	{8'd173,8'd172} : s = 345;
	{8'd173,8'd173} : s = 346;
	{8'd173,8'd174} : s = 347;
	{8'd173,8'd175} : s = 348;
	{8'd173,8'd176} : s = 349;
	{8'd173,8'd177} : s = 350;
	{8'd173,8'd178} : s = 351;
	{8'd173,8'd179} : s = 352;
	{8'd173,8'd180} : s = 353;
	{8'd173,8'd181} : s = 354;
	{8'd173,8'd182} : s = 355;
	{8'd173,8'd183} : s = 356;
	{8'd173,8'd184} : s = 357;
	{8'd173,8'd185} : s = 358;
	{8'd173,8'd186} : s = 359;
	{8'd173,8'd187} : s = 360;
	{8'd173,8'd188} : s = 361;
	{8'd173,8'd189} : s = 362;
	{8'd173,8'd190} : s = 363;
	{8'd173,8'd191} : s = 364;
	{8'd173,8'd192} : s = 365;
	{8'd173,8'd193} : s = 366;
	{8'd173,8'd194} : s = 367;
	{8'd173,8'd195} : s = 368;
	{8'd173,8'd196} : s = 369;
	{8'd173,8'd197} : s = 370;
	{8'd173,8'd198} : s = 371;
	{8'd173,8'd199} : s = 372;
	{8'd173,8'd200} : s = 373;
	{8'd173,8'd201} : s = 374;
	{8'd173,8'd202} : s = 375;
	{8'd173,8'd203} : s = 376;
	{8'd173,8'd204} : s = 377;
	{8'd173,8'd205} : s = 378;
	{8'd173,8'd206} : s = 379;
	{8'd173,8'd207} : s = 380;
	{8'd173,8'd208} : s = 381;
	{8'd173,8'd209} : s = 382;
	{8'd173,8'd210} : s = 383;
	{8'd173,8'd211} : s = 384;
	{8'd173,8'd212} : s = 385;
	{8'd173,8'd213} : s = 386;
	{8'd173,8'd214} : s = 387;
	{8'd173,8'd215} : s = 388;
	{8'd173,8'd216} : s = 389;
	{8'd173,8'd217} : s = 390;
	{8'd173,8'd218} : s = 391;
	{8'd173,8'd219} : s = 392;
	{8'd173,8'd220} : s = 393;
	{8'd173,8'd221} : s = 394;
	{8'd173,8'd222} : s = 395;
	{8'd173,8'd223} : s = 396;
	{8'd173,8'd224} : s = 397;
	{8'd173,8'd225} : s = 398;
	{8'd173,8'd226} : s = 399;
	{8'd173,8'd227} : s = 400;
	{8'd173,8'd228} : s = 401;
	{8'd173,8'd229} : s = 402;
	{8'd173,8'd230} : s = 403;
	{8'd173,8'd231} : s = 404;
	{8'd173,8'd232} : s = 405;
	{8'd173,8'd233} : s = 406;
	{8'd173,8'd234} : s = 407;
	{8'd173,8'd235} : s = 408;
	{8'd173,8'd236} : s = 409;
	{8'd173,8'd237} : s = 410;
	{8'd173,8'd238} : s = 411;
	{8'd173,8'd239} : s = 412;
	{8'd173,8'd240} : s = 413;
	{8'd173,8'd241} : s = 414;
	{8'd173,8'd242} : s = 415;
	{8'd173,8'd243} : s = 416;
	{8'd173,8'd244} : s = 417;
	{8'd173,8'd245} : s = 418;
	{8'd173,8'd246} : s = 419;
	{8'd173,8'd247} : s = 420;
	{8'd173,8'd248} : s = 421;
	{8'd173,8'd249} : s = 422;
	{8'd173,8'd250} : s = 423;
	{8'd173,8'd251} : s = 424;
	{8'd173,8'd252} : s = 425;
	{8'd173,8'd253} : s = 426;
	{8'd173,8'd254} : s = 427;
	{8'd173,8'd255} : s = 428;
	{8'd174,8'd0} : s = 174;
	{8'd174,8'd1} : s = 175;
	{8'd174,8'd2} : s = 176;
	{8'd174,8'd3} : s = 177;
	{8'd174,8'd4} : s = 178;
	{8'd174,8'd5} : s = 179;
	{8'd174,8'd6} : s = 180;
	{8'd174,8'd7} : s = 181;
	{8'd174,8'd8} : s = 182;
	{8'd174,8'd9} : s = 183;
	{8'd174,8'd10} : s = 184;
	{8'd174,8'd11} : s = 185;
	{8'd174,8'd12} : s = 186;
	{8'd174,8'd13} : s = 187;
	{8'd174,8'd14} : s = 188;
	{8'd174,8'd15} : s = 189;
	{8'd174,8'd16} : s = 190;
	{8'd174,8'd17} : s = 191;
	{8'd174,8'd18} : s = 192;
	{8'd174,8'd19} : s = 193;
	{8'd174,8'd20} : s = 194;
	{8'd174,8'd21} : s = 195;
	{8'd174,8'd22} : s = 196;
	{8'd174,8'd23} : s = 197;
	{8'd174,8'd24} : s = 198;
	{8'd174,8'd25} : s = 199;
	{8'd174,8'd26} : s = 200;
	{8'd174,8'd27} : s = 201;
	{8'd174,8'd28} : s = 202;
	{8'd174,8'd29} : s = 203;
	{8'd174,8'd30} : s = 204;
	{8'd174,8'd31} : s = 205;
	{8'd174,8'd32} : s = 206;
	{8'd174,8'd33} : s = 207;
	{8'd174,8'd34} : s = 208;
	{8'd174,8'd35} : s = 209;
	{8'd174,8'd36} : s = 210;
	{8'd174,8'd37} : s = 211;
	{8'd174,8'd38} : s = 212;
	{8'd174,8'd39} : s = 213;
	{8'd174,8'd40} : s = 214;
	{8'd174,8'd41} : s = 215;
	{8'd174,8'd42} : s = 216;
	{8'd174,8'd43} : s = 217;
	{8'd174,8'd44} : s = 218;
	{8'd174,8'd45} : s = 219;
	{8'd174,8'd46} : s = 220;
	{8'd174,8'd47} : s = 221;
	{8'd174,8'd48} : s = 222;
	{8'd174,8'd49} : s = 223;
	{8'd174,8'd50} : s = 224;
	{8'd174,8'd51} : s = 225;
	{8'd174,8'd52} : s = 226;
	{8'd174,8'd53} : s = 227;
	{8'd174,8'd54} : s = 228;
	{8'd174,8'd55} : s = 229;
	{8'd174,8'd56} : s = 230;
	{8'd174,8'd57} : s = 231;
	{8'd174,8'd58} : s = 232;
	{8'd174,8'd59} : s = 233;
	{8'd174,8'd60} : s = 234;
	{8'd174,8'd61} : s = 235;
	{8'd174,8'd62} : s = 236;
	{8'd174,8'd63} : s = 237;
	{8'd174,8'd64} : s = 238;
	{8'd174,8'd65} : s = 239;
	{8'd174,8'd66} : s = 240;
	{8'd174,8'd67} : s = 241;
	{8'd174,8'd68} : s = 242;
	{8'd174,8'd69} : s = 243;
	{8'd174,8'd70} : s = 244;
	{8'd174,8'd71} : s = 245;
	{8'd174,8'd72} : s = 246;
	{8'd174,8'd73} : s = 247;
	{8'd174,8'd74} : s = 248;
	{8'd174,8'd75} : s = 249;
	{8'd174,8'd76} : s = 250;
	{8'd174,8'd77} : s = 251;
	{8'd174,8'd78} : s = 252;
	{8'd174,8'd79} : s = 253;
	{8'd174,8'd80} : s = 254;
	{8'd174,8'd81} : s = 255;
	{8'd174,8'd82} : s = 256;
	{8'd174,8'd83} : s = 257;
	{8'd174,8'd84} : s = 258;
	{8'd174,8'd85} : s = 259;
	{8'd174,8'd86} : s = 260;
	{8'd174,8'd87} : s = 261;
	{8'd174,8'd88} : s = 262;
	{8'd174,8'd89} : s = 263;
	{8'd174,8'd90} : s = 264;
	{8'd174,8'd91} : s = 265;
	{8'd174,8'd92} : s = 266;
	{8'd174,8'd93} : s = 267;
	{8'd174,8'd94} : s = 268;
	{8'd174,8'd95} : s = 269;
	{8'd174,8'd96} : s = 270;
	{8'd174,8'd97} : s = 271;
	{8'd174,8'd98} : s = 272;
	{8'd174,8'd99} : s = 273;
	{8'd174,8'd100} : s = 274;
	{8'd174,8'd101} : s = 275;
	{8'd174,8'd102} : s = 276;
	{8'd174,8'd103} : s = 277;
	{8'd174,8'd104} : s = 278;
	{8'd174,8'd105} : s = 279;
	{8'd174,8'd106} : s = 280;
	{8'd174,8'd107} : s = 281;
	{8'd174,8'd108} : s = 282;
	{8'd174,8'd109} : s = 283;
	{8'd174,8'd110} : s = 284;
	{8'd174,8'd111} : s = 285;
	{8'd174,8'd112} : s = 286;
	{8'd174,8'd113} : s = 287;
	{8'd174,8'd114} : s = 288;
	{8'd174,8'd115} : s = 289;
	{8'd174,8'd116} : s = 290;
	{8'd174,8'd117} : s = 291;
	{8'd174,8'd118} : s = 292;
	{8'd174,8'd119} : s = 293;
	{8'd174,8'd120} : s = 294;
	{8'd174,8'd121} : s = 295;
	{8'd174,8'd122} : s = 296;
	{8'd174,8'd123} : s = 297;
	{8'd174,8'd124} : s = 298;
	{8'd174,8'd125} : s = 299;
	{8'd174,8'd126} : s = 300;
	{8'd174,8'd127} : s = 301;
	{8'd174,8'd128} : s = 302;
	{8'd174,8'd129} : s = 303;
	{8'd174,8'd130} : s = 304;
	{8'd174,8'd131} : s = 305;
	{8'd174,8'd132} : s = 306;
	{8'd174,8'd133} : s = 307;
	{8'd174,8'd134} : s = 308;
	{8'd174,8'd135} : s = 309;
	{8'd174,8'd136} : s = 310;
	{8'd174,8'd137} : s = 311;
	{8'd174,8'd138} : s = 312;
	{8'd174,8'd139} : s = 313;
	{8'd174,8'd140} : s = 314;
	{8'd174,8'd141} : s = 315;
	{8'd174,8'd142} : s = 316;
	{8'd174,8'd143} : s = 317;
	{8'd174,8'd144} : s = 318;
	{8'd174,8'd145} : s = 319;
	{8'd174,8'd146} : s = 320;
	{8'd174,8'd147} : s = 321;
	{8'd174,8'd148} : s = 322;
	{8'd174,8'd149} : s = 323;
	{8'd174,8'd150} : s = 324;
	{8'd174,8'd151} : s = 325;
	{8'd174,8'd152} : s = 326;
	{8'd174,8'd153} : s = 327;
	{8'd174,8'd154} : s = 328;
	{8'd174,8'd155} : s = 329;
	{8'd174,8'd156} : s = 330;
	{8'd174,8'd157} : s = 331;
	{8'd174,8'd158} : s = 332;
	{8'd174,8'd159} : s = 333;
	{8'd174,8'd160} : s = 334;
	{8'd174,8'd161} : s = 335;
	{8'd174,8'd162} : s = 336;
	{8'd174,8'd163} : s = 337;
	{8'd174,8'd164} : s = 338;
	{8'd174,8'd165} : s = 339;
	{8'd174,8'd166} : s = 340;
	{8'd174,8'd167} : s = 341;
	{8'd174,8'd168} : s = 342;
	{8'd174,8'd169} : s = 343;
	{8'd174,8'd170} : s = 344;
	{8'd174,8'd171} : s = 345;
	{8'd174,8'd172} : s = 346;
	{8'd174,8'd173} : s = 347;
	{8'd174,8'd174} : s = 348;
	{8'd174,8'd175} : s = 349;
	{8'd174,8'd176} : s = 350;
	{8'd174,8'd177} : s = 351;
	{8'd174,8'd178} : s = 352;
	{8'd174,8'd179} : s = 353;
	{8'd174,8'd180} : s = 354;
	{8'd174,8'd181} : s = 355;
	{8'd174,8'd182} : s = 356;
	{8'd174,8'd183} : s = 357;
	{8'd174,8'd184} : s = 358;
	{8'd174,8'd185} : s = 359;
	{8'd174,8'd186} : s = 360;
	{8'd174,8'd187} : s = 361;
	{8'd174,8'd188} : s = 362;
	{8'd174,8'd189} : s = 363;
	{8'd174,8'd190} : s = 364;
	{8'd174,8'd191} : s = 365;
	{8'd174,8'd192} : s = 366;
	{8'd174,8'd193} : s = 367;
	{8'd174,8'd194} : s = 368;
	{8'd174,8'd195} : s = 369;
	{8'd174,8'd196} : s = 370;
	{8'd174,8'd197} : s = 371;
	{8'd174,8'd198} : s = 372;
	{8'd174,8'd199} : s = 373;
	{8'd174,8'd200} : s = 374;
	{8'd174,8'd201} : s = 375;
	{8'd174,8'd202} : s = 376;
	{8'd174,8'd203} : s = 377;
	{8'd174,8'd204} : s = 378;
	{8'd174,8'd205} : s = 379;
	{8'd174,8'd206} : s = 380;
	{8'd174,8'd207} : s = 381;
	{8'd174,8'd208} : s = 382;
	{8'd174,8'd209} : s = 383;
	{8'd174,8'd210} : s = 384;
	{8'd174,8'd211} : s = 385;
	{8'd174,8'd212} : s = 386;
	{8'd174,8'd213} : s = 387;
	{8'd174,8'd214} : s = 388;
	{8'd174,8'd215} : s = 389;
	{8'd174,8'd216} : s = 390;
	{8'd174,8'd217} : s = 391;
	{8'd174,8'd218} : s = 392;
	{8'd174,8'd219} : s = 393;
	{8'd174,8'd220} : s = 394;
	{8'd174,8'd221} : s = 395;
	{8'd174,8'd222} : s = 396;
	{8'd174,8'd223} : s = 397;
	{8'd174,8'd224} : s = 398;
	{8'd174,8'd225} : s = 399;
	{8'd174,8'd226} : s = 400;
	{8'd174,8'd227} : s = 401;
	{8'd174,8'd228} : s = 402;
	{8'd174,8'd229} : s = 403;
	{8'd174,8'd230} : s = 404;
	{8'd174,8'd231} : s = 405;
	{8'd174,8'd232} : s = 406;
	{8'd174,8'd233} : s = 407;
	{8'd174,8'd234} : s = 408;
	{8'd174,8'd235} : s = 409;
	{8'd174,8'd236} : s = 410;
	{8'd174,8'd237} : s = 411;
	{8'd174,8'd238} : s = 412;
	{8'd174,8'd239} : s = 413;
	{8'd174,8'd240} : s = 414;
	{8'd174,8'd241} : s = 415;
	{8'd174,8'd242} : s = 416;
	{8'd174,8'd243} : s = 417;
	{8'd174,8'd244} : s = 418;
	{8'd174,8'd245} : s = 419;
	{8'd174,8'd246} : s = 420;
	{8'd174,8'd247} : s = 421;
	{8'd174,8'd248} : s = 422;
	{8'd174,8'd249} : s = 423;
	{8'd174,8'd250} : s = 424;
	{8'd174,8'd251} : s = 425;
	{8'd174,8'd252} : s = 426;
	{8'd174,8'd253} : s = 427;
	{8'd174,8'd254} : s = 428;
	{8'd174,8'd255} : s = 429;
	{8'd175,8'd0} : s = 175;
	{8'd175,8'd1} : s = 176;
	{8'd175,8'd2} : s = 177;
	{8'd175,8'd3} : s = 178;
	{8'd175,8'd4} : s = 179;
	{8'd175,8'd5} : s = 180;
	{8'd175,8'd6} : s = 181;
	{8'd175,8'd7} : s = 182;
	{8'd175,8'd8} : s = 183;
	{8'd175,8'd9} : s = 184;
	{8'd175,8'd10} : s = 185;
	{8'd175,8'd11} : s = 186;
	{8'd175,8'd12} : s = 187;
	{8'd175,8'd13} : s = 188;
	{8'd175,8'd14} : s = 189;
	{8'd175,8'd15} : s = 190;
	{8'd175,8'd16} : s = 191;
	{8'd175,8'd17} : s = 192;
	{8'd175,8'd18} : s = 193;
	{8'd175,8'd19} : s = 194;
	{8'd175,8'd20} : s = 195;
	{8'd175,8'd21} : s = 196;
	{8'd175,8'd22} : s = 197;
	{8'd175,8'd23} : s = 198;
	{8'd175,8'd24} : s = 199;
	{8'd175,8'd25} : s = 200;
	{8'd175,8'd26} : s = 201;
	{8'd175,8'd27} : s = 202;
	{8'd175,8'd28} : s = 203;
	{8'd175,8'd29} : s = 204;
	{8'd175,8'd30} : s = 205;
	{8'd175,8'd31} : s = 206;
	{8'd175,8'd32} : s = 207;
	{8'd175,8'd33} : s = 208;
	{8'd175,8'd34} : s = 209;
	{8'd175,8'd35} : s = 210;
	{8'd175,8'd36} : s = 211;
	{8'd175,8'd37} : s = 212;
	{8'd175,8'd38} : s = 213;
	{8'd175,8'd39} : s = 214;
	{8'd175,8'd40} : s = 215;
	{8'd175,8'd41} : s = 216;
	{8'd175,8'd42} : s = 217;
	{8'd175,8'd43} : s = 218;
	{8'd175,8'd44} : s = 219;
	{8'd175,8'd45} : s = 220;
	{8'd175,8'd46} : s = 221;
	{8'd175,8'd47} : s = 222;
	{8'd175,8'd48} : s = 223;
	{8'd175,8'd49} : s = 224;
	{8'd175,8'd50} : s = 225;
	{8'd175,8'd51} : s = 226;
	{8'd175,8'd52} : s = 227;
	{8'd175,8'd53} : s = 228;
	{8'd175,8'd54} : s = 229;
	{8'd175,8'd55} : s = 230;
	{8'd175,8'd56} : s = 231;
	{8'd175,8'd57} : s = 232;
	{8'd175,8'd58} : s = 233;
	{8'd175,8'd59} : s = 234;
	{8'd175,8'd60} : s = 235;
	{8'd175,8'd61} : s = 236;
	{8'd175,8'd62} : s = 237;
	{8'd175,8'd63} : s = 238;
	{8'd175,8'd64} : s = 239;
	{8'd175,8'd65} : s = 240;
	{8'd175,8'd66} : s = 241;
	{8'd175,8'd67} : s = 242;
	{8'd175,8'd68} : s = 243;
	{8'd175,8'd69} : s = 244;
	{8'd175,8'd70} : s = 245;
	{8'd175,8'd71} : s = 246;
	{8'd175,8'd72} : s = 247;
	{8'd175,8'd73} : s = 248;
	{8'd175,8'd74} : s = 249;
	{8'd175,8'd75} : s = 250;
	{8'd175,8'd76} : s = 251;
	{8'd175,8'd77} : s = 252;
	{8'd175,8'd78} : s = 253;
	{8'd175,8'd79} : s = 254;
	{8'd175,8'd80} : s = 255;
	{8'd175,8'd81} : s = 256;
	{8'd175,8'd82} : s = 257;
	{8'd175,8'd83} : s = 258;
	{8'd175,8'd84} : s = 259;
	{8'd175,8'd85} : s = 260;
	{8'd175,8'd86} : s = 261;
	{8'd175,8'd87} : s = 262;
	{8'd175,8'd88} : s = 263;
	{8'd175,8'd89} : s = 264;
	{8'd175,8'd90} : s = 265;
	{8'd175,8'd91} : s = 266;
	{8'd175,8'd92} : s = 267;
	{8'd175,8'd93} : s = 268;
	{8'd175,8'd94} : s = 269;
	{8'd175,8'd95} : s = 270;
	{8'd175,8'd96} : s = 271;
	{8'd175,8'd97} : s = 272;
	{8'd175,8'd98} : s = 273;
	{8'd175,8'd99} : s = 274;
	{8'd175,8'd100} : s = 275;
	{8'd175,8'd101} : s = 276;
	{8'd175,8'd102} : s = 277;
	{8'd175,8'd103} : s = 278;
	{8'd175,8'd104} : s = 279;
	{8'd175,8'd105} : s = 280;
	{8'd175,8'd106} : s = 281;
	{8'd175,8'd107} : s = 282;
	{8'd175,8'd108} : s = 283;
	{8'd175,8'd109} : s = 284;
	{8'd175,8'd110} : s = 285;
	{8'd175,8'd111} : s = 286;
	{8'd175,8'd112} : s = 287;
	{8'd175,8'd113} : s = 288;
	{8'd175,8'd114} : s = 289;
	{8'd175,8'd115} : s = 290;
	{8'd175,8'd116} : s = 291;
	{8'd175,8'd117} : s = 292;
	{8'd175,8'd118} : s = 293;
	{8'd175,8'd119} : s = 294;
	{8'd175,8'd120} : s = 295;
	{8'd175,8'd121} : s = 296;
	{8'd175,8'd122} : s = 297;
	{8'd175,8'd123} : s = 298;
	{8'd175,8'd124} : s = 299;
	{8'd175,8'd125} : s = 300;
	{8'd175,8'd126} : s = 301;
	{8'd175,8'd127} : s = 302;
	{8'd175,8'd128} : s = 303;
	{8'd175,8'd129} : s = 304;
	{8'd175,8'd130} : s = 305;
	{8'd175,8'd131} : s = 306;
	{8'd175,8'd132} : s = 307;
	{8'd175,8'd133} : s = 308;
	{8'd175,8'd134} : s = 309;
	{8'd175,8'd135} : s = 310;
	{8'd175,8'd136} : s = 311;
	{8'd175,8'd137} : s = 312;
	{8'd175,8'd138} : s = 313;
	{8'd175,8'd139} : s = 314;
	{8'd175,8'd140} : s = 315;
	{8'd175,8'd141} : s = 316;
	{8'd175,8'd142} : s = 317;
	{8'd175,8'd143} : s = 318;
	{8'd175,8'd144} : s = 319;
	{8'd175,8'd145} : s = 320;
	{8'd175,8'd146} : s = 321;
	{8'd175,8'd147} : s = 322;
	{8'd175,8'd148} : s = 323;
	{8'd175,8'd149} : s = 324;
	{8'd175,8'd150} : s = 325;
	{8'd175,8'd151} : s = 326;
	{8'd175,8'd152} : s = 327;
	{8'd175,8'd153} : s = 328;
	{8'd175,8'd154} : s = 329;
	{8'd175,8'd155} : s = 330;
	{8'd175,8'd156} : s = 331;
	{8'd175,8'd157} : s = 332;
	{8'd175,8'd158} : s = 333;
	{8'd175,8'd159} : s = 334;
	{8'd175,8'd160} : s = 335;
	{8'd175,8'd161} : s = 336;
	{8'd175,8'd162} : s = 337;
	{8'd175,8'd163} : s = 338;
	{8'd175,8'd164} : s = 339;
	{8'd175,8'd165} : s = 340;
	{8'd175,8'd166} : s = 341;
	{8'd175,8'd167} : s = 342;
	{8'd175,8'd168} : s = 343;
	{8'd175,8'd169} : s = 344;
	{8'd175,8'd170} : s = 345;
	{8'd175,8'd171} : s = 346;
	{8'd175,8'd172} : s = 347;
	{8'd175,8'd173} : s = 348;
	{8'd175,8'd174} : s = 349;
	{8'd175,8'd175} : s = 350;
	{8'd175,8'd176} : s = 351;
	{8'd175,8'd177} : s = 352;
	{8'd175,8'd178} : s = 353;
	{8'd175,8'd179} : s = 354;
	{8'd175,8'd180} : s = 355;
	{8'd175,8'd181} : s = 356;
	{8'd175,8'd182} : s = 357;
	{8'd175,8'd183} : s = 358;
	{8'd175,8'd184} : s = 359;
	{8'd175,8'd185} : s = 360;
	{8'd175,8'd186} : s = 361;
	{8'd175,8'd187} : s = 362;
	{8'd175,8'd188} : s = 363;
	{8'd175,8'd189} : s = 364;
	{8'd175,8'd190} : s = 365;
	{8'd175,8'd191} : s = 366;
	{8'd175,8'd192} : s = 367;
	{8'd175,8'd193} : s = 368;
	{8'd175,8'd194} : s = 369;
	{8'd175,8'd195} : s = 370;
	{8'd175,8'd196} : s = 371;
	{8'd175,8'd197} : s = 372;
	{8'd175,8'd198} : s = 373;
	{8'd175,8'd199} : s = 374;
	{8'd175,8'd200} : s = 375;
	{8'd175,8'd201} : s = 376;
	{8'd175,8'd202} : s = 377;
	{8'd175,8'd203} : s = 378;
	{8'd175,8'd204} : s = 379;
	{8'd175,8'd205} : s = 380;
	{8'd175,8'd206} : s = 381;
	{8'd175,8'd207} : s = 382;
	{8'd175,8'd208} : s = 383;
	{8'd175,8'd209} : s = 384;
	{8'd175,8'd210} : s = 385;
	{8'd175,8'd211} : s = 386;
	{8'd175,8'd212} : s = 387;
	{8'd175,8'd213} : s = 388;
	{8'd175,8'd214} : s = 389;
	{8'd175,8'd215} : s = 390;
	{8'd175,8'd216} : s = 391;
	{8'd175,8'd217} : s = 392;
	{8'd175,8'd218} : s = 393;
	{8'd175,8'd219} : s = 394;
	{8'd175,8'd220} : s = 395;
	{8'd175,8'd221} : s = 396;
	{8'd175,8'd222} : s = 397;
	{8'd175,8'd223} : s = 398;
	{8'd175,8'd224} : s = 399;
	{8'd175,8'd225} : s = 400;
	{8'd175,8'd226} : s = 401;
	{8'd175,8'd227} : s = 402;
	{8'd175,8'd228} : s = 403;
	{8'd175,8'd229} : s = 404;
	{8'd175,8'd230} : s = 405;
	{8'd175,8'd231} : s = 406;
	{8'd175,8'd232} : s = 407;
	{8'd175,8'd233} : s = 408;
	{8'd175,8'd234} : s = 409;
	{8'd175,8'd235} : s = 410;
	{8'd175,8'd236} : s = 411;
	{8'd175,8'd237} : s = 412;
	{8'd175,8'd238} : s = 413;
	{8'd175,8'd239} : s = 414;
	{8'd175,8'd240} : s = 415;
	{8'd175,8'd241} : s = 416;
	{8'd175,8'd242} : s = 417;
	{8'd175,8'd243} : s = 418;
	{8'd175,8'd244} : s = 419;
	{8'd175,8'd245} : s = 420;
	{8'd175,8'd246} : s = 421;
	{8'd175,8'd247} : s = 422;
	{8'd175,8'd248} : s = 423;
	{8'd175,8'd249} : s = 424;
	{8'd175,8'd250} : s = 425;
	{8'd175,8'd251} : s = 426;
	{8'd175,8'd252} : s = 427;
	{8'd175,8'd253} : s = 428;
	{8'd175,8'd254} : s = 429;
	{8'd175,8'd255} : s = 430;
	{8'd176,8'd0} : s = 176;
	{8'd176,8'd1} : s = 177;
	{8'd176,8'd2} : s = 178;
	{8'd176,8'd3} : s = 179;
	{8'd176,8'd4} : s = 180;
	{8'd176,8'd5} : s = 181;
	{8'd176,8'd6} : s = 182;
	{8'd176,8'd7} : s = 183;
	{8'd176,8'd8} : s = 184;
	{8'd176,8'd9} : s = 185;
	{8'd176,8'd10} : s = 186;
	{8'd176,8'd11} : s = 187;
	{8'd176,8'd12} : s = 188;
	{8'd176,8'd13} : s = 189;
	{8'd176,8'd14} : s = 190;
	{8'd176,8'd15} : s = 191;
	{8'd176,8'd16} : s = 192;
	{8'd176,8'd17} : s = 193;
	{8'd176,8'd18} : s = 194;
	{8'd176,8'd19} : s = 195;
	{8'd176,8'd20} : s = 196;
	{8'd176,8'd21} : s = 197;
	{8'd176,8'd22} : s = 198;
	{8'd176,8'd23} : s = 199;
	{8'd176,8'd24} : s = 200;
	{8'd176,8'd25} : s = 201;
	{8'd176,8'd26} : s = 202;
	{8'd176,8'd27} : s = 203;
	{8'd176,8'd28} : s = 204;
	{8'd176,8'd29} : s = 205;
	{8'd176,8'd30} : s = 206;
	{8'd176,8'd31} : s = 207;
	{8'd176,8'd32} : s = 208;
	{8'd176,8'd33} : s = 209;
	{8'd176,8'd34} : s = 210;
	{8'd176,8'd35} : s = 211;
	{8'd176,8'd36} : s = 212;
	{8'd176,8'd37} : s = 213;
	{8'd176,8'd38} : s = 214;
	{8'd176,8'd39} : s = 215;
	{8'd176,8'd40} : s = 216;
	{8'd176,8'd41} : s = 217;
	{8'd176,8'd42} : s = 218;
	{8'd176,8'd43} : s = 219;
	{8'd176,8'd44} : s = 220;
	{8'd176,8'd45} : s = 221;
	{8'd176,8'd46} : s = 222;
	{8'd176,8'd47} : s = 223;
	{8'd176,8'd48} : s = 224;
	{8'd176,8'd49} : s = 225;
	{8'd176,8'd50} : s = 226;
	{8'd176,8'd51} : s = 227;
	{8'd176,8'd52} : s = 228;
	{8'd176,8'd53} : s = 229;
	{8'd176,8'd54} : s = 230;
	{8'd176,8'd55} : s = 231;
	{8'd176,8'd56} : s = 232;
	{8'd176,8'd57} : s = 233;
	{8'd176,8'd58} : s = 234;
	{8'd176,8'd59} : s = 235;
	{8'd176,8'd60} : s = 236;
	{8'd176,8'd61} : s = 237;
	{8'd176,8'd62} : s = 238;
	{8'd176,8'd63} : s = 239;
	{8'd176,8'd64} : s = 240;
	{8'd176,8'd65} : s = 241;
	{8'd176,8'd66} : s = 242;
	{8'd176,8'd67} : s = 243;
	{8'd176,8'd68} : s = 244;
	{8'd176,8'd69} : s = 245;
	{8'd176,8'd70} : s = 246;
	{8'd176,8'd71} : s = 247;
	{8'd176,8'd72} : s = 248;
	{8'd176,8'd73} : s = 249;
	{8'd176,8'd74} : s = 250;
	{8'd176,8'd75} : s = 251;
	{8'd176,8'd76} : s = 252;
	{8'd176,8'd77} : s = 253;
	{8'd176,8'd78} : s = 254;
	{8'd176,8'd79} : s = 255;
	{8'd176,8'd80} : s = 256;
	{8'd176,8'd81} : s = 257;
	{8'd176,8'd82} : s = 258;
	{8'd176,8'd83} : s = 259;
	{8'd176,8'd84} : s = 260;
	{8'd176,8'd85} : s = 261;
	{8'd176,8'd86} : s = 262;
	{8'd176,8'd87} : s = 263;
	{8'd176,8'd88} : s = 264;
	{8'd176,8'd89} : s = 265;
	{8'd176,8'd90} : s = 266;
	{8'd176,8'd91} : s = 267;
	{8'd176,8'd92} : s = 268;
	{8'd176,8'd93} : s = 269;
	{8'd176,8'd94} : s = 270;
	{8'd176,8'd95} : s = 271;
	{8'd176,8'd96} : s = 272;
	{8'd176,8'd97} : s = 273;
	{8'd176,8'd98} : s = 274;
	{8'd176,8'd99} : s = 275;
	{8'd176,8'd100} : s = 276;
	{8'd176,8'd101} : s = 277;
	{8'd176,8'd102} : s = 278;
	{8'd176,8'd103} : s = 279;
	{8'd176,8'd104} : s = 280;
	{8'd176,8'd105} : s = 281;
	{8'd176,8'd106} : s = 282;
	{8'd176,8'd107} : s = 283;
	{8'd176,8'd108} : s = 284;
	{8'd176,8'd109} : s = 285;
	{8'd176,8'd110} : s = 286;
	{8'd176,8'd111} : s = 287;
	{8'd176,8'd112} : s = 288;
	{8'd176,8'd113} : s = 289;
	{8'd176,8'd114} : s = 290;
	{8'd176,8'd115} : s = 291;
	{8'd176,8'd116} : s = 292;
	{8'd176,8'd117} : s = 293;
	{8'd176,8'd118} : s = 294;
	{8'd176,8'd119} : s = 295;
	{8'd176,8'd120} : s = 296;
	{8'd176,8'd121} : s = 297;
	{8'd176,8'd122} : s = 298;
	{8'd176,8'd123} : s = 299;
	{8'd176,8'd124} : s = 300;
	{8'd176,8'd125} : s = 301;
	{8'd176,8'd126} : s = 302;
	{8'd176,8'd127} : s = 303;
	{8'd176,8'd128} : s = 304;
	{8'd176,8'd129} : s = 305;
	{8'd176,8'd130} : s = 306;
	{8'd176,8'd131} : s = 307;
	{8'd176,8'd132} : s = 308;
	{8'd176,8'd133} : s = 309;
	{8'd176,8'd134} : s = 310;
	{8'd176,8'd135} : s = 311;
	{8'd176,8'd136} : s = 312;
	{8'd176,8'd137} : s = 313;
	{8'd176,8'd138} : s = 314;
	{8'd176,8'd139} : s = 315;
	{8'd176,8'd140} : s = 316;
	{8'd176,8'd141} : s = 317;
	{8'd176,8'd142} : s = 318;
	{8'd176,8'd143} : s = 319;
	{8'd176,8'd144} : s = 320;
	{8'd176,8'd145} : s = 321;
	{8'd176,8'd146} : s = 322;
	{8'd176,8'd147} : s = 323;
	{8'd176,8'd148} : s = 324;
	{8'd176,8'd149} : s = 325;
	{8'd176,8'd150} : s = 326;
	{8'd176,8'd151} : s = 327;
	{8'd176,8'd152} : s = 328;
	{8'd176,8'd153} : s = 329;
	{8'd176,8'd154} : s = 330;
	{8'd176,8'd155} : s = 331;
	{8'd176,8'd156} : s = 332;
	{8'd176,8'd157} : s = 333;
	{8'd176,8'd158} : s = 334;
	{8'd176,8'd159} : s = 335;
	{8'd176,8'd160} : s = 336;
	{8'd176,8'd161} : s = 337;
	{8'd176,8'd162} : s = 338;
	{8'd176,8'd163} : s = 339;
	{8'd176,8'd164} : s = 340;
	{8'd176,8'd165} : s = 341;
	{8'd176,8'd166} : s = 342;
	{8'd176,8'd167} : s = 343;
	{8'd176,8'd168} : s = 344;
	{8'd176,8'd169} : s = 345;
	{8'd176,8'd170} : s = 346;
	{8'd176,8'd171} : s = 347;
	{8'd176,8'd172} : s = 348;
	{8'd176,8'd173} : s = 349;
	{8'd176,8'd174} : s = 350;
	{8'd176,8'd175} : s = 351;
	{8'd176,8'd176} : s = 352;
	{8'd176,8'd177} : s = 353;
	{8'd176,8'd178} : s = 354;
	{8'd176,8'd179} : s = 355;
	{8'd176,8'd180} : s = 356;
	{8'd176,8'd181} : s = 357;
	{8'd176,8'd182} : s = 358;
	{8'd176,8'd183} : s = 359;
	{8'd176,8'd184} : s = 360;
	{8'd176,8'd185} : s = 361;
	{8'd176,8'd186} : s = 362;
	{8'd176,8'd187} : s = 363;
	{8'd176,8'd188} : s = 364;
	{8'd176,8'd189} : s = 365;
	{8'd176,8'd190} : s = 366;
	{8'd176,8'd191} : s = 367;
	{8'd176,8'd192} : s = 368;
	{8'd176,8'd193} : s = 369;
	{8'd176,8'd194} : s = 370;
	{8'd176,8'd195} : s = 371;
	{8'd176,8'd196} : s = 372;
	{8'd176,8'd197} : s = 373;
	{8'd176,8'd198} : s = 374;
	{8'd176,8'd199} : s = 375;
	{8'd176,8'd200} : s = 376;
	{8'd176,8'd201} : s = 377;
	{8'd176,8'd202} : s = 378;
	{8'd176,8'd203} : s = 379;
	{8'd176,8'd204} : s = 380;
	{8'd176,8'd205} : s = 381;
	{8'd176,8'd206} : s = 382;
	{8'd176,8'd207} : s = 383;
	{8'd176,8'd208} : s = 384;
	{8'd176,8'd209} : s = 385;
	{8'd176,8'd210} : s = 386;
	{8'd176,8'd211} : s = 387;
	{8'd176,8'd212} : s = 388;
	{8'd176,8'd213} : s = 389;
	{8'd176,8'd214} : s = 390;
	{8'd176,8'd215} : s = 391;
	{8'd176,8'd216} : s = 392;
	{8'd176,8'd217} : s = 393;
	{8'd176,8'd218} : s = 394;
	{8'd176,8'd219} : s = 395;
	{8'd176,8'd220} : s = 396;
	{8'd176,8'd221} : s = 397;
	{8'd176,8'd222} : s = 398;
	{8'd176,8'd223} : s = 399;
	{8'd176,8'd224} : s = 400;
	{8'd176,8'd225} : s = 401;
	{8'd176,8'd226} : s = 402;
	{8'd176,8'd227} : s = 403;
	{8'd176,8'd228} : s = 404;
	{8'd176,8'd229} : s = 405;
	{8'd176,8'd230} : s = 406;
	{8'd176,8'd231} : s = 407;
	{8'd176,8'd232} : s = 408;
	{8'd176,8'd233} : s = 409;
	{8'd176,8'd234} : s = 410;
	{8'd176,8'd235} : s = 411;
	{8'd176,8'd236} : s = 412;
	{8'd176,8'd237} : s = 413;
	{8'd176,8'd238} : s = 414;
	{8'd176,8'd239} : s = 415;
	{8'd176,8'd240} : s = 416;
	{8'd176,8'd241} : s = 417;
	{8'd176,8'd242} : s = 418;
	{8'd176,8'd243} : s = 419;
	{8'd176,8'd244} : s = 420;
	{8'd176,8'd245} : s = 421;
	{8'd176,8'd246} : s = 422;
	{8'd176,8'd247} : s = 423;
	{8'd176,8'd248} : s = 424;
	{8'd176,8'd249} : s = 425;
	{8'd176,8'd250} : s = 426;
	{8'd176,8'd251} : s = 427;
	{8'd176,8'd252} : s = 428;
	{8'd176,8'd253} : s = 429;
	{8'd176,8'd254} : s = 430;
	{8'd176,8'd255} : s = 431;
	{8'd177,8'd0} : s = 177;
	{8'd177,8'd1} : s = 178;
	{8'd177,8'd2} : s = 179;
	{8'd177,8'd3} : s = 180;
	{8'd177,8'd4} : s = 181;
	{8'd177,8'd5} : s = 182;
	{8'd177,8'd6} : s = 183;
	{8'd177,8'd7} : s = 184;
	{8'd177,8'd8} : s = 185;
	{8'd177,8'd9} : s = 186;
	{8'd177,8'd10} : s = 187;
	{8'd177,8'd11} : s = 188;
	{8'd177,8'd12} : s = 189;
	{8'd177,8'd13} : s = 190;
	{8'd177,8'd14} : s = 191;
	{8'd177,8'd15} : s = 192;
	{8'd177,8'd16} : s = 193;
	{8'd177,8'd17} : s = 194;
	{8'd177,8'd18} : s = 195;
	{8'd177,8'd19} : s = 196;
	{8'd177,8'd20} : s = 197;
	{8'd177,8'd21} : s = 198;
	{8'd177,8'd22} : s = 199;
	{8'd177,8'd23} : s = 200;
	{8'd177,8'd24} : s = 201;
	{8'd177,8'd25} : s = 202;
	{8'd177,8'd26} : s = 203;
	{8'd177,8'd27} : s = 204;
	{8'd177,8'd28} : s = 205;
	{8'd177,8'd29} : s = 206;
	{8'd177,8'd30} : s = 207;
	{8'd177,8'd31} : s = 208;
	{8'd177,8'd32} : s = 209;
	{8'd177,8'd33} : s = 210;
	{8'd177,8'd34} : s = 211;
	{8'd177,8'd35} : s = 212;
	{8'd177,8'd36} : s = 213;
	{8'd177,8'd37} : s = 214;
	{8'd177,8'd38} : s = 215;
	{8'd177,8'd39} : s = 216;
	{8'd177,8'd40} : s = 217;
	{8'd177,8'd41} : s = 218;
	{8'd177,8'd42} : s = 219;
	{8'd177,8'd43} : s = 220;
	{8'd177,8'd44} : s = 221;
	{8'd177,8'd45} : s = 222;
	{8'd177,8'd46} : s = 223;
	{8'd177,8'd47} : s = 224;
	{8'd177,8'd48} : s = 225;
	{8'd177,8'd49} : s = 226;
	{8'd177,8'd50} : s = 227;
	{8'd177,8'd51} : s = 228;
	{8'd177,8'd52} : s = 229;
	{8'd177,8'd53} : s = 230;
	{8'd177,8'd54} : s = 231;
	{8'd177,8'd55} : s = 232;
	{8'd177,8'd56} : s = 233;
	{8'd177,8'd57} : s = 234;
	{8'd177,8'd58} : s = 235;
	{8'd177,8'd59} : s = 236;
	{8'd177,8'd60} : s = 237;
	{8'd177,8'd61} : s = 238;
	{8'd177,8'd62} : s = 239;
	{8'd177,8'd63} : s = 240;
	{8'd177,8'd64} : s = 241;
	{8'd177,8'd65} : s = 242;
	{8'd177,8'd66} : s = 243;
	{8'd177,8'd67} : s = 244;
	{8'd177,8'd68} : s = 245;
	{8'd177,8'd69} : s = 246;
	{8'd177,8'd70} : s = 247;
	{8'd177,8'd71} : s = 248;
	{8'd177,8'd72} : s = 249;
	{8'd177,8'd73} : s = 250;
	{8'd177,8'd74} : s = 251;
	{8'd177,8'd75} : s = 252;
	{8'd177,8'd76} : s = 253;
	{8'd177,8'd77} : s = 254;
	{8'd177,8'd78} : s = 255;
	{8'd177,8'd79} : s = 256;
	{8'd177,8'd80} : s = 257;
	{8'd177,8'd81} : s = 258;
	{8'd177,8'd82} : s = 259;
	{8'd177,8'd83} : s = 260;
	{8'd177,8'd84} : s = 261;
	{8'd177,8'd85} : s = 262;
	{8'd177,8'd86} : s = 263;
	{8'd177,8'd87} : s = 264;
	{8'd177,8'd88} : s = 265;
	{8'd177,8'd89} : s = 266;
	{8'd177,8'd90} : s = 267;
	{8'd177,8'd91} : s = 268;
	{8'd177,8'd92} : s = 269;
	{8'd177,8'd93} : s = 270;
	{8'd177,8'd94} : s = 271;
	{8'd177,8'd95} : s = 272;
	{8'd177,8'd96} : s = 273;
	{8'd177,8'd97} : s = 274;
	{8'd177,8'd98} : s = 275;
	{8'd177,8'd99} : s = 276;
	{8'd177,8'd100} : s = 277;
	{8'd177,8'd101} : s = 278;
	{8'd177,8'd102} : s = 279;
	{8'd177,8'd103} : s = 280;
	{8'd177,8'd104} : s = 281;
	{8'd177,8'd105} : s = 282;
	{8'd177,8'd106} : s = 283;
	{8'd177,8'd107} : s = 284;
	{8'd177,8'd108} : s = 285;
	{8'd177,8'd109} : s = 286;
	{8'd177,8'd110} : s = 287;
	{8'd177,8'd111} : s = 288;
	{8'd177,8'd112} : s = 289;
	{8'd177,8'd113} : s = 290;
	{8'd177,8'd114} : s = 291;
	{8'd177,8'd115} : s = 292;
	{8'd177,8'd116} : s = 293;
	{8'd177,8'd117} : s = 294;
	{8'd177,8'd118} : s = 295;
	{8'd177,8'd119} : s = 296;
	{8'd177,8'd120} : s = 297;
	{8'd177,8'd121} : s = 298;
	{8'd177,8'd122} : s = 299;
	{8'd177,8'd123} : s = 300;
	{8'd177,8'd124} : s = 301;
	{8'd177,8'd125} : s = 302;
	{8'd177,8'd126} : s = 303;
	{8'd177,8'd127} : s = 304;
	{8'd177,8'd128} : s = 305;
	{8'd177,8'd129} : s = 306;
	{8'd177,8'd130} : s = 307;
	{8'd177,8'd131} : s = 308;
	{8'd177,8'd132} : s = 309;
	{8'd177,8'd133} : s = 310;
	{8'd177,8'd134} : s = 311;
	{8'd177,8'd135} : s = 312;
	{8'd177,8'd136} : s = 313;
	{8'd177,8'd137} : s = 314;
	{8'd177,8'd138} : s = 315;
	{8'd177,8'd139} : s = 316;
	{8'd177,8'd140} : s = 317;
	{8'd177,8'd141} : s = 318;
	{8'd177,8'd142} : s = 319;
	{8'd177,8'd143} : s = 320;
	{8'd177,8'd144} : s = 321;
	{8'd177,8'd145} : s = 322;
	{8'd177,8'd146} : s = 323;
	{8'd177,8'd147} : s = 324;
	{8'd177,8'd148} : s = 325;
	{8'd177,8'd149} : s = 326;
	{8'd177,8'd150} : s = 327;
	{8'd177,8'd151} : s = 328;
	{8'd177,8'd152} : s = 329;
	{8'd177,8'd153} : s = 330;
	{8'd177,8'd154} : s = 331;
	{8'd177,8'd155} : s = 332;
	{8'd177,8'd156} : s = 333;
	{8'd177,8'd157} : s = 334;
	{8'd177,8'd158} : s = 335;
	{8'd177,8'd159} : s = 336;
	{8'd177,8'd160} : s = 337;
	{8'd177,8'd161} : s = 338;
	{8'd177,8'd162} : s = 339;
	{8'd177,8'd163} : s = 340;
	{8'd177,8'd164} : s = 341;
	{8'd177,8'd165} : s = 342;
	{8'd177,8'd166} : s = 343;
	{8'd177,8'd167} : s = 344;
	{8'd177,8'd168} : s = 345;
	{8'd177,8'd169} : s = 346;
	{8'd177,8'd170} : s = 347;
	{8'd177,8'd171} : s = 348;
	{8'd177,8'd172} : s = 349;
	{8'd177,8'd173} : s = 350;
	{8'd177,8'd174} : s = 351;
	{8'd177,8'd175} : s = 352;
	{8'd177,8'd176} : s = 353;
	{8'd177,8'd177} : s = 354;
	{8'd177,8'd178} : s = 355;
	{8'd177,8'd179} : s = 356;
	{8'd177,8'd180} : s = 357;
	{8'd177,8'd181} : s = 358;
	{8'd177,8'd182} : s = 359;
	{8'd177,8'd183} : s = 360;
	{8'd177,8'd184} : s = 361;
	{8'd177,8'd185} : s = 362;
	{8'd177,8'd186} : s = 363;
	{8'd177,8'd187} : s = 364;
	{8'd177,8'd188} : s = 365;
	{8'd177,8'd189} : s = 366;
	{8'd177,8'd190} : s = 367;
	{8'd177,8'd191} : s = 368;
	{8'd177,8'd192} : s = 369;
	{8'd177,8'd193} : s = 370;
	{8'd177,8'd194} : s = 371;
	{8'd177,8'd195} : s = 372;
	{8'd177,8'd196} : s = 373;
	{8'd177,8'd197} : s = 374;
	{8'd177,8'd198} : s = 375;
	{8'd177,8'd199} : s = 376;
	{8'd177,8'd200} : s = 377;
	{8'd177,8'd201} : s = 378;
	{8'd177,8'd202} : s = 379;
	{8'd177,8'd203} : s = 380;
	{8'd177,8'd204} : s = 381;
	{8'd177,8'd205} : s = 382;
	{8'd177,8'd206} : s = 383;
	{8'd177,8'd207} : s = 384;
	{8'd177,8'd208} : s = 385;
	{8'd177,8'd209} : s = 386;
	{8'd177,8'd210} : s = 387;
	{8'd177,8'd211} : s = 388;
	{8'd177,8'd212} : s = 389;
	{8'd177,8'd213} : s = 390;
	{8'd177,8'd214} : s = 391;
	{8'd177,8'd215} : s = 392;
	{8'd177,8'd216} : s = 393;
	{8'd177,8'd217} : s = 394;
	{8'd177,8'd218} : s = 395;
	{8'd177,8'd219} : s = 396;
	{8'd177,8'd220} : s = 397;
	{8'd177,8'd221} : s = 398;
	{8'd177,8'd222} : s = 399;
	{8'd177,8'd223} : s = 400;
	{8'd177,8'd224} : s = 401;
	{8'd177,8'd225} : s = 402;
	{8'd177,8'd226} : s = 403;
	{8'd177,8'd227} : s = 404;
	{8'd177,8'd228} : s = 405;
	{8'd177,8'd229} : s = 406;
	{8'd177,8'd230} : s = 407;
	{8'd177,8'd231} : s = 408;
	{8'd177,8'd232} : s = 409;
	{8'd177,8'd233} : s = 410;
	{8'd177,8'd234} : s = 411;
	{8'd177,8'd235} : s = 412;
	{8'd177,8'd236} : s = 413;
	{8'd177,8'd237} : s = 414;
	{8'd177,8'd238} : s = 415;
	{8'd177,8'd239} : s = 416;
	{8'd177,8'd240} : s = 417;
	{8'd177,8'd241} : s = 418;
	{8'd177,8'd242} : s = 419;
	{8'd177,8'd243} : s = 420;
	{8'd177,8'd244} : s = 421;
	{8'd177,8'd245} : s = 422;
	{8'd177,8'd246} : s = 423;
	{8'd177,8'd247} : s = 424;
	{8'd177,8'd248} : s = 425;
	{8'd177,8'd249} : s = 426;
	{8'd177,8'd250} : s = 427;
	{8'd177,8'd251} : s = 428;
	{8'd177,8'd252} : s = 429;
	{8'd177,8'd253} : s = 430;
	{8'd177,8'd254} : s = 431;
	{8'd177,8'd255} : s = 432;
	{8'd178,8'd0} : s = 178;
	{8'd178,8'd1} : s = 179;
	{8'd178,8'd2} : s = 180;
	{8'd178,8'd3} : s = 181;
	{8'd178,8'd4} : s = 182;
	{8'd178,8'd5} : s = 183;
	{8'd178,8'd6} : s = 184;
	{8'd178,8'd7} : s = 185;
	{8'd178,8'd8} : s = 186;
	{8'd178,8'd9} : s = 187;
	{8'd178,8'd10} : s = 188;
	{8'd178,8'd11} : s = 189;
	{8'd178,8'd12} : s = 190;
	{8'd178,8'd13} : s = 191;
	{8'd178,8'd14} : s = 192;
	{8'd178,8'd15} : s = 193;
	{8'd178,8'd16} : s = 194;
	{8'd178,8'd17} : s = 195;
	{8'd178,8'd18} : s = 196;
	{8'd178,8'd19} : s = 197;
	{8'd178,8'd20} : s = 198;
	{8'd178,8'd21} : s = 199;
	{8'd178,8'd22} : s = 200;
	{8'd178,8'd23} : s = 201;
	{8'd178,8'd24} : s = 202;
	{8'd178,8'd25} : s = 203;
	{8'd178,8'd26} : s = 204;
	{8'd178,8'd27} : s = 205;
	{8'd178,8'd28} : s = 206;
	{8'd178,8'd29} : s = 207;
	{8'd178,8'd30} : s = 208;
	{8'd178,8'd31} : s = 209;
	{8'd178,8'd32} : s = 210;
	{8'd178,8'd33} : s = 211;
	{8'd178,8'd34} : s = 212;
	{8'd178,8'd35} : s = 213;
	{8'd178,8'd36} : s = 214;
	{8'd178,8'd37} : s = 215;
	{8'd178,8'd38} : s = 216;
	{8'd178,8'd39} : s = 217;
	{8'd178,8'd40} : s = 218;
	{8'd178,8'd41} : s = 219;
	{8'd178,8'd42} : s = 220;
	{8'd178,8'd43} : s = 221;
	{8'd178,8'd44} : s = 222;
	{8'd178,8'd45} : s = 223;
	{8'd178,8'd46} : s = 224;
	{8'd178,8'd47} : s = 225;
	{8'd178,8'd48} : s = 226;
	{8'd178,8'd49} : s = 227;
	{8'd178,8'd50} : s = 228;
	{8'd178,8'd51} : s = 229;
	{8'd178,8'd52} : s = 230;
	{8'd178,8'd53} : s = 231;
	{8'd178,8'd54} : s = 232;
	{8'd178,8'd55} : s = 233;
	{8'd178,8'd56} : s = 234;
	{8'd178,8'd57} : s = 235;
	{8'd178,8'd58} : s = 236;
	{8'd178,8'd59} : s = 237;
	{8'd178,8'd60} : s = 238;
	{8'd178,8'd61} : s = 239;
	{8'd178,8'd62} : s = 240;
	{8'd178,8'd63} : s = 241;
	{8'd178,8'd64} : s = 242;
	{8'd178,8'd65} : s = 243;
	{8'd178,8'd66} : s = 244;
	{8'd178,8'd67} : s = 245;
	{8'd178,8'd68} : s = 246;
	{8'd178,8'd69} : s = 247;
	{8'd178,8'd70} : s = 248;
	{8'd178,8'd71} : s = 249;
	{8'd178,8'd72} : s = 250;
	{8'd178,8'd73} : s = 251;
	{8'd178,8'd74} : s = 252;
	{8'd178,8'd75} : s = 253;
	{8'd178,8'd76} : s = 254;
	{8'd178,8'd77} : s = 255;
	{8'd178,8'd78} : s = 256;
	{8'd178,8'd79} : s = 257;
	{8'd178,8'd80} : s = 258;
	{8'd178,8'd81} : s = 259;
	{8'd178,8'd82} : s = 260;
	{8'd178,8'd83} : s = 261;
	{8'd178,8'd84} : s = 262;
	{8'd178,8'd85} : s = 263;
	{8'd178,8'd86} : s = 264;
	{8'd178,8'd87} : s = 265;
	{8'd178,8'd88} : s = 266;
	{8'd178,8'd89} : s = 267;
	{8'd178,8'd90} : s = 268;
	{8'd178,8'd91} : s = 269;
	{8'd178,8'd92} : s = 270;
	{8'd178,8'd93} : s = 271;
	{8'd178,8'd94} : s = 272;
	{8'd178,8'd95} : s = 273;
	{8'd178,8'd96} : s = 274;
	{8'd178,8'd97} : s = 275;
	{8'd178,8'd98} : s = 276;
	{8'd178,8'd99} : s = 277;
	{8'd178,8'd100} : s = 278;
	{8'd178,8'd101} : s = 279;
	{8'd178,8'd102} : s = 280;
	{8'd178,8'd103} : s = 281;
	{8'd178,8'd104} : s = 282;
	{8'd178,8'd105} : s = 283;
	{8'd178,8'd106} : s = 284;
	{8'd178,8'd107} : s = 285;
	{8'd178,8'd108} : s = 286;
	{8'd178,8'd109} : s = 287;
	{8'd178,8'd110} : s = 288;
	{8'd178,8'd111} : s = 289;
	{8'd178,8'd112} : s = 290;
	{8'd178,8'd113} : s = 291;
	{8'd178,8'd114} : s = 292;
	{8'd178,8'd115} : s = 293;
	{8'd178,8'd116} : s = 294;
	{8'd178,8'd117} : s = 295;
	{8'd178,8'd118} : s = 296;
	{8'd178,8'd119} : s = 297;
	{8'd178,8'd120} : s = 298;
	{8'd178,8'd121} : s = 299;
	{8'd178,8'd122} : s = 300;
	{8'd178,8'd123} : s = 301;
	{8'd178,8'd124} : s = 302;
	{8'd178,8'd125} : s = 303;
	{8'd178,8'd126} : s = 304;
	{8'd178,8'd127} : s = 305;
	{8'd178,8'd128} : s = 306;
	{8'd178,8'd129} : s = 307;
	{8'd178,8'd130} : s = 308;
	{8'd178,8'd131} : s = 309;
	{8'd178,8'd132} : s = 310;
	{8'd178,8'd133} : s = 311;
	{8'd178,8'd134} : s = 312;
	{8'd178,8'd135} : s = 313;
	{8'd178,8'd136} : s = 314;
	{8'd178,8'd137} : s = 315;
	{8'd178,8'd138} : s = 316;
	{8'd178,8'd139} : s = 317;
	{8'd178,8'd140} : s = 318;
	{8'd178,8'd141} : s = 319;
	{8'd178,8'd142} : s = 320;
	{8'd178,8'd143} : s = 321;
	{8'd178,8'd144} : s = 322;
	{8'd178,8'd145} : s = 323;
	{8'd178,8'd146} : s = 324;
	{8'd178,8'd147} : s = 325;
	{8'd178,8'd148} : s = 326;
	{8'd178,8'd149} : s = 327;
	{8'd178,8'd150} : s = 328;
	{8'd178,8'd151} : s = 329;
	{8'd178,8'd152} : s = 330;
	{8'd178,8'd153} : s = 331;
	{8'd178,8'd154} : s = 332;
	{8'd178,8'd155} : s = 333;
	{8'd178,8'd156} : s = 334;
	{8'd178,8'd157} : s = 335;
	{8'd178,8'd158} : s = 336;
	{8'd178,8'd159} : s = 337;
	{8'd178,8'd160} : s = 338;
	{8'd178,8'd161} : s = 339;
	{8'd178,8'd162} : s = 340;
	{8'd178,8'd163} : s = 341;
	{8'd178,8'd164} : s = 342;
	{8'd178,8'd165} : s = 343;
	{8'd178,8'd166} : s = 344;
	{8'd178,8'd167} : s = 345;
	{8'd178,8'd168} : s = 346;
	{8'd178,8'd169} : s = 347;
	{8'd178,8'd170} : s = 348;
	{8'd178,8'd171} : s = 349;
	{8'd178,8'd172} : s = 350;
	{8'd178,8'd173} : s = 351;
	{8'd178,8'd174} : s = 352;
	{8'd178,8'd175} : s = 353;
	{8'd178,8'd176} : s = 354;
	{8'd178,8'd177} : s = 355;
	{8'd178,8'd178} : s = 356;
	{8'd178,8'd179} : s = 357;
	{8'd178,8'd180} : s = 358;
	{8'd178,8'd181} : s = 359;
	{8'd178,8'd182} : s = 360;
	{8'd178,8'd183} : s = 361;
	{8'd178,8'd184} : s = 362;
	{8'd178,8'd185} : s = 363;
	{8'd178,8'd186} : s = 364;
	{8'd178,8'd187} : s = 365;
	{8'd178,8'd188} : s = 366;
	{8'd178,8'd189} : s = 367;
	{8'd178,8'd190} : s = 368;
	{8'd178,8'd191} : s = 369;
	{8'd178,8'd192} : s = 370;
	{8'd178,8'd193} : s = 371;
	{8'd178,8'd194} : s = 372;
	{8'd178,8'd195} : s = 373;
	{8'd178,8'd196} : s = 374;
	{8'd178,8'd197} : s = 375;
	{8'd178,8'd198} : s = 376;
	{8'd178,8'd199} : s = 377;
	{8'd178,8'd200} : s = 378;
	{8'd178,8'd201} : s = 379;
	{8'd178,8'd202} : s = 380;
	{8'd178,8'd203} : s = 381;
	{8'd178,8'd204} : s = 382;
	{8'd178,8'd205} : s = 383;
	{8'd178,8'd206} : s = 384;
	{8'd178,8'd207} : s = 385;
	{8'd178,8'd208} : s = 386;
	{8'd178,8'd209} : s = 387;
	{8'd178,8'd210} : s = 388;
	{8'd178,8'd211} : s = 389;
	{8'd178,8'd212} : s = 390;
	{8'd178,8'd213} : s = 391;
	{8'd178,8'd214} : s = 392;
	{8'd178,8'd215} : s = 393;
	{8'd178,8'd216} : s = 394;
	{8'd178,8'd217} : s = 395;
	{8'd178,8'd218} : s = 396;
	{8'd178,8'd219} : s = 397;
	{8'd178,8'd220} : s = 398;
	{8'd178,8'd221} : s = 399;
	{8'd178,8'd222} : s = 400;
	{8'd178,8'd223} : s = 401;
	{8'd178,8'd224} : s = 402;
	{8'd178,8'd225} : s = 403;
	{8'd178,8'd226} : s = 404;
	{8'd178,8'd227} : s = 405;
	{8'd178,8'd228} : s = 406;
	{8'd178,8'd229} : s = 407;
	{8'd178,8'd230} : s = 408;
	{8'd178,8'd231} : s = 409;
	{8'd178,8'd232} : s = 410;
	{8'd178,8'd233} : s = 411;
	{8'd178,8'd234} : s = 412;
	{8'd178,8'd235} : s = 413;
	{8'd178,8'd236} : s = 414;
	{8'd178,8'd237} : s = 415;
	{8'd178,8'd238} : s = 416;
	{8'd178,8'd239} : s = 417;
	{8'd178,8'd240} : s = 418;
	{8'd178,8'd241} : s = 419;
	{8'd178,8'd242} : s = 420;
	{8'd178,8'd243} : s = 421;
	{8'd178,8'd244} : s = 422;
	{8'd178,8'd245} : s = 423;
	{8'd178,8'd246} : s = 424;
	{8'd178,8'd247} : s = 425;
	{8'd178,8'd248} : s = 426;
	{8'd178,8'd249} : s = 427;
	{8'd178,8'd250} : s = 428;
	{8'd178,8'd251} : s = 429;
	{8'd178,8'd252} : s = 430;
	{8'd178,8'd253} : s = 431;
	{8'd178,8'd254} : s = 432;
	{8'd178,8'd255} : s = 433;
	{8'd179,8'd0} : s = 179;
	{8'd179,8'd1} : s = 180;
	{8'd179,8'd2} : s = 181;
	{8'd179,8'd3} : s = 182;
	{8'd179,8'd4} : s = 183;
	{8'd179,8'd5} : s = 184;
	{8'd179,8'd6} : s = 185;
	{8'd179,8'd7} : s = 186;
	{8'd179,8'd8} : s = 187;
	{8'd179,8'd9} : s = 188;
	{8'd179,8'd10} : s = 189;
	{8'd179,8'd11} : s = 190;
	{8'd179,8'd12} : s = 191;
	{8'd179,8'd13} : s = 192;
	{8'd179,8'd14} : s = 193;
	{8'd179,8'd15} : s = 194;
	{8'd179,8'd16} : s = 195;
	{8'd179,8'd17} : s = 196;
	{8'd179,8'd18} : s = 197;
	{8'd179,8'd19} : s = 198;
	{8'd179,8'd20} : s = 199;
	{8'd179,8'd21} : s = 200;
	{8'd179,8'd22} : s = 201;
	{8'd179,8'd23} : s = 202;
	{8'd179,8'd24} : s = 203;
	{8'd179,8'd25} : s = 204;
	{8'd179,8'd26} : s = 205;
	{8'd179,8'd27} : s = 206;
	{8'd179,8'd28} : s = 207;
	{8'd179,8'd29} : s = 208;
	{8'd179,8'd30} : s = 209;
	{8'd179,8'd31} : s = 210;
	{8'd179,8'd32} : s = 211;
	{8'd179,8'd33} : s = 212;
	{8'd179,8'd34} : s = 213;
	{8'd179,8'd35} : s = 214;
	{8'd179,8'd36} : s = 215;
	{8'd179,8'd37} : s = 216;
	{8'd179,8'd38} : s = 217;
	{8'd179,8'd39} : s = 218;
	{8'd179,8'd40} : s = 219;
	{8'd179,8'd41} : s = 220;
	{8'd179,8'd42} : s = 221;
	{8'd179,8'd43} : s = 222;
	{8'd179,8'd44} : s = 223;
	{8'd179,8'd45} : s = 224;
	{8'd179,8'd46} : s = 225;
	{8'd179,8'd47} : s = 226;
	{8'd179,8'd48} : s = 227;
	{8'd179,8'd49} : s = 228;
	{8'd179,8'd50} : s = 229;
	{8'd179,8'd51} : s = 230;
	{8'd179,8'd52} : s = 231;
	{8'd179,8'd53} : s = 232;
	{8'd179,8'd54} : s = 233;
	{8'd179,8'd55} : s = 234;
	{8'd179,8'd56} : s = 235;
	{8'd179,8'd57} : s = 236;
	{8'd179,8'd58} : s = 237;
	{8'd179,8'd59} : s = 238;
	{8'd179,8'd60} : s = 239;
	{8'd179,8'd61} : s = 240;
	{8'd179,8'd62} : s = 241;
	{8'd179,8'd63} : s = 242;
	{8'd179,8'd64} : s = 243;
	{8'd179,8'd65} : s = 244;
	{8'd179,8'd66} : s = 245;
	{8'd179,8'd67} : s = 246;
	{8'd179,8'd68} : s = 247;
	{8'd179,8'd69} : s = 248;
	{8'd179,8'd70} : s = 249;
	{8'd179,8'd71} : s = 250;
	{8'd179,8'd72} : s = 251;
	{8'd179,8'd73} : s = 252;
	{8'd179,8'd74} : s = 253;
	{8'd179,8'd75} : s = 254;
	{8'd179,8'd76} : s = 255;
	{8'd179,8'd77} : s = 256;
	{8'd179,8'd78} : s = 257;
	{8'd179,8'd79} : s = 258;
	{8'd179,8'd80} : s = 259;
	{8'd179,8'd81} : s = 260;
	{8'd179,8'd82} : s = 261;
	{8'd179,8'd83} : s = 262;
	{8'd179,8'd84} : s = 263;
	{8'd179,8'd85} : s = 264;
	{8'd179,8'd86} : s = 265;
	{8'd179,8'd87} : s = 266;
	{8'd179,8'd88} : s = 267;
	{8'd179,8'd89} : s = 268;
	{8'd179,8'd90} : s = 269;
	{8'd179,8'd91} : s = 270;
	{8'd179,8'd92} : s = 271;
	{8'd179,8'd93} : s = 272;
	{8'd179,8'd94} : s = 273;
	{8'd179,8'd95} : s = 274;
	{8'd179,8'd96} : s = 275;
	{8'd179,8'd97} : s = 276;
	{8'd179,8'd98} : s = 277;
	{8'd179,8'd99} : s = 278;
	{8'd179,8'd100} : s = 279;
	{8'd179,8'd101} : s = 280;
	{8'd179,8'd102} : s = 281;
	{8'd179,8'd103} : s = 282;
	{8'd179,8'd104} : s = 283;
	{8'd179,8'd105} : s = 284;
	{8'd179,8'd106} : s = 285;
	{8'd179,8'd107} : s = 286;
	{8'd179,8'd108} : s = 287;
	{8'd179,8'd109} : s = 288;
	{8'd179,8'd110} : s = 289;
	{8'd179,8'd111} : s = 290;
	{8'd179,8'd112} : s = 291;
	{8'd179,8'd113} : s = 292;
	{8'd179,8'd114} : s = 293;
	{8'd179,8'd115} : s = 294;
	{8'd179,8'd116} : s = 295;
	{8'd179,8'd117} : s = 296;
	{8'd179,8'd118} : s = 297;
	{8'd179,8'd119} : s = 298;
	{8'd179,8'd120} : s = 299;
	{8'd179,8'd121} : s = 300;
	{8'd179,8'd122} : s = 301;
	{8'd179,8'd123} : s = 302;
	{8'd179,8'd124} : s = 303;
	{8'd179,8'd125} : s = 304;
	{8'd179,8'd126} : s = 305;
	{8'd179,8'd127} : s = 306;
	{8'd179,8'd128} : s = 307;
	{8'd179,8'd129} : s = 308;
	{8'd179,8'd130} : s = 309;
	{8'd179,8'd131} : s = 310;
	{8'd179,8'd132} : s = 311;
	{8'd179,8'd133} : s = 312;
	{8'd179,8'd134} : s = 313;
	{8'd179,8'd135} : s = 314;
	{8'd179,8'd136} : s = 315;
	{8'd179,8'd137} : s = 316;
	{8'd179,8'd138} : s = 317;
	{8'd179,8'd139} : s = 318;
	{8'd179,8'd140} : s = 319;
	{8'd179,8'd141} : s = 320;
	{8'd179,8'd142} : s = 321;
	{8'd179,8'd143} : s = 322;
	{8'd179,8'd144} : s = 323;
	{8'd179,8'd145} : s = 324;
	{8'd179,8'd146} : s = 325;
	{8'd179,8'd147} : s = 326;
	{8'd179,8'd148} : s = 327;
	{8'd179,8'd149} : s = 328;
	{8'd179,8'd150} : s = 329;
	{8'd179,8'd151} : s = 330;
	{8'd179,8'd152} : s = 331;
	{8'd179,8'd153} : s = 332;
	{8'd179,8'd154} : s = 333;
	{8'd179,8'd155} : s = 334;
	{8'd179,8'd156} : s = 335;
	{8'd179,8'd157} : s = 336;
	{8'd179,8'd158} : s = 337;
	{8'd179,8'd159} : s = 338;
	{8'd179,8'd160} : s = 339;
	{8'd179,8'd161} : s = 340;
	{8'd179,8'd162} : s = 341;
	{8'd179,8'd163} : s = 342;
	{8'd179,8'd164} : s = 343;
	{8'd179,8'd165} : s = 344;
	{8'd179,8'd166} : s = 345;
	{8'd179,8'd167} : s = 346;
	{8'd179,8'd168} : s = 347;
	{8'd179,8'd169} : s = 348;
	{8'd179,8'd170} : s = 349;
	{8'd179,8'd171} : s = 350;
	{8'd179,8'd172} : s = 351;
	{8'd179,8'd173} : s = 352;
	{8'd179,8'd174} : s = 353;
	{8'd179,8'd175} : s = 354;
	{8'd179,8'd176} : s = 355;
	{8'd179,8'd177} : s = 356;
	{8'd179,8'd178} : s = 357;
	{8'd179,8'd179} : s = 358;
	{8'd179,8'd180} : s = 359;
	{8'd179,8'd181} : s = 360;
	{8'd179,8'd182} : s = 361;
	{8'd179,8'd183} : s = 362;
	{8'd179,8'd184} : s = 363;
	{8'd179,8'd185} : s = 364;
	{8'd179,8'd186} : s = 365;
	{8'd179,8'd187} : s = 366;
	{8'd179,8'd188} : s = 367;
	{8'd179,8'd189} : s = 368;
	{8'd179,8'd190} : s = 369;
	{8'd179,8'd191} : s = 370;
	{8'd179,8'd192} : s = 371;
	{8'd179,8'd193} : s = 372;
	{8'd179,8'd194} : s = 373;
	{8'd179,8'd195} : s = 374;
	{8'd179,8'd196} : s = 375;
	{8'd179,8'd197} : s = 376;
	{8'd179,8'd198} : s = 377;
	{8'd179,8'd199} : s = 378;
	{8'd179,8'd200} : s = 379;
	{8'd179,8'd201} : s = 380;
	{8'd179,8'd202} : s = 381;
	{8'd179,8'd203} : s = 382;
	{8'd179,8'd204} : s = 383;
	{8'd179,8'd205} : s = 384;
	{8'd179,8'd206} : s = 385;
	{8'd179,8'd207} : s = 386;
	{8'd179,8'd208} : s = 387;
	{8'd179,8'd209} : s = 388;
	{8'd179,8'd210} : s = 389;
	{8'd179,8'd211} : s = 390;
	{8'd179,8'd212} : s = 391;
	{8'd179,8'd213} : s = 392;
	{8'd179,8'd214} : s = 393;
	{8'd179,8'd215} : s = 394;
	{8'd179,8'd216} : s = 395;
	{8'd179,8'd217} : s = 396;
	{8'd179,8'd218} : s = 397;
	{8'd179,8'd219} : s = 398;
	{8'd179,8'd220} : s = 399;
	{8'd179,8'd221} : s = 400;
	{8'd179,8'd222} : s = 401;
	{8'd179,8'd223} : s = 402;
	{8'd179,8'd224} : s = 403;
	{8'd179,8'd225} : s = 404;
	{8'd179,8'd226} : s = 405;
	{8'd179,8'd227} : s = 406;
	{8'd179,8'd228} : s = 407;
	{8'd179,8'd229} : s = 408;
	{8'd179,8'd230} : s = 409;
	{8'd179,8'd231} : s = 410;
	{8'd179,8'd232} : s = 411;
	{8'd179,8'd233} : s = 412;
	{8'd179,8'd234} : s = 413;
	{8'd179,8'd235} : s = 414;
	{8'd179,8'd236} : s = 415;
	{8'd179,8'd237} : s = 416;
	{8'd179,8'd238} : s = 417;
	{8'd179,8'd239} : s = 418;
	{8'd179,8'd240} : s = 419;
	{8'd179,8'd241} : s = 420;
	{8'd179,8'd242} : s = 421;
	{8'd179,8'd243} : s = 422;
	{8'd179,8'd244} : s = 423;
	{8'd179,8'd245} : s = 424;
	{8'd179,8'd246} : s = 425;
	{8'd179,8'd247} : s = 426;
	{8'd179,8'd248} : s = 427;
	{8'd179,8'd249} : s = 428;
	{8'd179,8'd250} : s = 429;
	{8'd179,8'd251} : s = 430;
	{8'd179,8'd252} : s = 431;
	{8'd179,8'd253} : s = 432;
	{8'd179,8'd254} : s = 433;
	{8'd179,8'd255} : s = 434;
	{8'd180,8'd0} : s = 180;
	{8'd180,8'd1} : s = 181;
	{8'd180,8'd2} : s = 182;
	{8'd180,8'd3} : s = 183;
	{8'd180,8'd4} : s = 184;
	{8'd180,8'd5} : s = 185;
	{8'd180,8'd6} : s = 186;
	{8'd180,8'd7} : s = 187;
	{8'd180,8'd8} : s = 188;
	{8'd180,8'd9} : s = 189;
	{8'd180,8'd10} : s = 190;
	{8'd180,8'd11} : s = 191;
	{8'd180,8'd12} : s = 192;
	{8'd180,8'd13} : s = 193;
	{8'd180,8'd14} : s = 194;
	{8'd180,8'd15} : s = 195;
	{8'd180,8'd16} : s = 196;
	{8'd180,8'd17} : s = 197;
	{8'd180,8'd18} : s = 198;
	{8'd180,8'd19} : s = 199;
	{8'd180,8'd20} : s = 200;
	{8'd180,8'd21} : s = 201;
	{8'd180,8'd22} : s = 202;
	{8'd180,8'd23} : s = 203;
	{8'd180,8'd24} : s = 204;
	{8'd180,8'd25} : s = 205;
	{8'd180,8'd26} : s = 206;
	{8'd180,8'd27} : s = 207;
	{8'd180,8'd28} : s = 208;
	{8'd180,8'd29} : s = 209;
	{8'd180,8'd30} : s = 210;
	{8'd180,8'd31} : s = 211;
	{8'd180,8'd32} : s = 212;
	{8'd180,8'd33} : s = 213;
	{8'd180,8'd34} : s = 214;
	{8'd180,8'd35} : s = 215;
	{8'd180,8'd36} : s = 216;
	{8'd180,8'd37} : s = 217;
	{8'd180,8'd38} : s = 218;
	{8'd180,8'd39} : s = 219;
	{8'd180,8'd40} : s = 220;
	{8'd180,8'd41} : s = 221;
	{8'd180,8'd42} : s = 222;
	{8'd180,8'd43} : s = 223;
	{8'd180,8'd44} : s = 224;
	{8'd180,8'd45} : s = 225;
	{8'd180,8'd46} : s = 226;
	{8'd180,8'd47} : s = 227;
	{8'd180,8'd48} : s = 228;
	{8'd180,8'd49} : s = 229;
	{8'd180,8'd50} : s = 230;
	{8'd180,8'd51} : s = 231;
	{8'd180,8'd52} : s = 232;
	{8'd180,8'd53} : s = 233;
	{8'd180,8'd54} : s = 234;
	{8'd180,8'd55} : s = 235;
	{8'd180,8'd56} : s = 236;
	{8'd180,8'd57} : s = 237;
	{8'd180,8'd58} : s = 238;
	{8'd180,8'd59} : s = 239;
	{8'd180,8'd60} : s = 240;
	{8'd180,8'd61} : s = 241;
	{8'd180,8'd62} : s = 242;
	{8'd180,8'd63} : s = 243;
	{8'd180,8'd64} : s = 244;
	{8'd180,8'd65} : s = 245;
	{8'd180,8'd66} : s = 246;
	{8'd180,8'd67} : s = 247;
	{8'd180,8'd68} : s = 248;
	{8'd180,8'd69} : s = 249;
	{8'd180,8'd70} : s = 250;
	{8'd180,8'd71} : s = 251;
	{8'd180,8'd72} : s = 252;
	{8'd180,8'd73} : s = 253;
	{8'd180,8'd74} : s = 254;
	{8'd180,8'd75} : s = 255;
	{8'd180,8'd76} : s = 256;
	{8'd180,8'd77} : s = 257;
	{8'd180,8'd78} : s = 258;
	{8'd180,8'd79} : s = 259;
	{8'd180,8'd80} : s = 260;
	{8'd180,8'd81} : s = 261;
	{8'd180,8'd82} : s = 262;
	{8'd180,8'd83} : s = 263;
	{8'd180,8'd84} : s = 264;
	{8'd180,8'd85} : s = 265;
	{8'd180,8'd86} : s = 266;
	{8'd180,8'd87} : s = 267;
	{8'd180,8'd88} : s = 268;
	{8'd180,8'd89} : s = 269;
	{8'd180,8'd90} : s = 270;
	{8'd180,8'd91} : s = 271;
	{8'd180,8'd92} : s = 272;
	{8'd180,8'd93} : s = 273;
	{8'd180,8'd94} : s = 274;
	{8'd180,8'd95} : s = 275;
	{8'd180,8'd96} : s = 276;
	{8'd180,8'd97} : s = 277;
	{8'd180,8'd98} : s = 278;
	{8'd180,8'd99} : s = 279;
	{8'd180,8'd100} : s = 280;
	{8'd180,8'd101} : s = 281;
	{8'd180,8'd102} : s = 282;
	{8'd180,8'd103} : s = 283;
	{8'd180,8'd104} : s = 284;
	{8'd180,8'd105} : s = 285;
	{8'd180,8'd106} : s = 286;
	{8'd180,8'd107} : s = 287;
	{8'd180,8'd108} : s = 288;
	{8'd180,8'd109} : s = 289;
	{8'd180,8'd110} : s = 290;
	{8'd180,8'd111} : s = 291;
	{8'd180,8'd112} : s = 292;
	{8'd180,8'd113} : s = 293;
	{8'd180,8'd114} : s = 294;
	{8'd180,8'd115} : s = 295;
	{8'd180,8'd116} : s = 296;
	{8'd180,8'd117} : s = 297;
	{8'd180,8'd118} : s = 298;
	{8'd180,8'd119} : s = 299;
	{8'd180,8'd120} : s = 300;
	{8'd180,8'd121} : s = 301;
	{8'd180,8'd122} : s = 302;
	{8'd180,8'd123} : s = 303;
	{8'd180,8'd124} : s = 304;
	{8'd180,8'd125} : s = 305;
	{8'd180,8'd126} : s = 306;
	{8'd180,8'd127} : s = 307;
	{8'd180,8'd128} : s = 308;
	{8'd180,8'd129} : s = 309;
	{8'd180,8'd130} : s = 310;
	{8'd180,8'd131} : s = 311;
	{8'd180,8'd132} : s = 312;
	{8'd180,8'd133} : s = 313;
	{8'd180,8'd134} : s = 314;
	{8'd180,8'd135} : s = 315;
	{8'd180,8'd136} : s = 316;
	{8'd180,8'd137} : s = 317;
	{8'd180,8'd138} : s = 318;
	{8'd180,8'd139} : s = 319;
	{8'd180,8'd140} : s = 320;
	{8'd180,8'd141} : s = 321;
	{8'd180,8'd142} : s = 322;
	{8'd180,8'd143} : s = 323;
	{8'd180,8'd144} : s = 324;
	{8'd180,8'd145} : s = 325;
	{8'd180,8'd146} : s = 326;
	{8'd180,8'd147} : s = 327;
	{8'd180,8'd148} : s = 328;
	{8'd180,8'd149} : s = 329;
	{8'd180,8'd150} : s = 330;
	{8'd180,8'd151} : s = 331;
	{8'd180,8'd152} : s = 332;
	{8'd180,8'd153} : s = 333;
	{8'd180,8'd154} : s = 334;
	{8'd180,8'd155} : s = 335;
	{8'd180,8'd156} : s = 336;
	{8'd180,8'd157} : s = 337;
	{8'd180,8'd158} : s = 338;
	{8'd180,8'd159} : s = 339;
	{8'd180,8'd160} : s = 340;
	{8'd180,8'd161} : s = 341;
	{8'd180,8'd162} : s = 342;
	{8'd180,8'd163} : s = 343;
	{8'd180,8'd164} : s = 344;
	{8'd180,8'd165} : s = 345;
	{8'd180,8'd166} : s = 346;
	{8'd180,8'd167} : s = 347;
	{8'd180,8'd168} : s = 348;
	{8'd180,8'd169} : s = 349;
	{8'd180,8'd170} : s = 350;
	{8'd180,8'd171} : s = 351;
	{8'd180,8'd172} : s = 352;
	{8'd180,8'd173} : s = 353;
	{8'd180,8'd174} : s = 354;
	{8'd180,8'd175} : s = 355;
	{8'd180,8'd176} : s = 356;
	{8'd180,8'd177} : s = 357;
	{8'd180,8'd178} : s = 358;
	{8'd180,8'd179} : s = 359;
	{8'd180,8'd180} : s = 360;
	{8'd180,8'd181} : s = 361;
	{8'd180,8'd182} : s = 362;
	{8'd180,8'd183} : s = 363;
	{8'd180,8'd184} : s = 364;
	{8'd180,8'd185} : s = 365;
	{8'd180,8'd186} : s = 366;
	{8'd180,8'd187} : s = 367;
	{8'd180,8'd188} : s = 368;
	{8'd180,8'd189} : s = 369;
	{8'd180,8'd190} : s = 370;
	{8'd180,8'd191} : s = 371;
	{8'd180,8'd192} : s = 372;
	{8'd180,8'd193} : s = 373;
	{8'd180,8'd194} : s = 374;
	{8'd180,8'd195} : s = 375;
	{8'd180,8'd196} : s = 376;
	{8'd180,8'd197} : s = 377;
	{8'd180,8'd198} : s = 378;
	{8'd180,8'd199} : s = 379;
	{8'd180,8'd200} : s = 380;
	{8'd180,8'd201} : s = 381;
	{8'd180,8'd202} : s = 382;
	{8'd180,8'd203} : s = 383;
	{8'd180,8'd204} : s = 384;
	{8'd180,8'd205} : s = 385;
	{8'd180,8'd206} : s = 386;
	{8'd180,8'd207} : s = 387;
	{8'd180,8'd208} : s = 388;
	{8'd180,8'd209} : s = 389;
	{8'd180,8'd210} : s = 390;
	{8'd180,8'd211} : s = 391;
	{8'd180,8'd212} : s = 392;
	{8'd180,8'd213} : s = 393;
	{8'd180,8'd214} : s = 394;
	{8'd180,8'd215} : s = 395;
	{8'd180,8'd216} : s = 396;
	{8'd180,8'd217} : s = 397;
	{8'd180,8'd218} : s = 398;
	{8'd180,8'd219} : s = 399;
	{8'd180,8'd220} : s = 400;
	{8'd180,8'd221} : s = 401;
	{8'd180,8'd222} : s = 402;
	{8'd180,8'd223} : s = 403;
	{8'd180,8'd224} : s = 404;
	{8'd180,8'd225} : s = 405;
	{8'd180,8'd226} : s = 406;
	{8'd180,8'd227} : s = 407;
	{8'd180,8'd228} : s = 408;
	{8'd180,8'd229} : s = 409;
	{8'd180,8'd230} : s = 410;
	{8'd180,8'd231} : s = 411;
	{8'd180,8'd232} : s = 412;
	{8'd180,8'd233} : s = 413;
	{8'd180,8'd234} : s = 414;
	{8'd180,8'd235} : s = 415;
	{8'd180,8'd236} : s = 416;
	{8'd180,8'd237} : s = 417;
	{8'd180,8'd238} : s = 418;
	{8'd180,8'd239} : s = 419;
	{8'd180,8'd240} : s = 420;
	{8'd180,8'd241} : s = 421;
	{8'd180,8'd242} : s = 422;
	{8'd180,8'd243} : s = 423;
	{8'd180,8'd244} : s = 424;
	{8'd180,8'd245} : s = 425;
	{8'd180,8'd246} : s = 426;
	{8'd180,8'd247} : s = 427;
	{8'd180,8'd248} : s = 428;
	{8'd180,8'd249} : s = 429;
	{8'd180,8'd250} : s = 430;
	{8'd180,8'd251} : s = 431;
	{8'd180,8'd252} : s = 432;
	{8'd180,8'd253} : s = 433;
	{8'd180,8'd254} : s = 434;
	{8'd180,8'd255} : s = 435;
	{8'd181,8'd0} : s = 181;
	{8'd181,8'd1} : s = 182;
	{8'd181,8'd2} : s = 183;
	{8'd181,8'd3} : s = 184;
	{8'd181,8'd4} : s = 185;
	{8'd181,8'd5} : s = 186;
	{8'd181,8'd6} : s = 187;
	{8'd181,8'd7} : s = 188;
	{8'd181,8'd8} : s = 189;
	{8'd181,8'd9} : s = 190;
	{8'd181,8'd10} : s = 191;
	{8'd181,8'd11} : s = 192;
	{8'd181,8'd12} : s = 193;
	{8'd181,8'd13} : s = 194;
	{8'd181,8'd14} : s = 195;
	{8'd181,8'd15} : s = 196;
	{8'd181,8'd16} : s = 197;
	{8'd181,8'd17} : s = 198;
	{8'd181,8'd18} : s = 199;
	{8'd181,8'd19} : s = 200;
	{8'd181,8'd20} : s = 201;
	{8'd181,8'd21} : s = 202;
	{8'd181,8'd22} : s = 203;
	{8'd181,8'd23} : s = 204;
	{8'd181,8'd24} : s = 205;
	{8'd181,8'd25} : s = 206;
	{8'd181,8'd26} : s = 207;
	{8'd181,8'd27} : s = 208;
	{8'd181,8'd28} : s = 209;
	{8'd181,8'd29} : s = 210;
	{8'd181,8'd30} : s = 211;
	{8'd181,8'd31} : s = 212;
	{8'd181,8'd32} : s = 213;
	{8'd181,8'd33} : s = 214;
	{8'd181,8'd34} : s = 215;
	{8'd181,8'd35} : s = 216;
	{8'd181,8'd36} : s = 217;
	{8'd181,8'd37} : s = 218;
	{8'd181,8'd38} : s = 219;
	{8'd181,8'd39} : s = 220;
	{8'd181,8'd40} : s = 221;
	{8'd181,8'd41} : s = 222;
	{8'd181,8'd42} : s = 223;
	{8'd181,8'd43} : s = 224;
	{8'd181,8'd44} : s = 225;
	{8'd181,8'd45} : s = 226;
	{8'd181,8'd46} : s = 227;
	{8'd181,8'd47} : s = 228;
	{8'd181,8'd48} : s = 229;
	{8'd181,8'd49} : s = 230;
	{8'd181,8'd50} : s = 231;
	{8'd181,8'd51} : s = 232;
	{8'd181,8'd52} : s = 233;
	{8'd181,8'd53} : s = 234;
	{8'd181,8'd54} : s = 235;
	{8'd181,8'd55} : s = 236;
	{8'd181,8'd56} : s = 237;
	{8'd181,8'd57} : s = 238;
	{8'd181,8'd58} : s = 239;
	{8'd181,8'd59} : s = 240;
	{8'd181,8'd60} : s = 241;
	{8'd181,8'd61} : s = 242;
	{8'd181,8'd62} : s = 243;
	{8'd181,8'd63} : s = 244;
	{8'd181,8'd64} : s = 245;
	{8'd181,8'd65} : s = 246;
	{8'd181,8'd66} : s = 247;
	{8'd181,8'd67} : s = 248;
	{8'd181,8'd68} : s = 249;
	{8'd181,8'd69} : s = 250;
	{8'd181,8'd70} : s = 251;
	{8'd181,8'd71} : s = 252;
	{8'd181,8'd72} : s = 253;
	{8'd181,8'd73} : s = 254;
	{8'd181,8'd74} : s = 255;
	{8'd181,8'd75} : s = 256;
	{8'd181,8'd76} : s = 257;
	{8'd181,8'd77} : s = 258;
	{8'd181,8'd78} : s = 259;
	{8'd181,8'd79} : s = 260;
	{8'd181,8'd80} : s = 261;
	{8'd181,8'd81} : s = 262;
	{8'd181,8'd82} : s = 263;
	{8'd181,8'd83} : s = 264;
	{8'd181,8'd84} : s = 265;
	{8'd181,8'd85} : s = 266;
	{8'd181,8'd86} : s = 267;
	{8'd181,8'd87} : s = 268;
	{8'd181,8'd88} : s = 269;
	{8'd181,8'd89} : s = 270;
	{8'd181,8'd90} : s = 271;
	{8'd181,8'd91} : s = 272;
	{8'd181,8'd92} : s = 273;
	{8'd181,8'd93} : s = 274;
	{8'd181,8'd94} : s = 275;
	{8'd181,8'd95} : s = 276;
	{8'd181,8'd96} : s = 277;
	{8'd181,8'd97} : s = 278;
	{8'd181,8'd98} : s = 279;
	{8'd181,8'd99} : s = 280;
	{8'd181,8'd100} : s = 281;
	{8'd181,8'd101} : s = 282;
	{8'd181,8'd102} : s = 283;
	{8'd181,8'd103} : s = 284;
	{8'd181,8'd104} : s = 285;
	{8'd181,8'd105} : s = 286;
	{8'd181,8'd106} : s = 287;
	{8'd181,8'd107} : s = 288;
	{8'd181,8'd108} : s = 289;
	{8'd181,8'd109} : s = 290;
	{8'd181,8'd110} : s = 291;
	{8'd181,8'd111} : s = 292;
	{8'd181,8'd112} : s = 293;
	{8'd181,8'd113} : s = 294;
	{8'd181,8'd114} : s = 295;
	{8'd181,8'd115} : s = 296;
	{8'd181,8'd116} : s = 297;
	{8'd181,8'd117} : s = 298;
	{8'd181,8'd118} : s = 299;
	{8'd181,8'd119} : s = 300;
	{8'd181,8'd120} : s = 301;
	{8'd181,8'd121} : s = 302;
	{8'd181,8'd122} : s = 303;
	{8'd181,8'd123} : s = 304;
	{8'd181,8'd124} : s = 305;
	{8'd181,8'd125} : s = 306;
	{8'd181,8'd126} : s = 307;
	{8'd181,8'd127} : s = 308;
	{8'd181,8'd128} : s = 309;
	{8'd181,8'd129} : s = 310;
	{8'd181,8'd130} : s = 311;
	{8'd181,8'd131} : s = 312;
	{8'd181,8'd132} : s = 313;
	{8'd181,8'd133} : s = 314;
	{8'd181,8'd134} : s = 315;
	{8'd181,8'd135} : s = 316;
	{8'd181,8'd136} : s = 317;
	{8'd181,8'd137} : s = 318;
	{8'd181,8'd138} : s = 319;
	{8'd181,8'd139} : s = 320;
	{8'd181,8'd140} : s = 321;
	{8'd181,8'd141} : s = 322;
	{8'd181,8'd142} : s = 323;
	{8'd181,8'd143} : s = 324;
	{8'd181,8'd144} : s = 325;
	{8'd181,8'd145} : s = 326;
	{8'd181,8'd146} : s = 327;
	{8'd181,8'd147} : s = 328;
	{8'd181,8'd148} : s = 329;
	{8'd181,8'd149} : s = 330;
	{8'd181,8'd150} : s = 331;
	{8'd181,8'd151} : s = 332;
	{8'd181,8'd152} : s = 333;
	{8'd181,8'd153} : s = 334;
	{8'd181,8'd154} : s = 335;
	{8'd181,8'd155} : s = 336;
	{8'd181,8'd156} : s = 337;
	{8'd181,8'd157} : s = 338;
	{8'd181,8'd158} : s = 339;
	{8'd181,8'd159} : s = 340;
	{8'd181,8'd160} : s = 341;
	{8'd181,8'd161} : s = 342;
	{8'd181,8'd162} : s = 343;
	{8'd181,8'd163} : s = 344;
	{8'd181,8'd164} : s = 345;
	{8'd181,8'd165} : s = 346;
	{8'd181,8'd166} : s = 347;
	{8'd181,8'd167} : s = 348;
	{8'd181,8'd168} : s = 349;
	{8'd181,8'd169} : s = 350;
	{8'd181,8'd170} : s = 351;
	{8'd181,8'd171} : s = 352;
	{8'd181,8'd172} : s = 353;
	{8'd181,8'd173} : s = 354;
	{8'd181,8'd174} : s = 355;
	{8'd181,8'd175} : s = 356;
	{8'd181,8'd176} : s = 357;
	{8'd181,8'd177} : s = 358;
	{8'd181,8'd178} : s = 359;
	{8'd181,8'd179} : s = 360;
	{8'd181,8'd180} : s = 361;
	{8'd181,8'd181} : s = 362;
	{8'd181,8'd182} : s = 363;
	{8'd181,8'd183} : s = 364;
	{8'd181,8'd184} : s = 365;
	{8'd181,8'd185} : s = 366;
	{8'd181,8'd186} : s = 367;
	{8'd181,8'd187} : s = 368;
	{8'd181,8'd188} : s = 369;
	{8'd181,8'd189} : s = 370;
	{8'd181,8'd190} : s = 371;
	{8'd181,8'd191} : s = 372;
	{8'd181,8'd192} : s = 373;
	{8'd181,8'd193} : s = 374;
	{8'd181,8'd194} : s = 375;
	{8'd181,8'd195} : s = 376;
	{8'd181,8'd196} : s = 377;
	{8'd181,8'd197} : s = 378;
	{8'd181,8'd198} : s = 379;
	{8'd181,8'd199} : s = 380;
	{8'd181,8'd200} : s = 381;
	{8'd181,8'd201} : s = 382;
	{8'd181,8'd202} : s = 383;
	{8'd181,8'd203} : s = 384;
	{8'd181,8'd204} : s = 385;
	{8'd181,8'd205} : s = 386;
	{8'd181,8'd206} : s = 387;
	{8'd181,8'd207} : s = 388;
	{8'd181,8'd208} : s = 389;
	{8'd181,8'd209} : s = 390;
	{8'd181,8'd210} : s = 391;
	{8'd181,8'd211} : s = 392;
	{8'd181,8'd212} : s = 393;
	{8'd181,8'd213} : s = 394;
	{8'd181,8'd214} : s = 395;
	{8'd181,8'd215} : s = 396;
	{8'd181,8'd216} : s = 397;
	{8'd181,8'd217} : s = 398;
	{8'd181,8'd218} : s = 399;
	{8'd181,8'd219} : s = 400;
	{8'd181,8'd220} : s = 401;
	{8'd181,8'd221} : s = 402;
	{8'd181,8'd222} : s = 403;
	{8'd181,8'd223} : s = 404;
	{8'd181,8'd224} : s = 405;
	{8'd181,8'd225} : s = 406;
	{8'd181,8'd226} : s = 407;
	{8'd181,8'd227} : s = 408;
	{8'd181,8'd228} : s = 409;
	{8'd181,8'd229} : s = 410;
	{8'd181,8'd230} : s = 411;
	{8'd181,8'd231} : s = 412;
	{8'd181,8'd232} : s = 413;
	{8'd181,8'd233} : s = 414;
	{8'd181,8'd234} : s = 415;
	{8'd181,8'd235} : s = 416;
	{8'd181,8'd236} : s = 417;
	{8'd181,8'd237} : s = 418;
	{8'd181,8'd238} : s = 419;
	{8'd181,8'd239} : s = 420;
	{8'd181,8'd240} : s = 421;
	{8'd181,8'd241} : s = 422;
	{8'd181,8'd242} : s = 423;
	{8'd181,8'd243} : s = 424;
	{8'd181,8'd244} : s = 425;
	{8'd181,8'd245} : s = 426;
	{8'd181,8'd246} : s = 427;
	{8'd181,8'd247} : s = 428;
	{8'd181,8'd248} : s = 429;
	{8'd181,8'd249} : s = 430;
	{8'd181,8'd250} : s = 431;
	{8'd181,8'd251} : s = 432;
	{8'd181,8'd252} : s = 433;
	{8'd181,8'd253} : s = 434;
	{8'd181,8'd254} : s = 435;
	{8'd181,8'd255} : s = 436;
	{8'd182,8'd0} : s = 182;
	{8'd182,8'd1} : s = 183;
	{8'd182,8'd2} : s = 184;
	{8'd182,8'd3} : s = 185;
	{8'd182,8'd4} : s = 186;
	{8'd182,8'd5} : s = 187;
	{8'd182,8'd6} : s = 188;
	{8'd182,8'd7} : s = 189;
	{8'd182,8'd8} : s = 190;
	{8'd182,8'd9} : s = 191;
	{8'd182,8'd10} : s = 192;
	{8'd182,8'd11} : s = 193;
	{8'd182,8'd12} : s = 194;
	{8'd182,8'd13} : s = 195;
	{8'd182,8'd14} : s = 196;
	{8'd182,8'd15} : s = 197;
	{8'd182,8'd16} : s = 198;
	{8'd182,8'd17} : s = 199;
	{8'd182,8'd18} : s = 200;
	{8'd182,8'd19} : s = 201;
	{8'd182,8'd20} : s = 202;
	{8'd182,8'd21} : s = 203;
	{8'd182,8'd22} : s = 204;
	{8'd182,8'd23} : s = 205;
	{8'd182,8'd24} : s = 206;
	{8'd182,8'd25} : s = 207;
	{8'd182,8'd26} : s = 208;
	{8'd182,8'd27} : s = 209;
	{8'd182,8'd28} : s = 210;
	{8'd182,8'd29} : s = 211;
	{8'd182,8'd30} : s = 212;
	{8'd182,8'd31} : s = 213;
	{8'd182,8'd32} : s = 214;
	{8'd182,8'd33} : s = 215;
	{8'd182,8'd34} : s = 216;
	{8'd182,8'd35} : s = 217;
	{8'd182,8'd36} : s = 218;
	{8'd182,8'd37} : s = 219;
	{8'd182,8'd38} : s = 220;
	{8'd182,8'd39} : s = 221;
	{8'd182,8'd40} : s = 222;
	{8'd182,8'd41} : s = 223;
	{8'd182,8'd42} : s = 224;
	{8'd182,8'd43} : s = 225;
	{8'd182,8'd44} : s = 226;
	{8'd182,8'd45} : s = 227;
	{8'd182,8'd46} : s = 228;
	{8'd182,8'd47} : s = 229;
	{8'd182,8'd48} : s = 230;
	{8'd182,8'd49} : s = 231;
	{8'd182,8'd50} : s = 232;
	{8'd182,8'd51} : s = 233;
	{8'd182,8'd52} : s = 234;
	{8'd182,8'd53} : s = 235;
	{8'd182,8'd54} : s = 236;
	{8'd182,8'd55} : s = 237;
	{8'd182,8'd56} : s = 238;
	{8'd182,8'd57} : s = 239;
	{8'd182,8'd58} : s = 240;
	{8'd182,8'd59} : s = 241;
	{8'd182,8'd60} : s = 242;
	{8'd182,8'd61} : s = 243;
	{8'd182,8'd62} : s = 244;
	{8'd182,8'd63} : s = 245;
	{8'd182,8'd64} : s = 246;
	{8'd182,8'd65} : s = 247;
	{8'd182,8'd66} : s = 248;
	{8'd182,8'd67} : s = 249;
	{8'd182,8'd68} : s = 250;
	{8'd182,8'd69} : s = 251;
	{8'd182,8'd70} : s = 252;
	{8'd182,8'd71} : s = 253;
	{8'd182,8'd72} : s = 254;
	{8'd182,8'd73} : s = 255;
	{8'd182,8'd74} : s = 256;
	{8'd182,8'd75} : s = 257;
	{8'd182,8'd76} : s = 258;
	{8'd182,8'd77} : s = 259;
	{8'd182,8'd78} : s = 260;
	{8'd182,8'd79} : s = 261;
	{8'd182,8'd80} : s = 262;
	{8'd182,8'd81} : s = 263;
	{8'd182,8'd82} : s = 264;
	{8'd182,8'd83} : s = 265;
	{8'd182,8'd84} : s = 266;
	{8'd182,8'd85} : s = 267;
	{8'd182,8'd86} : s = 268;
	{8'd182,8'd87} : s = 269;
	{8'd182,8'd88} : s = 270;
	{8'd182,8'd89} : s = 271;
	{8'd182,8'd90} : s = 272;
	{8'd182,8'd91} : s = 273;
	{8'd182,8'd92} : s = 274;
	{8'd182,8'd93} : s = 275;
	{8'd182,8'd94} : s = 276;
	{8'd182,8'd95} : s = 277;
	{8'd182,8'd96} : s = 278;
	{8'd182,8'd97} : s = 279;
	{8'd182,8'd98} : s = 280;
	{8'd182,8'd99} : s = 281;
	{8'd182,8'd100} : s = 282;
	{8'd182,8'd101} : s = 283;
	{8'd182,8'd102} : s = 284;
	{8'd182,8'd103} : s = 285;
	{8'd182,8'd104} : s = 286;
	{8'd182,8'd105} : s = 287;
	{8'd182,8'd106} : s = 288;
	{8'd182,8'd107} : s = 289;
	{8'd182,8'd108} : s = 290;
	{8'd182,8'd109} : s = 291;
	{8'd182,8'd110} : s = 292;
	{8'd182,8'd111} : s = 293;
	{8'd182,8'd112} : s = 294;
	{8'd182,8'd113} : s = 295;
	{8'd182,8'd114} : s = 296;
	{8'd182,8'd115} : s = 297;
	{8'd182,8'd116} : s = 298;
	{8'd182,8'd117} : s = 299;
	{8'd182,8'd118} : s = 300;
	{8'd182,8'd119} : s = 301;
	{8'd182,8'd120} : s = 302;
	{8'd182,8'd121} : s = 303;
	{8'd182,8'd122} : s = 304;
	{8'd182,8'd123} : s = 305;
	{8'd182,8'd124} : s = 306;
	{8'd182,8'd125} : s = 307;
	{8'd182,8'd126} : s = 308;
	{8'd182,8'd127} : s = 309;
	{8'd182,8'd128} : s = 310;
	{8'd182,8'd129} : s = 311;
	{8'd182,8'd130} : s = 312;
	{8'd182,8'd131} : s = 313;
	{8'd182,8'd132} : s = 314;
	{8'd182,8'd133} : s = 315;
	{8'd182,8'd134} : s = 316;
	{8'd182,8'd135} : s = 317;
	{8'd182,8'd136} : s = 318;
	{8'd182,8'd137} : s = 319;
	{8'd182,8'd138} : s = 320;
	{8'd182,8'd139} : s = 321;
	{8'd182,8'd140} : s = 322;
	{8'd182,8'd141} : s = 323;
	{8'd182,8'd142} : s = 324;
	{8'd182,8'd143} : s = 325;
	{8'd182,8'd144} : s = 326;
	{8'd182,8'd145} : s = 327;
	{8'd182,8'd146} : s = 328;
	{8'd182,8'd147} : s = 329;
	{8'd182,8'd148} : s = 330;
	{8'd182,8'd149} : s = 331;
	{8'd182,8'd150} : s = 332;
	{8'd182,8'd151} : s = 333;
	{8'd182,8'd152} : s = 334;
	{8'd182,8'd153} : s = 335;
	{8'd182,8'd154} : s = 336;
	{8'd182,8'd155} : s = 337;
	{8'd182,8'd156} : s = 338;
	{8'd182,8'd157} : s = 339;
	{8'd182,8'd158} : s = 340;
	{8'd182,8'd159} : s = 341;
	{8'd182,8'd160} : s = 342;
	{8'd182,8'd161} : s = 343;
	{8'd182,8'd162} : s = 344;
	{8'd182,8'd163} : s = 345;
	{8'd182,8'd164} : s = 346;
	{8'd182,8'd165} : s = 347;
	{8'd182,8'd166} : s = 348;
	{8'd182,8'd167} : s = 349;
	{8'd182,8'd168} : s = 350;
	{8'd182,8'd169} : s = 351;
	{8'd182,8'd170} : s = 352;
	{8'd182,8'd171} : s = 353;
	{8'd182,8'd172} : s = 354;
	{8'd182,8'd173} : s = 355;
	{8'd182,8'd174} : s = 356;
	{8'd182,8'd175} : s = 357;
	{8'd182,8'd176} : s = 358;
	{8'd182,8'd177} : s = 359;
	{8'd182,8'd178} : s = 360;
	{8'd182,8'd179} : s = 361;
	{8'd182,8'd180} : s = 362;
	{8'd182,8'd181} : s = 363;
	{8'd182,8'd182} : s = 364;
	{8'd182,8'd183} : s = 365;
	{8'd182,8'd184} : s = 366;
	{8'd182,8'd185} : s = 367;
	{8'd182,8'd186} : s = 368;
	{8'd182,8'd187} : s = 369;
	{8'd182,8'd188} : s = 370;
	{8'd182,8'd189} : s = 371;
	{8'd182,8'd190} : s = 372;
	{8'd182,8'd191} : s = 373;
	{8'd182,8'd192} : s = 374;
	{8'd182,8'd193} : s = 375;
	{8'd182,8'd194} : s = 376;
	{8'd182,8'd195} : s = 377;
	{8'd182,8'd196} : s = 378;
	{8'd182,8'd197} : s = 379;
	{8'd182,8'd198} : s = 380;
	{8'd182,8'd199} : s = 381;
	{8'd182,8'd200} : s = 382;
	{8'd182,8'd201} : s = 383;
	{8'd182,8'd202} : s = 384;
	{8'd182,8'd203} : s = 385;
	{8'd182,8'd204} : s = 386;
	{8'd182,8'd205} : s = 387;
	{8'd182,8'd206} : s = 388;
	{8'd182,8'd207} : s = 389;
	{8'd182,8'd208} : s = 390;
	{8'd182,8'd209} : s = 391;
	{8'd182,8'd210} : s = 392;
	{8'd182,8'd211} : s = 393;
	{8'd182,8'd212} : s = 394;
	{8'd182,8'd213} : s = 395;
	{8'd182,8'd214} : s = 396;
	{8'd182,8'd215} : s = 397;
	{8'd182,8'd216} : s = 398;
	{8'd182,8'd217} : s = 399;
	{8'd182,8'd218} : s = 400;
	{8'd182,8'd219} : s = 401;
	{8'd182,8'd220} : s = 402;
	{8'd182,8'd221} : s = 403;
	{8'd182,8'd222} : s = 404;
	{8'd182,8'd223} : s = 405;
	{8'd182,8'd224} : s = 406;
	{8'd182,8'd225} : s = 407;
	{8'd182,8'd226} : s = 408;
	{8'd182,8'd227} : s = 409;
	{8'd182,8'd228} : s = 410;
	{8'd182,8'd229} : s = 411;
	{8'd182,8'd230} : s = 412;
	{8'd182,8'd231} : s = 413;
	{8'd182,8'd232} : s = 414;
	{8'd182,8'd233} : s = 415;
	{8'd182,8'd234} : s = 416;
	{8'd182,8'd235} : s = 417;
	{8'd182,8'd236} : s = 418;
	{8'd182,8'd237} : s = 419;
	{8'd182,8'd238} : s = 420;
	{8'd182,8'd239} : s = 421;
	{8'd182,8'd240} : s = 422;
	{8'd182,8'd241} : s = 423;
	{8'd182,8'd242} : s = 424;
	{8'd182,8'd243} : s = 425;
	{8'd182,8'd244} : s = 426;
	{8'd182,8'd245} : s = 427;
	{8'd182,8'd246} : s = 428;
	{8'd182,8'd247} : s = 429;
	{8'd182,8'd248} : s = 430;
	{8'd182,8'd249} : s = 431;
	{8'd182,8'd250} : s = 432;
	{8'd182,8'd251} : s = 433;
	{8'd182,8'd252} : s = 434;
	{8'd182,8'd253} : s = 435;
	{8'd182,8'd254} : s = 436;
	{8'd182,8'd255} : s = 437;
	{8'd183,8'd0} : s = 183;
	{8'd183,8'd1} : s = 184;
	{8'd183,8'd2} : s = 185;
	{8'd183,8'd3} : s = 186;
	{8'd183,8'd4} : s = 187;
	{8'd183,8'd5} : s = 188;
	{8'd183,8'd6} : s = 189;
	{8'd183,8'd7} : s = 190;
	{8'd183,8'd8} : s = 191;
	{8'd183,8'd9} : s = 192;
	{8'd183,8'd10} : s = 193;
	{8'd183,8'd11} : s = 194;
	{8'd183,8'd12} : s = 195;
	{8'd183,8'd13} : s = 196;
	{8'd183,8'd14} : s = 197;
	{8'd183,8'd15} : s = 198;
	{8'd183,8'd16} : s = 199;
	{8'd183,8'd17} : s = 200;
	{8'd183,8'd18} : s = 201;
	{8'd183,8'd19} : s = 202;
	{8'd183,8'd20} : s = 203;
	{8'd183,8'd21} : s = 204;
	{8'd183,8'd22} : s = 205;
	{8'd183,8'd23} : s = 206;
	{8'd183,8'd24} : s = 207;
	{8'd183,8'd25} : s = 208;
	{8'd183,8'd26} : s = 209;
	{8'd183,8'd27} : s = 210;
	{8'd183,8'd28} : s = 211;
	{8'd183,8'd29} : s = 212;
	{8'd183,8'd30} : s = 213;
	{8'd183,8'd31} : s = 214;
	{8'd183,8'd32} : s = 215;
	{8'd183,8'd33} : s = 216;
	{8'd183,8'd34} : s = 217;
	{8'd183,8'd35} : s = 218;
	{8'd183,8'd36} : s = 219;
	{8'd183,8'd37} : s = 220;
	{8'd183,8'd38} : s = 221;
	{8'd183,8'd39} : s = 222;
	{8'd183,8'd40} : s = 223;
	{8'd183,8'd41} : s = 224;
	{8'd183,8'd42} : s = 225;
	{8'd183,8'd43} : s = 226;
	{8'd183,8'd44} : s = 227;
	{8'd183,8'd45} : s = 228;
	{8'd183,8'd46} : s = 229;
	{8'd183,8'd47} : s = 230;
	{8'd183,8'd48} : s = 231;
	{8'd183,8'd49} : s = 232;
	{8'd183,8'd50} : s = 233;
	{8'd183,8'd51} : s = 234;
	{8'd183,8'd52} : s = 235;
	{8'd183,8'd53} : s = 236;
	{8'd183,8'd54} : s = 237;
	{8'd183,8'd55} : s = 238;
	{8'd183,8'd56} : s = 239;
	{8'd183,8'd57} : s = 240;
	{8'd183,8'd58} : s = 241;
	{8'd183,8'd59} : s = 242;
	{8'd183,8'd60} : s = 243;
	{8'd183,8'd61} : s = 244;
	{8'd183,8'd62} : s = 245;
	{8'd183,8'd63} : s = 246;
	{8'd183,8'd64} : s = 247;
	{8'd183,8'd65} : s = 248;
	{8'd183,8'd66} : s = 249;
	{8'd183,8'd67} : s = 250;
	{8'd183,8'd68} : s = 251;
	{8'd183,8'd69} : s = 252;
	{8'd183,8'd70} : s = 253;
	{8'd183,8'd71} : s = 254;
	{8'd183,8'd72} : s = 255;
	{8'd183,8'd73} : s = 256;
	{8'd183,8'd74} : s = 257;
	{8'd183,8'd75} : s = 258;
	{8'd183,8'd76} : s = 259;
	{8'd183,8'd77} : s = 260;
	{8'd183,8'd78} : s = 261;
	{8'd183,8'd79} : s = 262;
	{8'd183,8'd80} : s = 263;
	{8'd183,8'd81} : s = 264;
	{8'd183,8'd82} : s = 265;
	{8'd183,8'd83} : s = 266;
	{8'd183,8'd84} : s = 267;
	{8'd183,8'd85} : s = 268;
	{8'd183,8'd86} : s = 269;
	{8'd183,8'd87} : s = 270;
	{8'd183,8'd88} : s = 271;
	{8'd183,8'd89} : s = 272;
	{8'd183,8'd90} : s = 273;
	{8'd183,8'd91} : s = 274;
	{8'd183,8'd92} : s = 275;
	{8'd183,8'd93} : s = 276;
	{8'd183,8'd94} : s = 277;
	{8'd183,8'd95} : s = 278;
	{8'd183,8'd96} : s = 279;
	{8'd183,8'd97} : s = 280;
	{8'd183,8'd98} : s = 281;
	{8'd183,8'd99} : s = 282;
	{8'd183,8'd100} : s = 283;
	{8'd183,8'd101} : s = 284;
	{8'd183,8'd102} : s = 285;
	{8'd183,8'd103} : s = 286;
	{8'd183,8'd104} : s = 287;
	{8'd183,8'd105} : s = 288;
	{8'd183,8'd106} : s = 289;
	{8'd183,8'd107} : s = 290;
	{8'd183,8'd108} : s = 291;
	{8'd183,8'd109} : s = 292;
	{8'd183,8'd110} : s = 293;
	{8'd183,8'd111} : s = 294;
	{8'd183,8'd112} : s = 295;
	{8'd183,8'd113} : s = 296;
	{8'd183,8'd114} : s = 297;
	{8'd183,8'd115} : s = 298;
	{8'd183,8'd116} : s = 299;
	{8'd183,8'd117} : s = 300;
	{8'd183,8'd118} : s = 301;
	{8'd183,8'd119} : s = 302;
	{8'd183,8'd120} : s = 303;
	{8'd183,8'd121} : s = 304;
	{8'd183,8'd122} : s = 305;
	{8'd183,8'd123} : s = 306;
	{8'd183,8'd124} : s = 307;
	{8'd183,8'd125} : s = 308;
	{8'd183,8'd126} : s = 309;
	{8'd183,8'd127} : s = 310;
	{8'd183,8'd128} : s = 311;
	{8'd183,8'd129} : s = 312;
	{8'd183,8'd130} : s = 313;
	{8'd183,8'd131} : s = 314;
	{8'd183,8'd132} : s = 315;
	{8'd183,8'd133} : s = 316;
	{8'd183,8'd134} : s = 317;
	{8'd183,8'd135} : s = 318;
	{8'd183,8'd136} : s = 319;
	{8'd183,8'd137} : s = 320;
	{8'd183,8'd138} : s = 321;
	{8'd183,8'd139} : s = 322;
	{8'd183,8'd140} : s = 323;
	{8'd183,8'd141} : s = 324;
	{8'd183,8'd142} : s = 325;
	{8'd183,8'd143} : s = 326;
	{8'd183,8'd144} : s = 327;
	{8'd183,8'd145} : s = 328;
	{8'd183,8'd146} : s = 329;
	{8'd183,8'd147} : s = 330;
	{8'd183,8'd148} : s = 331;
	{8'd183,8'd149} : s = 332;
	{8'd183,8'd150} : s = 333;
	{8'd183,8'd151} : s = 334;
	{8'd183,8'd152} : s = 335;
	{8'd183,8'd153} : s = 336;
	{8'd183,8'd154} : s = 337;
	{8'd183,8'd155} : s = 338;
	{8'd183,8'd156} : s = 339;
	{8'd183,8'd157} : s = 340;
	{8'd183,8'd158} : s = 341;
	{8'd183,8'd159} : s = 342;
	{8'd183,8'd160} : s = 343;
	{8'd183,8'd161} : s = 344;
	{8'd183,8'd162} : s = 345;
	{8'd183,8'd163} : s = 346;
	{8'd183,8'd164} : s = 347;
	{8'd183,8'd165} : s = 348;
	{8'd183,8'd166} : s = 349;
	{8'd183,8'd167} : s = 350;
	{8'd183,8'd168} : s = 351;
	{8'd183,8'd169} : s = 352;
	{8'd183,8'd170} : s = 353;
	{8'd183,8'd171} : s = 354;
	{8'd183,8'd172} : s = 355;
	{8'd183,8'd173} : s = 356;
	{8'd183,8'd174} : s = 357;
	{8'd183,8'd175} : s = 358;
	{8'd183,8'd176} : s = 359;
	{8'd183,8'd177} : s = 360;
	{8'd183,8'd178} : s = 361;
	{8'd183,8'd179} : s = 362;
	{8'd183,8'd180} : s = 363;
	{8'd183,8'd181} : s = 364;
	{8'd183,8'd182} : s = 365;
	{8'd183,8'd183} : s = 366;
	{8'd183,8'd184} : s = 367;
	{8'd183,8'd185} : s = 368;
	{8'd183,8'd186} : s = 369;
	{8'd183,8'd187} : s = 370;
	{8'd183,8'd188} : s = 371;
	{8'd183,8'd189} : s = 372;
	{8'd183,8'd190} : s = 373;
	{8'd183,8'd191} : s = 374;
	{8'd183,8'd192} : s = 375;
	{8'd183,8'd193} : s = 376;
	{8'd183,8'd194} : s = 377;
	{8'd183,8'd195} : s = 378;
	{8'd183,8'd196} : s = 379;
	{8'd183,8'd197} : s = 380;
	{8'd183,8'd198} : s = 381;
	{8'd183,8'd199} : s = 382;
	{8'd183,8'd200} : s = 383;
	{8'd183,8'd201} : s = 384;
	{8'd183,8'd202} : s = 385;
	{8'd183,8'd203} : s = 386;
	{8'd183,8'd204} : s = 387;
	{8'd183,8'd205} : s = 388;
	{8'd183,8'd206} : s = 389;
	{8'd183,8'd207} : s = 390;
	{8'd183,8'd208} : s = 391;
	{8'd183,8'd209} : s = 392;
	{8'd183,8'd210} : s = 393;
	{8'd183,8'd211} : s = 394;
	{8'd183,8'd212} : s = 395;
	{8'd183,8'd213} : s = 396;
	{8'd183,8'd214} : s = 397;
	{8'd183,8'd215} : s = 398;
	{8'd183,8'd216} : s = 399;
	{8'd183,8'd217} : s = 400;
	{8'd183,8'd218} : s = 401;
	{8'd183,8'd219} : s = 402;
	{8'd183,8'd220} : s = 403;
	{8'd183,8'd221} : s = 404;
	{8'd183,8'd222} : s = 405;
	{8'd183,8'd223} : s = 406;
	{8'd183,8'd224} : s = 407;
	{8'd183,8'd225} : s = 408;
	{8'd183,8'd226} : s = 409;
	{8'd183,8'd227} : s = 410;
	{8'd183,8'd228} : s = 411;
	{8'd183,8'd229} : s = 412;
	{8'd183,8'd230} : s = 413;
	{8'd183,8'd231} : s = 414;
	{8'd183,8'd232} : s = 415;
	{8'd183,8'd233} : s = 416;
	{8'd183,8'd234} : s = 417;
	{8'd183,8'd235} : s = 418;
	{8'd183,8'd236} : s = 419;
	{8'd183,8'd237} : s = 420;
	{8'd183,8'd238} : s = 421;
	{8'd183,8'd239} : s = 422;
	{8'd183,8'd240} : s = 423;
	{8'd183,8'd241} : s = 424;
	{8'd183,8'd242} : s = 425;
	{8'd183,8'd243} : s = 426;
	{8'd183,8'd244} : s = 427;
	{8'd183,8'd245} : s = 428;
	{8'd183,8'd246} : s = 429;
	{8'd183,8'd247} : s = 430;
	{8'd183,8'd248} : s = 431;
	{8'd183,8'd249} : s = 432;
	{8'd183,8'd250} : s = 433;
	{8'd183,8'd251} : s = 434;
	{8'd183,8'd252} : s = 435;
	{8'd183,8'd253} : s = 436;
	{8'd183,8'd254} : s = 437;
	{8'd183,8'd255} : s = 438;
	{8'd184,8'd0} : s = 184;
	{8'd184,8'd1} : s = 185;
	{8'd184,8'd2} : s = 186;
	{8'd184,8'd3} : s = 187;
	{8'd184,8'd4} : s = 188;
	{8'd184,8'd5} : s = 189;
	{8'd184,8'd6} : s = 190;
	{8'd184,8'd7} : s = 191;
	{8'd184,8'd8} : s = 192;
	{8'd184,8'd9} : s = 193;
	{8'd184,8'd10} : s = 194;
	{8'd184,8'd11} : s = 195;
	{8'd184,8'd12} : s = 196;
	{8'd184,8'd13} : s = 197;
	{8'd184,8'd14} : s = 198;
	{8'd184,8'd15} : s = 199;
	{8'd184,8'd16} : s = 200;
	{8'd184,8'd17} : s = 201;
	{8'd184,8'd18} : s = 202;
	{8'd184,8'd19} : s = 203;
	{8'd184,8'd20} : s = 204;
	{8'd184,8'd21} : s = 205;
	{8'd184,8'd22} : s = 206;
	{8'd184,8'd23} : s = 207;
	{8'd184,8'd24} : s = 208;
	{8'd184,8'd25} : s = 209;
	{8'd184,8'd26} : s = 210;
	{8'd184,8'd27} : s = 211;
	{8'd184,8'd28} : s = 212;
	{8'd184,8'd29} : s = 213;
	{8'd184,8'd30} : s = 214;
	{8'd184,8'd31} : s = 215;
	{8'd184,8'd32} : s = 216;
	{8'd184,8'd33} : s = 217;
	{8'd184,8'd34} : s = 218;
	{8'd184,8'd35} : s = 219;
	{8'd184,8'd36} : s = 220;
	{8'd184,8'd37} : s = 221;
	{8'd184,8'd38} : s = 222;
	{8'd184,8'd39} : s = 223;
	{8'd184,8'd40} : s = 224;
	{8'd184,8'd41} : s = 225;
	{8'd184,8'd42} : s = 226;
	{8'd184,8'd43} : s = 227;
	{8'd184,8'd44} : s = 228;
	{8'd184,8'd45} : s = 229;
	{8'd184,8'd46} : s = 230;
	{8'd184,8'd47} : s = 231;
	{8'd184,8'd48} : s = 232;
	{8'd184,8'd49} : s = 233;
	{8'd184,8'd50} : s = 234;
	{8'd184,8'd51} : s = 235;
	{8'd184,8'd52} : s = 236;
	{8'd184,8'd53} : s = 237;
	{8'd184,8'd54} : s = 238;
	{8'd184,8'd55} : s = 239;
	{8'd184,8'd56} : s = 240;
	{8'd184,8'd57} : s = 241;
	{8'd184,8'd58} : s = 242;
	{8'd184,8'd59} : s = 243;
	{8'd184,8'd60} : s = 244;
	{8'd184,8'd61} : s = 245;
	{8'd184,8'd62} : s = 246;
	{8'd184,8'd63} : s = 247;
	{8'd184,8'd64} : s = 248;
	{8'd184,8'd65} : s = 249;
	{8'd184,8'd66} : s = 250;
	{8'd184,8'd67} : s = 251;
	{8'd184,8'd68} : s = 252;
	{8'd184,8'd69} : s = 253;
	{8'd184,8'd70} : s = 254;
	{8'd184,8'd71} : s = 255;
	{8'd184,8'd72} : s = 256;
	{8'd184,8'd73} : s = 257;
	{8'd184,8'd74} : s = 258;
	{8'd184,8'd75} : s = 259;
	{8'd184,8'd76} : s = 260;
	{8'd184,8'd77} : s = 261;
	{8'd184,8'd78} : s = 262;
	{8'd184,8'd79} : s = 263;
	{8'd184,8'd80} : s = 264;
	{8'd184,8'd81} : s = 265;
	{8'd184,8'd82} : s = 266;
	{8'd184,8'd83} : s = 267;
	{8'd184,8'd84} : s = 268;
	{8'd184,8'd85} : s = 269;
	{8'd184,8'd86} : s = 270;
	{8'd184,8'd87} : s = 271;
	{8'd184,8'd88} : s = 272;
	{8'd184,8'd89} : s = 273;
	{8'd184,8'd90} : s = 274;
	{8'd184,8'd91} : s = 275;
	{8'd184,8'd92} : s = 276;
	{8'd184,8'd93} : s = 277;
	{8'd184,8'd94} : s = 278;
	{8'd184,8'd95} : s = 279;
	{8'd184,8'd96} : s = 280;
	{8'd184,8'd97} : s = 281;
	{8'd184,8'd98} : s = 282;
	{8'd184,8'd99} : s = 283;
	{8'd184,8'd100} : s = 284;
	{8'd184,8'd101} : s = 285;
	{8'd184,8'd102} : s = 286;
	{8'd184,8'd103} : s = 287;
	{8'd184,8'd104} : s = 288;
	{8'd184,8'd105} : s = 289;
	{8'd184,8'd106} : s = 290;
	{8'd184,8'd107} : s = 291;
	{8'd184,8'd108} : s = 292;
	{8'd184,8'd109} : s = 293;
	{8'd184,8'd110} : s = 294;
	{8'd184,8'd111} : s = 295;
	{8'd184,8'd112} : s = 296;
	{8'd184,8'd113} : s = 297;
	{8'd184,8'd114} : s = 298;
	{8'd184,8'd115} : s = 299;
	{8'd184,8'd116} : s = 300;
	{8'd184,8'd117} : s = 301;
	{8'd184,8'd118} : s = 302;
	{8'd184,8'd119} : s = 303;
	{8'd184,8'd120} : s = 304;
	{8'd184,8'd121} : s = 305;
	{8'd184,8'd122} : s = 306;
	{8'd184,8'd123} : s = 307;
	{8'd184,8'd124} : s = 308;
	{8'd184,8'd125} : s = 309;
	{8'd184,8'd126} : s = 310;
	{8'd184,8'd127} : s = 311;
	{8'd184,8'd128} : s = 312;
	{8'd184,8'd129} : s = 313;
	{8'd184,8'd130} : s = 314;
	{8'd184,8'd131} : s = 315;
	{8'd184,8'd132} : s = 316;
	{8'd184,8'd133} : s = 317;
	{8'd184,8'd134} : s = 318;
	{8'd184,8'd135} : s = 319;
	{8'd184,8'd136} : s = 320;
	{8'd184,8'd137} : s = 321;
	{8'd184,8'd138} : s = 322;
	{8'd184,8'd139} : s = 323;
	{8'd184,8'd140} : s = 324;
	{8'd184,8'd141} : s = 325;
	{8'd184,8'd142} : s = 326;
	{8'd184,8'd143} : s = 327;
	{8'd184,8'd144} : s = 328;
	{8'd184,8'd145} : s = 329;
	{8'd184,8'd146} : s = 330;
	{8'd184,8'd147} : s = 331;
	{8'd184,8'd148} : s = 332;
	{8'd184,8'd149} : s = 333;
	{8'd184,8'd150} : s = 334;
	{8'd184,8'd151} : s = 335;
	{8'd184,8'd152} : s = 336;
	{8'd184,8'd153} : s = 337;
	{8'd184,8'd154} : s = 338;
	{8'd184,8'd155} : s = 339;
	{8'd184,8'd156} : s = 340;
	{8'd184,8'd157} : s = 341;
	{8'd184,8'd158} : s = 342;
	{8'd184,8'd159} : s = 343;
	{8'd184,8'd160} : s = 344;
	{8'd184,8'd161} : s = 345;
	{8'd184,8'd162} : s = 346;
	{8'd184,8'd163} : s = 347;
	{8'd184,8'd164} : s = 348;
	{8'd184,8'd165} : s = 349;
	{8'd184,8'd166} : s = 350;
	{8'd184,8'd167} : s = 351;
	{8'd184,8'd168} : s = 352;
	{8'd184,8'd169} : s = 353;
	{8'd184,8'd170} : s = 354;
	{8'd184,8'd171} : s = 355;
	{8'd184,8'd172} : s = 356;
	{8'd184,8'd173} : s = 357;
	{8'd184,8'd174} : s = 358;
	{8'd184,8'd175} : s = 359;
	{8'd184,8'd176} : s = 360;
	{8'd184,8'd177} : s = 361;
	{8'd184,8'd178} : s = 362;
	{8'd184,8'd179} : s = 363;
	{8'd184,8'd180} : s = 364;
	{8'd184,8'd181} : s = 365;
	{8'd184,8'd182} : s = 366;
	{8'd184,8'd183} : s = 367;
	{8'd184,8'd184} : s = 368;
	{8'd184,8'd185} : s = 369;
	{8'd184,8'd186} : s = 370;
	{8'd184,8'd187} : s = 371;
	{8'd184,8'd188} : s = 372;
	{8'd184,8'd189} : s = 373;
	{8'd184,8'd190} : s = 374;
	{8'd184,8'd191} : s = 375;
	{8'd184,8'd192} : s = 376;
	{8'd184,8'd193} : s = 377;
	{8'd184,8'd194} : s = 378;
	{8'd184,8'd195} : s = 379;
	{8'd184,8'd196} : s = 380;
	{8'd184,8'd197} : s = 381;
	{8'd184,8'd198} : s = 382;
	{8'd184,8'd199} : s = 383;
	{8'd184,8'd200} : s = 384;
	{8'd184,8'd201} : s = 385;
	{8'd184,8'd202} : s = 386;
	{8'd184,8'd203} : s = 387;
	{8'd184,8'd204} : s = 388;
	{8'd184,8'd205} : s = 389;
	{8'd184,8'd206} : s = 390;
	{8'd184,8'd207} : s = 391;
	{8'd184,8'd208} : s = 392;
	{8'd184,8'd209} : s = 393;
	{8'd184,8'd210} : s = 394;
	{8'd184,8'd211} : s = 395;
	{8'd184,8'd212} : s = 396;
	{8'd184,8'd213} : s = 397;
	{8'd184,8'd214} : s = 398;
	{8'd184,8'd215} : s = 399;
	{8'd184,8'd216} : s = 400;
	{8'd184,8'd217} : s = 401;
	{8'd184,8'd218} : s = 402;
	{8'd184,8'd219} : s = 403;
	{8'd184,8'd220} : s = 404;
	{8'd184,8'd221} : s = 405;
	{8'd184,8'd222} : s = 406;
	{8'd184,8'd223} : s = 407;
	{8'd184,8'd224} : s = 408;
	{8'd184,8'd225} : s = 409;
	{8'd184,8'd226} : s = 410;
	{8'd184,8'd227} : s = 411;
	{8'd184,8'd228} : s = 412;
	{8'd184,8'd229} : s = 413;
	{8'd184,8'd230} : s = 414;
	{8'd184,8'd231} : s = 415;
	{8'd184,8'd232} : s = 416;
	{8'd184,8'd233} : s = 417;
	{8'd184,8'd234} : s = 418;
	{8'd184,8'd235} : s = 419;
	{8'd184,8'd236} : s = 420;
	{8'd184,8'd237} : s = 421;
	{8'd184,8'd238} : s = 422;
	{8'd184,8'd239} : s = 423;
	{8'd184,8'd240} : s = 424;
	{8'd184,8'd241} : s = 425;
	{8'd184,8'd242} : s = 426;
	{8'd184,8'd243} : s = 427;
	{8'd184,8'd244} : s = 428;
	{8'd184,8'd245} : s = 429;
	{8'd184,8'd246} : s = 430;
	{8'd184,8'd247} : s = 431;
	{8'd184,8'd248} : s = 432;
	{8'd184,8'd249} : s = 433;
	{8'd184,8'd250} : s = 434;
	{8'd184,8'd251} : s = 435;
	{8'd184,8'd252} : s = 436;
	{8'd184,8'd253} : s = 437;
	{8'd184,8'd254} : s = 438;
	{8'd184,8'd255} : s = 439;
	{8'd185,8'd0} : s = 185;
	{8'd185,8'd1} : s = 186;
	{8'd185,8'd2} : s = 187;
	{8'd185,8'd3} : s = 188;
	{8'd185,8'd4} : s = 189;
	{8'd185,8'd5} : s = 190;
	{8'd185,8'd6} : s = 191;
	{8'd185,8'd7} : s = 192;
	{8'd185,8'd8} : s = 193;
	{8'd185,8'd9} : s = 194;
	{8'd185,8'd10} : s = 195;
	{8'd185,8'd11} : s = 196;
	{8'd185,8'd12} : s = 197;
	{8'd185,8'd13} : s = 198;
	{8'd185,8'd14} : s = 199;
	{8'd185,8'd15} : s = 200;
	{8'd185,8'd16} : s = 201;
	{8'd185,8'd17} : s = 202;
	{8'd185,8'd18} : s = 203;
	{8'd185,8'd19} : s = 204;
	{8'd185,8'd20} : s = 205;
	{8'd185,8'd21} : s = 206;
	{8'd185,8'd22} : s = 207;
	{8'd185,8'd23} : s = 208;
	{8'd185,8'd24} : s = 209;
	{8'd185,8'd25} : s = 210;
	{8'd185,8'd26} : s = 211;
	{8'd185,8'd27} : s = 212;
	{8'd185,8'd28} : s = 213;
	{8'd185,8'd29} : s = 214;
	{8'd185,8'd30} : s = 215;
	{8'd185,8'd31} : s = 216;
	{8'd185,8'd32} : s = 217;
	{8'd185,8'd33} : s = 218;
	{8'd185,8'd34} : s = 219;
	{8'd185,8'd35} : s = 220;
	{8'd185,8'd36} : s = 221;
	{8'd185,8'd37} : s = 222;
	{8'd185,8'd38} : s = 223;
	{8'd185,8'd39} : s = 224;
	{8'd185,8'd40} : s = 225;
	{8'd185,8'd41} : s = 226;
	{8'd185,8'd42} : s = 227;
	{8'd185,8'd43} : s = 228;
	{8'd185,8'd44} : s = 229;
	{8'd185,8'd45} : s = 230;
	{8'd185,8'd46} : s = 231;
	{8'd185,8'd47} : s = 232;
	{8'd185,8'd48} : s = 233;
	{8'd185,8'd49} : s = 234;
	{8'd185,8'd50} : s = 235;
	{8'd185,8'd51} : s = 236;
	{8'd185,8'd52} : s = 237;
	{8'd185,8'd53} : s = 238;
	{8'd185,8'd54} : s = 239;
	{8'd185,8'd55} : s = 240;
	{8'd185,8'd56} : s = 241;
	{8'd185,8'd57} : s = 242;
	{8'd185,8'd58} : s = 243;
	{8'd185,8'd59} : s = 244;
	{8'd185,8'd60} : s = 245;
	{8'd185,8'd61} : s = 246;
	{8'd185,8'd62} : s = 247;
	{8'd185,8'd63} : s = 248;
	{8'd185,8'd64} : s = 249;
	{8'd185,8'd65} : s = 250;
	{8'd185,8'd66} : s = 251;
	{8'd185,8'd67} : s = 252;
	{8'd185,8'd68} : s = 253;
	{8'd185,8'd69} : s = 254;
	{8'd185,8'd70} : s = 255;
	{8'd185,8'd71} : s = 256;
	{8'd185,8'd72} : s = 257;
	{8'd185,8'd73} : s = 258;
	{8'd185,8'd74} : s = 259;
	{8'd185,8'd75} : s = 260;
	{8'd185,8'd76} : s = 261;
	{8'd185,8'd77} : s = 262;
	{8'd185,8'd78} : s = 263;
	{8'd185,8'd79} : s = 264;
	{8'd185,8'd80} : s = 265;
	{8'd185,8'd81} : s = 266;
	{8'd185,8'd82} : s = 267;
	{8'd185,8'd83} : s = 268;
	{8'd185,8'd84} : s = 269;
	{8'd185,8'd85} : s = 270;
	{8'd185,8'd86} : s = 271;
	{8'd185,8'd87} : s = 272;
	{8'd185,8'd88} : s = 273;
	{8'd185,8'd89} : s = 274;
	{8'd185,8'd90} : s = 275;
	{8'd185,8'd91} : s = 276;
	{8'd185,8'd92} : s = 277;
	{8'd185,8'd93} : s = 278;
	{8'd185,8'd94} : s = 279;
	{8'd185,8'd95} : s = 280;
	{8'd185,8'd96} : s = 281;
	{8'd185,8'd97} : s = 282;
	{8'd185,8'd98} : s = 283;
	{8'd185,8'd99} : s = 284;
	{8'd185,8'd100} : s = 285;
	{8'd185,8'd101} : s = 286;
	{8'd185,8'd102} : s = 287;
	{8'd185,8'd103} : s = 288;
	{8'd185,8'd104} : s = 289;
	{8'd185,8'd105} : s = 290;
	{8'd185,8'd106} : s = 291;
	{8'd185,8'd107} : s = 292;
	{8'd185,8'd108} : s = 293;
	{8'd185,8'd109} : s = 294;
	{8'd185,8'd110} : s = 295;
	{8'd185,8'd111} : s = 296;
	{8'd185,8'd112} : s = 297;
	{8'd185,8'd113} : s = 298;
	{8'd185,8'd114} : s = 299;
	{8'd185,8'd115} : s = 300;
	{8'd185,8'd116} : s = 301;
	{8'd185,8'd117} : s = 302;
	{8'd185,8'd118} : s = 303;
	{8'd185,8'd119} : s = 304;
	{8'd185,8'd120} : s = 305;
	{8'd185,8'd121} : s = 306;
	{8'd185,8'd122} : s = 307;
	{8'd185,8'd123} : s = 308;
	{8'd185,8'd124} : s = 309;
	{8'd185,8'd125} : s = 310;
	{8'd185,8'd126} : s = 311;
	{8'd185,8'd127} : s = 312;
	{8'd185,8'd128} : s = 313;
	{8'd185,8'd129} : s = 314;
	{8'd185,8'd130} : s = 315;
	{8'd185,8'd131} : s = 316;
	{8'd185,8'd132} : s = 317;
	{8'd185,8'd133} : s = 318;
	{8'd185,8'd134} : s = 319;
	{8'd185,8'd135} : s = 320;
	{8'd185,8'd136} : s = 321;
	{8'd185,8'd137} : s = 322;
	{8'd185,8'd138} : s = 323;
	{8'd185,8'd139} : s = 324;
	{8'd185,8'd140} : s = 325;
	{8'd185,8'd141} : s = 326;
	{8'd185,8'd142} : s = 327;
	{8'd185,8'd143} : s = 328;
	{8'd185,8'd144} : s = 329;
	{8'd185,8'd145} : s = 330;
	{8'd185,8'd146} : s = 331;
	{8'd185,8'd147} : s = 332;
	{8'd185,8'd148} : s = 333;
	{8'd185,8'd149} : s = 334;
	{8'd185,8'd150} : s = 335;
	{8'd185,8'd151} : s = 336;
	{8'd185,8'd152} : s = 337;
	{8'd185,8'd153} : s = 338;
	{8'd185,8'd154} : s = 339;
	{8'd185,8'd155} : s = 340;
	{8'd185,8'd156} : s = 341;
	{8'd185,8'd157} : s = 342;
	{8'd185,8'd158} : s = 343;
	{8'd185,8'd159} : s = 344;
	{8'd185,8'd160} : s = 345;
	{8'd185,8'd161} : s = 346;
	{8'd185,8'd162} : s = 347;
	{8'd185,8'd163} : s = 348;
	{8'd185,8'd164} : s = 349;
	{8'd185,8'd165} : s = 350;
	{8'd185,8'd166} : s = 351;
	{8'd185,8'd167} : s = 352;
	{8'd185,8'd168} : s = 353;
	{8'd185,8'd169} : s = 354;
	{8'd185,8'd170} : s = 355;
	{8'd185,8'd171} : s = 356;
	{8'd185,8'd172} : s = 357;
	{8'd185,8'd173} : s = 358;
	{8'd185,8'd174} : s = 359;
	{8'd185,8'd175} : s = 360;
	{8'd185,8'd176} : s = 361;
	{8'd185,8'd177} : s = 362;
	{8'd185,8'd178} : s = 363;
	{8'd185,8'd179} : s = 364;
	{8'd185,8'd180} : s = 365;
	{8'd185,8'd181} : s = 366;
	{8'd185,8'd182} : s = 367;
	{8'd185,8'd183} : s = 368;
	{8'd185,8'd184} : s = 369;
	{8'd185,8'd185} : s = 370;
	{8'd185,8'd186} : s = 371;
	{8'd185,8'd187} : s = 372;
	{8'd185,8'd188} : s = 373;
	{8'd185,8'd189} : s = 374;
	{8'd185,8'd190} : s = 375;
	{8'd185,8'd191} : s = 376;
	{8'd185,8'd192} : s = 377;
	{8'd185,8'd193} : s = 378;
	{8'd185,8'd194} : s = 379;
	{8'd185,8'd195} : s = 380;
	{8'd185,8'd196} : s = 381;
	{8'd185,8'd197} : s = 382;
	{8'd185,8'd198} : s = 383;
	{8'd185,8'd199} : s = 384;
	{8'd185,8'd200} : s = 385;
	{8'd185,8'd201} : s = 386;
	{8'd185,8'd202} : s = 387;
	{8'd185,8'd203} : s = 388;
	{8'd185,8'd204} : s = 389;
	{8'd185,8'd205} : s = 390;
	{8'd185,8'd206} : s = 391;
	{8'd185,8'd207} : s = 392;
	{8'd185,8'd208} : s = 393;
	{8'd185,8'd209} : s = 394;
	{8'd185,8'd210} : s = 395;
	{8'd185,8'd211} : s = 396;
	{8'd185,8'd212} : s = 397;
	{8'd185,8'd213} : s = 398;
	{8'd185,8'd214} : s = 399;
	{8'd185,8'd215} : s = 400;
	{8'd185,8'd216} : s = 401;
	{8'd185,8'd217} : s = 402;
	{8'd185,8'd218} : s = 403;
	{8'd185,8'd219} : s = 404;
	{8'd185,8'd220} : s = 405;
	{8'd185,8'd221} : s = 406;
	{8'd185,8'd222} : s = 407;
	{8'd185,8'd223} : s = 408;
	{8'd185,8'd224} : s = 409;
	{8'd185,8'd225} : s = 410;
	{8'd185,8'd226} : s = 411;
	{8'd185,8'd227} : s = 412;
	{8'd185,8'd228} : s = 413;
	{8'd185,8'd229} : s = 414;
	{8'd185,8'd230} : s = 415;
	{8'd185,8'd231} : s = 416;
	{8'd185,8'd232} : s = 417;
	{8'd185,8'd233} : s = 418;
	{8'd185,8'd234} : s = 419;
	{8'd185,8'd235} : s = 420;
	{8'd185,8'd236} : s = 421;
	{8'd185,8'd237} : s = 422;
	{8'd185,8'd238} : s = 423;
	{8'd185,8'd239} : s = 424;
	{8'd185,8'd240} : s = 425;
	{8'd185,8'd241} : s = 426;
	{8'd185,8'd242} : s = 427;
	{8'd185,8'd243} : s = 428;
	{8'd185,8'd244} : s = 429;
	{8'd185,8'd245} : s = 430;
	{8'd185,8'd246} : s = 431;
	{8'd185,8'd247} : s = 432;
	{8'd185,8'd248} : s = 433;
	{8'd185,8'd249} : s = 434;
	{8'd185,8'd250} : s = 435;
	{8'd185,8'd251} : s = 436;
	{8'd185,8'd252} : s = 437;
	{8'd185,8'd253} : s = 438;
	{8'd185,8'd254} : s = 439;
	{8'd185,8'd255} : s = 440;
	{8'd186,8'd0} : s = 186;
	{8'd186,8'd1} : s = 187;
	{8'd186,8'd2} : s = 188;
	{8'd186,8'd3} : s = 189;
	{8'd186,8'd4} : s = 190;
	{8'd186,8'd5} : s = 191;
	{8'd186,8'd6} : s = 192;
	{8'd186,8'd7} : s = 193;
	{8'd186,8'd8} : s = 194;
	{8'd186,8'd9} : s = 195;
	{8'd186,8'd10} : s = 196;
	{8'd186,8'd11} : s = 197;
	{8'd186,8'd12} : s = 198;
	{8'd186,8'd13} : s = 199;
	{8'd186,8'd14} : s = 200;
	{8'd186,8'd15} : s = 201;
	{8'd186,8'd16} : s = 202;
	{8'd186,8'd17} : s = 203;
	{8'd186,8'd18} : s = 204;
	{8'd186,8'd19} : s = 205;
	{8'd186,8'd20} : s = 206;
	{8'd186,8'd21} : s = 207;
	{8'd186,8'd22} : s = 208;
	{8'd186,8'd23} : s = 209;
	{8'd186,8'd24} : s = 210;
	{8'd186,8'd25} : s = 211;
	{8'd186,8'd26} : s = 212;
	{8'd186,8'd27} : s = 213;
	{8'd186,8'd28} : s = 214;
	{8'd186,8'd29} : s = 215;
	{8'd186,8'd30} : s = 216;
	{8'd186,8'd31} : s = 217;
	{8'd186,8'd32} : s = 218;
	{8'd186,8'd33} : s = 219;
	{8'd186,8'd34} : s = 220;
	{8'd186,8'd35} : s = 221;
	{8'd186,8'd36} : s = 222;
	{8'd186,8'd37} : s = 223;
	{8'd186,8'd38} : s = 224;
	{8'd186,8'd39} : s = 225;
	{8'd186,8'd40} : s = 226;
	{8'd186,8'd41} : s = 227;
	{8'd186,8'd42} : s = 228;
	{8'd186,8'd43} : s = 229;
	{8'd186,8'd44} : s = 230;
	{8'd186,8'd45} : s = 231;
	{8'd186,8'd46} : s = 232;
	{8'd186,8'd47} : s = 233;
	{8'd186,8'd48} : s = 234;
	{8'd186,8'd49} : s = 235;
	{8'd186,8'd50} : s = 236;
	{8'd186,8'd51} : s = 237;
	{8'd186,8'd52} : s = 238;
	{8'd186,8'd53} : s = 239;
	{8'd186,8'd54} : s = 240;
	{8'd186,8'd55} : s = 241;
	{8'd186,8'd56} : s = 242;
	{8'd186,8'd57} : s = 243;
	{8'd186,8'd58} : s = 244;
	{8'd186,8'd59} : s = 245;
	{8'd186,8'd60} : s = 246;
	{8'd186,8'd61} : s = 247;
	{8'd186,8'd62} : s = 248;
	{8'd186,8'd63} : s = 249;
	{8'd186,8'd64} : s = 250;
	{8'd186,8'd65} : s = 251;
	{8'd186,8'd66} : s = 252;
	{8'd186,8'd67} : s = 253;
	{8'd186,8'd68} : s = 254;
	{8'd186,8'd69} : s = 255;
	{8'd186,8'd70} : s = 256;
	{8'd186,8'd71} : s = 257;
	{8'd186,8'd72} : s = 258;
	{8'd186,8'd73} : s = 259;
	{8'd186,8'd74} : s = 260;
	{8'd186,8'd75} : s = 261;
	{8'd186,8'd76} : s = 262;
	{8'd186,8'd77} : s = 263;
	{8'd186,8'd78} : s = 264;
	{8'd186,8'd79} : s = 265;
	{8'd186,8'd80} : s = 266;
	{8'd186,8'd81} : s = 267;
	{8'd186,8'd82} : s = 268;
	{8'd186,8'd83} : s = 269;
	{8'd186,8'd84} : s = 270;
	{8'd186,8'd85} : s = 271;
	{8'd186,8'd86} : s = 272;
	{8'd186,8'd87} : s = 273;
	{8'd186,8'd88} : s = 274;
	{8'd186,8'd89} : s = 275;
	{8'd186,8'd90} : s = 276;
	{8'd186,8'd91} : s = 277;
	{8'd186,8'd92} : s = 278;
	{8'd186,8'd93} : s = 279;
	{8'd186,8'd94} : s = 280;
	{8'd186,8'd95} : s = 281;
	{8'd186,8'd96} : s = 282;
	{8'd186,8'd97} : s = 283;
	{8'd186,8'd98} : s = 284;
	{8'd186,8'd99} : s = 285;
	{8'd186,8'd100} : s = 286;
	{8'd186,8'd101} : s = 287;
	{8'd186,8'd102} : s = 288;
	{8'd186,8'd103} : s = 289;
	{8'd186,8'd104} : s = 290;
	{8'd186,8'd105} : s = 291;
	{8'd186,8'd106} : s = 292;
	{8'd186,8'd107} : s = 293;
	{8'd186,8'd108} : s = 294;
	{8'd186,8'd109} : s = 295;
	{8'd186,8'd110} : s = 296;
	{8'd186,8'd111} : s = 297;
	{8'd186,8'd112} : s = 298;
	{8'd186,8'd113} : s = 299;
	{8'd186,8'd114} : s = 300;
	{8'd186,8'd115} : s = 301;
	{8'd186,8'd116} : s = 302;
	{8'd186,8'd117} : s = 303;
	{8'd186,8'd118} : s = 304;
	{8'd186,8'd119} : s = 305;
	{8'd186,8'd120} : s = 306;
	{8'd186,8'd121} : s = 307;
	{8'd186,8'd122} : s = 308;
	{8'd186,8'd123} : s = 309;
	{8'd186,8'd124} : s = 310;
	{8'd186,8'd125} : s = 311;
	{8'd186,8'd126} : s = 312;
	{8'd186,8'd127} : s = 313;
	{8'd186,8'd128} : s = 314;
	{8'd186,8'd129} : s = 315;
	{8'd186,8'd130} : s = 316;
	{8'd186,8'd131} : s = 317;
	{8'd186,8'd132} : s = 318;
	{8'd186,8'd133} : s = 319;
	{8'd186,8'd134} : s = 320;
	{8'd186,8'd135} : s = 321;
	{8'd186,8'd136} : s = 322;
	{8'd186,8'd137} : s = 323;
	{8'd186,8'd138} : s = 324;
	{8'd186,8'd139} : s = 325;
	{8'd186,8'd140} : s = 326;
	{8'd186,8'd141} : s = 327;
	{8'd186,8'd142} : s = 328;
	{8'd186,8'd143} : s = 329;
	{8'd186,8'd144} : s = 330;
	{8'd186,8'd145} : s = 331;
	{8'd186,8'd146} : s = 332;
	{8'd186,8'd147} : s = 333;
	{8'd186,8'd148} : s = 334;
	{8'd186,8'd149} : s = 335;
	{8'd186,8'd150} : s = 336;
	{8'd186,8'd151} : s = 337;
	{8'd186,8'd152} : s = 338;
	{8'd186,8'd153} : s = 339;
	{8'd186,8'd154} : s = 340;
	{8'd186,8'd155} : s = 341;
	{8'd186,8'd156} : s = 342;
	{8'd186,8'd157} : s = 343;
	{8'd186,8'd158} : s = 344;
	{8'd186,8'd159} : s = 345;
	{8'd186,8'd160} : s = 346;
	{8'd186,8'd161} : s = 347;
	{8'd186,8'd162} : s = 348;
	{8'd186,8'd163} : s = 349;
	{8'd186,8'd164} : s = 350;
	{8'd186,8'd165} : s = 351;
	{8'd186,8'd166} : s = 352;
	{8'd186,8'd167} : s = 353;
	{8'd186,8'd168} : s = 354;
	{8'd186,8'd169} : s = 355;
	{8'd186,8'd170} : s = 356;
	{8'd186,8'd171} : s = 357;
	{8'd186,8'd172} : s = 358;
	{8'd186,8'd173} : s = 359;
	{8'd186,8'd174} : s = 360;
	{8'd186,8'd175} : s = 361;
	{8'd186,8'd176} : s = 362;
	{8'd186,8'd177} : s = 363;
	{8'd186,8'd178} : s = 364;
	{8'd186,8'd179} : s = 365;
	{8'd186,8'd180} : s = 366;
	{8'd186,8'd181} : s = 367;
	{8'd186,8'd182} : s = 368;
	{8'd186,8'd183} : s = 369;
	{8'd186,8'd184} : s = 370;
	{8'd186,8'd185} : s = 371;
	{8'd186,8'd186} : s = 372;
	{8'd186,8'd187} : s = 373;
	{8'd186,8'd188} : s = 374;
	{8'd186,8'd189} : s = 375;
	{8'd186,8'd190} : s = 376;
	{8'd186,8'd191} : s = 377;
	{8'd186,8'd192} : s = 378;
	{8'd186,8'd193} : s = 379;
	{8'd186,8'd194} : s = 380;
	{8'd186,8'd195} : s = 381;
	{8'd186,8'd196} : s = 382;
	{8'd186,8'd197} : s = 383;
	{8'd186,8'd198} : s = 384;
	{8'd186,8'd199} : s = 385;
	{8'd186,8'd200} : s = 386;
	{8'd186,8'd201} : s = 387;
	{8'd186,8'd202} : s = 388;
	{8'd186,8'd203} : s = 389;
	{8'd186,8'd204} : s = 390;
	{8'd186,8'd205} : s = 391;
	{8'd186,8'd206} : s = 392;
	{8'd186,8'd207} : s = 393;
	{8'd186,8'd208} : s = 394;
	{8'd186,8'd209} : s = 395;
	{8'd186,8'd210} : s = 396;
	{8'd186,8'd211} : s = 397;
	{8'd186,8'd212} : s = 398;
	{8'd186,8'd213} : s = 399;
	{8'd186,8'd214} : s = 400;
	{8'd186,8'd215} : s = 401;
	{8'd186,8'd216} : s = 402;
	{8'd186,8'd217} : s = 403;
	{8'd186,8'd218} : s = 404;
	{8'd186,8'd219} : s = 405;
	{8'd186,8'd220} : s = 406;
	{8'd186,8'd221} : s = 407;
	{8'd186,8'd222} : s = 408;
	{8'd186,8'd223} : s = 409;
	{8'd186,8'd224} : s = 410;
	{8'd186,8'd225} : s = 411;
	{8'd186,8'd226} : s = 412;
	{8'd186,8'd227} : s = 413;
	{8'd186,8'd228} : s = 414;
	{8'd186,8'd229} : s = 415;
	{8'd186,8'd230} : s = 416;
	{8'd186,8'd231} : s = 417;
	{8'd186,8'd232} : s = 418;
	{8'd186,8'd233} : s = 419;
	{8'd186,8'd234} : s = 420;
	{8'd186,8'd235} : s = 421;
	{8'd186,8'd236} : s = 422;
	{8'd186,8'd237} : s = 423;
	{8'd186,8'd238} : s = 424;
	{8'd186,8'd239} : s = 425;
	{8'd186,8'd240} : s = 426;
	{8'd186,8'd241} : s = 427;
	{8'd186,8'd242} : s = 428;
	{8'd186,8'd243} : s = 429;
	{8'd186,8'd244} : s = 430;
	{8'd186,8'd245} : s = 431;
	{8'd186,8'd246} : s = 432;
	{8'd186,8'd247} : s = 433;
	{8'd186,8'd248} : s = 434;
	{8'd186,8'd249} : s = 435;
	{8'd186,8'd250} : s = 436;
	{8'd186,8'd251} : s = 437;
	{8'd186,8'd252} : s = 438;
	{8'd186,8'd253} : s = 439;
	{8'd186,8'd254} : s = 440;
	{8'd186,8'd255} : s = 441;
	{8'd187,8'd0} : s = 187;
	{8'd187,8'd1} : s = 188;
	{8'd187,8'd2} : s = 189;
	{8'd187,8'd3} : s = 190;
	{8'd187,8'd4} : s = 191;
	{8'd187,8'd5} : s = 192;
	{8'd187,8'd6} : s = 193;
	{8'd187,8'd7} : s = 194;
	{8'd187,8'd8} : s = 195;
	{8'd187,8'd9} : s = 196;
	{8'd187,8'd10} : s = 197;
	{8'd187,8'd11} : s = 198;
	{8'd187,8'd12} : s = 199;
	{8'd187,8'd13} : s = 200;
	{8'd187,8'd14} : s = 201;
	{8'd187,8'd15} : s = 202;
	{8'd187,8'd16} : s = 203;
	{8'd187,8'd17} : s = 204;
	{8'd187,8'd18} : s = 205;
	{8'd187,8'd19} : s = 206;
	{8'd187,8'd20} : s = 207;
	{8'd187,8'd21} : s = 208;
	{8'd187,8'd22} : s = 209;
	{8'd187,8'd23} : s = 210;
	{8'd187,8'd24} : s = 211;
	{8'd187,8'd25} : s = 212;
	{8'd187,8'd26} : s = 213;
	{8'd187,8'd27} : s = 214;
	{8'd187,8'd28} : s = 215;
	{8'd187,8'd29} : s = 216;
	{8'd187,8'd30} : s = 217;
	{8'd187,8'd31} : s = 218;
	{8'd187,8'd32} : s = 219;
	{8'd187,8'd33} : s = 220;
	{8'd187,8'd34} : s = 221;
	{8'd187,8'd35} : s = 222;
	{8'd187,8'd36} : s = 223;
	{8'd187,8'd37} : s = 224;
	{8'd187,8'd38} : s = 225;
	{8'd187,8'd39} : s = 226;
	{8'd187,8'd40} : s = 227;
	{8'd187,8'd41} : s = 228;
	{8'd187,8'd42} : s = 229;
	{8'd187,8'd43} : s = 230;
	{8'd187,8'd44} : s = 231;
	{8'd187,8'd45} : s = 232;
	{8'd187,8'd46} : s = 233;
	{8'd187,8'd47} : s = 234;
	{8'd187,8'd48} : s = 235;
	{8'd187,8'd49} : s = 236;
	{8'd187,8'd50} : s = 237;
	{8'd187,8'd51} : s = 238;
	{8'd187,8'd52} : s = 239;
	{8'd187,8'd53} : s = 240;
	{8'd187,8'd54} : s = 241;
	{8'd187,8'd55} : s = 242;
	{8'd187,8'd56} : s = 243;
	{8'd187,8'd57} : s = 244;
	{8'd187,8'd58} : s = 245;
	{8'd187,8'd59} : s = 246;
	{8'd187,8'd60} : s = 247;
	{8'd187,8'd61} : s = 248;
	{8'd187,8'd62} : s = 249;
	{8'd187,8'd63} : s = 250;
	{8'd187,8'd64} : s = 251;
	{8'd187,8'd65} : s = 252;
	{8'd187,8'd66} : s = 253;
	{8'd187,8'd67} : s = 254;
	{8'd187,8'd68} : s = 255;
	{8'd187,8'd69} : s = 256;
	{8'd187,8'd70} : s = 257;
	{8'd187,8'd71} : s = 258;
	{8'd187,8'd72} : s = 259;
	{8'd187,8'd73} : s = 260;
	{8'd187,8'd74} : s = 261;
	{8'd187,8'd75} : s = 262;
	{8'd187,8'd76} : s = 263;
	{8'd187,8'd77} : s = 264;
	{8'd187,8'd78} : s = 265;
	{8'd187,8'd79} : s = 266;
	{8'd187,8'd80} : s = 267;
	{8'd187,8'd81} : s = 268;
	{8'd187,8'd82} : s = 269;
	{8'd187,8'd83} : s = 270;
	{8'd187,8'd84} : s = 271;
	{8'd187,8'd85} : s = 272;
	{8'd187,8'd86} : s = 273;
	{8'd187,8'd87} : s = 274;
	{8'd187,8'd88} : s = 275;
	{8'd187,8'd89} : s = 276;
	{8'd187,8'd90} : s = 277;
	{8'd187,8'd91} : s = 278;
	{8'd187,8'd92} : s = 279;
	{8'd187,8'd93} : s = 280;
	{8'd187,8'd94} : s = 281;
	{8'd187,8'd95} : s = 282;
	{8'd187,8'd96} : s = 283;
	{8'd187,8'd97} : s = 284;
	{8'd187,8'd98} : s = 285;
	{8'd187,8'd99} : s = 286;
	{8'd187,8'd100} : s = 287;
	{8'd187,8'd101} : s = 288;
	{8'd187,8'd102} : s = 289;
	{8'd187,8'd103} : s = 290;
	{8'd187,8'd104} : s = 291;
	{8'd187,8'd105} : s = 292;
	{8'd187,8'd106} : s = 293;
	{8'd187,8'd107} : s = 294;
	{8'd187,8'd108} : s = 295;
	{8'd187,8'd109} : s = 296;
	{8'd187,8'd110} : s = 297;
	{8'd187,8'd111} : s = 298;
	{8'd187,8'd112} : s = 299;
	{8'd187,8'd113} : s = 300;
	{8'd187,8'd114} : s = 301;
	{8'd187,8'd115} : s = 302;
	{8'd187,8'd116} : s = 303;
	{8'd187,8'd117} : s = 304;
	{8'd187,8'd118} : s = 305;
	{8'd187,8'd119} : s = 306;
	{8'd187,8'd120} : s = 307;
	{8'd187,8'd121} : s = 308;
	{8'd187,8'd122} : s = 309;
	{8'd187,8'd123} : s = 310;
	{8'd187,8'd124} : s = 311;
	{8'd187,8'd125} : s = 312;
	{8'd187,8'd126} : s = 313;
	{8'd187,8'd127} : s = 314;
	{8'd187,8'd128} : s = 315;
	{8'd187,8'd129} : s = 316;
	{8'd187,8'd130} : s = 317;
	{8'd187,8'd131} : s = 318;
	{8'd187,8'd132} : s = 319;
	{8'd187,8'd133} : s = 320;
	{8'd187,8'd134} : s = 321;
	{8'd187,8'd135} : s = 322;
	{8'd187,8'd136} : s = 323;
	{8'd187,8'd137} : s = 324;
	{8'd187,8'd138} : s = 325;
	{8'd187,8'd139} : s = 326;
	{8'd187,8'd140} : s = 327;
	{8'd187,8'd141} : s = 328;
	{8'd187,8'd142} : s = 329;
	{8'd187,8'd143} : s = 330;
	{8'd187,8'd144} : s = 331;
	{8'd187,8'd145} : s = 332;
	{8'd187,8'd146} : s = 333;
	{8'd187,8'd147} : s = 334;
	{8'd187,8'd148} : s = 335;
	{8'd187,8'd149} : s = 336;
	{8'd187,8'd150} : s = 337;
	{8'd187,8'd151} : s = 338;
	{8'd187,8'd152} : s = 339;
	{8'd187,8'd153} : s = 340;
	{8'd187,8'd154} : s = 341;
	{8'd187,8'd155} : s = 342;
	{8'd187,8'd156} : s = 343;
	{8'd187,8'd157} : s = 344;
	{8'd187,8'd158} : s = 345;
	{8'd187,8'd159} : s = 346;
	{8'd187,8'd160} : s = 347;
	{8'd187,8'd161} : s = 348;
	{8'd187,8'd162} : s = 349;
	{8'd187,8'd163} : s = 350;
	{8'd187,8'd164} : s = 351;
	{8'd187,8'd165} : s = 352;
	{8'd187,8'd166} : s = 353;
	{8'd187,8'd167} : s = 354;
	{8'd187,8'd168} : s = 355;
	{8'd187,8'd169} : s = 356;
	{8'd187,8'd170} : s = 357;
	{8'd187,8'd171} : s = 358;
	{8'd187,8'd172} : s = 359;
	{8'd187,8'd173} : s = 360;
	{8'd187,8'd174} : s = 361;
	{8'd187,8'd175} : s = 362;
	{8'd187,8'd176} : s = 363;
	{8'd187,8'd177} : s = 364;
	{8'd187,8'd178} : s = 365;
	{8'd187,8'd179} : s = 366;
	{8'd187,8'd180} : s = 367;
	{8'd187,8'd181} : s = 368;
	{8'd187,8'd182} : s = 369;
	{8'd187,8'd183} : s = 370;
	{8'd187,8'd184} : s = 371;
	{8'd187,8'd185} : s = 372;
	{8'd187,8'd186} : s = 373;
	{8'd187,8'd187} : s = 374;
	{8'd187,8'd188} : s = 375;
	{8'd187,8'd189} : s = 376;
	{8'd187,8'd190} : s = 377;
	{8'd187,8'd191} : s = 378;
	{8'd187,8'd192} : s = 379;
	{8'd187,8'd193} : s = 380;
	{8'd187,8'd194} : s = 381;
	{8'd187,8'd195} : s = 382;
	{8'd187,8'd196} : s = 383;
	{8'd187,8'd197} : s = 384;
	{8'd187,8'd198} : s = 385;
	{8'd187,8'd199} : s = 386;
	{8'd187,8'd200} : s = 387;
	{8'd187,8'd201} : s = 388;
	{8'd187,8'd202} : s = 389;
	{8'd187,8'd203} : s = 390;
	{8'd187,8'd204} : s = 391;
	{8'd187,8'd205} : s = 392;
	{8'd187,8'd206} : s = 393;
	{8'd187,8'd207} : s = 394;
	{8'd187,8'd208} : s = 395;
	{8'd187,8'd209} : s = 396;
	{8'd187,8'd210} : s = 397;
	{8'd187,8'd211} : s = 398;
	{8'd187,8'd212} : s = 399;
	{8'd187,8'd213} : s = 400;
	{8'd187,8'd214} : s = 401;
	{8'd187,8'd215} : s = 402;
	{8'd187,8'd216} : s = 403;
	{8'd187,8'd217} : s = 404;
	{8'd187,8'd218} : s = 405;
	{8'd187,8'd219} : s = 406;
	{8'd187,8'd220} : s = 407;
	{8'd187,8'd221} : s = 408;
	{8'd187,8'd222} : s = 409;
	{8'd187,8'd223} : s = 410;
	{8'd187,8'd224} : s = 411;
	{8'd187,8'd225} : s = 412;
	{8'd187,8'd226} : s = 413;
	{8'd187,8'd227} : s = 414;
	{8'd187,8'd228} : s = 415;
	{8'd187,8'd229} : s = 416;
	{8'd187,8'd230} : s = 417;
	{8'd187,8'd231} : s = 418;
	{8'd187,8'd232} : s = 419;
	{8'd187,8'd233} : s = 420;
	{8'd187,8'd234} : s = 421;
	{8'd187,8'd235} : s = 422;
	{8'd187,8'd236} : s = 423;
	{8'd187,8'd237} : s = 424;
	{8'd187,8'd238} : s = 425;
	{8'd187,8'd239} : s = 426;
	{8'd187,8'd240} : s = 427;
	{8'd187,8'd241} : s = 428;
	{8'd187,8'd242} : s = 429;
	{8'd187,8'd243} : s = 430;
	{8'd187,8'd244} : s = 431;
	{8'd187,8'd245} : s = 432;
	{8'd187,8'd246} : s = 433;
	{8'd187,8'd247} : s = 434;
	{8'd187,8'd248} : s = 435;
	{8'd187,8'd249} : s = 436;
	{8'd187,8'd250} : s = 437;
	{8'd187,8'd251} : s = 438;
	{8'd187,8'd252} : s = 439;
	{8'd187,8'd253} : s = 440;
	{8'd187,8'd254} : s = 441;
	{8'd187,8'd255} : s = 442;
	{8'd188,8'd0} : s = 188;
	{8'd188,8'd1} : s = 189;
	{8'd188,8'd2} : s = 190;
	{8'd188,8'd3} : s = 191;
	{8'd188,8'd4} : s = 192;
	{8'd188,8'd5} : s = 193;
	{8'd188,8'd6} : s = 194;
	{8'd188,8'd7} : s = 195;
	{8'd188,8'd8} : s = 196;
	{8'd188,8'd9} : s = 197;
	{8'd188,8'd10} : s = 198;
	{8'd188,8'd11} : s = 199;
	{8'd188,8'd12} : s = 200;
	{8'd188,8'd13} : s = 201;
	{8'd188,8'd14} : s = 202;
	{8'd188,8'd15} : s = 203;
	{8'd188,8'd16} : s = 204;
	{8'd188,8'd17} : s = 205;
	{8'd188,8'd18} : s = 206;
	{8'd188,8'd19} : s = 207;
	{8'd188,8'd20} : s = 208;
	{8'd188,8'd21} : s = 209;
	{8'd188,8'd22} : s = 210;
	{8'd188,8'd23} : s = 211;
	{8'd188,8'd24} : s = 212;
	{8'd188,8'd25} : s = 213;
	{8'd188,8'd26} : s = 214;
	{8'd188,8'd27} : s = 215;
	{8'd188,8'd28} : s = 216;
	{8'd188,8'd29} : s = 217;
	{8'd188,8'd30} : s = 218;
	{8'd188,8'd31} : s = 219;
	{8'd188,8'd32} : s = 220;
	{8'd188,8'd33} : s = 221;
	{8'd188,8'd34} : s = 222;
	{8'd188,8'd35} : s = 223;
	{8'd188,8'd36} : s = 224;
	{8'd188,8'd37} : s = 225;
	{8'd188,8'd38} : s = 226;
	{8'd188,8'd39} : s = 227;
	{8'd188,8'd40} : s = 228;
	{8'd188,8'd41} : s = 229;
	{8'd188,8'd42} : s = 230;
	{8'd188,8'd43} : s = 231;
	{8'd188,8'd44} : s = 232;
	{8'd188,8'd45} : s = 233;
	{8'd188,8'd46} : s = 234;
	{8'd188,8'd47} : s = 235;
	{8'd188,8'd48} : s = 236;
	{8'd188,8'd49} : s = 237;
	{8'd188,8'd50} : s = 238;
	{8'd188,8'd51} : s = 239;
	{8'd188,8'd52} : s = 240;
	{8'd188,8'd53} : s = 241;
	{8'd188,8'd54} : s = 242;
	{8'd188,8'd55} : s = 243;
	{8'd188,8'd56} : s = 244;
	{8'd188,8'd57} : s = 245;
	{8'd188,8'd58} : s = 246;
	{8'd188,8'd59} : s = 247;
	{8'd188,8'd60} : s = 248;
	{8'd188,8'd61} : s = 249;
	{8'd188,8'd62} : s = 250;
	{8'd188,8'd63} : s = 251;
	{8'd188,8'd64} : s = 252;
	{8'd188,8'd65} : s = 253;
	{8'd188,8'd66} : s = 254;
	{8'd188,8'd67} : s = 255;
	{8'd188,8'd68} : s = 256;
	{8'd188,8'd69} : s = 257;
	{8'd188,8'd70} : s = 258;
	{8'd188,8'd71} : s = 259;
	{8'd188,8'd72} : s = 260;
	{8'd188,8'd73} : s = 261;
	{8'd188,8'd74} : s = 262;
	{8'd188,8'd75} : s = 263;
	{8'd188,8'd76} : s = 264;
	{8'd188,8'd77} : s = 265;
	{8'd188,8'd78} : s = 266;
	{8'd188,8'd79} : s = 267;
	{8'd188,8'd80} : s = 268;
	{8'd188,8'd81} : s = 269;
	{8'd188,8'd82} : s = 270;
	{8'd188,8'd83} : s = 271;
	{8'd188,8'd84} : s = 272;
	{8'd188,8'd85} : s = 273;
	{8'd188,8'd86} : s = 274;
	{8'd188,8'd87} : s = 275;
	{8'd188,8'd88} : s = 276;
	{8'd188,8'd89} : s = 277;
	{8'd188,8'd90} : s = 278;
	{8'd188,8'd91} : s = 279;
	{8'd188,8'd92} : s = 280;
	{8'd188,8'd93} : s = 281;
	{8'd188,8'd94} : s = 282;
	{8'd188,8'd95} : s = 283;
	{8'd188,8'd96} : s = 284;
	{8'd188,8'd97} : s = 285;
	{8'd188,8'd98} : s = 286;
	{8'd188,8'd99} : s = 287;
	{8'd188,8'd100} : s = 288;
	{8'd188,8'd101} : s = 289;
	{8'd188,8'd102} : s = 290;
	{8'd188,8'd103} : s = 291;
	{8'd188,8'd104} : s = 292;
	{8'd188,8'd105} : s = 293;
	{8'd188,8'd106} : s = 294;
	{8'd188,8'd107} : s = 295;
	{8'd188,8'd108} : s = 296;
	{8'd188,8'd109} : s = 297;
	{8'd188,8'd110} : s = 298;
	{8'd188,8'd111} : s = 299;
	{8'd188,8'd112} : s = 300;
	{8'd188,8'd113} : s = 301;
	{8'd188,8'd114} : s = 302;
	{8'd188,8'd115} : s = 303;
	{8'd188,8'd116} : s = 304;
	{8'd188,8'd117} : s = 305;
	{8'd188,8'd118} : s = 306;
	{8'd188,8'd119} : s = 307;
	{8'd188,8'd120} : s = 308;
	{8'd188,8'd121} : s = 309;
	{8'd188,8'd122} : s = 310;
	{8'd188,8'd123} : s = 311;
	{8'd188,8'd124} : s = 312;
	{8'd188,8'd125} : s = 313;
	{8'd188,8'd126} : s = 314;
	{8'd188,8'd127} : s = 315;
	{8'd188,8'd128} : s = 316;
	{8'd188,8'd129} : s = 317;
	{8'd188,8'd130} : s = 318;
	{8'd188,8'd131} : s = 319;
	{8'd188,8'd132} : s = 320;
	{8'd188,8'd133} : s = 321;
	{8'd188,8'd134} : s = 322;
	{8'd188,8'd135} : s = 323;
	{8'd188,8'd136} : s = 324;
	{8'd188,8'd137} : s = 325;
	{8'd188,8'd138} : s = 326;
	{8'd188,8'd139} : s = 327;
	{8'd188,8'd140} : s = 328;
	{8'd188,8'd141} : s = 329;
	{8'd188,8'd142} : s = 330;
	{8'd188,8'd143} : s = 331;
	{8'd188,8'd144} : s = 332;
	{8'd188,8'd145} : s = 333;
	{8'd188,8'd146} : s = 334;
	{8'd188,8'd147} : s = 335;
	{8'd188,8'd148} : s = 336;
	{8'd188,8'd149} : s = 337;
	{8'd188,8'd150} : s = 338;
	{8'd188,8'd151} : s = 339;
	{8'd188,8'd152} : s = 340;
	{8'd188,8'd153} : s = 341;
	{8'd188,8'd154} : s = 342;
	{8'd188,8'd155} : s = 343;
	{8'd188,8'd156} : s = 344;
	{8'd188,8'd157} : s = 345;
	{8'd188,8'd158} : s = 346;
	{8'd188,8'd159} : s = 347;
	{8'd188,8'd160} : s = 348;
	{8'd188,8'd161} : s = 349;
	{8'd188,8'd162} : s = 350;
	{8'd188,8'd163} : s = 351;
	{8'd188,8'd164} : s = 352;
	{8'd188,8'd165} : s = 353;
	{8'd188,8'd166} : s = 354;
	{8'd188,8'd167} : s = 355;
	{8'd188,8'd168} : s = 356;
	{8'd188,8'd169} : s = 357;
	{8'd188,8'd170} : s = 358;
	{8'd188,8'd171} : s = 359;
	{8'd188,8'd172} : s = 360;
	{8'd188,8'd173} : s = 361;
	{8'd188,8'd174} : s = 362;
	{8'd188,8'd175} : s = 363;
	{8'd188,8'd176} : s = 364;
	{8'd188,8'd177} : s = 365;
	{8'd188,8'd178} : s = 366;
	{8'd188,8'd179} : s = 367;
	{8'd188,8'd180} : s = 368;
	{8'd188,8'd181} : s = 369;
	{8'd188,8'd182} : s = 370;
	{8'd188,8'd183} : s = 371;
	{8'd188,8'd184} : s = 372;
	{8'd188,8'd185} : s = 373;
	{8'd188,8'd186} : s = 374;
	{8'd188,8'd187} : s = 375;
	{8'd188,8'd188} : s = 376;
	{8'd188,8'd189} : s = 377;
	{8'd188,8'd190} : s = 378;
	{8'd188,8'd191} : s = 379;
	{8'd188,8'd192} : s = 380;
	{8'd188,8'd193} : s = 381;
	{8'd188,8'd194} : s = 382;
	{8'd188,8'd195} : s = 383;
	{8'd188,8'd196} : s = 384;
	{8'd188,8'd197} : s = 385;
	{8'd188,8'd198} : s = 386;
	{8'd188,8'd199} : s = 387;
	{8'd188,8'd200} : s = 388;
	{8'd188,8'd201} : s = 389;
	{8'd188,8'd202} : s = 390;
	{8'd188,8'd203} : s = 391;
	{8'd188,8'd204} : s = 392;
	{8'd188,8'd205} : s = 393;
	{8'd188,8'd206} : s = 394;
	{8'd188,8'd207} : s = 395;
	{8'd188,8'd208} : s = 396;
	{8'd188,8'd209} : s = 397;
	{8'd188,8'd210} : s = 398;
	{8'd188,8'd211} : s = 399;
	{8'd188,8'd212} : s = 400;
	{8'd188,8'd213} : s = 401;
	{8'd188,8'd214} : s = 402;
	{8'd188,8'd215} : s = 403;
	{8'd188,8'd216} : s = 404;
	{8'd188,8'd217} : s = 405;
	{8'd188,8'd218} : s = 406;
	{8'd188,8'd219} : s = 407;
	{8'd188,8'd220} : s = 408;
	{8'd188,8'd221} : s = 409;
	{8'd188,8'd222} : s = 410;
	{8'd188,8'd223} : s = 411;
	{8'd188,8'd224} : s = 412;
	{8'd188,8'd225} : s = 413;
	{8'd188,8'd226} : s = 414;
	{8'd188,8'd227} : s = 415;
	{8'd188,8'd228} : s = 416;
	{8'd188,8'd229} : s = 417;
	{8'd188,8'd230} : s = 418;
	{8'd188,8'd231} : s = 419;
	{8'd188,8'd232} : s = 420;
	{8'd188,8'd233} : s = 421;
	{8'd188,8'd234} : s = 422;
	{8'd188,8'd235} : s = 423;
	{8'd188,8'd236} : s = 424;
	{8'd188,8'd237} : s = 425;
	{8'd188,8'd238} : s = 426;
	{8'd188,8'd239} : s = 427;
	{8'd188,8'd240} : s = 428;
	{8'd188,8'd241} : s = 429;
	{8'd188,8'd242} : s = 430;
	{8'd188,8'd243} : s = 431;
	{8'd188,8'd244} : s = 432;
	{8'd188,8'd245} : s = 433;
	{8'd188,8'd246} : s = 434;
	{8'd188,8'd247} : s = 435;
	{8'd188,8'd248} : s = 436;
	{8'd188,8'd249} : s = 437;
	{8'd188,8'd250} : s = 438;
	{8'd188,8'd251} : s = 439;
	{8'd188,8'd252} : s = 440;
	{8'd188,8'd253} : s = 441;
	{8'd188,8'd254} : s = 442;
	{8'd188,8'd255} : s = 443;
	{8'd189,8'd0} : s = 189;
	{8'd189,8'd1} : s = 190;
	{8'd189,8'd2} : s = 191;
	{8'd189,8'd3} : s = 192;
	{8'd189,8'd4} : s = 193;
	{8'd189,8'd5} : s = 194;
	{8'd189,8'd6} : s = 195;
	{8'd189,8'd7} : s = 196;
	{8'd189,8'd8} : s = 197;
	{8'd189,8'd9} : s = 198;
	{8'd189,8'd10} : s = 199;
	{8'd189,8'd11} : s = 200;
	{8'd189,8'd12} : s = 201;
	{8'd189,8'd13} : s = 202;
	{8'd189,8'd14} : s = 203;
	{8'd189,8'd15} : s = 204;
	{8'd189,8'd16} : s = 205;
	{8'd189,8'd17} : s = 206;
	{8'd189,8'd18} : s = 207;
	{8'd189,8'd19} : s = 208;
	{8'd189,8'd20} : s = 209;
	{8'd189,8'd21} : s = 210;
	{8'd189,8'd22} : s = 211;
	{8'd189,8'd23} : s = 212;
	{8'd189,8'd24} : s = 213;
	{8'd189,8'd25} : s = 214;
	{8'd189,8'd26} : s = 215;
	{8'd189,8'd27} : s = 216;
	{8'd189,8'd28} : s = 217;
	{8'd189,8'd29} : s = 218;
	{8'd189,8'd30} : s = 219;
	{8'd189,8'd31} : s = 220;
	{8'd189,8'd32} : s = 221;
	{8'd189,8'd33} : s = 222;
	{8'd189,8'd34} : s = 223;
	{8'd189,8'd35} : s = 224;
	{8'd189,8'd36} : s = 225;
	{8'd189,8'd37} : s = 226;
	{8'd189,8'd38} : s = 227;
	{8'd189,8'd39} : s = 228;
	{8'd189,8'd40} : s = 229;
	{8'd189,8'd41} : s = 230;
	{8'd189,8'd42} : s = 231;
	{8'd189,8'd43} : s = 232;
	{8'd189,8'd44} : s = 233;
	{8'd189,8'd45} : s = 234;
	{8'd189,8'd46} : s = 235;
	{8'd189,8'd47} : s = 236;
	{8'd189,8'd48} : s = 237;
	{8'd189,8'd49} : s = 238;
	{8'd189,8'd50} : s = 239;
	{8'd189,8'd51} : s = 240;
	{8'd189,8'd52} : s = 241;
	{8'd189,8'd53} : s = 242;
	{8'd189,8'd54} : s = 243;
	{8'd189,8'd55} : s = 244;
	{8'd189,8'd56} : s = 245;
	{8'd189,8'd57} : s = 246;
	{8'd189,8'd58} : s = 247;
	{8'd189,8'd59} : s = 248;
	{8'd189,8'd60} : s = 249;
	{8'd189,8'd61} : s = 250;
	{8'd189,8'd62} : s = 251;
	{8'd189,8'd63} : s = 252;
	{8'd189,8'd64} : s = 253;
	{8'd189,8'd65} : s = 254;
	{8'd189,8'd66} : s = 255;
	{8'd189,8'd67} : s = 256;
	{8'd189,8'd68} : s = 257;
	{8'd189,8'd69} : s = 258;
	{8'd189,8'd70} : s = 259;
	{8'd189,8'd71} : s = 260;
	{8'd189,8'd72} : s = 261;
	{8'd189,8'd73} : s = 262;
	{8'd189,8'd74} : s = 263;
	{8'd189,8'd75} : s = 264;
	{8'd189,8'd76} : s = 265;
	{8'd189,8'd77} : s = 266;
	{8'd189,8'd78} : s = 267;
	{8'd189,8'd79} : s = 268;
	{8'd189,8'd80} : s = 269;
	{8'd189,8'd81} : s = 270;
	{8'd189,8'd82} : s = 271;
	{8'd189,8'd83} : s = 272;
	{8'd189,8'd84} : s = 273;
	{8'd189,8'd85} : s = 274;
	{8'd189,8'd86} : s = 275;
	{8'd189,8'd87} : s = 276;
	{8'd189,8'd88} : s = 277;
	{8'd189,8'd89} : s = 278;
	{8'd189,8'd90} : s = 279;
	{8'd189,8'd91} : s = 280;
	{8'd189,8'd92} : s = 281;
	{8'd189,8'd93} : s = 282;
	{8'd189,8'd94} : s = 283;
	{8'd189,8'd95} : s = 284;
	{8'd189,8'd96} : s = 285;
	{8'd189,8'd97} : s = 286;
	{8'd189,8'd98} : s = 287;
	{8'd189,8'd99} : s = 288;
	{8'd189,8'd100} : s = 289;
	{8'd189,8'd101} : s = 290;
	{8'd189,8'd102} : s = 291;
	{8'd189,8'd103} : s = 292;
	{8'd189,8'd104} : s = 293;
	{8'd189,8'd105} : s = 294;
	{8'd189,8'd106} : s = 295;
	{8'd189,8'd107} : s = 296;
	{8'd189,8'd108} : s = 297;
	{8'd189,8'd109} : s = 298;
	{8'd189,8'd110} : s = 299;
	{8'd189,8'd111} : s = 300;
	{8'd189,8'd112} : s = 301;
	{8'd189,8'd113} : s = 302;
	{8'd189,8'd114} : s = 303;
	{8'd189,8'd115} : s = 304;
	{8'd189,8'd116} : s = 305;
	{8'd189,8'd117} : s = 306;
	{8'd189,8'd118} : s = 307;
	{8'd189,8'd119} : s = 308;
	{8'd189,8'd120} : s = 309;
	{8'd189,8'd121} : s = 310;
	{8'd189,8'd122} : s = 311;
	{8'd189,8'd123} : s = 312;
	{8'd189,8'd124} : s = 313;
	{8'd189,8'd125} : s = 314;
	{8'd189,8'd126} : s = 315;
	{8'd189,8'd127} : s = 316;
	{8'd189,8'd128} : s = 317;
	{8'd189,8'd129} : s = 318;
	{8'd189,8'd130} : s = 319;
	{8'd189,8'd131} : s = 320;
	{8'd189,8'd132} : s = 321;
	{8'd189,8'd133} : s = 322;
	{8'd189,8'd134} : s = 323;
	{8'd189,8'd135} : s = 324;
	{8'd189,8'd136} : s = 325;
	{8'd189,8'd137} : s = 326;
	{8'd189,8'd138} : s = 327;
	{8'd189,8'd139} : s = 328;
	{8'd189,8'd140} : s = 329;
	{8'd189,8'd141} : s = 330;
	{8'd189,8'd142} : s = 331;
	{8'd189,8'd143} : s = 332;
	{8'd189,8'd144} : s = 333;
	{8'd189,8'd145} : s = 334;
	{8'd189,8'd146} : s = 335;
	{8'd189,8'd147} : s = 336;
	{8'd189,8'd148} : s = 337;
	{8'd189,8'd149} : s = 338;
	{8'd189,8'd150} : s = 339;
	{8'd189,8'd151} : s = 340;
	{8'd189,8'd152} : s = 341;
	{8'd189,8'd153} : s = 342;
	{8'd189,8'd154} : s = 343;
	{8'd189,8'd155} : s = 344;
	{8'd189,8'd156} : s = 345;
	{8'd189,8'd157} : s = 346;
	{8'd189,8'd158} : s = 347;
	{8'd189,8'd159} : s = 348;
	{8'd189,8'd160} : s = 349;
	{8'd189,8'd161} : s = 350;
	{8'd189,8'd162} : s = 351;
	{8'd189,8'd163} : s = 352;
	{8'd189,8'd164} : s = 353;
	{8'd189,8'd165} : s = 354;
	{8'd189,8'd166} : s = 355;
	{8'd189,8'd167} : s = 356;
	{8'd189,8'd168} : s = 357;
	{8'd189,8'd169} : s = 358;
	{8'd189,8'd170} : s = 359;
	{8'd189,8'd171} : s = 360;
	{8'd189,8'd172} : s = 361;
	{8'd189,8'd173} : s = 362;
	{8'd189,8'd174} : s = 363;
	{8'd189,8'd175} : s = 364;
	{8'd189,8'd176} : s = 365;
	{8'd189,8'd177} : s = 366;
	{8'd189,8'd178} : s = 367;
	{8'd189,8'd179} : s = 368;
	{8'd189,8'd180} : s = 369;
	{8'd189,8'd181} : s = 370;
	{8'd189,8'd182} : s = 371;
	{8'd189,8'd183} : s = 372;
	{8'd189,8'd184} : s = 373;
	{8'd189,8'd185} : s = 374;
	{8'd189,8'd186} : s = 375;
	{8'd189,8'd187} : s = 376;
	{8'd189,8'd188} : s = 377;
	{8'd189,8'd189} : s = 378;
	{8'd189,8'd190} : s = 379;
	{8'd189,8'd191} : s = 380;
	{8'd189,8'd192} : s = 381;
	{8'd189,8'd193} : s = 382;
	{8'd189,8'd194} : s = 383;
	{8'd189,8'd195} : s = 384;
	{8'd189,8'd196} : s = 385;
	{8'd189,8'd197} : s = 386;
	{8'd189,8'd198} : s = 387;
	{8'd189,8'd199} : s = 388;
	{8'd189,8'd200} : s = 389;
	{8'd189,8'd201} : s = 390;
	{8'd189,8'd202} : s = 391;
	{8'd189,8'd203} : s = 392;
	{8'd189,8'd204} : s = 393;
	{8'd189,8'd205} : s = 394;
	{8'd189,8'd206} : s = 395;
	{8'd189,8'd207} : s = 396;
	{8'd189,8'd208} : s = 397;
	{8'd189,8'd209} : s = 398;
	{8'd189,8'd210} : s = 399;
	{8'd189,8'd211} : s = 400;
	{8'd189,8'd212} : s = 401;
	{8'd189,8'd213} : s = 402;
	{8'd189,8'd214} : s = 403;
	{8'd189,8'd215} : s = 404;
	{8'd189,8'd216} : s = 405;
	{8'd189,8'd217} : s = 406;
	{8'd189,8'd218} : s = 407;
	{8'd189,8'd219} : s = 408;
	{8'd189,8'd220} : s = 409;
	{8'd189,8'd221} : s = 410;
	{8'd189,8'd222} : s = 411;
	{8'd189,8'd223} : s = 412;
	{8'd189,8'd224} : s = 413;
	{8'd189,8'd225} : s = 414;
	{8'd189,8'd226} : s = 415;
	{8'd189,8'd227} : s = 416;
	{8'd189,8'd228} : s = 417;
	{8'd189,8'd229} : s = 418;
	{8'd189,8'd230} : s = 419;
	{8'd189,8'd231} : s = 420;
	{8'd189,8'd232} : s = 421;
	{8'd189,8'd233} : s = 422;
	{8'd189,8'd234} : s = 423;
	{8'd189,8'd235} : s = 424;
	{8'd189,8'd236} : s = 425;
	{8'd189,8'd237} : s = 426;
	{8'd189,8'd238} : s = 427;
	{8'd189,8'd239} : s = 428;
	{8'd189,8'd240} : s = 429;
	{8'd189,8'd241} : s = 430;
	{8'd189,8'd242} : s = 431;
	{8'd189,8'd243} : s = 432;
	{8'd189,8'd244} : s = 433;
	{8'd189,8'd245} : s = 434;
	{8'd189,8'd246} : s = 435;
	{8'd189,8'd247} : s = 436;
	{8'd189,8'd248} : s = 437;
	{8'd189,8'd249} : s = 438;
	{8'd189,8'd250} : s = 439;
	{8'd189,8'd251} : s = 440;
	{8'd189,8'd252} : s = 441;
	{8'd189,8'd253} : s = 442;
	{8'd189,8'd254} : s = 443;
	{8'd189,8'd255} : s = 444;
	{8'd190,8'd0} : s = 190;
	{8'd190,8'd1} : s = 191;
	{8'd190,8'd2} : s = 192;
	{8'd190,8'd3} : s = 193;
	{8'd190,8'd4} : s = 194;
	{8'd190,8'd5} : s = 195;
	{8'd190,8'd6} : s = 196;
	{8'd190,8'd7} : s = 197;
	{8'd190,8'd8} : s = 198;
	{8'd190,8'd9} : s = 199;
	{8'd190,8'd10} : s = 200;
	{8'd190,8'd11} : s = 201;
	{8'd190,8'd12} : s = 202;
	{8'd190,8'd13} : s = 203;
	{8'd190,8'd14} : s = 204;
	{8'd190,8'd15} : s = 205;
	{8'd190,8'd16} : s = 206;
	{8'd190,8'd17} : s = 207;
	{8'd190,8'd18} : s = 208;
	{8'd190,8'd19} : s = 209;
	{8'd190,8'd20} : s = 210;
	{8'd190,8'd21} : s = 211;
	{8'd190,8'd22} : s = 212;
	{8'd190,8'd23} : s = 213;
	{8'd190,8'd24} : s = 214;
	{8'd190,8'd25} : s = 215;
	{8'd190,8'd26} : s = 216;
	{8'd190,8'd27} : s = 217;
	{8'd190,8'd28} : s = 218;
	{8'd190,8'd29} : s = 219;
	{8'd190,8'd30} : s = 220;
	{8'd190,8'd31} : s = 221;
	{8'd190,8'd32} : s = 222;
	{8'd190,8'd33} : s = 223;
	{8'd190,8'd34} : s = 224;
	{8'd190,8'd35} : s = 225;
	{8'd190,8'd36} : s = 226;
	{8'd190,8'd37} : s = 227;
	{8'd190,8'd38} : s = 228;
	{8'd190,8'd39} : s = 229;
	{8'd190,8'd40} : s = 230;
	{8'd190,8'd41} : s = 231;
	{8'd190,8'd42} : s = 232;
	{8'd190,8'd43} : s = 233;
	{8'd190,8'd44} : s = 234;
	{8'd190,8'd45} : s = 235;
	{8'd190,8'd46} : s = 236;
	{8'd190,8'd47} : s = 237;
	{8'd190,8'd48} : s = 238;
	{8'd190,8'd49} : s = 239;
	{8'd190,8'd50} : s = 240;
	{8'd190,8'd51} : s = 241;
	{8'd190,8'd52} : s = 242;
	{8'd190,8'd53} : s = 243;
	{8'd190,8'd54} : s = 244;
	{8'd190,8'd55} : s = 245;
	{8'd190,8'd56} : s = 246;
	{8'd190,8'd57} : s = 247;
	{8'd190,8'd58} : s = 248;
	{8'd190,8'd59} : s = 249;
	{8'd190,8'd60} : s = 250;
	{8'd190,8'd61} : s = 251;
	{8'd190,8'd62} : s = 252;
	{8'd190,8'd63} : s = 253;
	{8'd190,8'd64} : s = 254;
	{8'd190,8'd65} : s = 255;
	{8'd190,8'd66} : s = 256;
	{8'd190,8'd67} : s = 257;
	{8'd190,8'd68} : s = 258;
	{8'd190,8'd69} : s = 259;
	{8'd190,8'd70} : s = 260;
	{8'd190,8'd71} : s = 261;
	{8'd190,8'd72} : s = 262;
	{8'd190,8'd73} : s = 263;
	{8'd190,8'd74} : s = 264;
	{8'd190,8'd75} : s = 265;
	{8'd190,8'd76} : s = 266;
	{8'd190,8'd77} : s = 267;
	{8'd190,8'd78} : s = 268;
	{8'd190,8'd79} : s = 269;
	{8'd190,8'd80} : s = 270;
	{8'd190,8'd81} : s = 271;
	{8'd190,8'd82} : s = 272;
	{8'd190,8'd83} : s = 273;
	{8'd190,8'd84} : s = 274;
	{8'd190,8'd85} : s = 275;
	{8'd190,8'd86} : s = 276;
	{8'd190,8'd87} : s = 277;
	{8'd190,8'd88} : s = 278;
	{8'd190,8'd89} : s = 279;
	{8'd190,8'd90} : s = 280;
	{8'd190,8'd91} : s = 281;
	{8'd190,8'd92} : s = 282;
	{8'd190,8'd93} : s = 283;
	{8'd190,8'd94} : s = 284;
	{8'd190,8'd95} : s = 285;
	{8'd190,8'd96} : s = 286;
	{8'd190,8'd97} : s = 287;
	{8'd190,8'd98} : s = 288;
	{8'd190,8'd99} : s = 289;
	{8'd190,8'd100} : s = 290;
	{8'd190,8'd101} : s = 291;
	{8'd190,8'd102} : s = 292;
	{8'd190,8'd103} : s = 293;
	{8'd190,8'd104} : s = 294;
	{8'd190,8'd105} : s = 295;
	{8'd190,8'd106} : s = 296;
	{8'd190,8'd107} : s = 297;
	{8'd190,8'd108} : s = 298;
	{8'd190,8'd109} : s = 299;
	{8'd190,8'd110} : s = 300;
	{8'd190,8'd111} : s = 301;
	{8'd190,8'd112} : s = 302;
	{8'd190,8'd113} : s = 303;
	{8'd190,8'd114} : s = 304;
	{8'd190,8'd115} : s = 305;
	{8'd190,8'd116} : s = 306;
	{8'd190,8'd117} : s = 307;
	{8'd190,8'd118} : s = 308;
	{8'd190,8'd119} : s = 309;
	{8'd190,8'd120} : s = 310;
	{8'd190,8'd121} : s = 311;
	{8'd190,8'd122} : s = 312;
	{8'd190,8'd123} : s = 313;
	{8'd190,8'd124} : s = 314;
	{8'd190,8'd125} : s = 315;
	{8'd190,8'd126} : s = 316;
	{8'd190,8'd127} : s = 317;
	{8'd190,8'd128} : s = 318;
	{8'd190,8'd129} : s = 319;
	{8'd190,8'd130} : s = 320;
	{8'd190,8'd131} : s = 321;
	{8'd190,8'd132} : s = 322;
	{8'd190,8'd133} : s = 323;
	{8'd190,8'd134} : s = 324;
	{8'd190,8'd135} : s = 325;
	{8'd190,8'd136} : s = 326;
	{8'd190,8'd137} : s = 327;
	{8'd190,8'd138} : s = 328;
	{8'd190,8'd139} : s = 329;
	{8'd190,8'd140} : s = 330;
	{8'd190,8'd141} : s = 331;
	{8'd190,8'd142} : s = 332;
	{8'd190,8'd143} : s = 333;
	{8'd190,8'd144} : s = 334;
	{8'd190,8'd145} : s = 335;
	{8'd190,8'd146} : s = 336;
	{8'd190,8'd147} : s = 337;
	{8'd190,8'd148} : s = 338;
	{8'd190,8'd149} : s = 339;
	{8'd190,8'd150} : s = 340;
	{8'd190,8'd151} : s = 341;
	{8'd190,8'd152} : s = 342;
	{8'd190,8'd153} : s = 343;
	{8'd190,8'd154} : s = 344;
	{8'd190,8'd155} : s = 345;
	{8'd190,8'd156} : s = 346;
	{8'd190,8'd157} : s = 347;
	{8'd190,8'd158} : s = 348;
	{8'd190,8'd159} : s = 349;
	{8'd190,8'd160} : s = 350;
	{8'd190,8'd161} : s = 351;
	{8'd190,8'd162} : s = 352;
	{8'd190,8'd163} : s = 353;
	{8'd190,8'd164} : s = 354;
	{8'd190,8'd165} : s = 355;
	{8'd190,8'd166} : s = 356;
	{8'd190,8'd167} : s = 357;
	{8'd190,8'd168} : s = 358;
	{8'd190,8'd169} : s = 359;
	{8'd190,8'd170} : s = 360;
	{8'd190,8'd171} : s = 361;
	{8'd190,8'd172} : s = 362;
	{8'd190,8'd173} : s = 363;
	{8'd190,8'd174} : s = 364;
	{8'd190,8'd175} : s = 365;
	{8'd190,8'd176} : s = 366;
	{8'd190,8'd177} : s = 367;
	{8'd190,8'd178} : s = 368;
	{8'd190,8'd179} : s = 369;
	{8'd190,8'd180} : s = 370;
	{8'd190,8'd181} : s = 371;
	{8'd190,8'd182} : s = 372;
	{8'd190,8'd183} : s = 373;
	{8'd190,8'd184} : s = 374;
	{8'd190,8'd185} : s = 375;
	{8'd190,8'd186} : s = 376;
	{8'd190,8'd187} : s = 377;
	{8'd190,8'd188} : s = 378;
	{8'd190,8'd189} : s = 379;
	{8'd190,8'd190} : s = 380;
	{8'd190,8'd191} : s = 381;
	{8'd190,8'd192} : s = 382;
	{8'd190,8'd193} : s = 383;
	{8'd190,8'd194} : s = 384;
	{8'd190,8'd195} : s = 385;
	{8'd190,8'd196} : s = 386;
	{8'd190,8'd197} : s = 387;
	{8'd190,8'd198} : s = 388;
	{8'd190,8'd199} : s = 389;
	{8'd190,8'd200} : s = 390;
	{8'd190,8'd201} : s = 391;
	{8'd190,8'd202} : s = 392;
	{8'd190,8'd203} : s = 393;
	{8'd190,8'd204} : s = 394;
	{8'd190,8'd205} : s = 395;
	{8'd190,8'd206} : s = 396;
	{8'd190,8'd207} : s = 397;
	{8'd190,8'd208} : s = 398;
	{8'd190,8'd209} : s = 399;
	{8'd190,8'd210} : s = 400;
	{8'd190,8'd211} : s = 401;
	{8'd190,8'd212} : s = 402;
	{8'd190,8'd213} : s = 403;
	{8'd190,8'd214} : s = 404;
	{8'd190,8'd215} : s = 405;
	{8'd190,8'd216} : s = 406;
	{8'd190,8'd217} : s = 407;
	{8'd190,8'd218} : s = 408;
	{8'd190,8'd219} : s = 409;
	{8'd190,8'd220} : s = 410;
	{8'd190,8'd221} : s = 411;
	{8'd190,8'd222} : s = 412;
	{8'd190,8'd223} : s = 413;
	{8'd190,8'd224} : s = 414;
	{8'd190,8'd225} : s = 415;
	{8'd190,8'd226} : s = 416;
	{8'd190,8'd227} : s = 417;
	{8'd190,8'd228} : s = 418;
	{8'd190,8'd229} : s = 419;
	{8'd190,8'd230} : s = 420;
	{8'd190,8'd231} : s = 421;
	{8'd190,8'd232} : s = 422;
	{8'd190,8'd233} : s = 423;
	{8'd190,8'd234} : s = 424;
	{8'd190,8'd235} : s = 425;
	{8'd190,8'd236} : s = 426;
	{8'd190,8'd237} : s = 427;
	{8'd190,8'd238} : s = 428;
	{8'd190,8'd239} : s = 429;
	{8'd190,8'd240} : s = 430;
	{8'd190,8'd241} : s = 431;
	{8'd190,8'd242} : s = 432;
	{8'd190,8'd243} : s = 433;
	{8'd190,8'd244} : s = 434;
	{8'd190,8'd245} : s = 435;
	{8'd190,8'd246} : s = 436;
	{8'd190,8'd247} : s = 437;
	{8'd190,8'd248} : s = 438;
	{8'd190,8'd249} : s = 439;
	{8'd190,8'd250} : s = 440;
	{8'd190,8'd251} : s = 441;
	{8'd190,8'd252} : s = 442;
	{8'd190,8'd253} : s = 443;
	{8'd190,8'd254} : s = 444;
	{8'd190,8'd255} : s = 445;
	{8'd191,8'd0} : s = 191;
	{8'd191,8'd1} : s = 192;
	{8'd191,8'd2} : s = 193;
	{8'd191,8'd3} : s = 194;
	{8'd191,8'd4} : s = 195;
	{8'd191,8'd5} : s = 196;
	{8'd191,8'd6} : s = 197;
	{8'd191,8'd7} : s = 198;
	{8'd191,8'd8} : s = 199;
	{8'd191,8'd9} : s = 200;
	{8'd191,8'd10} : s = 201;
	{8'd191,8'd11} : s = 202;
	{8'd191,8'd12} : s = 203;
	{8'd191,8'd13} : s = 204;
	{8'd191,8'd14} : s = 205;
	{8'd191,8'd15} : s = 206;
	{8'd191,8'd16} : s = 207;
	{8'd191,8'd17} : s = 208;
	{8'd191,8'd18} : s = 209;
	{8'd191,8'd19} : s = 210;
	{8'd191,8'd20} : s = 211;
	{8'd191,8'd21} : s = 212;
	{8'd191,8'd22} : s = 213;
	{8'd191,8'd23} : s = 214;
	{8'd191,8'd24} : s = 215;
	{8'd191,8'd25} : s = 216;
	{8'd191,8'd26} : s = 217;
	{8'd191,8'd27} : s = 218;
	{8'd191,8'd28} : s = 219;
	{8'd191,8'd29} : s = 220;
	{8'd191,8'd30} : s = 221;
	{8'd191,8'd31} : s = 222;
	{8'd191,8'd32} : s = 223;
	{8'd191,8'd33} : s = 224;
	{8'd191,8'd34} : s = 225;
	{8'd191,8'd35} : s = 226;
	{8'd191,8'd36} : s = 227;
	{8'd191,8'd37} : s = 228;
	{8'd191,8'd38} : s = 229;
	{8'd191,8'd39} : s = 230;
	{8'd191,8'd40} : s = 231;
	{8'd191,8'd41} : s = 232;
	{8'd191,8'd42} : s = 233;
	{8'd191,8'd43} : s = 234;
	{8'd191,8'd44} : s = 235;
	{8'd191,8'd45} : s = 236;
	{8'd191,8'd46} : s = 237;
	{8'd191,8'd47} : s = 238;
	{8'd191,8'd48} : s = 239;
	{8'd191,8'd49} : s = 240;
	{8'd191,8'd50} : s = 241;
	{8'd191,8'd51} : s = 242;
	{8'd191,8'd52} : s = 243;
	{8'd191,8'd53} : s = 244;
	{8'd191,8'd54} : s = 245;
	{8'd191,8'd55} : s = 246;
	{8'd191,8'd56} : s = 247;
	{8'd191,8'd57} : s = 248;
	{8'd191,8'd58} : s = 249;
	{8'd191,8'd59} : s = 250;
	{8'd191,8'd60} : s = 251;
	{8'd191,8'd61} : s = 252;
	{8'd191,8'd62} : s = 253;
	{8'd191,8'd63} : s = 254;
	{8'd191,8'd64} : s = 255;
	{8'd191,8'd65} : s = 256;
	{8'd191,8'd66} : s = 257;
	{8'd191,8'd67} : s = 258;
	{8'd191,8'd68} : s = 259;
	{8'd191,8'd69} : s = 260;
	{8'd191,8'd70} : s = 261;
	{8'd191,8'd71} : s = 262;
	{8'd191,8'd72} : s = 263;
	{8'd191,8'd73} : s = 264;
	{8'd191,8'd74} : s = 265;
	{8'd191,8'd75} : s = 266;
	{8'd191,8'd76} : s = 267;
	{8'd191,8'd77} : s = 268;
	{8'd191,8'd78} : s = 269;
	{8'd191,8'd79} : s = 270;
	{8'd191,8'd80} : s = 271;
	{8'd191,8'd81} : s = 272;
	{8'd191,8'd82} : s = 273;
	{8'd191,8'd83} : s = 274;
	{8'd191,8'd84} : s = 275;
	{8'd191,8'd85} : s = 276;
	{8'd191,8'd86} : s = 277;
	{8'd191,8'd87} : s = 278;
	{8'd191,8'd88} : s = 279;
	{8'd191,8'd89} : s = 280;
	{8'd191,8'd90} : s = 281;
	{8'd191,8'd91} : s = 282;
	{8'd191,8'd92} : s = 283;
	{8'd191,8'd93} : s = 284;
	{8'd191,8'd94} : s = 285;
	{8'd191,8'd95} : s = 286;
	{8'd191,8'd96} : s = 287;
	{8'd191,8'd97} : s = 288;
	{8'd191,8'd98} : s = 289;
	{8'd191,8'd99} : s = 290;
	{8'd191,8'd100} : s = 291;
	{8'd191,8'd101} : s = 292;
	{8'd191,8'd102} : s = 293;
	{8'd191,8'd103} : s = 294;
	{8'd191,8'd104} : s = 295;
	{8'd191,8'd105} : s = 296;
	{8'd191,8'd106} : s = 297;
	{8'd191,8'd107} : s = 298;
	{8'd191,8'd108} : s = 299;
	{8'd191,8'd109} : s = 300;
	{8'd191,8'd110} : s = 301;
	{8'd191,8'd111} : s = 302;
	{8'd191,8'd112} : s = 303;
	{8'd191,8'd113} : s = 304;
	{8'd191,8'd114} : s = 305;
	{8'd191,8'd115} : s = 306;
	{8'd191,8'd116} : s = 307;
	{8'd191,8'd117} : s = 308;
	{8'd191,8'd118} : s = 309;
	{8'd191,8'd119} : s = 310;
	{8'd191,8'd120} : s = 311;
	{8'd191,8'd121} : s = 312;
	{8'd191,8'd122} : s = 313;
	{8'd191,8'd123} : s = 314;
	{8'd191,8'd124} : s = 315;
	{8'd191,8'd125} : s = 316;
	{8'd191,8'd126} : s = 317;
	{8'd191,8'd127} : s = 318;
	{8'd191,8'd128} : s = 319;
	{8'd191,8'd129} : s = 320;
	{8'd191,8'd130} : s = 321;
	{8'd191,8'd131} : s = 322;
	{8'd191,8'd132} : s = 323;
	{8'd191,8'd133} : s = 324;
	{8'd191,8'd134} : s = 325;
	{8'd191,8'd135} : s = 326;
	{8'd191,8'd136} : s = 327;
	{8'd191,8'd137} : s = 328;
	{8'd191,8'd138} : s = 329;
	{8'd191,8'd139} : s = 330;
	{8'd191,8'd140} : s = 331;
	{8'd191,8'd141} : s = 332;
	{8'd191,8'd142} : s = 333;
	{8'd191,8'd143} : s = 334;
	{8'd191,8'd144} : s = 335;
	{8'd191,8'd145} : s = 336;
	{8'd191,8'd146} : s = 337;
	{8'd191,8'd147} : s = 338;
	{8'd191,8'd148} : s = 339;
	{8'd191,8'd149} : s = 340;
	{8'd191,8'd150} : s = 341;
	{8'd191,8'd151} : s = 342;
	{8'd191,8'd152} : s = 343;
	{8'd191,8'd153} : s = 344;
	{8'd191,8'd154} : s = 345;
	{8'd191,8'd155} : s = 346;
	{8'd191,8'd156} : s = 347;
	{8'd191,8'd157} : s = 348;
	{8'd191,8'd158} : s = 349;
	{8'd191,8'd159} : s = 350;
	{8'd191,8'd160} : s = 351;
	{8'd191,8'd161} : s = 352;
	{8'd191,8'd162} : s = 353;
	{8'd191,8'd163} : s = 354;
	{8'd191,8'd164} : s = 355;
	{8'd191,8'd165} : s = 356;
	{8'd191,8'd166} : s = 357;
	{8'd191,8'd167} : s = 358;
	{8'd191,8'd168} : s = 359;
	{8'd191,8'd169} : s = 360;
	{8'd191,8'd170} : s = 361;
	{8'd191,8'd171} : s = 362;
	{8'd191,8'd172} : s = 363;
	{8'd191,8'd173} : s = 364;
	{8'd191,8'd174} : s = 365;
	{8'd191,8'd175} : s = 366;
	{8'd191,8'd176} : s = 367;
	{8'd191,8'd177} : s = 368;
	{8'd191,8'd178} : s = 369;
	{8'd191,8'd179} : s = 370;
	{8'd191,8'd180} : s = 371;
	{8'd191,8'd181} : s = 372;
	{8'd191,8'd182} : s = 373;
	{8'd191,8'd183} : s = 374;
	{8'd191,8'd184} : s = 375;
	{8'd191,8'd185} : s = 376;
	{8'd191,8'd186} : s = 377;
	{8'd191,8'd187} : s = 378;
	{8'd191,8'd188} : s = 379;
	{8'd191,8'd189} : s = 380;
	{8'd191,8'd190} : s = 381;
	{8'd191,8'd191} : s = 382;
	{8'd191,8'd192} : s = 383;
	{8'd191,8'd193} : s = 384;
	{8'd191,8'd194} : s = 385;
	{8'd191,8'd195} : s = 386;
	{8'd191,8'd196} : s = 387;
	{8'd191,8'd197} : s = 388;
	{8'd191,8'd198} : s = 389;
	{8'd191,8'd199} : s = 390;
	{8'd191,8'd200} : s = 391;
	{8'd191,8'd201} : s = 392;
	{8'd191,8'd202} : s = 393;
	{8'd191,8'd203} : s = 394;
	{8'd191,8'd204} : s = 395;
	{8'd191,8'd205} : s = 396;
	{8'd191,8'd206} : s = 397;
	{8'd191,8'd207} : s = 398;
	{8'd191,8'd208} : s = 399;
	{8'd191,8'd209} : s = 400;
	{8'd191,8'd210} : s = 401;
	{8'd191,8'd211} : s = 402;
	{8'd191,8'd212} : s = 403;
	{8'd191,8'd213} : s = 404;
	{8'd191,8'd214} : s = 405;
	{8'd191,8'd215} : s = 406;
	{8'd191,8'd216} : s = 407;
	{8'd191,8'd217} : s = 408;
	{8'd191,8'd218} : s = 409;
	{8'd191,8'd219} : s = 410;
	{8'd191,8'd220} : s = 411;
	{8'd191,8'd221} : s = 412;
	{8'd191,8'd222} : s = 413;
	{8'd191,8'd223} : s = 414;
	{8'd191,8'd224} : s = 415;
	{8'd191,8'd225} : s = 416;
	{8'd191,8'd226} : s = 417;
	{8'd191,8'd227} : s = 418;
	{8'd191,8'd228} : s = 419;
	{8'd191,8'd229} : s = 420;
	{8'd191,8'd230} : s = 421;
	{8'd191,8'd231} : s = 422;
	{8'd191,8'd232} : s = 423;
	{8'd191,8'd233} : s = 424;
	{8'd191,8'd234} : s = 425;
	{8'd191,8'd235} : s = 426;
	{8'd191,8'd236} : s = 427;
	{8'd191,8'd237} : s = 428;
	{8'd191,8'd238} : s = 429;
	{8'd191,8'd239} : s = 430;
	{8'd191,8'd240} : s = 431;
	{8'd191,8'd241} : s = 432;
	{8'd191,8'd242} : s = 433;
	{8'd191,8'd243} : s = 434;
	{8'd191,8'd244} : s = 435;
	{8'd191,8'd245} : s = 436;
	{8'd191,8'd246} : s = 437;
	{8'd191,8'd247} : s = 438;
	{8'd191,8'd248} : s = 439;
	{8'd191,8'd249} : s = 440;
	{8'd191,8'd250} : s = 441;
	{8'd191,8'd251} : s = 442;
	{8'd191,8'd252} : s = 443;
	{8'd191,8'd253} : s = 444;
	{8'd191,8'd254} : s = 445;
	{8'd191,8'd255} : s = 446;
	{8'd192,8'd0} : s = 192;
	{8'd192,8'd1} : s = 193;
	{8'd192,8'd2} : s = 194;
	{8'd192,8'd3} : s = 195;
	{8'd192,8'd4} : s = 196;
	{8'd192,8'd5} : s = 197;
	{8'd192,8'd6} : s = 198;
	{8'd192,8'd7} : s = 199;
	{8'd192,8'd8} : s = 200;
	{8'd192,8'd9} : s = 201;
	{8'd192,8'd10} : s = 202;
	{8'd192,8'd11} : s = 203;
	{8'd192,8'd12} : s = 204;
	{8'd192,8'd13} : s = 205;
	{8'd192,8'd14} : s = 206;
	{8'd192,8'd15} : s = 207;
	{8'd192,8'd16} : s = 208;
	{8'd192,8'd17} : s = 209;
	{8'd192,8'd18} : s = 210;
	{8'd192,8'd19} : s = 211;
	{8'd192,8'd20} : s = 212;
	{8'd192,8'd21} : s = 213;
	{8'd192,8'd22} : s = 214;
	{8'd192,8'd23} : s = 215;
	{8'd192,8'd24} : s = 216;
	{8'd192,8'd25} : s = 217;
	{8'd192,8'd26} : s = 218;
	{8'd192,8'd27} : s = 219;
	{8'd192,8'd28} : s = 220;
	{8'd192,8'd29} : s = 221;
	{8'd192,8'd30} : s = 222;
	{8'd192,8'd31} : s = 223;
	{8'd192,8'd32} : s = 224;
	{8'd192,8'd33} : s = 225;
	{8'd192,8'd34} : s = 226;
	{8'd192,8'd35} : s = 227;
	{8'd192,8'd36} : s = 228;
	{8'd192,8'd37} : s = 229;
	{8'd192,8'd38} : s = 230;
	{8'd192,8'd39} : s = 231;
	{8'd192,8'd40} : s = 232;
	{8'd192,8'd41} : s = 233;
	{8'd192,8'd42} : s = 234;
	{8'd192,8'd43} : s = 235;
	{8'd192,8'd44} : s = 236;
	{8'd192,8'd45} : s = 237;
	{8'd192,8'd46} : s = 238;
	{8'd192,8'd47} : s = 239;
	{8'd192,8'd48} : s = 240;
	{8'd192,8'd49} : s = 241;
	{8'd192,8'd50} : s = 242;
	{8'd192,8'd51} : s = 243;
	{8'd192,8'd52} : s = 244;
	{8'd192,8'd53} : s = 245;
	{8'd192,8'd54} : s = 246;
	{8'd192,8'd55} : s = 247;
	{8'd192,8'd56} : s = 248;
	{8'd192,8'd57} : s = 249;
	{8'd192,8'd58} : s = 250;
	{8'd192,8'd59} : s = 251;
	{8'd192,8'd60} : s = 252;
	{8'd192,8'd61} : s = 253;
	{8'd192,8'd62} : s = 254;
	{8'd192,8'd63} : s = 255;
	{8'd192,8'd64} : s = 256;
	{8'd192,8'd65} : s = 257;
	{8'd192,8'd66} : s = 258;
	{8'd192,8'd67} : s = 259;
	{8'd192,8'd68} : s = 260;
	{8'd192,8'd69} : s = 261;
	{8'd192,8'd70} : s = 262;
	{8'd192,8'd71} : s = 263;
	{8'd192,8'd72} : s = 264;
	{8'd192,8'd73} : s = 265;
	{8'd192,8'd74} : s = 266;
	{8'd192,8'd75} : s = 267;
	{8'd192,8'd76} : s = 268;
	{8'd192,8'd77} : s = 269;
	{8'd192,8'd78} : s = 270;
	{8'd192,8'd79} : s = 271;
	{8'd192,8'd80} : s = 272;
	{8'd192,8'd81} : s = 273;
	{8'd192,8'd82} : s = 274;
	{8'd192,8'd83} : s = 275;
	{8'd192,8'd84} : s = 276;
	{8'd192,8'd85} : s = 277;
	{8'd192,8'd86} : s = 278;
	{8'd192,8'd87} : s = 279;
	{8'd192,8'd88} : s = 280;
	{8'd192,8'd89} : s = 281;
	{8'd192,8'd90} : s = 282;
	{8'd192,8'd91} : s = 283;
	{8'd192,8'd92} : s = 284;
	{8'd192,8'd93} : s = 285;
	{8'd192,8'd94} : s = 286;
	{8'd192,8'd95} : s = 287;
	{8'd192,8'd96} : s = 288;
	{8'd192,8'd97} : s = 289;
	{8'd192,8'd98} : s = 290;
	{8'd192,8'd99} : s = 291;
	{8'd192,8'd100} : s = 292;
	{8'd192,8'd101} : s = 293;
	{8'd192,8'd102} : s = 294;
	{8'd192,8'd103} : s = 295;
	{8'd192,8'd104} : s = 296;
	{8'd192,8'd105} : s = 297;
	{8'd192,8'd106} : s = 298;
	{8'd192,8'd107} : s = 299;
	{8'd192,8'd108} : s = 300;
	{8'd192,8'd109} : s = 301;
	{8'd192,8'd110} : s = 302;
	{8'd192,8'd111} : s = 303;
	{8'd192,8'd112} : s = 304;
	{8'd192,8'd113} : s = 305;
	{8'd192,8'd114} : s = 306;
	{8'd192,8'd115} : s = 307;
	{8'd192,8'd116} : s = 308;
	{8'd192,8'd117} : s = 309;
	{8'd192,8'd118} : s = 310;
	{8'd192,8'd119} : s = 311;
	{8'd192,8'd120} : s = 312;
	{8'd192,8'd121} : s = 313;
	{8'd192,8'd122} : s = 314;
	{8'd192,8'd123} : s = 315;
	{8'd192,8'd124} : s = 316;
	{8'd192,8'd125} : s = 317;
	{8'd192,8'd126} : s = 318;
	{8'd192,8'd127} : s = 319;
	{8'd192,8'd128} : s = 320;
	{8'd192,8'd129} : s = 321;
	{8'd192,8'd130} : s = 322;
	{8'd192,8'd131} : s = 323;
	{8'd192,8'd132} : s = 324;
	{8'd192,8'd133} : s = 325;
	{8'd192,8'd134} : s = 326;
	{8'd192,8'd135} : s = 327;
	{8'd192,8'd136} : s = 328;
	{8'd192,8'd137} : s = 329;
	{8'd192,8'd138} : s = 330;
	{8'd192,8'd139} : s = 331;
	{8'd192,8'd140} : s = 332;
	{8'd192,8'd141} : s = 333;
	{8'd192,8'd142} : s = 334;
	{8'd192,8'd143} : s = 335;
	{8'd192,8'd144} : s = 336;
	{8'd192,8'd145} : s = 337;
	{8'd192,8'd146} : s = 338;
	{8'd192,8'd147} : s = 339;
	{8'd192,8'd148} : s = 340;
	{8'd192,8'd149} : s = 341;
	{8'd192,8'd150} : s = 342;
	{8'd192,8'd151} : s = 343;
	{8'd192,8'd152} : s = 344;
	{8'd192,8'd153} : s = 345;
	{8'd192,8'd154} : s = 346;
	{8'd192,8'd155} : s = 347;
	{8'd192,8'd156} : s = 348;
	{8'd192,8'd157} : s = 349;
	{8'd192,8'd158} : s = 350;
	{8'd192,8'd159} : s = 351;
	{8'd192,8'd160} : s = 352;
	{8'd192,8'd161} : s = 353;
	{8'd192,8'd162} : s = 354;
	{8'd192,8'd163} : s = 355;
	{8'd192,8'd164} : s = 356;
	{8'd192,8'd165} : s = 357;
	{8'd192,8'd166} : s = 358;
	{8'd192,8'd167} : s = 359;
	{8'd192,8'd168} : s = 360;
	{8'd192,8'd169} : s = 361;
	{8'd192,8'd170} : s = 362;
	{8'd192,8'd171} : s = 363;
	{8'd192,8'd172} : s = 364;
	{8'd192,8'd173} : s = 365;
	{8'd192,8'd174} : s = 366;
	{8'd192,8'd175} : s = 367;
	{8'd192,8'd176} : s = 368;
	{8'd192,8'd177} : s = 369;
	{8'd192,8'd178} : s = 370;
	{8'd192,8'd179} : s = 371;
	{8'd192,8'd180} : s = 372;
	{8'd192,8'd181} : s = 373;
	{8'd192,8'd182} : s = 374;
	{8'd192,8'd183} : s = 375;
	{8'd192,8'd184} : s = 376;
	{8'd192,8'd185} : s = 377;
	{8'd192,8'd186} : s = 378;
	{8'd192,8'd187} : s = 379;
	{8'd192,8'd188} : s = 380;
	{8'd192,8'd189} : s = 381;
	{8'd192,8'd190} : s = 382;
	{8'd192,8'd191} : s = 383;
	{8'd192,8'd192} : s = 384;
	{8'd192,8'd193} : s = 385;
	{8'd192,8'd194} : s = 386;
	{8'd192,8'd195} : s = 387;
	{8'd192,8'd196} : s = 388;
	{8'd192,8'd197} : s = 389;
	{8'd192,8'd198} : s = 390;
	{8'd192,8'd199} : s = 391;
	{8'd192,8'd200} : s = 392;
	{8'd192,8'd201} : s = 393;
	{8'd192,8'd202} : s = 394;
	{8'd192,8'd203} : s = 395;
	{8'd192,8'd204} : s = 396;
	{8'd192,8'd205} : s = 397;
	{8'd192,8'd206} : s = 398;
	{8'd192,8'd207} : s = 399;
	{8'd192,8'd208} : s = 400;
	{8'd192,8'd209} : s = 401;
	{8'd192,8'd210} : s = 402;
	{8'd192,8'd211} : s = 403;
	{8'd192,8'd212} : s = 404;
	{8'd192,8'd213} : s = 405;
	{8'd192,8'd214} : s = 406;
	{8'd192,8'd215} : s = 407;
	{8'd192,8'd216} : s = 408;
	{8'd192,8'd217} : s = 409;
	{8'd192,8'd218} : s = 410;
	{8'd192,8'd219} : s = 411;
	{8'd192,8'd220} : s = 412;
	{8'd192,8'd221} : s = 413;
	{8'd192,8'd222} : s = 414;
	{8'd192,8'd223} : s = 415;
	{8'd192,8'd224} : s = 416;
	{8'd192,8'd225} : s = 417;
	{8'd192,8'd226} : s = 418;
	{8'd192,8'd227} : s = 419;
	{8'd192,8'd228} : s = 420;
	{8'd192,8'd229} : s = 421;
	{8'd192,8'd230} : s = 422;
	{8'd192,8'd231} : s = 423;
	{8'd192,8'd232} : s = 424;
	{8'd192,8'd233} : s = 425;
	{8'd192,8'd234} : s = 426;
	{8'd192,8'd235} : s = 427;
	{8'd192,8'd236} : s = 428;
	{8'd192,8'd237} : s = 429;
	{8'd192,8'd238} : s = 430;
	{8'd192,8'd239} : s = 431;
	{8'd192,8'd240} : s = 432;
	{8'd192,8'd241} : s = 433;
	{8'd192,8'd242} : s = 434;
	{8'd192,8'd243} : s = 435;
	{8'd192,8'd244} : s = 436;
	{8'd192,8'd245} : s = 437;
	{8'd192,8'd246} : s = 438;
	{8'd192,8'd247} : s = 439;
	{8'd192,8'd248} : s = 440;
	{8'd192,8'd249} : s = 441;
	{8'd192,8'd250} : s = 442;
	{8'd192,8'd251} : s = 443;
	{8'd192,8'd252} : s = 444;
	{8'd192,8'd253} : s = 445;
	{8'd192,8'd254} : s = 446;
	{8'd192,8'd255} : s = 447;
	{8'd193,8'd0} : s = 193;
	{8'd193,8'd1} : s = 194;
	{8'd193,8'd2} : s = 195;
	{8'd193,8'd3} : s = 196;
	{8'd193,8'd4} : s = 197;
	{8'd193,8'd5} : s = 198;
	{8'd193,8'd6} : s = 199;
	{8'd193,8'd7} : s = 200;
	{8'd193,8'd8} : s = 201;
	{8'd193,8'd9} : s = 202;
	{8'd193,8'd10} : s = 203;
	{8'd193,8'd11} : s = 204;
	{8'd193,8'd12} : s = 205;
	{8'd193,8'd13} : s = 206;
	{8'd193,8'd14} : s = 207;
	{8'd193,8'd15} : s = 208;
	{8'd193,8'd16} : s = 209;
	{8'd193,8'd17} : s = 210;
	{8'd193,8'd18} : s = 211;
	{8'd193,8'd19} : s = 212;
	{8'd193,8'd20} : s = 213;
	{8'd193,8'd21} : s = 214;
	{8'd193,8'd22} : s = 215;
	{8'd193,8'd23} : s = 216;
	{8'd193,8'd24} : s = 217;
	{8'd193,8'd25} : s = 218;
	{8'd193,8'd26} : s = 219;
	{8'd193,8'd27} : s = 220;
	{8'd193,8'd28} : s = 221;
	{8'd193,8'd29} : s = 222;
	{8'd193,8'd30} : s = 223;
	{8'd193,8'd31} : s = 224;
	{8'd193,8'd32} : s = 225;
	{8'd193,8'd33} : s = 226;
	{8'd193,8'd34} : s = 227;
	{8'd193,8'd35} : s = 228;
	{8'd193,8'd36} : s = 229;
	{8'd193,8'd37} : s = 230;
	{8'd193,8'd38} : s = 231;
	{8'd193,8'd39} : s = 232;
	{8'd193,8'd40} : s = 233;
	{8'd193,8'd41} : s = 234;
	{8'd193,8'd42} : s = 235;
	{8'd193,8'd43} : s = 236;
	{8'd193,8'd44} : s = 237;
	{8'd193,8'd45} : s = 238;
	{8'd193,8'd46} : s = 239;
	{8'd193,8'd47} : s = 240;
	{8'd193,8'd48} : s = 241;
	{8'd193,8'd49} : s = 242;
	{8'd193,8'd50} : s = 243;
	{8'd193,8'd51} : s = 244;
	{8'd193,8'd52} : s = 245;
	{8'd193,8'd53} : s = 246;
	{8'd193,8'd54} : s = 247;
	{8'd193,8'd55} : s = 248;
	{8'd193,8'd56} : s = 249;
	{8'd193,8'd57} : s = 250;
	{8'd193,8'd58} : s = 251;
	{8'd193,8'd59} : s = 252;
	{8'd193,8'd60} : s = 253;
	{8'd193,8'd61} : s = 254;
	{8'd193,8'd62} : s = 255;
	{8'd193,8'd63} : s = 256;
	{8'd193,8'd64} : s = 257;
	{8'd193,8'd65} : s = 258;
	{8'd193,8'd66} : s = 259;
	{8'd193,8'd67} : s = 260;
	{8'd193,8'd68} : s = 261;
	{8'd193,8'd69} : s = 262;
	{8'd193,8'd70} : s = 263;
	{8'd193,8'd71} : s = 264;
	{8'd193,8'd72} : s = 265;
	{8'd193,8'd73} : s = 266;
	{8'd193,8'd74} : s = 267;
	{8'd193,8'd75} : s = 268;
	{8'd193,8'd76} : s = 269;
	{8'd193,8'd77} : s = 270;
	{8'd193,8'd78} : s = 271;
	{8'd193,8'd79} : s = 272;
	{8'd193,8'd80} : s = 273;
	{8'd193,8'd81} : s = 274;
	{8'd193,8'd82} : s = 275;
	{8'd193,8'd83} : s = 276;
	{8'd193,8'd84} : s = 277;
	{8'd193,8'd85} : s = 278;
	{8'd193,8'd86} : s = 279;
	{8'd193,8'd87} : s = 280;
	{8'd193,8'd88} : s = 281;
	{8'd193,8'd89} : s = 282;
	{8'd193,8'd90} : s = 283;
	{8'd193,8'd91} : s = 284;
	{8'd193,8'd92} : s = 285;
	{8'd193,8'd93} : s = 286;
	{8'd193,8'd94} : s = 287;
	{8'd193,8'd95} : s = 288;
	{8'd193,8'd96} : s = 289;
	{8'd193,8'd97} : s = 290;
	{8'd193,8'd98} : s = 291;
	{8'd193,8'd99} : s = 292;
	{8'd193,8'd100} : s = 293;
	{8'd193,8'd101} : s = 294;
	{8'd193,8'd102} : s = 295;
	{8'd193,8'd103} : s = 296;
	{8'd193,8'd104} : s = 297;
	{8'd193,8'd105} : s = 298;
	{8'd193,8'd106} : s = 299;
	{8'd193,8'd107} : s = 300;
	{8'd193,8'd108} : s = 301;
	{8'd193,8'd109} : s = 302;
	{8'd193,8'd110} : s = 303;
	{8'd193,8'd111} : s = 304;
	{8'd193,8'd112} : s = 305;
	{8'd193,8'd113} : s = 306;
	{8'd193,8'd114} : s = 307;
	{8'd193,8'd115} : s = 308;
	{8'd193,8'd116} : s = 309;
	{8'd193,8'd117} : s = 310;
	{8'd193,8'd118} : s = 311;
	{8'd193,8'd119} : s = 312;
	{8'd193,8'd120} : s = 313;
	{8'd193,8'd121} : s = 314;
	{8'd193,8'd122} : s = 315;
	{8'd193,8'd123} : s = 316;
	{8'd193,8'd124} : s = 317;
	{8'd193,8'd125} : s = 318;
	{8'd193,8'd126} : s = 319;
	{8'd193,8'd127} : s = 320;
	{8'd193,8'd128} : s = 321;
	{8'd193,8'd129} : s = 322;
	{8'd193,8'd130} : s = 323;
	{8'd193,8'd131} : s = 324;
	{8'd193,8'd132} : s = 325;
	{8'd193,8'd133} : s = 326;
	{8'd193,8'd134} : s = 327;
	{8'd193,8'd135} : s = 328;
	{8'd193,8'd136} : s = 329;
	{8'd193,8'd137} : s = 330;
	{8'd193,8'd138} : s = 331;
	{8'd193,8'd139} : s = 332;
	{8'd193,8'd140} : s = 333;
	{8'd193,8'd141} : s = 334;
	{8'd193,8'd142} : s = 335;
	{8'd193,8'd143} : s = 336;
	{8'd193,8'd144} : s = 337;
	{8'd193,8'd145} : s = 338;
	{8'd193,8'd146} : s = 339;
	{8'd193,8'd147} : s = 340;
	{8'd193,8'd148} : s = 341;
	{8'd193,8'd149} : s = 342;
	{8'd193,8'd150} : s = 343;
	{8'd193,8'd151} : s = 344;
	{8'd193,8'd152} : s = 345;
	{8'd193,8'd153} : s = 346;
	{8'd193,8'd154} : s = 347;
	{8'd193,8'd155} : s = 348;
	{8'd193,8'd156} : s = 349;
	{8'd193,8'd157} : s = 350;
	{8'd193,8'd158} : s = 351;
	{8'd193,8'd159} : s = 352;
	{8'd193,8'd160} : s = 353;
	{8'd193,8'd161} : s = 354;
	{8'd193,8'd162} : s = 355;
	{8'd193,8'd163} : s = 356;
	{8'd193,8'd164} : s = 357;
	{8'd193,8'd165} : s = 358;
	{8'd193,8'd166} : s = 359;
	{8'd193,8'd167} : s = 360;
	{8'd193,8'd168} : s = 361;
	{8'd193,8'd169} : s = 362;
	{8'd193,8'd170} : s = 363;
	{8'd193,8'd171} : s = 364;
	{8'd193,8'd172} : s = 365;
	{8'd193,8'd173} : s = 366;
	{8'd193,8'd174} : s = 367;
	{8'd193,8'd175} : s = 368;
	{8'd193,8'd176} : s = 369;
	{8'd193,8'd177} : s = 370;
	{8'd193,8'd178} : s = 371;
	{8'd193,8'd179} : s = 372;
	{8'd193,8'd180} : s = 373;
	{8'd193,8'd181} : s = 374;
	{8'd193,8'd182} : s = 375;
	{8'd193,8'd183} : s = 376;
	{8'd193,8'd184} : s = 377;
	{8'd193,8'd185} : s = 378;
	{8'd193,8'd186} : s = 379;
	{8'd193,8'd187} : s = 380;
	{8'd193,8'd188} : s = 381;
	{8'd193,8'd189} : s = 382;
	{8'd193,8'd190} : s = 383;
	{8'd193,8'd191} : s = 384;
	{8'd193,8'd192} : s = 385;
	{8'd193,8'd193} : s = 386;
	{8'd193,8'd194} : s = 387;
	{8'd193,8'd195} : s = 388;
	{8'd193,8'd196} : s = 389;
	{8'd193,8'd197} : s = 390;
	{8'd193,8'd198} : s = 391;
	{8'd193,8'd199} : s = 392;
	{8'd193,8'd200} : s = 393;
	{8'd193,8'd201} : s = 394;
	{8'd193,8'd202} : s = 395;
	{8'd193,8'd203} : s = 396;
	{8'd193,8'd204} : s = 397;
	{8'd193,8'd205} : s = 398;
	{8'd193,8'd206} : s = 399;
	{8'd193,8'd207} : s = 400;
	{8'd193,8'd208} : s = 401;
	{8'd193,8'd209} : s = 402;
	{8'd193,8'd210} : s = 403;
	{8'd193,8'd211} : s = 404;
	{8'd193,8'd212} : s = 405;
	{8'd193,8'd213} : s = 406;
	{8'd193,8'd214} : s = 407;
	{8'd193,8'd215} : s = 408;
	{8'd193,8'd216} : s = 409;
	{8'd193,8'd217} : s = 410;
	{8'd193,8'd218} : s = 411;
	{8'd193,8'd219} : s = 412;
	{8'd193,8'd220} : s = 413;
	{8'd193,8'd221} : s = 414;
	{8'd193,8'd222} : s = 415;
	{8'd193,8'd223} : s = 416;
	{8'd193,8'd224} : s = 417;
	{8'd193,8'd225} : s = 418;
	{8'd193,8'd226} : s = 419;
	{8'd193,8'd227} : s = 420;
	{8'd193,8'd228} : s = 421;
	{8'd193,8'd229} : s = 422;
	{8'd193,8'd230} : s = 423;
	{8'd193,8'd231} : s = 424;
	{8'd193,8'd232} : s = 425;
	{8'd193,8'd233} : s = 426;
	{8'd193,8'd234} : s = 427;
	{8'd193,8'd235} : s = 428;
	{8'd193,8'd236} : s = 429;
	{8'd193,8'd237} : s = 430;
	{8'd193,8'd238} : s = 431;
	{8'd193,8'd239} : s = 432;
	{8'd193,8'd240} : s = 433;
	{8'd193,8'd241} : s = 434;
	{8'd193,8'd242} : s = 435;
	{8'd193,8'd243} : s = 436;
	{8'd193,8'd244} : s = 437;
	{8'd193,8'd245} : s = 438;
	{8'd193,8'd246} : s = 439;
	{8'd193,8'd247} : s = 440;
	{8'd193,8'd248} : s = 441;
	{8'd193,8'd249} : s = 442;
	{8'd193,8'd250} : s = 443;
	{8'd193,8'd251} : s = 444;
	{8'd193,8'd252} : s = 445;
	{8'd193,8'd253} : s = 446;
	{8'd193,8'd254} : s = 447;
	{8'd193,8'd255} : s = 448;
	{8'd194,8'd0} : s = 194;
	{8'd194,8'd1} : s = 195;
	{8'd194,8'd2} : s = 196;
	{8'd194,8'd3} : s = 197;
	{8'd194,8'd4} : s = 198;
	{8'd194,8'd5} : s = 199;
	{8'd194,8'd6} : s = 200;
	{8'd194,8'd7} : s = 201;
	{8'd194,8'd8} : s = 202;
	{8'd194,8'd9} : s = 203;
	{8'd194,8'd10} : s = 204;
	{8'd194,8'd11} : s = 205;
	{8'd194,8'd12} : s = 206;
	{8'd194,8'd13} : s = 207;
	{8'd194,8'd14} : s = 208;
	{8'd194,8'd15} : s = 209;
	{8'd194,8'd16} : s = 210;
	{8'd194,8'd17} : s = 211;
	{8'd194,8'd18} : s = 212;
	{8'd194,8'd19} : s = 213;
	{8'd194,8'd20} : s = 214;
	{8'd194,8'd21} : s = 215;
	{8'd194,8'd22} : s = 216;
	{8'd194,8'd23} : s = 217;
	{8'd194,8'd24} : s = 218;
	{8'd194,8'd25} : s = 219;
	{8'd194,8'd26} : s = 220;
	{8'd194,8'd27} : s = 221;
	{8'd194,8'd28} : s = 222;
	{8'd194,8'd29} : s = 223;
	{8'd194,8'd30} : s = 224;
	{8'd194,8'd31} : s = 225;
	{8'd194,8'd32} : s = 226;
	{8'd194,8'd33} : s = 227;
	{8'd194,8'd34} : s = 228;
	{8'd194,8'd35} : s = 229;
	{8'd194,8'd36} : s = 230;
	{8'd194,8'd37} : s = 231;
	{8'd194,8'd38} : s = 232;
	{8'd194,8'd39} : s = 233;
	{8'd194,8'd40} : s = 234;
	{8'd194,8'd41} : s = 235;
	{8'd194,8'd42} : s = 236;
	{8'd194,8'd43} : s = 237;
	{8'd194,8'd44} : s = 238;
	{8'd194,8'd45} : s = 239;
	{8'd194,8'd46} : s = 240;
	{8'd194,8'd47} : s = 241;
	{8'd194,8'd48} : s = 242;
	{8'd194,8'd49} : s = 243;
	{8'd194,8'd50} : s = 244;
	{8'd194,8'd51} : s = 245;
	{8'd194,8'd52} : s = 246;
	{8'd194,8'd53} : s = 247;
	{8'd194,8'd54} : s = 248;
	{8'd194,8'd55} : s = 249;
	{8'd194,8'd56} : s = 250;
	{8'd194,8'd57} : s = 251;
	{8'd194,8'd58} : s = 252;
	{8'd194,8'd59} : s = 253;
	{8'd194,8'd60} : s = 254;
	{8'd194,8'd61} : s = 255;
	{8'd194,8'd62} : s = 256;
	{8'd194,8'd63} : s = 257;
	{8'd194,8'd64} : s = 258;
	{8'd194,8'd65} : s = 259;
	{8'd194,8'd66} : s = 260;
	{8'd194,8'd67} : s = 261;
	{8'd194,8'd68} : s = 262;
	{8'd194,8'd69} : s = 263;
	{8'd194,8'd70} : s = 264;
	{8'd194,8'd71} : s = 265;
	{8'd194,8'd72} : s = 266;
	{8'd194,8'd73} : s = 267;
	{8'd194,8'd74} : s = 268;
	{8'd194,8'd75} : s = 269;
	{8'd194,8'd76} : s = 270;
	{8'd194,8'd77} : s = 271;
	{8'd194,8'd78} : s = 272;
	{8'd194,8'd79} : s = 273;
	{8'd194,8'd80} : s = 274;
	{8'd194,8'd81} : s = 275;
	{8'd194,8'd82} : s = 276;
	{8'd194,8'd83} : s = 277;
	{8'd194,8'd84} : s = 278;
	{8'd194,8'd85} : s = 279;
	{8'd194,8'd86} : s = 280;
	{8'd194,8'd87} : s = 281;
	{8'd194,8'd88} : s = 282;
	{8'd194,8'd89} : s = 283;
	{8'd194,8'd90} : s = 284;
	{8'd194,8'd91} : s = 285;
	{8'd194,8'd92} : s = 286;
	{8'd194,8'd93} : s = 287;
	{8'd194,8'd94} : s = 288;
	{8'd194,8'd95} : s = 289;
	{8'd194,8'd96} : s = 290;
	{8'd194,8'd97} : s = 291;
	{8'd194,8'd98} : s = 292;
	{8'd194,8'd99} : s = 293;
	{8'd194,8'd100} : s = 294;
	{8'd194,8'd101} : s = 295;
	{8'd194,8'd102} : s = 296;
	{8'd194,8'd103} : s = 297;
	{8'd194,8'd104} : s = 298;
	{8'd194,8'd105} : s = 299;
	{8'd194,8'd106} : s = 300;
	{8'd194,8'd107} : s = 301;
	{8'd194,8'd108} : s = 302;
	{8'd194,8'd109} : s = 303;
	{8'd194,8'd110} : s = 304;
	{8'd194,8'd111} : s = 305;
	{8'd194,8'd112} : s = 306;
	{8'd194,8'd113} : s = 307;
	{8'd194,8'd114} : s = 308;
	{8'd194,8'd115} : s = 309;
	{8'd194,8'd116} : s = 310;
	{8'd194,8'd117} : s = 311;
	{8'd194,8'd118} : s = 312;
	{8'd194,8'd119} : s = 313;
	{8'd194,8'd120} : s = 314;
	{8'd194,8'd121} : s = 315;
	{8'd194,8'd122} : s = 316;
	{8'd194,8'd123} : s = 317;
	{8'd194,8'd124} : s = 318;
	{8'd194,8'd125} : s = 319;
	{8'd194,8'd126} : s = 320;
	{8'd194,8'd127} : s = 321;
	{8'd194,8'd128} : s = 322;
	{8'd194,8'd129} : s = 323;
	{8'd194,8'd130} : s = 324;
	{8'd194,8'd131} : s = 325;
	{8'd194,8'd132} : s = 326;
	{8'd194,8'd133} : s = 327;
	{8'd194,8'd134} : s = 328;
	{8'd194,8'd135} : s = 329;
	{8'd194,8'd136} : s = 330;
	{8'd194,8'd137} : s = 331;
	{8'd194,8'd138} : s = 332;
	{8'd194,8'd139} : s = 333;
	{8'd194,8'd140} : s = 334;
	{8'd194,8'd141} : s = 335;
	{8'd194,8'd142} : s = 336;
	{8'd194,8'd143} : s = 337;
	{8'd194,8'd144} : s = 338;
	{8'd194,8'd145} : s = 339;
	{8'd194,8'd146} : s = 340;
	{8'd194,8'd147} : s = 341;
	{8'd194,8'd148} : s = 342;
	{8'd194,8'd149} : s = 343;
	{8'd194,8'd150} : s = 344;
	{8'd194,8'd151} : s = 345;
	{8'd194,8'd152} : s = 346;
	{8'd194,8'd153} : s = 347;
	{8'd194,8'd154} : s = 348;
	{8'd194,8'd155} : s = 349;
	{8'd194,8'd156} : s = 350;
	{8'd194,8'd157} : s = 351;
	{8'd194,8'd158} : s = 352;
	{8'd194,8'd159} : s = 353;
	{8'd194,8'd160} : s = 354;
	{8'd194,8'd161} : s = 355;
	{8'd194,8'd162} : s = 356;
	{8'd194,8'd163} : s = 357;
	{8'd194,8'd164} : s = 358;
	{8'd194,8'd165} : s = 359;
	{8'd194,8'd166} : s = 360;
	{8'd194,8'd167} : s = 361;
	{8'd194,8'd168} : s = 362;
	{8'd194,8'd169} : s = 363;
	{8'd194,8'd170} : s = 364;
	{8'd194,8'd171} : s = 365;
	{8'd194,8'd172} : s = 366;
	{8'd194,8'd173} : s = 367;
	{8'd194,8'd174} : s = 368;
	{8'd194,8'd175} : s = 369;
	{8'd194,8'd176} : s = 370;
	{8'd194,8'd177} : s = 371;
	{8'd194,8'd178} : s = 372;
	{8'd194,8'd179} : s = 373;
	{8'd194,8'd180} : s = 374;
	{8'd194,8'd181} : s = 375;
	{8'd194,8'd182} : s = 376;
	{8'd194,8'd183} : s = 377;
	{8'd194,8'd184} : s = 378;
	{8'd194,8'd185} : s = 379;
	{8'd194,8'd186} : s = 380;
	{8'd194,8'd187} : s = 381;
	{8'd194,8'd188} : s = 382;
	{8'd194,8'd189} : s = 383;
	{8'd194,8'd190} : s = 384;
	{8'd194,8'd191} : s = 385;
	{8'd194,8'd192} : s = 386;
	{8'd194,8'd193} : s = 387;
	{8'd194,8'd194} : s = 388;
	{8'd194,8'd195} : s = 389;
	{8'd194,8'd196} : s = 390;
	{8'd194,8'd197} : s = 391;
	{8'd194,8'd198} : s = 392;
	{8'd194,8'd199} : s = 393;
	{8'd194,8'd200} : s = 394;
	{8'd194,8'd201} : s = 395;
	{8'd194,8'd202} : s = 396;
	{8'd194,8'd203} : s = 397;
	{8'd194,8'd204} : s = 398;
	{8'd194,8'd205} : s = 399;
	{8'd194,8'd206} : s = 400;
	{8'd194,8'd207} : s = 401;
	{8'd194,8'd208} : s = 402;
	{8'd194,8'd209} : s = 403;
	{8'd194,8'd210} : s = 404;
	{8'd194,8'd211} : s = 405;
	{8'd194,8'd212} : s = 406;
	{8'd194,8'd213} : s = 407;
	{8'd194,8'd214} : s = 408;
	{8'd194,8'd215} : s = 409;
	{8'd194,8'd216} : s = 410;
	{8'd194,8'd217} : s = 411;
	{8'd194,8'd218} : s = 412;
	{8'd194,8'd219} : s = 413;
	{8'd194,8'd220} : s = 414;
	{8'd194,8'd221} : s = 415;
	{8'd194,8'd222} : s = 416;
	{8'd194,8'd223} : s = 417;
	{8'd194,8'd224} : s = 418;
	{8'd194,8'd225} : s = 419;
	{8'd194,8'd226} : s = 420;
	{8'd194,8'd227} : s = 421;
	{8'd194,8'd228} : s = 422;
	{8'd194,8'd229} : s = 423;
	{8'd194,8'd230} : s = 424;
	{8'd194,8'd231} : s = 425;
	{8'd194,8'd232} : s = 426;
	{8'd194,8'd233} : s = 427;
	{8'd194,8'd234} : s = 428;
	{8'd194,8'd235} : s = 429;
	{8'd194,8'd236} : s = 430;
	{8'd194,8'd237} : s = 431;
	{8'd194,8'd238} : s = 432;
	{8'd194,8'd239} : s = 433;
	{8'd194,8'd240} : s = 434;
	{8'd194,8'd241} : s = 435;
	{8'd194,8'd242} : s = 436;
	{8'd194,8'd243} : s = 437;
	{8'd194,8'd244} : s = 438;
	{8'd194,8'd245} : s = 439;
	{8'd194,8'd246} : s = 440;
	{8'd194,8'd247} : s = 441;
	{8'd194,8'd248} : s = 442;
	{8'd194,8'd249} : s = 443;
	{8'd194,8'd250} : s = 444;
	{8'd194,8'd251} : s = 445;
	{8'd194,8'd252} : s = 446;
	{8'd194,8'd253} : s = 447;
	{8'd194,8'd254} : s = 448;
	{8'd194,8'd255} : s = 449;
	{8'd195,8'd0} : s = 195;
	{8'd195,8'd1} : s = 196;
	{8'd195,8'd2} : s = 197;
	{8'd195,8'd3} : s = 198;
	{8'd195,8'd4} : s = 199;
	{8'd195,8'd5} : s = 200;
	{8'd195,8'd6} : s = 201;
	{8'd195,8'd7} : s = 202;
	{8'd195,8'd8} : s = 203;
	{8'd195,8'd9} : s = 204;
	{8'd195,8'd10} : s = 205;
	{8'd195,8'd11} : s = 206;
	{8'd195,8'd12} : s = 207;
	{8'd195,8'd13} : s = 208;
	{8'd195,8'd14} : s = 209;
	{8'd195,8'd15} : s = 210;
	{8'd195,8'd16} : s = 211;
	{8'd195,8'd17} : s = 212;
	{8'd195,8'd18} : s = 213;
	{8'd195,8'd19} : s = 214;
	{8'd195,8'd20} : s = 215;
	{8'd195,8'd21} : s = 216;
	{8'd195,8'd22} : s = 217;
	{8'd195,8'd23} : s = 218;
	{8'd195,8'd24} : s = 219;
	{8'd195,8'd25} : s = 220;
	{8'd195,8'd26} : s = 221;
	{8'd195,8'd27} : s = 222;
	{8'd195,8'd28} : s = 223;
	{8'd195,8'd29} : s = 224;
	{8'd195,8'd30} : s = 225;
	{8'd195,8'd31} : s = 226;
	{8'd195,8'd32} : s = 227;
	{8'd195,8'd33} : s = 228;
	{8'd195,8'd34} : s = 229;
	{8'd195,8'd35} : s = 230;
	{8'd195,8'd36} : s = 231;
	{8'd195,8'd37} : s = 232;
	{8'd195,8'd38} : s = 233;
	{8'd195,8'd39} : s = 234;
	{8'd195,8'd40} : s = 235;
	{8'd195,8'd41} : s = 236;
	{8'd195,8'd42} : s = 237;
	{8'd195,8'd43} : s = 238;
	{8'd195,8'd44} : s = 239;
	{8'd195,8'd45} : s = 240;
	{8'd195,8'd46} : s = 241;
	{8'd195,8'd47} : s = 242;
	{8'd195,8'd48} : s = 243;
	{8'd195,8'd49} : s = 244;
	{8'd195,8'd50} : s = 245;
	{8'd195,8'd51} : s = 246;
	{8'd195,8'd52} : s = 247;
	{8'd195,8'd53} : s = 248;
	{8'd195,8'd54} : s = 249;
	{8'd195,8'd55} : s = 250;
	{8'd195,8'd56} : s = 251;
	{8'd195,8'd57} : s = 252;
	{8'd195,8'd58} : s = 253;
	{8'd195,8'd59} : s = 254;
	{8'd195,8'd60} : s = 255;
	{8'd195,8'd61} : s = 256;
	{8'd195,8'd62} : s = 257;
	{8'd195,8'd63} : s = 258;
	{8'd195,8'd64} : s = 259;
	{8'd195,8'd65} : s = 260;
	{8'd195,8'd66} : s = 261;
	{8'd195,8'd67} : s = 262;
	{8'd195,8'd68} : s = 263;
	{8'd195,8'd69} : s = 264;
	{8'd195,8'd70} : s = 265;
	{8'd195,8'd71} : s = 266;
	{8'd195,8'd72} : s = 267;
	{8'd195,8'd73} : s = 268;
	{8'd195,8'd74} : s = 269;
	{8'd195,8'd75} : s = 270;
	{8'd195,8'd76} : s = 271;
	{8'd195,8'd77} : s = 272;
	{8'd195,8'd78} : s = 273;
	{8'd195,8'd79} : s = 274;
	{8'd195,8'd80} : s = 275;
	{8'd195,8'd81} : s = 276;
	{8'd195,8'd82} : s = 277;
	{8'd195,8'd83} : s = 278;
	{8'd195,8'd84} : s = 279;
	{8'd195,8'd85} : s = 280;
	{8'd195,8'd86} : s = 281;
	{8'd195,8'd87} : s = 282;
	{8'd195,8'd88} : s = 283;
	{8'd195,8'd89} : s = 284;
	{8'd195,8'd90} : s = 285;
	{8'd195,8'd91} : s = 286;
	{8'd195,8'd92} : s = 287;
	{8'd195,8'd93} : s = 288;
	{8'd195,8'd94} : s = 289;
	{8'd195,8'd95} : s = 290;
	{8'd195,8'd96} : s = 291;
	{8'd195,8'd97} : s = 292;
	{8'd195,8'd98} : s = 293;
	{8'd195,8'd99} : s = 294;
	{8'd195,8'd100} : s = 295;
	{8'd195,8'd101} : s = 296;
	{8'd195,8'd102} : s = 297;
	{8'd195,8'd103} : s = 298;
	{8'd195,8'd104} : s = 299;
	{8'd195,8'd105} : s = 300;
	{8'd195,8'd106} : s = 301;
	{8'd195,8'd107} : s = 302;
	{8'd195,8'd108} : s = 303;
	{8'd195,8'd109} : s = 304;
	{8'd195,8'd110} : s = 305;
	{8'd195,8'd111} : s = 306;
	{8'd195,8'd112} : s = 307;
	{8'd195,8'd113} : s = 308;
	{8'd195,8'd114} : s = 309;
	{8'd195,8'd115} : s = 310;
	{8'd195,8'd116} : s = 311;
	{8'd195,8'd117} : s = 312;
	{8'd195,8'd118} : s = 313;
	{8'd195,8'd119} : s = 314;
	{8'd195,8'd120} : s = 315;
	{8'd195,8'd121} : s = 316;
	{8'd195,8'd122} : s = 317;
	{8'd195,8'd123} : s = 318;
	{8'd195,8'd124} : s = 319;
	{8'd195,8'd125} : s = 320;
	{8'd195,8'd126} : s = 321;
	{8'd195,8'd127} : s = 322;
	{8'd195,8'd128} : s = 323;
	{8'd195,8'd129} : s = 324;
	{8'd195,8'd130} : s = 325;
	{8'd195,8'd131} : s = 326;
	{8'd195,8'd132} : s = 327;
	{8'd195,8'd133} : s = 328;
	{8'd195,8'd134} : s = 329;
	{8'd195,8'd135} : s = 330;
	{8'd195,8'd136} : s = 331;
	{8'd195,8'd137} : s = 332;
	{8'd195,8'd138} : s = 333;
	{8'd195,8'd139} : s = 334;
	{8'd195,8'd140} : s = 335;
	{8'd195,8'd141} : s = 336;
	{8'd195,8'd142} : s = 337;
	{8'd195,8'd143} : s = 338;
	{8'd195,8'd144} : s = 339;
	{8'd195,8'd145} : s = 340;
	{8'd195,8'd146} : s = 341;
	{8'd195,8'd147} : s = 342;
	{8'd195,8'd148} : s = 343;
	{8'd195,8'd149} : s = 344;
	{8'd195,8'd150} : s = 345;
	{8'd195,8'd151} : s = 346;
	{8'd195,8'd152} : s = 347;
	{8'd195,8'd153} : s = 348;
	{8'd195,8'd154} : s = 349;
	{8'd195,8'd155} : s = 350;
	{8'd195,8'd156} : s = 351;
	{8'd195,8'd157} : s = 352;
	{8'd195,8'd158} : s = 353;
	{8'd195,8'd159} : s = 354;
	{8'd195,8'd160} : s = 355;
	{8'd195,8'd161} : s = 356;
	{8'd195,8'd162} : s = 357;
	{8'd195,8'd163} : s = 358;
	{8'd195,8'd164} : s = 359;
	{8'd195,8'd165} : s = 360;
	{8'd195,8'd166} : s = 361;
	{8'd195,8'd167} : s = 362;
	{8'd195,8'd168} : s = 363;
	{8'd195,8'd169} : s = 364;
	{8'd195,8'd170} : s = 365;
	{8'd195,8'd171} : s = 366;
	{8'd195,8'd172} : s = 367;
	{8'd195,8'd173} : s = 368;
	{8'd195,8'd174} : s = 369;
	{8'd195,8'd175} : s = 370;
	{8'd195,8'd176} : s = 371;
	{8'd195,8'd177} : s = 372;
	{8'd195,8'd178} : s = 373;
	{8'd195,8'd179} : s = 374;
	{8'd195,8'd180} : s = 375;
	{8'd195,8'd181} : s = 376;
	{8'd195,8'd182} : s = 377;
	{8'd195,8'd183} : s = 378;
	{8'd195,8'd184} : s = 379;
	{8'd195,8'd185} : s = 380;
	{8'd195,8'd186} : s = 381;
	{8'd195,8'd187} : s = 382;
	{8'd195,8'd188} : s = 383;
	{8'd195,8'd189} : s = 384;
	{8'd195,8'd190} : s = 385;
	{8'd195,8'd191} : s = 386;
	{8'd195,8'd192} : s = 387;
	{8'd195,8'd193} : s = 388;
	{8'd195,8'd194} : s = 389;
	{8'd195,8'd195} : s = 390;
	{8'd195,8'd196} : s = 391;
	{8'd195,8'd197} : s = 392;
	{8'd195,8'd198} : s = 393;
	{8'd195,8'd199} : s = 394;
	{8'd195,8'd200} : s = 395;
	{8'd195,8'd201} : s = 396;
	{8'd195,8'd202} : s = 397;
	{8'd195,8'd203} : s = 398;
	{8'd195,8'd204} : s = 399;
	{8'd195,8'd205} : s = 400;
	{8'd195,8'd206} : s = 401;
	{8'd195,8'd207} : s = 402;
	{8'd195,8'd208} : s = 403;
	{8'd195,8'd209} : s = 404;
	{8'd195,8'd210} : s = 405;
	{8'd195,8'd211} : s = 406;
	{8'd195,8'd212} : s = 407;
	{8'd195,8'd213} : s = 408;
	{8'd195,8'd214} : s = 409;
	{8'd195,8'd215} : s = 410;
	{8'd195,8'd216} : s = 411;
	{8'd195,8'd217} : s = 412;
	{8'd195,8'd218} : s = 413;
	{8'd195,8'd219} : s = 414;
	{8'd195,8'd220} : s = 415;
	{8'd195,8'd221} : s = 416;
	{8'd195,8'd222} : s = 417;
	{8'd195,8'd223} : s = 418;
	{8'd195,8'd224} : s = 419;
	{8'd195,8'd225} : s = 420;
	{8'd195,8'd226} : s = 421;
	{8'd195,8'd227} : s = 422;
	{8'd195,8'd228} : s = 423;
	{8'd195,8'd229} : s = 424;
	{8'd195,8'd230} : s = 425;
	{8'd195,8'd231} : s = 426;
	{8'd195,8'd232} : s = 427;
	{8'd195,8'd233} : s = 428;
	{8'd195,8'd234} : s = 429;
	{8'd195,8'd235} : s = 430;
	{8'd195,8'd236} : s = 431;
	{8'd195,8'd237} : s = 432;
	{8'd195,8'd238} : s = 433;
	{8'd195,8'd239} : s = 434;
	{8'd195,8'd240} : s = 435;
	{8'd195,8'd241} : s = 436;
	{8'd195,8'd242} : s = 437;
	{8'd195,8'd243} : s = 438;
	{8'd195,8'd244} : s = 439;
	{8'd195,8'd245} : s = 440;
	{8'd195,8'd246} : s = 441;
	{8'd195,8'd247} : s = 442;
	{8'd195,8'd248} : s = 443;
	{8'd195,8'd249} : s = 444;
	{8'd195,8'd250} : s = 445;
	{8'd195,8'd251} : s = 446;
	{8'd195,8'd252} : s = 447;
	{8'd195,8'd253} : s = 448;
	{8'd195,8'd254} : s = 449;
	{8'd195,8'd255} : s = 450;
	{8'd196,8'd0} : s = 196;
	{8'd196,8'd1} : s = 197;
	{8'd196,8'd2} : s = 198;
	{8'd196,8'd3} : s = 199;
	{8'd196,8'd4} : s = 200;
	{8'd196,8'd5} : s = 201;
	{8'd196,8'd6} : s = 202;
	{8'd196,8'd7} : s = 203;
	{8'd196,8'd8} : s = 204;
	{8'd196,8'd9} : s = 205;
	{8'd196,8'd10} : s = 206;
	{8'd196,8'd11} : s = 207;
	{8'd196,8'd12} : s = 208;
	{8'd196,8'd13} : s = 209;
	{8'd196,8'd14} : s = 210;
	{8'd196,8'd15} : s = 211;
	{8'd196,8'd16} : s = 212;
	{8'd196,8'd17} : s = 213;
	{8'd196,8'd18} : s = 214;
	{8'd196,8'd19} : s = 215;
	{8'd196,8'd20} : s = 216;
	{8'd196,8'd21} : s = 217;
	{8'd196,8'd22} : s = 218;
	{8'd196,8'd23} : s = 219;
	{8'd196,8'd24} : s = 220;
	{8'd196,8'd25} : s = 221;
	{8'd196,8'd26} : s = 222;
	{8'd196,8'd27} : s = 223;
	{8'd196,8'd28} : s = 224;
	{8'd196,8'd29} : s = 225;
	{8'd196,8'd30} : s = 226;
	{8'd196,8'd31} : s = 227;
	{8'd196,8'd32} : s = 228;
	{8'd196,8'd33} : s = 229;
	{8'd196,8'd34} : s = 230;
	{8'd196,8'd35} : s = 231;
	{8'd196,8'd36} : s = 232;
	{8'd196,8'd37} : s = 233;
	{8'd196,8'd38} : s = 234;
	{8'd196,8'd39} : s = 235;
	{8'd196,8'd40} : s = 236;
	{8'd196,8'd41} : s = 237;
	{8'd196,8'd42} : s = 238;
	{8'd196,8'd43} : s = 239;
	{8'd196,8'd44} : s = 240;
	{8'd196,8'd45} : s = 241;
	{8'd196,8'd46} : s = 242;
	{8'd196,8'd47} : s = 243;
	{8'd196,8'd48} : s = 244;
	{8'd196,8'd49} : s = 245;
	{8'd196,8'd50} : s = 246;
	{8'd196,8'd51} : s = 247;
	{8'd196,8'd52} : s = 248;
	{8'd196,8'd53} : s = 249;
	{8'd196,8'd54} : s = 250;
	{8'd196,8'd55} : s = 251;
	{8'd196,8'd56} : s = 252;
	{8'd196,8'd57} : s = 253;
	{8'd196,8'd58} : s = 254;
	{8'd196,8'd59} : s = 255;
	{8'd196,8'd60} : s = 256;
	{8'd196,8'd61} : s = 257;
	{8'd196,8'd62} : s = 258;
	{8'd196,8'd63} : s = 259;
	{8'd196,8'd64} : s = 260;
	{8'd196,8'd65} : s = 261;
	{8'd196,8'd66} : s = 262;
	{8'd196,8'd67} : s = 263;
	{8'd196,8'd68} : s = 264;
	{8'd196,8'd69} : s = 265;
	{8'd196,8'd70} : s = 266;
	{8'd196,8'd71} : s = 267;
	{8'd196,8'd72} : s = 268;
	{8'd196,8'd73} : s = 269;
	{8'd196,8'd74} : s = 270;
	{8'd196,8'd75} : s = 271;
	{8'd196,8'd76} : s = 272;
	{8'd196,8'd77} : s = 273;
	{8'd196,8'd78} : s = 274;
	{8'd196,8'd79} : s = 275;
	{8'd196,8'd80} : s = 276;
	{8'd196,8'd81} : s = 277;
	{8'd196,8'd82} : s = 278;
	{8'd196,8'd83} : s = 279;
	{8'd196,8'd84} : s = 280;
	{8'd196,8'd85} : s = 281;
	{8'd196,8'd86} : s = 282;
	{8'd196,8'd87} : s = 283;
	{8'd196,8'd88} : s = 284;
	{8'd196,8'd89} : s = 285;
	{8'd196,8'd90} : s = 286;
	{8'd196,8'd91} : s = 287;
	{8'd196,8'd92} : s = 288;
	{8'd196,8'd93} : s = 289;
	{8'd196,8'd94} : s = 290;
	{8'd196,8'd95} : s = 291;
	{8'd196,8'd96} : s = 292;
	{8'd196,8'd97} : s = 293;
	{8'd196,8'd98} : s = 294;
	{8'd196,8'd99} : s = 295;
	{8'd196,8'd100} : s = 296;
	{8'd196,8'd101} : s = 297;
	{8'd196,8'd102} : s = 298;
	{8'd196,8'd103} : s = 299;
	{8'd196,8'd104} : s = 300;
	{8'd196,8'd105} : s = 301;
	{8'd196,8'd106} : s = 302;
	{8'd196,8'd107} : s = 303;
	{8'd196,8'd108} : s = 304;
	{8'd196,8'd109} : s = 305;
	{8'd196,8'd110} : s = 306;
	{8'd196,8'd111} : s = 307;
	{8'd196,8'd112} : s = 308;
	{8'd196,8'd113} : s = 309;
	{8'd196,8'd114} : s = 310;
	{8'd196,8'd115} : s = 311;
	{8'd196,8'd116} : s = 312;
	{8'd196,8'd117} : s = 313;
	{8'd196,8'd118} : s = 314;
	{8'd196,8'd119} : s = 315;
	{8'd196,8'd120} : s = 316;
	{8'd196,8'd121} : s = 317;
	{8'd196,8'd122} : s = 318;
	{8'd196,8'd123} : s = 319;
	{8'd196,8'd124} : s = 320;
	{8'd196,8'd125} : s = 321;
	{8'd196,8'd126} : s = 322;
	{8'd196,8'd127} : s = 323;
	{8'd196,8'd128} : s = 324;
	{8'd196,8'd129} : s = 325;
	{8'd196,8'd130} : s = 326;
	{8'd196,8'd131} : s = 327;
	{8'd196,8'd132} : s = 328;
	{8'd196,8'd133} : s = 329;
	{8'd196,8'd134} : s = 330;
	{8'd196,8'd135} : s = 331;
	{8'd196,8'd136} : s = 332;
	{8'd196,8'd137} : s = 333;
	{8'd196,8'd138} : s = 334;
	{8'd196,8'd139} : s = 335;
	{8'd196,8'd140} : s = 336;
	{8'd196,8'd141} : s = 337;
	{8'd196,8'd142} : s = 338;
	{8'd196,8'd143} : s = 339;
	{8'd196,8'd144} : s = 340;
	{8'd196,8'd145} : s = 341;
	{8'd196,8'd146} : s = 342;
	{8'd196,8'd147} : s = 343;
	{8'd196,8'd148} : s = 344;
	{8'd196,8'd149} : s = 345;
	{8'd196,8'd150} : s = 346;
	{8'd196,8'd151} : s = 347;
	{8'd196,8'd152} : s = 348;
	{8'd196,8'd153} : s = 349;
	{8'd196,8'd154} : s = 350;
	{8'd196,8'd155} : s = 351;
	{8'd196,8'd156} : s = 352;
	{8'd196,8'd157} : s = 353;
	{8'd196,8'd158} : s = 354;
	{8'd196,8'd159} : s = 355;
	{8'd196,8'd160} : s = 356;
	{8'd196,8'd161} : s = 357;
	{8'd196,8'd162} : s = 358;
	{8'd196,8'd163} : s = 359;
	{8'd196,8'd164} : s = 360;
	{8'd196,8'd165} : s = 361;
	{8'd196,8'd166} : s = 362;
	{8'd196,8'd167} : s = 363;
	{8'd196,8'd168} : s = 364;
	{8'd196,8'd169} : s = 365;
	{8'd196,8'd170} : s = 366;
	{8'd196,8'd171} : s = 367;
	{8'd196,8'd172} : s = 368;
	{8'd196,8'd173} : s = 369;
	{8'd196,8'd174} : s = 370;
	{8'd196,8'd175} : s = 371;
	{8'd196,8'd176} : s = 372;
	{8'd196,8'd177} : s = 373;
	{8'd196,8'd178} : s = 374;
	{8'd196,8'd179} : s = 375;
	{8'd196,8'd180} : s = 376;
	{8'd196,8'd181} : s = 377;
	{8'd196,8'd182} : s = 378;
	{8'd196,8'd183} : s = 379;
	{8'd196,8'd184} : s = 380;
	{8'd196,8'd185} : s = 381;
	{8'd196,8'd186} : s = 382;
	{8'd196,8'd187} : s = 383;
	{8'd196,8'd188} : s = 384;
	{8'd196,8'd189} : s = 385;
	{8'd196,8'd190} : s = 386;
	{8'd196,8'd191} : s = 387;
	{8'd196,8'd192} : s = 388;
	{8'd196,8'd193} : s = 389;
	{8'd196,8'd194} : s = 390;
	{8'd196,8'd195} : s = 391;
	{8'd196,8'd196} : s = 392;
	{8'd196,8'd197} : s = 393;
	{8'd196,8'd198} : s = 394;
	{8'd196,8'd199} : s = 395;
	{8'd196,8'd200} : s = 396;
	{8'd196,8'd201} : s = 397;
	{8'd196,8'd202} : s = 398;
	{8'd196,8'd203} : s = 399;
	{8'd196,8'd204} : s = 400;
	{8'd196,8'd205} : s = 401;
	{8'd196,8'd206} : s = 402;
	{8'd196,8'd207} : s = 403;
	{8'd196,8'd208} : s = 404;
	{8'd196,8'd209} : s = 405;
	{8'd196,8'd210} : s = 406;
	{8'd196,8'd211} : s = 407;
	{8'd196,8'd212} : s = 408;
	{8'd196,8'd213} : s = 409;
	{8'd196,8'd214} : s = 410;
	{8'd196,8'd215} : s = 411;
	{8'd196,8'd216} : s = 412;
	{8'd196,8'd217} : s = 413;
	{8'd196,8'd218} : s = 414;
	{8'd196,8'd219} : s = 415;
	{8'd196,8'd220} : s = 416;
	{8'd196,8'd221} : s = 417;
	{8'd196,8'd222} : s = 418;
	{8'd196,8'd223} : s = 419;
	{8'd196,8'd224} : s = 420;
	{8'd196,8'd225} : s = 421;
	{8'd196,8'd226} : s = 422;
	{8'd196,8'd227} : s = 423;
	{8'd196,8'd228} : s = 424;
	{8'd196,8'd229} : s = 425;
	{8'd196,8'd230} : s = 426;
	{8'd196,8'd231} : s = 427;
	{8'd196,8'd232} : s = 428;
	{8'd196,8'd233} : s = 429;
	{8'd196,8'd234} : s = 430;
	{8'd196,8'd235} : s = 431;
	{8'd196,8'd236} : s = 432;
	{8'd196,8'd237} : s = 433;
	{8'd196,8'd238} : s = 434;
	{8'd196,8'd239} : s = 435;
	{8'd196,8'd240} : s = 436;
	{8'd196,8'd241} : s = 437;
	{8'd196,8'd242} : s = 438;
	{8'd196,8'd243} : s = 439;
	{8'd196,8'd244} : s = 440;
	{8'd196,8'd245} : s = 441;
	{8'd196,8'd246} : s = 442;
	{8'd196,8'd247} : s = 443;
	{8'd196,8'd248} : s = 444;
	{8'd196,8'd249} : s = 445;
	{8'd196,8'd250} : s = 446;
	{8'd196,8'd251} : s = 447;
	{8'd196,8'd252} : s = 448;
	{8'd196,8'd253} : s = 449;
	{8'd196,8'd254} : s = 450;
	{8'd196,8'd255} : s = 451;
	{8'd197,8'd0} : s = 197;
	{8'd197,8'd1} : s = 198;
	{8'd197,8'd2} : s = 199;
	{8'd197,8'd3} : s = 200;
	{8'd197,8'd4} : s = 201;
	{8'd197,8'd5} : s = 202;
	{8'd197,8'd6} : s = 203;
	{8'd197,8'd7} : s = 204;
	{8'd197,8'd8} : s = 205;
	{8'd197,8'd9} : s = 206;
	{8'd197,8'd10} : s = 207;
	{8'd197,8'd11} : s = 208;
	{8'd197,8'd12} : s = 209;
	{8'd197,8'd13} : s = 210;
	{8'd197,8'd14} : s = 211;
	{8'd197,8'd15} : s = 212;
	{8'd197,8'd16} : s = 213;
	{8'd197,8'd17} : s = 214;
	{8'd197,8'd18} : s = 215;
	{8'd197,8'd19} : s = 216;
	{8'd197,8'd20} : s = 217;
	{8'd197,8'd21} : s = 218;
	{8'd197,8'd22} : s = 219;
	{8'd197,8'd23} : s = 220;
	{8'd197,8'd24} : s = 221;
	{8'd197,8'd25} : s = 222;
	{8'd197,8'd26} : s = 223;
	{8'd197,8'd27} : s = 224;
	{8'd197,8'd28} : s = 225;
	{8'd197,8'd29} : s = 226;
	{8'd197,8'd30} : s = 227;
	{8'd197,8'd31} : s = 228;
	{8'd197,8'd32} : s = 229;
	{8'd197,8'd33} : s = 230;
	{8'd197,8'd34} : s = 231;
	{8'd197,8'd35} : s = 232;
	{8'd197,8'd36} : s = 233;
	{8'd197,8'd37} : s = 234;
	{8'd197,8'd38} : s = 235;
	{8'd197,8'd39} : s = 236;
	{8'd197,8'd40} : s = 237;
	{8'd197,8'd41} : s = 238;
	{8'd197,8'd42} : s = 239;
	{8'd197,8'd43} : s = 240;
	{8'd197,8'd44} : s = 241;
	{8'd197,8'd45} : s = 242;
	{8'd197,8'd46} : s = 243;
	{8'd197,8'd47} : s = 244;
	{8'd197,8'd48} : s = 245;
	{8'd197,8'd49} : s = 246;
	{8'd197,8'd50} : s = 247;
	{8'd197,8'd51} : s = 248;
	{8'd197,8'd52} : s = 249;
	{8'd197,8'd53} : s = 250;
	{8'd197,8'd54} : s = 251;
	{8'd197,8'd55} : s = 252;
	{8'd197,8'd56} : s = 253;
	{8'd197,8'd57} : s = 254;
	{8'd197,8'd58} : s = 255;
	{8'd197,8'd59} : s = 256;
	{8'd197,8'd60} : s = 257;
	{8'd197,8'd61} : s = 258;
	{8'd197,8'd62} : s = 259;
	{8'd197,8'd63} : s = 260;
	{8'd197,8'd64} : s = 261;
	{8'd197,8'd65} : s = 262;
	{8'd197,8'd66} : s = 263;
	{8'd197,8'd67} : s = 264;
	{8'd197,8'd68} : s = 265;
	{8'd197,8'd69} : s = 266;
	{8'd197,8'd70} : s = 267;
	{8'd197,8'd71} : s = 268;
	{8'd197,8'd72} : s = 269;
	{8'd197,8'd73} : s = 270;
	{8'd197,8'd74} : s = 271;
	{8'd197,8'd75} : s = 272;
	{8'd197,8'd76} : s = 273;
	{8'd197,8'd77} : s = 274;
	{8'd197,8'd78} : s = 275;
	{8'd197,8'd79} : s = 276;
	{8'd197,8'd80} : s = 277;
	{8'd197,8'd81} : s = 278;
	{8'd197,8'd82} : s = 279;
	{8'd197,8'd83} : s = 280;
	{8'd197,8'd84} : s = 281;
	{8'd197,8'd85} : s = 282;
	{8'd197,8'd86} : s = 283;
	{8'd197,8'd87} : s = 284;
	{8'd197,8'd88} : s = 285;
	{8'd197,8'd89} : s = 286;
	{8'd197,8'd90} : s = 287;
	{8'd197,8'd91} : s = 288;
	{8'd197,8'd92} : s = 289;
	{8'd197,8'd93} : s = 290;
	{8'd197,8'd94} : s = 291;
	{8'd197,8'd95} : s = 292;
	{8'd197,8'd96} : s = 293;
	{8'd197,8'd97} : s = 294;
	{8'd197,8'd98} : s = 295;
	{8'd197,8'd99} : s = 296;
	{8'd197,8'd100} : s = 297;
	{8'd197,8'd101} : s = 298;
	{8'd197,8'd102} : s = 299;
	{8'd197,8'd103} : s = 300;
	{8'd197,8'd104} : s = 301;
	{8'd197,8'd105} : s = 302;
	{8'd197,8'd106} : s = 303;
	{8'd197,8'd107} : s = 304;
	{8'd197,8'd108} : s = 305;
	{8'd197,8'd109} : s = 306;
	{8'd197,8'd110} : s = 307;
	{8'd197,8'd111} : s = 308;
	{8'd197,8'd112} : s = 309;
	{8'd197,8'd113} : s = 310;
	{8'd197,8'd114} : s = 311;
	{8'd197,8'd115} : s = 312;
	{8'd197,8'd116} : s = 313;
	{8'd197,8'd117} : s = 314;
	{8'd197,8'd118} : s = 315;
	{8'd197,8'd119} : s = 316;
	{8'd197,8'd120} : s = 317;
	{8'd197,8'd121} : s = 318;
	{8'd197,8'd122} : s = 319;
	{8'd197,8'd123} : s = 320;
	{8'd197,8'd124} : s = 321;
	{8'd197,8'd125} : s = 322;
	{8'd197,8'd126} : s = 323;
	{8'd197,8'd127} : s = 324;
	{8'd197,8'd128} : s = 325;
	{8'd197,8'd129} : s = 326;
	{8'd197,8'd130} : s = 327;
	{8'd197,8'd131} : s = 328;
	{8'd197,8'd132} : s = 329;
	{8'd197,8'd133} : s = 330;
	{8'd197,8'd134} : s = 331;
	{8'd197,8'd135} : s = 332;
	{8'd197,8'd136} : s = 333;
	{8'd197,8'd137} : s = 334;
	{8'd197,8'd138} : s = 335;
	{8'd197,8'd139} : s = 336;
	{8'd197,8'd140} : s = 337;
	{8'd197,8'd141} : s = 338;
	{8'd197,8'd142} : s = 339;
	{8'd197,8'd143} : s = 340;
	{8'd197,8'd144} : s = 341;
	{8'd197,8'd145} : s = 342;
	{8'd197,8'd146} : s = 343;
	{8'd197,8'd147} : s = 344;
	{8'd197,8'd148} : s = 345;
	{8'd197,8'd149} : s = 346;
	{8'd197,8'd150} : s = 347;
	{8'd197,8'd151} : s = 348;
	{8'd197,8'd152} : s = 349;
	{8'd197,8'd153} : s = 350;
	{8'd197,8'd154} : s = 351;
	{8'd197,8'd155} : s = 352;
	{8'd197,8'd156} : s = 353;
	{8'd197,8'd157} : s = 354;
	{8'd197,8'd158} : s = 355;
	{8'd197,8'd159} : s = 356;
	{8'd197,8'd160} : s = 357;
	{8'd197,8'd161} : s = 358;
	{8'd197,8'd162} : s = 359;
	{8'd197,8'd163} : s = 360;
	{8'd197,8'd164} : s = 361;
	{8'd197,8'd165} : s = 362;
	{8'd197,8'd166} : s = 363;
	{8'd197,8'd167} : s = 364;
	{8'd197,8'd168} : s = 365;
	{8'd197,8'd169} : s = 366;
	{8'd197,8'd170} : s = 367;
	{8'd197,8'd171} : s = 368;
	{8'd197,8'd172} : s = 369;
	{8'd197,8'd173} : s = 370;
	{8'd197,8'd174} : s = 371;
	{8'd197,8'd175} : s = 372;
	{8'd197,8'd176} : s = 373;
	{8'd197,8'd177} : s = 374;
	{8'd197,8'd178} : s = 375;
	{8'd197,8'd179} : s = 376;
	{8'd197,8'd180} : s = 377;
	{8'd197,8'd181} : s = 378;
	{8'd197,8'd182} : s = 379;
	{8'd197,8'd183} : s = 380;
	{8'd197,8'd184} : s = 381;
	{8'd197,8'd185} : s = 382;
	{8'd197,8'd186} : s = 383;
	{8'd197,8'd187} : s = 384;
	{8'd197,8'd188} : s = 385;
	{8'd197,8'd189} : s = 386;
	{8'd197,8'd190} : s = 387;
	{8'd197,8'd191} : s = 388;
	{8'd197,8'd192} : s = 389;
	{8'd197,8'd193} : s = 390;
	{8'd197,8'd194} : s = 391;
	{8'd197,8'd195} : s = 392;
	{8'd197,8'd196} : s = 393;
	{8'd197,8'd197} : s = 394;
	{8'd197,8'd198} : s = 395;
	{8'd197,8'd199} : s = 396;
	{8'd197,8'd200} : s = 397;
	{8'd197,8'd201} : s = 398;
	{8'd197,8'd202} : s = 399;
	{8'd197,8'd203} : s = 400;
	{8'd197,8'd204} : s = 401;
	{8'd197,8'd205} : s = 402;
	{8'd197,8'd206} : s = 403;
	{8'd197,8'd207} : s = 404;
	{8'd197,8'd208} : s = 405;
	{8'd197,8'd209} : s = 406;
	{8'd197,8'd210} : s = 407;
	{8'd197,8'd211} : s = 408;
	{8'd197,8'd212} : s = 409;
	{8'd197,8'd213} : s = 410;
	{8'd197,8'd214} : s = 411;
	{8'd197,8'd215} : s = 412;
	{8'd197,8'd216} : s = 413;
	{8'd197,8'd217} : s = 414;
	{8'd197,8'd218} : s = 415;
	{8'd197,8'd219} : s = 416;
	{8'd197,8'd220} : s = 417;
	{8'd197,8'd221} : s = 418;
	{8'd197,8'd222} : s = 419;
	{8'd197,8'd223} : s = 420;
	{8'd197,8'd224} : s = 421;
	{8'd197,8'd225} : s = 422;
	{8'd197,8'd226} : s = 423;
	{8'd197,8'd227} : s = 424;
	{8'd197,8'd228} : s = 425;
	{8'd197,8'd229} : s = 426;
	{8'd197,8'd230} : s = 427;
	{8'd197,8'd231} : s = 428;
	{8'd197,8'd232} : s = 429;
	{8'd197,8'd233} : s = 430;
	{8'd197,8'd234} : s = 431;
	{8'd197,8'd235} : s = 432;
	{8'd197,8'd236} : s = 433;
	{8'd197,8'd237} : s = 434;
	{8'd197,8'd238} : s = 435;
	{8'd197,8'd239} : s = 436;
	{8'd197,8'd240} : s = 437;
	{8'd197,8'd241} : s = 438;
	{8'd197,8'd242} : s = 439;
	{8'd197,8'd243} : s = 440;
	{8'd197,8'd244} : s = 441;
	{8'd197,8'd245} : s = 442;
	{8'd197,8'd246} : s = 443;
	{8'd197,8'd247} : s = 444;
	{8'd197,8'd248} : s = 445;
	{8'd197,8'd249} : s = 446;
	{8'd197,8'd250} : s = 447;
	{8'd197,8'd251} : s = 448;
	{8'd197,8'd252} : s = 449;
	{8'd197,8'd253} : s = 450;
	{8'd197,8'd254} : s = 451;
	{8'd197,8'd255} : s = 452;
	{8'd198,8'd0} : s = 198;
	{8'd198,8'd1} : s = 199;
	{8'd198,8'd2} : s = 200;
	{8'd198,8'd3} : s = 201;
	{8'd198,8'd4} : s = 202;
	{8'd198,8'd5} : s = 203;
	{8'd198,8'd6} : s = 204;
	{8'd198,8'd7} : s = 205;
	{8'd198,8'd8} : s = 206;
	{8'd198,8'd9} : s = 207;
	{8'd198,8'd10} : s = 208;
	{8'd198,8'd11} : s = 209;
	{8'd198,8'd12} : s = 210;
	{8'd198,8'd13} : s = 211;
	{8'd198,8'd14} : s = 212;
	{8'd198,8'd15} : s = 213;
	{8'd198,8'd16} : s = 214;
	{8'd198,8'd17} : s = 215;
	{8'd198,8'd18} : s = 216;
	{8'd198,8'd19} : s = 217;
	{8'd198,8'd20} : s = 218;
	{8'd198,8'd21} : s = 219;
	{8'd198,8'd22} : s = 220;
	{8'd198,8'd23} : s = 221;
	{8'd198,8'd24} : s = 222;
	{8'd198,8'd25} : s = 223;
	{8'd198,8'd26} : s = 224;
	{8'd198,8'd27} : s = 225;
	{8'd198,8'd28} : s = 226;
	{8'd198,8'd29} : s = 227;
	{8'd198,8'd30} : s = 228;
	{8'd198,8'd31} : s = 229;
	{8'd198,8'd32} : s = 230;
	{8'd198,8'd33} : s = 231;
	{8'd198,8'd34} : s = 232;
	{8'd198,8'd35} : s = 233;
	{8'd198,8'd36} : s = 234;
	{8'd198,8'd37} : s = 235;
	{8'd198,8'd38} : s = 236;
	{8'd198,8'd39} : s = 237;
	{8'd198,8'd40} : s = 238;
	{8'd198,8'd41} : s = 239;
	{8'd198,8'd42} : s = 240;
	{8'd198,8'd43} : s = 241;
	{8'd198,8'd44} : s = 242;
	{8'd198,8'd45} : s = 243;
	{8'd198,8'd46} : s = 244;
	{8'd198,8'd47} : s = 245;
	{8'd198,8'd48} : s = 246;
	{8'd198,8'd49} : s = 247;
	{8'd198,8'd50} : s = 248;
	{8'd198,8'd51} : s = 249;
	{8'd198,8'd52} : s = 250;
	{8'd198,8'd53} : s = 251;
	{8'd198,8'd54} : s = 252;
	{8'd198,8'd55} : s = 253;
	{8'd198,8'd56} : s = 254;
	{8'd198,8'd57} : s = 255;
	{8'd198,8'd58} : s = 256;
	{8'd198,8'd59} : s = 257;
	{8'd198,8'd60} : s = 258;
	{8'd198,8'd61} : s = 259;
	{8'd198,8'd62} : s = 260;
	{8'd198,8'd63} : s = 261;
	{8'd198,8'd64} : s = 262;
	{8'd198,8'd65} : s = 263;
	{8'd198,8'd66} : s = 264;
	{8'd198,8'd67} : s = 265;
	{8'd198,8'd68} : s = 266;
	{8'd198,8'd69} : s = 267;
	{8'd198,8'd70} : s = 268;
	{8'd198,8'd71} : s = 269;
	{8'd198,8'd72} : s = 270;
	{8'd198,8'd73} : s = 271;
	{8'd198,8'd74} : s = 272;
	{8'd198,8'd75} : s = 273;
	{8'd198,8'd76} : s = 274;
	{8'd198,8'd77} : s = 275;
	{8'd198,8'd78} : s = 276;
	{8'd198,8'd79} : s = 277;
	{8'd198,8'd80} : s = 278;
	{8'd198,8'd81} : s = 279;
	{8'd198,8'd82} : s = 280;
	{8'd198,8'd83} : s = 281;
	{8'd198,8'd84} : s = 282;
	{8'd198,8'd85} : s = 283;
	{8'd198,8'd86} : s = 284;
	{8'd198,8'd87} : s = 285;
	{8'd198,8'd88} : s = 286;
	{8'd198,8'd89} : s = 287;
	{8'd198,8'd90} : s = 288;
	{8'd198,8'd91} : s = 289;
	{8'd198,8'd92} : s = 290;
	{8'd198,8'd93} : s = 291;
	{8'd198,8'd94} : s = 292;
	{8'd198,8'd95} : s = 293;
	{8'd198,8'd96} : s = 294;
	{8'd198,8'd97} : s = 295;
	{8'd198,8'd98} : s = 296;
	{8'd198,8'd99} : s = 297;
	{8'd198,8'd100} : s = 298;
	{8'd198,8'd101} : s = 299;
	{8'd198,8'd102} : s = 300;
	{8'd198,8'd103} : s = 301;
	{8'd198,8'd104} : s = 302;
	{8'd198,8'd105} : s = 303;
	{8'd198,8'd106} : s = 304;
	{8'd198,8'd107} : s = 305;
	{8'd198,8'd108} : s = 306;
	{8'd198,8'd109} : s = 307;
	{8'd198,8'd110} : s = 308;
	{8'd198,8'd111} : s = 309;
	{8'd198,8'd112} : s = 310;
	{8'd198,8'd113} : s = 311;
	{8'd198,8'd114} : s = 312;
	{8'd198,8'd115} : s = 313;
	{8'd198,8'd116} : s = 314;
	{8'd198,8'd117} : s = 315;
	{8'd198,8'd118} : s = 316;
	{8'd198,8'd119} : s = 317;
	{8'd198,8'd120} : s = 318;
	{8'd198,8'd121} : s = 319;
	{8'd198,8'd122} : s = 320;
	{8'd198,8'd123} : s = 321;
	{8'd198,8'd124} : s = 322;
	{8'd198,8'd125} : s = 323;
	{8'd198,8'd126} : s = 324;
	{8'd198,8'd127} : s = 325;
	{8'd198,8'd128} : s = 326;
	{8'd198,8'd129} : s = 327;
	{8'd198,8'd130} : s = 328;
	{8'd198,8'd131} : s = 329;
	{8'd198,8'd132} : s = 330;
	{8'd198,8'd133} : s = 331;
	{8'd198,8'd134} : s = 332;
	{8'd198,8'd135} : s = 333;
	{8'd198,8'd136} : s = 334;
	{8'd198,8'd137} : s = 335;
	{8'd198,8'd138} : s = 336;
	{8'd198,8'd139} : s = 337;
	{8'd198,8'd140} : s = 338;
	{8'd198,8'd141} : s = 339;
	{8'd198,8'd142} : s = 340;
	{8'd198,8'd143} : s = 341;
	{8'd198,8'd144} : s = 342;
	{8'd198,8'd145} : s = 343;
	{8'd198,8'd146} : s = 344;
	{8'd198,8'd147} : s = 345;
	{8'd198,8'd148} : s = 346;
	{8'd198,8'd149} : s = 347;
	{8'd198,8'd150} : s = 348;
	{8'd198,8'd151} : s = 349;
	{8'd198,8'd152} : s = 350;
	{8'd198,8'd153} : s = 351;
	{8'd198,8'd154} : s = 352;
	{8'd198,8'd155} : s = 353;
	{8'd198,8'd156} : s = 354;
	{8'd198,8'd157} : s = 355;
	{8'd198,8'd158} : s = 356;
	{8'd198,8'd159} : s = 357;
	{8'd198,8'd160} : s = 358;
	{8'd198,8'd161} : s = 359;
	{8'd198,8'd162} : s = 360;
	{8'd198,8'd163} : s = 361;
	{8'd198,8'd164} : s = 362;
	{8'd198,8'd165} : s = 363;
	{8'd198,8'd166} : s = 364;
	{8'd198,8'd167} : s = 365;
	{8'd198,8'd168} : s = 366;
	{8'd198,8'd169} : s = 367;
	{8'd198,8'd170} : s = 368;
	{8'd198,8'd171} : s = 369;
	{8'd198,8'd172} : s = 370;
	{8'd198,8'd173} : s = 371;
	{8'd198,8'd174} : s = 372;
	{8'd198,8'd175} : s = 373;
	{8'd198,8'd176} : s = 374;
	{8'd198,8'd177} : s = 375;
	{8'd198,8'd178} : s = 376;
	{8'd198,8'd179} : s = 377;
	{8'd198,8'd180} : s = 378;
	{8'd198,8'd181} : s = 379;
	{8'd198,8'd182} : s = 380;
	{8'd198,8'd183} : s = 381;
	{8'd198,8'd184} : s = 382;
	{8'd198,8'd185} : s = 383;
	{8'd198,8'd186} : s = 384;
	{8'd198,8'd187} : s = 385;
	{8'd198,8'd188} : s = 386;
	{8'd198,8'd189} : s = 387;
	{8'd198,8'd190} : s = 388;
	{8'd198,8'd191} : s = 389;
	{8'd198,8'd192} : s = 390;
	{8'd198,8'd193} : s = 391;
	{8'd198,8'd194} : s = 392;
	{8'd198,8'd195} : s = 393;
	{8'd198,8'd196} : s = 394;
	{8'd198,8'd197} : s = 395;
	{8'd198,8'd198} : s = 396;
	{8'd198,8'd199} : s = 397;
	{8'd198,8'd200} : s = 398;
	{8'd198,8'd201} : s = 399;
	{8'd198,8'd202} : s = 400;
	{8'd198,8'd203} : s = 401;
	{8'd198,8'd204} : s = 402;
	{8'd198,8'd205} : s = 403;
	{8'd198,8'd206} : s = 404;
	{8'd198,8'd207} : s = 405;
	{8'd198,8'd208} : s = 406;
	{8'd198,8'd209} : s = 407;
	{8'd198,8'd210} : s = 408;
	{8'd198,8'd211} : s = 409;
	{8'd198,8'd212} : s = 410;
	{8'd198,8'd213} : s = 411;
	{8'd198,8'd214} : s = 412;
	{8'd198,8'd215} : s = 413;
	{8'd198,8'd216} : s = 414;
	{8'd198,8'd217} : s = 415;
	{8'd198,8'd218} : s = 416;
	{8'd198,8'd219} : s = 417;
	{8'd198,8'd220} : s = 418;
	{8'd198,8'd221} : s = 419;
	{8'd198,8'd222} : s = 420;
	{8'd198,8'd223} : s = 421;
	{8'd198,8'd224} : s = 422;
	{8'd198,8'd225} : s = 423;
	{8'd198,8'd226} : s = 424;
	{8'd198,8'd227} : s = 425;
	{8'd198,8'd228} : s = 426;
	{8'd198,8'd229} : s = 427;
	{8'd198,8'd230} : s = 428;
	{8'd198,8'd231} : s = 429;
	{8'd198,8'd232} : s = 430;
	{8'd198,8'd233} : s = 431;
	{8'd198,8'd234} : s = 432;
	{8'd198,8'd235} : s = 433;
	{8'd198,8'd236} : s = 434;
	{8'd198,8'd237} : s = 435;
	{8'd198,8'd238} : s = 436;
	{8'd198,8'd239} : s = 437;
	{8'd198,8'd240} : s = 438;
	{8'd198,8'd241} : s = 439;
	{8'd198,8'd242} : s = 440;
	{8'd198,8'd243} : s = 441;
	{8'd198,8'd244} : s = 442;
	{8'd198,8'd245} : s = 443;
	{8'd198,8'd246} : s = 444;
	{8'd198,8'd247} : s = 445;
	{8'd198,8'd248} : s = 446;
	{8'd198,8'd249} : s = 447;
	{8'd198,8'd250} : s = 448;
	{8'd198,8'd251} : s = 449;
	{8'd198,8'd252} : s = 450;
	{8'd198,8'd253} : s = 451;
	{8'd198,8'd254} : s = 452;
	{8'd198,8'd255} : s = 453;
	{8'd199,8'd0} : s = 199;
	{8'd199,8'd1} : s = 200;
	{8'd199,8'd2} : s = 201;
	{8'd199,8'd3} : s = 202;
	{8'd199,8'd4} : s = 203;
	{8'd199,8'd5} : s = 204;
	{8'd199,8'd6} : s = 205;
	{8'd199,8'd7} : s = 206;
	{8'd199,8'd8} : s = 207;
	{8'd199,8'd9} : s = 208;
	{8'd199,8'd10} : s = 209;
	{8'd199,8'd11} : s = 210;
	{8'd199,8'd12} : s = 211;
	{8'd199,8'd13} : s = 212;
	{8'd199,8'd14} : s = 213;
	{8'd199,8'd15} : s = 214;
	{8'd199,8'd16} : s = 215;
	{8'd199,8'd17} : s = 216;
	{8'd199,8'd18} : s = 217;
	{8'd199,8'd19} : s = 218;
	{8'd199,8'd20} : s = 219;
	{8'd199,8'd21} : s = 220;
	{8'd199,8'd22} : s = 221;
	{8'd199,8'd23} : s = 222;
	{8'd199,8'd24} : s = 223;
	{8'd199,8'd25} : s = 224;
	{8'd199,8'd26} : s = 225;
	{8'd199,8'd27} : s = 226;
	{8'd199,8'd28} : s = 227;
	{8'd199,8'd29} : s = 228;
	{8'd199,8'd30} : s = 229;
	{8'd199,8'd31} : s = 230;
	{8'd199,8'd32} : s = 231;
	{8'd199,8'd33} : s = 232;
	{8'd199,8'd34} : s = 233;
	{8'd199,8'd35} : s = 234;
	{8'd199,8'd36} : s = 235;
	{8'd199,8'd37} : s = 236;
	{8'd199,8'd38} : s = 237;
	{8'd199,8'd39} : s = 238;
	{8'd199,8'd40} : s = 239;
	{8'd199,8'd41} : s = 240;
	{8'd199,8'd42} : s = 241;
	{8'd199,8'd43} : s = 242;
	{8'd199,8'd44} : s = 243;
	{8'd199,8'd45} : s = 244;
	{8'd199,8'd46} : s = 245;
	{8'd199,8'd47} : s = 246;
	{8'd199,8'd48} : s = 247;
	{8'd199,8'd49} : s = 248;
	{8'd199,8'd50} : s = 249;
	{8'd199,8'd51} : s = 250;
	{8'd199,8'd52} : s = 251;
	{8'd199,8'd53} : s = 252;
	{8'd199,8'd54} : s = 253;
	{8'd199,8'd55} : s = 254;
	{8'd199,8'd56} : s = 255;
	{8'd199,8'd57} : s = 256;
	{8'd199,8'd58} : s = 257;
	{8'd199,8'd59} : s = 258;
	{8'd199,8'd60} : s = 259;
	{8'd199,8'd61} : s = 260;
	{8'd199,8'd62} : s = 261;
	{8'd199,8'd63} : s = 262;
	{8'd199,8'd64} : s = 263;
	{8'd199,8'd65} : s = 264;
	{8'd199,8'd66} : s = 265;
	{8'd199,8'd67} : s = 266;
	{8'd199,8'd68} : s = 267;
	{8'd199,8'd69} : s = 268;
	{8'd199,8'd70} : s = 269;
	{8'd199,8'd71} : s = 270;
	{8'd199,8'd72} : s = 271;
	{8'd199,8'd73} : s = 272;
	{8'd199,8'd74} : s = 273;
	{8'd199,8'd75} : s = 274;
	{8'd199,8'd76} : s = 275;
	{8'd199,8'd77} : s = 276;
	{8'd199,8'd78} : s = 277;
	{8'd199,8'd79} : s = 278;
	{8'd199,8'd80} : s = 279;
	{8'd199,8'd81} : s = 280;
	{8'd199,8'd82} : s = 281;
	{8'd199,8'd83} : s = 282;
	{8'd199,8'd84} : s = 283;
	{8'd199,8'd85} : s = 284;
	{8'd199,8'd86} : s = 285;
	{8'd199,8'd87} : s = 286;
	{8'd199,8'd88} : s = 287;
	{8'd199,8'd89} : s = 288;
	{8'd199,8'd90} : s = 289;
	{8'd199,8'd91} : s = 290;
	{8'd199,8'd92} : s = 291;
	{8'd199,8'd93} : s = 292;
	{8'd199,8'd94} : s = 293;
	{8'd199,8'd95} : s = 294;
	{8'd199,8'd96} : s = 295;
	{8'd199,8'd97} : s = 296;
	{8'd199,8'd98} : s = 297;
	{8'd199,8'd99} : s = 298;
	{8'd199,8'd100} : s = 299;
	{8'd199,8'd101} : s = 300;
	{8'd199,8'd102} : s = 301;
	{8'd199,8'd103} : s = 302;
	{8'd199,8'd104} : s = 303;
	{8'd199,8'd105} : s = 304;
	{8'd199,8'd106} : s = 305;
	{8'd199,8'd107} : s = 306;
	{8'd199,8'd108} : s = 307;
	{8'd199,8'd109} : s = 308;
	{8'd199,8'd110} : s = 309;
	{8'd199,8'd111} : s = 310;
	{8'd199,8'd112} : s = 311;
	{8'd199,8'd113} : s = 312;
	{8'd199,8'd114} : s = 313;
	{8'd199,8'd115} : s = 314;
	{8'd199,8'd116} : s = 315;
	{8'd199,8'd117} : s = 316;
	{8'd199,8'd118} : s = 317;
	{8'd199,8'd119} : s = 318;
	{8'd199,8'd120} : s = 319;
	{8'd199,8'd121} : s = 320;
	{8'd199,8'd122} : s = 321;
	{8'd199,8'd123} : s = 322;
	{8'd199,8'd124} : s = 323;
	{8'd199,8'd125} : s = 324;
	{8'd199,8'd126} : s = 325;
	{8'd199,8'd127} : s = 326;
	{8'd199,8'd128} : s = 327;
	{8'd199,8'd129} : s = 328;
	{8'd199,8'd130} : s = 329;
	{8'd199,8'd131} : s = 330;
	{8'd199,8'd132} : s = 331;
	{8'd199,8'd133} : s = 332;
	{8'd199,8'd134} : s = 333;
	{8'd199,8'd135} : s = 334;
	{8'd199,8'd136} : s = 335;
	{8'd199,8'd137} : s = 336;
	{8'd199,8'd138} : s = 337;
	{8'd199,8'd139} : s = 338;
	{8'd199,8'd140} : s = 339;
	{8'd199,8'd141} : s = 340;
	{8'd199,8'd142} : s = 341;
	{8'd199,8'd143} : s = 342;
	{8'd199,8'd144} : s = 343;
	{8'd199,8'd145} : s = 344;
	{8'd199,8'd146} : s = 345;
	{8'd199,8'd147} : s = 346;
	{8'd199,8'd148} : s = 347;
	{8'd199,8'd149} : s = 348;
	{8'd199,8'd150} : s = 349;
	{8'd199,8'd151} : s = 350;
	{8'd199,8'd152} : s = 351;
	{8'd199,8'd153} : s = 352;
	{8'd199,8'd154} : s = 353;
	{8'd199,8'd155} : s = 354;
	{8'd199,8'd156} : s = 355;
	{8'd199,8'd157} : s = 356;
	{8'd199,8'd158} : s = 357;
	{8'd199,8'd159} : s = 358;
	{8'd199,8'd160} : s = 359;
	{8'd199,8'd161} : s = 360;
	{8'd199,8'd162} : s = 361;
	{8'd199,8'd163} : s = 362;
	{8'd199,8'd164} : s = 363;
	{8'd199,8'd165} : s = 364;
	{8'd199,8'd166} : s = 365;
	{8'd199,8'd167} : s = 366;
	{8'd199,8'd168} : s = 367;
	{8'd199,8'd169} : s = 368;
	{8'd199,8'd170} : s = 369;
	{8'd199,8'd171} : s = 370;
	{8'd199,8'd172} : s = 371;
	{8'd199,8'd173} : s = 372;
	{8'd199,8'd174} : s = 373;
	{8'd199,8'd175} : s = 374;
	{8'd199,8'd176} : s = 375;
	{8'd199,8'd177} : s = 376;
	{8'd199,8'd178} : s = 377;
	{8'd199,8'd179} : s = 378;
	{8'd199,8'd180} : s = 379;
	{8'd199,8'd181} : s = 380;
	{8'd199,8'd182} : s = 381;
	{8'd199,8'd183} : s = 382;
	{8'd199,8'd184} : s = 383;
	{8'd199,8'd185} : s = 384;
	{8'd199,8'd186} : s = 385;
	{8'd199,8'd187} : s = 386;
	{8'd199,8'd188} : s = 387;
	{8'd199,8'd189} : s = 388;
	{8'd199,8'd190} : s = 389;
	{8'd199,8'd191} : s = 390;
	{8'd199,8'd192} : s = 391;
	{8'd199,8'd193} : s = 392;
	{8'd199,8'd194} : s = 393;
	{8'd199,8'd195} : s = 394;
	{8'd199,8'd196} : s = 395;
	{8'd199,8'd197} : s = 396;
	{8'd199,8'd198} : s = 397;
	{8'd199,8'd199} : s = 398;
	{8'd199,8'd200} : s = 399;
	{8'd199,8'd201} : s = 400;
	{8'd199,8'd202} : s = 401;
	{8'd199,8'd203} : s = 402;
	{8'd199,8'd204} : s = 403;
	{8'd199,8'd205} : s = 404;
	{8'd199,8'd206} : s = 405;
	{8'd199,8'd207} : s = 406;
	{8'd199,8'd208} : s = 407;
	{8'd199,8'd209} : s = 408;
	{8'd199,8'd210} : s = 409;
	{8'd199,8'd211} : s = 410;
	{8'd199,8'd212} : s = 411;
	{8'd199,8'd213} : s = 412;
	{8'd199,8'd214} : s = 413;
	{8'd199,8'd215} : s = 414;
	{8'd199,8'd216} : s = 415;
	{8'd199,8'd217} : s = 416;
	{8'd199,8'd218} : s = 417;
	{8'd199,8'd219} : s = 418;
	{8'd199,8'd220} : s = 419;
	{8'd199,8'd221} : s = 420;
	{8'd199,8'd222} : s = 421;
	{8'd199,8'd223} : s = 422;
	{8'd199,8'd224} : s = 423;
	{8'd199,8'd225} : s = 424;
	{8'd199,8'd226} : s = 425;
	{8'd199,8'd227} : s = 426;
	{8'd199,8'd228} : s = 427;
	{8'd199,8'd229} : s = 428;
	{8'd199,8'd230} : s = 429;
	{8'd199,8'd231} : s = 430;
	{8'd199,8'd232} : s = 431;
	{8'd199,8'd233} : s = 432;
	{8'd199,8'd234} : s = 433;
	{8'd199,8'd235} : s = 434;
	{8'd199,8'd236} : s = 435;
	{8'd199,8'd237} : s = 436;
	{8'd199,8'd238} : s = 437;
	{8'd199,8'd239} : s = 438;
	{8'd199,8'd240} : s = 439;
	{8'd199,8'd241} : s = 440;
	{8'd199,8'd242} : s = 441;
	{8'd199,8'd243} : s = 442;
	{8'd199,8'd244} : s = 443;
	{8'd199,8'd245} : s = 444;
	{8'd199,8'd246} : s = 445;
	{8'd199,8'd247} : s = 446;
	{8'd199,8'd248} : s = 447;
	{8'd199,8'd249} : s = 448;
	{8'd199,8'd250} : s = 449;
	{8'd199,8'd251} : s = 450;
	{8'd199,8'd252} : s = 451;
	{8'd199,8'd253} : s = 452;
	{8'd199,8'd254} : s = 453;
	{8'd199,8'd255} : s = 454;
	{8'd200,8'd0} : s = 200;
	{8'd200,8'd1} : s = 201;
	{8'd200,8'd2} : s = 202;
	{8'd200,8'd3} : s = 203;
	{8'd200,8'd4} : s = 204;
	{8'd200,8'd5} : s = 205;
	{8'd200,8'd6} : s = 206;
	{8'd200,8'd7} : s = 207;
	{8'd200,8'd8} : s = 208;
	{8'd200,8'd9} : s = 209;
	{8'd200,8'd10} : s = 210;
	{8'd200,8'd11} : s = 211;
	{8'd200,8'd12} : s = 212;
	{8'd200,8'd13} : s = 213;
	{8'd200,8'd14} : s = 214;
	{8'd200,8'd15} : s = 215;
	{8'd200,8'd16} : s = 216;
	{8'd200,8'd17} : s = 217;
	{8'd200,8'd18} : s = 218;
	{8'd200,8'd19} : s = 219;
	{8'd200,8'd20} : s = 220;
	{8'd200,8'd21} : s = 221;
	{8'd200,8'd22} : s = 222;
	{8'd200,8'd23} : s = 223;
	{8'd200,8'd24} : s = 224;
	{8'd200,8'd25} : s = 225;
	{8'd200,8'd26} : s = 226;
	{8'd200,8'd27} : s = 227;
	{8'd200,8'd28} : s = 228;
	{8'd200,8'd29} : s = 229;
	{8'd200,8'd30} : s = 230;
	{8'd200,8'd31} : s = 231;
	{8'd200,8'd32} : s = 232;
	{8'd200,8'd33} : s = 233;
	{8'd200,8'd34} : s = 234;
	{8'd200,8'd35} : s = 235;
	{8'd200,8'd36} : s = 236;
	{8'd200,8'd37} : s = 237;
	{8'd200,8'd38} : s = 238;
	{8'd200,8'd39} : s = 239;
	{8'd200,8'd40} : s = 240;
	{8'd200,8'd41} : s = 241;
	{8'd200,8'd42} : s = 242;
	{8'd200,8'd43} : s = 243;
	{8'd200,8'd44} : s = 244;
	{8'd200,8'd45} : s = 245;
	{8'd200,8'd46} : s = 246;
	{8'd200,8'd47} : s = 247;
	{8'd200,8'd48} : s = 248;
	{8'd200,8'd49} : s = 249;
	{8'd200,8'd50} : s = 250;
	{8'd200,8'd51} : s = 251;
	{8'd200,8'd52} : s = 252;
	{8'd200,8'd53} : s = 253;
	{8'd200,8'd54} : s = 254;
	{8'd200,8'd55} : s = 255;
	{8'd200,8'd56} : s = 256;
	{8'd200,8'd57} : s = 257;
	{8'd200,8'd58} : s = 258;
	{8'd200,8'd59} : s = 259;
	{8'd200,8'd60} : s = 260;
	{8'd200,8'd61} : s = 261;
	{8'd200,8'd62} : s = 262;
	{8'd200,8'd63} : s = 263;
	{8'd200,8'd64} : s = 264;
	{8'd200,8'd65} : s = 265;
	{8'd200,8'd66} : s = 266;
	{8'd200,8'd67} : s = 267;
	{8'd200,8'd68} : s = 268;
	{8'd200,8'd69} : s = 269;
	{8'd200,8'd70} : s = 270;
	{8'd200,8'd71} : s = 271;
	{8'd200,8'd72} : s = 272;
	{8'd200,8'd73} : s = 273;
	{8'd200,8'd74} : s = 274;
	{8'd200,8'd75} : s = 275;
	{8'd200,8'd76} : s = 276;
	{8'd200,8'd77} : s = 277;
	{8'd200,8'd78} : s = 278;
	{8'd200,8'd79} : s = 279;
	{8'd200,8'd80} : s = 280;
	{8'd200,8'd81} : s = 281;
	{8'd200,8'd82} : s = 282;
	{8'd200,8'd83} : s = 283;
	{8'd200,8'd84} : s = 284;
	{8'd200,8'd85} : s = 285;
	{8'd200,8'd86} : s = 286;
	{8'd200,8'd87} : s = 287;
	{8'd200,8'd88} : s = 288;
	{8'd200,8'd89} : s = 289;
	{8'd200,8'd90} : s = 290;
	{8'd200,8'd91} : s = 291;
	{8'd200,8'd92} : s = 292;
	{8'd200,8'd93} : s = 293;
	{8'd200,8'd94} : s = 294;
	{8'd200,8'd95} : s = 295;
	{8'd200,8'd96} : s = 296;
	{8'd200,8'd97} : s = 297;
	{8'd200,8'd98} : s = 298;
	{8'd200,8'd99} : s = 299;
	{8'd200,8'd100} : s = 300;
	{8'd200,8'd101} : s = 301;
	{8'd200,8'd102} : s = 302;
	{8'd200,8'd103} : s = 303;
	{8'd200,8'd104} : s = 304;
	{8'd200,8'd105} : s = 305;
	{8'd200,8'd106} : s = 306;
	{8'd200,8'd107} : s = 307;
	{8'd200,8'd108} : s = 308;
	{8'd200,8'd109} : s = 309;
	{8'd200,8'd110} : s = 310;
	{8'd200,8'd111} : s = 311;
	{8'd200,8'd112} : s = 312;
	{8'd200,8'd113} : s = 313;
	{8'd200,8'd114} : s = 314;
	{8'd200,8'd115} : s = 315;
	{8'd200,8'd116} : s = 316;
	{8'd200,8'd117} : s = 317;
	{8'd200,8'd118} : s = 318;
	{8'd200,8'd119} : s = 319;
	{8'd200,8'd120} : s = 320;
	{8'd200,8'd121} : s = 321;
	{8'd200,8'd122} : s = 322;
	{8'd200,8'd123} : s = 323;
	{8'd200,8'd124} : s = 324;
	{8'd200,8'd125} : s = 325;
	{8'd200,8'd126} : s = 326;
	{8'd200,8'd127} : s = 327;
	{8'd200,8'd128} : s = 328;
	{8'd200,8'd129} : s = 329;
	{8'd200,8'd130} : s = 330;
	{8'd200,8'd131} : s = 331;
	{8'd200,8'd132} : s = 332;
	{8'd200,8'd133} : s = 333;
	{8'd200,8'd134} : s = 334;
	{8'd200,8'd135} : s = 335;
	{8'd200,8'd136} : s = 336;
	{8'd200,8'd137} : s = 337;
	{8'd200,8'd138} : s = 338;
	{8'd200,8'd139} : s = 339;
	{8'd200,8'd140} : s = 340;
	{8'd200,8'd141} : s = 341;
	{8'd200,8'd142} : s = 342;
	{8'd200,8'd143} : s = 343;
	{8'd200,8'd144} : s = 344;
	{8'd200,8'd145} : s = 345;
	{8'd200,8'd146} : s = 346;
	{8'd200,8'd147} : s = 347;
	{8'd200,8'd148} : s = 348;
	{8'd200,8'd149} : s = 349;
	{8'd200,8'd150} : s = 350;
	{8'd200,8'd151} : s = 351;
	{8'd200,8'd152} : s = 352;
	{8'd200,8'd153} : s = 353;
	{8'd200,8'd154} : s = 354;
	{8'd200,8'd155} : s = 355;
	{8'd200,8'd156} : s = 356;
	{8'd200,8'd157} : s = 357;
	{8'd200,8'd158} : s = 358;
	{8'd200,8'd159} : s = 359;
	{8'd200,8'd160} : s = 360;
	{8'd200,8'd161} : s = 361;
	{8'd200,8'd162} : s = 362;
	{8'd200,8'd163} : s = 363;
	{8'd200,8'd164} : s = 364;
	{8'd200,8'd165} : s = 365;
	{8'd200,8'd166} : s = 366;
	{8'd200,8'd167} : s = 367;
	{8'd200,8'd168} : s = 368;
	{8'd200,8'd169} : s = 369;
	{8'd200,8'd170} : s = 370;
	{8'd200,8'd171} : s = 371;
	{8'd200,8'd172} : s = 372;
	{8'd200,8'd173} : s = 373;
	{8'd200,8'd174} : s = 374;
	{8'd200,8'd175} : s = 375;
	{8'd200,8'd176} : s = 376;
	{8'd200,8'd177} : s = 377;
	{8'd200,8'd178} : s = 378;
	{8'd200,8'd179} : s = 379;
	{8'd200,8'd180} : s = 380;
	{8'd200,8'd181} : s = 381;
	{8'd200,8'd182} : s = 382;
	{8'd200,8'd183} : s = 383;
	{8'd200,8'd184} : s = 384;
	{8'd200,8'd185} : s = 385;
	{8'd200,8'd186} : s = 386;
	{8'd200,8'd187} : s = 387;
	{8'd200,8'd188} : s = 388;
	{8'd200,8'd189} : s = 389;
	{8'd200,8'd190} : s = 390;
	{8'd200,8'd191} : s = 391;
	{8'd200,8'd192} : s = 392;
	{8'd200,8'd193} : s = 393;
	{8'd200,8'd194} : s = 394;
	{8'd200,8'd195} : s = 395;
	{8'd200,8'd196} : s = 396;
	{8'd200,8'd197} : s = 397;
	{8'd200,8'd198} : s = 398;
	{8'd200,8'd199} : s = 399;
	{8'd200,8'd200} : s = 400;
	{8'd200,8'd201} : s = 401;
	{8'd200,8'd202} : s = 402;
	{8'd200,8'd203} : s = 403;
	{8'd200,8'd204} : s = 404;
	{8'd200,8'd205} : s = 405;
	{8'd200,8'd206} : s = 406;
	{8'd200,8'd207} : s = 407;
	{8'd200,8'd208} : s = 408;
	{8'd200,8'd209} : s = 409;
	{8'd200,8'd210} : s = 410;
	{8'd200,8'd211} : s = 411;
	{8'd200,8'd212} : s = 412;
	{8'd200,8'd213} : s = 413;
	{8'd200,8'd214} : s = 414;
	{8'd200,8'd215} : s = 415;
	{8'd200,8'd216} : s = 416;
	{8'd200,8'd217} : s = 417;
	{8'd200,8'd218} : s = 418;
	{8'd200,8'd219} : s = 419;
	{8'd200,8'd220} : s = 420;
	{8'd200,8'd221} : s = 421;
	{8'd200,8'd222} : s = 422;
	{8'd200,8'd223} : s = 423;
	{8'd200,8'd224} : s = 424;
	{8'd200,8'd225} : s = 425;
	{8'd200,8'd226} : s = 426;
	{8'd200,8'd227} : s = 427;
	{8'd200,8'd228} : s = 428;
	{8'd200,8'd229} : s = 429;
	{8'd200,8'd230} : s = 430;
	{8'd200,8'd231} : s = 431;
	{8'd200,8'd232} : s = 432;
	{8'd200,8'd233} : s = 433;
	{8'd200,8'd234} : s = 434;
	{8'd200,8'd235} : s = 435;
	{8'd200,8'd236} : s = 436;
	{8'd200,8'd237} : s = 437;
	{8'd200,8'd238} : s = 438;
	{8'd200,8'd239} : s = 439;
	{8'd200,8'd240} : s = 440;
	{8'd200,8'd241} : s = 441;
	{8'd200,8'd242} : s = 442;
	{8'd200,8'd243} : s = 443;
	{8'd200,8'd244} : s = 444;
	{8'd200,8'd245} : s = 445;
	{8'd200,8'd246} : s = 446;
	{8'd200,8'd247} : s = 447;
	{8'd200,8'd248} : s = 448;
	{8'd200,8'd249} : s = 449;
	{8'd200,8'd250} : s = 450;
	{8'd200,8'd251} : s = 451;
	{8'd200,8'd252} : s = 452;
	{8'd200,8'd253} : s = 453;
	{8'd200,8'd254} : s = 454;
	{8'd200,8'd255} : s = 455;
	{8'd201,8'd0} : s = 201;
	{8'd201,8'd1} : s = 202;
	{8'd201,8'd2} : s = 203;
	{8'd201,8'd3} : s = 204;
	{8'd201,8'd4} : s = 205;
	{8'd201,8'd5} : s = 206;
	{8'd201,8'd6} : s = 207;
	{8'd201,8'd7} : s = 208;
	{8'd201,8'd8} : s = 209;
	{8'd201,8'd9} : s = 210;
	{8'd201,8'd10} : s = 211;
	{8'd201,8'd11} : s = 212;
	{8'd201,8'd12} : s = 213;
	{8'd201,8'd13} : s = 214;
	{8'd201,8'd14} : s = 215;
	{8'd201,8'd15} : s = 216;
	{8'd201,8'd16} : s = 217;
	{8'd201,8'd17} : s = 218;
	{8'd201,8'd18} : s = 219;
	{8'd201,8'd19} : s = 220;
	{8'd201,8'd20} : s = 221;
	{8'd201,8'd21} : s = 222;
	{8'd201,8'd22} : s = 223;
	{8'd201,8'd23} : s = 224;
	{8'd201,8'd24} : s = 225;
	{8'd201,8'd25} : s = 226;
	{8'd201,8'd26} : s = 227;
	{8'd201,8'd27} : s = 228;
	{8'd201,8'd28} : s = 229;
	{8'd201,8'd29} : s = 230;
	{8'd201,8'd30} : s = 231;
	{8'd201,8'd31} : s = 232;
	{8'd201,8'd32} : s = 233;
	{8'd201,8'd33} : s = 234;
	{8'd201,8'd34} : s = 235;
	{8'd201,8'd35} : s = 236;
	{8'd201,8'd36} : s = 237;
	{8'd201,8'd37} : s = 238;
	{8'd201,8'd38} : s = 239;
	{8'd201,8'd39} : s = 240;
	{8'd201,8'd40} : s = 241;
	{8'd201,8'd41} : s = 242;
	{8'd201,8'd42} : s = 243;
	{8'd201,8'd43} : s = 244;
	{8'd201,8'd44} : s = 245;
	{8'd201,8'd45} : s = 246;
	{8'd201,8'd46} : s = 247;
	{8'd201,8'd47} : s = 248;
	{8'd201,8'd48} : s = 249;
	{8'd201,8'd49} : s = 250;
	{8'd201,8'd50} : s = 251;
	{8'd201,8'd51} : s = 252;
	{8'd201,8'd52} : s = 253;
	{8'd201,8'd53} : s = 254;
	{8'd201,8'd54} : s = 255;
	{8'd201,8'd55} : s = 256;
	{8'd201,8'd56} : s = 257;
	{8'd201,8'd57} : s = 258;
	{8'd201,8'd58} : s = 259;
	{8'd201,8'd59} : s = 260;
	{8'd201,8'd60} : s = 261;
	{8'd201,8'd61} : s = 262;
	{8'd201,8'd62} : s = 263;
	{8'd201,8'd63} : s = 264;
	{8'd201,8'd64} : s = 265;
	{8'd201,8'd65} : s = 266;
	{8'd201,8'd66} : s = 267;
	{8'd201,8'd67} : s = 268;
	{8'd201,8'd68} : s = 269;
	{8'd201,8'd69} : s = 270;
	{8'd201,8'd70} : s = 271;
	{8'd201,8'd71} : s = 272;
	{8'd201,8'd72} : s = 273;
	{8'd201,8'd73} : s = 274;
	{8'd201,8'd74} : s = 275;
	{8'd201,8'd75} : s = 276;
	{8'd201,8'd76} : s = 277;
	{8'd201,8'd77} : s = 278;
	{8'd201,8'd78} : s = 279;
	{8'd201,8'd79} : s = 280;
	{8'd201,8'd80} : s = 281;
	{8'd201,8'd81} : s = 282;
	{8'd201,8'd82} : s = 283;
	{8'd201,8'd83} : s = 284;
	{8'd201,8'd84} : s = 285;
	{8'd201,8'd85} : s = 286;
	{8'd201,8'd86} : s = 287;
	{8'd201,8'd87} : s = 288;
	{8'd201,8'd88} : s = 289;
	{8'd201,8'd89} : s = 290;
	{8'd201,8'd90} : s = 291;
	{8'd201,8'd91} : s = 292;
	{8'd201,8'd92} : s = 293;
	{8'd201,8'd93} : s = 294;
	{8'd201,8'd94} : s = 295;
	{8'd201,8'd95} : s = 296;
	{8'd201,8'd96} : s = 297;
	{8'd201,8'd97} : s = 298;
	{8'd201,8'd98} : s = 299;
	{8'd201,8'd99} : s = 300;
	{8'd201,8'd100} : s = 301;
	{8'd201,8'd101} : s = 302;
	{8'd201,8'd102} : s = 303;
	{8'd201,8'd103} : s = 304;
	{8'd201,8'd104} : s = 305;
	{8'd201,8'd105} : s = 306;
	{8'd201,8'd106} : s = 307;
	{8'd201,8'd107} : s = 308;
	{8'd201,8'd108} : s = 309;
	{8'd201,8'd109} : s = 310;
	{8'd201,8'd110} : s = 311;
	{8'd201,8'd111} : s = 312;
	{8'd201,8'd112} : s = 313;
	{8'd201,8'd113} : s = 314;
	{8'd201,8'd114} : s = 315;
	{8'd201,8'd115} : s = 316;
	{8'd201,8'd116} : s = 317;
	{8'd201,8'd117} : s = 318;
	{8'd201,8'd118} : s = 319;
	{8'd201,8'd119} : s = 320;
	{8'd201,8'd120} : s = 321;
	{8'd201,8'd121} : s = 322;
	{8'd201,8'd122} : s = 323;
	{8'd201,8'd123} : s = 324;
	{8'd201,8'd124} : s = 325;
	{8'd201,8'd125} : s = 326;
	{8'd201,8'd126} : s = 327;
	{8'd201,8'd127} : s = 328;
	{8'd201,8'd128} : s = 329;
	{8'd201,8'd129} : s = 330;
	{8'd201,8'd130} : s = 331;
	{8'd201,8'd131} : s = 332;
	{8'd201,8'd132} : s = 333;
	{8'd201,8'd133} : s = 334;
	{8'd201,8'd134} : s = 335;
	{8'd201,8'd135} : s = 336;
	{8'd201,8'd136} : s = 337;
	{8'd201,8'd137} : s = 338;
	{8'd201,8'd138} : s = 339;
	{8'd201,8'd139} : s = 340;
	{8'd201,8'd140} : s = 341;
	{8'd201,8'd141} : s = 342;
	{8'd201,8'd142} : s = 343;
	{8'd201,8'd143} : s = 344;
	{8'd201,8'd144} : s = 345;
	{8'd201,8'd145} : s = 346;
	{8'd201,8'd146} : s = 347;
	{8'd201,8'd147} : s = 348;
	{8'd201,8'd148} : s = 349;
	{8'd201,8'd149} : s = 350;
	{8'd201,8'd150} : s = 351;
	{8'd201,8'd151} : s = 352;
	{8'd201,8'd152} : s = 353;
	{8'd201,8'd153} : s = 354;
	{8'd201,8'd154} : s = 355;
	{8'd201,8'd155} : s = 356;
	{8'd201,8'd156} : s = 357;
	{8'd201,8'd157} : s = 358;
	{8'd201,8'd158} : s = 359;
	{8'd201,8'd159} : s = 360;
	{8'd201,8'd160} : s = 361;
	{8'd201,8'd161} : s = 362;
	{8'd201,8'd162} : s = 363;
	{8'd201,8'd163} : s = 364;
	{8'd201,8'd164} : s = 365;
	{8'd201,8'd165} : s = 366;
	{8'd201,8'd166} : s = 367;
	{8'd201,8'd167} : s = 368;
	{8'd201,8'd168} : s = 369;
	{8'd201,8'd169} : s = 370;
	{8'd201,8'd170} : s = 371;
	{8'd201,8'd171} : s = 372;
	{8'd201,8'd172} : s = 373;
	{8'd201,8'd173} : s = 374;
	{8'd201,8'd174} : s = 375;
	{8'd201,8'd175} : s = 376;
	{8'd201,8'd176} : s = 377;
	{8'd201,8'd177} : s = 378;
	{8'd201,8'd178} : s = 379;
	{8'd201,8'd179} : s = 380;
	{8'd201,8'd180} : s = 381;
	{8'd201,8'd181} : s = 382;
	{8'd201,8'd182} : s = 383;
	{8'd201,8'd183} : s = 384;
	{8'd201,8'd184} : s = 385;
	{8'd201,8'd185} : s = 386;
	{8'd201,8'd186} : s = 387;
	{8'd201,8'd187} : s = 388;
	{8'd201,8'd188} : s = 389;
	{8'd201,8'd189} : s = 390;
	{8'd201,8'd190} : s = 391;
	{8'd201,8'd191} : s = 392;
	{8'd201,8'd192} : s = 393;
	{8'd201,8'd193} : s = 394;
	{8'd201,8'd194} : s = 395;
	{8'd201,8'd195} : s = 396;
	{8'd201,8'd196} : s = 397;
	{8'd201,8'd197} : s = 398;
	{8'd201,8'd198} : s = 399;
	{8'd201,8'd199} : s = 400;
	{8'd201,8'd200} : s = 401;
	{8'd201,8'd201} : s = 402;
	{8'd201,8'd202} : s = 403;
	{8'd201,8'd203} : s = 404;
	{8'd201,8'd204} : s = 405;
	{8'd201,8'd205} : s = 406;
	{8'd201,8'd206} : s = 407;
	{8'd201,8'd207} : s = 408;
	{8'd201,8'd208} : s = 409;
	{8'd201,8'd209} : s = 410;
	{8'd201,8'd210} : s = 411;
	{8'd201,8'd211} : s = 412;
	{8'd201,8'd212} : s = 413;
	{8'd201,8'd213} : s = 414;
	{8'd201,8'd214} : s = 415;
	{8'd201,8'd215} : s = 416;
	{8'd201,8'd216} : s = 417;
	{8'd201,8'd217} : s = 418;
	{8'd201,8'd218} : s = 419;
	{8'd201,8'd219} : s = 420;
	{8'd201,8'd220} : s = 421;
	{8'd201,8'd221} : s = 422;
	{8'd201,8'd222} : s = 423;
	{8'd201,8'd223} : s = 424;
	{8'd201,8'd224} : s = 425;
	{8'd201,8'd225} : s = 426;
	{8'd201,8'd226} : s = 427;
	{8'd201,8'd227} : s = 428;
	{8'd201,8'd228} : s = 429;
	{8'd201,8'd229} : s = 430;
	{8'd201,8'd230} : s = 431;
	{8'd201,8'd231} : s = 432;
	{8'd201,8'd232} : s = 433;
	{8'd201,8'd233} : s = 434;
	{8'd201,8'd234} : s = 435;
	{8'd201,8'd235} : s = 436;
	{8'd201,8'd236} : s = 437;
	{8'd201,8'd237} : s = 438;
	{8'd201,8'd238} : s = 439;
	{8'd201,8'd239} : s = 440;
	{8'd201,8'd240} : s = 441;
	{8'd201,8'd241} : s = 442;
	{8'd201,8'd242} : s = 443;
	{8'd201,8'd243} : s = 444;
	{8'd201,8'd244} : s = 445;
	{8'd201,8'd245} : s = 446;
	{8'd201,8'd246} : s = 447;
	{8'd201,8'd247} : s = 448;
	{8'd201,8'd248} : s = 449;
	{8'd201,8'd249} : s = 450;
	{8'd201,8'd250} : s = 451;
	{8'd201,8'd251} : s = 452;
	{8'd201,8'd252} : s = 453;
	{8'd201,8'd253} : s = 454;
	{8'd201,8'd254} : s = 455;
	{8'd201,8'd255} : s = 456;
	{8'd202,8'd0} : s = 202;
	{8'd202,8'd1} : s = 203;
	{8'd202,8'd2} : s = 204;
	{8'd202,8'd3} : s = 205;
	{8'd202,8'd4} : s = 206;
	{8'd202,8'd5} : s = 207;
	{8'd202,8'd6} : s = 208;
	{8'd202,8'd7} : s = 209;
	{8'd202,8'd8} : s = 210;
	{8'd202,8'd9} : s = 211;
	{8'd202,8'd10} : s = 212;
	{8'd202,8'd11} : s = 213;
	{8'd202,8'd12} : s = 214;
	{8'd202,8'd13} : s = 215;
	{8'd202,8'd14} : s = 216;
	{8'd202,8'd15} : s = 217;
	{8'd202,8'd16} : s = 218;
	{8'd202,8'd17} : s = 219;
	{8'd202,8'd18} : s = 220;
	{8'd202,8'd19} : s = 221;
	{8'd202,8'd20} : s = 222;
	{8'd202,8'd21} : s = 223;
	{8'd202,8'd22} : s = 224;
	{8'd202,8'd23} : s = 225;
	{8'd202,8'd24} : s = 226;
	{8'd202,8'd25} : s = 227;
	{8'd202,8'd26} : s = 228;
	{8'd202,8'd27} : s = 229;
	{8'd202,8'd28} : s = 230;
	{8'd202,8'd29} : s = 231;
	{8'd202,8'd30} : s = 232;
	{8'd202,8'd31} : s = 233;
	{8'd202,8'd32} : s = 234;
	{8'd202,8'd33} : s = 235;
	{8'd202,8'd34} : s = 236;
	{8'd202,8'd35} : s = 237;
	{8'd202,8'd36} : s = 238;
	{8'd202,8'd37} : s = 239;
	{8'd202,8'd38} : s = 240;
	{8'd202,8'd39} : s = 241;
	{8'd202,8'd40} : s = 242;
	{8'd202,8'd41} : s = 243;
	{8'd202,8'd42} : s = 244;
	{8'd202,8'd43} : s = 245;
	{8'd202,8'd44} : s = 246;
	{8'd202,8'd45} : s = 247;
	{8'd202,8'd46} : s = 248;
	{8'd202,8'd47} : s = 249;
	{8'd202,8'd48} : s = 250;
	{8'd202,8'd49} : s = 251;
	{8'd202,8'd50} : s = 252;
	{8'd202,8'd51} : s = 253;
	{8'd202,8'd52} : s = 254;
	{8'd202,8'd53} : s = 255;
	{8'd202,8'd54} : s = 256;
	{8'd202,8'd55} : s = 257;
	{8'd202,8'd56} : s = 258;
	{8'd202,8'd57} : s = 259;
	{8'd202,8'd58} : s = 260;
	{8'd202,8'd59} : s = 261;
	{8'd202,8'd60} : s = 262;
	{8'd202,8'd61} : s = 263;
	{8'd202,8'd62} : s = 264;
	{8'd202,8'd63} : s = 265;
	{8'd202,8'd64} : s = 266;
	{8'd202,8'd65} : s = 267;
	{8'd202,8'd66} : s = 268;
	{8'd202,8'd67} : s = 269;
	{8'd202,8'd68} : s = 270;
	{8'd202,8'd69} : s = 271;
	{8'd202,8'd70} : s = 272;
	{8'd202,8'd71} : s = 273;
	{8'd202,8'd72} : s = 274;
	{8'd202,8'd73} : s = 275;
	{8'd202,8'd74} : s = 276;
	{8'd202,8'd75} : s = 277;
	{8'd202,8'd76} : s = 278;
	{8'd202,8'd77} : s = 279;
	{8'd202,8'd78} : s = 280;
	{8'd202,8'd79} : s = 281;
	{8'd202,8'd80} : s = 282;
	{8'd202,8'd81} : s = 283;
	{8'd202,8'd82} : s = 284;
	{8'd202,8'd83} : s = 285;
	{8'd202,8'd84} : s = 286;
	{8'd202,8'd85} : s = 287;
	{8'd202,8'd86} : s = 288;
	{8'd202,8'd87} : s = 289;
	{8'd202,8'd88} : s = 290;
	{8'd202,8'd89} : s = 291;
	{8'd202,8'd90} : s = 292;
	{8'd202,8'd91} : s = 293;
	{8'd202,8'd92} : s = 294;
	{8'd202,8'd93} : s = 295;
	{8'd202,8'd94} : s = 296;
	{8'd202,8'd95} : s = 297;
	{8'd202,8'd96} : s = 298;
	{8'd202,8'd97} : s = 299;
	{8'd202,8'd98} : s = 300;
	{8'd202,8'd99} : s = 301;
	{8'd202,8'd100} : s = 302;
	{8'd202,8'd101} : s = 303;
	{8'd202,8'd102} : s = 304;
	{8'd202,8'd103} : s = 305;
	{8'd202,8'd104} : s = 306;
	{8'd202,8'd105} : s = 307;
	{8'd202,8'd106} : s = 308;
	{8'd202,8'd107} : s = 309;
	{8'd202,8'd108} : s = 310;
	{8'd202,8'd109} : s = 311;
	{8'd202,8'd110} : s = 312;
	{8'd202,8'd111} : s = 313;
	{8'd202,8'd112} : s = 314;
	{8'd202,8'd113} : s = 315;
	{8'd202,8'd114} : s = 316;
	{8'd202,8'd115} : s = 317;
	{8'd202,8'd116} : s = 318;
	{8'd202,8'd117} : s = 319;
	{8'd202,8'd118} : s = 320;
	{8'd202,8'd119} : s = 321;
	{8'd202,8'd120} : s = 322;
	{8'd202,8'd121} : s = 323;
	{8'd202,8'd122} : s = 324;
	{8'd202,8'd123} : s = 325;
	{8'd202,8'd124} : s = 326;
	{8'd202,8'd125} : s = 327;
	{8'd202,8'd126} : s = 328;
	{8'd202,8'd127} : s = 329;
	{8'd202,8'd128} : s = 330;
	{8'd202,8'd129} : s = 331;
	{8'd202,8'd130} : s = 332;
	{8'd202,8'd131} : s = 333;
	{8'd202,8'd132} : s = 334;
	{8'd202,8'd133} : s = 335;
	{8'd202,8'd134} : s = 336;
	{8'd202,8'd135} : s = 337;
	{8'd202,8'd136} : s = 338;
	{8'd202,8'd137} : s = 339;
	{8'd202,8'd138} : s = 340;
	{8'd202,8'd139} : s = 341;
	{8'd202,8'd140} : s = 342;
	{8'd202,8'd141} : s = 343;
	{8'd202,8'd142} : s = 344;
	{8'd202,8'd143} : s = 345;
	{8'd202,8'd144} : s = 346;
	{8'd202,8'd145} : s = 347;
	{8'd202,8'd146} : s = 348;
	{8'd202,8'd147} : s = 349;
	{8'd202,8'd148} : s = 350;
	{8'd202,8'd149} : s = 351;
	{8'd202,8'd150} : s = 352;
	{8'd202,8'd151} : s = 353;
	{8'd202,8'd152} : s = 354;
	{8'd202,8'd153} : s = 355;
	{8'd202,8'd154} : s = 356;
	{8'd202,8'd155} : s = 357;
	{8'd202,8'd156} : s = 358;
	{8'd202,8'd157} : s = 359;
	{8'd202,8'd158} : s = 360;
	{8'd202,8'd159} : s = 361;
	{8'd202,8'd160} : s = 362;
	{8'd202,8'd161} : s = 363;
	{8'd202,8'd162} : s = 364;
	{8'd202,8'd163} : s = 365;
	{8'd202,8'd164} : s = 366;
	{8'd202,8'd165} : s = 367;
	{8'd202,8'd166} : s = 368;
	{8'd202,8'd167} : s = 369;
	{8'd202,8'd168} : s = 370;
	{8'd202,8'd169} : s = 371;
	{8'd202,8'd170} : s = 372;
	{8'd202,8'd171} : s = 373;
	{8'd202,8'd172} : s = 374;
	{8'd202,8'd173} : s = 375;
	{8'd202,8'd174} : s = 376;
	{8'd202,8'd175} : s = 377;
	{8'd202,8'd176} : s = 378;
	{8'd202,8'd177} : s = 379;
	{8'd202,8'd178} : s = 380;
	{8'd202,8'd179} : s = 381;
	{8'd202,8'd180} : s = 382;
	{8'd202,8'd181} : s = 383;
	{8'd202,8'd182} : s = 384;
	{8'd202,8'd183} : s = 385;
	{8'd202,8'd184} : s = 386;
	{8'd202,8'd185} : s = 387;
	{8'd202,8'd186} : s = 388;
	{8'd202,8'd187} : s = 389;
	{8'd202,8'd188} : s = 390;
	{8'd202,8'd189} : s = 391;
	{8'd202,8'd190} : s = 392;
	{8'd202,8'd191} : s = 393;
	{8'd202,8'd192} : s = 394;
	{8'd202,8'd193} : s = 395;
	{8'd202,8'd194} : s = 396;
	{8'd202,8'd195} : s = 397;
	{8'd202,8'd196} : s = 398;
	{8'd202,8'd197} : s = 399;
	{8'd202,8'd198} : s = 400;
	{8'd202,8'd199} : s = 401;
	{8'd202,8'd200} : s = 402;
	{8'd202,8'd201} : s = 403;
	{8'd202,8'd202} : s = 404;
	{8'd202,8'd203} : s = 405;
	{8'd202,8'd204} : s = 406;
	{8'd202,8'd205} : s = 407;
	{8'd202,8'd206} : s = 408;
	{8'd202,8'd207} : s = 409;
	{8'd202,8'd208} : s = 410;
	{8'd202,8'd209} : s = 411;
	{8'd202,8'd210} : s = 412;
	{8'd202,8'd211} : s = 413;
	{8'd202,8'd212} : s = 414;
	{8'd202,8'd213} : s = 415;
	{8'd202,8'd214} : s = 416;
	{8'd202,8'd215} : s = 417;
	{8'd202,8'd216} : s = 418;
	{8'd202,8'd217} : s = 419;
	{8'd202,8'd218} : s = 420;
	{8'd202,8'd219} : s = 421;
	{8'd202,8'd220} : s = 422;
	{8'd202,8'd221} : s = 423;
	{8'd202,8'd222} : s = 424;
	{8'd202,8'd223} : s = 425;
	{8'd202,8'd224} : s = 426;
	{8'd202,8'd225} : s = 427;
	{8'd202,8'd226} : s = 428;
	{8'd202,8'd227} : s = 429;
	{8'd202,8'd228} : s = 430;
	{8'd202,8'd229} : s = 431;
	{8'd202,8'd230} : s = 432;
	{8'd202,8'd231} : s = 433;
	{8'd202,8'd232} : s = 434;
	{8'd202,8'd233} : s = 435;
	{8'd202,8'd234} : s = 436;
	{8'd202,8'd235} : s = 437;
	{8'd202,8'd236} : s = 438;
	{8'd202,8'd237} : s = 439;
	{8'd202,8'd238} : s = 440;
	{8'd202,8'd239} : s = 441;
	{8'd202,8'd240} : s = 442;
	{8'd202,8'd241} : s = 443;
	{8'd202,8'd242} : s = 444;
	{8'd202,8'd243} : s = 445;
	{8'd202,8'd244} : s = 446;
	{8'd202,8'd245} : s = 447;
	{8'd202,8'd246} : s = 448;
	{8'd202,8'd247} : s = 449;
	{8'd202,8'd248} : s = 450;
	{8'd202,8'd249} : s = 451;
	{8'd202,8'd250} : s = 452;
	{8'd202,8'd251} : s = 453;
	{8'd202,8'd252} : s = 454;
	{8'd202,8'd253} : s = 455;
	{8'd202,8'd254} : s = 456;
	{8'd202,8'd255} : s = 457;
	{8'd203,8'd0} : s = 203;
	{8'd203,8'd1} : s = 204;
	{8'd203,8'd2} : s = 205;
	{8'd203,8'd3} : s = 206;
	{8'd203,8'd4} : s = 207;
	{8'd203,8'd5} : s = 208;
	{8'd203,8'd6} : s = 209;
	{8'd203,8'd7} : s = 210;
	{8'd203,8'd8} : s = 211;
	{8'd203,8'd9} : s = 212;
	{8'd203,8'd10} : s = 213;
	{8'd203,8'd11} : s = 214;
	{8'd203,8'd12} : s = 215;
	{8'd203,8'd13} : s = 216;
	{8'd203,8'd14} : s = 217;
	{8'd203,8'd15} : s = 218;
	{8'd203,8'd16} : s = 219;
	{8'd203,8'd17} : s = 220;
	{8'd203,8'd18} : s = 221;
	{8'd203,8'd19} : s = 222;
	{8'd203,8'd20} : s = 223;
	{8'd203,8'd21} : s = 224;
	{8'd203,8'd22} : s = 225;
	{8'd203,8'd23} : s = 226;
	{8'd203,8'd24} : s = 227;
	{8'd203,8'd25} : s = 228;
	{8'd203,8'd26} : s = 229;
	{8'd203,8'd27} : s = 230;
	{8'd203,8'd28} : s = 231;
	{8'd203,8'd29} : s = 232;
	{8'd203,8'd30} : s = 233;
	{8'd203,8'd31} : s = 234;
	{8'd203,8'd32} : s = 235;
	{8'd203,8'd33} : s = 236;
	{8'd203,8'd34} : s = 237;
	{8'd203,8'd35} : s = 238;
	{8'd203,8'd36} : s = 239;
	{8'd203,8'd37} : s = 240;
	{8'd203,8'd38} : s = 241;
	{8'd203,8'd39} : s = 242;
	{8'd203,8'd40} : s = 243;
	{8'd203,8'd41} : s = 244;
	{8'd203,8'd42} : s = 245;
	{8'd203,8'd43} : s = 246;
	{8'd203,8'd44} : s = 247;
	{8'd203,8'd45} : s = 248;
	{8'd203,8'd46} : s = 249;
	{8'd203,8'd47} : s = 250;
	{8'd203,8'd48} : s = 251;
	{8'd203,8'd49} : s = 252;
	{8'd203,8'd50} : s = 253;
	{8'd203,8'd51} : s = 254;
	{8'd203,8'd52} : s = 255;
	{8'd203,8'd53} : s = 256;
	{8'd203,8'd54} : s = 257;
	{8'd203,8'd55} : s = 258;
	{8'd203,8'd56} : s = 259;
	{8'd203,8'd57} : s = 260;
	{8'd203,8'd58} : s = 261;
	{8'd203,8'd59} : s = 262;
	{8'd203,8'd60} : s = 263;
	{8'd203,8'd61} : s = 264;
	{8'd203,8'd62} : s = 265;
	{8'd203,8'd63} : s = 266;
	{8'd203,8'd64} : s = 267;
	{8'd203,8'd65} : s = 268;
	{8'd203,8'd66} : s = 269;
	{8'd203,8'd67} : s = 270;
	{8'd203,8'd68} : s = 271;
	{8'd203,8'd69} : s = 272;
	{8'd203,8'd70} : s = 273;
	{8'd203,8'd71} : s = 274;
	{8'd203,8'd72} : s = 275;
	{8'd203,8'd73} : s = 276;
	{8'd203,8'd74} : s = 277;
	{8'd203,8'd75} : s = 278;
	{8'd203,8'd76} : s = 279;
	{8'd203,8'd77} : s = 280;
	{8'd203,8'd78} : s = 281;
	{8'd203,8'd79} : s = 282;
	{8'd203,8'd80} : s = 283;
	{8'd203,8'd81} : s = 284;
	{8'd203,8'd82} : s = 285;
	{8'd203,8'd83} : s = 286;
	{8'd203,8'd84} : s = 287;
	{8'd203,8'd85} : s = 288;
	{8'd203,8'd86} : s = 289;
	{8'd203,8'd87} : s = 290;
	{8'd203,8'd88} : s = 291;
	{8'd203,8'd89} : s = 292;
	{8'd203,8'd90} : s = 293;
	{8'd203,8'd91} : s = 294;
	{8'd203,8'd92} : s = 295;
	{8'd203,8'd93} : s = 296;
	{8'd203,8'd94} : s = 297;
	{8'd203,8'd95} : s = 298;
	{8'd203,8'd96} : s = 299;
	{8'd203,8'd97} : s = 300;
	{8'd203,8'd98} : s = 301;
	{8'd203,8'd99} : s = 302;
	{8'd203,8'd100} : s = 303;
	{8'd203,8'd101} : s = 304;
	{8'd203,8'd102} : s = 305;
	{8'd203,8'd103} : s = 306;
	{8'd203,8'd104} : s = 307;
	{8'd203,8'd105} : s = 308;
	{8'd203,8'd106} : s = 309;
	{8'd203,8'd107} : s = 310;
	{8'd203,8'd108} : s = 311;
	{8'd203,8'd109} : s = 312;
	{8'd203,8'd110} : s = 313;
	{8'd203,8'd111} : s = 314;
	{8'd203,8'd112} : s = 315;
	{8'd203,8'd113} : s = 316;
	{8'd203,8'd114} : s = 317;
	{8'd203,8'd115} : s = 318;
	{8'd203,8'd116} : s = 319;
	{8'd203,8'd117} : s = 320;
	{8'd203,8'd118} : s = 321;
	{8'd203,8'd119} : s = 322;
	{8'd203,8'd120} : s = 323;
	{8'd203,8'd121} : s = 324;
	{8'd203,8'd122} : s = 325;
	{8'd203,8'd123} : s = 326;
	{8'd203,8'd124} : s = 327;
	{8'd203,8'd125} : s = 328;
	{8'd203,8'd126} : s = 329;
	{8'd203,8'd127} : s = 330;
	{8'd203,8'd128} : s = 331;
	{8'd203,8'd129} : s = 332;
	{8'd203,8'd130} : s = 333;
	{8'd203,8'd131} : s = 334;
	{8'd203,8'd132} : s = 335;
	{8'd203,8'd133} : s = 336;
	{8'd203,8'd134} : s = 337;
	{8'd203,8'd135} : s = 338;
	{8'd203,8'd136} : s = 339;
	{8'd203,8'd137} : s = 340;
	{8'd203,8'd138} : s = 341;
	{8'd203,8'd139} : s = 342;
	{8'd203,8'd140} : s = 343;
	{8'd203,8'd141} : s = 344;
	{8'd203,8'd142} : s = 345;
	{8'd203,8'd143} : s = 346;
	{8'd203,8'd144} : s = 347;
	{8'd203,8'd145} : s = 348;
	{8'd203,8'd146} : s = 349;
	{8'd203,8'd147} : s = 350;
	{8'd203,8'd148} : s = 351;
	{8'd203,8'd149} : s = 352;
	{8'd203,8'd150} : s = 353;
	{8'd203,8'd151} : s = 354;
	{8'd203,8'd152} : s = 355;
	{8'd203,8'd153} : s = 356;
	{8'd203,8'd154} : s = 357;
	{8'd203,8'd155} : s = 358;
	{8'd203,8'd156} : s = 359;
	{8'd203,8'd157} : s = 360;
	{8'd203,8'd158} : s = 361;
	{8'd203,8'd159} : s = 362;
	{8'd203,8'd160} : s = 363;
	{8'd203,8'd161} : s = 364;
	{8'd203,8'd162} : s = 365;
	{8'd203,8'd163} : s = 366;
	{8'd203,8'd164} : s = 367;
	{8'd203,8'd165} : s = 368;
	{8'd203,8'd166} : s = 369;
	{8'd203,8'd167} : s = 370;
	{8'd203,8'd168} : s = 371;
	{8'd203,8'd169} : s = 372;
	{8'd203,8'd170} : s = 373;
	{8'd203,8'd171} : s = 374;
	{8'd203,8'd172} : s = 375;
	{8'd203,8'd173} : s = 376;
	{8'd203,8'd174} : s = 377;
	{8'd203,8'd175} : s = 378;
	{8'd203,8'd176} : s = 379;
	{8'd203,8'd177} : s = 380;
	{8'd203,8'd178} : s = 381;
	{8'd203,8'd179} : s = 382;
	{8'd203,8'd180} : s = 383;
	{8'd203,8'd181} : s = 384;
	{8'd203,8'd182} : s = 385;
	{8'd203,8'd183} : s = 386;
	{8'd203,8'd184} : s = 387;
	{8'd203,8'd185} : s = 388;
	{8'd203,8'd186} : s = 389;
	{8'd203,8'd187} : s = 390;
	{8'd203,8'd188} : s = 391;
	{8'd203,8'd189} : s = 392;
	{8'd203,8'd190} : s = 393;
	{8'd203,8'd191} : s = 394;
	{8'd203,8'd192} : s = 395;
	{8'd203,8'd193} : s = 396;
	{8'd203,8'd194} : s = 397;
	{8'd203,8'd195} : s = 398;
	{8'd203,8'd196} : s = 399;
	{8'd203,8'd197} : s = 400;
	{8'd203,8'd198} : s = 401;
	{8'd203,8'd199} : s = 402;
	{8'd203,8'd200} : s = 403;
	{8'd203,8'd201} : s = 404;
	{8'd203,8'd202} : s = 405;
	{8'd203,8'd203} : s = 406;
	{8'd203,8'd204} : s = 407;
	{8'd203,8'd205} : s = 408;
	{8'd203,8'd206} : s = 409;
	{8'd203,8'd207} : s = 410;
	{8'd203,8'd208} : s = 411;
	{8'd203,8'd209} : s = 412;
	{8'd203,8'd210} : s = 413;
	{8'd203,8'd211} : s = 414;
	{8'd203,8'd212} : s = 415;
	{8'd203,8'd213} : s = 416;
	{8'd203,8'd214} : s = 417;
	{8'd203,8'd215} : s = 418;
	{8'd203,8'd216} : s = 419;
	{8'd203,8'd217} : s = 420;
	{8'd203,8'd218} : s = 421;
	{8'd203,8'd219} : s = 422;
	{8'd203,8'd220} : s = 423;
	{8'd203,8'd221} : s = 424;
	{8'd203,8'd222} : s = 425;
	{8'd203,8'd223} : s = 426;
	{8'd203,8'd224} : s = 427;
	{8'd203,8'd225} : s = 428;
	{8'd203,8'd226} : s = 429;
	{8'd203,8'd227} : s = 430;
	{8'd203,8'd228} : s = 431;
	{8'd203,8'd229} : s = 432;
	{8'd203,8'd230} : s = 433;
	{8'd203,8'd231} : s = 434;
	{8'd203,8'd232} : s = 435;
	{8'd203,8'd233} : s = 436;
	{8'd203,8'd234} : s = 437;
	{8'd203,8'd235} : s = 438;
	{8'd203,8'd236} : s = 439;
	{8'd203,8'd237} : s = 440;
	{8'd203,8'd238} : s = 441;
	{8'd203,8'd239} : s = 442;
	{8'd203,8'd240} : s = 443;
	{8'd203,8'd241} : s = 444;
	{8'd203,8'd242} : s = 445;
	{8'd203,8'd243} : s = 446;
	{8'd203,8'd244} : s = 447;
	{8'd203,8'd245} : s = 448;
	{8'd203,8'd246} : s = 449;
	{8'd203,8'd247} : s = 450;
	{8'd203,8'd248} : s = 451;
	{8'd203,8'd249} : s = 452;
	{8'd203,8'd250} : s = 453;
	{8'd203,8'd251} : s = 454;
	{8'd203,8'd252} : s = 455;
	{8'd203,8'd253} : s = 456;
	{8'd203,8'd254} : s = 457;
	{8'd203,8'd255} : s = 458;
	{8'd204,8'd0} : s = 204;
	{8'd204,8'd1} : s = 205;
	{8'd204,8'd2} : s = 206;
	{8'd204,8'd3} : s = 207;
	{8'd204,8'd4} : s = 208;
	{8'd204,8'd5} : s = 209;
	{8'd204,8'd6} : s = 210;
	{8'd204,8'd7} : s = 211;
	{8'd204,8'd8} : s = 212;
	{8'd204,8'd9} : s = 213;
	{8'd204,8'd10} : s = 214;
	{8'd204,8'd11} : s = 215;
	{8'd204,8'd12} : s = 216;
	{8'd204,8'd13} : s = 217;
	{8'd204,8'd14} : s = 218;
	{8'd204,8'd15} : s = 219;
	{8'd204,8'd16} : s = 220;
	{8'd204,8'd17} : s = 221;
	{8'd204,8'd18} : s = 222;
	{8'd204,8'd19} : s = 223;
	{8'd204,8'd20} : s = 224;
	{8'd204,8'd21} : s = 225;
	{8'd204,8'd22} : s = 226;
	{8'd204,8'd23} : s = 227;
	{8'd204,8'd24} : s = 228;
	{8'd204,8'd25} : s = 229;
	{8'd204,8'd26} : s = 230;
	{8'd204,8'd27} : s = 231;
	{8'd204,8'd28} : s = 232;
	{8'd204,8'd29} : s = 233;
	{8'd204,8'd30} : s = 234;
	{8'd204,8'd31} : s = 235;
	{8'd204,8'd32} : s = 236;
	{8'd204,8'd33} : s = 237;
	{8'd204,8'd34} : s = 238;
	{8'd204,8'd35} : s = 239;
	{8'd204,8'd36} : s = 240;
	{8'd204,8'd37} : s = 241;
	{8'd204,8'd38} : s = 242;
	{8'd204,8'd39} : s = 243;
	{8'd204,8'd40} : s = 244;
	{8'd204,8'd41} : s = 245;
	{8'd204,8'd42} : s = 246;
	{8'd204,8'd43} : s = 247;
	{8'd204,8'd44} : s = 248;
	{8'd204,8'd45} : s = 249;
	{8'd204,8'd46} : s = 250;
	{8'd204,8'd47} : s = 251;
	{8'd204,8'd48} : s = 252;
	{8'd204,8'd49} : s = 253;
	{8'd204,8'd50} : s = 254;
	{8'd204,8'd51} : s = 255;
	{8'd204,8'd52} : s = 256;
	{8'd204,8'd53} : s = 257;
	{8'd204,8'd54} : s = 258;
	{8'd204,8'd55} : s = 259;
	{8'd204,8'd56} : s = 260;
	{8'd204,8'd57} : s = 261;
	{8'd204,8'd58} : s = 262;
	{8'd204,8'd59} : s = 263;
	{8'd204,8'd60} : s = 264;
	{8'd204,8'd61} : s = 265;
	{8'd204,8'd62} : s = 266;
	{8'd204,8'd63} : s = 267;
	{8'd204,8'd64} : s = 268;
	{8'd204,8'd65} : s = 269;
	{8'd204,8'd66} : s = 270;
	{8'd204,8'd67} : s = 271;
	{8'd204,8'd68} : s = 272;
	{8'd204,8'd69} : s = 273;
	{8'd204,8'd70} : s = 274;
	{8'd204,8'd71} : s = 275;
	{8'd204,8'd72} : s = 276;
	{8'd204,8'd73} : s = 277;
	{8'd204,8'd74} : s = 278;
	{8'd204,8'd75} : s = 279;
	{8'd204,8'd76} : s = 280;
	{8'd204,8'd77} : s = 281;
	{8'd204,8'd78} : s = 282;
	{8'd204,8'd79} : s = 283;
	{8'd204,8'd80} : s = 284;
	{8'd204,8'd81} : s = 285;
	{8'd204,8'd82} : s = 286;
	{8'd204,8'd83} : s = 287;
	{8'd204,8'd84} : s = 288;
	{8'd204,8'd85} : s = 289;
	{8'd204,8'd86} : s = 290;
	{8'd204,8'd87} : s = 291;
	{8'd204,8'd88} : s = 292;
	{8'd204,8'd89} : s = 293;
	{8'd204,8'd90} : s = 294;
	{8'd204,8'd91} : s = 295;
	{8'd204,8'd92} : s = 296;
	{8'd204,8'd93} : s = 297;
	{8'd204,8'd94} : s = 298;
	{8'd204,8'd95} : s = 299;
	{8'd204,8'd96} : s = 300;
	{8'd204,8'd97} : s = 301;
	{8'd204,8'd98} : s = 302;
	{8'd204,8'd99} : s = 303;
	{8'd204,8'd100} : s = 304;
	{8'd204,8'd101} : s = 305;
	{8'd204,8'd102} : s = 306;
	{8'd204,8'd103} : s = 307;
	{8'd204,8'd104} : s = 308;
	{8'd204,8'd105} : s = 309;
	{8'd204,8'd106} : s = 310;
	{8'd204,8'd107} : s = 311;
	{8'd204,8'd108} : s = 312;
	{8'd204,8'd109} : s = 313;
	{8'd204,8'd110} : s = 314;
	{8'd204,8'd111} : s = 315;
	{8'd204,8'd112} : s = 316;
	{8'd204,8'd113} : s = 317;
	{8'd204,8'd114} : s = 318;
	{8'd204,8'd115} : s = 319;
	{8'd204,8'd116} : s = 320;
	{8'd204,8'd117} : s = 321;
	{8'd204,8'd118} : s = 322;
	{8'd204,8'd119} : s = 323;
	{8'd204,8'd120} : s = 324;
	{8'd204,8'd121} : s = 325;
	{8'd204,8'd122} : s = 326;
	{8'd204,8'd123} : s = 327;
	{8'd204,8'd124} : s = 328;
	{8'd204,8'd125} : s = 329;
	{8'd204,8'd126} : s = 330;
	{8'd204,8'd127} : s = 331;
	{8'd204,8'd128} : s = 332;
	{8'd204,8'd129} : s = 333;
	{8'd204,8'd130} : s = 334;
	{8'd204,8'd131} : s = 335;
	{8'd204,8'd132} : s = 336;
	{8'd204,8'd133} : s = 337;
	{8'd204,8'd134} : s = 338;
	{8'd204,8'd135} : s = 339;
	{8'd204,8'd136} : s = 340;
	{8'd204,8'd137} : s = 341;
	{8'd204,8'd138} : s = 342;
	{8'd204,8'd139} : s = 343;
	{8'd204,8'd140} : s = 344;
	{8'd204,8'd141} : s = 345;
	{8'd204,8'd142} : s = 346;
	{8'd204,8'd143} : s = 347;
	{8'd204,8'd144} : s = 348;
	{8'd204,8'd145} : s = 349;
	{8'd204,8'd146} : s = 350;
	{8'd204,8'd147} : s = 351;
	{8'd204,8'd148} : s = 352;
	{8'd204,8'd149} : s = 353;
	{8'd204,8'd150} : s = 354;
	{8'd204,8'd151} : s = 355;
	{8'd204,8'd152} : s = 356;
	{8'd204,8'd153} : s = 357;
	{8'd204,8'd154} : s = 358;
	{8'd204,8'd155} : s = 359;
	{8'd204,8'd156} : s = 360;
	{8'd204,8'd157} : s = 361;
	{8'd204,8'd158} : s = 362;
	{8'd204,8'd159} : s = 363;
	{8'd204,8'd160} : s = 364;
	{8'd204,8'd161} : s = 365;
	{8'd204,8'd162} : s = 366;
	{8'd204,8'd163} : s = 367;
	{8'd204,8'd164} : s = 368;
	{8'd204,8'd165} : s = 369;
	{8'd204,8'd166} : s = 370;
	{8'd204,8'd167} : s = 371;
	{8'd204,8'd168} : s = 372;
	{8'd204,8'd169} : s = 373;
	{8'd204,8'd170} : s = 374;
	{8'd204,8'd171} : s = 375;
	{8'd204,8'd172} : s = 376;
	{8'd204,8'd173} : s = 377;
	{8'd204,8'd174} : s = 378;
	{8'd204,8'd175} : s = 379;
	{8'd204,8'd176} : s = 380;
	{8'd204,8'd177} : s = 381;
	{8'd204,8'd178} : s = 382;
	{8'd204,8'd179} : s = 383;
	{8'd204,8'd180} : s = 384;
	{8'd204,8'd181} : s = 385;
	{8'd204,8'd182} : s = 386;
	{8'd204,8'd183} : s = 387;
	{8'd204,8'd184} : s = 388;
	{8'd204,8'd185} : s = 389;
	{8'd204,8'd186} : s = 390;
	{8'd204,8'd187} : s = 391;
	{8'd204,8'd188} : s = 392;
	{8'd204,8'd189} : s = 393;
	{8'd204,8'd190} : s = 394;
	{8'd204,8'd191} : s = 395;
	{8'd204,8'd192} : s = 396;
	{8'd204,8'd193} : s = 397;
	{8'd204,8'd194} : s = 398;
	{8'd204,8'd195} : s = 399;
	{8'd204,8'd196} : s = 400;
	{8'd204,8'd197} : s = 401;
	{8'd204,8'd198} : s = 402;
	{8'd204,8'd199} : s = 403;
	{8'd204,8'd200} : s = 404;
	{8'd204,8'd201} : s = 405;
	{8'd204,8'd202} : s = 406;
	{8'd204,8'd203} : s = 407;
	{8'd204,8'd204} : s = 408;
	{8'd204,8'd205} : s = 409;
	{8'd204,8'd206} : s = 410;
	{8'd204,8'd207} : s = 411;
	{8'd204,8'd208} : s = 412;
	{8'd204,8'd209} : s = 413;
	{8'd204,8'd210} : s = 414;
	{8'd204,8'd211} : s = 415;
	{8'd204,8'd212} : s = 416;
	{8'd204,8'd213} : s = 417;
	{8'd204,8'd214} : s = 418;
	{8'd204,8'd215} : s = 419;
	{8'd204,8'd216} : s = 420;
	{8'd204,8'd217} : s = 421;
	{8'd204,8'd218} : s = 422;
	{8'd204,8'd219} : s = 423;
	{8'd204,8'd220} : s = 424;
	{8'd204,8'd221} : s = 425;
	{8'd204,8'd222} : s = 426;
	{8'd204,8'd223} : s = 427;
	{8'd204,8'd224} : s = 428;
	{8'd204,8'd225} : s = 429;
	{8'd204,8'd226} : s = 430;
	{8'd204,8'd227} : s = 431;
	{8'd204,8'd228} : s = 432;
	{8'd204,8'd229} : s = 433;
	{8'd204,8'd230} : s = 434;
	{8'd204,8'd231} : s = 435;
	{8'd204,8'd232} : s = 436;
	{8'd204,8'd233} : s = 437;
	{8'd204,8'd234} : s = 438;
	{8'd204,8'd235} : s = 439;
	{8'd204,8'd236} : s = 440;
	{8'd204,8'd237} : s = 441;
	{8'd204,8'd238} : s = 442;
	{8'd204,8'd239} : s = 443;
	{8'd204,8'd240} : s = 444;
	{8'd204,8'd241} : s = 445;
	{8'd204,8'd242} : s = 446;
	{8'd204,8'd243} : s = 447;
	{8'd204,8'd244} : s = 448;
	{8'd204,8'd245} : s = 449;
	{8'd204,8'd246} : s = 450;
	{8'd204,8'd247} : s = 451;
	{8'd204,8'd248} : s = 452;
	{8'd204,8'd249} : s = 453;
	{8'd204,8'd250} : s = 454;
	{8'd204,8'd251} : s = 455;
	{8'd204,8'd252} : s = 456;
	{8'd204,8'd253} : s = 457;
	{8'd204,8'd254} : s = 458;
	{8'd204,8'd255} : s = 459;
	{8'd205,8'd0} : s = 205;
	{8'd205,8'd1} : s = 206;
	{8'd205,8'd2} : s = 207;
	{8'd205,8'd3} : s = 208;
	{8'd205,8'd4} : s = 209;
	{8'd205,8'd5} : s = 210;
	{8'd205,8'd6} : s = 211;
	{8'd205,8'd7} : s = 212;
	{8'd205,8'd8} : s = 213;
	{8'd205,8'd9} : s = 214;
	{8'd205,8'd10} : s = 215;
	{8'd205,8'd11} : s = 216;
	{8'd205,8'd12} : s = 217;
	{8'd205,8'd13} : s = 218;
	{8'd205,8'd14} : s = 219;
	{8'd205,8'd15} : s = 220;
	{8'd205,8'd16} : s = 221;
	{8'd205,8'd17} : s = 222;
	{8'd205,8'd18} : s = 223;
	{8'd205,8'd19} : s = 224;
	{8'd205,8'd20} : s = 225;
	{8'd205,8'd21} : s = 226;
	{8'd205,8'd22} : s = 227;
	{8'd205,8'd23} : s = 228;
	{8'd205,8'd24} : s = 229;
	{8'd205,8'd25} : s = 230;
	{8'd205,8'd26} : s = 231;
	{8'd205,8'd27} : s = 232;
	{8'd205,8'd28} : s = 233;
	{8'd205,8'd29} : s = 234;
	{8'd205,8'd30} : s = 235;
	{8'd205,8'd31} : s = 236;
	{8'd205,8'd32} : s = 237;
	{8'd205,8'd33} : s = 238;
	{8'd205,8'd34} : s = 239;
	{8'd205,8'd35} : s = 240;
	{8'd205,8'd36} : s = 241;
	{8'd205,8'd37} : s = 242;
	{8'd205,8'd38} : s = 243;
	{8'd205,8'd39} : s = 244;
	{8'd205,8'd40} : s = 245;
	{8'd205,8'd41} : s = 246;
	{8'd205,8'd42} : s = 247;
	{8'd205,8'd43} : s = 248;
	{8'd205,8'd44} : s = 249;
	{8'd205,8'd45} : s = 250;
	{8'd205,8'd46} : s = 251;
	{8'd205,8'd47} : s = 252;
	{8'd205,8'd48} : s = 253;
	{8'd205,8'd49} : s = 254;
	{8'd205,8'd50} : s = 255;
	{8'd205,8'd51} : s = 256;
	{8'd205,8'd52} : s = 257;
	{8'd205,8'd53} : s = 258;
	{8'd205,8'd54} : s = 259;
	{8'd205,8'd55} : s = 260;
	{8'd205,8'd56} : s = 261;
	{8'd205,8'd57} : s = 262;
	{8'd205,8'd58} : s = 263;
	{8'd205,8'd59} : s = 264;
	{8'd205,8'd60} : s = 265;
	{8'd205,8'd61} : s = 266;
	{8'd205,8'd62} : s = 267;
	{8'd205,8'd63} : s = 268;
	{8'd205,8'd64} : s = 269;
	{8'd205,8'd65} : s = 270;
	{8'd205,8'd66} : s = 271;
	{8'd205,8'd67} : s = 272;
	{8'd205,8'd68} : s = 273;
	{8'd205,8'd69} : s = 274;
	{8'd205,8'd70} : s = 275;
	{8'd205,8'd71} : s = 276;
	{8'd205,8'd72} : s = 277;
	{8'd205,8'd73} : s = 278;
	{8'd205,8'd74} : s = 279;
	{8'd205,8'd75} : s = 280;
	{8'd205,8'd76} : s = 281;
	{8'd205,8'd77} : s = 282;
	{8'd205,8'd78} : s = 283;
	{8'd205,8'd79} : s = 284;
	{8'd205,8'd80} : s = 285;
	{8'd205,8'd81} : s = 286;
	{8'd205,8'd82} : s = 287;
	{8'd205,8'd83} : s = 288;
	{8'd205,8'd84} : s = 289;
	{8'd205,8'd85} : s = 290;
	{8'd205,8'd86} : s = 291;
	{8'd205,8'd87} : s = 292;
	{8'd205,8'd88} : s = 293;
	{8'd205,8'd89} : s = 294;
	{8'd205,8'd90} : s = 295;
	{8'd205,8'd91} : s = 296;
	{8'd205,8'd92} : s = 297;
	{8'd205,8'd93} : s = 298;
	{8'd205,8'd94} : s = 299;
	{8'd205,8'd95} : s = 300;
	{8'd205,8'd96} : s = 301;
	{8'd205,8'd97} : s = 302;
	{8'd205,8'd98} : s = 303;
	{8'd205,8'd99} : s = 304;
	{8'd205,8'd100} : s = 305;
	{8'd205,8'd101} : s = 306;
	{8'd205,8'd102} : s = 307;
	{8'd205,8'd103} : s = 308;
	{8'd205,8'd104} : s = 309;
	{8'd205,8'd105} : s = 310;
	{8'd205,8'd106} : s = 311;
	{8'd205,8'd107} : s = 312;
	{8'd205,8'd108} : s = 313;
	{8'd205,8'd109} : s = 314;
	{8'd205,8'd110} : s = 315;
	{8'd205,8'd111} : s = 316;
	{8'd205,8'd112} : s = 317;
	{8'd205,8'd113} : s = 318;
	{8'd205,8'd114} : s = 319;
	{8'd205,8'd115} : s = 320;
	{8'd205,8'd116} : s = 321;
	{8'd205,8'd117} : s = 322;
	{8'd205,8'd118} : s = 323;
	{8'd205,8'd119} : s = 324;
	{8'd205,8'd120} : s = 325;
	{8'd205,8'd121} : s = 326;
	{8'd205,8'd122} : s = 327;
	{8'd205,8'd123} : s = 328;
	{8'd205,8'd124} : s = 329;
	{8'd205,8'd125} : s = 330;
	{8'd205,8'd126} : s = 331;
	{8'd205,8'd127} : s = 332;
	{8'd205,8'd128} : s = 333;
	{8'd205,8'd129} : s = 334;
	{8'd205,8'd130} : s = 335;
	{8'd205,8'd131} : s = 336;
	{8'd205,8'd132} : s = 337;
	{8'd205,8'd133} : s = 338;
	{8'd205,8'd134} : s = 339;
	{8'd205,8'd135} : s = 340;
	{8'd205,8'd136} : s = 341;
	{8'd205,8'd137} : s = 342;
	{8'd205,8'd138} : s = 343;
	{8'd205,8'd139} : s = 344;
	{8'd205,8'd140} : s = 345;
	{8'd205,8'd141} : s = 346;
	{8'd205,8'd142} : s = 347;
	{8'd205,8'd143} : s = 348;
	{8'd205,8'd144} : s = 349;
	{8'd205,8'd145} : s = 350;
	{8'd205,8'd146} : s = 351;
	{8'd205,8'd147} : s = 352;
	{8'd205,8'd148} : s = 353;
	{8'd205,8'd149} : s = 354;
	{8'd205,8'd150} : s = 355;
	{8'd205,8'd151} : s = 356;
	{8'd205,8'd152} : s = 357;
	{8'd205,8'd153} : s = 358;
	{8'd205,8'd154} : s = 359;
	{8'd205,8'd155} : s = 360;
	{8'd205,8'd156} : s = 361;
	{8'd205,8'd157} : s = 362;
	{8'd205,8'd158} : s = 363;
	{8'd205,8'd159} : s = 364;
	{8'd205,8'd160} : s = 365;
	{8'd205,8'd161} : s = 366;
	{8'd205,8'd162} : s = 367;
	{8'd205,8'd163} : s = 368;
	{8'd205,8'd164} : s = 369;
	{8'd205,8'd165} : s = 370;
	{8'd205,8'd166} : s = 371;
	{8'd205,8'd167} : s = 372;
	{8'd205,8'd168} : s = 373;
	{8'd205,8'd169} : s = 374;
	{8'd205,8'd170} : s = 375;
	{8'd205,8'd171} : s = 376;
	{8'd205,8'd172} : s = 377;
	{8'd205,8'd173} : s = 378;
	{8'd205,8'd174} : s = 379;
	{8'd205,8'd175} : s = 380;
	{8'd205,8'd176} : s = 381;
	{8'd205,8'd177} : s = 382;
	{8'd205,8'd178} : s = 383;
	{8'd205,8'd179} : s = 384;
	{8'd205,8'd180} : s = 385;
	{8'd205,8'd181} : s = 386;
	{8'd205,8'd182} : s = 387;
	{8'd205,8'd183} : s = 388;
	{8'd205,8'd184} : s = 389;
	{8'd205,8'd185} : s = 390;
	{8'd205,8'd186} : s = 391;
	{8'd205,8'd187} : s = 392;
	{8'd205,8'd188} : s = 393;
	{8'd205,8'd189} : s = 394;
	{8'd205,8'd190} : s = 395;
	{8'd205,8'd191} : s = 396;
	{8'd205,8'd192} : s = 397;
	{8'd205,8'd193} : s = 398;
	{8'd205,8'd194} : s = 399;
	{8'd205,8'd195} : s = 400;
	{8'd205,8'd196} : s = 401;
	{8'd205,8'd197} : s = 402;
	{8'd205,8'd198} : s = 403;
	{8'd205,8'd199} : s = 404;
	{8'd205,8'd200} : s = 405;
	{8'd205,8'd201} : s = 406;
	{8'd205,8'd202} : s = 407;
	{8'd205,8'd203} : s = 408;
	{8'd205,8'd204} : s = 409;
	{8'd205,8'd205} : s = 410;
	{8'd205,8'd206} : s = 411;
	{8'd205,8'd207} : s = 412;
	{8'd205,8'd208} : s = 413;
	{8'd205,8'd209} : s = 414;
	{8'd205,8'd210} : s = 415;
	{8'd205,8'd211} : s = 416;
	{8'd205,8'd212} : s = 417;
	{8'd205,8'd213} : s = 418;
	{8'd205,8'd214} : s = 419;
	{8'd205,8'd215} : s = 420;
	{8'd205,8'd216} : s = 421;
	{8'd205,8'd217} : s = 422;
	{8'd205,8'd218} : s = 423;
	{8'd205,8'd219} : s = 424;
	{8'd205,8'd220} : s = 425;
	{8'd205,8'd221} : s = 426;
	{8'd205,8'd222} : s = 427;
	{8'd205,8'd223} : s = 428;
	{8'd205,8'd224} : s = 429;
	{8'd205,8'd225} : s = 430;
	{8'd205,8'd226} : s = 431;
	{8'd205,8'd227} : s = 432;
	{8'd205,8'd228} : s = 433;
	{8'd205,8'd229} : s = 434;
	{8'd205,8'd230} : s = 435;
	{8'd205,8'd231} : s = 436;
	{8'd205,8'd232} : s = 437;
	{8'd205,8'd233} : s = 438;
	{8'd205,8'd234} : s = 439;
	{8'd205,8'd235} : s = 440;
	{8'd205,8'd236} : s = 441;
	{8'd205,8'd237} : s = 442;
	{8'd205,8'd238} : s = 443;
	{8'd205,8'd239} : s = 444;
	{8'd205,8'd240} : s = 445;
	{8'd205,8'd241} : s = 446;
	{8'd205,8'd242} : s = 447;
	{8'd205,8'd243} : s = 448;
	{8'd205,8'd244} : s = 449;
	{8'd205,8'd245} : s = 450;
	{8'd205,8'd246} : s = 451;
	{8'd205,8'd247} : s = 452;
	{8'd205,8'd248} : s = 453;
	{8'd205,8'd249} : s = 454;
	{8'd205,8'd250} : s = 455;
	{8'd205,8'd251} : s = 456;
	{8'd205,8'd252} : s = 457;
	{8'd205,8'd253} : s = 458;
	{8'd205,8'd254} : s = 459;
	{8'd205,8'd255} : s = 460;
	{8'd206,8'd0} : s = 206;
	{8'd206,8'd1} : s = 207;
	{8'd206,8'd2} : s = 208;
	{8'd206,8'd3} : s = 209;
	{8'd206,8'd4} : s = 210;
	{8'd206,8'd5} : s = 211;
	{8'd206,8'd6} : s = 212;
	{8'd206,8'd7} : s = 213;
	{8'd206,8'd8} : s = 214;
	{8'd206,8'd9} : s = 215;
	{8'd206,8'd10} : s = 216;
	{8'd206,8'd11} : s = 217;
	{8'd206,8'd12} : s = 218;
	{8'd206,8'd13} : s = 219;
	{8'd206,8'd14} : s = 220;
	{8'd206,8'd15} : s = 221;
	{8'd206,8'd16} : s = 222;
	{8'd206,8'd17} : s = 223;
	{8'd206,8'd18} : s = 224;
	{8'd206,8'd19} : s = 225;
	{8'd206,8'd20} : s = 226;
	{8'd206,8'd21} : s = 227;
	{8'd206,8'd22} : s = 228;
	{8'd206,8'd23} : s = 229;
	{8'd206,8'd24} : s = 230;
	{8'd206,8'd25} : s = 231;
	{8'd206,8'd26} : s = 232;
	{8'd206,8'd27} : s = 233;
	{8'd206,8'd28} : s = 234;
	{8'd206,8'd29} : s = 235;
	{8'd206,8'd30} : s = 236;
	{8'd206,8'd31} : s = 237;
	{8'd206,8'd32} : s = 238;
	{8'd206,8'd33} : s = 239;
	{8'd206,8'd34} : s = 240;
	{8'd206,8'd35} : s = 241;
	{8'd206,8'd36} : s = 242;
	{8'd206,8'd37} : s = 243;
	{8'd206,8'd38} : s = 244;
	{8'd206,8'd39} : s = 245;
	{8'd206,8'd40} : s = 246;
	{8'd206,8'd41} : s = 247;
	{8'd206,8'd42} : s = 248;
	{8'd206,8'd43} : s = 249;
	{8'd206,8'd44} : s = 250;
	{8'd206,8'd45} : s = 251;
	{8'd206,8'd46} : s = 252;
	{8'd206,8'd47} : s = 253;
	{8'd206,8'd48} : s = 254;
	{8'd206,8'd49} : s = 255;
	{8'd206,8'd50} : s = 256;
	{8'd206,8'd51} : s = 257;
	{8'd206,8'd52} : s = 258;
	{8'd206,8'd53} : s = 259;
	{8'd206,8'd54} : s = 260;
	{8'd206,8'd55} : s = 261;
	{8'd206,8'd56} : s = 262;
	{8'd206,8'd57} : s = 263;
	{8'd206,8'd58} : s = 264;
	{8'd206,8'd59} : s = 265;
	{8'd206,8'd60} : s = 266;
	{8'd206,8'd61} : s = 267;
	{8'd206,8'd62} : s = 268;
	{8'd206,8'd63} : s = 269;
	{8'd206,8'd64} : s = 270;
	{8'd206,8'd65} : s = 271;
	{8'd206,8'd66} : s = 272;
	{8'd206,8'd67} : s = 273;
	{8'd206,8'd68} : s = 274;
	{8'd206,8'd69} : s = 275;
	{8'd206,8'd70} : s = 276;
	{8'd206,8'd71} : s = 277;
	{8'd206,8'd72} : s = 278;
	{8'd206,8'd73} : s = 279;
	{8'd206,8'd74} : s = 280;
	{8'd206,8'd75} : s = 281;
	{8'd206,8'd76} : s = 282;
	{8'd206,8'd77} : s = 283;
	{8'd206,8'd78} : s = 284;
	{8'd206,8'd79} : s = 285;
	{8'd206,8'd80} : s = 286;
	{8'd206,8'd81} : s = 287;
	{8'd206,8'd82} : s = 288;
	{8'd206,8'd83} : s = 289;
	{8'd206,8'd84} : s = 290;
	{8'd206,8'd85} : s = 291;
	{8'd206,8'd86} : s = 292;
	{8'd206,8'd87} : s = 293;
	{8'd206,8'd88} : s = 294;
	{8'd206,8'd89} : s = 295;
	{8'd206,8'd90} : s = 296;
	{8'd206,8'd91} : s = 297;
	{8'd206,8'd92} : s = 298;
	{8'd206,8'd93} : s = 299;
	{8'd206,8'd94} : s = 300;
	{8'd206,8'd95} : s = 301;
	{8'd206,8'd96} : s = 302;
	{8'd206,8'd97} : s = 303;
	{8'd206,8'd98} : s = 304;
	{8'd206,8'd99} : s = 305;
	{8'd206,8'd100} : s = 306;
	{8'd206,8'd101} : s = 307;
	{8'd206,8'd102} : s = 308;
	{8'd206,8'd103} : s = 309;
	{8'd206,8'd104} : s = 310;
	{8'd206,8'd105} : s = 311;
	{8'd206,8'd106} : s = 312;
	{8'd206,8'd107} : s = 313;
	{8'd206,8'd108} : s = 314;
	{8'd206,8'd109} : s = 315;
	{8'd206,8'd110} : s = 316;
	{8'd206,8'd111} : s = 317;
	{8'd206,8'd112} : s = 318;
	{8'd206,8'd113} : s = 319;
	{8'd206,8'd114} : s = 320;
	{8'd206,8'd115} : s = 321;
	{8'd206,8'd116} : s = 322;
	{8'd206,8'd117} : s = 323;
	{8'd206,8'd118} : s = 324;
	{8'd206,8'd119} : s = 325;
	{8'd206,8'd120} : s = 326;
	{8'd206,8'd121} : s = 327;
	{8'd206,8'd122} : s = 328;
	{8'd206,8'd123} : s = 329;
	{8'd206,8'd124} : s = 330;
	{8'd206,8'd125} : s = 331;
	{8'd206,8'd126} : s = 332;
	{8'd206,8'd127} : s = 333;
	{8'd206,8'd128} : s = 334;
	{8'd206,8'd129} : s = 335;
	{8'd206,8'd130} : s = 336;
	{8'd206,8'd131} : s = 337;
	{8'd206,8'd132} : s = 338;
	{8'd206,8'd133} : s = 339;
	{8'd206,8'd134} : s = 340;
	{8'd206,8'd135} : s = 341;
	{8'd206,8'd136} : s = 342;
	{8'd206,8'd137} : s = 343;
	{8'd206,8'd138} : s = 344;
	{8'd206,8'd139} : s = 345;
	{8'd206,8'd140} : s = 346;
	{8'd206,8'd141} : s = 347;
	{8'd206,8'd142} : s = 348;
	{8'd206,8'd143} : s = 349;
	{8'd206,8'd144} : s = 350;
	{8'd206,8'd145} : s = 351;
	{8'd206,8'd146} : s = 352;
	{8'd206,8'd147} : s = 353;
	{8'd206,8'd148} : s = 354;
	{8'd206,8'd149} : s = 355;
	{8'd206,8'd150} : s = 356;
	{8'd206,8'd151} : s = 357;
	{8'd206,8'd152} : s = 358;
	{8'd206,8'd153} : s = 359;
	{8'd206,8'd154} : s = 360;
	{8'd206,8'd155} : s = 361;
	{8'd206,8'd156} : s = 362;
	{8'd206,8'd157} : s = 363;
	{8'd206,8'd158} : s = 364;
	{8'd206,8'd159} : s = 365;
	{8'd206,8'd160} : s = 366;
	{8'd206,8'd161} : s = 367;
	{8'd206,8'd162} : s = 368;
	{8'd206,8'd163} : s = 369;
	{8'd206,8'd164} : s = 370;
	{8'd206,8'd165} : s = 371;
	{8'd206,8'd166} : s = 372;
	{8'd206,8'd167} : s = 373;
	{8'd206,8'd168} : s = 374;
	{8'd206,8'd169} : s = 375;
	{8'd206,8'd170} : s = 376;
	{8'd206,8'd171} : s = 377;
	{8'd206,8'd172} : s = 378;
	{8'd206,8'd173} : s = 379;
	{8'd206,8'd174} : s = 380;
	{8'd206,8'd175} : s = 381;
	{8'd206,8'd176} : s = 382;
	{8'd206,8'd177} : s = 383;
	{8'd206,8'd178} : s = 384;
	{8'd206,8'd179} : s = 385;
	{8'd206,8'd180} : s = 386;
	{8'd206,8'd181} : s = 387;
	{8'd206,8'd182} : s = 388;
	{8'd206,8'd183} : s = 389;
	{8'd206,8'd184} : s = 390;
	{8'd206,8'd185} : s = 391;
	{8'd206,8'd186} : s = 392;
	{8'd206,8'd187} : s = 393;
	{8'd206,8'd188} : s = 394;
	{8'd206,8'd189} : s = 395;
	{8'd206,8'd190} : s = 396;
	{8'd206,8'd191} : s = 397;
	{8'd206,8'd192} : s = 398;
	{8'd206,8'd193} : s = 399;
	{8'd206,8'd194} : s = 400;
	{8'd206,8'd195} : s = 401;
	{8'd206,8'd196} : s = 402;
	{8'd206,8'd197} : s = 403;
	{8'd206,8'd198} : s = 404;
	{8'd206,8'd199} : s = 405;
	{8'd206,8'd200} : s = 406;
	{8'd206,8'd201} : s = 407;
	{8'd206,8'd202} : s = 408;
	{8'd206,8'd203} : s = 409;
	{8'd206,8'd204} : s = 410;
	{8'd206,8'd205} : s = 411;
	{8'd206,8'd206} : s = 412;
	{8'd206,8'd207} : s = 413;
	{8'd206,8'd208} : s = 414;
	{8'd206,8'd209} : s = 415;
	{8'd206,8'd210} : s = 416;
	{8'd206,8'd211} : s = 417;
	{8'd206,8'd212} : s = 418;
	{8'd206,8'd213} : s = 419;
	{8'd206,8'd214} : s = 420;
	{8'd206,8'd215} : s = 421;
	{8'd206,8'd216} : s = 422;
	{8'd206,8'd217} : s = 423;
	{8'd206,8'd218} : s = 424;
	{8'd206,8'd219} : s = 425;
	{8'd206,8'd220} : s = 426;
	{8'd206,8'd221} : s = 427;
	{8'd206,8'd222} : s = 428;
	{8'd206,8'd223} : s = 429;
	{8'd206,8'd224} : s = 430;
	{8'd206,8'd225} : s = 431;
	{8'd206,8'd226} : s = 432;
	{8'd206,8'd227} : s = 433;
	{8'd206,8'd228} : s = 434;
	{8'd206,8'd229} : s = 435;
	{8'd206,8'd230} : s = 436;
	{8'd206,8'd231} : s = 437;
	{8'd206,8'd232} : s = 438;
	{8'd206,8'd233} : s = 439;
	{8'd206,8'd234} : s = 440;
	{8'd206,8'd235} : s = 441;
	{8'd206,8'd236} : s = 442;
	{8'd206,8'd237} : s = 443;
	{8'd206,8'd238} : s = 444;
	{8'd206,8'd239} : s = 445;
	{8'd206,8'd240} : s = 446;
	{8'd206,8'd241} : s = 447;
	{8'd206,8'd242} : s = 448;
	{8'd206,8'd243} : s = 449;
	{8'd206,8'd244} : s = 450;
	{8'd206,8'd245} : s = 451;
	{8'd206,8'd246} : s = 452;
	{8'd206,8'd247} : s = 453;
	{8'd206,8'd248} : s = 454;
	{8'd206,8'd249} : s = 455;
	{8'd206,8'd250} : s = 456;
	{8'd206,8'd251} : s = 457;
	{8'd206,8'd252} : s = 458;
	{8'd206,8'd253} : s = 459;
	{8'd206,8'd254} : s = 460;
	{8'd206,8'd255} : s = 461;
	{8'd207,8'd0} : s = 207;
	{8'd207,8'd1} : s = 208;
	{8'd207,8'd2} : s = 209;
	{8'd207,8'd3} : s = 210;
	{8'd207,8'd4} : s = 211;
	{8'd207,8'd5} : s = 212;
	{8'd207,8'd6} : s = 213;
	{8'd207,8'd7} : s = 214;
	{8'd207,8'd8} : s = 215;
	{8'd207,8'd9} : s = 216;
	{8'd207,8'd10} : s = 217;
	{8'd207,8'd11} : s = 218;
	{8'd207,8'd12} : s = 219;
	{8'd207,8'd13} : s = 220;
	{8'd207,8'd14} : s = 221;
	{8'd207,8'd15} : s = 222;
	{8'd207,8'd16} : s = 223;
	{8'd207,8'd17} : s = 224;
	{8'd207,8'd18} : s = 225;
	{8'd207,8'd19} : s = 226;
	{8'd207,8'd20} : s = 227;
	{8'd207,8'd21} : s = 228;
	{8'd207,8'd22} : s = 229;
	{8'd207,8'd23} : s = 230;
	{8'd207,8'd24} : s = 231;
	{8'd207,8'd25} : s = 232;
	{8'd207,8'd26} : s = 233;
	{8'd207,8'd27} : s = 234;
	{8'd207,8'd28} : s = 235;
	{8'd207,8'd29} : s = 236;
	{8'd207,8'd30} : s = 237;
	{8'd207,8'd31} : s = 238;
	{8'd207,8'd32} : s = 239;
	{8'd207,8'd33} : s = 240;
	{8'd207,8'd34} : s = 241;
	{8'd207,8'd35} : s = 242;
	{8'd207,8'd36} : s = 243;
	{8'd207,8'd37} : s = 244;
	{8'd207,8'd38} : s = 245;
	{8'd207,8'd39} : s = 246;
	{8'd207,8'd40} : s = 247;
	{8'd207,8'd41} : s = 248;
	{8'd207,8'd42} : s = 249;
	{8'd207,8'd43} : s = 250;
	{8'd207,8'd44} : s = 251;
	{8'd207,8'd45} : s = 252;
	{8'd207,8'd46} : s = 253;
	{8'd207,8'd47} : s = 254;
	{8'd207,8'd48} : s = 255;
	{8'd207,8'd49} : s = 256;
	{8'd207,8'd50} : s = 257;
	{8'd207,8'd51} : s = 258;
	{8'd207,8'd52} : s = 259;
	{8'd207,8'd53} : s = 260;
	{8'd207,8'd54} : s = 261;
	{8'd207,8'd55} : s = 262;
	{8'd207,8'd56} : s = 263;
	{8'd207,8'd57} : s = 264;
	{8'd207,8'd58} : s = 265;
	{8'd207,8'd59} : s = 266;
	{8'd207,8'd60} : s = 267;
	{8'd207,8'd61} : s = 268;
	{8'd207,8'd62} : s = 269;
	{8'd207,8'd63} : s = 270;
	{8'd207,8'd64} : s = 271;
	{8'd207,8'd65} : s = 272;
	{8'd207,8'd66} : s = 273;
	{8'd207,8'd67} : s = 274;
	{8'd207,8'd68} : s = 275;
	{8'd207,8'd69} : s = 276;
	{8'd207,8'd70} : s = 277;
	{8'd207,8'd71} : s = 278;
	{8'd207,8'd72} : s = 279;
	{8'd207,8'd73} : s = 280;
	{8'd207,8'd74} : s = 281;
	{8'd207,8'd75} : s = 282;
	{8'd207,8'd76} : s = 283;
	{8'd207,8'd77} : s = 284;
	{8'd207,8'd78} : s = 285;
	{8'd207,8'd79} : s = 286;
	{8'd207,8'd80} : s = 287;
	{8'd207,8'd81} : s = 288;
	{8'd207,8'd82} : s = 289;
	{8'd207,8'd83} : s = 290;
	{8'd207,8'd84} : s = 291;
	{8'd207,8'd85} : s = 292;
	{8'd207,8'd86} : s = 293;
	{8'd207,8'd87} : s = 294;
	{8'd207,8'd88} : s = 295;
	{8'd207,8'd89} : s = 296;
	{8'd207,8'd90} : s = 297;
	{8'd207,8'd91} : s = 298;
	{8'd207,8'd92} : s = 299;
	{8'd207,8'd93} : s = 300;
	{8'd207,8'd94} : s = 301;
	{8'd207,8'd95} : s = 302;
	{8'd207,8'd96} : s = 303;
	{8'd207,8'd97} : s = 304;
	{8'd207,8'd98} : s = 305;
	{8'd207,8'd99} : s = 306;
	{8'd207,8'd100} : s = 307;
	{8'd207,8'd101} : s = 308;
	{8'd207,8'd102} : s = 309;
	{8'd207,8'd103} : s = 310;
	{8'd207,8'd104} : s = 311;
	{8'd207,8'd105} : s = 312;
	{8'd207,8'd106} : s = 313;
	{8'd207,8'd107} : s = 314;
	{8'd207,8'd108} : s = 315;
	{8'd207,8'd109} : s = 316;
	{8'd207,8'd110} : s = 317;
	{8'd207,8'd111} : s = 318;
	{8'd207,8'd112} : s = 319;
	{8'd207,8'd113} : s = 320;
	{8'd207,8'd114} : s = 321;
	{8'd207,8'd115} : s = 322;
	{8'd207,8'd116} : s = 323;
	{8'd207,8'd117} : s = 324;
	{8'd207,8'd118} : s = 325;
	{8'd207,8'd119} : s = 326;
	{8'd207,8'd120} : s = 327;
	{8'd207,8'd121} : s = 328;
	{8'd207,8'd122} : s = 329;
	{8'd207,8'd123} : s = 330;
	{8'd207,8'd124} : s = 331;
	{8'd207,8'd125} : s = 332;
	{8'd207,8'd126} : s = 333;
	{8'd207,8'd127} : s = 334;
	{8'd207,8'd128} : s = 335;
	{8'd207,8'd129} : s = 336;
	{8'd207,8'd130} : s = 337;
	{8'd207,8'd131} : s = 338;
	{8'd207,8'd132} : s = 339;
	{8'd207,8'd133} : s = 340;
	{8'd207,8'd134} : s = 341;
	{8'd207,8'd135} : s = 342;
	{8'd207,8'd136} : s = 343;
	{8'd207,8'd137} : s = 344;
	{8'd207,8'd138} : s = 345;
	{8'd207,8'd139} : s = 346;
	{8'd207,8'd140} : s = 347;
	{8'd207,8'd141} : s = 348;
	{8'd207,8'd142} : s = 349;
	{8'd207,8'd143} : s = 350;
	{8'd207,8'd144} : s = 351;
	{8'd207,8'd145} : s = 352;
	{8'd207,8'd146} : s = 353;
	{8'd207,8'd147} : s = 354;
	{8'd207,8'd148} : s = 355;
	{8'd207,8'd149} : s = 356;
	{8'd207,8'd150} : s = 357;
	{8'd207,8'd151} : s = 358;
	{8'd207,8'd152} : s = 359;
	{8'd207,8'd153} : s = 360;
	{8'd207,8'd154} : s = 361;
	{8'd207,8'd155} : s = 362;
	{8'd207,8'd156} : s = 363;
	{8'd207,8'd157} : s = 364;
	{8'd207,8'd158} : s = 365;
	{8'd207,8'd159} : s = 366;
	{8'd207,8'd160} : s = 367;
	{8'd207,8'd161} : s = 368;
	{8'd207,8'd162} : s = 369;
	{8'd207,8'd163} : s = 370;
	{8'd207,8'd164} : s = 371;
	{8'd207,8'd165} : s = 372;
	{8'd207,8'd166} : s = 373;
	{8'd207,8'd167} : s = 374;
	{8'd207,8'd168} : s = 375;
	{8'd207,8'd169} : s = 376;
	{8'd207,8'd170} : s = 377;
	{8'd207,8'd171} : s = 378;
	{8'd207,8'd172} : s = 379;
	{8'd207,8'd173} : s = 380;
	{8'd207,8'd174} : s = 381;
	{8'd207,8'd175} : s = 382;
	{8'd207,8'd176} : s = 383;
	{8'd207,8'd177} : s = 384;
	{8'd207,8'd178} : s = 385;
	{8'd207,8'd179} : s = 386;
	{8'd207,8'd180} : s = 387;
	{8'd207,8'd181} : s = 388;
	{8'd207,8'd182} : s = 389;
	{8'd207,8'd183} : s = 390;
	{8'd207,8'd184} : s = 391;
	{8'd207,8'd185} : s = 392;
	{8'd207,8'd186} : s = 393;
	{8'd207,8'd187} : s = 394;
	{8'd207,8'd188} : s = 395;
	{8'd207,8'd189} : s = 396;
	{8'd207,8'd190} : s = 397;
	{8'd207,8'd191} : s = 398;
	{8'd207,8'd192} : s = 399;
	{8'd207,8'd193} : s = 400;
	{8'd207,8'd194} : s = 401;
	{8'd207,8'd195} : s = 402;
	{8'd207,8'd196} : s = 403;
	{8'd207,8'd197} : s = 404;
	{8'd207,8'd198} : s = 405;
	{8'd207,8'd199} : s = 406;
	{8'd207,8'd200} : s = 407;
	{8'd207,8'd201} : s = 408;
	{8'd207,8'd202} : s = 409;
	{8'd207,8'd203} : s = 410;
	{8'd207,8'd204} : s = 411;
	{8'd207,8'd205} : s = 412;
	{8'd207,8'd206} : s = 413;
	{8'd207,8'd207} : s = 414;
	{8'd207,8'd208} : s = 415;
	{8'd207,8'd209} : s = 416;
	{8'd207,8'd210} : s = 417;
	{8'd207,8'd211} : s = 418;
	{8'd207,8'd212} : s = 419;
	{8'd207,8'd213} : s = 420;
	{8'd207,8'd214} : s = 421;
	{8'd207,8'd215} : s = 422;
	{8'd207,8'd216} : s = 423;
	{8'd207,8'd217} : s = 424;
	{8'd207,8'd218} : s = 425;
	{8'd207,8'd219} : s = 426;
	{8'd207,8'd220} : s = 427;
	{8'd207,8'd221} : s = 428;
	{8'd207,8'd222} : s = 429;
	{8'd207,8'd223} : s = 430;
	{8'd207,8'd224} : s = 431;
	{8'd207,8'd225} : s = 432;
	{8'd207,8'd226} : s = 433;
	{8'd207,8'd227} : s = 434;
	{8'd207,8'd228} : s = 435;
	{8'd207,8'd229} : s = 436;
	{8'd207,8'd230} : s = 437;
	{8'd207,8'd231} : s = 438;
	{8'd207,8'd232} : s = 439;
	{8'd207,8'd233} : s = 440;
	{8'd207,8'd234} : s = 441;
	{8'd207,8'd235} : s = 442;
	{8'd207,8'd236} : s = 443;
	{8'd207,8'd237} : s = 444;
	{8'd207,8'd238} : s = 445;
	{8'd207,8'd239} : s = 446;
	{8'd207,8'd240} : s = 447;
	{8'd207,8'd241} : s = 448;
	{8'd207,8'd242} : s = 449;
	{8'd207,8'd243} : s = 450;
	{8'd207,8'd244} : s = 451;
	{8'd207,8'd245} : s = 452;
	{8'd207,8'd246} : s = 453;
	{8'd207,8'd247} : s = 454;
	{8'd207,8'd248} : s = 455;
	{8'd207,8'd249} : s = 456;
	{8'd207,8'd250} : s = 457;
	{8'd207,8'd251} : s = 458;
	{8'd207,8'd252} : s = 459;
	{8'd207,8'd253} : s = 460;
	{8'd207,8'd254} : s = 461;
	{8'd207,8'd255} : s = 462;
	{8'd208,8'd0} : s = 208;
	{8'd208,8'd1} : s = 209;
	{8'd208,8'd2} : s = 210;
	{8'd208,8'd3} : s = 211;
	{8'd208,8'd4} : s = 212;
	{8'd208,8'd5} : s = 213;
	{8'd208,8'd6} : s = 214;
	{8'd208,8'd7} : s = 215;
	{8'd208,8'd8} : s = 216;
	{8'd208,8'd9} : s = 217;
	{8'd208,8'd10} : s = 218;
	{8'd208,8'd11} : s = 219;
	{8'd208,8'd12} : s = 220;
	{8'd208,8'd13} : s = 221;
	{8'd208,8'd14} : s = 222;
	{8'd208,8'd15} : s = 223;
	{8'd208,8'd16} : s = 224;
	{8'd208,8'd17} : s = 225;
	{8'd208,8'd18} : s = 226;
	{8'd208,8'd19} : s = 227;
	{8'd208,8'd20} : s = 228;
	{8'd208,8'd21} : s = 229;
	{8'd208,8'd22} : s = 230;
	{8'd208,8'd23} : s = 231;
	{8'd208,8'd24} : s = 232;
	{8'd208,8'd25} : s = 233;
	{8'd208,8'd26} : s = 234;
	{8'd208,8'd27} : s = 235;
	{8'd208,8'd28} : s = 236;
	{8'd208,8'd29} : s = 237;
	{8'd208,8'd30} : s = 238;
	{8'd208,8'd31} : s = 239;
	{8'd208,8'd32} : s = 240;
	{8'd208,8'd33} : s = 241;
	{8'd208,8'd34} : s = 242;
	{8'd208,8'd35} : s = 243;
	{8'd208,8'd36} : s = 244;
	{8'd208,8'd37} : s = 245;
	{8'd208,8'd38} : s = 246;
	{8'd208,8'd39} : s = 247;
	{8'd208,8'd40} : s = 248;
	{8'd208,8'd41} : s = 249;
	{8'd208,8'd42} : s = 250;
	{8'd208,8'd43} : s = 251;
	{8'd208,8'd44} : s = 252;
	{8'd208,8'd45} : s = 253;
	{8'd208,8'd46} : s = 254;
	{8'd208,8'd47} : s = 255;
	{8'd208,8'd48} : s = 256;
	{8'd208,8'd49} : s = 257;
	{8'd208,8'd50} : s = 258;
	{8'd208,8'd51} : s = 259;
	{8'd208,8'd52} : s = 260;
	{8'd208,8'd53} : s = 261;
	{8'd208,8'd54} : s = 262;
	{8'd208,8'd55} : s = 263;
	{8'd208,8'd56} : s = 264;
	{8'd208,8'd57} : s = 265;
	{8'd208,8'd58} : s = 266;
	{8'd208,8'd59} : s = 267;
	{8'd208,8'd60} : s = 268;
	{8'd208,8'd61} : s = 269;
	{8'd208,8'd62} : s = 270;
	{8'd208,8'd63} : s = 271;
	{8'd208,8'd64} : s = 272;
	{8'd208,8'd65} : s = 273;
	{8'd208,8'd66} : s = 274;
	{8'd208,8'd67} : s = 275;
	{8'd208,8'd68} : s = 276;
	{8'd208,8'd69} : s = 277;
	{8'd208,8'd70} : s = 278;
	{8'd208,8'd71} : s = 279;
	{8'd208,8'd72} : s = 280;
	{8'd208,8'd73} : s = 281;
	{8'd208,8'd74} : s = 282;
	{8'd208,8'd75} : s = 283;
	{8'd208,8'd76} : s = 284;
	{8'd208,8'd77} : s = 285;
	{8'd208,8'd78} : s = 286;
	{8'd208,8'd79} : s = 287;
	{8'd208,8'd80} : s = 288;
	{8'd208,8'd81} : s = 289;
	{8'd208,8'd82} : s = 290;
	{8'd208,8'd83} : s = 291;
	{8'd208,8'd84} : s = 292;
	{8'd208,8'd85} : s = 293;
	{8'd208,8'd86} : s = 294;
	{8'd208,8'd87} : s = 295;
	{8'd208,8'd88} : s = 296;
	{8'd208,8'd89} : s = 297;
	{8'd208,8'd90} : s = 298;
	{8'd208,8'd91} : s = 299;
	{8'd208,8'd92} : s = 300;
	{8'd208,8'd93} : s = 301;
	{8'd208,8'd94} : s = 302;
	{8'd208,8'd95} : s = 303;
	{8'd208,8'd96} : s = 304;
	{8'd208,8'd97} : s = 305;
	{8'd208,8'd98} : s = 306;
	{8'd208,8'd99} : s = 307;
	{8'd208,8'd100} : s = 308;
	{8'd208,8'd101} : s = 309;
	{8'd208,8'd102} : s = 310;
	{8'd208,8'd103} : s = 311;
	{8'd208,8'd104} : s = 312;
	{8'd208,8'd105} : s = 313;
	{8'd208,8'd106} : s = 314;
	{8'd208,8'd107} : s = 315;
	{8'd208,8'd108} : s = 316;
	{8'd208,8'd109} : s = 317;
	{8'd208,8'd110} : s = 318;
	{8'd208,8'd111} : s = 319;
	{8'd208,8'd112} : s = 320;
	{8'd208,8'd113} : s = 321;
	{8'd208,8'd114} : s = 322;
	{8'd208,8'd115} : s = 323;
	{8'd208,8'd116} : s = 324;
	{8'd208,8'd117} : s = 325;
	{8'd208,8'd118} : s = 326;
	{8'd208,8'd119} : s = 327;
	{8'd208,8'd120} : s = 328;
	{8'd208,8'd121} : s = 329;
	{8'd208,8'd122} : s = 330;
	{8'd208,8'd123} : s = 331;
	{8'd208,8'd124} : s = 332;
	{8'd208,8'd125} : s = 333;
	{8'd208,8'd126} : s = 334;
	{8'd208,8'd127} : s = 335;
	{8'd208,8'd128} : s = 336;
	{8'd208,8'd129} : s = 337;
	{8'd208,8'd130} : s = 338;
	{8'd208,8'd131} : s = 339;
	{8'd208,8'd132} : s = 340;
	{8'd208,8'd133} : s = 341;
	{8'd208,8'd134} : s = 342;
	{8'd208,8'd135} : s = 343;
	{8'd208,8'd136} : s = 344;
	{8'd208,8'd137} : s = 345;
	{8'd208,8'd138} : s = 346;
	{8'd208,8'd139} : s = 347;
	{8'd208,8'd140} : s = 348;
	{8'd208,8'd141} : s = 349;
	{8'd208,8'd142} : s = 350;
	{8'd208,8'd143} : s = 351;
	{8'd208,8'd144} : s = 352;
	{8'd208,8'd145} : s = 353;
	{8'd208,8'd146} : s = 354;
	{8'd208,8'd147} : s = 355;
	{8'd208,8'd148} : s = 356;
	{8'd208,8'd149} : s = 357;
	{8'd208,8'd150} : s = 358;
	{8'd208,8'd151} : s = 359;
	{8'd208,8'd152} : s = 360;
	{8'd208,8'd153} : s = 361;
	{8'd208,8'd154} : s = 362;
	{8'd208,8'd155} : s = 363;
	{8'd208,8'd156} : s = 364;
	{8'd208,8'd157} : s = 365;
	{8'd208,8'd158} : s = 366;
	{8'd208,8'd159} : s = 367;
	{8'd208,8'd160} : s = 368;
	{8'd208,8'd161} : s = 369;
	{8'd208,8'd162} : s = 370;
	{8'd208,8'd163} : s = 371;
	{8'd208,8'd164} : s = 372;
	{8'd208,8'd165} : s = 373;
	{8'd208,8'd166} : s = 374;
	{8'd208,8'd167} : s = 375;
	{8'd208,8'd168} : s = 376;
	{8'd208,8'd169} : s = 377;
	{8'd208,8'd170} : s = 378;
	{8'd208,8'd171} : s = 379;
	{8'd208,8'd172} : s = 380;
	{8'd208,8'd173} : s = 381;
	{8'd208,8'd174} : s = 382;
	{8'd208,8'd175} : s = 383;
	{8'd208,8'd176} : s = 384;
	{8'd208,8'd177} : s = 385;
	{8'd208,8'd178} : s = 386;
	{8'd208,8'd179} : s = 387;
	{8'd208,8'd180} : s = 388;
	{8'd208,8'd181} : s = 389;
	{8'd208,8'd182} : s = 390;
	{8'd208,8'd183} : s = 391;
	{8'd208,8'd184} : s = 392;
	{8'd208,8'd185} : s = 393;
	{8'd208,8'd186} : s = 394;
	{8'd208,8'd187} : s = 395;
	{8'd208,8'd188} : s = 396;
	{8'd208,8'd189} : s = 397;
	{8'd208,8'd190} : s = 398;
	{8'd208,8'd191} : s = 399;
	{8'd208,8'd192} : s = 400;
	{8'd208,8'd193} : s = 401;
	{8'd208,8'd194} : s = 402;
	{8'd208,8'd195} : s = 403;
	{8'd208,8'd196} : s = 404;
	{8'd208,8'd197} : s = 405;
	{8'd208,8'd198} : s = 406;
	{8'd208,8'd199} : s = 407;
	{8'd208,8'd200} : s = 408;
	{8'd208,8'd201} : s = 409;
	{8'd208,8'd202} : s = 410;
	{8'd208,8'd203} : s = 411;
	{8'd208,8'd204} : s = 412;
	{8'd208,8'd205} : s = 413;
	{8'd208,8'd206} : s = 414;
	{8'd208,8'd207} : s = 415;
	{8'd208,8'd208} : s = 416;
	{8'd208,8'd209} : s = 417;
	{8'd208,8'd210} : s = 418;
	{8'd208,8'd211} : s = 419;
	{8'd208,8'd212} : s = 420;
	{8'd208,8'd213} : s = 421;
	{8'd208,8'd214} : s = 422;
	{8'd208,8'd215} : s = 423;
	{8'd208,8'd216} : s = 424;
	{8'd208,8'd217} : s = 425;
	{8'd208,8'd218} : s = 426;
	{8'd208,8'd219} : s = 427;
	{8'd208,8'd220} : s = 428;
	{8'd208,8'd221} : s = 429;
	{8'd208,8'd222} : s = 430;
	{8'd208,8'd223} : s = 431;
	{8'd208,8'd224} : s = 432;
	{8'd208,8'd225} : s = 433;
	{8'd208,8'd226} : s = 434;
	{8'd208,8'd227} : s = 435;
	{8'd208,8'd228} : s = 436;
	{8'd208,8'd229} : s = 437;
	{8'd208,8'd230} : s = 438;
	{8'd208,8'd231} : s = 439;
	{8'd208,8'd232} : s = 440;
	{8'd208,8'd233} : s = 441;
	{8'd208,8'd234} : s = 442;
	{8'd208,8'd235} : s = 443;
	{8'd208,8'd236} : s = 444;
	{8'd208,8'd237} : s = 445;
	{8'd208,8'd238} : s = 446;
	{8'd208,8'd239} : s = 447;
	{8'd208,8'd240} : s = 448;
	{8'd208,8'd241} : s = 449;
	{8'd208,8'd242} : s = 450;
	{8'd208,8'd243} : s = 451;
	{8'd208,8'd244} : s = 452;
	{8'd208,8'd245} : s = 453;
	{8'd208,8'd246} : s = 454;
	{8'd208,8'd247} : s = 455;
	{8'd208,8'd248} : s = 456;
	{8'd208,8'd249} : s = 457;
	{8'd208,8'd250} : s = 458;
	{8'd208,8'd251} : s = 459;
	{8'd208,8'd252} : s = 460;
	{8'd208,8'd253} : s = 461;
	{8'd208,8'd254} : s = 462;
	{8'd208,8'd255} : s = 463;
	{8'd209,8'd0} : s = 209;
	{8'd209,8'd1} : s = 210;
	{8'd209,8'd2} : s = 211;
	{8'd209,8'd3} : s = 212;
	{8'd209,8'd4} : s = 213;
	{8'd209,8'd5} : s = 214;
	{8'd209,8'd6} : s = 215;
	{8'd209,8'd7} : s = 216;
	{8'd209,8'd8} : s = 217;
	{8'd209,8'd9} : s = 218;
	{8'd209,8'd10} : s = 219;
	{8'd209,8'd11} : s = 220;
	{8'd209,8'd12} : s = 221;
	{8'd209,8'd13} : s = 222;
	{8'd209,8'd14} : s = 223;
	{8'd209,8'd15} : s = 224;
	{8'd209,8'd16} : s = 225;
	{8'd209,8'd17} : s = 226;
	{8'd209,8'd18} : s = 227;
	{8'd209,8'd19} : s = 228;
	{8'd209,8'd20} : s = 229;
	{8'd209,8'd21} : s = 230;
	{8'd209,8'd22} : s = 231;
	{8'd209,8'd23} : s = 232;
	{8'd209,8'd24} : s = 233;
	{8'd209,8'd25} : s = 234;
	{8'd209,8'd26} : s = 235;
	{8'd209,8'd27} : s = 236;
	{8'd209,8'd28} : s = 237;
	{8'd209,8'd29} : s = 238;
	{8'd209,8'd30} : s = 239;
	{8'd209,8'd31} : s = 240;
	{8'd209,8'd32} : s = 241;
	{8'd209,8'd33} : s = 242;
	{8'd209,8'd34} : s = 243;
	{8'd209,8'd35} : s = 244;
	{8'd209,8'd36} : s = 245;
	{8'd209,8'd37} : s = 246;
	{8'd209,8'd38} : s = 247;
	{8'd209,8'd39} : s = 248;
	{8'd209,8'd40} : s = 249;
	{8'd209,8'd41} : s = 250;
	{8'd209,8'd42} : s = 251;
	{8'd209,8'd43} : s = 252;
	{8'd209,8'd44} : s = 253;
	{8'd209,8'd45} : s = 254;
	{8'd209,8'd46} : s = 255;
	{8'd209,8'd47} : s = 256;
	{8'd209,8'd48} : s = 257;
	{8'd209,8'd49} : s = 258;
	{8'd209,8'd50} : s = 259;
	{8'd209,8'd51} : s = 260;
	{8'd209,8'd52} : s = 261;
	{8'd209,8'd53} : s = 262;
	{8'd209,8'd54} : s = 263;
	{8'd209,8'd55} : s = 264;
	{8'd209,8'd56} : s = 265;
	{8'd209,8'd57} : s = 266;
	{8'd209,8'd58} : s = 267;
	{8'd209,8'd59} : s = 268;
	{8'd209,8'd60} : s = 269;
	{8'd209,8'd61} : s = 270;
	{8'd209,8'd62} : s = 271;
	{8'd209,8'd63} : s = 272;
	{8'd209,8'd64} : s = 273;
	{8'd209,8'd65} : s = 274;
	{8'd209,8'd66} : s = 275;
	{8'd209,8'd67} : s = 276;
	{8'd209,8'd68} : s = 277;
	{8'd209,8'd69} : s = 278;
	{8'd209,8'd70} : s = 279;
	{8'd209,8'd71} : s = 280;
	{8'd209,8'd72} : s = 281;
	{8'd209,8'd73} : s = 282;
	{8'd209,8'd74} : s = 283;
	{8'd209,8'd75} : s = 284;
	{8'd209,8'd76} : s = 285;
	{8'd209,8'd77} : s = 286;
	{8'd209,8'd78} : s = 287;
	{8'd209,8'd79} : s = 288;
	{8'd209,8'd80} : s = 289;
	{8'd209,8'd81} : s = 290;
	{8'd209,8'd82} : s = 291;
	{8'd209,8'd83} : s = 292;
	{8'd209,8'd84} : s = 293;
	{8'd209,8'd85} : s = 294;
	{8'd209,8'd86} : s = 295;
	{8'd209,8'd87} : s = 296;
	{8'd209,8'd88} : s = 297;
	{8'd209,8'd89} : s = 298;
	{8'd209,8'd90} : s = 299;
	{8'd209,8'd91} : s = 300;
	{8'd209,8'd92} : s = 301;
	{8'd209,8'd93} : s = 302;
	{8'd209,8'd94} : s = 303;
	{8'd209,8'd95} : s = 304;
	{8'd209,8'd96} : s = 305;
	{8'd209,8'd97} : s = 306;
	{8'd209,8'd98} : s = 307;
	{8'd209,8'd99} : s = 308;
	{8'd209,8'd100} : s = 309;
	{8'd209,8'd101} : s = 310;
	{8'd209,8'd102} : s = 311;
	{8'd209,8'd103} : s = 312;
	{8'd209,8'd104} : s = 313;
	{8'd209,8'd105} : s = 314;
	{8'd209,8'd106} : s = 315;
	{8'd209,8'd107} : s = 316;
	{8'd209,8'd108} : s = 317;
	{8'd209,8'd109} : s = 318;
	{8'd209,8'd110} : s = 319;
	{8'd209,8'd111} : s = 320;
	{8'd209,8'd112} : s = 321;
	{8'd209,8'd113} : s = 322;
	{8'd209,8'd114} : s = 323;
	{8'd209,8'd115} : s = 324;
	{8'd209,8'd116} : s = 325;
	{8'd209,8'd117} : s = 326;
	{8'd209,8'd118} : s = 327;
	{8'd209,8'd119} : s = 328;
	{8'd209,8'd120} : s = 329;
	{8'd209,8'd121} : s = 330;
	{8'd209,8'd122} : s = 331;
	{8'd209,8'd123} : s = 332;
	{8'd209,8'd124} : s = 333;
	{8'd209,8'd125} : s = 334;
	{8'd209,8'd126} : s = 335;
	{8'd209,8'd127} : s = 336;
	{8'd209,8'd128} : s = 337;
	{8'd209,8'd129} : s = 338;
	{8'd209,8'd130} : s = 339;
	{8'd209,8'd131} : s = 340;
	{8'd209,8'd132} : s = 341;
	{8'd209,8'd133} : s = 342;
	{8'd209,8'd134} : s = 343;
	{8'd209,8'd135} : s = 344;
	{8'd209,8'd136} : s = 345;
	{8'd209,8'd137} : s = 346;
	{8'd209,8'd138} : s = 347;
	{8'd209,8'd139} : s = 348;
	{8'd209,8'd140} : s = 349;
	{8'd209,8'd141} : s = 350;
	{8'd209,8'd142} : s = 351;
	{8'd209,8'd143} : s = 352;
	{8'd209,8'd144} : s = 353;
	{8'd209,8'd145} : s = 354;
	{8'd209,8'd146} : s = 355;
	{8'd209,8'd147} : s = 356;
	{8'd209,8'd148} : s = 357;
	{8'd209,8'd149} : s = 358;
	{8'd209,8'd150} : s = 359;
	{8'd209,8'd151} : s = 360;
	{8'd209,8'd152} : s = 361;
	{8'd209,8'd153} : s = 362;
	{8'd209,8'd154} : s = 363;
	{8'd209,8'd155} : s = 364;
	{8'd209,8'd156} : s = 365;
	{8'd209,8'd157} : s = 366;
	{8'd209,8'd158} : s = 367;
	{8'd209,8'd159} : s = 368;
	{8'd209,8'd160} : s = 369;
	{8'd209,8'd161} : s = 370;
	{8'd209,8'd162} : s = 371;
	{8'd209,8'd163} : s = 372;
	{8'd209,8'd164} : s = 373;
	{8'd209,8'd165} : s = 374;
	{8'd209,8'd166} : s = 375;
	{8'd209,8'd167} : s = 376;
	{8'd209,8'd168} : s = 377;
	{8'd209,8'd169} : s = 378;
	{8'd209,8'd170} : s = 379;
	{8'd209,8'd171} : s = 380;
	{8'd209,8'd172} : s = 381;
	{8'd209,8'd173} : s = 382;
	{8'd209,8'd174} : s = 383;
	{8'd209,8'd175} : s = 384;
	{8'd209,8'd176} : s = 385;
	{8'd209,8'd177} : s = 386;
	{8'd209,8'd178} : s = 387;
	{8'd209,8'd179} : s = 388;
	{8'd209,8'd180} : s = 389;
	{8'd209,8'd181} : s = 390;
	{8'd209,8'd182} : s = 391;
	{8'd209,8'd183} : s = 392;
	{8'd209,8'd184} : s = 393;
	{8'd209,8'd185} : s = 394;
	{8'd209,8'd186} : s = 395;
	{8'd209,8'd187} : s = 396;
	{8'd209,8'd188} : s = 397;
	{8'd209,8'd189} : s = 398;
	{8'd209,8'd190} : s = 399;
	{8'd209,8'd191} : s = 400;
	{8'd209,8'd192} : s = 401;
	{8'd209,8'd193} : s = 402;
	{8'd209,8'd194} : s = 403;
	{8'd209,8'd195} : s = 404;
	{8'd209,8'd196} : s = 405;
	{8'd209,8'd197} : s = 406;
	{8'd209,8'd198} : s = 407;
	{8'd209,8'd199} : s = 408;
	{8'd209,8'd200} : s = 409;
	{8'd209,8'd201} : s = 410;
	{8'd209,8'd202} : s = 411;
	{8'd209,8'd203} : s = 412;
	{8'd209,8'd204} : s = 413;
	{8'd209,8'd205} : s = 414;
	{8'd209,8'd206} : s = 415;
	{8'd209,8'd207} : s = 416;
	{8'd209,8'd208} : s = 417;
	{8'd209,8'd209} : s = 418;
	{8'd209,8'd210} : s = 419;
	{8'd209,8'd211} : s = 420;
	{8'd209,8'd212} : s = 421;
	{8'd209,8'd213} : s = 422;
	{8'd209,8'd214} : s = 423;
	{8'd209,8'd215} : s = 424;
	{8'd209,8'd216} : s = 425;
	{8'd209,8'd217} : s = 426;
	{8'd209,8'd218} : s = 427;
	{8'd209,8'd219} : s = 428;
	{8'd209,8'd220} : s = 429;
	{8'd209,8'd221} : s = 430;
	{8'd209,8'd222} : s = 431;
	{8'd209,8'd223} : s = 432;
	{8'd209,8'd224} : s = 433;
	{8'd209,8'd225} : s = 434;
	{8'd209,8'd226} : s = 435;
	{8'd209,8'd227} : s = 436;
	{8'd209,8'd228} : s = 437;
	{8'd209,8'd229} : s = 438;
	{8'd209,8'd230} : s = 439;
	{8'd209,8'd231} : s = 440;
	{8'd209,8'd232} : s = 441;
	{8'd209,8'd233} : s = 442;
	{8'd209,8'd234} : s = 443;
	{8'd209,8'd235} : s = 444;
	{8'd209,8'd236} : s = 445;
	{8'd209,8'd237} : s = 446;
	{8'd209,8'd238} : s = 447;
	{8'd209,8'd239} : s = 448;
	{8'd209,8'd240} : s = 449;
	{8'd209,8'd241} : s = 450;
	{8'd209,8'd242} : s = 451;
	{8'd209,8'd243} : s = 452;
	{8'd209,8'd244} : s = 453;
	{8'd209,8'd245} : s = 454;
	{8'd209,8'd246} : s = 455;
	{8'd209,8'd247} : s = 456;
	{8'd209,8'd248} : s = 457;
	{8'd209,8'd249} : s = 458;
	{8'd209,8'd250} : s = 459;
	{8'd209,8'd251} : s = 460;
	{8'd209,8'd252} : s = 461;
	{8'd209,8'd253} : s = 462;
	{8'd209,8'd254} : s = 463;
	{8'd209,8'd255} : s = 464;
	{8'd210,8'd0} : s = 210;
	{8'd210,8'd1} : s = 211;
	{8'd210,8'd2} : s = 212;
	{8'd210,8'd3} : s = 213;
	{8'd210,8'd4} : s = 214;
	{8'd210,8'd5} : s = 215;
	{8'd210,8'd6} : s = 216;
	{8'd210,8'd7} : s = 217;
	{8'd210,8'd8} : s = 218;
	{8'd210,8'd9} : s = 219;
	{8'd210,8'd10} : s = 220;
	{8'd210,8'd11} : s = 221;
	{8'd210,8'd12} : s = 222;
	{8'd210,8'd13} : s = 223;
	{8'd210,8'd14} : s = 224;
	{8'd210,8'd15} : s = 225;
	{8'd210,8'd16} : s = 226;
	{8'd210,8'd17} : s = 227;
	{8'd210,8'd18} : s = 228;
	{8'd210,8'd19} : s = 229;
	{8'd210,8'd20} : s = 230;
	{8'd210,8'd21} : s = 231;
	{8'd210,8'd22} : s = 232;
	{8'd210,8'd23} : s = 233;
	{8'd210,8'd24} : s = 234;
	{8'd210,8'd25} : s = 235;
	{8'd210,8'd26} : s = 236;
	{8'd210,8'd27} : s = 237;
	{8'd210,8'd28} : s = 238;
	{8'd210,8'd29} : s = 239;
	{8'd210,8'd30} : s = 240;
	{8'd210,8'd31} : s = 241;
	{8'd210,8'd32} : s = 242;
	{8'd210,8'd33} : s = 243;
	{8'd210,8'd34} : s = 244;
	{8'd210,8'd35} : s = 245;
	{8'd210,8'd36} : s = 246;
	{8'd210,8'd37} : s = 247;
	{8'd210,8'd38} : s = 248;
	{8'd210,8'd39} : s = 249;
	{8'd210,8'd40} : s = 250;
	{8'd210,8'd41} : s = 251;
	{8'd210,8'd42} : s = 252;
	{8'd210,8'd43} : s = 253;
	{8'd210,8'd44} : s = 254;
	{8'd210,8'd45} : s = 255;
	{8'd210,8'd46} : s = 256;
	{8'd210,8'd47} : s = 257;
	{8'd210,8'd48} : s = 258;
	{8'd210,8'd49} : s = 259;
	{8'd210,8'd50} : s = 260;
	{8'd210,8'd51} : s = 261;
	{8'd210,8'd52} : s = 262;
	{8'd210,8'd53} : s = 263;
	{8'd210,8'd54} : s = 264;
	{8'd210,8'd55} : s = 265;
	{8'd210,8'd56} : s = 266;
	{8'd210,8'd57} : s = 267;
	{8'd210,8'd58} : s = 268;
	{8'd210,8'd59} : s = 269;
	{8'd210,8'd60} : s = 270;
	{8'd210,8'd61} : s = 271;
	{8'd210,8'd62} : s = 272;
	{8'd210,8'd63} : s = 273;
	{8'd210,8'd64} : s = 274;
	{8'd210,8'd65} : s = 275;
	{8'd210,8'd66} : s = 276;
	{8'd210,8'd67} : s = 277;
	{8'd210,8'd68} : s = 278;
	{8'd210,8'd69} : s = 279;
	{8'd210,8'd70} : s = 280;
	{8'd210,8'd71} : s = 281;
	{8'd210,8'd72} : s = 282;
	{8'd210,8'd73} : s = 283;
	{8'd210,8'd74} : s = 284;
	{8'd210,8'd75} : s = 285;
	{8'd210,8'd76} : s = 286;
	{8'd210,8'd77} : s = 287;
	{8'd210,8'd78} : s = 288;
	{8'd210,8'd79} : s = 289;
	{8'd210,8'd80} : s = 290;
	{8'd210,8'd81} : s = 291;
	{8'd210,8'd82} : s = 292;
	{8'd210,8'd83} : s = 293;
	{8'd210,8'd84} : s = 294;
	{8'd210,8'd85} : s = 295;
	{8'd210,8'd86} : s = 296;
	{8'd210,8'd87} : s = 297;
	{8'd210,8'd88} : s = 298;
	{8'd210,8'd89} : s = 299;
	{8'd210,8'd90} : s = 300;
	{8'd210,8'd91} : s = 301;
	{8'd210,8'd92} : s = 302;
	{8'd210,8'd93} : s = 303;
	{8'd210,8'd94} : s = 304;
	{8'd210,8'd95} : s = 305;
	{8'd210,8'd96} : s = 306;
	{8'd210,8'd97} : s = 307;
	{8'd210,8'd98} : s = 308;
	{8'd210,8'd99} : s = 309;
	{8'd210,8'd100} : s = 310;
	{8'd210,8'd101} : s = 311;
	{8'd210,8'd102} : s = 312;
	{8'd210,8'd103} : s = 313;
	{8'd210,8'd104} : s = 314;
	{8'd210,8'd105} : s = 315;
	{8'd210,8'd106} : s = 316;
	{8'd210,8'd107} : s = 317;
	{8'd210,8'd108} : s = 318;
	{8'd210,8'd109} : s = 319;
	{8'd210,8'd110} : s = 320;
	{8'd210,8'd111} : s = 321;
	{8'd210,8'd112} : s = 322;
	{8'd210,8'd113} : s = 323;
	{8'd210,8'd114} : s = 324;
	{8'd210,8'd115} : s = 325;
	{8'd210,8'd116} : s = 326;
	{8'd210,8'd117} : s = 327;
	{8'd210,8'd118} : s = 328;
	{8'd210,8'd119} : s = 329;
	{8'd210,8'd120} : s = 330;
	{8'd210,8'd121} : s = 331;
	{8'd210,8'd122} : s = 332;
	{8'd210,8'd123} : s = 333;
	{8'd210,8'd124} : s = 334;
	{8'd210,8'd125} : s = 335;
	{8'd210,8'd126} : s = 336;
	{8'd210,8'd127} : s = 337;
	{8'd210,8'd128} : s = 338;
	{8'd210,8'd129} : s = 339;
	{8'd210,8'd130} : s = 340;
	{8'd210,8'd131} : s = 341;
	{8'd210,8'd132} : s = 342;
	{8'd210,8'd133} : s = 343;
	{8'd210,8'd134} : s = 344;
	{8'd210,8'd135} : s = 345;
	{8'd210,8'd136} : s = 346;
	{8'd210,8'd137} : s = 347;
	{8'd210,8'd138} : s = 348;
	{8'd210,8'd139} : s = 349;
	{8'd210,8'd140} : s = 350;
	{8'd210,8'd141} : s = 351;
	{8'd210,8'd142} : s = 352;
	{8'd210,8'd143} : s = 353;
	{8'd210,8'd144} : s = 354;
	{8'd210,8'd145} : s = 355;
	{8'd210,8'd146} : s = 356;
	{8'd210,8'd147} : s = 357;
	{8'd210,8'd148} : s = 358;
	{8'd210,8'd149} : s = 359;
	{8'd210,8'd150} : s = 360;
	{8'd210,8'd151} : s = 361;
	{8'd210,8'd152} : s = 362;
	{8'd210,8'd153} : s = 363;
	{8'd210,8'd154} : s = 364;
	{8'd210,8'd155} : s = 365;
	{8'd210,8'd156} : s = 366;
	{8'd210,8'd157} : s = 367;
	{8'd210,8'd158} : s = 368;
	{8'd210,8'd159} : s = 369;
	{8'd210,8'd160} : s = 370;
	{8'd210,8'd161} : s = 371;
	{8'd210,8'd162} : s = 372;
	{8'd210,8'd163} : s = 373;
	{8'd210,8'd164} : s = 374;
	{8'd210,8'd165} : s = 375;
	{8'd210,8'd166} : s = 376;
	{8'd210,8'd167} : s = 377;
	{8'd210,8'd168} : s = 378;
	{8'd210,8'd169} : s = 379;
	{8'd210,8'd170} : s = 380;
	{8'd210,8'd171} : s = 381;
	{8'd210,8'd172} : s = 382;
	{8'd210,8'd173} : s = 383;
	{8'd210,8'd174} : s = 384;
	{8'd210,8'd175} : s = 385;
	{8'd210,8'd176} : s = 386;
	{8'd210,8'd177} : s = 387;
	{8'd210,8'd178} : s = 388;
	{8'd210,8'd179} : s = 389;
	{8'd210,8'd180} : s = 390;
	{8'd210,8'd181} : s = 391;
	{8'd210,8'd182} : s = 392;
	{8'd210,8'd183} : s = 393;
	{8'd210,8'd184} : s = 394;
	{8'd210,8'd185} : s = 395;
	{8'd210,8'd186} : s = 396;
	{8'd210,8'd187} : s = 397;
	{8'd210,8'd188} : s = 398;
	{8'd210,8'd189} : s = 399;
	{8'd210,8'd190} : s = 400;
	{8'd210,8'd191} : s = 401;
	{8'd210,8'd192} : s = 402;
	{8'd210,8'd193} : s = 403;
	{8'd210,8'd194} : s = 404;
	{8'd210,8'd195} : s = 405;
	{8'd210,8'd196} : s = 406;
	{8'd210,8'd197} : s = 407;
	{8'd210,8'd198} : s = 408;
	{8'd210,8'd199} : s = 409;
	{8'd210,8'd200} : s = 410;
	{8'd210,8'd201} : s = 411;
	{8'd210,8'd202} : s = 412;
	{8'd210,8'd203} : s = 413;
	{8'd210,8'd204} : s = 414;
	{8'd210,8'd205} : s = 415;
	{8'd210,8'd206} : s = 416;
	{8'd210,8'd207} : s = 417;
	{8'd210,8'd208} : s = 418;
	{8'd210,8'd209} : s = 419;
	{8'd210,8'd210} : s = 420;
	{8'd210,8'd211} : s = 421;
	{8'd210,8'd212} : s = 422;
	{8'd210,8'd213} : s = 423;
	{8'd210,8'd214} : s = 424;
	{8'd210,8'd215} : s = 425;
	{8'd210,8'd216} : s = 426;
	{8'd210,8'd217} : s = 427;
	{8'd210,8'd218} : s = 428;
	{8'd210,8'd219} : s = 429;
	{8'd210,8'd220} : s = 430;
	{8'd210,8'd221} : s = 431;
	{8'd210,8'd222} : s = 432;
	{8'd210,8'd223} : s = 433;
	{8'd210,8'd224} : s = 434;
	{8'd210,8'd225} : s = 435;
	{8'd210,8'd226} : s = 436;
	{8'd210,8'd227} : s = 437;
	{8'd210,8'd228} : s = 438;
	{8'd210,8'd229} : s = 439;
	{8'd210,8'd230} : s = 440;
	{8'd210,8'd231} : s = 441;
	{8'd210,8'd232} : s = 442;
	{8'd210,8'd233} : s = 443;
	{8'd210,8'd234} : s = 444;
	{8'd210,8'd235} : s = 445;
	{8'd210,8'd236} : s = 446;
	{8'd210,8'd237} : s = 447;
	{8'd210,8'd238} : s = 448;
	{8'd210,8'd239} : s = 449;
	{8'd210,8'd240} : s = 450;
	{8'd210,8'd241} : s = 451;
	{8'd210,8'd242} : s = 452;
	{8'd210,8'd243} : s = 453;
	{8'd210,8'd244} : s = 454;
	{8'd210,8'd245} : s = 455;
	{8'd210,8'd246} : s = 456;
	{8'd210,8'd247} : s = 457;
	{8'd210,8'd248} : s = 458;
	{8'd210,8'd249} : s = 459;
	{8'd210,8'd250} : s = 460;
	{8'd210,8'd251} : s = 461;
	{8'd210,8'd252} : s = 462;
	{8'd210,8'd253} : s = 463;
	{8'd210,8'd254} : s = 464;
	{8'd210,8'd255} : s = 465;
	{8'd211,8'd0} : s = 211;
	{8'd211,8'd1} : s = 212;
	{8'd211,8'd2} : s = 213;
	{8'd211,8'd3} : s = 214;
	{8'd211,8'd4} : s = 215;
	{8'd211,8'd5} : s = 216;
	{8'd211,8'd6} : s = 217;
	{8'd211,8'd7} : s = 218;
	{8'd211,8'd8} : s = 219;
	{8'd211,8'd9} : s = 220;
	{8'd211,8'd10} : s = 221;
	{8'd211,8'd11} : s = 222;
	{8'd211,8'd12} : s = 223;
	{8'd211,8'd13} : s = 224;
	{8'd211,8'd14} : s = 225;
	{8'd211,8'd15} : s = 226;
	{8'd211,8'd16} : s = 227;
	{8'd211,8'd17} : s = 228;
	{8'd211,8'd18} : s = 229;
	{8'd211,8'd19} : s = 230;
	{8'd211,8'd20} : s = 231;
	{8'd211,8'd21} : s = 232;
	{8'd211,8'd22} : s = 233;
	{8'd211,8'd23} : s = 234;
	{8'd211,8'd24} : s = 235;
	{8'd211,8'd25} : s = 236;
	{8'd211,8'd26} : s = 237;
	{8'd211,8'd27} : s = 238;
	{8'd211,8'd28} : s = 239;
	{8'd211,8'd29} : s = 240;
	{8'd211,8'd30} : s = 241;
	{8'd211,8'd31} : s = 242;
	{8'd211,8'd32} : s = 243;
	{8'd211,8'd33} : s = 244;
	{8'd211,8'd34} : s = 245;
	{8'd211,8'd35} : s = 246;
	{8'd211,8'd36} : s = 247;
	{8'd211,8'd37} : s = 248;
	{8'd211,8'd38} : s = 249;
	{8'd211,8'd39} : s = 250;
	{8'd211,8'd40} : s = 251;
	{8'd211,8'd41} : s = 252;
	{8'd211,8'd42} : s = 253;
	{8'd211,8'd43} : s = 254;
	{8'd211,8'd44} : s = 255;
	{8'd211,8'd45} : s = 256;
	{8'd211,8'd46} : s = 257;
	{8'd211,8'd47} : s = 258;
	{8'd211,8'd48} : s = 259;
	{8'd211,8'd49} : s = 260;
	{8'd211,8'd50} : s = 261;
	{8'd211,8'd51} : s = 262;
	{8'd211,8'd52} : s = 263;
	{8'd211,8'd53} : s = 264;
	{8'd211,8'd54} : s = 265;
	{8'd211,8'd55} : s = 266;
	{8'd211,8'd56} : s = 267;
	{8'd211,8'd57} : s = 268;
	{8'd211,8'd58} : s = 269;
	{8'd211,8'd59} : s = 270;
	{8'd211,8'd60} : s = 271;
	{8'd211,8'd61} : s = 272;
	{8'd211,8'd62} : s = 273;
	{8'd211,8'd63} : s = 274;
	{8'd211,8'd64} : s = 275;
	{8'd211,8'd65} : s = 276;
	{8'd211,8'd66} : s = 277;
	{8'd211,8'd67} : s = 278;
	{8'd211,8'd68} : s = 279;
	{8'd211,8'd69} : s = 280;
	{8'd211,8'd70} : s = 281;
	{8'd211,8'd71} : s = 282;
	{8'd211,8'd72} : s = 283;
	{8'd211,8'd73} : s = 284;
	{8'd211,8'd74} : s = 285;
	{8'd211,8'd75} : s = 286;
	{8'd211,8'd76} : s = 287;
	{8'd211,8'd77} : s = 288;
	{8'd211,8'd78} : s = 289;
	{8'd211,8'd79} : s = 290;
	{8'd211,8'd80} : s = 291;
	{8'd211,8'd81} : s = 292;
	{8'd211,8'd82} : s = 293;
	{8'd211,8'd83} : s = 294;
	{8'd211,8'd84} : s = 295;
	{8'd211,8'd85} : s = 296;
	{8'd211,8'd86} : s = 297;
	{8'd211,8'd87} : s = 298;
	{8'd211,8'd88} : s = 299;
	{8'd211,8'd89} : s = 300;
	{8'd211,8'd90} : s = 301;
	{8'd211,8'd91} : s = 302;
	{8'd211,8'd92} : s = 303;
	{8'd211,8'd93} : s = 304;
	{8'd211,8'd94} : s = 305;
	{8'd211,8'd95} : s = 306;
	{8'd211,8'd96} : s = 307;
	{8'd211,8'd97} : s = 308;
	{8'd211,8'd98} : s = 309;
	{8'd211,8'd99} : s = 310;
	{8'd211,8'd100} : s = 311;
	{8'd211,8'd101} : s = 312;
	{8'd211,8'd102} : s = 313;
	{8'd211,8'd103} : s = 314;
	{8'd211,8'd104} : s = 315;
	{8'd211,8'd105} : s = 316;
	{8'd211,8'd106} : s = 317;
	{8'd211,8'd107} : s = 318;
	{8'd211,8'd108} : s = 319;
	{8'd211,8'd109} : s = 320;
	{8'd211,8'd110} : s = 321;
	{8'd211,8'd111} : s = 322;
	{8'd211,8'd112} : s = 323;
	{8'd211,8'd113} : s = 324;
	{8'd211,8'd114} : s = 325;
	{8'd211,8'd115} : s = 326;
	{8'd211,8'd116} : s = 327;
	{8'd211,8'd117} : s = 328;
	{8'd211,8'd118} : s = 329;
	{8'd211,8'd119} : s = 330;
	{8'd211,8'd120} : s = 331;
	{8'd211,8'd121} : s = 332;
	{8'd211,8'd122} : s = 333;
	{8'd211,8'd123} : s = 334;
	{8'd211,8'd124} : s = 335;
	{8'd211,8'd125} : s = 336;
	{8'd211,8'd126} : s = 337;
	{8'd211,8'd127} : s = 338;
	{8'd211,8'd128} : s = 339;
	{8'd211,8'd129} : s = 340;
	{8'd211,8'd130} : s = 341;
	{8'd211,8'd131} : s = 342;
	{8'd211,8'd132} : s = 343;
	{8'd211,8'd133} : s = 344;
	{8'd211,8'd134} : s = 345;
	{8'd211,8'd135} : s = 346;
	{8'd211,8'd136} : s = 347;
	{8'd211,8'd137} : s = 348;
	{8'd211,8'd138} : s = 349;
	{8'd211,8'd139} : s = 350;
	{8'd211,8'd140} : s = 351;
	{8'd211,8'd141} : s = 352;
	{8'd211,8'd142} : s = 353;
	{8'd211,8'd143} : s = 354;
	{8'd211,8'd144} : s = 355;
	{8'd211,8'd145} : s = 356;
	{8'd211,8'd146} : s = 357;
	{8'd211,8'd147} : s = 358;
	{8'd211,8'd148} : s = 359;
	{8'd211,8'd149} : s = 360;
	{8'd211,8'd150} : s = 361;
	{8'd211,8'd151} : s = 362;
	{8'd211,8'd152} : s = 363;
	{8'd211,8'd153} : s = 364;
	{8'd211,8'd154} : s = 365;
	{8'd211,8'd155} : s = 366;
	{8'd211,8'd156} : s = 367;
	{8'd211,8'd157} : s = 368;
	{8'd211,8'd158} : s = 369;
	{8'd211,8'd159} : s = 370;
	{8'd211,8'd160} : s = 371;
	{8'd211,8'd161} : s = 372;
	{8'd211,8'd162} : s = 373;
	{8'd211,8'd163} : s = 374;
	{8'd211,8'd164} : s = 375;
	{8'd211,8'd165} : s = 376;
	{8'd211,8'd166} : s = 377;
	{8'd211,8'd167} : s = 378;
	{8'd211,8'd168} : s = 379;
	{8'd211,8'd169} : s = 380;
	{8'd211,8'd170} : s = 381;
	{8'd211,8'd171} : s = 382;
	{8'd211,8'd172} : s = 383;
	{8'd211,8'd173} : s = 384;
	{8'd211,8'd174} : s = 385;
	{8'd211,8'd175} : s = 386;
	{8'd211,8'd176} : s = 387;
	{8'd211,8'd177} : s = 388;
	{8'd211,8'd178} : s = 389;
	{8'd211,8'd179} : s = 390;
	{8'd211,8'd180} : s = 391;
	{8'd211,8'd181} : s = 392;
	{8'd211,8'd182} : s = 393;
	{8'd211,8'd183} : s = 394;
	{8'd211,8'd184} : s = 395;
	{8'd211,8'd185} : s = 396;
	{8'd211,8'd186} : s = 397;
	{8'd211,8'd187} : s = 398;
	{8'd211,8'd188} : s = 399;
	{8'd211,8'd189} : s = 400;
	{8'd211,8'd190} : s = 401;
	{8'd211,8'd191} : s = 402;
	{8'd211,8'd192} : s = 403;
	{8'd211,8'd193} : s = 404;
	{8'd211,8'd194} : s = 405;
	{8'd211,8'd195} : s = 406;
	{8'd211,8'd196} : s = 407;
	{8'd211,8'd197} : s = 408;
	{8'd211,8'd198} : s = 409;
	{8'd211,8'd199} : s = 410;
	{8'd211,8'd200} : s = 411;
	{8'd211,8'd201} : s = 412;
	{8'd211,8'd202} : s = 413;
	{8'd211,8'd203} : s = 414;
	{8'd211,8'd204} : s = 415;
	{8'd211,8'd205} : s = 416;
	{8'd211,8'd206} : s = 417;
	{8'd211,8'd207} : s = 418;
	{8'd211,8'd208} : s = 419;
	{8'd211,8'd209} : s = 420;
	{8'd211,8'd210} : s = 421;
	{8'd211,8'd211} : s = 422;
	{8'd211,8'd212} : s = 423;
	{8'd211,8'd213} : s = 424;
	{8'd211,8'd214} : s = 425;
	{8'd211,8'd215} : s = 426;
	{8'd211,8'd216} : s = 427;
	{8'd211,8'd217} : s = 428;
	{8'd211,8'd218} : s = 429;
	{8'd211,8'd219} : s = 430;
	{8'd211,8'd220} : s = 431;
	{8'd211,8'd221} : s = 432;
	{8'd211,8'd222} : s = 433;
	{8'd211,8'd223} : s = 434;
	{8'd211,8'd224} : s = 435;
	{8'd211,8'd225} : s = 436;
	{8'd211,8'd226} : s = 437;
	{8'd211,8'd227} : s = 438;
	{8'd211,8'd228} : s = 439;
	{8'd211,8'd229} : s = 440;
	{8'd211,8'd230} : s = 441;
	{8'd211,8'd231} : s = 442;
	{8'd211,8'd232} : s = 443;
	{8'd211,8'd233} : s = 444;
	{8'd211,8'd234} : s = 445;
	{8'd211,8'd235} : s = 446;
	{8'd211,8'd236} : s = 447;
	{8'd211,8'd237} : s = 448;
	{8'd211,8'd238} : s = 449;
	{8'd211,8'd239} : s = 450;
	{8'd211,8'd240} : s = 451;
	{8'd211,8'd241} : s = 452;
	{8'd211,8'd242} : s = 453;
	{8'd211,8'd243} : s = 454;
	{8'd211,8'd244} : s = 455;
	{8'd211,8'd245} : s = 456;
	{8'd211,8'd246} : s = 457;
	{8'd211,8'd247} : s = 458;
	{8'd211,8'd248} : s = 459;
	{8'd211,8'd249} : s = 460;
	{8'd211,8'd250} : s = 461;
	{8'd211,8'd251} : s = 462;
	{8'd211,8'd252} : s = 463;
	{8'd211,8'd253} : s = 464;
	{8'd211,8'd254} : s = 465;
	{8'd211,8'd255} : s = 466;
	{8'd212,8'd0} : s = 212;
	{8'd212,8'd1} : s = 213;
	{8'd212,8'd2} : s = 214;
	{8'd212,8'd3} : s = 215;
	{8'd212,8'd4} : s = 216;
	{8'd212,8'd5} : s = 217;
	{8'd212,8'd6} : s = 218;
	{8'd212,8'd7} : s = 219;
	{8'd212,8'd8} : s = 220;
	{8'd212,8'd9} : s = 221;
	{8'd212,8'd10} : s = 222;
	{8'd212,8'd11} : s = 223;
	{8'd212,8'd12} : s = 224;
	{8'd212,8'd13} : s = 225;
	{8'd212,8'd14} : s = 226;
	{8'd212,8'd15} : s = 227;
	{8'd212,8'd16} : s = 228;
	{8'd212,8'd17} : s = 229;
	{8'd212,8'd18} : s = 230;
	{8'd212,8'd19} : s = 231;
	{8'd212,8'd20} : s = 232;
	{8'd212,8'd21} : s = 233;
	{8'd212,8'd22} : s = 234;
	{8'd212,8'd23} : s = 235;
	{8'd212,8'd24} : s = 236;
	{8'd212,8'd25} : s = 237;
	{8'd212,8'd26} : s = 238;
	{8'd212,8'd27} : s = 239;
	{8'd212,8'd28} : s = 240;
	{8'd212,8'd29} : s = 241;
	{8'd212,8'd30} : s = 242;
	{8'd212,8'd31} : s = 243;
	{8'd212,8'd32} : s = 244;
	{8'd212,8'd33} : s = 245;
	{8'd212,8'd34} : s = 246;
	{8'd212,8'd35} : s = 247;
	{8'd212,8'd36} : s = 248;
	{8'd212,8'd37} : s = 249;
	{8'd212,8'd38} : s = 250;
	{8'd212,8'd39} : s = 251;
	{8'd212,8'd40} : s = 252;
	{8'd212,8'd41} : s = 253;
	{8'd212,8'd42} : s = 254;
	{8'd212,8'd43} : s = 255;
	{8'd212,8'd44} : s = 256;
	{8'd212,8'd45} : s = 257;
	{8'd212,8'd46} : s = 258;
	{8'd212,8'd47} : s = 259;
	{8'd212,8'd48} : s = 260;
	{8'd212,8'd49} : s = 261;
	{8'd212,8'd50} : s = 262;
	{8'd212,8'd51} : s = 263;
	{8'd212,8'd52} : s = 264;
	{8'd212,8'd53} : s = 265;
	{8'd212,8'd54} : s = 266;
	{8'd212,8'd55} : s = 267;
	{8'd212,8'd56} : s = 268;
	{8'd212,8'd57} : s = 269;
	{8'd212,8'd58} : s = 270;
	{8'd212,8'd59} : s = 271;
	{8'd212,8'd60} : s = 272;
	{8'd212,8'd61} : s = 273;
	{8'd212,8'd62} : s = 274;
	{8'd212,8'd63} : s = 275;
	{8'd212,8'd64} : s = 276;
	{8'd212,8'd65} : s = 277;
	{8'd212,8'd66} : s = 278;
	{8'd212,8'd67} : s = 279;
	{8'd212,8'd68} : s = 280;
	{8'd212,8'd69} : s = 281;
	{8'd212,8'd70} : s = 282;
	{8'd212,8'd71} : s = 283;
	{8'd212,8'd72} : s = 284;
	{8'd212,8'd73} : s = 285;
	{8'd212,8'd74} : s = 286;
	{8'd212,8'd75} : s = 287;
	{8'd212,8'd76} : s = 288;
	{8'd212,8'd77} : s = 289;
	{8'd212,8'd78} : s = 290;
	{8'd212,8'd79} : s = 291;
	{8'd212,8'd80} : s = 292;
	{8'd212,8'd81} : s = 293;
	{8'd212,8'd82} : s = 294;
	{8'd212,8'd83} : s = 295;
	{8'd212,8'd84} : s = 296;
	{8'd212,8'd85} : s = 297;
	{8'd212,8'd86} : s = 298;
	{8'd212,8'd87} : s = 299;
	{8'd212,8'd88} : s = 300;
	{8'd212,8'd89} : s = 301;
	{8'd212,8'd90} : s = 302;
	{8'd212,8'd91} : s = 303;
	{8'd212,8'd92} : s = 304;
	{8'd212,8'd93} : s = 305;
	{8'd212,8'd94} : s = 306;
	{8'd212,8'd95} : s = 307;
	{8'd212,8'd96} : s = 308;
	{8'd212,8'd97} : s = 309;
	{8'd212,8'd98} : s = 310;
	{8'd212,8'd99} : s = 311;
	{8'd212,8'd100} : s = 312;
	{8'd212,8'd101} : s = 313;
	{8'd212,8'd102} : s = 314;
	{8'd212,8'd103} : s = 315;
	{8'd212,8'd104} : s = 316;
	{8'd212,8'd105} : s = 317;
	{8'd212,8'd106} : s = 318;
	{8'd212,8'd107} : s = 319;
	{8'd212,8'd108} : s = 320;
	{8'd212,8'd109} : s = 321;
	{8'd212,8'd110} : s = 322;
	{8'd212,8'd111} : s = 323;
	{8'd212,8'd112} : s = 324;
	{8'd212,8'd113} : s = 325;
	{8'd212,8'd114} : s = 326;
	{8'd212,8'd115} : s = 327;
	{8'd212,8'd116} : s = 328;
	{8'd212,8'd117} : s = 329;
	{8'd212,8'd118} : s = 330;
	{8'd212,8'd119} : s = 331;
	{8'd212,8'd120} : s = 332;
	{8'd212,8'd121} : s = 333;
	{8'd212,8'd122} : s = 334;
	{8'd212,8'd123} : s = 335;
	{8'd212,8'd124} : s = 336;
	{8'd212,8'd125} : s = 337;
	{8'd212,8'd126} : s = 338;
	{8'd212,8'd127} : s = 339;
	{8'd212,8'd128} : s = 340;
	{8'd212,8'd129} : s = 341;
	{8'd212,8'd130} : s = 342;
	{8'd212,8'd131} : s = 343;
	{8'd212,8'd132} : s = 344;
	{8'd212,8'd133} : s = 345;
	{8'd212,8'd134} : s = 346;
	{8'd212,8'd135} : s = 347;
	{8'd212,8'd136} : s = 348;
	{8'd212,8'd137} : s = 349;
	{8'd212,8'd138} : s = 350;
	{8'd212,8'd139} : s = 351;
	{8'd212,8'd140} : s = 352;
	{8'd212,8'd141} : s = 353;
	{8'd212,8'd142} : s = 354;
	{8'd212,8'd143} : s = 355;
	{8'd212,8'd144} : s = 356;
	{8'd212,8'd145} : s = 357;
	{8'd212,8'd146} : s = 358;
	{8'd212,8'd147} : s = 359;
	{8'd212,8'd148} : s = 360;
	{8'd212,8'd149} : s = 361;
	{8'd212,8'd150} : s = 362;
	{8'd212,8'd151} : s = 363;
	{8'd212,8'd152} : s = 364;
	{8'd212,8'd153} : s = 365;
	{8'd212,8'd154} : s = 366;
	{8'd212,8'd155} : s = 367;
	{8'd212,8'd156} : s = 368;
	{8'd212,8'd157} : s = 369;
	{8'd212,8'd158} : s = 370;
	{8'd212,8'd159} : s = 371;
	{8'd212,8'd160} : s = 372;
	{8'd212,8'd161} : s = 373;
	{8'd212,8'd162} : s = 374;
	{8'd212,8'd163} : s = 375;
	{8'd212,8'd164} : s = 376;
	{8'd212,8'd165} : s = 377;
	{8'd212,8'd166} : s = 378;
	{8'd212,8'd167} : s = 379;
	{8'd212,8'd168} : s = 380;
	{8'd212,8'd169} : s = 381;
	{8'd212,8'd170} : s = 382;
	{8'd212,8'd171} : s = 383;
	{8'd212,8'd172} : s = 384;
	{8'd212,8'd173} : s = 385;
	{8'd212,8'd174} : s = 386;
	{8'd212,8'd175} : s = 387;
	{8'd212,8'd176} : s = 388;
	{8'd212,8'd177} : s = 389;
	{8'd212,8'd178} : s = 390;
	{8'd212,8'd179} : s = 391;
	{8'd212,8'd180} : s = 392;
	{8'd212,8'd181} : s = 393;
	{8'd212,8'd182} : s = 394;
	{8'd212,8'd183} : s = 395;
	{8'd212,8'd184} : s = 396;
	{8'd212,8'd185} : s = 397;
	{8'd212,8'd186} : s = 398;
	{8'd212,8'd187} : s = 399;
	{8'd212,8'd188} : s = 400;
	{8'd212,8'd189} : s = 401;
	{8'd212,8'd190} : s = 402;
	{8'd212,8'd191} : s = 403;
	{8'd212,8'd192} : s = 404;
	{8'd212,8'd193} : s = 405;
	{8'd212,8'd194} : s = 406;
	{8'd212,8'd195} : s = 407;
	{8'd212,8'd196} : s = 408;
	{8'd212,8'd197} : s = 409;
	{8'd212,8'd198} : s = 410;
	{8'd212,8'd199} : s = 411;
	{8'd212,8'd200} : s = 412;
	{8'd212,8'd201} : s = 413;
	{8'd212,8'd202} : s = 414;
	{8'd212,8'd203} : s = 415;
	{8'd212,8'd204} : s = 416;
	{8'd212,8'd205} : s = 417;
	{8'd212,8'd206} : s = 418;
	{8'd212,8'd207} : s = 419;
	{8'd212,8'd208} : s = 420;
	{8'd212,8'd209} : s = 421;
	{8'd212,8'd210} : s = 422;
	{8'd212,8'd211} : s = 423;
	{8'd212,8'd212} : s = 424;
	{8'd212,8'd213} : s = 425;
	{8'd212,8'd214} : s = 426;
	{8'd212,8'd215} : s = 427;
	{8'd212,8'd216} : s = 428;
	{8'd212,8'd217} : s = 429;
	{8'd212,8'd218} : s = 430;
	{8'd212,8'd219} : s = 431;
	{8'd212,8'd220} : s = 432;
	{8'd212,8'd221} : s = 433;
	{8'd212,8'd222} : s = 434;
	{8'd212,8'd223} : s = 435;
	{8'd212,8'd224} : s = 436;
	{8'd212,8'd225} : s = 437;
	{8'd212,8'd226} : s = 438;
	{8'd212,8'd227} : s = 439;
	{8'd212,8'd228} : s = 440;
	{8'd212,8'd229} : s = 441;
	{8'd212,8'd230} : s = 442;
	{8'd212,8'd231} : s = 443;
	{8'd212,8'd232} : s = 444;
	{8'd212,8'd233} : s = 445;
	{8'd212,8'd234} : s = 446;
	{8'd212,8'd235} : s = 447;
	{8'd212,8'd236} : s = 448;
	{8'd212,8'd237} : s = 449;
	{8'd212,8'd238} : s = 450;
	{8'd212,8'd239} : s = 451;
	{8'd212,8'd240} : s = 452;
	{8'd212,8'd241} : s = 453;
	{8'd212,8'd242} : s = 454;
	{8'd212,8'd243} : s = 455;
	{8'd212,8'd244} : s = 456;
	{8'd212,8'd245} : s = 457;
	{8'd212,8'd246} : s = 458;
	{8'd212,8'd247} : s = 459;
	{8'd212,8'd248} : s = 460;
	{8'd212,8'd249} : s = 461;
	{8'd212,8'd250} : s = 462;
	{8'd212,8'd251} : s = 463;
	{8'd212,8'd252} : s = 464;
	{8'd212,8'd253} : s = 465;
	{8'd212,8'd254} : s = 466;
	{8'd212,8'd255} : s = 467;
	{8'd213,8'd0} : s = 213;
	{8'd213,8'd1} : s = 214;
	{8'd213,8'd2} : s = 215;
	{8'd213,8'd3} : s = 216;
	{8'd213,8'd4} : s = 217;
	{8'd213,8'd5} : s = 218;
	{8'd213,8'd6} : s = 219;
	{8'd213,8'd7} : s = 220;
	{8'd213,8'd8} : s = 221;
	{8'd213,8'd9} : s = 222;
	{8'd213,8'd10} : s = 223;
	{8'd213,8'd11} : s = 224;
	{8'd213,8'd12} : s = 225;
	{8'd213,8'd13} : s = 226;
	{8'd213,8'd14} : s = 227;
	{8'd213,8'd15} : s = 228;
	{8'd213,8'd16} : s = 229;
	{8'd213,8'd17} : s = 230;
	{8'd213,8'd18} : s = 231;
	{8'd213,8'd19} : s = 232;
	{8'd213,8'd20} : s = 233;
	{8'd213,8'd21} : s = 234;
	{8'd213,8'd22} : s = 235;
	{8'd213,8'd23} : s = 236;
	{8'd213,8'd24} : s = 237;
	{8'd213,8'd25} : s = 238;
	{8'd213,8'd26} : s = 239;
	{8'd213,8'd27} : s = 240;
	{8'd213,8'd28} : s = 241;
	{8'd213,8'd29} : s = 242;
	{8'd213,8'd30} : s = 243;
	{8'd213,8'd31} : s = 244;
	{8'd213,8'd32} : s = 245;
	{8'd213,8'd33} : s = 246;
	{8'd213,8'd34} : s = 247;
	{8'd213,8'd35} : s = 248;
	{8'd213,8'd36} : s = 249;
	{8'd213,8'd37} : s = 250;
	{8'd213,8'd38} : s = 251;
	{8'd213,8'd39} : s = 252;
	{8'd213,8'd40} : s = 253;
	{8'd213,8'd41} : s = 254;
	{8'd213,8'd42} : s = 255;
	{8'd213,8'd43} : s = 256;
	{8'd213,8'd44} : s = 257;
	{8'd213,8'd45} : s = 258;
	{8'd213,8'd46} : s = 259;
	{8'd213,8'd47} : s = 260;
	{8'd213,8'd48} : s = 261;
	{8'd213,8'd49} : s = 262;
	{8'd213,8'd50} : s = 263;
	{8'd213,8'd51} : s = 264;
	{8'd213,8'd52} : s = 265;
	{8'd213,8'd53} : s = 266;
	{8'd213,8'd54} : s = 267;
	{8'd213,8'd55} : s = 268;
	{8'd213,8'd56} : s = 269;
	{8'd213,8'd57} : s = 270;
	{8'd213,8'd58} : s = 271;
	{8'd213,8'd59} : s = 272;
	{8'd213,8'd60} : s = 273;
	{8'd213,8'd61} : s = 274;
	{8'd213,8'd62} : s = 275;
	{8'd213,8'd63} : s = 276;
	{8'd213,8'd64} : s = 277;
	{8'd213,8'd65} : s = 278;
	{8'd213,8'd66} : s = 279;
	{8'd213,8'd67} : s = 280;
	{8'd213,8'd68} : s = 281;
	{8'd213,8'd69} : s = 282;
	{8'd213,8'd70} : s = 283;
	{8'd213,8'd71} : s = 284;
	{8'd213,8'd72} : s = 285;
	{8'd213,8'd73} : s = 286;
	{8'd213,8'd74} : s = 287;
	{8'd213,8'd75} : s = 288;
	{8'd213,8'd76} : s = 289;
	{8'd213,8'd77} : s = 290;
	{8'd213,8'd78} : s = 291;
	{8'd213,8'd79} : s = 292;
	{8'd213,8'd80} : s = 293;
	{8'd213,8'd81} : s = 294;
	{8'd213,8'd82} : s = 295;
	{8'd213,8'd83} : s = 296;
	{8'd213,8'd84} : s = 297;
	{8'd213,8'd85} : s = 298;
	{8'd213,8'd86} : s = 299;
	{8'd213,8'd87} : s = 300;
	{8'd213,8'd88} : s = 301;
	{8'd213,8'd89} : s = 302;
	{8'd213,8'd90} : s = 303;
	{8'd213,8'd91} : s = 304;
	{8'd213,8'd92} : s = 305;
	{8'd213,8'd93} : s = 306;
	{8'd213,8'd94} : s = 307;
	{8'd213,8'd95} : s = 308;
	{8'd213,8'd96} : s = 309;
	{8'd213,8'd97} : s = 310;
	{8'd213,8'd98} : s = 311;
	{8'd213,8'd99} : s = 312;
	{8'd213,8'd100} : s = 313;
	{8'd213,8'd101} : s = 314;
	{8'd213,8'd102} : s = 315;
	{8'd213,8'd103} : s = 316;
	{8'd213,8'd104} : s = 317;
	{8'd213,8'd105} : s = 318;
	{8'd213,8'd106} : s = 319;
	{8'd213,8'd107} : s = 320;
	{8'd213,8'd108} : s = 321;
	{8'd213,8'd109} : s = 322;
	{8'd213,8'd110} : s = 323;
	{8'd213,8'd111} : s = 324;
	{8'd213,8'd112} : s = 325;
	{8'd213,8'd113} : s = 326;
	{8'd213,8'd114} : s = 327;
	{8'd213,8'd115} : s = 328;
	{8'd213,8'd116} : s = 329;
	{8'd213,8'd117} : s = 330;
	{8'd213,8'd118} : s = 331;
	{8'd213,8'd119} : s = 332;
	{8'd213,8'd120} : s = 333;
	{8'd213,8'd121} : s = 334;
	{8'd213,8'd122} : s = 335;
	{8'd213,8'd123} : s = 336;
	{8'd213,8'd124} : s = 337;
	{8'd213,8'd125} : s = 338;
	{8'd213,8'd126} : s = 339;
	{8'd213,8'd127} : s = 340;
	{8'd213,8'd128} : s = 341;
	{8'd213,8'd129} : s = 342;
	{8'd213,8'd130} : s = 343;
	{8'd213,8'd131} : s = 344;
	{8'd213,8'd132} : s = 345;
	{8'd213,8'd133} : s = 346;
	{8'd213,8'd134} : s = 347;
	{8'd213,8'd135} : s = 348;
	{8'd213,8'd136} : s = 349;
	{8'd213,8'd137} : s = 350;
	{8'd213,8'd138} : s = 351;
	{8'd213,8'd139} : s = 352;
	{8'd213,8'd140} : s = 353;
	{8'd213,8'd141} : s = 354;
	{8'd213,8'd142} : s = 355;
	{8'd213,8'd143} : s = 356;
	{8'd213,8'd144} : s = 357;
	{8'd213,8'd145} : s = 358;
	{8'd213,8'd146} : s = 359;
	{8'd213,8'd147} : s = 360;
	{8'd213,8'd148} : s = 361;
	{8'd213,8'd149} : s = 362;
	{8'd213,8'd150} : s = 363;
	{8'd213,8'd151} : s = 364;
	{8'd213,8'd152} : s = 365;
	{8'd213,8'd153} : s = 366;
	{8'd213,8'd154} : s = 367;
	{8'd213,8'd155} : s = 368;
	{8'd213,8'd156} : s = 369;
	{8'd213,8'd157} : s = 370;
	{8'd213,8'd158} : s = 371;
	{8'd213,8'd159} : s = 372;
	{8'd213,8'd160} : s = 373;
	{8'd213,8'd161} : s = 374;
	{8'd213,8'd162} : s = 375;
	{8'd213,8'd163} : s = 376;
	{8'd213,8'd164} : s = 377;
	{8'd213,8'd165} : s = 378;
	{8'd213,8'd166} : s = 379;
	{8'd213,8'd167} : s = 380;
	{8'd213,8'd168} : s = 381;
	{8'd213,8'd169} : s = 382;
	{8'd213,8'd170} : s = 383;
	{8'd213,8'd171} : s = 384;
	{8'd213,8'd172} : s = 385;
	{8'd213,8'd173} : s = 386;
	{8'd213,8'd174} : s = 387;
	{8'd213,8'd175} : s = 388;
	{8'd213,8'd176} : s = 389;
	{8'd213,8'd177} : s = 390;
	{8'd213,8'd178} : s = 391;
	{8'd213,8'd179} : s = 392;
	{8'd213,8'd180} : s = 393;
	{8'd213,8'd181} : s = 394;
	{8'd213,8'd182} : s = 395;
	{8'd213,8'd183} : s = 396;
	{8'd213,8'd184} : s = 397;
	{8'd213,8'd185} : s = 398;
	{8'd213,8'd186} : s = 399;
	{8'd213,8'd187} : s = 400;
	{8'd213,8'd188} : s = 401;
	{8'd213,8'd189} : s = 402;
	{8'd213,8'd190} : s = 403;
	{8'd213,8'd191} : s = 404;
	{8'd213,8'd192} : s = 405;
	{8'd213,8'd193} : s = 406;
	{8'd213,8'd194} : s = 407;
	{8'd213,8'd195} : s = 408;
	{8'd213,8'd196} : s = 409;
	{8'd213,8'd197} : s = 410;
	{8'd213,8'd198} : s = 411;
	{8'd213,8'd199} : s = 412;
	{8'd213,8'd200} : s = 413;
	{8'd213,8'd201} : s = 414;
	{8'd213,8'd202} : s = 415;
	{8'd213,8'd203} : s = 416;
	{8'd213,8'd204} : s = 417;
	{8'd213,8'd205} : s = 418;
	{8'd213,8'd206} : s = 419;
	{8'd213,8'd207} : s = 420;
	{8'd213,8'd208} : s = 421;
	{8'd213,8'd209} : s = 422;
	{8'd213,8'd210} : s = 423;
	{8'd213,8'd211} : s = 424;
	{8'd213,8'd212} : s = 425;
	{8'd213,8'd213} : s = 426;
	{8'd213,8'd214} : s = 427;
	{8'd213,8'd215} : s = 428;
	{8'd213,8'd216} : s = 429;
	{8'd213,8'd217} : s = 430;
	{8'd213,8'd218} : s = 431;
	{8'd213,8'd219} : s = 432;
	{8'd213,8'd220} : s = 433;
	{8'd213,8'd221} : s = 434;
	{8'd213,8'd222} : s = 435;
	{8'd213,8'd223} : s = 436;
	{8'd213,8'd224} : s = 437;
	{8'd213,8'd225} : s = 438;
	{8'd213,8'd226} : s = 439;
	{8'd213,8'd227} : s = 440;
	{8'd213,8'd228} : s = 441;
	{8'd213,8'd229} : s = 442;
	{8'd213,8'd230} : s = 443;
	{8'd213,8'd231} : s = 444;
	{8'd213,8'd232} : s = 445;
	{8'd213,8'd233} : s = 446;
	{8'd213,8'd234} : s = 447;
	{8'd213,8'd235} : s = 448;
	{8'd213,8'd236} : s = 449;
	{8'd213,8'd237} : s = 450;
	{8'd213,8'd238} : s = 451;
	{8'd213,8'd239} : s = 452;
	{8'd213,8'd240} : s = 453;
	{8'd213,8'd241} : s = 454;
	{8'd213,8'd242} : s = 455;
	{8'd213,8'd243} : s = 456;
	{8'd213,8'd244} : s = 457;
	{8'd213,8'd245} : s = 458;
	{8'd213,8'd246} : s = 459;
	{8'd213,8'd247} : s = 460;
	{8'd213,8'd248} : s = 461;
	{8'd213,8'd249} : s = 462;
	{8'd213,8'd250} : s = 463;
	{8'd213,8'd251} : s = 464;
	{8'd213,8'd252} : s = 465;
	{8'd213,8'd253} : s = 466;
	{8'd213,8'd254} : s = 467;
	{8'd213,8'd255} : s = 468;
	{8'd214,8'd0} : s = 214;
	{8'd214,8'd1} : s = 215;
	{8'd214,8'd2} : s = 216;
	{8'd214,8'd3} : s = 217;
	{8'd214,8'd4} : s = 218;
	{8'd214,8'd5} : s = 219;
	{8'd214,8'd6} : s = 220;
	{8'd214,8'd7} : s = 221;
	{8'd214,8'd8} : s = 222;
	{8'd214,8'd9} : s = 223;
	{8'd214,8'd10} : s = 224;
	{8'd214,8'd11} : s = 225;
	{8'd214,8'd12} : s = 226;
	{8'd214,8'd13} : s = 227;
	{8'd214,8'd14} : s = 228;
	{8'd214,8'd15} : s = 229;
	{8'd214,8'd16} : s = 230;
	{8'd214,8'd17} : s = 231;
	{8'd214,8'd18} : s = 232;
	{8'd214,8'd19} : s = 233;
	{8'd214,8'd20} : s = 234;
	{8'd214,8'd21} : s = 235;
	{8'd214,8'd22} : s = 236;
	{8'd214,8'd23} : s = 237;
	{8'd214,8'd24} : s = 238;
	{8'd214,8'd25} : s = 239;
	{8'd214,8'd26} : s = 240;
	{8'd214,8'd27} : s = 241;
	{8'd214,8'd28} : s = 242;
	{8'd214,8'd29} : s = 243;
	{8'd214,8'd30} : s = 244;
	{8'd214,8'd31} : s = 245;
	{8'd214,8'd32} : s = 246;
	{8'd214,8'd33} : s = 247;
	{8'd214,8'd34} : s = 248;
	{8'd214,8'd35} : s = 249;
	{8'd214,8'd36} : s = 250;
	{8'd214,8'd37} : s = 251;
	{8'd214,8'd38} : s = 252;
	{8'd214,8'd39} : s = 253;
	{8'd214,8'd40} : s = 254;
	{8'd214,8'd41} : s = 255;
	{8'd214,8'd42} : s = 256;
	{8'd214,8'd43} : s = 257;
	{8'd214,8'd44} : s = 258;
	{8'd214,8'd45} : s = 259;
	{8'd214,8'd46} : s = 260;
	{8'd214,8'd47} : s = 261;
	{8'd214,8'd48} : s = 262;
	{8'd214,8'd49} : s = 263;
	{8'd214,8'd50} : s = 264;
	{8'd214,8'd51} : s = 265;
	{8'd214,8'd52} : s = 266;
	{8'd214,8'd53} : s = 267;
	{8'd214,8'd54} : s = 268;
	{8'd214,8'd55} : s = 269;
	{8'd214,8'd56} : s = 270;
	{8'd214,8'd57} : s = 271;
	{8'd214,8'd58} : s = 272;
	{8'd214,8'd59} : s = 273;
	{8'd214,8'd60} : s = 274;
	{8'd214,8'd61} : s = 275;
	{8'd214,8'd62} : s = 276;
	{8'd214,8'd63} : s = 277;
	{8'd214,8'd64} : s = 278;
	{8'd214,8'd65} : s = 279;
	{8'd214,8'd66} : s = 280;
	{8'd214,8'd67} : s = 281;
	{8'd214,8'd68} : s = 282;
	{8'd214,8'd69} : s = 283;
	{8'd214,8'd70} : s = 284;
	{8'd214,8'd71} : s = 285;
	{8'd214,8'd72} : s = 286;
	{8'd214,8'd73} : s = 287;
	{8'd214,8'd74} : s = 288;
	{8'd214,8'd75} : s = 289;
	{8'd214,8'd76} : s = 290;
	{8'd214,8'd77} : s = 291;
	{8'd214,8'd78} : s = 292;
	{8'd214,8'd79} : s = 293;
	{8'd214,8'd80} : s = 294;
	{8'd214,8'd81} : s = 295;
	{8'd214,8'd82} : s = 296;
	{8'd214,8'd83} : s = 297;
	{8'd214,8'd84} : s = 298;
	{8'd214,8'd85} : s = 299;
	{8'd214,8'd86} : s = 300;
	{8'd214,8'd87} : s = 301;
	{8'd214,8'd88} : s = 302;
	{8'd214,8'd89} : s = 303;
	{8'd214,8'd90} : s = 304;
	{8'd214,8'd91} : s = 305;
	{8'd214,8'd92} : s = 306;
	{8'd214,8'd93} : s = 307;
	{8'd214,8'd94} : s = 308;
	{8'd214,8'd95} : s = 309;
	{8'd214,8'd96} : s = 310;
	{8'd214,8'd97} : s = 311;
	{8'd214,8'd98} : s = 312;
	{8'd214,8'd99} : s = 313;
	{8'd214,8'd100} : s = 314;
	{8'd214,8'd101} : s = 315;
	{8'd214,8'd102} : s = 316;
	{8'd214,8'd103} : s = 317;
	{8'd214,8'd104} : s = 318;
	{8'd214,8'd105} : s = 319;
	{8'd214,8'd106} : s = 320;
	{8'd214,8'd107} : s = 321;
	{8'd214,8'd108} : s = 322;
	{8'd214,8'd109} : s = 323;
	{8'd214,8'd110} : s = 324;
	{8'd214,8'd111} : s = 325;
	{8'd214,8'd112} : s = 326;
	{8'd214,8'd113} : s = 327;
	{8'd214,8'd114} : s = 328;
	{8'd214,8'd115} : s = 329;
	{8'd214,8'd116} : s = 330;
	{8'd214,8'd117} : s = 331;
	{8'd214,8'd118} : s = 332;
	{8'd214,8'd119} : s = 333;
	{8'd214,8'd120} : s = 334;
	{8'd214,8'd121} : s = 335;
	{8'd214,8'd122} : s = 336;
	{8'd214,8'd123} : s = 337;
	{8'd214,8'd124} : s = 338;
	{8'd214,8'd125} : s = 339;
	{8'd214,8'd126} : s = 340;
	{8'd214,8'd127} : s = 341;
	{8'd214,8'd128} : s = 342;
	{8'd214,8'd129} : s = 343;
	{8'd214,8'd130} : s = 344;
	{8'd214,8'd131} : s = 345;
	{8'd214,8'd132} : s = 346;
	{8'd214,8'd133} : s = 347;
	{8'd214,8'd134} : s = 348;
	{8'd214,8'd135} : s = 349;
	{8'd214,8'd136} : s = 350;
	{8'd214,8'd137} : s = 351;
	{8'd214,8'd138} : s = 352;
	{8'd214,8'd139} : s = 353;
	{8'd214,8'd140} : s = 354;
	{8'd214,8'd141} : s = 355;
	{8'd214,8'd142} : s = 356;
	{8'd214,8'd143} : s = 357;
	{8'd214,8'd144} : s = 358;
	{8'd214,8'd145} : s = 359;
	{8'd214,8'd146} : s = 360;
	{8'd214,8'd147} : s = 361;
	{8'd214,8'd148} : s = 362;
	{8'd214,8'd149} : s = 363;
	{8'd214,8'd150} : s = 364;
	{8'd214,8'd151} : s = 365;
	{8'd214,8'd152} : s = 366;
	{8'd214,8'd153} : s = 367;
	{8'd214,8'd154} : s = 368;
	{8'd214,8'd155} : s = 369;
	{8'd214,8'd156} : s = 370;
	{8'd214,8'd157} : s = 371;
	{8'd214,8'd158} : s = 372;
	{8'd214,8'd159} : s = 373;
	{8'd214,8'd160} : s = 374;
	{8'd214,8'd161} : s = 375;
	{8'd214,8'd162} : s = 376;
	{8'd214,8'd163} : s = 377;
	{8'd214,8'd164} : s = 378;
	{8'd214,8'd165} : s = 379;
	{8'd214,8'd166} : s = 380;
	{8'd214,8'd167} : s = 381;
	{8'd214,8'd168} : s = 382;
	{8'd214,8'd169} : s = 383;
	{8'd214,8'd170} : s = 384;
	{8'd214,8'd171} : s = 385;
	{8'd214,8'd172} : s = 386;
	{8'd214,8'd173} : s = 387;
	{8'd214,8'd174} : s = 388;
	{8'd214,8'd175} : s = 389;
	{8'd214,8'd176} : s = 390;
	{8'd214,8'd177} : s = 391;
	{8'd214,8'd178} : s = 392;
	{8'd214,8'd179} : s = 393;
	{8'd214,8'd180} : s = 394;
	{8'd214,8'd181} : s = 395;
	{8'd214,8'd182} : s = 396;
	{8'd214,8'd183} : s = 397;
	{8'd214,8'd184} : s = 398;
	{8'd214,8'd185} : s = 399;
	{8'd214,8'd186} : s = 400;
	{8'd214,8'd187} : s = 401;
	{8'd214,8'd188} : s = 402;
	{8'd214,8'd189} : s = 403;
	{8'd214,8'd190} : s = 404;
	{8'd214,8'd191} : s = 405;
	{8'd214,8'd192} : s = 406;
	{8'd214,8'd193} : s = 407;
	{8'd214,8'd194} : s = 408;
	{8'd214,8'd195} : s = 409;
	{8'd214,8'd196} : s = 410;
	{8'd214,8'd197} : s = 411;
	{8'd214,8'd198} : s = 412;
	{8'd214,8'd199} : s = 413;
	{8'd214,8'd200} : s = 414;
	{8'd214,8'd201} : s = 415;
	{8'd214,8'd202} : s = 416;
	{8'd214,8'd203} : s = 417;
	{8'd214,8'd204} : s = 418;
	{8'd214,8'd205} : s = 419;
	{8'd214,8'd206} : s = 420;
	{8'd214,8'd207} : s = 421;
	{8'd214,8'd208} : s = 422;
	{8'd214,8'd209} : s = 423;
	{8'd214,8'd210} : s = 424;
	{8'd214,8'd211} : s = 425;
	{8'd214,8'd212} : s = 426;
	{8'd214,8'd213} : s = 427;
	{8'd214,8'd214} : s = 428;
	{8'd214,8'd215} : s = 429;
	{8'd214,8'd216} : s = 430;
	{8'd214,8'd217} : s = 431;
	{8'd214,8'd218} : s = 432;
	{8'd214,8'd219} : s = 433;
	{8'd214,8'd220} : s = 434;
	{8'd214,8'd221} : s = 435;
	{8'd214,8'd222} : s = 436;
	{8'd214,8'd223} : s = 437;
	{8'd214,8'd224} : s = 438;
	{8'd214,8'd225} : s = 439;
	{8'd214,8'd226} : s = 440;
	{8'd214,8'd227} : s = 441;
	{8'd214,8'd228} : s = 442;
	{8'd214,8'd229} : s = 443;
	{8'd214,8'd230} : s = 444;
	{8'd214,8'd231} : s = 445;
	{8'd214,8'd232} : s = 446;
	{8'd214,8'd233} : s = 447;
	{8'd214,8'd234} : s = 448;
	{8'd214,8'd235} : s = 449;
	{8'd214,8'd236} : s = 450;
	{8'd214,8'd237} : s = 451;
	{8'd214,8'd238} : s = 452;
	{8'd214,8'd239} : s = 453;
	{8'd214,8'd240} : s = 454;
	{8'd214,8'd241} : s = 455;
	{8'd214,8'd242} : s = 456;
	{8'd214,8'd243} : s = 457;
	{8'd214,8'd244} : s = 458;
	{8'd214,8'd245} : s = 459;
	{8'd214,8'd246} : s = 460;
	{8'd214,8'd247} : s = 461;
	{8'd214,8'd248} : s = 462;
	{8'd214,8'd249} : s = 463;
	{8'd214,8'd250} : s = 464;
	{8'd214,8'd251} : s = 465;
	{8'd214,8'd252} : s = 466;
	{8'd214,8'd253} : s = 467;
	{8'd214,8'd254} : s = 468;
	{8'd214,8'd255} : s = 469;
	{8'd215,8'd0} : s = 215;
	{8'd215,8'd1} : s = 216;
	{8'd215,8'd2} : s = 217;
	{8'd215,8'd3} : s = 218;
	{8'd215,8'd4} : s = 219;
	{8'd215,8'd5} : s = 220;
	{8'd215,8'd6} : s = 221;
	{8'd215,8'd7} : s = 222;
	{8'd215,8'd8} : s = 223;
	{8'd215,8'd9} : s = 224;
	{8'd215,8'd10} : s = 225;
	{8'd215,8'd11} : s = 226;
	{8'd215,8'd12} : s = 227;
	{8'd215,8'd13} : s = 228;
	{8'd215,8'd14} : s = 229;
	{8'd215,8'd15} : s = 230;
	{8'd215,8'd16} : s = 231;
	{8'd215,8'd17} : s = 232;
	{8'd215,8'd18} : s = 233;
	{8'd215,8'd19} : s = 234;
	{8'd215,8'd20} : s = 235;
	{8'd215,8'd21} : s = 236;
	{8'd215,8'd22} : s = 237;
	{8'd215,8'd23} : s = 238;
	{8'd215,8'd24} : s = 239;
	{8'd215,8'd25} : s = 240;
	{8'd215,8'd26} : s = 241;
	{8'd215,8'd27} : s = 242;
	{8'd215,8'd28} : s = 243;
	{8'd215,8'd29} : s = 244;
	{8'd215,8'd30} : s = 245;
	{8'd215,8'd31} : s = 246;
	{8'd215,8'd32} : s = 247;
	{8'd215,8'd33} : s = 248;
	{8'd215,8'd34} : s = 249;
	{8'd215,8'd35} : s = 250;
	{8'd215,8'd36} : s = 251;
	{8'd215,8'd37} : s = 252;
	{8'd215,8'd38} : s = 253;
	{8'd215,8'd39} : s = 254;
	{8'd215,8'd40} : s = 255;
	{8'd215,8'd41} : s = 256;
	{8'd215,8'd42} : s = 257;
	{8'd215,8'd43} : s = 258;
	{8'd215,8'd44} : s = 259;
	{8'd215,8'd45} : s = 260;
	{8'd215,8'd46} : s = 261;
	{8'd215,8'd47} : s = 262;
	{8'd215,8'd48} : s = 263;
	{8'd215,8'd49} : s = 264;
	{8'd215,8'd50} : s = 265;
	{8'd215,8'd51} : s = 266;
	{8'd215,8'd52} : s = 267;
	{8'd215,8'd53} : s = 268;
	{8'd215,8'd54} : s = 269;
	{8'd215,8'd55} : s = 270;
	{8'd215,8'd56} : s = 271;
	{8'd215,8'd57} : s = 272;
	{8'd215,8'd58} : s = 273;
	{8'd215,8'd59} : s = 274;
	{8'd215,8'd60} : s = 275;
	{8'd215,8'd61} : s = 276;
	{8'd215,8'd62} : s = 277;
	{8'd215,8'd63} : s = 278;
	{8'd215,8'd64} : s = 279;
	{8'd215,8'd65} : s = 280;
	{8'd215,8'd66} : s = 281;
	{8'd215,8'd67} : s = 282;
	{8'd215,8'd68} : s = 283;
	{8'd215,8'd69} : s = 284;
	{8'd215,8'd70} : s = 285;
	{8'd215,8'd71} : s = 286;
	{8'd215,8'd72} : s = 287;
	{8'd215,8'd73} : s = 288;
	{8'd215,8'd74} : s = 289;
	{8'd215,8'd75} : s = 290;
	{8'd215,8'd76} : s = 291;
	{8'd215,8'd77} : s = 292;
	{8'd215,8'd78} : s = 293;
	{8'd215,8'd79} : s = 294;
	{8'd215,8'd80} : s = 295;
	{8'd215,8'd81} : s = 296;
	{8'd215,8'd82} : s = 297;
	{8'd215,8'd83} : s = 298;
	{8'd215,8'd84} : s = 299;
	{8'd215,8'd85} : s = 300;
	{8'd215,8'd86} : s = 301;
	{8'd215,8'd87} : s = 302;
	{8'd215,8'd88} : s = 303;
	{8'd215,8'd89} : s = 304;
	{8'd215,8'd90} : s = 305;
	{8'd215,8'd91} : s = 306;
	{8'd215,8'd92} : s = 307;
	{8'd215,8'd93} : s = 308;
	{8'd215,8'd94} : s = 309;
	{8'd215,8'd95} : s = 310;
	{8'd215,8'd96} : s = 311;
	{8'd215,8'd97} : s = 312;
	{8'd215,8'd98} : s = 313;
	{8'd215,8'd99} : s = 314;
	{8'd215,8'd100} : s = 315;
	{8'd215,8'd101} : s = 316;
	{8'd215,8'd102} : s = 317;
	{8'd215,8'd103} : s = 318;
	{8'd215,8'd104} : s = 319;
	{8'd215,8'd105} : s = 320;
	{8'd215,8'd106} : s = 321;
	{8'd215,8'd107} : s = 322;
	{8'd215,8'd108} : s = 323;
	{8'd215,8'd109} : s = 324;
	{8'd215,8'd110} : s = 325;
	{8'd215,8'd111} : s = 326;
	{8'd215,8'd112} : s = 327;
	{8'd215,8'd113} : s = 328;
	{8'd215,8'd114} : s = 329;
	{8'd215,8'd115} : s = 330;
	{8'd215,8'd116} : s = 331;
	{8'd215,8'd117} : s = 332;
	{8'd215,8'd118} : s = 333;
	{8'd215,8'd119} : s = 334;
	{8'd215,8'd120} : s = 335;
	{8'd215,8'd121} : s = 336;
	{8'd215,8'd122} : s = 337;
	{8'd215,8'd123} : s = 338;
	{8'd215,8'd124} : s = 339;
	{8'd215,8'd125} : s = 340;
	{8'd215,8'd126} : s = 341;
	{8'd215,8'd127} : s = 342;
	{8'd215,8'd128} : s = 343;
	{8'd215,8'd129} : s = 344;
	{8'd215,8'd130} : s = 345;
	{8'd215,8'd131} : s = 346;
	{8'd215,8'd132} : s = 347;
	{8'd215,8'd133} : s = 348;
	{8'd215,8'd134} : s = 349;
	{8'd215,8'd135} : s = 350;
	{8'd215,8'd136} : s = 351;
	{8'd215,8'd137} : s = 352;
	{8'd215,8'd138} : s = 353;
	{8'd215,8'd139} : s = 354;
	{8'd215,8'd140} : s = 355;
	{8'd215,8'd141} : s = 356;
	{8'd215,8'd142} : s = 357;
	{8'd215,8'd143} : s = 358;
	{8'd215,8'd144} : s = 359;
	{8'd215,8'd145} : s = 360;
	{8'd215,8'd146} : s = 361;
	{8'd215,8'd147} : s = 362;
	{8'd215,8'd148} : s = 363;
	{8'd215,8'd149} : s = 364;
	{8'd215,8'd150} : s = 365;
	{8'd215,8'd151} : s = 366;
	{8'd215,8'd152} : s = 367;
	{8'd215,8'd153} : s = 368;
	{8'd215,8'd154} : s = 369;
	{8'd215,8'd155} : s = 370;
	{8'd215,8'd156} : s = 371;
	{8'd215,8'd157} : s = 372;
	{8'd215,8'd158} : s = 373;
	{8'd215,8'd159} : s = 374;
	{8'd215,8'd160} : s = 375;
	{8'd215,8'd161} : s = 376;
	{8'd215,8'd162} : s = 377;
	{8'd215,8'd163} : s = 378;
	{8'd215,8'd164} : s = 379;
	{8'd215,8'd165} : s = 380;
	{8'd215,8'd166} : s = 381;
	{8'd215,8'd167} : s = 382;
	{8'd215,8'd168} : s = 383;
	{8'd215,8'd169} : s = 384;
	{8'd215,8'd170} : s = 385;
	{8'd215,8'd171} : s = 386;
	{8'd215,8'd172} : s = 387;
	{8'd215,8'd173} : s = 388;
	{8'd215,8'd174} : s = 389;
	{8'd215,8'd175} : s = 390;
	{8'd215,8'd176} : s = 391;
	{8'd215,8'd177} : s = 392;
	{8'd215,8'd178} : s = 393;
	{8'd215,8'd179} : s = 394;
	{8'd215,8'd180} : s = 395;
	{8'd215,8'd181} : s = 396;
	{8'd215,8'd182} : s = 397;
	{8'd215,8'd183} : s = 398;
	{8'd215,8'd184} : s = 399;
	{8'd215,8'd185} : s = 400;
	{8'd215,8'd186} : s = 401;
	{8'd215,8'd187} : s = 402;
	{8'd215,8'd188} : s = 403;
	{8'd215,8'd189} : s = 404;
	{8'd215,8'd190} : s = 405;
	{8'd215,8'd191} : s = 406;
	{8'd215,8'd192} : s = 407;
	{8'd215,8'd193} : s = 408;
	{8'd215,8'd194} : s = 409;
	{8'd215,8'd195} : s = 410;
	{8'd215,8'd196} : s = 411;
	{8'd215,8'd197} : s = 412;
	{8'd215,8'd198} : s = 413;
	{8'd215,8'd199} : s = 414;
	{8'd215,8'd200} : s = 415;
	{8'd215,8'd201} : s = 416;
	{8'd215,8'd202} : s = 417;
	{8'd215,8'd203} : s = 418;
	{8'd215,8'd204} : s = 419;
	{8'd215,8'd205} : s = 420;
	{8'd215,8'd206} : s = 421;
	{8'd215,8'd207} : s = 422;
	{8'd215,8'd208} : s = 423;
	{8'd215,8'd209} : s = 424;
	{8'd215,8'd210} : s = 425;
	{8'd215,8'd211} : s = 426;
	{8'd215,8'd212} : s = 427;
	{8'd215,8'd213} : s = 428;
	{8'd215,8'd214} : s = 429;
	{8'd215,8'd215} : s = 430;
	{8'd215,8'd216} : s = 431;
	{8'd215,8'd217} : s = 432;
	{8'd215,8'd218} : s = 433;
	{8'd215,8'd219} : s = 434;
	{8'd215,8'd220} : s = 435;
	{8'd215,8'd221} : s = 436;
	{8'd215,8'd222} : s = 437;
	{8'd215,8'd223} : s = 438;
	{8'd215,8'd224} : s = 439;
	{8'd215,8'd225} : s = 440;
	{8'd215,8'd226} : s = 441;
	{8'd215,8'd227} : s = 442;
	{8'd215,8'd228} : s = 443;
	{8'd215,8'd229} : s = 444;
	{8'd215,8'd230} : s = 445;
	{8'd215,8'd231} : s = 446;
	{8'd215,8'd232} : s = 447;
	{8'd215,8'd233} : s = 448;
	{8'd215,8'd234} : s = 449;
	{8'd215,8'd235} : s = 450;
	{8'd215,8'd236} : s = 451;
	{8'd215,8'd237} : s = 452;
	{8'd215,8'd238} : s = 453;
	{8'd215,8'd239} : s = 454;
	{8'd215,8'd240} : s = 455;
	{8'd215,8'd241} : s = 456;
	{8'd215,8'd242} : s = 457;
	{8'd215,8'd243} : s = 458;
	{8'd215,8'd244} : s = 459;
	{8'd215,8'd245} : s = 460;
	{8'd215,8'd246} : s = 461;
	{8'd215,8'd247} : s = 462;
	{8'd215,8'd248} : s = 463;
	{8'd215,8'd249} : s = 464;
	{8'd215,8'd250} : s = 465;
	{8'd215,8'd251} : s = 466;
	{8'd215,8'd252} : s = 467;
	{8'd215,8'd253} : s = 468;
	{8'd215,8'd254} : s = 469;
	{8'd215,8'd255} : s = 470;
	{8'd216,8'd0} : s = 216;
	{8'd216,8'd1} : s = 217;
	{8'd216,8'd2} : s = 218;
	{8'd216,8'd3} : s = 219;
	{8'd216,8'd4} : s = 220;
	{8'd216,8'd5} : s = 221;
	{8'd216,8'd6} : s = 222;
	{8'd216,8'd7} : s = 223;
	{8'd216,8'd8} : s = 224;
	{8'd216,8'd9} : s = 225;
	{8'd216,8'd10} : s = 226;
	{8'd216,8'd11} : s = 227;
	{8'd216,8'd12} : s = 228;
	{8'd216,8'd13} : s = 229;
	{8'd216,8'd14} : s = 230;
	{8'd216,8'd15} : s = 231;
	{8'd216,8'd16} : s = 232;
	{8'd216,8'd17} : s = 233;
	{8'd216,8'd18} : s = 234;
	{8'd216,8'd19} : s = 235;
	{8'd216,8'd20} : s = 236;
	{8'd216,8'd21} : s = 237;
	{8'd216,8'd22} : s = 238;
	{8'd216,8'd23} : s = 239;
	{8'd216,8'd24} : s = 240;
	{8'd216,8'd25} : s = 241;
	{8'd216,8'd26} : s = 242;
	{8'd216,8'd27} : s = 243;
	{8'd216,8'd28} : s = 244;
	{8'd216,8'd29} : s = 245;
	{8'd216,8'd30} : s = 246;
	{8'd216,8'd31} : s = 247;
	{8'd216,8'd32} : s = 248;
	{8'd216,8'd33} : s = 249;
	{8'd216,8'd34} : s = 250;
	{8'd216,8'd35} : s = 251;
	{8'd216,8'd36} : s = 252;
	{8'd216,8'd37} : s = 253;
	{8'd216,8'd38} : s = 254;
	{8'd216,8'd39} : s = 255;
	{8'd216,8'd40} : s = 256;
	{8'd216,8'd41} : s = 257;
	{8'd216,8'd42} : s = 258;
	{8'd216,8'd43} : s = 259;
	{8'd216,8'd44} : s = 260;
	{8'd216,8'd45} : s = 261;
	{8'd216,8'd46} : s = 262;
	{8'd216,8'd47} : s = 263;
	{8'd216,8'd48} : s = 264;
	{8'd216,8'd49} : s = 265;
	{8'd216,8'd50} : s = 266;
	{8'd216,8'd51} : s = 267;
	{8'd216,8'd52} : s = 268;
	{8'd216,8'd53} : s = 269;
	{8'd216,8'd54} : s = 270;
	{8'd216,8'd55} : s = 271;
	{8'd216,8'd56} : s = 272;
	{8'd216,8'd57} : s = 273;
	{8'd216,8'd58} : s = 274;
	{8'd216,8'd59} : s = 275;
	{8'd216,8'd60} : s = 276;
	{8'd216,8'd61} : s = 277;
	{8'd216,8'd62} : s = 278;
	{8'd216,8'd63} : s = 279;
	{8'd216,8'd64} : s = 280;
	{8'd216,8'd65} : s = 281;
	{8'd216,8'd66} : s = 282;
	{8'd216,8'd67} : s = 283;
	{8'd216,8'd68} : s = 284;
	{8'd216,8'd69} : s = 285;
	{8'd216,8'd70} : s = 286;
	{8'd216,8'd71} : s = 287;
	{8'd216,8'd72} : s = 288;
	{8'd216,8'd73} : s = 289;
	{8'd216,8'd74} : s = 290;
	{8'd216,8'd75} : s = 291;
	{8'd216,8'd76} : s = 292;
	{8'd216,8'd77} : s = 293;
	{8'd216,8'd78} : s = 294;
	{8'd216,8'd79} : s = 295;
	{8'd216,8'd80} : s = 296;
	{8'd216,8'd81} : s = 297;
	{8'd216,8'd82} : s = 298;
	{8'd216,8'd83} : s = 299;
	{8'd216,8'd84} : s = 300;
	{8'd216,8'd85} : s = 301;
	{8'd216,8'd86} : s = 302;
	{8'd216,8'd87} : s = 303;
	{8'd216,8'd88} : s = 304;
	{8'd216,8'd89} : s = 305;
	{8'd216,8'd90} : s = 306;
	{8'd216,8'd91} : s = 307;
	{8'd216,8'd92} : s = 308;
	{8'd216,8'd93} : s = 309;
	{8'd216,8'd94} : s = 310;
	{8'd216,8'd95} : s = 311;
	{8'd216,8'd96} : s = 312;
	{8'd216,8'd97} : s = 313;
	{8'd216,8'd98} : s = 314;
	{8'd216,8'd99} : s = 315;
	{8'd216,8'd100} : s = 316;
	{8'd216,8'd101} : s = 317;
	{8'd216,8'd102} : s = 318;
	{8'd216,8'd103} : s = 319;
	{8'd216,8'd104} : s = 320;
	{8'd216,8'd105} : s = 321;
	{8'd216,8'd106} : s = 322;
	{8'd216,8'd107} : s = 323;
	{8'd216,8'd108} : s = 324;
	{8'd216,8'd109} : s = 325;
	{8'd216,8'd110} : s = 326;
	{8'd216,8'd111} : s = 327;
	{8'd216,8'd112} : s = 328;
	{8'd216,8'd113} : s = 329;
	{8'd216,8'd114} : s = 330;
	{8'd216,8'd115} : s = 331;
	{8'd216,8'd116} : s = 332;
	{8'd216,8'd117} : s = 333;
	{8'd216,8'd118} : s = 334;
	{8'd216,8'd119} : s = 335;
	{8'd216,8'd120} : s = 336;
	{8'd216,8'd121} : s = 337;
	{8'd216,8'd122} : s = 338;
	{8'd216,8'd123} : s = 339;
	{8'd216,8'd124} : s = 340;
	{8'd216,8'd125} : s = 341;
	{8'd216,8'd126} : s = 342;
	{8'd216,8'd127} : s = 343;
	{8'd216,8'd128} : s = 344;
	{8'd216,8'd129} : s = 345;
	{8'd216,8'd130} : s = 346;
	{8'd216,8'd131} : s = 347;
	{8'd216,8'd132} : s = 348;
	{8'd216,8'd133} : s = 349;
	{8'd216,8'd134} : s = 350;
	{8'd216,8'd135} : s = 351;
	{8'd216,8'd136} : s = 352;
	{8'd216,8'd137} : s = 353;
	{8'd216,8'd138} : s = 354;
	{8'd216,8'd139} : s = 355;
	{8'd216,8'd140} : s = 356;
	{8'd216,8'd141} : s = 357;
	{8'd216,8'd142} : s = 358;
	{8'd216,8'd143} : s = 359;
	{8'd216,8'd144} : s = 360;
	{8'd216,8'd145} : s = 361;
	{8'd216,8'd146} : s = 362;
	{8'd216,8'd147} : s = 363;
	{8'd216,8'd148} : s = 364;
	{8'd216,8'd149} : s = 365;
	{8'd216,8'd150} : s = 366;
	{8'd216,8'd151} : s = 367;
	{8'd216,8'd152} : s = 368;
	{8'd216,8'd153} : s = 369;
	{8'd216,8'd154} : s = 370;
	{8'd216,8'd155} : s = 371;
	{8'd216,8'd156} : s = 372;
	{8'd216,8'd157} : s = 373;
	{8'd216,8'd158} : s = 374;
	{8'd216,8'd159} : s = 375;
	{8'd216,8'd160} : s = 376;
	{8'd216,8'd161} : s = 377;
	{8'd216,8'd162} : s = 378;
	{8'd216,8'd163} : s = 379;
	{8'd216,8'd164} : s = 380;
	{8'd216,8'd165} : s = 381;
	{8'd216,8'd166} : s = 382;
	{8'd216,8'd167} : s = 383;
	{8'd216,8'd168} : s = 384;
	{8'd216,8'd169} : s = 385;
	{8'd216,8'd170} : s = 386;
	{8'd216,8'd171} : s = 387;
	{8'd216,8'd172} : s = 388;
	{8'd216,8'd173} : s = 389;
	{8'd216,8'd174} : s = 390;
	{8'd216,8'd175} : s = 391;
	{8'd216,8'd176} : s = 392;
	{8'd216,8'd177} : s = 393;
	{8'd216,8'd178} : s = 394;
	{8'd216,8'd179} : s = 395;
	{8'd216,8'd180} : s = 396;
	{8'd216,8'd181} : s = 397;
	{8'd216,8'd182} : s = 398;
	{8'd216,8'd183} : s = 399;
	{8'd216,8'd184} : s = 400;
	{8'd216,8'd185} : s = 401;
	{8'd216,8'd186} : s = 402;
	{8'd216,8'd187} : s = 403;
	{8'd216,8'd188} : s = 404;
	{8'd216,8'd189} : s = 405;
	{8'd216,8'd190} : s = 406;
	{8'd216,8'd191} : s = 407;
	{8'd216,8'd192} : s = 408;
	{8'd216,8'd193} : s = 409;
	{8'd216,8'd194} : s = 410;
	{8'd216,8'd195} : s = 411;
	{8'd216,8'd196} : s = 412;
	{8'd216,8'd197} : s = 413;
	{8'd216,8'd198} : s = 414;
	{8'd216,8'd199} : s = 415;
	{8'd216,8'd200} : s = 416;
	{8'd216,8'd201} : s = 417;
	{8'd216,8'd202} : s = 418;
	{8'd216,8'd203} : s = 419;
	{8'd216,8'd204} : s = 420;
	{8'd216,8'd205} : s = 421;
	{8'd216,8'd206} : s = 422;
	{8'd216,8'd207} : s = 423;
	{8'd216,8'd208} : s = 424;
	{8'd216,8'd209} : s = 425;
	{8'd216,8'd210} : s = 426;
	{8'd216,8'd211} : s = 427;
	{8'd216,8'd212} : s = 428;
	{8'd216,8'd213} : s = 429;
	{8'd216,8'd214} : s = 430;
	{8'd216,8'd215} : s = 431;
	{8'd216,8'd216} : s = 432;
	{8'd216,8'd217} : s = 433;
	{8'd216,8'd218} : s = 434;
	{8'd216,8'd219} : s = 435;
	{8'd216,8'd220} : s = 436;
	{8'd216,8'd221} : s = 437;
	{8'd216,8'd222} : s = 438;
	{8'd216,8'd223} : s = 439;
	{8'd216,8'd224} : s = 440;
	{8'd216,8'd225} : s = 441;
	{8'd216,8'd226} : s = 442;
	{8'd216,8'd227} : s = 443;
	{8'd216,8'd228} : s = 444;
	{8'd216,8'd229} : s = 445;
	{8'd216,8'd230} : s = 446;
	{8'd216,8'd231} : s = 447;
	{8'd216,8'd232} : s = 448;
	{8'd216,8'd233} : s = 449;
	{8'd216,8'd234} : s = 450;
	{8'd216,8'd235} : s = 451;
	{8'd216,8'd236} : s = 452;
	{8'd216,8'd237} : s = 453;
	{8'd216,8'd238} : s = 454;
	{8'd216,8'd239} : s = 455;
	{8'd216,8'd240} : s = 456;
	{8'd216,8'd241} : s = 457;
	{8'd216,8'd242} : s = 458;
	{8'd216,8'd243} : s = 459;
	{8'd216,8'd244} : s = 460;
	{8'd216,8'd245} : s = 461;
	{8'd216,8'd246} : s = 462;
	{8'd216,8'd247} : s = 463;
	{8'd216,8'd248} : s = 464;
	{8'd216,8'd249} : s = 465;
	{8'd216,8'd250} : s = 466;
	{8'd216,8'd251} : s = 467;
	{8'd216,8'd252} : s = 468;
	{8'd216,8'd253} : s = 469;
	{8'd216,8'd254} : s = 470;
	{8'd216,8'd255} : s = 471;
	{8'd217,8'd0} : s = 217;
	{8'd217,8'd1} : s = 218;
	{8'd217,8'd2} : s = 219;
	{8'd217,8'd3} : s = 220;
	{8'd217,8'd4} : s = 221;
	{8'd217,8'd5} : s = 222;
	{8'd217,8'd6} : s = 223;
	{8'd217,8'd7} : s = 224;
	{8'd217,8'd8} : s = 225;
	{8'd217,8'd9} : s = 226;
	{8'd217,8'd10} : s = 227;
	{8'd217,8'd11} : s = 228;
	{8'd217,8'd12} : s = 229;
	{8'd217,8'd13} : s = 230;
	{8'd217,8'd14} : s = 231;
	{8'd217,8'd15} : s = 232;
	{8'd217,8'd16} : s = 233;
	{8'd217,8'd17} : s = 234;
	{8'd217,8'd18} : s = 235;
	{8'd217,8'd19} : s = 236;
	{8'd217,8'd20} : s = 237;
	{8'd217,8'd21} : s = 238;
	{8'd217,8'd22} : s = 239;
	{8'd217,8'd23} : s = 240;
	{8'd217,8'd24} : s = 241;
	{8'd217,8'd25} : s = 242;
	{8'd217,8'd26} : s = 243;
	{8'd217,8'd27} : s = 244;
	{8'd217,8'd28} : s = 245;
	{8'd217,8'd29} : s = 246;
	{8'd217,8'd30} : s = 247;
	{8'd217,8'd31} : s = 248;
	{8'd217,8'd32} : s = 249;
	{8'd217,8'd33} : s = 250;
	{8'd217,8'd34} : s = 251;
	{8'd217,8'd35} : s = 252;
	{8'd217,8'd36} : s = 253;
	{8'd217,8'd37} : s = 254;
	{8'd217,8'd38} : s = 255;
	{8'd217,8'd39} : s = 256;
	{8'd217,8'd40} : s = 257;
	{8'd217,8'd41} : s = 258;
	{8'd217,8'd42} : s = 259;
	{8'd217,8'd43} : s = 260;
	{8'd217,8'd44} : s = 261;
	{8'd217,8'd45} : s = 262;
	{8'd217,8'd46} : s = 263;
	{8'd217,8'd47} : s = 264;
	{8'd217,8'd48} : s = 265;
	{8'd217,8'd49} : s = 266;
	{8'd217,8'd50} : s = 267;
	{8'd217,8'd51} : s = 268;
	{8'd217,8'd52} : s = 269;
	{8'd217,8'd53} : s = 270;
	{8'd217,8'd54} : s = 271;
	{8'd217,8'd55} : s = 272;
	{8'd217,8'd56} : s = 273;
	{8'd217,8'd57} : s = 274;
	{8'd217,8'd58} : s = 275;
	{8'd217,8'd59} : s = 276;
	{8'd217,8'd60} : s = 277;
	{8'd217,8'd61} : s = 278;
	{8'd217,8'd62} : s = 279;
	{8'd217,8'd63} : s = 280;
	{8'd217,8'd64} : s = 281;
	{8'd217,8'd65} : s = 282;
	{8'd217,8'd66} : s = 283;
	{8'd217,8'd67} : s = 284;
	{8'd217,8'd68} : s = 285;
	{8'd217,8'd69} : s = 286;
	{8'd217,8'd70} : s = 287;
	{8'd217,8'd71} : s = 288;
	{8'd217,8'd72} : s = 289;
	{8'd217,8'd73} : s = 290;
	{8'd217,8'd74} : s = 291;
	{8'd217,8'd75} : s = 292;
	{8'd217,8'd76} : s = 293;
	{8'd217,8'd77} : s = 294;
	{8'd217,8'd78} : s = 295;
	{8'd217,8'd79} : s = 296;
	{8'd217,8'd80} : s = 297;
	{8'd217,8'd81} : s = 298;
	{8'd217,8'd82} : s = 299;
	{8'd217,8'd83} : s = 300;
	{8'd217,8'd84} : s = 301;
	{8'd217,8'd85} : s = 302;
	{8'd217,8'd86} : s = 303;
	{8'd217,8'd87} : s = 304;
	{8'd217,8'd88} : s = 305;
	{8'd217,8'd89} : s = 306;
	{8'd217,8'd90} : s = 307;
	{8'd217,8'd91} : s = 308;
	{8'd217,8'd92} : s = 309;
	{8'd217,8'd93} : s = 310;
	{8'd217,8'd94} : s = 311;
	{8'd217,8'd95} : s = 312;
	{8'd217,8'd96} : s = 313;
	{8'd217,8'd97} : s = 314;
	{8'd217,8'd98} : s = 315;
	{8'd217,8'd99} : s = 316;
	{8'd217,8'd100} : s = 317;
	{8'd217,8'd101} : s = 318;
	{8'd217,8'd102} : s = 319;
	{8'd217,8'd103} : s = 320;
	{8'd217,8'd104} : s = 321;
	{8'd217,8'd105} : s = 322;
	{8'd217,8'd106} : s = 323;
	{8'd217,8'd107} : s = 324;
	{8'd217,8'd108} : s = 325;
	{8'd217,8'd109} : s = 326;
	{8'd217,8'd110} : s = 327;
	{8'd217,8'd111} : s = 328;
	{8'd217,8'd112} : s = 329;
	{8'd217,8'd113} : s = 330;
	{8'd217,8'd114} : s = 331;
	{8'd217,8'd115} : s = 332;
	{8'd217,8'd116} : s = 333;
	{8'd217,8'd117} : s = 334;
	{8'd217,8'd118} : s = 335;
	{8'd217,8'd119} : s = 336;
	{8'd217,8'd120} : s = 337;
	{8'd217,8'd121} : s = 338;
	{8'd217,8'd122} : s = 339;
	{8'd217,8'd123} : s = 340;
	{8'd217,8'd124} : s = 341;
	{8'd217,8'd125} : s = 342;
	{8'd217,8'd126} : s = 343;
	{8'd217,8'd127} : s = 344;
	{8'd217,8'd128} : s = 345;
	{8'd217,8'd129} : s = 346;
	{8'd217,8'd130} : s = 347;
	{8'd217,8'd131} : s = 348;
	{8'd217,8'd132} : s = 349;
	{8'd217,8'd133} : s = 350;
	{8'd217,8'd134} : s = 351;
	{8'd217,8'd135} : s = 352;
	{8'd217,8'd136} : s = 353;
	{8'd217,8'd137} : s = 354;
	{8'd217,8'd138} : s = 355;
	{8'd217,8'd139} : s = 356;
	{8'd217,8'd140} : s = 357;
	{8'd217,8'd141} : s = 358;
	{8'd217,8'd142} : s = 359;
	{8'd217,8'd143} : s = 360;
	{8'd217,8'd144} : s = 361;
	{8'd217,8'd145} : s = 362;
	{8'd217,8'd146} : s = 363;
	{8'd217,8'd147} : s = 364;
	{8'd217,8'd148} : s = 365;
	{8'd217,8'd149} : s = 366;
	{8'd217,8'd150} : s = 367;
	{8'd217,8'd151} : s = 368;
	{8'd217,8'd152} : s = 369;
	{8'd217,8'd153} : s = 370;
	{8'd217,8'd154} : s = 371;
	{8'd217,8'd155} : s = 372;
	{8'd217,8'd156} : s = 373;
	{8'd217,8'd157} : s = 374;
	{8'd217,8'd158} : s = 375;
	{8'd217,8'd159} : s = 376;
	{8'd217,8'd160} : s = 377;
	{8'd217,8'd161} : s = 378;
	{8'd217,8'd162} : s = 379;
	{8'd217,8'd163} : s = 380;
	{8'd217,8'd164} : s = 381;
	{8'd217,8'd165} : s = 382;
	{8'd217,8'd166} : s = 383;
	{8'd217,8'd167} : s = 384;
	{8'd217,8'd168} : s = 385;
	{8'd217,8'd169} : s = 386;
	{8'd217,8'd170} : s = 387;
	{8'd217,8'd171} : s = 388;
	{8'd217,8'd172} : s = 389;
	{8'd217,8'd173} : s = 390;
	{8'd217,8'd174} : s = 391;
	{8'd217,8'd175} : s = 392;
	{8'd217,8'd176} : s = 393;
	{8'd217,8'd177} : s = 394;
	{8'd217,8'd178} : s = 395;
	{8'd217,8'd179} : s = 396;
	{8'd217,8'd180} : s = 397;
	{8'd217,8'd181} : s = 398;
	{8'd217,8'd182} : s = 399;
	{8'd217,8'd183} : s = 400;
	{8'd217,8'd184} : s = 401;
	{8'd217,8'd185} : s = 402;
	{8'd217,8'd186} : s = 403;
	{8'd217,8'd187} : s = 404;
	{8'd217,8'd188} : s = 405;
	{8'd217,8'd189} : s = 406;
	{8'd217,8'd190} : s = 407;
	{8'd217,8'd191} : s = 408;
	{8'd217,8'd192} : s = 409;
	{8'd217,8'd193} : s = 410;
	{8'd217,8'd194} : s = 411;
	{8'd217,8'd195} : s = 412;
	{8'd217,8'd196} : s = 413;
	{8'd217,8'd197} : s = 414;
	{8'd217,8'd198} : s = 415;
	{8'd217,8'd199} : s = 416;
	{8'd217,8'd200} : s = 417;
	{8'd217,8'd201} : s = 418;
	{8'd217,8'd202} : s = 419;
	{8'd217,8'd203} : s = 420;
	{8'd217,8'd204} : s = 421;
	{8'd217,8'd205} : s = 422;
	{8'd217,8'd206} : s = 423;
	{8'd217,8'd207} : s = 424;
	{8'd217,8'd208} : s = 425;
	{8'd217,8'd209} : s = 426;
	{8'd217,8'd210} : s = 427;
	{8'd217,8'd211} : s = 428;
	{8'd217,8'd212} : s = 429;
	{8'd217,8'd213} : s = 430;
	{8'd217,8'd214} : s = 431;
	{8'd217,8'd215} : s = 432;
	{8'd217,8'd216} : s = 433;
	{8'd217,8'd217} : s = 434;
	{8'd217,8'd218} : s = 435;
	{8'd217,8'd219} : s = 436;
	{8'd217,8'd220} : s = 437;
	{8'd217,8'd221} : s = 438;
	{8'd217,8'd222} : s = 439;
	{8'd217,8'd223} : s = 440;
	{8'd217,8'd224} : s = 441;
	{8'd217,8'd225} : s = 442;
	{8'd217,8'd226} : s = 443;
	{8'd217,8'd227} : s = 444;
	{8'd217,8'd228} : s = 445;
	{8'd217,8'd229} : s = 446;
	{8'd217,8'd230} : s = 447;
	{8'd217,8'd231} : s = 448;
	{8'd217,8'd232} : s = 449;
	{8'd217,8'd233} : s = 450;
	{8'd217,8'd234} : s = 451;
	{8'd217,8'd235} : s = 452;
	{8'd217,8'd236} : s = 453;
	{8'd217,8'd237} : s = 454;
	{8'd217,8'd238} : s = 455;
	{8'd217,8'd239} : s = 456;
	{8'd217,8'd240} : s = 457;
	{8'd217,8'd241} : s = 458;
	{8'd217,8'd242} : s = 459;
	{8'd217,8'd243} : s = 460;
	{8'd217,8'd244} : s = 461;
	{8'd217,8'd245} : s = 462;
	{8'd217,8'd246} : s = 463;
	{8'd217,8'd247} : s = 464;
	{8'd217,8'd248} : s = 465;
	{8'd217,8'd249} : s = 466;
	{8'd217,8'd250} : s = 467;
	{8'd217,8'd251} : s = 468;
	{8'd217,8'd252} : s = 469;
	{8'd217,8'd253} : s = 470;
	{8'd217,8'd254} : s = 471;
	{8'd217,8'd255} : s = 472;
	{8'd218,8'd0} : s = 218;
	{8'd218,8'd1} : s = 219;
	{8'd218,8'd2} : s = 220;
	{8'd218,8'd3} : s = 221;
	{8'd218,8'd4} : s = 222;
	{8'd218,8'd5} : s = 223;
	{8'd218,8'd6} : s = 224;
	{8'd218,8'd7} : s = 225;
	{8'd218,8'd8} : s = 226;
	{8'd218,8'd9} : s = 227;
	{8'd218,8'd10} : s = 228;
	{8'd218,8'd11} : s = 229;
	{8'd218,8'd12} : s = 230;
	{8'd218,8'd13} : s = 231;
	{8'd218,8'd14} : s = 232;
	{8'd218,8'd15} : s = 233;
	{8'd218,8'd16} : s = 234;
	{8'd218,8'd17} : s = 235;
	{8'd218,8'd18} : s = 236;
	{8'd218,8'd19} : s = 237;
	{8'd218,8'd20} : s = 238;
	{8'd218,8'd21} : s = 239;
	{8'd218,8'd22} : s = 240;
	{8'd218,8'd23} : s = 241;
	{8'd218,8'd24} : s = 242;
	{8'd218,8'd25} : s = 243;
	{8'd218,8'd26} : s = 244;
	{8'd218,8'd27} : s = 245;
	{8'd218,8'd28} : s = 246;
	{8'd218,8'd29} : s = 247;
	{8'd218,8'd30} : s = 248;
	{8'd218,8'd31} : s = 249;
	{8'd218,8'd32} : s = 250;
	{8'd218,8'd33} : s = 251;
	{8'd218,8'd34} : s = 252;
	{8'd218,8'd35} : s = 253;
	{8'd218,8'd36} : s = 254;
	{8'd218,8'd37} : s = 255;
	{8'd218,8'd38} : s = 256;
	{8'd218,8'd39} : s = 257;
	{8'd218,8'd40} : s = 258;
	{8'd218,8'd41} : s = 259;
	{8'd218,8'd42} : s = 260;
	{8'd218,8'd43} : s = 261;
	{8'd218,8'd44} : s = 262;
	{8'd218,8'd45} : s = 263;
	{8'd218,8'd46} : s = 264;
	{8'd218,8'd47} : s = 265;
	{8'd218,8'd48} : s = 266;
	{8'd218,8'd49} : s = 267;
	{8'd218,8'd50} : s = 268;
	{8'd218,8'd51} : s = 269;
	{8'd218,8'd52} : s = 270;
	{8'd218,8'd53} : s = 271;
	{8'd218,8'd54} : s = 272;
	{8'd218,8'd55} : s = 273;
	{8'd218,8'd56} : s = 274;
	{8'd218,8'd57} : s = 275;
	{8'd218,8'd58} : s = 276;
	{8'd218,8'd59} : s = 277;
	{8'd218,8'd60} : s = 278;
	{8'd218,8'd61} : s = 279;
	{8'd218,8'd62} : s = 280;
	{8'd218,8'd63} : s = 281;
	{8'd218,8'd64} : s = 282;
	{8'd218,8'd65} : s = 283;
	{8'd218,8'd66} : s = 284;
	{8'd218,8'd67} : s = 285;
	{8'd218,8'd68} : s = 286;
	{8'd218,8'd69} : s = 287;
	{8'd218,8'd70} : s = 288;
	{8'd218,8'd71} : s = 289;
	{8'd218,8'd72} : s = 290;
	{8'd218,8'd73} : s = 291;
	{8'd218,8'd74} : s = 292;
	{8'd218,8'd75} : s = 293;
	{8'd218,8'd76} : s = 294;
	{8'd218,8'd77} : s = 295;
	{8'd218,8'd78} : s = 296;
	{8'd218,8'd79} : s = 297;
	{8'd218,8'd80} : s = 298;
	{8'd218,8'd81} : s = 299;
	{8'd218,8'd82} : s = 300;
	{8'd218,8'd83} : s = 301;
	{8'd218,8'd84} : s = 302;
	{8'd218,8'd85} : s = 303;
	{8'd218,8'd86} : s = 304;
	{8'd218,8'd87} : s = 305;
	{8'd218,8'd88} : s = 306;
	{8'd218,8'd89} : s = 307;
	{8'd218,8'd90} : s = 308;
	{8'd218,8'd91} : s = 309;
	{8'd218,8'd92} : s = 310;
	{8'd218,8'd93} : s = 311;
	{8'd218,8'd94} : s = 312;
	{8'd218,8'd95} : s = 313;
	{8'd218,8'd96} : s = 314;
	{8'd218,8'd97} : s = 315;
	{8'd218,8'd98} : s = 316;
	{8'd218,8'd99} : s = 317;
	{8'd218,8'd100} : s = 318;
	{8'd218,8'd101} : s = 319;
	{8'd218,8'd102} : s = 320;
	{8'd218,8'd103} : s = 321;
	{8'd218,8'd104} : s = 322;
	{8'd218,8'd105} : s = 323;
	{8'd218,8'd106} : s = 324;
	{8'd218,8'd107} : s = 325;
	{8'd218,8'd108} : s = 326;
	{8'd218,8'd109} : s = 327;
	{8'd218,8'd110} : s = 328;
	{8'd218,8'd111} : s = 329;
	{8'd218,8'd112} : s = 330;
	{8'd218,8'd113} : s = 331;
	{8'd218,8'd114} : s = 332;
	{8'd218,8'd115} : s = 333;
	{8'd218,8'd116} : s = 334;
	{8'd218,8'd117} : s = 335;
	{8'd218,8'd118} : s = 336;
	{8'd218,8'd119} : s = 337;
	{8'd218,8'd120} : s = 338;
	{8'd218,8'd121} : s = 339;
	{8'd218,8'd122} : s = 340;
	{8'd218,8'd123} : s = 341;
	{8'd218,8'd124} : s = 342;
	{8'd218,8'd125} : s = 343;
	{8'd218,8'd126} : s = 344;
	{8'd218,8'd127} : s = 345;
	{8'd218,8'd128} : s = 346;
	{8'd218,8'd129} : s = 347;
	{8'd218,8'd130} : s = 348;
	{8'd218,8'd131} : s = 349;
	{8'd218,8'd132} : s = 350;
	{8'd218,8'd133} : s = 351;
	{8'd218,8'd134} : s = 352;
	{8'd218,8'd135} : s = 353;
	{8'd218,8'd136} : s = 354;
	{8'd218,8'd137} : s = 355;
	{8'd218,8'd138} : s = 356;
	{8'd218,8'd139} : s = 357;
	{8'd218,8'd140} : s = 358;
	{8'd218,8'd141} : s = 359;
	{8'd218,8'd142} : s = 360;
	{8'd218,8'd143} : s = 361;
	{8'd218,8'd144} : s = 362;
	{8'd218,8'd145} : s = 363;
	{8'd218,8'd146} : s = 364;
	{8'd218,8'd147} : s = 365;
	{8'd218,8'd148} : s = 366;
	{8'd218,8'd149} : s = 367;
	{8'd218,8'd150} : s = 368;
	{8'd218,8'd151} : s = 369;
	{8'd218,8'd152} : s = 370;
	{8'd218,8'd153} : s = 371;
	{8'd218,8'd154} : s = 372;
	{8'd218,8'd155} : s = 373;
	{8'd218,8'd156} : s = 374;
	{8'd218,8'd157} : s = 375;
	{8'd218,8'd158} : s = 376;
	{8'd218,8'd159} : s = 377;
	{8'd218,8'd160} : s = 378;
	{8'd218,8'd161} : s = 379;
	{8'd218,8'd162} : s = 380;
	{8'd218,8'd163} : s = 381;
	{8'd218,8'd164} : s = 382;
	{8'd218,8'd165} : s = 383;
	{8'd218,8'd166} : s = 384;
	{8'd218,8'd167} : s = 385;
	{8'd218,8'd168} : s = 386;
	{8'd218,8'd169} : s = 387;
	{8'd218,8'd170} : s = 388;
	{8'd218,8'd171} : s = 389;
	{8'd218,8'd172} : s = 390;
	{8'd218,8'd173} : s = 391;
	{8'd218,8'd174} : s = 392;
	{8'd218,8'd175} : s = 393;
	{8'd218,8'd176} : s = 394;
	{8'd218,8'd177} : s = 395;
	{8'd218,8'd178} : s = 396;
	{8'd218,8'd179} : s = 397;
	{8'd218,8'd180} : s = 398;
	{8'd218,8'd181} : s = 399;
	{8'd218,8'd182} : s = 400;
	{8'd218,8'd183} : s = 401;
	{8'd218,8'd184} : s = 402;
	{8'd218,8'd185} : s = 403;
	{8'd218,8'd186} : s = 404;
	{8'd218,8'd187} : s = 405;
	{8'd218,8'd188} : s = 406;
	{8'd218,8'd189} : s = 407;
	{8'd218,8'd190} : s = 408;
	{8'd218,8'd191} : s = 409;
	{8'd218,8'd192} : s = 410;
	{8'd218,8'd193} : s = 411;
	{8'd218,8'd194} : s = 412;
	{8'd218,8'd195} : s = 413;
	{8'd218,8'd196} : s = 414;
	{8'd218,8'd197} : s = 415;
	{8'd218,8'd198} : s = 416;
	{8'd218,8'd199} : s = 417;
	{8'd218,8'd200} : s = 418;
	{8'd218,8'd201} : s = 419;
	{8'd218,8'd202} : s = 420;
	{8'd218,8'd203} : s = 421;
	{8'd218,8'd204} : s = 422;
	{8'd218,8'd205} : s = 423;
	{8'd218,8'd206} : s = 424;
	{8'd218,8'd207} : s = 425;
	{8'd218,8'd208} : s = 426;
	{8'd218,8'd209} : s = 427;
	{8'd218,8'd210} : s = 428;
	{8'd218,8'd211} : s = 429;
	{8'd218,8'd212} : s = 430;
	{8'd218,8'd213} : s = 431;
	{8'd218,8'd214} : s = 432;
	{8'd218,8'd215} : s = 433;
	{8'd218,8'd216} : s = 434;
	{8'd218,8'd217} : s = 435;
	{8'd218,8'd218} : s = 436;
	{8'd218,8'd219} : s = 437;
	{8'd218,8'd220} : s = 438;
	{8'd218,8'd221} : s = 439;
	{8'd218,8'd222} : s = 440;
	{8'd218,8'd223} : s = 441;
	{8'd218,8'd224} : s = 442;
	{8'd218,8'd225} : s = 443;
	{8'd218,8'd226} : s = 444;
	{8'd218,8'd227} : s = 445;
	{8'd218,8'd228} : s = 446;
	{8'd218,8'd229} : s = 447;
	{8'd218,8'd230} : s = 448;
	{8'd218,8'd231} : s = 449;
	{8'd218,8'd232} : s = 450;
	{8'd218,8'd233} : s = 451;
	{8'd218,8'd234} : s = 452;
	{8'd218,8'd235} : s = 453;
	{8'd218,8'd236} : s = 454;
	{8'd218,8'd237} : s = 455;
	{8'd218,8'd238} : s = 456;
	{8'd218,8'd239} : s = 457;
	{8'd218,8'd240} : s = 458;
	{8'd218,8'd241} : s = 459;
	{8'd218,8'd242} : s = 460;
	{8'd218,8'd243} : s = 461;
	{8'd218,8'd244} : s = 462;
	{8'd218,8'd245} : s = 463;
	{8'd218,8'd246} : s = 464;
	{8'd218,8'd247} : s = 465;
	{8'd218,8'd248} : s = 466;
	{8'd218,8'd249} : s = 467;
	{8'd218,8'd250} : s = 468;
	{8'd218,8'd251} : s = 469;
	{8'd218,8'd252} : s = 470;
	{8'd218,8'd253} : s = 471;
	{8'd218,8'd254} : s = 472;
	{8'd218,8'd255} : s = 473;
	{8'd219,8'd0} : s = 219;
	{8'd219,8'd1} : s = 220;
	{8'd219,8'd2} : s = 221;
	{8'd219,8'd3} : s = 222;
	{8'd219,8'd4} : s = 223;
	{8'd219,8'd5} : s = 224;
	{8'd219,8'd6} : s = 225;
	{8'd219,8'd7} : s = 226;
	{8'd219,8'd8} : s = 227;
	{8'd219,8'd9} : s = 228;
	{8'd219,8'd10} : s = 229;
	{8'd219,8'd11} : s = 230;
	{8'd219,8'd12} : s = 231;
	{8'd219,8'd13} : s = 232;
	{8'd219,8'd14} : s = 233;
	{8'd219,8'd15} : s = 234;
	{8'd219,8'd16} : s = 235;
	{8'd219,8'd17} : s = 236;
	{8'd219,8'd18} : s = 237;
	{8'd219,8'd19} : s = 238;
	{8'd219,8'd20} : s = 239;
	{8'd219,8'd21} : s = 240;
	{8'd219,8'd22} : s = 241;
	{8'd219,8'd23} : s = 242;
	{8'd219,8'd24} : s = 243;
	{8'd219,8'd25} : s = 244;
	{8'd219,8'd26} : s = 245;
	{8'd219,8'd27} : s = 246;
	{8'd219,8'd28} : s = 247;
	{8'd219,8'd29} : s = 248;
	{8'd219,8'd30} : s = 249;
	{8'd219,8'd31} : s = 250;
	{8'd219,8'd32} : s = 251;
	{8'd219,8'd33} : s = 252;
	{8'd219,8'd34} : s = 253;
	{8'd219,8'd35} : s = 254;
	{8'd219,8'd36} : s = 255;
	{8'd219,8'd37} : s = 256;
	{8'd219,8'd38} : s = 257;
	{8'd219,8'd39} : s = 258;
	{8'd219,8'd40} : s = 259;
	{8'd219,8'd41} : s = 260;
	{8'd219,8'd42} : s = 261;
	{8'd219,8'd43} : s = 262;
	{8'd219,8'd44} : s = 263;
	{8'd219,8'd45} : s = 264;
	{8'd219,8'd46} : s = 265;
	{8'd219,8'd47} : s = 266;
	{8'd219,8'd48} : s = 267;
	{8'd219,8'd49} : s = 268;
	{8'd219,8'd50} : s = 269;
	{8'd219,8'd51} : s = 270;
	{8'd219,8'd52} : s = 271;
	{8'd219,8'd53} : s = 272;
	{8'd219,8'd54} : s = 273;
	{8'd219,8'd55} : s = 274;
	{8'd219,8'd56} : s = 275;
	{8'd219,8'd57} : s = 276;
	{8'd219,8'd58} : s = 277;
	{8'd219,8'd59} : s = 278;
	{8'd219,8'd60} : s = 279;
	{8'd219,8'd61} : s = 280;
	{8'd219,8'd62} : s = 281;
	{8'd219,8'd63} : s = 282;
	{8'd219,8'd64} : s = 283;
	{8'd219,8'd65} : s = 284;
	{8'd219,8'd66} : s = 285;
	{8'd219,8'd67} : s = 286;
	{8'd219,8'd68} : s = 287;
	{8'd219,8'd69} : s = 288;
	{8'd219,8'd70} : s = 289;
	{8'd219,8'd71} : s = 290;
	{8'd219,8'd72} : s = 291;
	{8'd219,8'd73} : s = 292;
	{8'd219,8'd74} : s = 293;
	{8'd219,8'd75} : s = 294;
	{8'd219,8'd76} : s = 295;
	{8'd219,8'd77} : s = 296;
	{8'd219,8'd78} : s = 297;
	{8'd219,8'd79} : s = 298;
	{8'd219,8'd80} : s = 299;
	{8'd219,8'd81} : s = 300;
	{8'd219,8'd82} : s = 301;
	{8'd219,8'd83} : s = 302;
	{8'd219,8'd84} : s = 303;
	{8'd219,8'd85} : s = 304;
	{8'd219,8'd86} : s = 305;
	{8'd219,8'd87} : s = 306;
	{8'd219,8'd88} : s = 307;
	{8'd219,8'd89} : s = 308;
	{8'd219,8'd90} : s = 309;
	{8'd219,8'd91} : s = 310;
	{8'd219,8'd92} : s = 311;
	{8'd219,8'd93} : s = 312;
	{8'd219,8'd94} : s = 313;
	{8'd219,8'd95} : s = 314;
	{8'd219,8'd96} : s = 315;
	{8'd219,8'd97} : s = 316;
	{8'd219,8'd98} : s = 317;
	{8'd219,8'd99} : s = 318;
	{8'd219,8'd100} : s = 319;
	{8'd219,8'd101} : s = 320;
	{8'd219,8'd102} : s = 321;
	{8'd219,8'd103} : s = 322;
	{8'd219,8'd104} : s = 323;
	{8'd219,8'd105} : s = 324;
	{8'd219,8'd106} : s = 325;
	{8'd219,8'd107} : s = 326;
	{8'd219,8'd108} : s = 327;
	{8'd219,8'd109} : s = 328;
	{8'd219,8'd110} : s = 329;
	{8'd219,8'd111} : s = 330;
	{8'd219,8'd112} : s = 331;
	{8'd219,8'd113} : s = 332;
	{8'd219,8'd114} : s = 333;
	{8'd219,8'd115} : s = 334;
	{8'd219,8'd116} : s = 335;
	{8'd219,8'd117} : s = 336;
	{8'd219,8'd118} : s = 337;
	{8'd219,8'd119} : s = 338;
	{8'd219,8'd120} : s = 339;
	{8'd219,8'd121} : s = 340;
	{8'd219,8'd122} : s = 341;
	{8'd219,8'd123} : s = 342;
	{8'd219,8'd124} : s = 343;
	{8'd219,8'd125} : s = 344;
	{8'd219,8'd126} : s = 345;
	{8'd219,8'd127} : s = 346;
	{8'd219,8'd128} : s = 347;
	{8'd219,8'd129} : s = 348;
	{8'd219,8'd130} : s = 349;
	{8'd219,8'd131} : s = 350;
	{8'd219,8'd132} : s = 351;
	{8'd219,8'd133} : s = 352;
	{8'd219,8'd134} : s = 353;
	{8'd219,8'd135} : s = 354;
	{8'd219,8'd136} : s = 355;
	{8'd219,8'd137} : s = 356;
	{8'd219,8'd138} : s = 357;
	{8'd219,8'd139} : s = 358;
	{8'd219,8'd140} : s = 359;
	{8'd219,8'd141} : s = 360;
	{8'd219,8'd142} : s = 361;
	{8'd219,8'd143} : s = 362;
	{8'd219,8'd144} : s = 363;
	{8'd219,8'd145} : s = 364;
	{8'd219,8'd146} : s = 365;
	{8'd219,8'd147} : s = 366;
	{8'd219,8'd148} : s = 367;
	{8'd219,8'd149} : s = 368;
	{8'd219,8'd150} : s = 369;
	{8'd219,8'd151} : s = 370;
	{8'd219,8'd152} : s = 371;
	{8'd219,8'd153} : s = 372;
	{8'd219,8'd154} : s = 373;
	{8'd219,8'd155} : s = 374;
	{8'd219,8'd156} : s = 375;
	{8'd219,8'd157} : s = 376;
	{8'd219,8'd158} : s = 377;
	{8'd219,8'd159} : s = 378;
	{8'd219,8'd160} : s = 379;
	{8'd219,8'd161} : s = 380;
	{8'd219,8'd162} : s = 381;
	{8'd219,8'd163} : s = 382;
	{8'd219,8'd164} : s = 383;
	{8'd219,8'd165} : s = 384;
	{8'd219,8'd166} : s = 385;
	{8'd219,8'd167} : s = 386;
	{8'd219,8'd168} : s = 387;
	{8'd219,8'd169} : s = 388;
	{8'd219,8'd170} : s = 389;
	{8'd219,8'd171} : s = 390;
	{8'd219,8'd172} : s = 391;
	{8'd219,8'd173} : s = 392;
	{8'd219,8'd174} : s = 393;
	{8'd219,8'd175} : s = 394;
	{8'd219,8'd176} : s = 395;
	{8'd219,8'd177} : s = 396;
	{8'd219,8'd178} : s = 397;
	{8'd219,8'd179} : s = 398;
	{8'd219,8'd180} : s = 399;
	{8'd219,8'd181} : s = 400;
	{8'd219,8'd182} : s = 401;
	{8'd219,8'd183} : s = 402;
	{8'd219,8'd184} : s = 403;
	{8'd219,8'd185} : s = 404;
	{8'd219,8'd186} : s = 405;
	{8'd219,8'd187} : s = 406;
	{8'd219,8'd188} : s = 407;
	{8'd219,8'd189} : s = 408;
	{8'd219,8'd190} : s = 409;
	{8'd219,8'd191} : s = 410;
	{8'd219,8'd192} : s = 411;
	{8'd219,8'd193} : s = 412;
	{8'd219,8'd194} : s = 413;
	{8'd219,8'd195} : s = 414;
	{8'd219,8'd196} : s = 415;
	{8'd219,8'd197} : s = 416;
	{8'd219,8'd198} : s = 417;
	{8'd219,8'd199} : s = 418;
	{8'd219,8'd200} : s = 419;
	{8'd219,8'd201} : s = 420;
	{8'd219,8'd202} : s = 421;
	{8'd219,8'd203} : s = 422;
	{8'd219,8'd204} : s = 423;
	{8'd219,8'd205} : s = 424;
	{8'd219,8'd206} : s = 425;
	{8'd219,8'd207} : s = 426;
	{8'd219,8'd208} : s = 427;
	{8'd219,8'd209} : s = 428;
	{8'd219,8'd210} : s = 429;
	{8'd219,8'd211} : s = 430;
	{8'd219,8'd212} : s = 431;
	{8'd219,8'd213} : s = 432;
	{8'd219,8'd214} : s = 433;
	{8'd219,8'd215} : s = 434;
	{8'd219,8'd216} : s = 435;
	{8'd219,8'd217} : s = 436;
	{8'd219,8'd218} : s = 437;
	{8'd219,8'd219} : s = 438;
	{8'd219,8'd220} : s = 439;
	{8'd219,8'd221} : s = 440;
	{8'd219,8'd222} : s = 441;
	{8'd219,8'd223} : s = 442;
	{8'd219,8'd224} : s = 443;
	{8'd219,8'd225} : s = 444;
	{8'd219,8'd226} : s = 445;
	{8'd219,8'd227} : s = 446;
	{8'd219,8'd228} : s = 447;
	{8'd219,8'd229} : s = 448;
	{8'd219,8'd230} : s = 449;
	{8'd219,8'd231} : s = 450;
	{8'd219,8'd232} : s = 451;
	{8'd219,8'd233} : s = 452;
	{8'd219,8'd234} : s = 453;
	{8'd219,8'd235} : s = 454;
	{8'd219,8'd236} : s = 455;
	{8'd219,8'd237} : s = 456;
	{8'd219,8'd238} : s = 457;
	{8'd219,8'd239} : s = 458;
	{8'd219,8'd240} : s = 459;
	{8'd219,8'd241} : s = 460;
	{8'd219,8'd242} : s = 461;
	{8'd219,8'd243} : s = 462;
	{8'd219,8'd244} : s = 463;
	{8'd219,8'd245} : s = 464;
	{8'd219,8'd246} : s = 465;
	{8'd219,8'd247} : s = 466;
	{8'd219,8'd248} : s = 467;
	{8'd219,8'd249} : s = 468;
	{8'd219,8'd250} : s = 469;
	{8'd219,8'd251} : s = 470;
	{8'd219,8'd252} : s = 471;
	{8'd219,8'd253} : s = 472;
	{8'd219,8'd254} : s = 473;
	{8'd219,8'd255} : s = 474;
	{8'd220,8'd0} : s = 220;
	{8'd220,8'd1} : s = 221;
	{8'd220,8'd2} : s = 222;
	{8'd220,8'd3} : s = 223;
	{8'd220,8'd4} : s = 224;
	{8'd220,8'd5} : s = 225;
	{8'd220,8'd6} : s = 226;
	{8'd220,8'd7} : s = 227;
	{8'd220,8'd8} : s = 228;
	{8'd220,8'd9} : s = 229;
	{8'd220,8'd10} : s = 230;
	{8'd220,8'd11} : s = 231;
	{8'd220,8'd12} : s = 232;
	{8'd220,8'd13} : s = 233;
	{8'd220,8'd14} : s = 234;
	{8'd220,8'd15} : s = 235;
	{8'd220,8'd16} : s = 236;
	{8'd220,8'd17} : s = 237;
	{8'd220,8'd18} : s = 238;
	{8'd220,8'd19} : s = 239;
	{8'd220,8'd20} : s = 240;
	{8'd220,8'd21} : s = 241;
	{8'd220,8'd22} : s = 242;
	{8'd220,8'd23} : s = 243;
	{8'd220,8'd24} : s = 244;
	{8'd220,8'd25} : s = 245;
	{8'd220,8'd26} : s = 246;
	{8'd220,8'd27} : s = 247;
	{8'd220,8'd28} : s = 248;
	{8'd220,8'd29} : s = 249;
	{8'd220,8'd30} : s = 250;
	{8'd220,8'd31} : s = 251;
	{8'd220,8'd32} : s = 252;
	{8'd220,8'd33} : s = 253;
	{8'd220,8'd34} : s = 254;
	{8'd220,8'd35} : s = 255;
	{8'd220,8'd36} : s = 256;
	{8'd220,8'd37} : s = 257;
	{8'd220,8'd38} : s = 258;
	{8'd220,8'd39} : s = 259;
	{8'd220,8'd40} : s = 260;
	{8'd220,8'd41} : s = 261;
	{8'd220,8'd42} : s = 262;
	{8'd220,8'd43} : s = 263;
	{8'd220,8'd44} : s = 264;
	{8'd220,8'd45} : s = 265;
	{8'd220,8'd46} : s = 266;
	{8'd220,8'd47} : s = 267;
	{8'd220,8'd48} : s = 268;
	{8'd220,8'd49} : s = 269;
	{8'd220,8'd50} : s = 270;
	{8'd220,8'd51} : s = 271;
	{8'd220,8'd52} : s = 272;
	{8'd220,8'd53} : s = 273;
	{8'd220,8'd54} : s = 274;
	{8'd220,8'd55} : s = 275;
	{8'd220,8'd56} : s = 276;
	{8'd220,8'd57} : s = 277;
	{8'd220,8'd58} : s = 278;
	{8'd220,8'd59} : s = 279;
	{8'd220,8'd60} : s = 280;
	{8'd220,8'd61} : s = 281;
	{8'd220,8'd62} : s = 282;
	{8'd220,8'd63} : s = 283;
	{8'd220,8'd64} : s = 284;
	{8'd220,8'd65} : s = 285;
	{8'd220,8'd66} : s = 286;
	{8'd220,8'd67} : s = 287;
	{8'd220,8'd68} : s = 288;
	{8'd220,8'd69} : s = 289;
	{8'd220,8'd70} : s = 290;
	{8'd220,8'd71} : s = 291;
	{8'd220,8'd72} : s = 292;
	{8'd220,8'd73} : s = 293;
	{8'd220,8'd74} : s = 294;
	{8'd220,8'd75} : s = 295;
	{8'd220,8'd76} : s = 296;
	{8'd220,8'd77} : s = 297;
	{8'd220,8'd78} : s = 298;
	{8'd220,8'd79} : s = 299;
	{8'd220,8'd80} : s = 300;
	{8'd220,8'd81} : s = 301;
	{8'd220,8'd82} : s = 302;
	{8'd220,8'd83} : s = 303;
	{8'd220,8'd84} : s = 304;
	{8'd220,8'd85} : s = 305;
	{8'd220,8'd86} : s = 306;
	{8'd220,8'd87} : s = 307;
	{8'd220,8'd88} : s = 308;
	{8'd220,8'd89} : s = 309;
	{8'd220,8'd90} : s = 310;
	{8'd220,8'd91} : s = 311;
	{8'd220,8'd92} : s = 312;
	{8'd220,8'd93} : s = 313;
	{8'd220,8'd94} : s = 314;
	{8'd220,8'd95} : s = 315;
	{8'd220,8'd96} : s = 316;
	{8'd220,8'd97} : s = 317;
	{8'd220,8'd98} : s = 318;
	{8'd220,8'd99} : s = 319;
	{8'd220,8'd100} : s = 320;
	{8'd220,8'd101} : s = 321;
	{8'd220,8'd102} : s = 322;
	{8'd220,8'd103} : s = 323;
	{8'd220,8'd104} : s = 324;
	{8'd220,8'd105} : s = 325;
	{8'd220,8'd106} : s = 326;
	{8'd220,8'd107} : s = 327;
	{8'd220,8'd108} : s = 328;
	{8'd220,8'd109} : s = 329;
	{8'd220,8'd110} : s = 330;
	{8'd220,8'd111} : s = 331;
	{8'd220,8'd112} : s = 332;
	{8'd220,8'd113} : s = 333;
	{8'd220,8'd114} : s = 334;
	{8'd220,8'd115} : s = 335;
	{8'd220,8'd116} : s = 336;
	{8'd220,8'd117} : s = 337;
	{8'd220,8'd118} : s = 338;
	{8'd220,8'd119} : s = 339;
	{8'd220,8'd120} : s = 340;
	{8'd220,8'd121} : s = 341;
	{8'd220,8'd122} : s = 342;
	{8'd220,8'd123} : s = 343;
	{8'd220,8'd124} : s = 344;
	{8'd220,8'd125} : s = 345;
	{8'd220,8'd126} : s = 346;
	{8'd220,8'd127} : s = 347;
	{8'd220,8'd128} : s = 348;
	{8'd220,8'd129} : s = 349;
	{8'd220,8'd130} : s = 350;
	{8'd220,8'd131} : s = 351;
	{8'd220,8'd132} : s = 352;
	{8'd220,8'd133} : s = 353;
	{8'd220,8'd134} : s = 354;
	{8'd220,8'd135} : s = 355;
	{8'd220,8'd136} : s = 356;
	{8'd220,8'd137} : s = 357;
	{8'd220,8'd138} : s = 358;
	{8'd220,8'd139} : s = 359;
	{8'd220,8'd140} : s = 360;
	{8'd220,8'd141} : s = 361;
	{8'd220,8'd142} : s = 362;
	{8'd220,8'd143} : s = 363;
	{8'd220,8'd144} : s = 364;
	{8'd220,8'd145} : s = 365;
	{8'd220,8'd146} : s = 366;
	{8'd220,8'd147} : s = 367;
	{8'd220,8'd148} : s = 368;
	{8'd220,8'd149} : s = 369;
	{8'd220,8'd150} : s = 370;
	{8'd220,8'd151} : s = 371;
	{8'd220,8'd152} : s = 372;
	{8'd220,8'd153} : s = 373;
	{8'd220,8'd154} : s = 374;
	{8'd220,8'd155} : s = 375;
	{8'd220,8'd156} : s = 376;
	{8'd220,8'd157} : s = 377;
	{8'd220,8'd158} : s = 378;
	{8'd220,8'd159} : s = 379;
	{8'd220,8'd160} : s = 380;
	{8'd220,8'd161} : s = 381;
	{8'd220,8'd162} : s = 382;
	{8'd220,8'd163} : s = 383;
	{8'd220,8'd164} : s = 384;
	{8'd220,8'd165} : s = 385;
	{8'd220,8'd166} : s = 386;
	{8'd220,8'd167} : s = 387;
	{8'd220,8'd168} : s = 388;
	{8'd220,8'd169} : s = 389;
	{8'd220,8'd170} : s = 390;
	{8'd220,8'd171} : s = 391;
	{8'd220,8'd172} : s = 392;
	{8'd220,8'd173} : s = 393;
	{8'd220,8'd174} : s = 394;
	{8'd220,8'd175} : s = 395;
	{8'd220,8'd176} : s = 396;
	{8'd220,8'd177} : s = 397;
	{8'd220,8'd178} : s = 398;
	{8'd220,8'd179} : s = 399;
	{8'd220,8'd180} : s = 400;
	{8'd220,8'd181} : s = 401;
	{8'd220,8'd182} : s = 402;
	{8'd220,8'd183} : s = 403;
	{8'd220,8'd184} : s = 404;
	{8'd220,8'd185} : s = 405;
	{8'd220,8'd186} : s = 406;
	{8'd220,8'd187} : s = 407;
	{8'd220,8'd188} : s = 408;
	{8'd220,8'd189} : s = 409;
	{8'd220,8'd190} : s = 410;
	{8'd220,8'd191} : s = 411;
	{8'd220,8'd192} : s = 412;
	{8'd220,8'd193} : s = 413;
	{8'd220,8'd194} : s = 414;
	{8'd220,8'd195} : s = 415;
	{8'd220,8'd196} : s = 416;
	{8'd220,8'd197} : s = 417;
	{8'd220,8'd198} : s = 418;
	{8'd220,8'd199} : s = 419;
	{8'd220,8'd200} : s = 420;
	{8'd220,8'd201} : s = 421;
	{8'd220,8'd202} : s = 422;
	{8'd220,8'd203} : s = 423;
	{8'd220,8'd204} : s = 424;
	{8'd220,8'd205} : s = 425;
	{8'd220,8'd206} : s = 426;
	{8'd220,8'd207} : s = 427;
	{8'd220,8'd208} : s = 428;
	{8'd220,8'd209} : s = 429;
	{8'd220,8'd210} : s = 430;
	{8'd220,8'd211} : s = 431;
	{8'd220,8'd212} : s = 432;
	{8'd220,8'd213} : s = 433;
	{8'd220,8'd214} : s = 434;
	{8'd220,8'd215} : s = 435;
	{8'd220,8'd216} : s = 436;
	{8'd220,8'd217} : s = 437;
	{8'd220,8'd218} : s = 438;
	{8'd220,8'd219} : s = 439;
	{8'd220,8'd220} : s = 440;
	{8'd220,8'd221} : s = 441;
	{8'd220,8'd222} : s = 442;
	{8'd220,8'd223} : s = 443;
	{8'd220,8'd224} : s = 444;
	{8'd220,8'd225} : s = 445;
	{8'd220,8'd226} : s = 446;
	{8'd220,8'd227} : s = 447;
	{8'd220,8'd228} : s = 448;
	{8'd220,8'd229} : s = 449;
	{8'd220,8'd230} : s = 450;
	{8'd220,8'd231} : s = 451;
	{8'd220,8'd232} : s = 452;
	{8'd220,8'd233} : s = 453;
	{8'd220,8'd234} : s = 454;
	{8'd220,8'd235} : s = 455;
	{8'd220,8'd236} : s = 456;
	{8'd220,8'd237} : s = 457;
	{8'd220,8'd238} : s = 458;
	{8'd220,8'd239} : s = 459;
	{8'd220,8'd240} : s = 460;
	{8'd220,8'd241} : s = 461;
	{8'd220,8'd242} : s = 462;
	{8'd220,8'd243} : s = 463;
	{8'd220,8'd244} : s = 464;
	{8'd220,8'd245} : s = 465;
	{8'd220,8'd246} : s = 466;
	{8'd220,8'd247} : s = 467;
	{8'd220,8'd248} : s = 468;
	{8'd220,8'd249} : s = 469;
	{8'd220,8'd250} : s = 470;
	{8'd220,8'd251} : s = 471;
	{8'd220,8'd252} : s = 472;
	{8'd220,8'd253} : s = 473;
	{8'd220,8'd254} : s = 474;
	{8'd220,8'd255} : s = 475;
	{8'd221,8'd0} : s = 221;
	{8'd221,8'd1} : s = 222;
	{8'd221,8'd2} : s = 223;
	{8'd221,8'd3} : s = 224;
	{8'd221,8'd4} : s = 225;
	{8'd221,8'd5} : s = 226;
	{8'd221,8'd6} : s = 227;
	{8'd221,8'd7} : s = 228;
	{8'd221,8'd8} : s = 229;
	{8'd221,8'd9} : s = 230;
	{8'd221,8'd10} : s = 231;
	{8'd221,8'd11} : s = 232;
	{8'd221,8'd12} : s = 233;
	{8'd221,8'd13} : s = 234;
	{8'd221,8'd14} : s = 235;
	{8'd221,8'd15} : s = 236;
	{8'd221,8'd16} : s = 237;
	{8'd221,8'd17} : s = 238;
	{8'd221,8'd18} : s = 239;
	{8'd221,8'd19} : s = 240;
	{8'd221,8'd20} : s = 241;
	{8'd221,8'd21} : s = 242;
	{8'd221,8'd22} : s = 243;
	{8'd221,8'd23} : s = 244;
	{8'd221,8'd24} : s = 245;
	{8'd221,8'd25} : s = 246;
	{8'd221,8'd26} : s = 247;
	{8'd221,8'd27} : s = 248;
	{8'd221,8'd28} : s = 249;
	{8'd221,8'd29} : s = 250;
	{8'd221,8'd30} : s = 251;
	{8'd221,8'd31} : s = 252;
	{8'd221,8'd32} : s = 253;
	{8'd221,8'd33} : s = 254;
	{8'd221,8'd34} : s = 255;
	{8'd221,8'd35} : s = 256;
	{8'd221,8'd36} : s = 257;
	{8'd221,8'd37} : s = 258;
	{8'd221,8'd38} : s = 259;
	{8'd221,8'd39} : s = 260;
	{8'd221,8'd40} : s = 261;
	{8'd221,8'd41} : s = 262;
	{8'd221,8'd42} : s = 263;
	{8'd221,8'd43} : s = 264;
	{8'd221,8'd44} : s = 265;
	{8'd221,8'd45} : s = 266;
	{8'd221,8'd46} : s = 267;
	{8'd221,8'd47} : s = 268;
	{8'd221,8'd48} : s = 269;
	{8'd221,8'd49} : s = 270;
	{8'd221,8'd50} : s = 271;
	{8'd221,8'd51} : s = 272;
	{8'd221,8'd52} : s = 273;
	{8'd221,8'd53} : s = 274;
	{8'd221,8'd54} : s = 275;
	{8'd221,8'd55} : s = 276;
	{8'd221,8'd56} : s = 277;
	{8'd221,8'd57} : s = 278;
	{8'd221,8'd58} : s = 279;
	{8'd221,8'd59} : s = 280;
	{8'd221,8'd60} : s = 281;
	{8'd221,8'd61} : s = 282;
	{8'd221,8'd62} : s = 283;
	{8'd221,8'd63} : s = 284;
	{8'd221,8'd64} : s = 285;
	{8'd221,8'd65} : s = 286;
	{8'd221,8'd66} : s = 287;
	{8'd221,8'd67} : s = 288;
	{8'd221,8'd68} : s = 289;
	{8'd221,8'd69} : s = 290;
	{8'd221,8'd70} : s = 291;
	{8'd221,8'd71} : s = 292;
	{8'd221,8'd72} : s = 293;
	{8'd221,8'd73} : s = 294;
	{8'd221,8'd74} : s = 295;
	{8'd221,8'd75} : s = 296;
	{8'd221,8'd76} : s = 297;
	{8'd221,8'd77} : s = 298;
	{8'd221,8'd78} : s = 299;
	{8'd221,8'd79} : s = 300;
	{8'd221,8'd80} : s = 301;
	{8'd221,8'd81} : s = 302;
	{8'd221,8'd82} : s = 303;
	{8'd221,8'd83} : s = 304;
	{8'd221,8'd84} : s = 305;
	{8'd221,8'd85} : s = 306;
	{8'd221,8'd86} : s = 307;
	{8'd221,8'd87} : s = 308;
	{8'd221,8'd88} : s = 309;
	{8'd221,8'd89} : s = 310;
	{8'd221,8'd90} : s = 311;
	{8'd221,8'd91} : s = 312;
	{8'd221,8'd92} : s = 313;
	{8'd221,8'd93} : s = 314;
	{8'd221,8'd94} : s = 315;
	{8'd221,8'd95} : s = 316;
	{8'd221,8'd96} : s = 317;
	{8'd221,8'd97} : s = 318;
	{8'd221,8'd98} : s = 319;
	{8'd221,8'd99} : s = 320;
	{8'd221,8'd100} : s = 321;
	{8'd221,8'd101} : s = 322;
	{8'd221,8'd102} : s = 323;
	{8'd221,8'd103} : s = 324;
	{8'd221,8'd104} : s = 325;
	{8'd221,8'd105} : s = 326;
	{8'd221,8'd106} : s = 327;
	{8'd221,8'd107} : s = 328;
	{8'd221,8'd108} : s = 329;
	{8'd221,8'd109} : s = 330;
	{8'd221,8'd110} : s = 331;
	{8'd221,8'd111} : s = 332;
	{8'd221,8'd112} : s = 333;
	{8'd221,8'd113} : s = 334;
	{8'd221,8'd114} : s = 335;
	{8'd221,8'd115} : s = 336;
	{8'd221,8'd116} : s = 337;
	{8'd221,8'd117} : s = 338;
	{8'd221,8'd118} : s = 339;
	{8'd221,8'd119} : s = 340;
	{8'd221,8'd120} : s = 341;
	{8'd221,8'd121} : s = 342;
	{8'd221,8'd122} : s = 343;
	{8'd221,8'd123} : s = 344;
	{8'd221,8'd124} : s = 345;
	{8'd221,8'd125} : s = 346;
	{8'd221,8'd126} : s = 347;
	{8'd221,8'd127} : s = 348;
	{8'd221,8'd128} : s = 349;
	{8'd221,8'd129} : s = 350;
	{8'd221,8'd130} : s = 351;
	{8'd221,8'd131} : s = 352;
	{8'd221,8'd132} : s = 353;
	{8'd221,8'd133} : s = 354;
	{8'd221,8'd134} : s = 355;
	{8'd221,8'd135} : s = 356;
	{8'd221,8'd136} : s = 357;
	{8'd221,8'd137} : s = 358;
	{8'd221,8'd138} : s = 359;
	{8'd221,8'd139} : s = 360;
	{8'd221,8'd140} : s = 361;
	{8'd221,8'd141} : s = 362;
	{8'd221,8'd142} : s = 363;
	{8'd221,8'd143} : s = 364;
	{8'd221,8'd144} : s = 365;
	{8'd221,8'd145} : s = 366;
	{8'd221,8'd146} : s = 367;
	{8'd221,8'd147} : s = 368;
	{8'd221,8'd148} : s = 369;
	{8'd221,8'd149} : s = 370;
	{8'd221,8'd150} : s = 371;
	{8'd221,8'd151} : s = 372;
	{8'd221,8'd152} : s = 373;
	{8'd221,8'd153} : s = 374;
	{8'd221,8'd154} : s = 375;
	{8'd221,8'd155} : s = 376;
	{8'd221,8'd156} : s = 377;
	{8'd221,8'd157} : s = 378;
	{8'd221,8'd158} : s = 379;
	{8'd221,8'd159} : s = 380;
	{8'd221,8'd160} : s = 381;
	{8'd221,8'd161} : s = 382;
	{8'd221,8'd162} : s = 383;
	{8'd221,8'd163} : s = 384;
	{8'd221,8'd164} : s = 385;
	{8'd221,8'd165} : s = 386;
	{8'd221,8'd166} : s = 387;
	{8'd221,8'd167} : s = 388;
	{8'd221,8'd168} : s = 389;
	{8'd221,8'd169} : s = 390;
	{8'd221,8'd170} : s = 391;
	{8'd221,8'd171} : s = 392;
	{8'd221,8'd172} : s = 393;
	{8'd221,8'd173} : s = 394;
	{8'd221,8'd174} : s = 395;
	{8'd221,8'd175} : s = 396;
	{8'd221,8'd176} : s = 397;
	{8'd221,8'd177} : s = 398;
	{8'd221,8'd178} : s = 399;
	{8'd221,8'd179} : s = 400;
	{8'd221,8'd180} : s = 401;
	{8'd221,8'd181} : s = 402;
	{8'd221,8'd182} : s = 403;
	{8'd221,8'd183} : s = 404;
	{8'd221,8'd184} : s = 405;
	{8'd221,8'd185} : s = 406;
	{8'd221,8'd186} : s = 407;
	{8'd221,8'd187} : s = 408;
	{8'd221,8'd188} : s = 409;
	{8'd221,8'd189} : s = 410;
	{8'd221,8'd190} : s = 411;
	{8'd221,8'd191} : s = 412;
	{8'd221,8'd192} : s = 413;
	{8'd221,8'd193} : s = 414;
	{8'd221,8'd194} : s = 415;
	{8'd221,8'd195} : s = 416;
	{8'd221,8'd196} : s = 417;
	{8'd221,8'd197} : s = 418;
	{8'd221,8'd198} : s = 419;
	{8'd221,8'd199} : s = 420;
	{8'd221,8'd200} : s = 421;
	{8'd221,8'd201} : s = 422;
	{8'd221,8'd202} : s = 423;
	{8'd221,8'd203} : s = 424;
	{8'd221,8'd204} : s = 425;
	{8'd221,8'd205} : s = 426;
	{8'd221,8'd206} : s = 427;
	{8'd221,8'd207} : s = 428;
	{8'd221,8'd208} : s = 429;
	{8'd221,8'd209} : s = 430;
	{8'd221,8'd210} : s = 431;
	{8'd221,8'd211} : s = 432;
	{8'd221,8'd212} : s = 433;
	{8'd221,8'd213} : s = 434;
	{8'd221,8'd214} : s = 435;
	{8'd221,8'd215} : s = 436;
	{8'd221,8'd216} : s = 437;
	{8'd221,8'd217} : s = 438;
	{8'd221,8'd218} : s = 439;
	{8'd221,8'd219} : s = 440;
	{8'd221,8'd220} : s = 441;
	{8'd221,8'd221} : s = 442;
	{8'd221,8'd222} : s = 443;
	{8'd221,8'd223} : s = 444;
	{8'd221,8'd224} : s = 445;
	{8'd221,8'd225} : s = 446;
	{8'd221,8'd226} : s = 447;
	{8'd221,8'd227} : s = 448;
	{8'd221,8'd228} : s = 449;
	{8'd221,8'd229} : s = 450;
	{8'd221,8'd230} : s = 451;
	{8'd221,8'd231} : s = 452;
	{8'd221,8'd232} : s = 453;
	{8'd221,8'd233} : s = 454;
	{8'd221,8'd234} : s = 455;
	{8'd221,8'd235} : s = 456;
	{8'd221,8'd236} : s = 457;
	{8'd221,8'd237} : s = 458;
	{8'd221,8'd238} : s = 459;
	{8'd221,8'd239} : s = 460;
	{8'd221,8'd240} : s = 461;
	{8'd221,8'd241} : s = 462;
	{8'd221,8'd242} : s = 463;
	{8'd221,8'd243} : s = 464;
	{8'd221,8'd244} : s = 465;
	{8'd221,8'd245} : s = 466;
	{8'd221,8'd246} : s = 467;
	{8'd221,8'd247} : s = 468;
	{8'd221,8'd248} : s = 469;
	{8'd221,8'd249} : s = 470;
	{8'd221,8'd250} : s = 471;
	{8'd221,8'd251} : s = 472;
	{8'd221,8'd252} : s = 473;
	{8'd221,8'd253} : s = 474;
	{8'd221,8'd254} : s = 475;
	{8'd221,8'd255} : s = 476;
	{8'd222,8'd0} : s = 222;
	{8'd222,8'd1} : s = 223;
	{8'd222,8'd2} : s = 224;
	{8'd222,8'd3} : s = 225;
	{8'd222,8'd4} : s = 226;
	{8'd222,8'd5} : s = 227;
	{8'd222,8'd6} : s = 228;
	{8'd222,8'd7} : s = 229;
	{8'd222,8'd8} : s = 230;
	{8'd222,8'd9} : s = 231;
	{8'd222,8'd10} : s = 232;
	{8'd222,8'd11} : s = 233;
	{8'd222,8'd12} : s = 234;
	{8'd222,8'd13} : s = 235;
	{8'd222,8'd14} : s = 236;
	{8'd222,8'd15} : s = 237;
	{8'd222,8'd16} : s = 238;
	{8'd222,8'd17} : s = 239;
	{8'd222,8'd18} : s = 240;
	{8'd222,8'd19} : s = 241;
	{8'd222,8'd20} : s = 242;
	{8'd222,8'd21} : s = 243;
	{8'd222,8'd22} : s = 244;
	{8'd222,8'd23} : s = 245;
	{8'd222,8'd24} : s = 246;
	{8'd222,8'd25} : s = 247;
	{8'd222,8'd26} : s = 248;
	{8'd222,8'd27} : s = 249;
	{8'd222,8'd28} : s = 250;
	{8'd222,8'd29} : s = 251;
	{8'd222,8'd30} : s = 252;
	{8'd222,8'd31} : s = 253;
	{8'd222,8'd32} : s = 254;
	{8'd222,8'd33} : s = 255;
	{8'd222,8'd34} : s = 256;
	{8'd222,8'd35} : s = 257;
	{8'd222,8'd36} : s = 258;
	{8'd222,8'd37} : s = 259;
	{8'd222,8'd38} : s = 260;
	{8'd222,8'd39} : s = 261;
	{8'd222,8'd40} : s = 262;
	{8'd222,8'd41} : s = 263;
	{8'd222,8'd42} : s = 264;
	{8'd222,8'd43} : s = 265;
	{8'd222,8'd44} : s = 266;
	{8'd222,8'd45} : s = 267;
	{8'd222,8'd46} : s = 268;
	{8'd222,8'd47} : s = 269;
	{8'd222,8'd48} : s = 270;
	{8'd222,8'd49} : s = 271;
	{8'd222,8'd50} : s = 272;
	{8'd222,8'd51} : s = 273;
	{8'd222,8'd52} : s = 274;
	{8'd222,8'd53} : s = 275;
	{8'd222,8'd54} : s = 276;
	{8'd222,8'd55} : s = 277;
	{8'd222,8'd56} : s = 278;
	{8'd222,8'd57} : s = 279;
	{8'd222,8'd58} : s = 280;
	{8'd222,8'd59} : s = 281;
	{8'd222,8'd60} : s = 282;
	{8'd222,8'd61} : s = 283;
	{8'd222,8'd62} : s = 284;
	{8'd222,8'd63} : s = 285;
	{8'd222,8'd64} : s = 286;
	{8'd222,8'd65} : s = 287;
	{8'd222,8'd66} : s = 288;
	{8'd222,8'd67} : s = 289;
	{8'd222,8'd68} : s = 290;
	{8'd222,8'd69} : s = 291;
	{8'd222,8'd70} : s = 292;
	{8'd222,8'd71} : s = 293;
	{8'd222,8'd72} : s = 294;
	{8'd222,8'd73} : s = 295;
	{8'd222,8'd74} : s = 296;
	{8'd222,8'd75} : s = 297;
	{8'd222,8'd76} : s = 298;
	{8'd222,8'd77} : s = 299;
	{8'd222,8'd78} : s = 300;
	{8'd222,8'd79} : s = 301;
	{8'd222,8'd80} : s = 302;
	{8'd222,8'd81} : s = 303;
	{8'd222,8'd82} : s = 304;
	{8'd222,8'd83} : s = 305;
	{8'd222,8'd84} : s = 306;
	{8'd222,8'd85} : s = 307;
	{8'd222,8'd86} : s = 308;
	{8'd222,8'd87} : s = 309;
	{8'd222,8'd88} : s = 310;
	{8'd222,8'd89} : s = 311;
	{8'd222,8'd90} : s = 312;
	{8'd222,8'd91} : s = 313;
	{8'd222,8'd92} : s = 314;
	{8'd222,8'd93} : s = 315;
	{8'd222,8'd94} : s = 316;
	{8'd222,8'd95} : s = 317;
	{8'd222,8'd96} : s = 318;
	{8'd222,8'd97} : s = 319;
	{8'd222,8'd98} : s = 320;
	{8'd222,8'd99} : s = 321;
	{8'd222,8'd100} : s = 322;
	{8'd222,8'd101} : s = 323;
	{8'd222,8'd102} : s = 324;
	{8'd222,8'd103} : s = 325;
	{8'd222,8'd104} : s = 326;
	{8'd222,8'd105} : s = 327;
	{8'd222,8'd106} : s = 328;
	{8'd222,8'd107} : s = 329;
	{8'd222,8'd108} : s = 330;
	{8'd222,8'd109} : s = 331;
	{8'd222,8'd110} : s = 332;
	{8'd222,8'd111} : s = 333;
	{8'd222,8'd112} : s = 334;
	{8'd222,8'd113} : s = 335;
	{8'd222,8'd114} : s = 336;
	{8'd222,8'd115} : s = 337;
	{8'd222,8'd116} : s = 338;
	{8'd222,8'd117} : s = 339;
	{8'd222,8'd118} : s = 340;
	{8'd222,8'd119} : s = 341;
	{8'd222,8'd120} : s = 342;
	{8'd222,8'd121} : s = 343;
	{8'd222,8'd122} : s = 344;
	{8'd222,8'd123} : s = 345;
	{8'd222,8'd124} : s = 346;
	{8'd222,8'd125} : s = 347;
	{8'd222,8'd126} : s = 348;
	{8'd222,8'd127} : s = 349;
	{8'd222,8'd128} : s = 350;
	{8'd222,8'd129} : s = 351;
	{8'd222,8'd130} : s = 352;
	{8'd222,8'd131} : s = 353;
	{8'd222,8'd132} : s = 354;
	{8'd222,8'd133} : s = 355;
	{8'd222,8'd134} : s = 356;
	{8'd222,8'd135} : s = 357;
	{8'd222,8'd136} : s = 358;
	{8'd222,8'd137} : s = 359;
	{8'd222,8'd138} : s = 360;
	{8'd222,8'd139} : s = 361;
	{8'd222,8'd140} : s = 362;
	{8'd222,8'd141} : s = 363;
	{8'd222,8'd142} : s = 364;
	{8'd222,8'd143} : s = 365;
	{8'd222,8'd144} : s = 366;
	{8'd222,8'd145} : s = 367;
	{8'd222,8'd146} : s = 368;
	{8'd222,8'd147} : s = 369;
	{8'd222,8'd148} : s = 370;
	{8'd222,8'd149} : s = 371;
	{8'd222,8'd150} : s = 372;
	{8'd222,8'd151} : s = 373;
	{8'd222,8'd152} : s = 374;
	{8'd222,8'd153} : s = 375;
	{8'd222,8'd154} : s = 376;
	{8'd222,8'd155} : s = 377;
	{8'd222,8'd156} : s = 378;
	{8'd222,8'd157} : s = 379;
	{8'd222,8'd158} : s = 380;
	{8'd222,8'd159} : s = 381;
	{8'd222,8'd160} : s = 382;
	{8'd222,8'd161} : s = 383;
	{8'd222,8'd162} : s = 384;
	{8'd222,8'd163} : s = 385;
	{8'd222,8'd164} : s = 386;
	{8'd222,8'd165} : s = 387;
	{8'd222,8'd166} : s = 388;
	{8'd222,8'd167} : s = 389;
	{8'd222,8'd168} : s = 390;
	{8'd222,8'd169} : s = 391;
	{8'd222,8'd170} : s = 392;
	{8'd222,8'd171} : s = 393;
	{8'd222,8'd172} : s = 394;
	{8'd222,8'd173} : s = 395;
	{8'd222,8'd174} : s = 396;
	{8'd222,8'd175} : s = 397;
	{8'd222,8'd176} : s = 398;
	{8'd222,8'd177} : s = 399;
	{8'd222,8'd178} : s = 400;
	{8'd222,8'd179} : s = 401;
	{8'd222,8'd180} : s = 402;
	{8'd222,8'd181} : s = 403;
	{8'd222,8'd182} : s = 404;
	{8'd222,8'd183} : s = 405;
	{8'd222,8'd184} : s = 406;
	{8'd222,8'd185} : s = 407;
	{8'd222,8'd186} : s = 408;
	{8'd222,8'd187} : s = 409;
	{8'd222,8'd188} : s = 410;
	{8'd222,8'd189} : s = 411;
	{8'd222,8'd190} : s = 412;
	{8'd222,8'd191} : s = 413;
	{8'd222,8'd192} : s = 414;
	{8'd222,8'd193} : s = 415;
	{8'd222,8'd194} : s = 416;
	{8'd222,8'd195} : s = 417;
	{8'd222,8'd196} : s = 418;
	{8'd222,8'd197} : s = 419;
	{8'd222,8'd198} : s = 420;
	{8'd222,8'd199} : s = 421;
	{8'd222,8'd200} : s = 422;
	{8'd222,8'd201} : s = 423;
	{8'd222,8'd202} : s = 424;
	{8'd222,8'd203} : s = 425;
	{8'd222,8'd204} : s = 426;
	{8'd222,8'd205} : s = 427;
	{8'd222,8'd206} : s = 428;
	{8'd222,8'd207} : s = 429;
	{8'd222,8'd208} : s = 430;
	{8'd222,8'd209} : s = 431;
	{8'd222,8'd210} : s = 432;
	{8'd222,8'd211} : s = 433;
	{8'd222,8'd212} : s = 434;
	{8'd222,8'd213} : s = 435;
	{8'd222,8'd214} : s = 436;
	{8'd222,8'd215} : s = 437;
	{8'd222,8'd216} : s = 438;
	{8'd222,8'd217} : s = 439;
	{8'd222,8'd218} : s = 440;
	{8'd222,8'd219} : s = 441;
	{8'd222,8'd220} : s = 442;
	{8'd222,8'd221} : s = 443;
	{8'd222,8'd222} : s = 444;
	{8'd222,8'd223} : s = 445;
	{8'd222,8'd224} : s = 446;
	{8'd222,8'd225} : s = 447;
	{8'd222,8'd226} : s = 448;
	{8'd222,8'd227} : s = 449;
	{8'd222,8'd228} : s = 450;
	{8'd222,8'd229} : s = 451;
	{8'd222,8'd230} : s = 452;
	{8'd222,8'd231} : s = 453;
	{8'd222,8'd232} : s = 454;
	{8'd222,8'd233} : s = 455;
	{8'd222,8'd234} : s = 456;
	{8'd222,8'd235} : s = 457;
	{8'd222,8'd236} : s = 458;
	{8'd222,8'd237} : s = 459;
	{8'd222,8'd238} : s = 460;
	{8'd222,8'd239} : s = 461;
	{8'd222,8'd240} : s = 462;
	{8'd222,8'd241} : s = 463;
	{8'd222,8'd242} : s = 464;
	{8'd222,8'd243} : s = 465;
	{8'd222,8'd244} : s = 466;
	{8'd222,8'd245} : s = 467;
	{8'd222,8'd246} : s = 468;
	{8'd222,8'd247} : s = 469;
	{8'd222,8'd248} : s = 470;
	{8'd222,8'd249} : s = 471;
	{8'd222,8'd250} : s = 472;
	{8'd222,8'd251} : s = 473;
	{8'd222,8'd252} : s = 474;
	{8'd222,8'd253} : s = 475;
	{8'd222,8'd254} : s = 476;
	{8'd222,8'd255} : s = 477;
	{8'd223,8'd0} : s = 223;
	{8'd223,8'd1} : s = 224;
	{8'd223,8'd2} : s = 225;
	{8'd223,8'd3} : s = 226;
	{8'd223,8'd4} : s = 227;
	{8'd223,8'd5} : s = 228;
	{8'd223,8'd6} : s = 229;
	{8'd223,8'd7} : s = 230;
	{8'd223,8'd8} : s = 231;
	{8'd223,8'd9} : s = 232;
	{8'd223,8'd10} : s = 233;
	{8'd223,8'd11} : s = 234;
	{8'd223,8'd12} : s = 235;
	{8'd223,8'd13} : s = 236;
	{8'd223,8'd14} : s = 237;
	{8'd223,8'd15} : s = 238;
	{8'd223,8'd16} : s = 239;
	{8'd223,8'd17} : s = 240;
	{8'd223,8'd18} : s = 241;
	{8'd223,8'd19} : s = 242;
	{8'd223,8'd20} : s = 243;
	{8'd223,8'd21} : s = 244;
	{8'd223,8'd22} : s = 245;
	{8'd223,8'd23} : s = 246;
	{8'd223,8'd24} : s = 247;
	{8'd223,8'd25} : s = 248;
	{8'd223,8'd26} : s = 249;
	{8'd223,8'd27} : s = 250;
	{8'd223,8'd28} : s = 251;
	{8'd223,8'd29} : s = 252;
	{8'd223,8'd30} : s = 253;
	{8'd223,8'd31} : s = 254;
	{8'd223,8'd32} : s = 255;
	{8'd223,8'd33} : s = 256;
	{8'd223,8'd34} : s = 257;
	{8'd223,8'd35} : s = 258;
	{8'd223,8'd36} : s = 259;
	{8'd223,8'd37} : s = 260;
	{8'd223,8'd38} : s = 261;
	{8'd223,8'd39} : s = 262;
	{8'd223,8'd40} : s = 263;
	{8'd223,8'd41} : s = 264;
	{8'd223,8'd42} : s = 265;
	{8'd223,8'd43} : s = 266;
	{8'd223,8'd44} : s = 267;
	{8'd223,8'd45} : s = 268;
	{8'd223,8'd46} : s = 269;
	{8'd223,8'd47} : s = 270;
	{8'd223,8'd48} : s = 271;
	{8'd223,8'd49} : s = 272;
	{8'd223,8'd50} : s = 273;
	{8'd223,8'd51} : s = 274;
	{8'd223,8'd52} : s = 275;
	{8'd223,8'd53} : s = 276;
	{8'd223,8'd54} : s = 277;
	{8'd223,8'd55} : s = 278;
	{8'd223,8'd56} : s = 279;
	{8'd223,8'd57} : s = 280;
	{8'd223,8'd58} : s = 281;
	{8'd223,8'd59} : s = 282;
	{8'd223,8'd60} : s = 283;
	{8'd223,8'd61} : s = 284;
	{8'd223,8'd62} : s = 285;
	{8'd223,8'd63} : s = 286;
	{8'd223,8'd64} : s = 287;
	{8'd223,8'd65} : s = 288;
	{8'd223,8'd66} : s = 289;
	{8'd223,8'd67} : s = 290;
	{8'd223,8'd68} : s = 291;
	{8'd223,8'd69} : s = 292;
	{8'd223,8'd70} : s = 293;
	{8'd223,8'd71} : s = 294;
	{8'd223,8'd72} : s = 295;
	{8'd223,8'd73} : s = 296;
	{8'd223,8'd74} : s = 297;
	{8'd223,8'd75} : s = 298;
	{8'd223,8'd76} : s = 299;
	{8'd223,8'd77} : s = 300;
	{8'd223,8'd78} : s = 301;
	{8'd223,8'd79} : s = 302;
	{8'd223,8'd80} : s = 303;
	{8'd223,8'd81} : s = 304;
	{8'd223,8'd82} : s = 305;
	{8'd223,8'd83} : s = 306;
	{8'd223,8'd84} : s = 307;
	{8'd223,8'd85} : s = 308;
	{8'd223,8'd86} : s = 309;
	{8'd223,8'd87} : s = 310;
	{8'd223,8'd88} : s = 311;
	{8'd223,8'd89} : s = 312;
	{8'd223,8'd90} : s = 313;
	{8'd223,8'd91} : s = 314;
	{8'd223,8'd92} : s = 315;
	{8'd223,8'd93} : s = 316;
	{8'd223,8'd94} : s = 317;
	{8'd223,8'd95} : s = 318;
	{8'd223,8'd96} : s = 319;
	{8'd223,8'd97} : s = 320;
	{8'd223,8'd98} : s = 321;
	{8'd223,8'd99} : s = 322;
	{8'd223,8'd100} : s = 323;
	{8'd223,8'd101} : s = 324;
	{8'd223,8'd102} : s = 325;
	{8'd223,8'd103} : s = 326;
	{8'd223,8'd104} : s = 327;
	{8'd223,8'd105} : s = 328;
	{8'd223,8'd106} : s = 329;
	{8'd223,8'd107} : s = 330;
	{8'd223,8'd108} : s = 331;
	{8'd223,8'd109} : s = 332;
	{8'd223,8'd110} : s = 333;
	{8'd223,8'd111} : s = 334;
	{8'd223,8'd112} : s = 335;
	{8'd223,8'd113} : s = 336;
	{8'd223,8'd114} : s = 337;
	{8'd223,8'd115} : s = 338;
	{8'd223,8'd116} : s = 339;
	{8'd223,8'd117} : s = 340;
	{8'd223,8'd118} : s = 341;
	{8'd223,8'd119} : s = 342;
	{8'd223,8'd120} : s = 343;
	{8'd223,8'd121} : s = 344;
	{8'd223,8'd122} : s = 345;
	{8'd223,8'd123} : s = 346;
	{8'd223,8'd124} : s = 347;
	{8'd223,8'd125} : s = 348;
	{8'd223,8'd126} : s = 349;
	{8'd223,8'd127} : s = 350;
	{8'd223,8'd128} : s = 351;
	{8'd223,8'd129} : s = 352;
	{8'd223,8'd130} : s = 353;
	{8'd223,8'd131} : s = 354;
	{8'd223,8'd132} : s = 355;
	{8'd223,8'd133} : s = 356;
	{8'd223,8'd134} : s = 357;
	{8'd223,8'd135} : s = 358;
	{8'd223,8'd136} : s = 359;
	{8'd223,8'd137} : s = 360;
	{8'd223,8'd138} : s = 361;
	{8'd223,8'd139} : s = 362;
	{8'd223,8'd140} : s = 363;
	{8'd223,8'd141} : s = 364;
	{8'd223,8'd142} : s = 365;
	{8'd223,8'd143} : s = 366;
	{8'd223,8'd144} : s = 367;
	{8'd223,8'd145} : s = 368;
	{8'd223,8'd146} : s = 369;
	{8'd223,8'd147} : s = 370;
	{8'd223,8'd148} : s = 371;
	{8'd223,8'd149} : s = 372;
	{8'd223,8'd150} : s = 373;
	{8'd223,8'd151} : s = 374;
	{8'd223,8'd152} : s = 375;
	{8'd223,8'd153} : s = 376;
	{8'd223,8'd154} : s = 377;
	{8'd223,8'd155} : s = 378;
	{8'd223,8'd156} : s = 379;
	{8'd223,8'd157} : s = 380;
	{8'd223,8'd158} : s = 381;
	{8'd223,8'd159} : s = 382;
	{8'd223,8'd160} : s = 383;
	{8'd223,8'd161} : s = 384;
	{8'd223,8'd162} : s = 385;
	{8'd223,8'd163} : s = 386;
	{8'd223,8'd164} : s = 387;
	{8'd223,8'd165} : s = 388;
	{8'd223,8'd166} : s = 389;
	{8'd223,8'd167} : s = 390;
	{8'd223,8'd168} : s = 391;
	{8'd223,8'd169} : s = 392;
	{8'd223,8'd170} : s = 393;
	{8'd223,8'd171} : s = 394;
	{8'd223,8'd172} : s = 395;
	{8'd223,8'd173} : s = 396;
	{8'd223,8'd174} : s = 397;
	{8'd223,8'd175} : s = 398;
	{8'd223,8'd176} : s = 399;
	{8'd223,8'd177} : s = 400;
	{8'd223,8'd178} : s = 401;
	{8'd223,8'd179} : s = 402;
	{8'd223,8'd180} : s = 403;
	{8'd223,8'd181} : s = 404;
	{8'd223,8'd182} : s = 405;
	{8'd223,8'd183} : s = 406;
	{8'd223,8'd184} : s = 407;
	{8'd223,8'd185} : s = 408;
	{8'd223,8'd186} : s = 409;
	{8'd223,8'd187} : s = 410;
	{8'd223,8'd188} : s = 411;
	{8'd223,8'd189} : s = 412;
	{8'd223,8'd190} : s = 413;
	{8'd223,8'd191} : s = 414;
	{8'd223,8'd192} : s = 415;
	{8'd223,8'd193} : s = 416;
	{8'd223,8'd194} : s = 417;
	{8'd223,8'd195} : s = 418;
	{8'd223,8'd196} : s = 419;
	{8'd223,8'd197} : s = 420;
	{8'd223,8'd198} : s = 421;
	{8'd223,8'd199} : s = 422;
	{8'd223,8'd200} : s = 423;
	{8'd223,8'd201} : s = 424;
	{8'd223,8'd202} : s = 425;
	{8'd223,8'd203} : s = 426;
	{8'd223,8'd204} : s = 427;
	{8'd223,8'd205} : s = 428;
	{8'd223,8'd206} : s = 429;
	{8'd223,8'd207} : s = 430;
	{8'd223,8'd208} : s = 431;
	{8'd223,8'd209} : s = 432;
	{8'd223,8'd210} : s = 433;
	{8'd223,8'd211} : s = 434;
	{8'd223,8'd212} : s = 435;
	{8'd223,8'd213} : s = 436;
	{8'd223,8'd214} : s = 437;
	{8'd223,8'd215} : s = 438;
	{8'd223,8'd216} : s = 439;
	{8'd223,8'd217} : s = 440;
	{8'd223,8'd218} : s = 441;
	{8'd223,8'd219} : s = 442;
	{8'd223,8'd220} : s = 443;
	{8'd223,8'd221} : s = 444;
	{8'd223,8'd222} : s = 445;
	{8'd223,8'd223} : s = 446;
	{8'd223,8'd224} : s = 447;
	{8'd223,8'd225} : s = 448;
	{8'd223,8'd226} : s = 449;
	{8'd223,8'd227} : s = 450;
	{8'd223,8'd228} : s = 451;
	{8'd223,8'd229} : s = 452;
	{8'd223,8'd230} : s = 453;
	{8'd223,8'd231} : s = 454;
	{8'd223,8'd232} : s = 455;
	{8'd223,8'd233} : s = 456;
	{8'd223,8'd234} : s = 457;
	{8'd223,8'd235} : s = 458;
	{8'd223,8'd236} : s = 459;
	{8'd223,8'd237} : s = 460;
	{8'd223,8'd238} : s = 461;
	{8'd223,8'd239} : s = 462;
	{8'd223,8'd240} : s = 463;
	{8'd223,8'd241} : s = 464;
	{8'd223,8'd242} : s = 465;
	{8'd223,8'd243} : s = 466;
	{8'd223,8'd244} : s = 467;
	{8'd223,8'd245} : s = 468;
	{8'd223,8'd246} : s = 469;
	{8'd223,8'd247} : s = 470;
	{8'd223,8'd248} : s = 471;
	{8'd223,8'd249} : s = 472;
	{8'd223,8'd250} : s = 473;
	{8'd223,8'd251} : s = 474;
	{8'd223,8'd252} : s = 475;
	{8'd223,8'd253} : s = 476;
	{8'd223,8'd254} : s = 477;
	{8'd223,8'd255} : s = 478;
	{8'd224,8'd0} : s = 224;
	{8'd224,8'd1} : s = 225;
	{8'd224,8'd2} : s = 226;
	{8'd224,8'd3} : s = 227;
	{8'd224,8'd4} : s = 228;
	{8'd224,8'd5} : s = 229;
	{8'd224,8'd6} : s = 230;
	{8'd224,8'd7} : s = 231;
	{8'd224,8'd8} : s = 232;
	{8'd224,8'd9} : s = 233;
	{8'd224,8'd10} : s = 234;
	{8'd224,8'd11} : s = 235;
	{8'd224,8'd12} : s = 236;
	{8'd224,8'd13} : s = 237;
	{8'd224,8'd14} : s = 238;
	{8'd224,8'd15} : s = 239;
	{8'd224,8'd16} : s = 240;
	{8'd224,8'd17} : s = 241;
	{8'd224,8'd18} : s = 242;
	{8'd224,8'd19} : s = 243;
	{8'd224,8'd20} : s = 244;
	{8'd224,8'd21} : s = 245;
	{8'd224,8'd22} : s = 246;
	{8'd224,8'd23} : s = 247;
	{8'd224,8'd24} : s = 248;
	{8'd224,8'd25} : s = 249;
	{8'd224,8'd26} : s = 250;
	{8'd224,8'd27} : s = 251;
	{8'd224,8'd28} : s = 252;
	{8'd224,8'd29} : s = 253;
	{8'd224,8'd30} : s = 254;
	{8'd224,8'd31} : s = 255;
	{8'd224,8'd32} : s = 256;
	{8'd224,8'd33} : s = 257;
	{8'd224,8'd34} : s = 258;
	{8'd224,8'd35} : s = 259;
	{8'd224,8'd36} : s = 260;
	{8'd224,8'd37} : s = 261;
	{8'd224,8'd38} : s = 262;
	{8'd224,8'd39} : s = 263;
	{8'd224,8'd40} : s = 264;
	{8'd224,8'd41} : s = 265;
	{8'd224,8'd42} : s = 266;
	{8'd224,8'd43} : s = 267;
	{8'd224,8'd44} : s = 268;
	{8'd224,8'd45} : s = 269;
	{8'd224,8'd46} : s = 270;
	{8'd224,8'd47} : s = 271;
	{8'd224,8'd48} : s = 272;
	{8'd224,8'd49} : s = 273;
	{8'd224,8'd50} : s = 274;
	{8'd224,8'd51} : s = 275;
	{8'd224,8'd52} : s = 276;
	{8'd224,8'd53} : s = 277;
	{8'd224,8'd54} : s = 278;
	{8'd224,8'd55} : s = 279;
	{8'd224,8'd56} : s = 280;
	{8'd224,8'd57} : s = 281;
	{8'd224,8'd58} : s = 282;
	{8'd224,8'd59} : s = 283;
	{8'd224,8'd60} : s = 284;
	{8'd224,8'd61} : s = 285;
	{8'd224,8'd62} : s = 286;
	{8'd224,8'd63} : s = 287;
	{8'd224,8'd64} : s = 288;
	{8'd224,8'd65} : s = 289;
	{8'd224,8'd66} : s = 290;
	{8'd224,8'd67} : s = 291;
	{8'd224,8'd68} : s = 292;
	{8'd224,8'd69} : s = 293;
	{8'd224,8'd70} : s = 294;
	{8'd224,8'd71} : s = 295;
	{8'd224,8'd72} : s = 296;
	{8'd224,8'd73} : s = 297;
	{8'd224,8'd74} : s = 298;
	{8'd224,8'd75} : s = 299;
	{8'd224,8'd76} : s = 300;
	{8'd224,8'd77} : s = 301;
	{8'd224,8'd78} : s = 302;
	{8'd224,8'd79} : s = 303;
	{8'd224,8'd80} : s = 304;
	{8'd224,8'd81} : s = 305;
	{8'd224,8'd82} : s = 306;
	{8'd224,8'd83} : s = 307;
	{8'd224,8'd84} : s = 308;
	{8'd224,8'd85} : s = 309;
	{8'd224,8'd86} : s = 310;
	{8'd224,8'd87} : s = 311;
	{8'd224,8'd88} : s = 312;
	{8'd224,8'd89} : s = 313;
	{8'd224,8'd90} : s = 314;
	{8'd224,8'd91} : s = 315;
	{8'd224,8'd92} : s = 316;
	{8'd224,8'd93} : s = 317;
	{8'd224,8'd94} : s = 318;
	{8'd224,8'd95} : s = 319;
	{8'd224,8'd96} : s = 320;
	{8'd224,8'd97} : s = 321;
	{8'd224,8'd98} : s = 322;
	{8'd224,8'd99} : s = 323;
	{8'd224,8'd100} : s = 324;
	{8'd224,8'd101} : s = 325;
	{8'd224,8'd102} : s = 326;
	{8'd224,8'd103} : s = 327;
	{8'd224,8'd104} : s = 328;
	{8'd224,8'd105} : s = 329;
	{8'd224,8'd106} : s = 330;
	{8'd224,8'd107} : s = 331;
	{8'd224,8'd108} : s = 332;
	{8'd224,8'd109} : s = 333;
	{8'd224,8'd110} : s = 334;
	{8'd224,8'd111} : s = 335;
	{8'd224,8'd112} : s = 336;
	{8'd224,8'd113} : s = 337;
	{8'd224,8'd114} : s = 338;
	{8'd224,8'd115} : s = 339;
	{8'd224,8'd116} : s = 340;
	{8'd224,8'd117} : s = 341;
	{8'd224,8'd118} : s = 342;
	{8'd224,8'd119} : s = 343;
	{8'd224,8'd120} : s = 344;
	{8'd224,8'd121} : s = 345;
	{8'd224,8'd122} : s = 346;
	{8'd224,8'd123} : s = 347;
	{8'd224,8'd124} : s = 348;
	{8'd224,8'd125} : s = 349;
	{8'd224,8'd126} : s = 350;
	{8'd224,8'd127} : s = 351;
	{8'd224,8'd128} : s = 352;
	{8'd224,8'd129} : s = 353;
	{8'd224,8'd130} : s = 354;
	{8'd224,8'd131} : s = 355;
	{8'd224,8'd132} : s = 356;
	{8'd224,8'd133} : s = 357;
	{8'd224,8'd134} : s = 358;
	{8'd224,8'd135} : s = 359;
	{8'd224,8'd136} : s = 360;
	{8'd224,8'd137} : s = 361;
	{8'd224,8'd138} : s = 362;
	{8'd224,8'd139} : s = 363;
	{8'd224,8'd140} : s = 364;
	{8'd224,8'd141} : s = 365;
	{8'd224,8'd142} : s = 366;
	{8'd224,8'd143} : s = 367;
	{8'd224,8'd144} : s = 368;
	{8'd224,8'd145} : s = 369;
	{8'd224,8'd146} : s = 370;
	{8'd224,8'd147} : s = 371;
	{8'd224,8'd148} : s = 372;
	{8'd224,8'd149} : s = 373;
	{8'd224,8'd150} : s = 374;
	{8'd224,8'd151} : s = 375;
	{8'd224,8'd152} : s = 376;
	{8'd224,8'd153} : s = 377;
	{8'd224,8'd154} : s = 378;
	{8'd224,8'd155} : s = 379;
	{8'd224,8'd156} : s = 380;
	{8'd224,8'd157} : s = 381;
	{8'd224,8'd158} : s = 382;
	{8'd224,8'd159} : s = 383;
	{8'd224,8'd160} : s = 384;
	{8'd224,8'd161} : s = 385;
	{8'd224,8'd162} : s = 386;
	{8'd224,8'd163} : s = 387;
	{8'd224,8'd164} : s = 388;
	{8'd224,8'd165} : s = 389;
	{8'd224,8'd166} : s = 390;
	{8'd224,8'd167} : s = 391;
	{8'd224,8'd168} : s = 392;
	{8'd224,8'd169} : s = 393;
	{8'd224,8'd170} : s = 394;
	{8'd224,8'd171} : s = 395;
	{8'd224,8'd172} : s = 396;
	{8'd224,8'd173} : s = 397;
	{8'd224,8'd174} : s = 398;
	{8'd224,8'd175} : s = 399;
	{8'd224,8'd176} : s = 400;
	{8'd224,8'd177} : s = 401;
	{8'd224,8'd178} : s = 402;
	{8'd224,8'd179} : s = 403;
	{8'd224,8'd180} : s = 404;
	{8'd224,8'd181} : s = 405;
	{8'd224,8'd182} : s = 406;
	{8'd224,8'd183} : s = 407;
	{8'd224,8'd184} : s = 408;
	{8'd224,8'd185} : s = 409;
	{8'd224,8'd186} : s = 410;
	{8'd224,8'd187} : s = 411;
	{8'd224,8'd188} : s = 412;
	{8'd224,8'd189} : s = 413;
	{8'd224,8'd190} : s = 414;
	{8'd224,8'd191} : s = 415;
	{8'd224,8'd192} : s = 416;
	{8'd224,8'd193} : s = 417;
	{8'd224,8'd194} : s = 418;
	{8'd224,8'd195} : s = 419;
	{8'd224,8'd196} : s = 420;
	{8'd224,8'd197} : s = 421;
	{8'd224,8'd198} : s = 422;
	{8'd224,8'd199} : s = 423;
	{8'd224,8'd200} : s = 424;
	{8'd224,8'd201} : s = 425;
	{8'd224,8'd202} : s = 426;
	{8'd224,8'd203} : s = 427;
	{8'd224,8'd204} : s = 428;
	{8'd224,8'd205} : s = 429;
	{8'd224,8'd206} : s = 430;
	{8'd224,8'd207} : s = 431;
	{8'd224,8'd208} : s = 432;
	{8'd224,8'd209} : s = 433;
	{8'd224,8'd210} : s = 434;
	{8'd224,8'd211} : s = 435;
	{8'd224,8'd212} : s = 436;
	{8'd224,8'd213} : s = 437;
	{8'd224,8'd214} : s = 438;
	{8'd224,8'd215} : s = 439;
	{8'd224,8'd216} : s = 440;
	{8'd224,8'd217} : s = 441;
	{8'd224,8'd218} : s = 442;
	{8'd224,8'd219} : s = 443;
	{8'd224,8'd220} : s = 444;
	{8'd224,8'd221} : s = 445;
	{8'd224,8'd222} : s = 446;
	{8'd224,8'd223} : s = 447;
	{8'd224,8'd224} : s = 448;
	{8'd224,8'd225} : s = 449;
	{8'd224,8'd226} : s = 450;
	{8'd224,8'd227} : s = 451;
	{8'd224,8'd228} : s = 452;
	{8'd224,8'd229} : s = 453;
	{8'd224,8'd230} : s = 454;
	{8'd224,8'd231} : s = 455;
	{8'd224,8'd232} : s = 456;
	{8'd224,8'd233} : s = 457;
	{8'd224,8'd234} : s = 458;
	{8'd224,8'd235} : s = 459;
	{8'd224,8'd236} : s = 460;
	{8'd224,8'd237} : s = 461;
	{8'd224,8'd238} : s = 462;
	{8'd224,8'd239} : s = 463;
	{8'd224,8'd240} : s = 464;
	{8'd224,8'd241} : s = 465;
	{8'd224,8'd242} : s = 466;
	{8'd224,8'd243} : s = 467;
	{8'd224,8'd244} : s = 468;
	{8'd224,8'd245} : s = 469;
	{8'd224,8'd246} : s = 470;
	{8'd224,8'd247} : s = 471;
	{8'd224,8'd248} : s = 472;
	{8'd224,8'd249} : s = 473;
	{8'd224,8'd250} : s = 474;
	{8'd224,8'd251} : s = 475;
	{8'd224,8'd252} : s = 476;
	{8'd224,8'd253} : s = 477;
	{8'd224,8'd254} : s = 478;
	{8'd224,8'd255} : s = 479;
	{8'd225,8'd0} : s = 225;
	{8'd225,8'd1} : s = 226;
	{8'd225,8'd2} : s = 227;
	{8'd225,8'd3} : s = 228;
	{8'd225,8'd4} : s = 229;
	{8'd225,8'd5} : s = 230;
	{8'd225,8'd6} : s = 231;
	{8'd225,8'd7} : s = 232;
	{8'd225,8'd8} : s = 233;
	{8'd225,8'd9} : s = 234;
	{8'd225,8'd10} : s = 235;
	{8'd225,8'd11} : s = 236;
	{8'd225,8'd12} : s = 237;
	{8'd225,8'd13} : s = 238;
	{8'd225,8'd14} : s = 239;
	{8'd225,8'd15} : s = 240;
	{8'd225,8'd16} : s = 241;
	{8'd225,8'd17} : s = 242;
	{8'd225,8'd18} : s = 243;
	{8'd225,8'd19} : s = 244;
	{8'd225,8'd20} : s = 245;
	{8'd225,8'd21} : s = 246;
	{8'd225,8'd22} : s = 247;
	{8'd225,8'd23} : s = 248;
	{8'd225,8'd24} : s = 249;
	{8'd225,8'd25} : s = 250;
	{8'd225,8'd26} : s = 251;
	{8'd225,8'd27} : s = 252;
	{8'd225,8'd28} : s = 253;
	{8'd225,8'd29} : s = 254;
	{8'd225,8'd30} : s = 255;
	{8'd225,8'd31} : s = 256;
	{8'd225,8'd32} : s = 257;
	{8'd225,8'd33} : s = 258;
	{8'd225,8'd34} : s = 259;
	{8'd225,8'd35} : s = 260;
	{8'd225,8'd36} : s = 261;
	{8'd225,8'd37} : s = 262;
	{8'd225,8'd38} : s = 263;
	{8'd225,8'd39} : s = 264;
	{8'd225,8'd40} : s = 265;
	{8'd225,8'd41} : s = 266;
	{8'd225,8'd42} : s = 267;
	{8'd225,8'd43} : s = 268;
	{8'd225,8'd44} : s = 269;
	{8'd225,8'd45} : s = 270;
	{8'd225,8'd46} : s = 271;
	{8'd225,8'd47} : s = 272;
	{8'd225,8'd48} : s = 273;
	{8'd225,8'd49} : s = 274;
	{8'd225,8'd50} : s = 275;
	{8'd225,8'd51} : s = 276;
	{8'd225,8'd52} : s = 277;
	{8'd225,8'd53} : s = 278;
	{8'd225,8'd54} : s = 279;
	{8'd225,8'd55} : s = 280;
	{8'd225,8'd56} : s = 281;
	{8'd225,8'd57} : s = 282;
	{8'd225,8'd58} : s = 283;
	{8'd225,8'd59} : s = 284;
	{8'd225,8'd60} : s = 285;
	{8'd225,8'd61} : s = 286;
	{8'd225,8'd62} : s = 287;
	{8'd225,8'd63} : s = 288;
	{8'd225,8'd64} : s = 289;
	{8'd225,8'd65} : s = 290;
	{8'd225,8'd66} : s = 291;
	{8'd225,8'd67} : s = 292;
	{8'd225,8'd68} : s = 293;
	{8'd225,8'd69} : s = 294;
	{8'd225,8'd70} : s = 295;
	{8'd225,8'd71} : s = 296;
	{8'd225,8'd72} : s = 297;
	{8'd225,8'd73} : s = 298;
	{8'd225,8'd74} : s = 299;
	{8'd225,8'd75} : s = 300;
	{8'd225,8'd76} : s = 301;
	{8'd225,8'd77} : s = 302;
	{8'd225,8'd78} : s = 303;
	{8'd225,8'd79} : s = 304;
	{8'd225,8'd80} : s = 305;
	{8'd225,8'd81} : s = 306;
	{8'd225,8'd82} : s = 307;
	{8'd225,8'd83} : s = 308;
	{8'd225,8'd84} : s = 309;
	{8'd225,8'd85} : s = 310;
	{8'd225,8'd86} : s = 311;
	{8'd225,8'd87} : s = 312;
	{8'd225,8'd88} : s = 313;
	{8'd225,8'd89} : s = 314;
	{8'd225,8'd90} : s = 315;
	{8'd225,8'd91} : s = 316;
	{8'd225,8'd92} : s = 317;
	{8'd225,8'd93} : s = 318;
	{8'd225,8'd94} : s = 319;
	{8'd225,8'd95} : s = 320;
	{8'd225,8'd96} : s = 321;
	{8'd225,8'd97} : s = 322;
	{8'd225,8'd98} : s = 323;
	{8'd225,8'd99} : s = 324;
	{8'd225,8'd100} : s = 325;
	{8'd225,8'd101} : s = 326;
	{8'd225,8'd102} : s = 327;
	{8'd225,8'd103} : s = 328;
	{8'd225,8'd104} : s = 329;
	{8'd225,8'd105} : s = 330;
	{8'd225,8'd106} : s = 331;
	{8'd225,8'd107} : s = 332;
	{8'd225,8'd108} : s = 333;
	{8'd225,8'd109} : s = 334;
	{8'd225,8'd110} : s = 335;
	{8'd225,8'd111} : s = 336;
	{8'd225,8'd112} : s = 337;
	{8'd225,8'd113} : s = 338;
	{8'd225,8'd114} : s = 339;
	{8'd225,8'd115} : s = 340;
	{8'd225,8'd116} : s = 341;
	{8'd225,8'd117} : s = 342;
	{8'd225,8'd118} : s = 343;
	{8'd225,8'd119} : s = 344;
	{8'd225,8'd120} : s = 345;
	{8'd225,8'd121} : s = 346;
	{8'd225,8'd122} : s = 347;
	{8'd225,8'd123} : s = 348;
	{8'd225,8'd124} : s = 349;
	{8'd225,8'd125} : s = 350;
	{8'd225,8'd126} : s = 351;
	{8'd225,8'd127} : s = 352;
	{8'd225,8'd128} : s = 353;
	{8'd225,8'd129} : s = 354;
	{8'd225,8'd130} : s = 355;
	{8'd225,8'd131} : s = 356;
	{8'd225,8'd132} : s = 357;
	{8'd225,8'd133} : s = 358;
	{8'd225,8'd134} : s = 359;
	{8'd225,8'd135} : s = 360;
	{8'd225,8'd136} : s = 361;
	{8'd225,8'd137} : s = 362;
	{8'd225,8'd138} : s = 363;
	{8'd225,8'd139} : s = 364;
	{8'd225,8'd140} : s = 365;
	{8'd225,8'd141} : s = 366;
	{8'd225,8'd142} : s = 367;
	{8'd225,8'd143} : s = 368;
	{8'd225,8'd144} : s = 369;
	{8'd225,8'd145} : s = 370;
	{8'd225,8'd146} : s = 371;
	{8'd225,8'd147} : s = 372;
	{8'd225,8'd148} : s = 373;
	{8'd225,8'd149} : s = 374;
	{8'd225,8'd150} : s = 375;
	{8'd225,8'd151} : s = 376;
	{8'd225,8'd152} : s = 377;
	{8'd225,8'd153} : s = 378;
	{8'd225,8'd154} : s = 379;
	{8'd225,8'd155} : s = 380;
	{8'd225,8'd156} : s = 381;
	{8'd225,8'd157} : s = 382;
	{8'd225,8'd158} : s = 383;
	{8'd225,8'd159} : s = 384;
	{8'd225,8'd160} : s = 385;
	{8'd225,8'd161} : s = 386;
	{8'd225,8'd162} : s = 387;
	{8'd225,8'd163} : s = 388;
	{8'd225,8'd164} : s = 389;
	{8'd225,8'd165} : s = 390;
	{8'd225,8'd166} : s = 391;
	{8'd225,8'd167} : s = 392;
	{8'd225,8'd168} : s = 393;
	{8'd225,8'd169} : s = 394;
	{8'd225,8'd170} : s = 395;
	{8'd225,8'd171} : s = 396;
	{8'd225,8'd172} : s = 397;
	{8'd225,8'd173} : s = 398;
	{8'd225,8'd174} : s = 399;
	{8'd225,8'd175} : s = 400;
	{8'd225,8'd176} : s = 401;
	{8'd225,8'd177} : s = 402;
	{8'd225,8'd178} : s = 403;
	{8'd225,8'd179} : s = 404;
	{8'd225,8'd180} : s = 405;
	{8'd225,8'd181} : s = 406;
	{8'd225,8'd182} : s = 407;
	{8'd225,8'd183} : s = 408;
	{8'd225,8'd184} : s = 409;
	{8'd225,8'd185} : s = 410;
	{8'd225,8'd186} : s = 411;
	{8'd225,8'd187} : s = 412;
	{8'd225,8'd188} : s = 413;
	{8'd225,8'd189} : s = 414;
	{8'd225,8'd190} : s = 415;
	{8'd225,8'd191} : s = 416;
	{8'd225,8'd192} : s = 417;
	{8'd225,8'd193} : s = 418;
	{8'd225,8'd194} : s = 419;
	{8'd225,8'd195} : s = 420;
	{8'd225,8'd196} : s = 421;
	{8'd225,8'd197} : s = 422;
	{8'd225,8'd198} : s = 423;
	{8'd225,8'd199} : s = 424;
	{8'd225,8'd200} : s = 425;
	{8'd225,8'd201} : s = 426;
	{8'd225,8'd202} : s = 427;
	{8'd225,8'd203} : s = 428;
	{8'd225,8'd204} : s = 429;
	{8'd225,8'd205} : s = 430;
	{8'd225,8'd206} : s = 431;
	{8'd225,8'd207} : s = 432;
	{8'd225,8'd208} : s = 433;
	{8'd225,8'd209} : s = 434;
	{8'd225,8'd210} : s = 435;
	{8'd225,8'd211} : s = 436;
	{8'd225,8'd212} : s = 437;
	{8'd225,8'd213} : s = 438;
	{8'd225,8'd214} : s = 439;
	{8'd225,8'd215} : s = 440;
	{8'd225,8'd216} : s = 441;
	{8'd225,8'd217} : s = 442;
	{8'd225,8'd218} : s = 443;
	{8'd225,8'd219} : s = 444;
	{8'd225,8'd220} : s = 445;
	{8'd225,8'd221} : s = 446;
	{8'd225,8'd222} : s = 447;
	{8'd225,8'd223} : s = 448;
	{8'd225,8'd224} : s = 449;
	{8'd225,8'd225} : s = 450;
	{8'd225,8'd226} : s = 451;
	{8'd225,8'd227} : s = 452;
	{8'd225,8'd228} : s = 453;
	{8'd225,8'd229} : s = 454;
	{8'd225,8'd230} : s = 455;
	{8'd225,8'd231} : s = 456;
	{8'd225,8'd232} : s = 457;
	{8'd225,8'd233} : s = 458;
	{8'd225,8'd234} : s = 459;
	{8'd225,8'd235} : s = 460;
	{8'd225,8'd236} : s = 461;
	{8'd225,8'd237} : s = 462;
	{8'd225,8'd238} : s = 463;
	{8'd225,8'd239} : s = 464;
	{8'd225,8'd240} : s = 465;
	{8'd225,8'd241} : s = 466;
	{8'd225,8'd242} : s = 467;
	{8'd225,8'd243} : s = 468;
	{8'd225,8'd244} : s = 469;
	{8'd225,8'd245} : s = 470;
	{8'd225,8'd246} : s = 471;
	{8'd225,8'd247} : s = 472;
	{8'd225,8'd248} : s = 473;
	{8'd225,8'd249} : s = 474;
	{8'd225,8'd250} : s = 475;
	{8'd225,8'd251} : s = 476;
	{8'd225,8'd252} : s = 477;
	{8'd225,8'd253} : s = 478;
	{8'd225,8'd254} : s = 479;
	{8'd225,8'd255} : s = 480;
	{8'd226,8'd0} : s = 226;
	{8'd226,8'd1} : s = 227;
	{8'd226,8'd2} : s = 228;
	{8'd226,8'd3} : s = 229;
	{8'd226,8'd4} : s = 230;
	{8'd226,8'd5} : s = 231;
	{8'd226,8'd6} : s = 232;
	{8'd226,8'd7} : s = 233;
	{8'd226,8'd8} : s = 234;
	{8'd226,8'd9} : s = 235;
	{8'd226,8'd10} : s = 236;
	{8'd226,8'd11} : s = 237;
	{8'd226,8'd12} : s = 238;
	{8'd226,8'd13} : s = 239;
	{8'd226,8'd14} : s = 240;
	{8'd226,8'd15} : s = 241;
	{8'd226,8'd16} : s = 242;
	{8'd226,8'd17} : s = 243;
	{8'd226,8'd18} : s = 244;
	{8'd226,8'd19} : s = 245;
	{8'd226,8'd20} : s = 246;
	{8'd226,8'd21} : s = 247;
	{8'd226,8'd22} : s = 248;
	{8'd226,8'd23} : s = 249;
	{8'd226,8'd24} : s = 250;
	{8'd226,8'd25} : s = 251;
	{8'd226,8'd26} : s = 252;
	{8'd226,8'd27} : s = 253;
	{8'd226,8'd28} : s = 254;
	{8'd226,8'd29} : s = 255;
	{8'd226,8'd30} : s = 256;
	{8'd226,8'd31} : s = 257;
	{8'd226,8'd32} : s = 258;
	{8'd226,8'd33} : s = 259;
	{8'd226,8'd34} : s = 260;
	{8'd226,8'd35} : s = 261;
	{8'd226,8'd36} : s = 262;
	{8'd226,8'd37} : s = 263;
	{8'd226,8'd38} : s = 264;
	{8'd226,8'd39} : s = 265;
	{8'd226,8'd40} : s = 266;
	{8'd226,8'd41} : s = 267;
	{8'd226,8'd42} : s = 268;
	{8'd226,8'd43} : s = 269;
	{8'd226,8'd44} : s = 270;
	{8'd226,8'd45} : s = 271;
	{8'd226,8'd46} : s = 272;
	{8'd226,8'd47} : s = 273;
	{8'd226,8'd48} : s = 274;
	{8'd226,8'd49} : s = 275;
	{8'd226,8'd50} : s = 276;
	{8'd226,8'd51} : s = 277;
	{8'd226,8'd52} : s = 278;
	{8'd226,8'd53} : s = 279;
	{8'd226,8'd54} : s = 280;
	{8'd226,8'd55} : s = 281;
	{8'd226,8'd56} : s = 282;
	{8'd226,8'd57} : s = 283;
	{8'd226,8'd58} : s = 284;
	{8'd226,8'd59} : s = 285;
	{8'd226,8'd60} : s = 286;
	{8'd226,8'd61} : s = 287;
	{8'd226,8'd62} : s = 288;
	{8'd226,8'd63} : s = 289;
	{8'd226,8'd64} : s = 290;
	{8'd226,8'd65} : s = 291;
	{8'd226,8'd66} : s = 292;
	{8'd226,8'd67} : s = 293;
	{8'd226,8'd68} : s = 294;
	{8'd226,8'd69} : s = 295;
	{8'd226,8'd70} : s = 296;
	{8'd226,8'd71} : s = 297;
	{8'd226,8'd72} : s = 298;
	{8'd226,8'd73} : s = 299;
	{8'd226,8'd74} : s = 300;
	{8'd226,8'd75} : s = 301;
	{8'd226,8'd76} : s = 302;
	{8'd226,8'd77} : s = 303;
	{8'd226,8'd78} : s = 304;
	{8'd226,8'd79} : s = 305;
	{8'd226,8'd80} : s = 306;
	{8'd226,8'd81} : s = 307;
	{8'd226,8'd82} : s = 308;
	{8'd226,8'd83} : s = 309;
	{8'd226,8'd84} : s = 310;
	{8'd226,8'd85} : s = 311;
	{8'd226,8'd86} : s = 312;
	{8'd226,8'd87} : s = 313;
	{8'd226,8'd88} : s = 314;
	{8'd226,8'd89} : s = 315;
	{8'd226,8'd90} : s = 316;
	{8'd226,8'd91} : s = 317;
	{8'd226,8'd92} : s = 318;
	{8'd226,8'd93} : s = 319;
	{8'd226,8'd94} : s = 320;
	{8'd226,8'd95} : s = 321;
	{8'd226,8'd96} : s = 322;
	{8'd226,8'd97} : s = 323;
	{8'd226,8'd98} : s = 324;
	{8'd226,8'd99} : s = 325;
	{8'd226,8'd100} : s = 326;
	{8'd226,8'd101} : s = 327;
	{8'd226,8'd102} : s = 328;
	{8'd226,8'd103} : s = 329;
	{8'd226,8'd104} : s = 330;
	{8'd226,8'd105} : s = 331;
	{8'd226,8'd106} : s = 332;
	{8'd226,8'd107} : s = 333;
	{8'd226,8'd108} : s = 334;
	{8'd226,8'd109} : s = 335;
	{8'd226,8'd110} : s = 336;
	{8'd226,8'd111} : s = 337;
	{8'd226,8'd112} : s = 338;
	{8'd226,8'd113} : s = 339;
	{8'd226,8'd114} : s = 340;
	{8'd226,8'd115} : s = 341;
	{8'd226,8'd116} : s = 342;
	{8'd226,8'd117} : s = 343;
	{8'd226,8'd118} : s = 344;
	{8'd226,8'd119} : s = 345;
	{8'd226,8'd120} : s = 346;
	{8'd226,8'd121} : s = 347;
	{8'd226,8'd122} : s = 348;
	{8'd226,8'd123} : s = 349;
	{8'd226,8'd124} : s = 350;
	{8'd226,8'd125} : s = 351;
	{8'd226,8'd126} : s = 352;
	{8'd226,8'd127} : s = 353;
	{8'd226,8'd128} : s = 354;
	{8'd226,8'd129} : s = 355;
	{8'd226,8'd130} : s = 356;
	{8'd226,8'd131} : s = 357;
	{8'd226,8'd132} : s = 358;
	{8'd226,8'd133} : s = 359;
	{8'd226,8'd134} : s = 360;
	{8'd226,8'd135} : s = 361;
	{8'd226,8'd136} : s = 362;
	{8'd226,8'd137} : s = 363;
	{8'd226,8'd138} : s = 364;
	{8'd226,8'd139} : s = 365;
	{8'd226,8'd140} : s = 366;
	{8'd226,8'd141} : s = 367;
	{8'd226,8'd142} : s = 368;
	{8'd226,8'd143} : s = 369;
	{8'd226,8'd144} : s = 370;
	{8'd226,8'd145} : s = 371;
	{8'd226,8'd146} : s = 372;
	{8'd226,8'd147} : s = 373;
	{8'd226,8'd148} : s = 374;
	{8'd226,8'd149} : s = 375;
	{8'd226,8'd150} : s = 376;
	{8'd226,8'd151} : s = 377;
	{8'd226,8'd152} : s = 378;
	{8'd226,8'd153} : s = 379;
	{8'd226,8'd154} : s = 380;
	{8'd226,8'd155} : s = 381;
	{8'd226,8'd156} : s = 382;
	{8'd226,8'd157} : s = 383;
	{8'd226,8'd158} : s = 384;
	{8'd226,8'd159} : s = 385;
	{8'd226,8'd160} : s = 386;
	{8'd226,8'd161} : s = 387;
	{8'd226,8'd162} : s = 388;
	{8'd226,8'd163} : s = 389;
	{8'd226,8'd164} : s = 390;
	{8'd226,8'd165} : s = 391;
	{8'd226,8'd166} : s = 392;
	{8'd226,8'd167} : s = 393;
	{8'd226,8'd168} : s = 394;
	{8'd226,8'd169} : s = 395;
	{8'd226,8'd170} : s = 396;
	{8'd226,8'd171} : s = 397;
	{8'd226,8'd172} : s = 398;
	{8'd226,8'd173} : s = 399;
	{8'd226,8'd174} : s = 400;
	{8'd226,8'd175} : s = 401;
	{8'd226,8'd176} : s = 402;
	{8'd226,8'd177} : s = 403;
	{8'd226,8'd178} : s = 404;
	{8'd226,8'd179} : s = 405;
	{8'd226,8'd180} : s = 406;
	{8'd226,8'd181} : s = 407;
	{8'd226,8'd182} : s = 408;
	{8'd226,8'd183} : s = 409;
	{8'd226,8'd184} : s = 410;
	{8'd226,8'd185} : s = 411;
	{8'd226,8'd186} : s = 412;
	{8'd226,8'd187} : s = 413;
	{8'd226,8'd188} : s = 414;
	{8'd226,8'd189} : s = 415;
	{8'd226,8'd190} : s = 416;
	{8'd226,8'd191} : s = 417;
	{8'd226,8'd192} : s = 418;
	{8'd226,8'd193} : s = 419;
	{8'd226,8'd194} : s = 420;
	{8'd226,8'd195} : s = 421;
	{8'd226,8'd196} : s = 422;
	{8'd226,8'd197} : s = 423;
	{8'd226,8'd198} : s = 424;
	{8'd226,8'd199} : s = 425;
	{8'd226,8'd200} : s = 426;
	{8'd226,8'd201} : s = 427;
	{8'd226,8'd202} : s = 428;
	{8'd226,8'd203} : s = 429;
	{8'd226,8'd204} : s = 430;
	{8'd226,8'd205} : s = 431;
	{8'd226,8'd206} : s = 432;
	{8'd226,8'd207} : s = 433;
	{8'd226,8'd208} : s = 434;
	{8'd226,8'd209} : s = 435;
	{8'd226,8'd210} : s = 436;
	{8'd226,8'd211} : s = 437;
	{8'd226,8'd212} : s = 438;
	{8'd226,8'd213} : s = 439;
	{8'd226,8'd214} : s = 440;
	{8'd226,8'd215} : s = 441;
	{8'd226,8'd216} : s = 442;
	{8'd226,8'd217} : s = 443;
	{8'd226,8'd218} : s = 444;
	{8'd226,8'd219} : s = 445;
	{8'd226,8'd220} : s = 446;
	{8'd226,8'd221} : s = 447;
	{8'd226,8'd222} : s = 448;
	{8'd226,8'd223} : s = 449;
	{8'd226,8'd224} : s = 450;
	{8'd226,8'd225} : s = 451;
	{8'd226,8'd226} : s = 452;
	{8'd226,8'd227} : s = 453;
	{8'd226,8'd228} : s = 454;
	{8'd226,8'd229} : s = 455;
	{8'd226,8'd230} : s = 456;
	{8'd226,8'd231} : s = 457;
	{8'd226,8'd232} : s = 458;
	{8'd226,8'd233} : s = 459;
	{8'd226,8'd234} : s = 460;
	{8'd226,8'd235} : s = 461;
	{8'd226,8'd236} : s = 462;
	{8'd226,8'd237} : s = 463;
	{8'd226,8'd238} : s = 464;
	{8'd226,8'd239} : s = 465;
	{8'd226,8'd240} : s = 466;
	{8'd226,8'd241} : s = 467;
	{8'd226,8'd242} : s = 468;
	{8'd226,8'd243} : s = 469;
	{8'd226,8'd244} : s = 470;
	{8'd226,8'd245} : s = 471;
	{8'd226,8'd246} : s = 472;
	{8'd226,8'd247} : s = 473;
	{8'd226,8'd248} : s = 474;
	{8'd226,8'd249} : s = 475;
	{8'd226,8'd250} : s = 476;
	{8'd226,8'd251} : s = 477;
	{8'd226,8'd252} : s = 478;
	{8'd226,8'd253} : s = 479;
	{8'd226,8'd254} : s = 480;
	{8'd226,8'd255} : s = 481;
	{8'd227,8'd0} : s = 227;
	{8'd227,8'd1} : s = 228;
	{8'd227,8'd2} : s = 229;
	{8'd227,8'd3} : s = 230;
	{8'd227,8'd4} : s = 231;
	{8'd227,8'd5} : s = 232;
	{8'd227,8'd6} : s = 233;
	{8'd227,8'd7} : s = 234;
	{8'd227,8'd8} : s = 235;
	{8'd227,8'd9} : s = 236;
	{8'd227,8'd10} : s = 237;
	{8'd227,8'd11} : s = 238;
	{8'd227,8'd12} : s = 239;
	{8'd227,8'd13} : s = 240;
	{8'd227,8'd14} : s = 241;
	{8'd227,8'd15} : s = 242;
	{8'd227,8'd16} : s = 243;
	{8'd227,8'd17} : s = 244;
	{8'd227,8'd18} : s = 245;
	{8'd227,8'd19} : s = 246;
	{8'd227,8'd20} : s = 247;
	{8'd227,8'd21} : s = 248;
	{8'd227,8'd22} : s = 249;
	{8'd227,8'd23} : s = 250;
	{8'd227,8'd24} : s = 251;
	{8'd227,8'd25} : s = 252;
	{8'd227,8'd26} : s = 253;
	{8'd227,8'd27} : s = 254;
	{8'd227,8'd28} : s = 255;
	{8'd227,8'd29} : s = 256;
	{8'd227,8'd30} : s = 257;
	{8'd227,8'd31} : s = 258;
	{8'd227,8'd32} : s = 259;
	{8'd227,8'd33} : s = 260;
	{8'd227,8'd34} : s = 261;
	{8'd227,8'd35} : s = 262;
	{8'd227,8'd36} : s = 263;
	{8'd227,8'd37} : s = 264;
	{8'd227,8'd38} : s = 265;
	{8'd227,8'd39} : s = 266;
	{8'd227,8'd40} : s = 267;
	{8'd227,8'd41} : s = 268;
	{8'd227,8'd42} : s = 269;
	{8'd227,8'd43} : s = 270;
	{8'd227,8'd44} : s = 271;
	{8'd227,8'd45} : s = 272;
	{8'd227,8'd46} : s = 273;
	{8'd227,8'd47} : s = 274;
	{8'd227,8'd48} : s = 275;
	{8'd227,8'd49} : s = 276;
	{8'd227,8'd50} : s = 277;
	{8'd227,8'd51} : s = 278;
	{8'd227,8'd52} : s = 279;
	{8'd227,8'd53} : s = 280;
	{8'd227,8'd54} : s = 281;
	{8'd227,8'd55} : s = 282;
	{8'd227,8'd56} : s = 283;
	{8'd227,8'd57} : s = 284;
	{8'd227,8'd58} : s = 285;
	{8'd227,8'd59} : s = 286;
	{8'd227,8'd60} : s = 287;
	{8'd227,8'd61} : s = 288;
	{8'd227,8'd62} : s = 289;
	{8'd227,8'd63} : s = 290;
	{8'd227,8'd64} : s = 291;
	{8'd227,8'd65} : s = 292;
	{8'd227,8'd66} : s = 293;
	{8'd227,8'd67} : s = 294;
	{8'd227,8'd68} : s = 295;
	{8'd227,8'd69} : s = 296;
	{8'd227,8'd70} : s = 297;
	{8'd227,8'd71} : s = 298;
	{8'd227,8'd72} : s = 299;
	{8'd227,8'd73} : s = 300;
	{8'd227,8'd74} : s = 301;
	{8'd227,8'd75} : s = 302;
	{8'd227,8'd76} : s = 303;
	{8'd227,8'd77} : s = 304;
	{8'd227,8'd78} : s = 305;
	{8'd227,8'd79} : s = 306;
	{8'd227,8'd80} : s = 307;
	{8'd227,8'd81} : s = 308;
	{8'd227,8'd82} : s = 309;
	{8'd227,8'd83} : s = 310;
	{8'd227,8'd84} : s = 311;
	{8'd227,8'd85} : s = 312;
	{8'd227,8'd86} : s = 313;
	{8'd227,8'd87} : s = 314;
	{8'd227,8'd88} : s = 315;
	{8'd227,8'd89} : s = 316;
	{8'd227,8'd90} : s = 317;
	{8'd227,8'd91} : s = 318;
	{8'd227,8'd92} : s = 319;
	{8'd227,8'd93} : s = 320;
	{8'd227,8'd94} : s = 321;
	{8'd227,8'd95} : s = 322;
	{8'd227,8'd96} : s = 323;
	{8'd227,8'd97} : s = 324;
	{8'd227,8'd98} : s = 325;
	{8'd227,8'd99} : s = 326;
	{8'd227,8'd100} : s = 327;
	{8'd227,8'd101} : s = 328;
	{8'd227,8'd102} : s = 329;
	{8'd227,8'd103} : s = 330;
	{8'd227,8'd104} : s = 331;
	{8'd227,8'd105} : s = 332;
	{8'd227,8'd106} : s = 333;
	{8'd227,8'd107} : s = 334;
	{8'd227,8'd108} : s = 335;
	{8'd227,8'd109} : s = 336;
	{8'd227,8'd110} : s = 337;
	{8'd227,8'd111} : s = 338;
	{8'd227,8'd112} : s = 339;
	{8'd227,8'd113} : s = 340;
	{8'd227,8'd114} : s = 341;
	{8'd227,8'd115} : s = 342;
	{8'd227,8'd116} : s = 343;
	{8'd227,8'd117} : s = 344;
	{8'd227,8'd118} : s = 345;
	{8'd227,8'd119} : s = 346;
	{8'd227,8'd120} : s = 347;
	{8'd227,8'd121} : s = 348;
	{8'd227,8'd122} : s = 349;
	{8'd227,8'd123} : s = 350;
	{8'd227,8'd124} : s = 351;
	{8'd227,8'd125} : s = 352;
	{8'd227,8'd126} : s = 353;
	{8'd227,8'd127} : s = 354;
	{8'd227,8'd128} : s = 355;
	{8'd227,8'd129} : s = 356;
	{8'd227,8'd130} : s = 357;
	{8'd227,8'd131} : s = 358;
	{8'd227,8'd132} : s = 359;
	{8'd227,8'd133} : s = 360;
	{8'd227,8'd134} : s = 361;
	{8'd227,8'd135} : s = 362;
	{8'd227,8'd136} : s = 363;
	{8'd227,8'd137} : s = 364;
	{8'd227,8'd138} : s = 365;
	{8'd227,8'd139} : s = 366;
	{8'd227,8'd140} : s = 367;
	{8'd227,8'd141} : s = 368;
	{8'd227,8'd142} : s = 369;
	{8'd227,8'd143} : s = 370;
	{8'd227,8'd144} : s = 371;
	{8'd227,8'd145} : s = 372;
	{8'd227,8'd146} : s = 373;
	{8'd227,8'd147} : s = 374;
	{8'd227,8'd148} : s = 375;
	{8'd227,8'd149} : s = 376;
	{8'd227,8'd150} : s = 377;
	{8'd227,8'd151} : s = 378;
	{8'd227,8'd152} : s = 379;
	{8'd227,8'd153} : s = 380;
	{8'd227,8'd154} : s = 381;
	{8'd227,8'd155} : s = 382;
	{8'd227,8'd156} : s = 383;
	{8'd227,8'd157} : s = 384;
	{8'd227,8'd158} : s = 385;
	{8'd227,8'd159} : s = 386;
	{8'd227,8'd160} : s = 387;
	{8'd227,8'd161} : s = 388;
	{8'd227,8'd162} : s = 389;
	{8'd227,8'd163} : s = 390;
	{8'd227,8'd164} : s = 391;
	{8'd227,8'd165} : s = 392;
	{8'd227,8'd166} : s = 393;
	{8'd227,8'd167} : s = 394;
	{8'd227,8'd168} : s = 395;
	{8'd227,8'd169} : s = 396;
	{8'd227,8'd170} : s = 397;
	{8'd227,8'd171} : s = 398;
	{8'd227,8'd172} : s = 399;
	{8'd227,8'd173} : s = 400;
	{8'd227,8'd174} : s = 401;
	{8'd227,8'd175} : s = 402;
	{8'd227,8'd176} : s = 403;
	{8'd227,8'd177} : s = 404;
	{8'd227,8'd178} : s = 405;
	{8'd227,8'd179} : s = 406;
	{8'd227,8'd180} : s = 407;
	{8'd227,8'd181} : s = 408;
	{8'd227,8'd182} : s = 409;
	{8'd227,8'd183} : s = 410;
	{8'd227,8'd184} : s = 411;
	{8'd227,8'd185} : s = 412;
	{8'd227,8'd186} : s = 413;
	{8'd227,8'd187} : s = 414;
	{8'd227,8'd188} : s = 415;
	{8'd227,8'd189} : s = 416;
	{8'd227,8'd190} : s = 417;
	{8'd227,8'd191} : s = 418;
	{8'd227,8'd192} : s = 419;
	{8'd227,8'd193} : s = 420;
	{8'd227,8'd194} : s = 421;
	{8'd227,8'd195} : s = 422;
	{8'd227,8'd196} : s = 423;
	{8'd227,8'd197} : s = 424;
	{8'd227,8'd198} : s = 425;
	{8'd227,8'd199} : s = 426;
	{8'd227,8'd200} : s = 427;
	{8'd227,8'd201} : s = 428;
	{8'd227,8'd202} : s = 429;
	{8'd227,8'd203} : s = 430;
	{8'd227,8'd204} : s = 431;
	{8'd227,8'd205} : s = 432;
	{8'd227,8'd206} : s = 433;
	{8'd227,8'd207} : s = 434;
	{8'd227,8'd208} : s = 435;
	{8'd227,8'd209} : s = 436;
	{8'd227,8'd210} : s = 437;
	{8'd227,8'd211} : s = 438;
	{8'd227,8'd212} : s = 439;
	{8'd227,8'd213} : s = 440;
	{8'd227,8'd214} : s = 441;
	{8'd227,8'd215} : s = 442;
	{8'd227,8'd216} : s = 443;
	{8'd227,8'd217} : s = 444;
	{8'd227,8'd218} : s = 445;
	{8'd227,8'd219} : s = 446;
	{8'd227,8'd220} : s = 447;
	{8'd227,8'd221} : s = 448;
	{8'd227,8'd222} : s = 449;
	{8'd227,8'd223} : s = 450;
	{8'd227,8'd224} : s = 451;
	{8'd227,8'd225} : s = 452;
	{8'd227,8'd226} : s = 453;
	{8'd227,8'd227} : s = 454;
	{8'd227,8'd228} : s = 455;
	{8'd227,8'd229} : s = 456;
	{8'd227,8'd230} : s = 457;
	{8'd227,8'd231} : s = 458;
	{8'd227,8'd232} : s = 459;
	{8'd227,8'd233} : s = 460;
	{8'd227,8'd234} : s = 461;
	{8'd227,8'd235} : s = 462;
	{8'd227,8'd236} : s = 463;
	{8'd227,8'd237} : s = 464;
	{8'd227,8'd238} : s = 465;
	{8'd227,8'd239} : s = 466;
	{8'd227,8'd240} : s = 467;
	{8'd227,8'd241} : s = 468;
	{8'd227,8'd242} : s = 469;
	{8'd227,8'd243} : s = 470;
	{8'd227,8'd244} : s = 471;
	{8'd227,8'd245} : s = 472;
	{8'd227,8'd246} : s = 473;
	{8'd227,8'd247} : s = 474;
	{8'd227,8'd248} : s = 475;
	{8'd227,8'd249} : s = 476;
	{8'd227,8'd250} : s = 477;
	{8'd227,8'd251} : s = 478;
	{8'd227,8'd252} : s = 479;
	{8'd227,8'd253} : s = 480;
	{8'd227,8'd254} : s = 481;
	{8'd227,8'd255} : s = 482;
	{8'd228,8'd0} : s = 228;
	{8'd228,8'd1} : s = 229;
	{8'd228,8'd2} : s = 230;
	{8'd228,8'd3} : s = 231;
	{8'd228,8'd4} : s = 232;
	{8'd228,8'd5} : s = 233;
	{8'd228,8'd6} : s = 234;
	{8'd228,8'd7} : s = 235;
	{8'd228,8'd8} : s = 236;
	{8'd228,8'd9} : s = 237;
	{8'd228,8'd10} : s = 238;
	{8'd228,8'd11} : s = 239;
	{8'd228,8'd12} : s = 240;
	{8'd228,8'd13} : s = 241;
	{8'd228,8'd14} : s = 242;
	{8'd228,8'd15} : s = 243;
	{8'd228,8'd16} : s = 244;
	{8'd228,8'd17} : s = 245;
	{8'd228,8'd18} : s = 246;
	{8'd228,8'd19} : s = 247;
	{8'd228,8'd20} : s = 248;
	{8'd228,8'd21} : s = 249;
	{8'd228,8'd22} : s = 250;
	{8'd228,8'd23} : s = 251;
	{8'd228,8'd24} : s = 252;
	{8'd228,8'd25} : s = 253;
	{8'd228,8'd26} : s = 254;
	{8'd228,8'd27} : s = 255;
	{8'd228,8'd28} : s = 256;
	{8'd228,8'd29} : s = 257;
	{8'd228,8'd30} : s = 258;
	{8'd228,8'd31} : s = 259;
	{8'd228,8'd32} : s = 260;
	{8'd228,8'd33} : s = 261;
	{8'd228,8'd34} : s = 262;
	{8'd228,8'd35} : s = 263;
	{8'd228,8'd36} : s = 264;
	{8'd228,8'd37} : s = 265;
	{8'd228,8'd38} : s = 266;
	{8'd228,8'd39} : s = 267;
	{8'd228,8'd40} : s = 268;
	{8'd228,8'd41} : s = 269;
	{8'd228,8'd42} : s = 270;
	{8'd228,8'd43} : s = 271;
	{8'd228,8'd44} : s = 272;
	{8'd228,8'd45} : s = 273;
	{8'd228,8'd46} : s = 274;
	{8'd228,8'd47} : s = 275;
	{8'd228,8'd48} : s = 276;
	{8'd228,8'd49} : s = 277;
	{8'd228,8'd50} : s = 278;
	{8'd228,8'd51} : s = 279;
	{8'd228,8'd52} : s = 280;
	{8'd228,8'd53} : s = 281;
	{8'd228,8'd54} : s = 282;
	{8'd228,8'd55} : s = 283;
	{8'd228,8'd56} : s = 284;
	{8'd228,8'd57} : s = 285;
	{8'd228,8'd58} : s = 286;
	{8'd228,8'd59} : s = 287;
	{8'd228,8'd60} : s = 288;
	{8'd228,8'd61} : s = 289;
	{8'd228,8'd62} : s = 290;
	{8'd228,8'd63} : s = 291;
	{8'd228,8'd64} : s = 292;
	{8'd228,8'd65} : s = 293;
	{8'd228,8'd66} : s = 294;
	{8'd228,8'd67} : s = 295;
	{8'd228,8'd68} : s = 296;
	{8'd228,8'd69} : s = 297;
	{8'd228,8'd70} : s = 298;
	{8'd228,8'd71} : s = 299;
	{8'd228,8'd72} : s = 300;
	{8'd228,8'd73} : s = 301;
	{8'd228,8'd74} : s = 302;
	{8'd228,8'd75} : s = 303;
	{8'd228,8'd76} : s = 304;
	{8'd228,8'd77} : s = 305;
	{8'd228,8'd78} : s = 306;
	{8'd228,8'd79} : s = 307;
	{8'd228,8'd80} : s = 308;
	{8'd228,8'd81} : s = 309;
	{8'd228,8'd82} : s = 310;
	{8'd228,8'd83} : s = 311;
	{8'd228,8'd84} : s = 312;
	{8'd228,8'd85} : s = 313;
	{8'd228,8'd86} : s = 314;
	{8'd228,8'd87} : s = 315;
	{8'd228,8'd88} : s = 316;
	{8'd228,8'd89} : s = 317;
	{8'd228,8'd90} : s = 318;
	{8'd228,8'd91} : s = 319;
	{8'd228,8'd92} : s = 320;
	{8'd228,8'd93} : s = 321;
	{8'd228,8'd94} : s = 322;
	{8'd228,8'd95} : s = 323;
	{8'd228,8'd96} : s = 324;
	{8'd228,8'd97} : s = 325;
	{8'd228,8'd98} : s = 326;
	{8'd228,8'd99} : s = 327;
	{8'd228,8'd100} : s = 328;
	{8'd228,8'd101} : s = 329;
	{8'd228,8'd102} : s = 330;
	{8'd228,8'd103} : s = 331;
	{8'd228,8'd104} : s = 332;
	{8'd228,8'd105} : s = 333;
	{8'd228,8'd106} : s = 334;
	{8'd228,8'd107} : s = 335;
	{8'd228,8'd108} : s = 336;
	{8'd228,8'd109} : s = 337;
	{8'd228,8'd110} : s = 338;
	{8'd228,8'd111} : s = 339;
	{8'd228,8'd112} : s = 340;
	{8'd228,8'd113} : s = 341;
	{8'd228,8'd114} : s = 342;
	{8'd228,8'd115} : s = 343;
	{8'd228,8'd116} : s = 344;
	{8'd228,8'd117} : s = 345;
	{8'd228,8'd118} : s = 346;
	{8'd228,8'd119} : s = 347;
	{8'd228,8'd120} : s = 348;
	{8'd228,8'd121} : s = 349;
	{8'd228,8'd122} : s = 350;
	{8'd228,8'd123} : s = 351;
	{8'd228,8'd124} : s = 352;
	{8'd228,8'd125} : s = 353;
	{8'd228,8'd126} : s = 354;
	{8'd228,8'd127} : s = 355;
	{8'd228,8'd128} : s = 356;
	{8'd228,8'd129} : s = 357;
	{8'd228,8'd130} : s = 358;
	{8'd228,8'd131} : s = 359;
	{8'd228,8'd132} : s = 360;
	{8'd228,8'd133} : s = 361;
	{8'd228,8'd134} : s = 362;
	{8'd228,8'd135} : s = 363;
	{8'd228,8'd136} : s = 364;
	{8'd228,8'd137} : s = 365;
	{8'd228,8'd138} : s = 366;
	{8'd228,8'd139} : s = 367;
	{8'd228,8'd140} : s = 368;
	{8'd228,8'd141} : s = 369;
	{8'd228,8'd142} : s = 370;
	{8'd228,8'd143} : s = 371;
	{8'd228,8'd144} : s = 372;
	{8'd228,8'd145} : s = 373;
	{8'd228,8'd146} : s = 374;
	{8'd228,8'd147} : s = 375;
	{8'd228,8'd148} : s = 376;
	{8'd228,8'd149} : s = 377;
	{8'd228,8'd150} : s = 378;
	{8'd228,8'd151} : s = 379;
	{8'd228,8'd152} : s = 380;
	{8'd228,8'd153} : s = 381;
	{8'd228,8'd154} : s = 382;
	{8'd228,8'd155} : s = 383;
	{8'd228,8'd156} : s = 384;
	{8'd228,8'd157} : s = 385;
	{8'd228,8'd158} : s = 386;
	{8'd228,8'd159} : s = 387;
	{8'd228,8'd160} : s = 388;
	{8'd228,8'd161} : s = 389;
	{8'd228,8'd162} : s = 390;
	{8'd228,8'd163} : s = 391;
	{8'd228,8'd164} : s = 392;
	{8'd228,8'd165} : s = 393;
	{8'd228,8'd166} : s = 394;
	{8'd228,8'd167} : s = 395;
	{8'd228,8'd168} : s = 396;
	{8'd228,8'd169} : s = 397;
	{8'd228,8'd170} : s = 398;
	{8'd228,8'd171} : s = 399;
	{8'd228,8'd172} : s = 400;
	{8'd228,8'd173} : s = 401;
	{8'd228,8'd174} : s = 402;
	{8'd228,8'd175} : s = 403;
	{8'd228,8'd176} : s = 404;
	{8'd228,8'd177} : s = 405;
	{8'd228,8'd178} : s = 406;
	{8'd228,8'd179} : s = 407;
	{8'd228,8'd180} : s = 408;
	{8'd228,8'd181} : s = 409;
	{8'd228,8'd182} : s = 410;
	{8'd228,8'd183} : s = 411;
	{8'd228,8'd184} : s = 412;
	{8'd228,8'd185} : s = 413;
	{8'd228,8'd186} : s = 414;
	{8'd228,8'd187} : s = 415;
	{8'd228,8'd188} : s = 416;
	{8'd228,8'd189} : s = 417;
	{8'd228,8'd190} : s = 418;
	{8'd228,8'd191} : s = 419;
	{8'd228,8'd192} : s = 420;
	{8'd228,8'd193} : s = 421;
	{8'd228,8'd194} : s = 422;
	{8'd228,8'd195} : s = 423;
	{8'd228,8'd196} : s = 424;
	{8'd228,8'd197} : s = 425;
	{8'd228,8'd198} : s = 426;
	{8'd228,8'd199} : s = 427;
	{8'd228,8'd200} : s = 428;
	{8'd228,8'd201} : s = 429;
	{8'd228,8'd202} : s = 430;
	{8'd228,8'd203} : s = 431;
	{8'd228,8'd204} : s = 432;
	{8'd228,8'd205} : s = 433;
	{8'd228,8'd206} : s = 434;
	{8'd228,8'd207} : s = 435;
	{8'd228,8'd208} : s = 436;
	{8'd228,8'd209} : s = 437;
	{8'd228,8'd210} : s = 438;
	{8'd228,8'd211} : s = 439;
	{8'd228,8'd212} : s = 440;
	{8'd228,8'd213} : s = 441;
	{8'd228,8'd214} : s = 442;
	{8'd228,8'd215} : s = 443;
	{8'd228,8'd216} : s = 444;
	{8'd228,8'd217} : s = 445;
	{8'd228,8'd218} : s = 446;
	{8'd228,8'd219} : s = 447;
	{8'd228,8'd220} : s = 448;
	{8'd228,8'd221} : s = 449;
	{8'd228,8'd222} : s = 450;
	{8'd228,8'd223} : s = 451;
	{8'd228,8'd224} : s = 452;
	{8'd228,8'd225} : s = 453;
	{8'd228,8'd226} : s = 454;
	{8'd228,8'd227} : s = 455;
	{8'd228,8'd228} : s = 456;
	{8'd228,8'd229} : s = 457;
	{8'd228,8'd230} : s = 458;
	{8'd228,8'd231} : s = 459;
	{8'd228,8'd232} : s = 460;
	{8'd228,8'd233} : s = 461;
	{8'd228,8'd234} : s = 462;
	{8'd228,8'd235} : s = 463;
	{8'd228,8'd236} : s = 464;
	{8'd228,8'd237} : s = 465;
	{8'd228,8'd238} : s = 466;
	{8'd228,8'd239} : s = 467;
	{8'd228,8'd240} : s = 468;
	{8'd228,8'd241} : s = 469;
	{8'd228,8'd242} : s = 470;
	{8'd228,8'd243} : s = 471;
	{8'd228,8'd244} : s = 472;
	{8'd228,8'd245} : s = 473;
	{8'd228,8'd246} : s = 474;
	{8'd228,8'd247} : s = 475;
	{8'd228,8'd248} : s = 476;
	{8'd228,8'd249} : s = 477;
	{8'd228,8'd250} : s = 478;
	{8'd228,8'd251} : s = 479;
	{8'd228,8'd252} : s = 480;
	{8'd228,8'd253} : s = 481;
	{8'd228,8'd254} : s = 482;
	{8'd228,8'd255} : s = 483;
	{8'd229,8'd0} : s = 229;
	{8'd229,8'd1} : s = 230;
	{8'd229,8'd2} : s = 231;
	{8'd229,8'd3} : s = 232;
	{8'd229,8'd4} : s = 233;
	{8'd229,8'd5} : s = 234;
	{8'd229,8'd6} : s = 235;
	{8'd229,8'd7} : s = 236;
	{8'd229,8'd8} : s = 237;
	{8'd229,8'd9} : s = 238;
	{8'd229,8'd10} : s = 239;
	{8'd229,8'd11} : s = 240;
	{8'd229,8'd12} : s = 241;
	{8'd229,8'd13} : s = 242;
	{8'd229,8'd14} : s = 243;
	{8'd229,8'd15} : s = 244;
	{8'd229,8'd16} : s = 245;
	{8'd229,8'd17} : s = 246;
	{8'd229,8'd18} : s = 247;
	{8'd229,8'd19} : s = 248;
	{8'd229,8'd20} : s = 249;
	{8'd229,8'd21} : s = 250;
	{8'd229,8'd22} : s = 251;
	{8'd229,8'd23} : s = 252;
	{8'd229,8'd24} : s = 253;
	{8'd229,8'd25} : s = 254;
	{8'd229,8'd26} : s = 255;
	{8'd229,8'd27} : s = 256;
	{8'd229,8'd28} : s = 257;
	{8'd229,8'd29} : s = 258;
	{8'd229,8'd30} : s = 259;
	{8'd229,8'd31} : s = 260;
	{8'd229,8'd32} : s = 261;
	{8'd229,8'd33} : s = 262;
	{8'd229,8'd34} : s = 263;
	{8'd229,8'd35} : s = 264;
	{8'd229,8'd36} : s = 265;
	{8'd229,8'd37} : s = 266;
	{8'd229,8'd38} : s = 267;
	{8'd229,8'd39} : s = 268;
	{8'd229,8'd40} : s = 269;
	{8'd229,8'd41} : s = 270;
	{8'd229,8'd42} : s = 271;
	{8'd229,8'd43} : s = 272;
	{8'd229,8'd44} : s = 273;
	{8'd229,8'd45} : s = 274;
	{8'd229,8'd46} : s = 275;
	{8'd229,8'd47} : s = 276;
	{8'd229,8'd48} : s = 277;
	{8'd229,8'd49} : s = 278;
	{8'd229,8'd50} : s = 279;
	{8'd229,8'd51} : s = 280;
	{8'd229,8'd52} : s = 281;
	{8'd229,8'd53} : s = 282;
	{8'd229,8'd54} : s = 283;
	{8'd229,8'd55} : s = 284;
	{8'd229,8'd56} : s = 285;
	{8'd229,8'd57} : s = 286;
	{8'd229,8'd58} : s = 287;
	{8'd229,8'd59} : s = 288;
	{8'd229,8'd60} : s = 289;
	{8'd229,8'd61} : s = 290;
	{8'd229,8'd62} : s = 291;
	{8'd229,8'd63} : s = 292;
	{8'd229,8'd64} : s = 293;
	{8'd229,8'd65} : s = 294;
	{8'd229,8'd66} : s = 295;
	{8'd229,8'd67} : s = 296;
	{8'd229,8'd68} : s = 297;
	{8'd229,8'd69} : s = 298;
	{8'd229,8'd70} : s = 299;
	{8'd229,8'd71} : s = 300;
	{8'd229,8'd72} : s = 301;
	{8'd229,8'd73} : s = 302;
	{8'd229,8'd74} : s = 303;
	{8'd229,8'd75} : s = 304;
	{8'd229,8'd76} : s = 305;
	{8'd229,8'd77} : s = 306;
	{8'd229,8'd78} : s = 307;
	{8'd229,8'd79} : s = 308;
	{8'd229,8'd80} : s = 309;
	{8'd229,8'd81} : s = 310;
	{8'd229,8'd82} : s = 311;
	{8'd229,8'd83} : s = 312;
	{8'd229,8'd84} : s = 313;
	{8'd229,8'd85} : s = 314;
	{8'd229,8'd86} : s = 315;
	{8'd229,8'd87} : s = 316;
	{8'd229,8'd88} : s = 317;
	{8'd229,8'd89} : s = 318;
	{8'd229,8'd90} : s = 319;
	{8'd229,8'd91} : s = 320;
	{8'd229,8'd92} : s = 321;
	{8'd229,8'd93} : s = 322;
	{8'd229,8'd94} : s = 323;
	{8'd229,8'd95} : s = 324;
	{8'd229,8'd96} : s = 325;
	{8'd229,8'd97} : s = 326;
	{8'd229,8'd98} : s = 327;
	{8'd229,8'd99} : s = 328;
	{8'd229,8'd100} : s = 329;
	{8'd229,8'd101} : s = 330;
	{8'd229,8'd102} : s = 331;
	{8'd229,8'd103} : s = 332;
	{8'd229,8'd104} : s = 333;
	{8'd229,8'd105} : s = 334;
	{8'd229,8'd106} : s = 335;
	{8'd229,8'd107} : s = 336;
	{8'd229,8'd108} : s = 337;
	{8'd229,8'd109} : s = 338;
	{8'd229,8'd110} : s = 339;
	{8'd229,8'd111} : s = 340;
	{8'd229,8'd112} : s = 341;
	{8'd229,8'd113} : s = 342;
	{8'd229,8'd114} : s = 343;
	{8'd229,8'd115} : s = 344;
	{8'd229,8'd116} : s = 345;
	{8'd229,8'd117} : s = 346;
	{8'd229,8'd118} : s = 347;
	{8'd229,8'd119} : s = 348;
	{8'd229,8'd120} : s = 349;
	{8'd229,8'd121} : s = 350;
	{8'd229,8'd122} : s = 351;
	{8'd229,8'd123} : s = 352;
	{8'd229,8'd124} : s = 353;
	{8'd229,8'd125} : s = 354;
	{8'd229,8'd126} : s = 355;
	{8'd229,8'd127} : s = 356;
	{8'd229,8'd128} : s = 357;
	{8'd229,8'd129} : s = 358;
	{8'd229,8'd130} : s = 359;
	{8'd229,8'd131} : s = 360;
	{8'd229,8'd132} : s = 361;
	{8'd229,8'd133} : s = 362;
	{8'd229,8'd134} : s = 363;
	{8'd229,8'd135} : s = 364;
	{8'd229,8'd136} : s = 365;
	{8'd229,8'd137} : s = 366;
	{8'd229,8'd138} : s = 367;
	{8'd229,8'd139} : s = 368;
	{8'd229,8'd140} : s = 369;
	{8'd229,8'd141} : s = 370;
	{8'd229,8'd142} : s = 371;
	{8'd229,8'd143} : s = 372;
	{8'd229,8'd144} : s = 373;
	{8'd229,8'd145} : s = 374;
	{8'd229,8'd146} : s = 375;
	{8'd229,8'd147} : s = 376;
	{8'd229,8'd148} : s = 377;
	{8'd229,8'd149} : s = 378;
	{8'd229,8'd150} : s = 379;
	{8'd229,8'd151} : s = 380;
	{8'd229,8'd152} : s = 381;
	{8'd229,8'd153} : s = 382;
	{8'd229,8'd154} : s = 383;
	{8'd229,8'd155} : s = 384;
	{8'd229,8'd156} : s = 385;
	{8'd229,8'd157} : s = 386;
	{8'd229,8'd158} : s = 387;
	{8'd229,8'd159} : s = 388;
	{8'd229,8'd160} : s = 389;
	{8'd229,8'd161} : s = 390;
	{8'd229,8'd162} : s = 391;
	{8'd229,8'd163} : s = 392;
	{8'd229,8'd164} : s = 393;
	{8'd229,8'd165} : s = 394;
	{8'd229,8'd166} : s = 395;
	{8'd229,8'd167} : s = 396;
	{8'd229,8'd168} : s = 397;
	{8'd229,8'd169} : s = 398;
	{8'd229,8'd170} : s = 399;
	{8'd229,8'd171} : s = 400;
	{8'd229,8'd172} : s = 401;
	{8'd229,8'd173} : s = 402;
	{8'd229,8'd174} : s = 403;
	{8'd229,8'd175} : s = 404;
	{8'd229,8'd176} : s = 405;
	{8'd229,8'd177} : s = 406;
	{8'd229,8'd178} : s = 407;
	{8'd229,8'd179} : s = 408;
	{8'd229,8'd180} : s = 409;
	{8'd229,8'd181} : s = 410;
	{8'd229,8'd182} : s = 411;
	{8'd229,8'd183} : s = 412;
	{8'd229,8'd184} : s = 413;
	{8'd229,8'd185} : s = 414;
	{8'd229,8'd186} : s = 415;
	{8'd229,8'd187} : s = 416;
	{8'd229,8'd188} : s = 417;
	{8'd229,8'd189} : s = 418;
	{8'd229,8'd190} : s = 419;
	{8'd229,8'd191} : s = 420;
	{8'd229,8'd192} : s = 421;
	{8'd229,8'd193} : s = 422;
	{8'd229,8'd194} : s = 423;
	{8'd229,8'd195} : s = 424;
	{8'd229,8'd196} : s = 425;
	{8'd229,8'd197} : s = 426;
	{8'd229,8'd198} : s = 427;
	{8'd229,8'd199} : s = 428;
	{8'd229,8'd200} : s = 429;
	{8'd229,8'd201} : s = 430;
	{8'd229,8'd202} : s = 431;
	{8'd229,8'd203} : s = 432;
	{8'd229,8'd204} : s = 433;
	{8'd229,8'd205} : s = 434;
	{8'd229,8'd206} : s = 435;
	{8'd229,8'd207} : s = 436;
	{8'd229,8'd208} : s = 437;
	{8'd229,8'd209} : s = 438;
	{8'd229,8'd210} : s = 439;
	{8'd229,8'd211} : s = 440;
	{8'd229,8'd212} : s = 441;
	{8'd229,8'd213} : s = 442;
	{8'd229,8'd214} : s = 443;
	{8'd229,8'd215} : s = 444;
	{8'd229,8'd216} : s = 445;
	{8'd229,8'd217} : s = 446;
	{8'd229,8'd218} : s = 447;
	{8'd229,8'd219} : s = 448;
	{8'd229,8'd220} : s = 449;
	{8'd229,8'd221} : s = 450;
	{8'd229,8'd222} : s = 451;
	{8'd229,8'd223} : s = 452;
	{8'd229,8'd224} : s = 453;
	{8'd229,8'd225} : s = 454;
	{8'd229,8'd226} : s = 455;
	{8'd229,8'd227} : s = 456;
	{8'd229,8'd228} : s = 457;
	{8'd229,8'd229} : s = 458;
	{8'd229,8'd230} : s = 459;
	{8'd229,8'd231} : s = 460;
	{8'd229,8'd232} : s = 461;
	{8'd229,8'd233} : s = 462;
	{8'd229,8'd234} : s = 463;
	{8'd229,8'd235} : s = 464;
	{8'd229,8'd236} : s = 465;
	{8'd229,8'd237} : s = 466;
	{8'd229,8'd238} : s = 467;
	{8'd229,8'd239} : s = 468;
	{8'd229,8'd240} : s = 469;
	{8'd229,8'd241} : s = 470;
	{8'd229,8'd242} : s = 471;
	{8'd229,8'd243} : s = 472;
	{8'd229,8'd244} : s = 473;
	{8'd229,8'd245} : s = 474;
	{8'd229,8'd246} : s = 475;
	{8'd229,8'd247} : s = 476;
	{8'd229,8'd248} : s = 477;
	{8'd229,8'd249} : s = 478;
	{8'd229,8'd250} : s = 479;
	{8'd229,8'd251} : s = 480;
	{8'd229,8'd252} : s = 481;
	{8'd229,8'd253} : s = 482;
	{8'd229,8'd254} : s = 483;
	{8'd229,8'd255} : s = 484;
	{8'd230,8'd0} : s = 230;
	{8'd230,8'd1} : s = 231;
	{8'd230,8'd2} : s = 232;
	{8'd230,8'd3} : s = 233;
	{8'd230,8'd4} : s = 234;
	{8'd230,8'd5} : s = 235;
	{8'd230,8'd6} : s = 236;
	{8'd230,8'd7} : s = 237;
	{8'd230,8'd8} : s = 238;
	{8'd230,8'd9} : s = 239;
	{8'd230,8'd10} : s = 240;
	{8'd230,8'd11} : s = 241;
	{8'd230,8'd12} : s = 242;
	{8'd230,8'd13} : s = 243;
	{8'd230,8'd14} : s = 244;
	{8'd230,8'd15} : s = 245;
	{8'd230,8'd16} : s = 246;
	{8'd230,8'd17} : s = 247;
	{8'd230,8'd18} : s = 248;
	{8'd230,8'd19} : s = 249;
	{8'd230,8'd20} : s = 250;
	{8'd230,8'd21} : s = 251;
	{8'd230,8'd22} : s = 252;
	{8'd230,8'd23} : s = 253;
	{8'd230,8'd24} : s = 254;
	{8'd230,8'd25} : s = 255;
	{8'd230,8'd26} : s = 256;
	{8'd230,8'd27} : s = 257;
	{8'd230,8'd28} : s = 258;
	{8'd230,8'd29} : s = 259;
	{8'd230,8'd30} : s = 260;
	{8'd230,8'd31} : s = 261;
	{8'd230,8'd32} : s = 262;
	{8'd230,8'd33} : s = 263;
	{8'd230,8'd34} : s = 264;
	{8'd230,8'd35} : s = 265;
	{8'd230,8'd36} : s = 266;
	{8'd230,8'd37} : s = 267;
	{8'd230,8'd38} : s = 268;
	{8'd230,8'd39} : s = 269;
	{8'd230,8'd40} : s = 270;
	{8'd230,8'd41} : s = 271;
	{8'd230,8'd42} : s = 272;
	{8'd230,8'd43} : s = 273;
	{8'd230,8'd44} : s = 274;
	{8'd230,8'd45} : s = 275;
	{8'd230,8'd46} : s = 276;
	{8'd230,8'd47} : s = 277;
	{8'd230,8'd48} : s = 278;
	{8'd230,8'd49} : s = 279;
	{8'd230,8'd50} : s = 280;
	{8'd230,8'd51} : s = 281;
	{8'd230,8'd52} : s = 282;
	{8'd230,8'd53} : s = 283;
	{8'd230,8'd54} : s = 284;
	{8'd230,8'd55} : s = 285;
	{8'd230,8'd56} : s = 286;
	{8'd230,8'd57} : s = 287;
	{8'd230,8'd58} : s = 288;
	{8'd230,8'd59} : s = 289;
	{8'd230,8'd60} : s = 290;
	{8'd230,8'd61} : s = 291;
	{8'd230,8'd62} : s = 292;
	{8'd230,8'd63} : s = 293;
	{8'd230,8'd64} : s = 294;
	{8'd230,8'd65} : s = 295;
	{8'd230,8'd66} : s = 296;
	{8'd230,8'd67} : s = 297;
	{8'd230,8'd68} : s = 298;
	{8'd230,8'd69} : s = 299;
	{8'd230,8'd70} : s = 300;
	{8'd230,8'd71} : s = 301;
	{8'd230,8'd72} : s = 302;
	{8'd230,8'd73} : s = 303;
	{8'd230,8'd74} : s = 304;
	{8'd230,8'd75} : s = 305;
	{8'd230,8'd76} : s = 306;
	{8'd230,8'd77} : s = 307;
	{8'd230,8'd78} : s = 308;
	{8'd230,8'd79} : s = 309;
	{8'd230,8'd80} : s = 310;
	{8'd230,8'd81} : s = 311;
	{8'd230,8'd82} : s = 312;
	{8'd230,8'd83} : s = 313;
	{8'd230,8'd84} : s = 314;
	{8'd230,8'd85} : s = 315;
	{8'd230,8'd86} : s = 316;
	{8'd230,8'd87} : s = 317;
	{8'd230,8'd88} : s = 318;
	{8'd230,8'd89} : s = 319;
	{8'd230,8'd90} : s = 320;
	{8'd230,8'd91} : s = 321;
	{8'd230,8'd92} : s = 322;
	{8'd230,8'd93} : s = 323;
	{8'd230,8'd94} : s = 324;
	{8'd230,8'd95} : s = 325;
	{8'd230,8'd96} : s = 326;
	{8'd230,8'd97} : s = 327;
	{8'd230,8'd98} : s = 328;
	{8'd230,8'd99} : s = 329;
	{8'd230,8'd100} : s = 330;
	{8'd230,8'd101} : s = 331;
	{8'd230,8'd102} : s = 332;
	{8'd230,8'd103} : s = 333;
	{8'd230,8'd104} : s = 334;
	{8'd230,8'd105} : s = 335;
	{8'd230,8'd106} : s = 336;
	{8'd230,8'd107} : s = 337;
	{8'd230,8'd108} : s = 338;
	{8'd230,8'd109} : s = 339;
	{8'd230,8'd110} : s = 340;
	{8'd230,8'd111} : s = 341;
	{8'd230,8'd112} : s = 342;
	{8'd230,8'd113} : s = 343;
	{8'd230,8'd114} : s = 344;
	{8'd230,8'd115} : s = 345;
	{8'd230,8'd116} : s = 346;
	{8'd230,8'd117} : s = 347;
	{8'd230,8'd118} : s = 348;
	{8'd230,8'd119} : s = 349;
	{8'd230,8'd120} : s = 350;
	{8'd230,8'd121} : s = 351;
	{8'd230,8'd122} : s = 352;
	{8'd230,8'd123} : s = 353;
	{8'd230,8'd124} : s = 354;
	{8'd230,8'd125} : s = 355;
	{8'd230,8'd126} : s = 356;
	{8'd230,8'd127} : s = 357;
	{8'd230,8'd128} : s = 358;
	{8'd230,8'd129} : s = 359;
	{8'd230,8'd130} : s = 360;
	{8'd230,8'd131} : s = 361;
	{8'd230,8'd132} : s = 362;
	{8'd230,8'd133} : s = 363;
	{8'd230,8'd134} : s = 364;
	{8'd230,8'd135} : s = 365;
	{8'd230,8'd136} : s = 366;
	{8'd230,8'd137} : s = 367;
	{8'd230,8'd138} : s = 368;
	{8'd230,8'd139} : s = 369;
	{8'd230,8'd140} : s = 370;
	{8'd230,8'd141} : s = 371;
	{8'd230,8'd142} : s = 372;
	{8'd230,8'd143} : s = 373;
	{8'd230,8'd144} : s = 374;
	{8'd230,8'd145} : s = 375;
	{8'd230,8'd146} : s = 376;
	{8'd230,8'd147} : s = 377;
	{8'd230,8'd148} : s = 378;
	{8'd230,8'd149} : s = 379;
	{8'd230,8'd150} : s = 380;
	{8'd230,8'd151} : s = 381;
	{8'd230,8'd152} : s = 382;
	{8'd230,8'd153} : s = 383;
	{8'd230,8'd154} : s = 384;
	{8'd230,8'd155} : s = 385;
	{8'd230,8'd156} : s = 386;
	{8'd230,8'd157} : s = 387;
	{8'd230,8'd158} : s = 388;
	{8'd230,8'd159} : s = 389;
	{8'd230,8'd160} : s = 390;
	{8'd230,8'd161} : s = 391;
	{8'd230,8'd162} : s = 392;
	{8'd230,8'd163} : s = 393;
	{8'd230,8'd164} : s = 394;
	{8'd230,8'd165} : s = 395;
	{8'd230,8'd166} : s = 396;
	{8'd230,8'd167} : s = 397;
	{8'd230,8'd168} : s = 398;
	{8'd230,8'd169} : s = 399;
	{8'd230,8'd170} : s = 400;
	{8'd230,8'd171} : s = 401;
	{8'd230,8'd172} : s = 402;
	{8'd230,8'd173} : s = 403;
	{8'd230,8'd174} : s = 404;
	{8'd230,8'd175} : s = 405;
	{8'd230,8'd176} : s = 406;
	{8'd230,8'd177} : s = 407;
	{8'd230,8'd178} : s = 408;
	{8'd230,8'd179} : s = 409;
	{8'd230,8'd180} : s = 410;
	{8'd230,8'd181} : s = 411;
	{8'd230,8'd182} : s = 412;
	{8'd230,8'd183} : s = 413;
	{8'd230,8'd184} : s = 414;
	{8'd230,8'd185} : s = 415;
	{8'd230,8'd186} : s = 416;
	{8'd230,8'd187} : s = 417;
	{8'd230,8'd188} : s = 418;
	{8'd230,8'd189} : s = 419;
	{8'd230,8'd190} : s = 420;
	{8'd230,8'd191} : s = 421;
	{8'd230,8'd192} : s = 422;
	{8'd230,8'd193} : s = 423;
	{8'd230,8'd194} : s = 424;
	{8'd230,8'd195} : s = 425;
	{8'd230,8'd196} : s = 426;
	{8'd230,8'd197} : s = 427;
	{8'd230,8'd198} : s = 428;
	{8'd230,8'd199} : s = 429;
	{8'd230,8'd200} : s = 430;
	{8'd230,8'd201} : s = 431;
	{8'd230,8'd202} : s = 432;
	{8'd230,8'd203} : s = 433;
	{8'd230,8'd204} : s = 434;
	{8'd230,8'd205} : s = 435;
	{8'd230,8'd206} : s = 436;
	{8'd230,8'd207} : s = 437;
	{8'd230,8'd208} : s = 438;
	{8'd230,8'd209} : s = 439;
	{8'd230,8'd210} : s = 440;
	{8'd230,8'd211} : s = 441;
	{8'd230,8'd212} : s = 442;
	{8'd230,8'd213} : s = 443;
	{8'd230,8'd214} : s = 444;
	{8'd230,8'd215} : s = 445;
	{8'd230,8'd216} : s = 446;
	{8'd230,8'd217} : s = 447;
	{8'd230,8'd218} : s = 448;
	{8'd230,8'd219} : s = 449;
	{8'd230,8'd220} : s = 450;
	{8'd230,8'd221} : s = 451;
	{8'd230,8'd222} : s = 452;
	{8'd230,8'd223} : s = 453;
	{8'd230,8'd224} : s = 454;
	{8'd230,8'd225} : s = 455;
	{8'd230,8'd226} : s = 456;
	{8'd230,8'd227} : s = 457;
	{8'd230,8'd228} : s = 458;
	{8'd230,8'd229} : s = 459;
	{8'd230,8'd230} : s = 460;
	{8'd230,8'd231} : s = 461;
	{8'd230,8'd232} : s = 462;
	{8'd230,8'd233} : s = 463;
	{8'd230,8'd234} : s = 464;
	{8'd230,8'd235} : s = 465;
	{8'd230,8'd236} : s = 466;
	{8'd230,8'd237} : s = 467;
	{8'd230,8'd238} : s = 468;
	{8'd230,8'd239} : s = 469;
	{8'd230,8'd240} : s = 470;
	{8'd230,8'd241} : s = 471;
	{8'd230,8'd242} : s = 472;
	{8'd230,8'd243} : s = 473;
	{8'd230,8'd244} : s = 474;
	{8'd230,8'd245} : s = 475;
	{8'd230,8'd246} : s = 476;
	{8'd230,8'd247} : s = 477;
	{8'd230,8'd248} : s = 478;
	{8'd230,8'd249} : s = 479;
	{8'd230,8'd250} : s = 480;
	{8'd230,8'd251} : s = 481;
	{8'd230,8'd252} : s = 482;
	{8'd230,8'd253} : s = 483;
	{8'd230,8'd254} : s = 484;
	{8'd230,8'd255} : s = 485;
	{8'd231,8'd0} : s = 231;
	{8'd231,8'd1} : s = 232;
	{8'd231,8'd2} : s = 233;
	{8'd231,8'd3} : s = 234;
	{8'd231,8'd4} : s = 235;
	{8'd231,8'd5} : s = 236;
	{8'd231,8'd6} : s = 237;
	{8'd231,8'd7} : s = 238;
	{8'd231,8'd8} : s = 239;
	{8'd231,8'd9} : s = 240;
	{8'd231,8'd10} : s = 241;
	{8'd231,8'd11} : s = 242;
	{8'd231,8'd12} : s = 243;
	{8'd231,8'd13} : s = 244;
	{8'd231,8'd14} : s = 245;
	{8'd231,8'd15} : s = 246;
	{8'd231,8'd16} : s = 247;
	{8'd231,8'd17} : s = 248;
	{8'd231,8'd18} : s = 249;
	{8'd231,8'd19} : s = 250;
	{8'd231,8'd20} : s = 251;
	{8'd231,8'd21} : s = 252;
	{8'd231,8'd22} : s = 253;
	{8'd231,8'd23} : s = 254;
	{8'd231,8'd24} : s = 255;
	{8'd231,8'd25} : s = 256;
	{8'd231,8'd26} : s = 257;
	{8'd231,8'd27} : s = 258;
	{8'd231,8'd28} : s = 259;
	{8'd231,8'd29} : s = 260;
	{8'd231,8'd30} : s = 261;
	{8'd231,8'd31} : s = 262;
	{8'd231,8'd32} : s = 263;
	{8'd231,8'd33} : s = 264;
	{8'd231,8'd34} : s = 265;
	{8'd231,8'd35} : s = 266;
	{8'd231,8'd36} : s = 267;
	{8'd231,8'd37} : s = 268;
	{8'd231,8'd38} : s = 269;
	{8'd231,8'd39} : s = 270;
	{8'd231,8'd40} : s = 271;
	{8'd231,8'd41} : s = 272;
	{8'd231,8'd42} : s = 273;
	{8'd231,8'd43} : s = 274;
	{8'd231,8'd44} : s = 275;
	{8'd231,8'd45} : s = 276;
	{8'd231,8'd46} : s = 277;
	{8'd231,8'd47} : s = 278;
	{8'd231,8'd48} : s = 279;
	{8'd231,8'd49} : s = 280;
	{8'd231,8'd50} : s = 281;
	{8'd231,8'd51} : s = 282;
	{8'd231,8'd52} : s = 283;
	{8'd231,8'd53} : s = 284;
	{8'd231,8'd54} : s = 285;
	{8'd231,8'd55} : s = 286;
	{8'd231,8'd56} : s = 287;
	{8'd231,8'd57} : s = 288;
	{8'd231,8'd58} : s = 289;
	{8'd231,8'd59} : s = 290;
	{8'd231,8'd60} : s = 291;
	{8'd231,8'd61} : s = 292;
	{8'd231,8'd62} : s = 293;
	{8'd231,8'd63} : s = 294;
	{8'd231,8'd64} : s = 295;
	{8'd231,8'd65} : s = 296;
	{8'd231,8'd66} : s = 297;
	{8'd231,8'd67} : s = 298;
	{8'd231,8'd68} : s = 299;
	{8'd231,8'd69} : s = 300;
	{8'd231,8'd70} : s = 301;
	{8'd231,8'd71} : s = 302;
	{8'd231,8'd72} : s = 303;
	{8'd231,8'd73} : s = 304;
	{8'd231,8'd74} : s = 305;
	{8'd231,8'd75} : s = 306;
	{8'd231,8'd76} : s = 307;
	{8'd231,8'd77} : s = 308;
	{8'd231,8'd78} : s = 309;
	{8'd231,8'd79} : s = 310;
	{8'd231,8'd80} : s = 311;
	{8'd231,8'd81} : s = 312;
	{8'd231,8'd82} : s = 313;
	{8'd231,8'd83} : s = 314;
	{8'd231,8'd84} : s = 315;
	{8'd231,8'd85} : s = 316;
	{8'd231,8'd86} : s = 317;
	{8'd231,8'd87} : s = 318;
	{8'd231,8'd88} : s = 319;
	{8'd231,8'd89} : s = 320;
	{8'd231,8'd90} : s = 321;
	{8'd231,8'd91} : s = 322;
	{8'd231,8'd92} : s = 323;
	{8'd231,8'd93} : s = 324;
	{8'd231,8'd94} : s = 325;
	{8'd231,8'd95} : s = 326;
	{8'd231,8'd96} : s = 327;
	{8'd231,8'd97} : s = 328;
	{8'd231,8'd98} : s = 329;
	{8'd231,8'd99} : s = 330;
	{8'd231,8'd100} : s = 331;
	{8'd231,8'd101} : s = 332;
	{8'd231,8'd102} : s = 333;
	{8'd231,8'd103} : s = 334;
	{8'd231,8'd104} : s = 335;
	{8'd231,8'd105} : s = 336;
	{8'd231,8'd106} : s = 337;
	{8'd231,8'd107} : s = 338;
	{8'd231,8'd108} : s = 339;
	{8'd231,8'd109} : s = 340;
	{8'd231,8'd110} : s = 341;
	{8'd231,8'd111} : s = 342;
	{8'd231,8'd112} : s = 343;
	{8'd231,8'd113} : s = 344;
	{8'd231,8'd114} : s = 345;
	{8'd231,8'd115} : s = 346;
	{8'd231,8'd116} : s = 347;
	{8'd231,8'd117} : s = 348;
	{8'd231,8'd118} : s = 349;
	{8'd231,8'd119} : s = 350;
	{8'd231,8'd120} : s = 351;
	{8'd231,8'd121} : s = 352;
	{8'd231,8'd122} : s = 353;
	{8'd231,8'd123} : s = 354;
	{8'd231,8'd124} : s = 355;
	{8'd231,8'd125} : s = 356;
	{8'd231,8'd126} : s = 357;
	{8'd231,8'd127} : s = 358;
	{8'd231,8'd128} : s = 359;
	{8'd231,8'd129} : s = 360;
	{8'd231,8'd130} : s = 361;
	{8'd231,8'd131} : s = 362;
	{8'd231,8'd132} : s = 363;
	{8'd231,8'd133} : s = 364;
	{8'd231,8'd134} : s = 365;
	{8'd231,8'd135} : s = 366;
	{8'd231,8'd136} : s = 367;
	{8'd231,8'd137} : s = 368;
	{8'd231,8'd138} : s = 369;
	{8'd231,8'd139} : s = 370;
	{8'd231,8'd140} : s = 371;
	{8'd231,8'd141} : s = 372;
	{8'd231,8'd142} : s = 373;
	{8'd231,8'd143} : s = 374;
	{8'd231,8'd144} : s = 375;
	{8'd231,8'd145} : s = 376;
	{8'd231,8'd146} : s = 377;
	{8'd231,8'd147} : s = 378;
	{8'd231,8'd148} : s = 379;
	{8'd231,8'd149} : s = 380;
	{8'd231,8'd150} : s = 381;
	{8'd231,8'd151} : s = 382;
	{8'd231,8'd152} : s = 383;
	{8'd231,8'd153} : s = 384;
	{8'd231,8'd154} : s = 385;
	{8'd231,8'd155} : s = 386;
	{8'd231,8'd156} : s = 387;
	{8'd231,8'd157} : s = 388;
	{8'd231,8'd158} : s = 389;
	{8'd231,8'd159} : s = 390;
	{8'd231,8'd160} : s = 391;
	{8'd231,8'd161} : s = 392;
	{8'd231,8'd162} : s = 393;
	{8'd231,8'd163} : s = 394;
	{8'd231,8'd164} : s = 395;
	{8'd231,8'd165} : s = 396;
	{8'd231,8'd166} : s = 397;
	{8'd231,8'd167} : s = 398;
	{8'd231,8'd168} : s = 399;
	{8'd231,8'd169} : s = 400;
	{8'd231,8'd170} : s = 401;
	{8'd231,8'd171} : s = 402;
	{8'd231,8'd172} : s = 403;
	{8'd231,8'd173} : s = 404;
	{8'd231,8'd174} : s = 405;
	{8'd231,8'd175} : s = 406;
	{8'd231,8'd176} : s = 407;
	{8'd231,8'd177} : s = 408;
	{8'd231,8'd178} : s = 409;
	{8'd231,8'd179} : s = 410;
	{8'd231,8'd180} : s = 411;
	{8'd231,8'd181} : s = 412;
	{8'd231,8'd182} : s = 413;
	{8'd231,8'd183} : s = 414;
	{8'd231,8'd184} : s = 415;
	{8'd231,8'd185} : s = 416;
	{8'd231,8'd186} : s = 417;
	{8'd231,8'd187} : s = 418;
	{8'd231,8'd188} : s = 419;
	{8'd231,8'd189} : s = 420;
	{8'd231,8'd190} : s = 421;
	{8'd231,8'd191} : s = 422;
	{8'd231,8'd192} : s = 423;
	{8'd231,8'd193} : s = 424;
	{8'd231,8'd194} : s = 425;
	{8'd231,8'd195} : s = 426;
	{8'd231,8'd196} : s = 427;
	{8'd231,8'd197} : s = 428;
	{8'd231,8'd198} : s = 429;
	{8'd231,8'd199} : s = 430;
	{8'd231,8'd200} : s = 431;
	{8'd231,8'd201} : s = 432;
	{8'd231,8'd202} : s = 433;
	{8'd231,8'd203} : s = 434;
	{8'd231,8'd204} : s = 435;
	{8'd231,8'd205} : s = 436;
	{8'd231,8'd206} : s = 437;
	{8'd231,8'd207} : s = 438;
	{8'd231,8'd208} : s = 439;
	{8'd231,8'd209} : s = 440;
	{8'd231,8'd210} : s = 441;
	{8'd231,8'd211} : s = 442;
	{8'd231,8'd212} : s = 443;
	{8'd231,8'd213} : s = 444;
	{8'd231,8'd214} : s = 445;
	{8'd231,8'd215} : s = 446;
	{8'd231,8'd216} : s = 447;
	{8'd231,8'd217} : s = 448;
	{8'd231,8'd218} : s = 449;
	{8'd231,8'd219} : s = 450;
	{8'd231,8'd220} : s = 451;
	{8'd231,8'd221} : s = 452;
	{8'd231,8'd222} : s = 453;
	{8'd231,8'd223} : s = 454;
	{8'd231,8'd224} : s = 455;
	{8'd231,8'd225} : s = 456;
	{8'd231,8'd226} : s = 457;
	{8'd231,8'd227} : s = 458;
	{8'd231,8'd228} : s = 459;
	{8'd231,8'd229} : s = 460;
	{8'd231,8'd230} : s = 461;
	{8'd231,8'd231} : s = 462;
	{8'd231,8'd232} : s = 463;
	{8'd231,8'd233} : s = 464;
	{8'd231,8'd234} : s = 465;
	{8'd231,8'd235} : s = 466;
	{8'd231,8'd236} : s = 467;
	{8'd231,8'd237} : s = 468;
	{8'd231,8'd238} : s = 469;
	{8'd231,8'd239} : s = 470;
	{8'd231,8'd240} : s = 471;
	{8'd231,8'd241} : s = 472;
	{8'd231,8'd242} : s = 473;
	{8'd231,8'd243} : s = 474;
	{8'd231,8'd244} : s = 475;
	{8'd231,8'd245} : s = 476;
	{8'd231,8'd246} : s = 477;
	{8'd231,8'd247} : s = 478;
	{8'd231,8'd248} : s = 479;
	{8'd231,8'd249} : s = 480;
	{8'd231,8'd250} : s = 481;
	{8'd231,8'd251} : s = 482;
	{8'd231,8'd252} : s = 483;
	{8'd231,8'd253} : s = 484;
	{8'd231,8'd254} : s = 485;
	{8'd231,8'd255} : s = 486;
	{8'd232,8'd0} : s = 232;
	{8'd232,8'd1} : s = 233;
	{8'd232,8'd2} : s = 234;
	{8'd232,8'd3} : s = 235;
	{8'd232,8'd4} : s = 236;
	{8'd232,8'd5} : s = 237;
	{8'd232,8'd6} : s = 238;
	{8'd232,8'd7} : s = 239;
	{8'd232,8'd8} : s = 240;
	{8'd232,8'd9} : s = 241;
	{8'd232,8'd10} : s = 242;
	{8'd232,8'd11} : s = 243;
	{8'd232,8'd12} : s = 244;
	{8'd232,8'd13} : s = 245;
	{8'd232,8'd14} : s = 246;
	{8'd232,8'd15} : s = 247;
	{8'd232,8'd16} : s = 248;
	{8'd232,8'd17} : s = 249;
	{8'd232,8'd18} : s = 250;
	{8'd232,8'd19} : s = 251;
	{8'd232,8'd20} : s = 252;
	{8'd232,8'd21} : s = 253;
	{8'd232,8'd22} : s = 254;
	{8'd232,8'd23} : s = 255;
	{8'd232,8'd24} : s = 256;
	{8'd232,8'd25} : s = 257;
	{8'd232,8'd26} : s = 258;
	{8'd232,8'd27} : s = 259;
	{8'd232,8'd28} : s = 260;
	{8'd232,8'd29} : s = 261;
	{8'd232,8'd30} : s = 262;
	{8'd232,8'd31} : s = 263;
	{8'd232,8'd32} : s = 264;
	{8'd232,8'd33} : s = 265;
	{8'd232,8'd34} : s = 266;
	{8'd232,8'd35} : s = 267;
	{8'd232,8'd36} : s = 268;
	{8'd232,8'd37} : s = 269;
	{8'd232,8'd38} : s = 270;
	{8'd232,8'd39} : s = 271;
	{8'd232,8'd40} : s = 272;
	{8'd232,8'd41} : s = 273;
	{8'd232,8'd42} : s = 274;
	{8'd232,8'd43} : s = 275;
	{8'd232,8'd44} : s = 276;
	{8'd232,8'd45} : s = 277;
	{8'd232,8'd46} : s = 278;
	{8'd232,8'd47} : s = 279;
	{8'd232,8'd48} : s = 280;
	{8'd232,8'd49} : s = 281;
	{8'd232,8'd50} : s = 282;
	{8'd232,8'd51} : s = 283;
	{8'd232,8'd52} : s = 284;
	{8'd232,8'd53} : s = 285;
	{8'd232,8'd54} : s = 286;
	{8'd232,8'd55} : s = 287;
	{8'd232,8'd56} : s = 288;
	{8'd232,8'd57} : s = 289;
	{8'd232,8'd58} : s = 290;
	{8'd232,8'd59} : s = 291;
	{8'd232,8'd60} : s = 292;
	{8'd232,8'd61} : s = 293;
	{8'd232,8'd62} : s = 294;
	{8'd232,8'd63} : s = 295;
	{8'd232,8'd64} : s = 296;
	{8'd232,8'd65} : s = 297;
	{8'd232,8'd66} : s = 298;
	{8'd232,8'd67} : s = 299;
	{8'd232,8'd68} : s = 300;
	{8'd232,8'd69} : s = 301;
	{8'd232,8'd70} : s = 302;
	{8'd232,8'd71} : s = 303;
	{8'd232,8'd72} : s = 304;
	{8'd232,8'd73} : s = 305;
	{8'd232,8'd74} : s = 306;
	{8'd232,8'd75} : s = 307;
	{8'd232,8'd76} : s = 308;
	{8'd232,8'd77} : s = 309;
	{8'd232,8'd78} : s = 310;
	{8'd232,8'd79} : s = 311;
	{8'd232,8'd80} : s = 312;
	{8'd232,8'd81} : s = 313;
	{8'd232,8'd82} : s = 314;
	{8'd232,8'd83} : s = 315;
	{8'd232,8'd84} : s = 316;
	{8'd232,8'd85} : s = 317;
	{8'd232,8'd86} : s = 318;
	{8'd232,8'd87} : s = 319;
	{8'd232,8'd88} : s = 320;
	{8'd232,8'd89} : s = 321;
	{8'd232,8'd90} : s = 322;
	{8'd232,8'd91} : s = 323;
	{8'd232,8'd92} : s = 324;
	{8'd232,8'd93} : s = 325;
	{8'd232,8'd94} : s = 326;
	{8'd232,8'd95} : s = 327;
	{8'd232,8'd96} : s = 328;
	{8'd232,8'd97} : s = 329;
	{8'd232,8'd98} : s = 330;
	{8'd232,8'd99} : s = 331;
	{8'd232,8'd100} : s = 332;
	{8'd232,8'd101} : s = 333;
	{8'd232,8'd102} : s = 334;
	{8'd232,8'd103} : s = 335;
	{8'd232,8'd104} : s = 336;
	{8'd232,8'd105} : s = 337;
	{8'd232,8'd106} : s = 338;
	{8'd232,8'd107} : s = 339;
	{8'd232,8'd108} : s = 340;
	{8'd232,8'd109} : s = 341;
	{8'd232,8'd110} : s = 342;
	{8'd232,8'd111} : s = 343;
	{8'd232,8'd112} : s = 344;
	{8'd232,8'd113} : s = 345;
	{8'd232,8'd114} : s = 346;
	{8'd232,8'd115} : s = 347;
	{8'd232,8'd116} : s = 348;
	{8'd232,8'd117} : s = 349;
	{8'd232,8'd118} : s = 350;
	{8'd232,8'd119} : s = 351;
	{8'd232,8'd120} : s = 352;
	{8'd232,8'd121} : s = 353;
	{8'd232,8'd122} : s = 354;
	{8'd232,8'd123} : s = 355;
	{8'd232,8'd124} : s = 356;
	{8'd232,8'd125} : s = 357;
	{8'd232,8'd126} : s = 358;
	{8'd232,8'd127} : s = 359;
	{8'd232,8'd128} : s = 360;
	{8'd232,8'd129} : s = 361;
	{8'd232,8'd130} : s = 362;
	{8'd232,8'd131} : s = 363;
	{8'd232,8'd132} : s = 364;
	{8'd232,8'd133} : s = 365;
	{8'd232,8'd134} : s = 366;
	{8'd232,8'd135} : s = 367;
	{8'd232,8'd136} : s = 368;
	{8'd232,8'd137} : s = 369;
	{8'd232,8'd138} : s = 370;
	{8'd232,8'd139} : s = 371;
	{8'd232,8'd140} : s = 372;
	{8'd232,8'd141} : s = 373;
	{8'd232,8'd142} : s = 374;
	{8'd232,8'd143} : s = 375;
	{8'd232,8'd144} : s = 376;
	{8'd232,8'd145} : s = 377;
	{8'd232,8'd146} : s = 378;
	{8'd232,8'd147} : s = 379;
	{8'd232,8'd148} : s = 380;
	{8'd232,8'd149} : s = 381;
	{8'd232,8'd150} : s = 382;
	{8'd232,8'd151} : s = 383;
	{8'd232,8'd152} : s = 384;
	{8'd232,8'd153} : s = 385;
	{8'd232,8'd154} : s = 386;
	{8'd232,8'd155} : s = 387;
	{8'd232,8'd156} : s = 388;
	{8'd232,8'd157} : s = 389;
	{8'd232,8'd158} : s = 390;
	{8'd232,8'd159} : s = 391;
	{8'd232,8'd160} : s = 392;
	{8'd232,8'd161} : s = 393;
	{8'd232,8'd162} : s = 394;
	{8'd232,8'd163} : s = 395;
	{8'd232,8'd164} : s = 396;
	{8'd232,8'd165} : s = 397;
	{8'd232,8'd166} : s = 398;
	{8'd232,8'd167} : s = 399;
	{8'd232,8'd168} : s = 400;
	{8'd232,8'd169} : s = 401;
	{8'd232,8'd170} : s = 402;
	{8'd232,8'd171} : s = 403;
	{8'd232,8'd172} : s = 404;
	{8'd232,8'd173} : s = 405;
	{8'd232,8'd174} : s = 406;
	{8'd232,8'd175} : s = 407;
	{8'd232,8'd176} : s = 408;
	{8'd232,8'd177} : s = 409;
	{8'd232,8'd178} : s = 410;
	{8'd232,8'd179} : s = 411;
	{8'd232,8'd180} : s = 412;
	{8'd232,8'd181} : s = 413;
	{8'd232,8'd182} : s = 414;
	{8'd232,8'd183} : s = 415;
	{8'd232,8'd184} : s = 416;
	{8'd232,8'd185} : s = 417;
	{8'd232,8'd186} : s = 418;
	{8'd232,8'd187} : s = 419;
	{8'd232,8'd188} : s = 420;
	{8'd232,8'd189} : s = 421;
	{8'd232,8'd190} : s = 422;
	{8'd232,8'd191} : s = 423;
	{8'd232,8'd192} : s = 424;
	{8'd232,8'd193} : s = 425;
	{8'd232,8'd194} : s = 426;
	{8'd232,8'd195} : s = 427;
	{8'd232,8'd196} : s = 428;
	{8'd232,8'd197} : s = 429;
	{8'd232,8'd198} : s = 430;
	{8'd232,8'd199} : s = 431;
	{8'd232,8'd200} : s = 432;
	{8'd232,8'd201} : s = 433;
	{8'd232,8'd202} : s = 434;
	{8'd232,8'd203} : s = 435;
	{8'd232,8'd204} : s = 436;
	{8'd232,8'd205} : s = 437;
	{8'd232,8'd206} : s = 438;
	{8'd232,8'd207} : s = 439;
	{8'd232,8'd208} : s = 440;
	{8'd232,8'd209} : s = 441;
	{8'd232,8'd210} : s = 442;
	{8'd232,8'd211} : s = 443;
	{8'd232,8'd212} : s = 444;
	{8'd232,8'd213} : s = 445;
	{8'd232,8'd214} : s = 446;
	{8'd232,8'd215} : s = 447;
	{8'd232,8'd216} : s = 448;
	{8'd232,8'd217} : s = 449;
	{8'd232,8'd218} : s = 450;
	{8'd232,8'd219} : s = 451;
	{8'd232,8'd220} : s = 452;
	{8'd232,8'd221} : s = 453;
	{8'd232,8'd222} : s = 454;
	{8'd232,8'd223} : s = 455;
	{8'd232,8'd224} : s = 456;
	{8'd232,8'd225} : s = 457;
	{8'd232,8'd226} : s = 458;
	{8'd232,8'd227} : s = 459;
	{8'd232,8'd228} : s = 460;
	{8'd232,8'd229} : s = 461;
	{8'd232,8'd230} : s = 462;
	{8'd232,8'd231} : s = 463;
	{8'd232,8'd232} : s = 464;
	{8'd232,8'd233} : s = 465;
	{8'd232,8'd234} : s = 466;
	{8'd232,8'd235} : s = 467;
	{8'd232,8'd236} : s = 468;
	{8'd232,8'd237} : s = 469;
	{8'd232,8'd238} : s = 470;
	{8'd232,8'd239} : s = 471;
	{8'd232,8'd240} : s = 472;
	{8'd232,8'd241} : s = 473;
	{8'd232,8'd242} : s = 474;
	{8'd232,8'd243} : s = 475;
	{8'd232,8'd244} : s = 476;
	{8'd232,8'd245} : s = 477;
	{8'd232,8'd246} : s = 478;
	{8'd232,8'd247} : s = 479;
	{8'd232,8'd248} : s = 480;
	{8'd232,8'd249} : s = 481;
	{8'd232,8'd250} : s = 482;
	{8'd232,8'd251} : s = 483;
	{8'd232,8'd252} : s = 484;
	{8'd232,8'd253} : s = 485;
	{8'd232,8'd254} : s = 486;
	{8'd232,8'd255} : s = 487;
	{8'd233,8'd0} : s = 233;
	{8'd233,8'd1} : s = 234;
	{8'd233,8'd2} : s = 235;
	{8'd233,8'd3} : s = 236;
	{8'd233,8'd4} : s = 237;
	{8'd233,8'd5} : s = 238;
	{8'd233,8'd6} : s = 239;
	{8'd233,8'd7} : s = 240;
	{8'd233,8'd8} : s = 241;
	{8'd233,8'd9} : s = 242;
	{8'd233,8'd10} : s = 243;
	{8'd233,8'd11} : s = 244;
	{8'd233,8'd12} : s = 245;
	{8'd233,8'd13} : s = 246;
	{8'd233,8'd14} : s = 247;
	{8'd233,8'd15} : s = 248;
	{8'd233,8'd16} : s = 249;
	{8'd233,8'd17} : s = 250;
	{8'd233,8'd18} : s = 251;
	{8'd233,8'd19} : s = 252;
	{8'd233,8'd20} : s = 253;
	{8'd233,8'd21} : s = 254;
	{8'd233,8'd22} : s = 255;
	{8'd233,8'd23} : s = 256;
	{8'd233,8'd24} : s = 257;
	{8'd233,8'd25} : s = 258;
	{8'd233,8'd26} : s = 259;
	{8'd233,8'd27} : s = 260;
	{8'd233,8'd28} : s = 261;
	{8'd233,8'd29} : s = 262;
	{8'd233,8'd30} : s = 263;
	{8'd233,8'd31} : s = 264;
	{8'd233,8'd32} : s = 265;
	{8'd233,8'd33} : s = 266;
	{8'd233,8'd34} : s = 267;
	{8'd233,8'd35} : s = 268;
	{8'd233,8'd36} : s = 269;
	{8'd233,8'd37} : s = 270;
	{8'd233,8'd38} : s = 271;
	{8'd233,8'd39} : s = 272;
	{8'd233,8'd40} : s = 273;
	{8'd233,8'd41} : s = 274;
	{8'd233,8'd42} : s = 275;
	{8'd233,8'd43} : s = 276;
	{8'd233,8'd44} : s = 277;
	{8'd233,8'd45} : s = 278;
	{8'd233,8'd46} : s = 279;
	{8'd233,8'd47} : s = 280;
	{8'd233,8'd48} : s = 281;
	{8'd233,8'd49} : s = 282;
	{8'd233,8'd50} : s = 283;
	{8'd233,8'd51} : s = 284;
	{8'd233,8'd52} : s = 285;
	{8'd233,8'd53} : s = 286;
	{8'd233,8'd54} : s = 287;
	{8'd233,8'd55} : s = 288;
	{8'd233,8'd56} : s = 289;
	{8'd233,8'd57} : s = 290;
	{8'd233,8'd58} : s = 291;
	{8'd233,8'd59} : s = 292;
	{8'd233,8'd60} : s = 293;
	{8'd233,8'd61} : s = 294;
	{8'd233,8'd62} : s = 295;
	{8'd233,8'd63} : s = 296;
	{8'd233,8'd64} : s = 297;
	{8'd233,8'd65} : s = 298;
	{8'd233,8'd66} : s = 299;
	{8'd233,8'd67} : s = 300;
	{8'd233,8'd68} : s = 301;
	{8'd233,8'd69} : s = 302;
	{8'd233,8'd70} : s = 303;
	{8'd233,8'd71} : s = 304;
	{8'd233,8'd72} : s = 305;
	{8'd233,8'd73} : s = 306;
	{8'd233,8'd74} : s = 307;
	{8'd233,8'd75} : s = 308;
	{8'd233,8'd76} : s = 309;
	{8'd233,8'd77} : s = 310;
	{8'd233,8'd78} : s = 311;
	{8'd233,8'd79} : s = 312;
	{8'd233,8'd80} : s = 313;
	{8'd233,8'd81} : s = 314;
	{8'd233,8'd82} : s = 315;
	{8'd233,8'd83} : s = 316;
	{8'd233,8'd84} : s = 317;
	{8'd233,8'd85} : s = 318;
	{8'd233,8'd86} : s = 319;
	{8'd233,8'd87} : s = 320;
	{8'd233,8'd88} : s = 321;
	{8'd233,8'd89} : s = 322;
	{8'd233,8'd90} : s = 323;
	{8'd233,8'd91} : s = 324;
	{8'd233,8'd92} : s = 325;
	{8'd233,8'd93} : s = 326;
	{8'd233,8'd94} : s = 327;
	{8'd233,8'd95} : s = 328;
	{8'd233,8'd96} : s = 329;
	{8'd233,8'd97} : s = 330;
	{8'd233,8'd98} : s = 331;
	{8'd233,8'd99} : s = 332;
	{8'd233,8'd100} : s = 333;
	{8'd233,8'd101} : s = 334;
	{8'd233,8'd102} : s = 335;
	{8'd233,8'd103} : s = 336;
	{8'd233,8'd104} : s = 337;
	{8'd233,8'd105} : s = 338;
	{8'd233,8'd106} : s = 339;
	{8'd233,8'd107} : s = 340;
	{8'd233,8'd108} : s = 341;
	{8'd233,8'd109} : s = 342;
	{8'd233,8'd110} : s = 343;
	{8'd233,8'd111} : s = 344;
	{8'd233,8'd112} : s = 345;
	{8'd233,8'd113} : s = 346;
	{8'd233,8'd114} : s = 347;
	{8'd233,8'd115} : s = 348;
	{8'd233,8'd116} : s = 349;
	{8'd233,8'd117} : s = 350;
	{8'd233,8'd118} : s = 351;
	{8'd233,8'd119} : s = 352;
	{8'd233,8'd120} : s = 353;
	{8'd233,8'd121} : s = 354;
	{8'd233,8'd122} : s = 355;
	{8'd233,8'd123} : s = 356;
	{8'd233,8'd124} : s = 357;
	{8'd233,8'd125} : s = 358;
	{8'd233,8'd126} : s = 359;
	{8'd233,8'd127} : s = 360;
	{8'd233,8'd128} : s = 361;
	{8'd233,8'd129} : s = 362;
	{8'd233,8'd130} : s = 363;
	{8'd233,8'd131} : s = 364;
	{8'd233,8'd132} : s = 365;
	{8'd233,8'd133} : s = 366;
	{8'd233,8'd134} : s = 367;
	{8'd233,8'd135} : s = 368;
	{8'd233,8'd136} : s = 369;
	{8'd233,8'd137} : s = 370;
	{8'd233,8'd138} : s = 371;
	{8'd233,8'd139} : s = 372;
	{8'd233,8'd140} : s = 373;
	{8'd233,8'd141} : s = 374;
	{8'd233,8'd142} : s = 375;
	{8'd233,8'd143} : s = 376;
	{8'd233,8'd144} : s = 377;
	{8'd233,8'd145} : s = 378;
	{8'd233,8'd146} : s = 379;
	{8'd233,8'd147} : s = 380;
	{8'd233,8'd148} : s = 381;
	{8'd233,8'd149} : s = 382;
	{8'd233,8'd150} : s = 383;
	{8'd233,8'd151} : s = 384;
	{8'd233,8'd152} : s = 385;
	{8'd233,8'd153} : s = 386;
	{8'd233,8'd154} : s = 387;
	{8'd233,8'd155} : s = 388;
	{8'd233,8'd156} : s = 389;
	{8'd233,8'd157} : s = 390;
	{8'd233,8'd158} : s = 391;
	{8'd233,8'd159} : s = 392;
	{8'd233,8'd160} : s = 393;
	{8'd233,8'd161} : s = 394;
	{8'd233,8'd162} : s = 395;
	{8'd233,8'd163} : s = 396;
	{8'd233,8'd164} : s = 397;
	{8'd233,8'd165} : s = 398;
	{8'd233,8'd166} : s = 399;
	{8'd233,8'd167} : s = 400;
	{8'd233,8'd168} : s = 401;
	{8'd233,8'd169} : s = 402;
	{8'd233,8'd170} : s = 403;
	{8'd233,8'd171} : s = 404;
	{8'd233,8'd172} : s = 405;
	{8'd233,8'd173} : s = 406;
	{8'd233,8'd174} : s = 407;
	{8'd233,8'd175} : s = 408;
	{8'd233,8'd176} : s = 409;
	{8'd233,8'd177} : s = 410;
	{8'd233,8'd178} : s = 411;
	{8'd233,8'd179} : s = 412;
	{8'd233,8'd180} : s = 413;
	{8'd233,8'd181} : s = 414;
	{8'd233,8'd182} : s = 415;
	{8'd233,8'd183} : s = 416;
	{8'd233,8'd184} : s = 417;
	{8'd233,8'd185} : s = 418;
	{8'd233,8'd186} : s = 419;
	{8'd233,8'd187} : s = 420;
	{8'd233,8'd188} : s = 421;
	{8'd233,8'd189} : s = 422;
	{8'd233,8'd190} : s = 423;
	{8'd233,8'd191} : s = 424;
	{8'd233,8'd192} : s = 425;
	{8'd233,8'd193} : s = 426;
	{8'd233,8'd194} : s = 427;
	{8'd233,8'd195} : s = 428;
	{8'd233,8'd196} : s = 429;
	{8'd233,8'd197} : s = 430;
	{8'd233,8'd198} : s = 431;
	{8'd233,8'd199} : s = 432;
	{8'd233,8'd200} : s = 433;
	{8'd233,8'd201} : s = 434;
	{8'd233,8'd202} : s = 435;
	{8'd233,8'd203} : s = 436;
	{8'd233,8'd204} : s = 437;
	{8'd233,8'd205} : s = 438;
	{8'd233,8'd206} : s = 439;
	{8'd233,8'd207} : s = 440;
	{8'd233,8'd208} : s = 441;
	{8'd233,8'd209} : s = 442;
	{8'd233,8'd210} : s = 443;
	{8'd233,8'd211} : s = 444;
	{8'd233,8'd212} : s = 445;
	{8'd233,8'd213} : s = 446;
	{8'd233,8'd214} : s = 447;
	{8'd233,8'd215} : s = 448;
	{8'd233,8'd216} : s = 449;
	{8'd233,8'd217} : s = 450;
	{8'd233,8'd218} : s = 451;
	{8'd233,8'd219} : s = 452;
	{8'd233,8'd220} : s = 453;
	{8'd233,8'd221} : s = 454;
	{8'd233,8'd222} : s = 455;
	{8'd233,8'd223} : s = 456;
	{8'd233,8'd224} : s = 457;
	{8'd233,8'd225} : s = 458;
	{8'd233,8'd226} : s = 459;
	{8'd233,8'd227} : s = 460;
	{8'd233,8'd228} : s = 461;
	{8'd233,8'd229} : s = 462;
	{8'd233,8'd230} : s = 463;
	{8'd233,8'd231} : s = 464;
	{8'd233,8'd232} : s = 465;
	{8'd233,8'd233} : s = 466;
	{8'd233,8'd234} : s = 467;
	{8'd233,8'd235} : s = 468;
	{8'd233,8'd236} : s = 469;
	{8'd233,8'd237} : s = 470;
	{8'd233,8'd238} : s = 471;
	{8'd233,8'd239} : s = 472;
	{8'd233,8'd240} : s = 473;
	{8'd233,8'd241} : s = 474;
	{8'd233,8'd242} : s = 475;
	{8'd233,8'd243} : s = 476;
	{8'd233,8'd244} : s = 477;
	{8'd233,8'd245} : s = 478;
	{8'd233,8'd246} : s = 479;
	{8'd233,8'd247} : s = 480;
	{8'd233,8'd248} : s = 481;
	{8'd233,8'd249} : s = 482;
	{8'd233,8'd250} : s = 483;
	{8'd233,8'd251} : s = 484;
	{8'd233,8'd252} : s = 485;
	{8'd233,8'd253} : s = 486;
	{8'd233,8'd254} : s = 487;
	{8'd233,8'd255} : s = 488;
	{8'd234,8'd0} : s = 234;
	{8'd234,8'd1} : s = 235;
	{8'd234,8'd2} : s = 236;
	{8'd234,8'd3} : s = 237;
	{8'd234,8'd4} : s = 238;
	{8'd234,8'd5} : s = 239;
	{8'd234,8'd6} : s = 240;
	{8'd234,8'd7} : s = 241;
	{8'd234,8'd8} : s = 242;
	{8'd234,8'd9} : s = 243;
	{8'd234,8'd10} : s = 244;
	{8'd234,8'd11} : s = 245;
	{8'd234,8'd12} : s = 246;
	{8'd234,8'd13} : s = 247;
	{8'd234,8'd14} : s = 248;
	{8'd234,8'd15} : s = 249;
	{8'd234,8'd16} : s = 250;
	{8'd234,8'd17} : s = 251;
	{8'd234,8'd18} : s = 252;
	{8'd234,8'd19} : s = 253;
	{8'd234,8'd20} : s = 254;
	{8'd234,8'd21} : s = 255;
	{8'd234,8'd22} : s = 256;
	{8'd234,8'd23} : s = 257;
	{8'd234,8'd24} : s = 258;
	{8'd234,8'd25} : s = 259;
	{8'd234,8'd26} : s = 260;
	{8'd234,8'd27} : s = 261;
	{8'd234,8'd28} : s = 262;
	{8'd234,8'd29} : s = 263;
	{8'd234,8'd30} : s = 264;
	{8'd234,8'd31} : s = 265;
	{8'd234,8'd32} : s = 266;
	{8'd234,8'd33} : s = 267;
	{8'd234,8'd34} : s = 268;
	{8'd234,8'd35} : s = 269;
	{8'd234,8'd36} : s = 270;
	{8'd234,8'd37} : s = 271;
	{8'd234,8'd38} : s = 272;
	{8'd234,8'd39} : s = 273;
	{8'd234,8'd40} : s = 274;
	{8'd234,8'd41} : s = 275;
	{8'd234,8'd42} : s = 276;
	{8'd234,8'd43} : s = 277;
	{8'd234,8'd44} : s = 278;
	{8'd234,8'd45} : s = 279;
	{8'd234,8'd46} : s = 280;
	{8'd234,8'd47} : s = 281;
	{8'd234,8'd48} : s = 282;
	{8'd234,8'd49} : s = 283;
	{8'd234,8'd50} : s = 284;
	{8'd234,8'd51} : s = 285;
	{8'd234,8'd52} : s = 286;
	{8'd234,8'd53} : s = 287;
	{8'd234,8'd54} : s = 288;
	{8'd234,8'd55} : s = 289;
	{8'd234,8'd56} : s = 290;
	{8'd234,8'd57} : s = 291;
	{8'd234,8'd58} : s = 292;
	{8'd234,8'd59} : s = 293;
	{8'd234,8'd60} : s = 294;
	{8'd234,8'd61} : s = 295;
	{8'd234,8'd62} : s = 296;
	{8'd234,8'd63} : s = 297;
	{8'd234,8'd64} : s = 298;
	{8'd234,8'd65} : s = 299;
	{8'd234,8'd66} : s = 300;
	{8'd234,8'd67} : s = 301;
	{8'd234,8'd68} : s = 302;
	{8'd234,8'd69} : s = 303;
	{8'd234,8'd70} : s = 304;
	{8'd234,8'd71} : s = 305;
	{8'd234,8'd72} : s = 306;
	{8'd234,8'd73} : s = 307;
	{8'd234,8'd74} : s = 308;
	{8'd234,8'd75} : s = 309;
	{8'd234,8'd76} : s = 310;
	{8'd234,8'd77} : s = 311;
	{8'd234,8'd78} : s = 312;
	{8'd234,8'd79} : s = 313;
	{8'd234,8'd80} : s = 314;
	{8'd234,8'd81} : s = 315;
	{8'd234,8'd82} : s = 316;
	{8'd234,8'd83} : s = 317;
	{8'd234,8'd84} : s = 318;
	{8'd234,8'd85} : s = 319;
	{8'd234,8'd86} : s = 320;
	{8'd234,8'd87} : s = 321;
	{8'd234,8'd88} : s = 322;
	{8'd234,8'd89} : s = 323;
	{8'd234,8'd90} : s = 324;
	{8'd234,8'd91} : s = 325;
	{8'd234,8'd92} : s = 326;
	{8'd234,8'd93} : s = 327;
	{8'd234,8'd94} : s = 328;
	{8'd234,8'd95} : s = 329;
	{8'd234,8'd96} : s = 330;
	{8'd234,8'd97} : s = 331;
	{8'd234,8'd98} : s = 332;
	{8'd234,8'd99} : s = 333;
	{8'd234,8'd100} : s = 334;
	{8'd234,8'd101} : s = 335;
	{8'd234,8'd102} : s = 336;
	{8'd234,8'd103} : s = 337;
	{8'd234,8'd104} : s = 338;
	{8'd234,8'd105} : s = 339;
	{8'd234,8'd106} : s = 340;
	{8'd234,8'd107} : s = 341;
	{8'd234,8'd108} : s = 342;
	{8'd234,8'd109} : s = 343;
	{8'd234,8'd110} : s = 344;
	{8'd234,8'd111} : s = 345;
	{8'd234,8'd112} : s = 346;
	{8'd234,8'd113} : s = 347;
	{8'd234,8'd114} : s = 348;
	{8'd234,8'd115} : s = 349;
	{8'd234,8'd116} : s = 350;
	{8'd234,8'd117} : s = 351;
	{8'd234,8'd118} : s = 352;
	{8'd234,8'd119} : s = 353;
	{8'd234,8'd120} : s = 354;
	{8'd234,8'd121} : s = 355;
	{8'd234,8'd122} : s = 356;
	{8'd234,8'd123} : s = 357;
	{8'd234,8'd124} : s = 358;
	{8'd234,8'd125} : s = 359;
	{8'd234,8'd126} : s = 360;
	{8'd234,8'd127} : s = 361;
	{8'd234,8'd128} : s = 362;
	{8'd234,8'd129} : s = 363;
	{8'd234,8'd130} : s = 364;
	{8'd234,8'd131} : s = 365;
	{8'd234,8'd132} : s = 366;
	{8'd234,8'd133} : s = 367;
	{8'd234,8'd134} : s = 368;
	{8'd234,8'd135} : s = 369;
	{8'd234,8'd136} : s = 370;
	{8'd234,8'd137} : s = 371;
	{8'd234,8'd138} : s = 372;
	{8'd234,8'd139} : s = 373;
	{8'd234,8'd140} : s = 374;
	{8'd234,8'd141} : s = 375;
	{8'd234,8'd142} : s = 376;
	{8'd234,8'd143} : s = 377;
	{8'd234,8'd144} : s = 378;
	{8'd234,8'd145} : s = 379;
	{8'd234,8'd146} : s = 380;
	{8'd234,8'd147} : s = 381;
	{8'd234,8'd148} : s = 382;
	{8'd234,8'd149} : s = 383;
	{8'd234,8'd150} : s = 384;
	{8'd234,8'd151} : s = 385;
	{8'd234,8'd152} : s = 386;
	{8'd234,8'd153} : s = 387;
	{8'd234,8'd154} : s = 388;
	{8'd234,8'd155} : s = 389;
	{8'd234,8'd156} : s = 390;
	{8'd234,8'd157} : s = 391;
	{8'd234,8'd158} : s = 392;
	{8'd234,8'd159} : s = 393;
	{8'd234,8'd160} : s = 394;
	{8'd234,8'd161} : s = 395;
	{8'd234,8'd162} : s = 396;
	{8'd234,8'd163} : s = 397;
	{8'd234,8'd164} : s = 398;
	{8'd234,8'd165} : s = 399;
	{8'd234,8'd166} : s = 400;
	{8'd234,8'd167} : s = 401;
	{8'd234,8'd168} : s = 402;
	{8'd234,8'd169} : s = 403;
	{8'd234,8'd170} : s = 404;
	{8'd234,8'd171} : s = 405;
	{8'd234,8'd172} : s = 406;
	{8'd234,8'd173} : s = 407;
	{8'd234,8'd174} : s = 408;
	{8'd234,8'd175} : s = 409;
	{8'd234,8'd176} : s = 410;
	{8'd234,8'd177} : s = 411;
	{8'd234,8'd178} : s = 412;
	{8'd234,8'd179} : s = 413;
	{8'd234,8'd180} : s = 414;
	{8'd234,8'd181} : s = 415;
	{8'd234,8'd182} : s = 416;
	{8'd234,8'd183} : s = 417;
	{8'd234,8'd184} : s = 418;
	{8'd234,8'd185} : s = 419;
	{8'd234,8'd186} : s = 420;
	{8'd234,8'd187} : s = 421;
	{8'd234,8'd188} : s = 422;
	{8'd234,8'd189} : s = 423;
	{8'd234,8'd190} : s = 424;
	{8'd234,8'd191} : s = 425;
	{8'd234,8'd192} : s = 426;
	{8'd234,8'd193} : s = 427;
	{8'd234,8'd194} : s = 428;
	{8'd234,8'd195} : s = 429;
	{8'd234,8'd196} : s = 430;
	{8'd234,8'd197} : s = 431;
	{8'd234,8'd198} : s = 432;
	{8'd234,8'd199} : s = 433;
	{8'd234,8'd200} : s = 434;
	{8'd234,8'd201} : s = 435;
	{8'd234,8'd202} : s = 436;
	{8'd234,8'd203} : s = 437;
	{8'd234,8'd204} : s = 438;
	{8'd234,8'd205} : s = 439;
	{8'd234,8'd206} : s = 440;
	{8'd234,8'd207} : s = 441;
	{8'd234,8'd208} : s = 442;
	{8'd234,8'd209} : s = 443;
	{8'd234,8'd210} : s = 444;
	{8'd234,8'd211} : s = 445;
	{8'd234,8'd212} : s = 446;
	{8'd234,8'd213} : s = 447;
	{8'd234,8'd214} : s = 448;
	{8'd234,8'd215} : s = 449;
	{8'd234,8'd216} : s = 450;
	{8'd234,8'd217} : s = 451;
	{8'd234,8'd218} : s = 452;
	{8'd234,8'd219} : s = 453;
	{8'd234,8'd220} : s = 454;
	{8'd234,8'd221} : s = 455;
	{8'd234,8'd222} : s = 456;
	{8'd234,8'd223} : s = 457;
	{8'd234,8'd224} : s = 458;
	{8'd234,8'd225} : s = 459;
	{8'd234,8'd226} : s = 460;
	{8'd234,8'd227} : s = 461;
	{8'd234,8'd228} : s = 462;
	{8'd234,8'd229} : s = 463;
	{8'd234,8'd230} : s = 464;
	{8'd234,8'd231} : s = 465;
	{8'd234,8'd232} : s = 466;
	{8'd234,8'd233} : s = 467;
	{8'd234,8'd234} : s = 468;
	{8'd234,8'd235} : s = 469;
	{8'd234,8'd236} : s = 470;
	{8'd234,8'd237} : s = 471;
	{8'd234,8'd238} : s = 472;
	{8'd234,8'd239} : s = 473;
	{8'd234,8'd240} : s = 474;
	{8'd234,8'd241} : s = 475;
	{8'd234,8'd242} : s = 476;
	{8'd234,8'd243} : s = 477;
	{8'd234,8'd244} : s = 478;
	{8'd234,8'd245} : s = 479;
	{8'd234,8'd246} : s = 480;
	{8'd234,8'd247} : s = 481;
	{8'd234,8'd248} : s = 482;
	{8'd234,8'd249} : s = 483;
	{8'd234,8'd250} : s = 484;
	{8'd234,8'd251} : s = 485;
	{8'd234,8'd252} : s = 486;
	{8'd234,8'd253} : s = 487;
	{8'd234,8'd254} : s = 488;
	{8'd234,8'd255} : s = 489;
	{8'd235,8'd0} : s = 235;
	{8'd235,8'd1} : s = 236;
	{8'd235,8'd2} : s = 237;
	{8'd235,8'd3} : s = 238;
	{8'd235,8'd4} : s = 239;
	{8'd235,8'd5} : s = 240;
	{8'd235,8'd6} : s = 241;
	{8'd235,8'd7} : s = 242;
	{8'd235,8'd8} : s = 243;
	{8'd235,8'd9} : s = 244;
	{8'd235,8'd10} : s = 245;
	{8'd235,8'd11} : s = 246;
	{8'd235,8'd12} : s = 247;
	{8'd235,8'd13} : s = 248;
	{8'd235,8'd14} : s = 249;
	{8'd235,8'd15} : s = 250;
	{8'd235,8'd16} : s = 251;
	{8'd235,8'd17} : s = 252;
	{8'd235,8'd18} : s = 253;
	{8'd235,8'd19} : s = 254;
	{8'd235,8'd20} : s = 255;
	{8'd235,8'd21} : s = 256;
	{8'd235,8'd22} : s = 257;
	{8'd235,8'd23} : s = 258;
	{8'd235,8'd24} : s = 259;
	{8'd235,8'd25} : s = 260;
	{8'd235,8'd26} : s = 261;
	{8'd235,8'd27} : s = 262;
	{8'd235,8'd28} : s = 263;
	{8'd235,8'd29} : s = 264;
	{8'd235,8'd30} : s = 265;
	{8'd235,8'd31} : s = 266;
	{8'd235,8'd32} : s = 267;
	{8'd235,8'd33} : s = 268;
	{8'd235,8'd34} : s = 269;
	{8'd235,8'd35} : s = 270;
	{8'd235,8'd36} : s = 271;
	{8'd235,8'd37} : s = 272;
	{8'd235,8'd38} : s = 273;
	{8'd235,8'd39} : s = 274;
	{8'd235,8'd40} : s = 275;
	{8'd235,8'd41} : s = 276;
	{8'd235,8'd42} : s = 277;
	{8'd235,8'd43} : s = 278;
	{8'd235,8'd44} : s = 279;
	{8'd235,8'd45} : s = 280;
	{8'd235,8'd46} : s = 281;
	{8'd235,8'd47} : s = 282;
	{8'd235,8'd48} : s = 283;
	{8'd235,8'd49} : s = 284;
	{8'd235,8'd50} : s = 285;
	{8'd235,8'd51} : s = 286;
	{8'd235,8'd52} : s = 287;
	{8'd235,8'd53} : s = 288;
	{8'd235,8'd54} : s = 289;
	{8'd235,8'd55} : s = 290;
	{8'd235,8'd56} : s = 291;
	{8'd235,8'd57} : s = 292;
	{8'd235,8'd58} : s = 293;
	{8'd235,8'd59} : s = 294;
	{8'd235,8'd60} : s = 295;
	{8'd235,8'd61} : s = 296;
	{8'd235,8'd62} : s = 297;
	{8'd235,8'd63} : s = 298;
	{8'd235,8'd64} : s = 299;
	{8'd235,8'd65} : s = 300;
	{8'd235,8'd66} : s = 301;
	{8'd235,8'd67} : s = 302;
	{8'd235,8'd68} : s = 303;
	{8'd235,8'd69} : s = 304;
	{8'd235,8'd70} : s = 305;
	{8'd235,8'd71} : s = 306;
	{8'd235,8'd72} : s = 307;
	{8'd235,8'd73} : s = 308;
	{8'd235,8'd74} : s = 309;
	{8'd235,8'd75} : s = 310;
	{8'd235,8'd76} : s = 311;
	{8'd235,8'd77} : s = 312;
	{8'd235,8'd78} : s = 313;
	{8'd235,8'd79} : s = 314;
	{8'd235,8'd80} : s = 315;
	{8'd235,8'd81} : s = 316;
	{8'd235,8'd82} : s = 317;
	{8'd235,8'd83} : s = 318;
	{8'd235,8'd84} : s = 319;
	{8'd235,8'd85} : s = 320;
	{8'd235,8'd86} : s = 321;
	{8'd235,8'd87} : s = 322;
	{8'd235,8'd88} : s = 323;
	{8'd235,8'd89} : s = 324;
	{8'd235,8'd90} : s = 325;
	{8'd235,8'd91} : s = 326;
	{8'd235,8'd92} : s = 327;
	{8'd235,8'd93} : s = 328;
	{8'd235,8'd94} : s = 329;
	{8'd235,8'd95} : s = 330;
	{8'd235,8'd96} : s = 331;
	{8'd235,8'd97} : s = 332;
	{8'd235,8'd98} : s = 333;
	{8'd235,8'd99} : s = 334;
	{8'd235,8'd100} : s = 335;
	{8'd235,8'd101} : s = 336;
	{8'd235,8'd102} : s = 337;
	{8'd235,8'd103} : s = 338;
	{8'd235,8'd104} : s = 339;
	{8'd235,8'd105} : s = 340;
	{8'd235,8'd106} : s = 341;
	{8'd235,8'd107} : s = 342;
	{8'd235,8'd108} : s = 343;
	{8'd235,8'd109} : s = 344;
	{8'd235,8'd110} : s = 345;
	{8'd235,8'd111} : s = 346;
	{8'd235,8'd112} : s = 347;
	{8'd235,8'd113} : s = 348;
	{8'd235,8'd114} : s = 349;
	{8'd235,8'd115} : s = 350;
	{8'd235,8'd116} : s = 351;
	{8'd235,8'd117} : s = 352;
	{8'd235,8'd118} : s = 353;
	{8'd235,8'd119} : s = 354;
	{8'd235,8'd120} : s = 355;
	{8'd235,8'd121} : s = 356;
	{8'd235,8'd122} : s = 357;
	{8'd235,8'd123} : s = 358;
	{8'd235,8'd124} : s = 359;
	{8'd235,8'd125} : s = 360;
	{8'd235,8'd126} : s = 361;
	{8'd235,8'd127} : s = 362;
	{8'd235,8'd128} : s = 363;
	{8'd235,8'd129} : s = 364;
	{8'd235,8'd130} : s = 365;
	{8'd235,8'd131} : s = 366;
	{8'd235,8'd132} : s = 367;
	{8'd235,8'd133} : s = 368;
	{8'd235,8'd134} : s = 369;
	{8'd235,8'd135} : s = 370;
	{8'd235,8'd136} : s = 371;
	{8'd235,8'd137} : s = 372;
	{8'd235,8'd138} : s = 373;
	{8'd235,8'd139} : s = 374;
	{8'd235,8'd140} : s = 375;
	{8'd235,8'd141} : s = 376;
	{8'd235,8'd142} : s = 377;
	{8'd235,8'd143} : s = 378;
	{8'd235,8'd144} : s = 379;
	{8'd235,8'd145} : s = 380;
	{8'd235,8'd146} : s = 381;
	{8'd235,8'd147} : s = 382;
	{8'd235,8'd148} : s = 383;
	{8'd235,8'd149} : s = 384;
	{8'd235,8'd150} : s = 385;
	{8'd235,8'd151} : s = 386;
	{8'd235,8'd152} : s = 387;
	{8'd235,8'd153} : s = 388;
	{8'd235,8'd154} : s = 389;
	{8'd235,8'd155} : s = 390;
	{8'd235,8'd156} : s = 391;
	{8'd235,8'd157} : s = 392;
	{8'd235,8'd158} : s = 393;
	{8'd235,8'd159} : s = 394;
	{8'd235,8'd160} : s = 395;
	{8'd235,8'd161} : s = 396;
	{8'd235,8'd162} : s = 397;
	{8'd235,8'd163} : s = 398;
	{8'd235,8'd164} : s = 399;
	{8'd235,8'd165} : s = 400;
	{8'd235,8'd166} : s = 401;
	{8'd235,8'd167} : s = 402;
	{8'd235,8'd168} : s = 403;
	{8'd235,8'd169} : s = 404;
	{8'd235,8'd170} : s = 405;
	{8'd235,8'd171} : s = 406;
	{8'd235,8'd172} : s = 407;
	{8'd235,8'd173} : s = 408;
	{8'd235,8'd174} : s = 409;
	{8'd235,8'd175} : s = 410;
	{8'd235,8'd176} : s = 411;
	{8'd235,8'd177} : s = 412;
	{8'd235,8'd178} : s = 413;
	{8'd235,8'd179} : s = 414;
	{8'd235,8'd180} : s = 415;
	{8'd235,8'd181} : s = 416;
	{8'd235,8'd182} : s = 417;
	{8'd235,8'd183} : s = 418;
	{8'd235,8'd184} : s = 419;
	{8'd235,8'd185} : s = 420;
	{8'd235,8'd186} : s = 421;
	{8'd235,8'd187} : s = 422;
	{8'd235,8'd188} : s = 423;
	{8'd235,8'd189} : s = 424;
	{8'd235,8'd190} : s = 425;
	{8'd235,8'd191} : s = 426;
	{8'd235,8'd192} : s = 427;
	{8'd235,8'd193} : s = 428;
	{8'd235,8'd194} : s = 429;
	{8'd235,8'd195} : s = 430;
	{8'd235,8'd196} : s = 431;
	{8'd235,8'd197} : s = 432;
	{8'd235,8'd198} : s = 433;
	{8'd235,8'd199} : s = 434;
	{8'd235,8'd200} : s = 435;
	{8'd235,8'd201} : s = 436;
	{8'd235,8'd202} : s = 437;
	{8'd235,8'd203} : s = 438;
	{8'd235,8'd204} : s = 439;
	{8'd235,8'd205} : s = 440;
	{8'd235,8'd206} : s = 441;
	{8'd235,8'd207} : s = 442;
	{8'd235,8'd208} : s = 443;
	{8'd235,8'd209} : s = 444;
	{8'd235,8'd210} : s = 445;
	{8'd235,8'd211} : s = 446;
	{8'd235,8'd212} : s = 447;
	{8'd235,8'd213} : s = 448;
	{8'd235,8'd214} : s = 449;
	{8'd235,8'd215} : s = 450;
	{8'd235,8'd216} : s = 451;
	{8'd235,8'd217} : s = 452;
	{8'd235,8'd218} : s = 453;
	{8'd235,8'd219} : s = 454;
	{8'd235,8'd220} : s = 455;
	{8'd235,8'd221} : s = 456;
	{8'd235,8'd222} : s = 457;
	{8'd235,8'd223} : s = 458;
	{8'd235,8'd224} : s = 459;
	{8'd235,8'd225} : s = 460;
	{8'd235,8'd226} : s = 461;
	{8'd235,8'd227} : s = 462;
	{8'd235,8'd228} : s = 463;
	{8'd235,8'd229} : s = 464;
	{8'd235,8'd230} : s = 465;
	{8'd235,8'd231} : s = 466;
	{8'd235,8'd232} : s = 467;
	{8'd235,8'd233} : s = 468;
	{8'd235,8'd234} : s = 469;
	{8'd235,8'd235} : s = 470;
	{8'd235,8'd236} : s = 471;
	{8'd235,8'd237} : s = 472;
	{8'd235,8'd238} : s = 473;
	{8'd235,8'd239} : s = 474;
	{8'd235,8'd240} : s = 475;
	{8'd235,8'd241} : s = 476;
	{8'd235,8'd242} : s = 477;
	{8'd235,8'd243} : s = 478;
	{8'd235,8'd244} : s = 479;
	{8'd235,8'd245} : s = 480;
	{8'd235,8'd246} : s = 481;
	{8'd235,8'd247} : s = 482;
	{8'd235,8'd248} : s = 483;
	{8'd235,8'd249} : s = 484;
	{8'd235,8'd250} : s = 485;
	{8'd235,8'd251} : s = 486;
	{8'd235,8'd252} : s = 487;
	{8'd235,8'd253} : s = 488;
	{8'd235,8'd254} : s = 489;
	{8'd235,8'd255} : s = 490;
	{8'd236,8'd0} : s = 236;
	{8'd236,8'd1} : s = 237;
	{8'd236,8'd2} : s = 238;
	{8'd236,8'd3} : s = 239;
	{8'd236,8'd4} : s = 240;
	{8'd236,8'd5} : s = 241;
	{8'd236,8'd6} : s = 242;
	{8'd236,8'd7} : s = 243;
	{8'd236,8'd8} : s = 244;
	{8'd236,8'd9} : s = 245;
	{8'd236,8'd10} : s = 246;
	{8'd236,8'd11} : s = 247;
	{8'd236,8'd12} : s = 248;
	{8'd236,8'd13} : s = 249;
	{8'd236,8'd14} : s = 250;
	{8'd236,8'd15} : s = 251;
	{8'd236,8'd16} : s = 252;
	{8'd236,8'd17} : s = 253;
	{8'd236,8'd18} : s = 254;
	{8'd236,8'd19} : s = 255;
	{8'd236,8'd20} : s = 256;
	{8'd236,8'd21} : s = 257;
	{8'd236,8'd22} : s = 258;
	{8'd236,8'd23} : s = 259;
	{8'd236,8'd24} : s = 260;
	{8'd236,8'd25} : s = 261;
	{8'd236,8'd26} : s = 262;
	{8'd236,8'd27} : s = 263;
	{8'd236,8'd28} : s = 264;
	{8'd236,8'd29} : s = 265;
	{8'd236,8'd30} : s = 266;
	{8'd236,8'd31} : s = 267;
	{8'd236,8'd32} : s = 268;
	{8'd236,8'd33} : s = 269;
	{8'd236,8'd34} : s = 270;
	{8'd236,8'd35} : s = 271;
	{8'd236,8'd36} : s = 272;
	{8'd236,8'd37} : s = 273;
	{8'd236,8'd38} : s = 274;
	{8'd236,8'd39} : s = 275;
	{8'd236,8'd40} : s = 276;
	{8'd236,8'd41} : s = 277;
	{8'd236,8'd42} : s = 278;
	{8'd236,8'd43} : s = 279;
	{8'd236,8'd44} : s = 280;
	{8'd236,8'd45} : s = 281;
	{8'd236,8'd46} : s = 282;
	{8'd236,8'd47} : s = 283;
	{8'd236,8'd48} : s = 284;
	{8'd236,8'd49} : s = 285;
	{8'd236,8'd50} : s = 286;
	{8'd236,8'd51} : s = 287;
	{8'd236,8'd52} : s = 288;
	{8'd236,8'd53} : s = 289;
	{8'd236,8'd54} : s = 290;
	{8'd236,8'd55} : s = 291;
	{8'd236,8'd56} : s = 292;
	{8'd236,8'd57} : s = 293;
	{8'd236,8'd58} : s = 294;
	{8'd236,8'd59} : s = 295;
	{8'd236,8'd60} : s = 296;
	{8'd236,8'd61} : s = 297;
	{8'd236,8'd62} : s = 298;
	{8'd236,8'd63} : s = 299;
	{8'd236,8'd64} : s = 300;
	{8'd236,8'd65} : s = 301;
	{8'd236,8'd66} : s = 302;
	{8'd236,8'd67} : s = 303;
	{8'd236,8'd68} : s = 304;
	{8'd236,8'd69} : s = 305;
	{8'd236,8'd70} : s = 306;
	{8'd236,8'd71} : s = 307;
	{8'd236,8'd72} : s = 308;
	{8'd236,8'd73} : s = 309;
	{8'd236,8'd74} : s = 310;
	{8'd236,8'd75} : s = 311;
	{8'd236,8'd76} : s = 312;
	{8'd236,8'd77} : s = 313;
	{8'd236,8'd78} : s = 314;
	{8'd236,8'd79} : s = 315;
	{8'd236,8'd80} : s = 316;
	{8'd236,8'd81} : s = 317;
	{8'd236,8'd82} : s = 318;
	{8'd236,8'd83} : s = 319;
	{8'd236,8'd84} : s = 320;
	{8'd236,8'd85} : s = 321;
	{8'd236,8'd86} : s = 322;
	{8'd236,8'd87} : s = 323;
	{8'd236,8'd88} : s = 324;
	{8'd236,8'd89} : s = 325;
	{8'd236,8'd90} : s = 326;
	{8'd236,8'd91} : s = 327;
	{8'd236,8'd92} : s = 328;
	{8'd236,8'd93} : s = 329;
	{8'd236,8'd94} : s = 330;
	{8'd236,8'd95} : s = 331;
	{8'd236,8'd96} : s = 332;
	{8'd236,8'd97} : s = 333;
	{8'd236,8'd98} : s = 334;
	{8'd236,8'd99} : s = 335;
	{8'd236,8'd100} : s = 336;
	{8'd236,8'd101} : s = 337;
	{8'd236,8'd102} : s = 338;
	{8'd236,8'd103} : s = 339;
	{8'd236,8'd104} : s = 340;
	{8'd236,8'd105} : s = 341;
	{8'd236,8'd106} : s = 342;
	{8'd236,8'd107} : s = 343;
	{8'd236,8'd108} : s = 344;
	{8'd236,8'd109} : s = 345;
	{8'd236,8'd110} : s = 346;
	{8'd236,8'd111} : s = 347;
	{8'd236,8'd112} : s = 348;
	{8'd236,8'd113} : s = 349;
	{8'd236,8'd114} : s = 350;
	{8'd236,8'd115} : s = 351;
	{8'd236,8'd116} : s = 352;
	{8'd236,8'd117} : s = 353;
	{8'd236,8'd118} : s = 354;
	{8'd236,8'd119} : s = 355;
	{8'd236,8'd120} : s = 356;
	{8'd236,8'd121} : s = 357;
	{8'd236,8'd122} : s = 358;
	{8'd236,8'd123} : s = 359;
	{8'd236,8'd124} : s = 360;
	{8'd236,8'd125} : s = 361;
	{8'd236,8'd126} : s = 362;
	{8'd236,8'd127} : s = 363;
	{8'd236,8'd128} : s = 364;
	{8'd236,8'd129} : s = 365;
	{8'd236,8'd130} : s = 366;
	{8'd236,8'd131} : s = 367;
	{8'd236,8'd132} : s = 368;
	{8'd236,8'd133} : s = 369;
	{8'd236,8'd134} : s = 370;
	{8'd236,8'd135} : s = 371;
	{8'd236,8'd136} : s = 372;
	{8'd236,8'd137} : s = 373;
	{8'd236,8'd138} : s = 374;
	{8'd236,8'd139} : s = 375;
	{8'd236,8'd140} : s = 376;
	{8'd236,8'd141} : s = 377;
	{8'd236,8'd142} : s = 378;
	{8'd236,8'd143} : s = 379;
	{8'd236,8'd144} : s = 380;
	{8'd236,8'd145} : s = 381;
	{8'd236,8'd146} : s = 382;
	{8'd236,8'd147} : s = 383;
	{8'd236,8'd148} : s = 384;
	{8'd236,8'd149} : s = 385;
	{8'd236,8'd150} : s = 386;
	{8'd236,8'd151} : s = 387;
	{8'd236,8'd152} : s = 388;
	{8'd236,8'd153} : s = 389;
	{8'd236,8'd154} : s = 390;
	{8'd236,8'd155} : s = 391;
	{8'd236,8'd156} : s = 392;
	{8'd236,8'd157} : s = 393;
	{8'd236,8'd158} : s = 394;
	{8'd236,8'd159} : s = 395;
	{8'd236,8'd160} : s = 396;
	{8'd236,8'd161} : s = 397;
	{8'd236,8'd162} : s = 398;
	{8'd236,8'd163} : s = 399;
	{8'd236,8'd164} : s = 400;
	{8'd236,8'd165} : s = 401;
	{8'd236,8'd166} : s = 402;
	{8'd236,8'd167} : s = 403;
	{8'd236,8'd168} : s = 404;
	{8'd236,8'd169} : s = 405;
	{8'd236,8'd170} : s = 406;
	{8'd236,8'd171} : s = 407;
	{8'd236,8'd172} : s = 408;
	{8'd236,8'd173} : s = 409;
	{8'd236,8'd174} : s = 410;
	{8'd236,8'd175} : s = 411;
	{8'd236,8'd176} : s = 412;
	{8'd236,8'd177} : s = 413;
	{8'd236,8'd178} : s = 414;
	{8'd236,8'd179} : s = 415;
	{8'd236,8'd180} : s = 416;
	{8'd236,8'd181} : s = 417;
	{8'd236,8'd182} : s = 418;
	{8'd236,8'd183} : s = 419;
	{8'd236,8'd184} : s = 420;
	{8'd236,8'd185} : s = 421;
	{8'd236,8'd186} : s = 422;
	{8'd236,8'd187} : s = 423;
	{8'd236,8'd188} : s = 424;
	{8'd236,8'd189} : s = 425;
	{8'd236,8'd190} : s = 426;
	{8'd236,8'd191} : s = 427;
	{8'd236,8'd192} : s = 428;
	{8'd236,8'd193} : s = 429;
	{8'd236,8'd194} : s = 430;
	{8'd236,8'd195} : s = 431;
	{8'd236,8'd196} : s = 432;
	{8'd236,8'd197} : s = 433;
	{8'd236,8'd198} : s = 434;
	{8'd236,8'd199} : s = 435;
	{8'd236,8'd200} : s = 436;
	{8'd236,8'd201} : s = 437;
	{8'd236,8'd202} : s = 438;
	{8'd236,8'd203} : s = 439;
	{8'd236,8'd204} : s = 440;
	{8'd236,8'd205} : s = 441;
	{8'd236,8'd206} : s = 442;
	{8'd236,8'd207} : s = 443;
	{8'd236,8'd208} : s = 444;
	{8'd236,8'd209} : s = 445;
	{8'd236,8'd210} : s = 446;
	{8'd236,8'd211} : s = 447;
	{8'd236,8'd212} : s = 448;
	{8'd236,8'd213} : s = 449;
	{8'd236,8'd214} : s = 450;
	{8'd236,8'd215} : s = 451;
	{8'd236,8'd216} : s = 452;
	{8'd236,8'd217} : s = 453;
	{8'd236,8'd218} : s = 454;
	{8'd236,8'd219} : s = 455;
	{8'd236,8'd220} : s = 456;
	{8'd236,8'd221} : s = 457;
	{8'd236,8'd222} : s = 458;
	{8'd236,8'd223} : s = 459;
	{8'd236,8'd224} : s = 460;
	{8'd236,8'd225} : s = 461;
	{8'd236,8'd226} : s = 462;
	{8'd236,8'd227} : s = 463;
	{8'd236,8'd228} : s = 464;
	{8'd236,8'd229} : s = 465;
	{8'd236,8'd230} : s = 466;
	{8'd236,8'd231} : s = 467;
	{8'd236,8'd232} : s = 468;
	{8'd236,8'd233} : s = 469;
	{8'd236,8'd234} : s = 470;
	{8'd236,8'd235} : s = 471;
	{8'd236,8'd236} : s = 472;
	{8'd236,8'd237} : s = 473;
	{8'd236,8'd238} : s = 474;
	{8'd236,8'd239} : s = 475;
	{8'd236,8'd240} : s = 476;
	{8'd236,8'd241} : s = 477;
	{8'd236,8'd242} : s = 478;
	{8'd236,8'd243} : s = 479;
	{8'd236,8'd244} : s = 480;
	{8'd236,8'd245} : s = 481;
	{8'd236,8'd246} : s = 482;
	{8'd236,8'd247} : s = 483;
	{8'd236,8'd248} : s = 484;
	{8'd236,8'd249} : s = 485;
	{8'd236,8'd250} : s = 486;
	{8'd236,8'd251} : s = 487;
	{8'd236,8'd252} : s = 488;
	{8'd236,8'd253} : s = 489;
	{8'd236,8'd254} : s = 490;
	{8'd236,8'd255} : s = 491;
	{8'd237,8'd0} : s = 237;
	{8'd237,8'd1} : s = 238;
	{8'd237,8'd2} : s = 239;
	{8'd237,8'd3} : s = 240;
	{8'd237,8'd4} : s = 241;
	{8'd237,8'd5} : s = 242;
	{8'd237,8'd6} : s = 243;
	{8'd237,8'd7} : s = 244;
	{8'd237,8'd8} : s = 245;
	{8'd237,8'd9} : s = 246;
	{8'd237,8'd10} : s = 247;
	{8'd237,8'd11} : s = 248;
	{8'd237,8'd12} : s = 249;
	{8'd237,8'd13} : s = 250;
	{8'd237,8'd14} : s = 251;
	{8'd237,8'd15} : s = 252;
	{8'd237,8'd16} : s = 253;
	{8'd237,8'd17} : s = 254;
	{8'd237,8'd18} : s = 255;
	{8'd237,8'd19} : s = 256;
	{8'd237,8'd20} : s = 257;
	{8'd237,8'd21} : s = 258;
	{8'd237,8'd22} : s = 259;
	{8'd237,8'd23} : s = 260;
	{8'd237,8'd24} : s = 261;
	{8'd237,8'd25} : s = 262;
	{8'd237,8'd26} : s = 263;
	{8'd237,8'd27} : s = 264;
	{8'd237,8'd28} : s = 265;
	{8'd237,8'd29} : s = 266;
	{8'd237,8'd30} : s = 267;
	{8'd237,8'd31} : s = 268;
	{8'd237,8'd32} : s = 269;
	{8'd237,8'd33} : s = 270;
	{8'd237,8'd34} : s = 271;
	{8'd237,8'd35} : s = 272;
	{8'd237,8'd36} : s = 273;
	{8'd237,8'd37} : s = 274;
	{8'd237,8'd38} : s = 275;
	{8'd237,8'd39} : s = 276;
	{8'd237,8'd40} : s = 277;
	{8'd237,8'd41} : s = 278;
	{8'd237,8'd42} : s = 279;
	{8'd237,8'd43} : s = 280;
	{8'd237,8'd44} : s = 281;
	{8'd237,8'd45} : s = 282;
	{8'd237,8'd46} : s = 283;
	{8'd237,8'd47} : s = 284;
	{8'd237,8'd48} : s = 285;
	{8'd237,8'd49} : s = 286;
	{8'd237,8'd50} : s = 287;
	{8'd237,8'd51} : s = 288;
	{8'd237,8'd52} : s = 289;
	{8'd237,8'd53} : s = 290;
	{8'd237,8'd54} : s = 291;
	{8'd237,8'd55} : s = 292;
	{8'd237,8'd56} : s = 293;
	{8'd237,8'd57} : s = 294;
	{8'd237,8'd58} : s = 295;
	{8'd237,8'd59} : s = 296;
	{8'd237,8'd60} : s = 297;
	{8'd237,8'd61} : s = 298;
	{8'd237,8'd62} : s = 299;
	{8'd237,8'd63} : s = 300;
	{8'd237,8'd64} : s = 301;
	{8'd237,8'd65} : s = 302;
	{8'd237,8'd66} : s = 303;
	{8'd237,8'd67} : s = 304;
	{8'd237,8'd68} : s = 305;
	{8'd237,8'd69} : s = 306;
	{8'd237,8'd70} : s = 307;
	{8'd237,8'd71} : s = 308;
	{8'd237,8'd72} : s = 309;
	{8'd237,8'd73} : s = 310;
	{8'd237,8'd74} : s = 311;
	{8'd237,8'd75} : s = 312;
	{8'd237,8'd76} : s = 313;
	{8'd237,8'd77} : s = 314;
	{8'd237,8'd78} : s = 315;
	{8'd237,8'd79} : s = 316;
	{8'd237,8'd80} : s = 317;
	{8'd237,8'd81} : s = 318;
	{8'd237,8'd82} : s = 319;
	{8'd237,8'd83} : s = 320;
	{8'd237,8'd84} : s = 321;
	{8'd237,8'd85} : s = 322;
	{8'd237,8'd86} : s = 323;
	{8'd237,8'd87} : s = 324;
	{8'd237,8'd88} : s = 325;
	{8'd237,8'd89} : s = 326;
	{8'd237,8'd90} : s = 327;
	{8'd237,8'd91} : s = 328;
	{8'd237,8'd92} : s = 329;
	{8'd237,8'd93} : s = 330;
	{8'd237,8'd94} : s = 331;
	{8'd237,8'd95} : s = 332;
	{8'd237,8'd96} : s = 333;
	{8'd237,8'd97} : s = 334;
	{8'd237,8'd98} : s = 335;
	{8'd237,8'd99} : s = 336;
	{8'd237,8'd100} : s = 337;
	{8'd237,8'd101} : s = 338;
	{8'd237,8'd102} : s = 339;
	{8'd237,8'd103} : s = 340;
	{8'd237,8'd104} : s = 341;
	{8'd237,8'd105} : s = 342;
	{8'd237,8'd106} : s = 343;
	{8'd237,8'd107} : s = 344;
	{8'd237,8'd108} : s = 345;
	{8'd237,8'd109} : s = 346;
	{8'd237,8'd110} : s = 347;
	{8'd237,8'd111} : s = 348;
	{8'd237,8'd112} : s = 349;
	{8'd237,8'd113} : s = 350;
	{8'd237,8'd114} : s = 351;
	{8'd237,8'd115} : s = 352;
	{8'd237,8'd116} : s = 353;
	{8'd237,8'd117} : s = 354;
	{8'd237,8'd118} : s = 355;
	{8'd237,8'd119} : s = 356;
	{8'd237,8'd120} : s = 357;
	{8'd237,8'd121} : s = 358;
	{8'd237,8'd122} : s = 359;
	{8'd237,8'd123} : s = 360;
	{8'd237,8'd124} : s = 361;
	{8'd237,8'd125} : s = 362;
	{8'd237,8'd126} : s = 363;
	{8'd237,8'd127} : s = 364;
	{8'd237,8'd128} : s = 365;
	{8'd237,8'd129} : s = 366;
	{8'd237,8'd130} : s = 367;
	{8'd237,8'd131} : s = 368;
	{8'd237,8'd132} : s = 369;
	{8'd237,8'd133} : s = 370;
	{8'd237,8'd134} : s = 371;
	{8'd237,8'd135} : s = 372;
	{8'd237,8'd136} : s = 373;
	{8'd237,8'd137} : s = 374;
	{8'd237,8'd138} : s = 375;
	{8'd237,8'd139} : s = 376;
	{8'd237,8'd140} : s = 377;
	{8'd237,8'd141} : s = 378;
	{8'd237,8'd142} : s = 379;
	{8'd237,8'd143} : s = 380;
	{8'd237,8'd144} : s = 381;
	{8'd237,8'd145} : s = 382;
	{8'd237,8'd146} : s = 383;
	{8'd237,8'd147} : s = 384;
	{8'd237,8'd148} : s = 385;
	{8'd237,8'd149} : s = 386;
	{8'd237,8'd150} : s = 387;
	{8'd237,8'd151} : s = 388;
	{8'd237,8'd152} : s = 389;
	{8'd237,8'd153} : s = 390;
	{8'd237,8'd154} : s = 391;
	{8'd237,8'd155} : s = 392;
	{8'd237,8'd156} : s = 393;
	{8'd237,8'd157} : s = 394;
	{8'd237,8'd158} : s = 395;
	{8'd237,8'd159} : s = 396;
	{8'd237,8'd160} : s = 397;
	{8'd237,8'd161} : s = 398;
	{8'd237,8'd162} : s = 399;
	{8'd237,8'd163} : s = 400;
	{8'd237,8'd164} : s = 401;
	{8'd237,8'd165} : s = 402;
	{8'd237,8'd166} : s = 403;
	{8'd237,8'd167} : s = 404;
	{8'd237,8'd168} : s = 405;
	{8'd237,8'd169} : s = 406;
	{8'd237,8'd170} : s = 407;
	{8'd237,8'd171} : s = 408;
	{8'd237,8'd172} : s = 409;
	{8'd237,8'd173} : s = 410;
	{8'd237,8'd174} : s = 411;
	{8'd237,8'd175} : s = 412;
	{8'd237,8'd176} : s = 413;
	{8'd237,8'd177} : s = 414;
	{8'd237,8'd178} : s = 415;
	{8'd237,8'd179} : s = 416;
	{8'd237,8'd180} : s = 417;
	{8'd237,8'd181} : s = 418;
	{8'd237,8'd182} : s = 419;
	{8'd237,8'd183} : s = 420;
	{8'd237,8'd184} : s = 421;
	{8'd237,8'd185} : s = 422;
	{8'd237,8'd186} : s = 423;
	{8'd237,8'd187} : s = 424;
	{8'd237,8'd188} : s = 425;
	{8'd237,8'd189} : s = 426;
	{8'd237,8'd190} : s = 427;
	{8'd237,8'd191} : s = 428;
	{8'd237,8'd192} : s = 429;
	{8'd237,8'd193} : s = 430;
	{8'd237,8'd194} : s = 431;
	{8'd237,8'd195} : s = 432;
	{8'd237,8'd196} : s = 433;
	{8'd237,8'd197} : s = 434;
	{8'd237,8'd198} : s = 435;
	{8'd237,8'd199} : s = 436;
	{8'd237,8'd200} : s = 437;
	{8'd237,8'd201} : s = 438;
	{8'd237,8'd202} : s = 439;
	{8'd237,8'd203} : s = 440;
	{8'd237,8'd204} : s = 441;
	{8'd237,8'd205} : s = 442;
	{8'd237,8'd206} : s = 443;
	{8'd237,8'd207} : s = 444;
	{8'd237,8'd208} : s = 445;
	{8'd237,8'd209} : s = 446;
	{8'd237,8'd210} : s = 447;
	{8'd237,8'd211} : s = 448;
	{8'd237,8'd212} : s = 449;
	{8'd237,8'd213} : s = 450;
	{8'd237,8'd214} : s = 451;
	{8'd237,8'd215} : s = 452;
	{8'd237,8'd216} : s = 453;
	{8'd237,8'd217} : s = 454;
	{8'd237,8'd218} : s = 455;
	{8'd237,8'd219} : s = 456;
	{8'd237,8'd220} : s = 457;
	{8'd237,8'd221} : s = 458;
	{8'd237,8'd222} : s = 459;
	{8'd237,8'd223} : s = 460;
	{8'd237,8'd224} : s = 461;
	{8'd237,8'd225} : s = 462;
	{8'd237,8'd226} : s = 463;
	{8'd237,8'd227} : s = 464;
	{8'd237,8'd228} : s = 465;
	{8'd237,8'd229} : s = 466;
	{8'd237,8'd230} : s = 467;
	{8'd237,8'd231} : s = 468;
	{8'd237,8'd232} : s = 469;
	{8'd237,8'd233} : s = 470;
	{8'd237,8'd234} : s = 471;
	{8'd237,8'd235} : s = 472;
	{8'd237,8'd236} : s = 473;
	{8'd237,8'd237} : s = 474;
	{8'd237,8'd238} : s = 475;
	{8'd237,8'd239} : s = 476;
	{8'd237,8'd240} : s = 477;
	{8'd237,8'd241} : s = 478;
	{8'd237,8'd242} : s = 479;
	{8'd237,8'd243} : s = 480;
	{8'd237,8'd244} : s = 481;
	{8'd237,8'd245} : s = 482;
	{8'd237,8'd246} : s = 483;
	{8'd237,8'd247} : s = 484;
	{8'd237,8'd248} : s = 485;
	{8'd237,8'd249} : s = 486;
	{8'd237,8'd250} : s = 487;
	{8'd237,8'd251} : s = 488;
	{8'd237,8'd252} : s = 489;
	{8'd237,8'd253} : s = 490;
	{8'd237,8'd254} : s = 491;
	{8'd237,8'd255} : s = 492;
	{8'd238,8'd0} : s = 238;
	{8'd238,8'd1} : s = 239;
	{8'd238,8'd2} : s = 240;
	{8'd238,8'd3} : s = 241;
	{8'd238,8'd4} : s = 242;
	{8'd238,8'd5} : s = 243;
	{8'd238,8'd6} : s = 244;
	{8'd238,8'd7} : s = 245;
	{8'd238,8'd8} : s = 246;
	{8'd238,8'd9} : s = 247;
	{8'd238,8'd10} : s = 248;
	{8'd238,8'd11} : s = 249;
	{8'd238,8'd12} : s = 250;
	{8'd238,8'd13} : s = 251;
	{8'd238,8'd14} : s = 252;
	{8'd238,8'd15} : s = 253;
	{8'd238,8'd16} : s = 254;
	{8'd238,8'd17} : s = 255;
	{8'd238,8'd18} : s = 256;
	{8'd238,8'd19} : s = 257;
	{8'd238,8'd20} : s = 258;
	{8'd238,8'd21} : s = 259;
	{8'd238,8'd22} : s = 260;
	{8'd238,8'd23} : s = 261;
	{8'd238,8'd24} : s = 262;
	{8'd238,8'd25} : s = 263;
	{8'd238,8'd26} : s = 264;
	{8'd238,8'd27} : s = 265;
	{8'd238,8'd28} : s = 266;
	{8'd238,8'd29} : s = 267;
	{8'd238,8'd30} : s = 268;
	{8'd238,8'd31} : s = 269;
	{8'd238,8'd32} : s = 270;
	{8'd238,8'd33} : s = 271;
	{8'd238,8'd34} : s = 272;
	{8'd238,8'd35} : s = 273;
	{8'd238,8'd36} : s = 274;
	{8'd238,8'd37} : s = 275;
	{8'd238,8'd38} : s = 276;
	{8'd238,8'd39} : s = 277;
	{8'd238,8'd40} : s = 278;
	{8'd238,8'd41} : s = 279;
	{8'd238,8'd42} : s = 280;
	{8'd238,8'd43} : s = 281;
	{8'd238,8'd44} : s = 282;
	{8'd238,8'd45} : s = 283;
	{8'd238,8'd46} : s = 284;
	{8'd238,8'd47} : s = 285;
	{8'd238,8'd48} : s = 286;
	{8'd238,8'd49} : s = 287;
	{8'd238,8'd50} : s = 288;
	{8'd238,8'd51} : s = 289;
	{8'd238,8'd52} : s = 290;
	{8'd238,8'd53} : s = 291;
	{8'd238,8'd54} : s = 292;
	{8'd238,8'd55} : s = 293;
	{8'd238,8'd56} : s = 294;
	{8'd238,8'd57} : s = 295;
	{8'd238,8'd58} : s = 296;
	{8'd238,8'd59} : s = 297;
	{8'd238,8'd60} : s = 298;
	{8'd238,8'd61} : s = 299;
	{8'd238,8'd62} : s = 300;
	{8'd238,8'd63} : s = 301;
	{8'd238,8'd64} : s = 302;
	{8'd238,8'd65} : s = 303;
	{8'd238,8'd66} : s = 304;
	{8'd238,8'd67} : s = 305;
	{8'd238,8'd68} : s = 306;
	{8'd238,8'd69} : s = 307;
	{8'd238,8'd70} : s = 308;
	{8'd238,8'd71} : s = 309;
	{8'd238,8'd72} : s = 310;
	{8'd238,8'd73} : s = 311;
	{8'd238,8'd74} : s = 312;
	{8'd238,8'd75} : s = 313;
	{8'd238,8'd76} : s = 314;
	{8'd238,8'd77} : s = 315;
	{8'd238,8'd78} : s = 316;
	{8'd238,8'd79} : s = 317;
	{8'd238,8'd80} : s = 318;
	{8'd238,8'd81} : s = 319;
	{8'd238,8'd82} : s = 320;
	{8'd238,8'd83} : s = 321;
	{8'd238,8'd84} : s = 322;
	{8'd238,8'd85} : s = 323;
	{8'd238,8'd86} : s = 324;
	{8'd238,8'd87} : s = 325;
	{8'd238,8'd88} : s = 326;
	{8'd238,8'd89} : s = 327;
	{8'd238,8'd90} : s = 328;
	{8'd238,8'd91} : s = 329;
	{8'd238,8'd92} : s = 330;
	{8'd238,8'd93} : s = 331;
	{8'd238,8'd94} : s = 332;
	{8'd238,8'd95} : s = 333;
	{8'd238,8'd96} : s = 334;
	{8'd238,8'd97} : s = 335;
	{8'd238,8'd98} : s = 336;
	{8'd238,8'd99} : s = 337;
	{8'd238,8'd100} : s = 338;
	{8'd238,8'd101} : s = 339;
	{8'd238,8'd102} : s = 340;
	{8'd238,8'd103} : s = 341;
	{8'd238,8'd104} : s = 342;
	{8'd238,8'd105} : s = 343;
	{8'd238,8'd106} : s = 344;
	{8'd238,8'd107} : s = 345;
	{8'd238,8'd108} : s = 346;
	{8'd238,8'd109} : s = 347;
	{8'd238,8'd110} : s = 348;
	{8'd238,8'd111} : s = 349;
	{8'd238,8'd112} : s = 350;
	{8'd238,8'd113} : s = 351;
	{8'd238,8'd114} : s = 352;
	{8'd238,8'd115} : s = 353;
	{8'd238,8'd116} : s = 354;
	{8'd238,8'd117} : s = 355;
	{8'd238,8'd118} : s = 356;
	{8'd238,8'd119} : s = 357;
	{8'd238,8'd120} : s = 358;
	{8'd238,8'd121} : s = 359;
	{8'd238,8'd122} : s = 360;
	{8'd238,8'd123} : s = 361;
	{8'd238,8'd124} : s = 362;
	{8'd238,8'd125} : s = 363;
	{8'd238,8'd126} : s = 364;
	{8'd238,8'd127} : s = 365;
	{8'd238,8'd128} : s = 366;
	{8'd238,8'd129} : s = 367;
	{8'd238,8'd130} : s = 368;
	{8'd238,8'd131} : s = 369;
	{8'd238,8'd132} : s = 370;
	{8'd238,8'd133} : s = 371;
	{8'd238,8'd134} : s = 372;
	{8'd238,8'd135} : s = 373;
	{8'd238,8'd136} : s = 374;
	{8'd238,8'd137} : s = 375;
	{8'd238,8'd138} : s = 376;
	{8'd238,8'd139} : s = 377;
	{8'd238,8'd140} : s = 378;
	{8'd238,8'd141} : s = 379;
	{8'd238,8'd142} : s = 380;
	{8'd238,8'd143} : s = 381;
	{8'd238,8'd144} : s = 382;
	{8'd238,8'd145} : s = 383;
	{8'd238,8'd146} : s = 384;
	{8'd238,8'd147} : s = 385;
	{8'd238,8'd148} : s = 386;
	{8'd238,8'd149} : s = 387;
	{8'd238,8'd150} : s = 388;
	{8'd238,8'd151} : s = 389;
	{8'd238,8'd152} : s = 390;
	{8'd238,8'd153} : s = 391;
	{8'd238,8'd154} : s = 392;
	{8'd238,8'd155} : s = 393;
	{8'd238,8'd156} : s = 394;
	{8'd238,8'd157} : s = 395;
	{8'd238,8'd158} : s = 396;
	{8'd238,8'd159} : s = 397;
	{8'd238,8'd160} : s = 398;
	{8'd238,8'd161} : s = 399;
	{8'd238,8'd162} : s = 400;
	{8'd238,8'd163} : s = 401;
	{8'd238,8'd164} : s = 402;
	{8'd238,8'd165} : s = 403;
	{8'd238,8'd166} : s = 404;
	{8'd238,8'd167} : s = 405;
	{8'd238,8'd168} : s = 406;
	{8'd238,8'd169} : s = 407;
	{8'd238,8'd170} : s = 408;
	{8'd238,8'd171} : s = 409;
	{8'd238,8'd172} : s = 410;
	{8'd238,8'd173} : s = 411;
	{8'd238,8'd174} : s = 412;
	{8'd238,8'd175} : s = 413;
	{8'd238,8'd176} : s = 414;
	{8'd238,8'd177} : s = 415;
	{8'd238,8'd178} : s = 416;
	{8'd238,8'd179} : s = 417;
	{8'd238,8'd180} : s = 418;
	{8'd238,8'd181} : s = 419;
	{8'd238,8'd182} : s = 420;
	{8'd238,8'd183} : s = 421;
	{8'd238,8'd184} : s = 422;
	{8'd238,8'd185} : s = 423;
	{8'd238,8'd186} : s = 424;
	{8'd238,8'd187} : s = 425;
	{8'd238,8'd188} : s = 426;
	{8'd238,8'd189} : s = 427;
	{8'd238,8'd190} : s = 428;
	{8'd238,8'd191} : s = 429;
	{8'd238,8'd192} : s = 430;
	{8'd238,8'd193} : s = 431;
	{8'd238,8'd194} : s = 432;
	{8'd238,8'd195} : s = 433;
	{8'd238,8'd196} : s = 434;
	{8'd238,8'd197} : s = 435;
	{8'd238,8'd198} : s = 436;
	{8'd238,8'd199} : s = 437;
	{8'd238,8'd200} : s = 438;
	{8'd238,8'd201} : s = 439;
	{8'd238,8'd202} : s = 440;
	{8'd238,8'd203} : s = 441;
	{8'd238,8'd204} : s = 442;
	{8'd238,8'd205} : s = 443;
	{8'd238,8'd206} : s = 444;
	{8'd238,8'd207} : s = 445;
	{8'd238,8'd208} : s = 446;
	{8'd238,8'd209} : s = 447;
	{8'd238,8'd210} : s = 448;
	{8'd238,8'd211} : s = 449;
	{8'd238,8'd212} : s = 450;
	{8'd238,8'd213} : s = 451;
	{8'd238,8'd214} : s = 452;
	{8'd238,8'd215} : s = 453;
	{8'd238,8'd216} : s = 454;
	{8'd238,8'd217} : s = 455;
	{8'd238,8'd218} : s = 456;
	{8'd238,8'd219} : s = 457;
	{8'd238,8'd220} : s = 458;
	{8'd238,8'd221} : s = 459;
	{8'd238,8'd222} : s = 460;
	{8'd238,8'd223} : s = 461;
	{8'd238,8'd224} : s = 462;
	{8'd238,8'd225} : s = 463;
	{8'd238,8'd226} : s = 464;
	{8'd238,8'd227} : s = 465;
	{8'd238,8'd228} : s = 466;
	{8'd238,8'd229} : s = 467;
	{8'd238,8'd230} : s = 468;
	{8'd238,8'd231} : s = 469;
	{8'd238,8'd232} : s = 470;
	{8'd238,8'd233} : s = 471;
	{8'd238,8'd234} : s = 472;
	{8'd238,8'd235} : s = 473;
	{8'd238,8'd236} : s = 474;
	{8'd238,8'd237} : s = 475;
	{8'd238,8'd238} : s = 476;
	{8'd238,8'd239} : s = 477;
	{8'd238,8'd240} : s = 478;
	{8'd238,8'd241} : s = 479;
	{8'd238,8'd242} : s = 480;
	{8'd238,8'd243} : s = 481;
	{8'd238,8'd244} : s = 482;
	{8'd238,8'd245} : s = 483;
	{8'd238,8'd246} : s = 484;
	{8'd238,8'd247} : s = 485;
	{8'd238,8'd248} : s = 486;
	{8'd238,8'd249} : s = 487;
	{8'd238,8'd250} : s = 488;
	{8'd238,8'd251} : s = 489;
	{8'd238,8'd252} : s = 490;
	{8'd238,8'd253} : s = 491;
	{8'd238,8'd254} : s = 492;
	{8'd238,8'd255} : s = 493;
	{8'd239,8'd0} : s = 239;
	{8'd239,8'd1} : s = 240;
	{8'd239,8'd2} : s = 241;
	{8'd239,8'd3} : s = 242;
	{8'd239,8'd4} : s = 243;
	{8'd239,8'd5} : s = 244;
	{8'd239,8'd6} : s = 245;
	{8'd239,8'd7} : s = 246;
	{8'd239,8'd8} : s = 247;
	{8'd239,8'd9} : s = 248;
	{8'd239,8'd10} : s = 249;
	{8'd239,8'd11} : s = 250;
	{8'd239,8'd12} : s = 251;
	{8'd239,8'd13} : s = 252;
	{8'd239,8'd14} : s = 253;
	{8'd239,8'd15} : s = 254;
	{8'd239,8'd16} : s = 255;
	{8'd239,8'd17} : s = 256;
	{8'd239,8'd18} : s = 257;
	{8'd239,8'd19} : s = 258;
	{8'd239,8'd20} : s = 259;
	{8'd239,8'd21} : s = 260;
	{8'd239,8'd22} : s = 261;
	{8'd239,8'd23} : s = 262;
	{8'd239,8'd24} : s = 263;
	{8'd239,8'd25} : s = 264;
	{8'd239,8'd26} : s = 265;
	{8'd239,8'd27} : s = 266;
	{8'd239,8'd28} : s = 267;
	{8'd239,8'd29} : s = 268;
	{8'd239,8'd30} : s = 269;
	{8'd239,8'd31} : s = 270;
	{8'd239,8'd32} : s = 271;
	{8'd239,8'd33} : s = 272;
	{8'd239,8'd34} : s = 273;
	{8'd239,8'd35} : s = 274;
	{8'd239,8'd36} : s = 275;
	{8'd239,8'd37} : s = 276;
	{8'd239,8'd38} : s = 277;
	{8'd239,8'd39} : s = 278;
	{8'd239,8'd40} : s = 279;
	{8'd239,8'd41} : s = 280;
	{8'd239,8'd42} : s = 281;
	{8'd239,8'd43} : s = 282;
	{8'd239,8'd44} : s = 283;
	{8'd239,8'd45} : s = 284;
	{8'd239,8'd46} : s = 285;
	{8'd239,8'd47} : s = 286;
	{8'd239,8'd48} : s = 287;
	{8'd239,8'd49} : s = 288;
	{8'd239,8'd50} : s = 289;
	{8'd239,8'd51} : s = 290;
	{8'd239,8'd52} : s = 291;
	{8'd239,8'd53} : s = 292;
	{8'd239,8'd54} : s = 293;
	{8'd239,8'd55} : s = 294;
	{8'd239,8'd56} : s = 295;
	{8'd239,8'd57} : s = 296;
	{8'd239,8'd58} : s = 297;
	{8'd239,8'd59} : s = 298;
	{8'd239,8'd60} : s = 299;
	{8'd239,8'd61} : s = 300;
	{8'd239,8'd62} : s = 301;
	{8'd239,8'd63} : s = 302;
	{8'd239,8'd64} : s = 303;
	{8'd239,8'd65} : s = 304;
	{8'd239,8'd66} : s = 305;
	{8'd239,8'd67} : s = 306;
	{8'd239,8'd68} : s = 307;
	{8'd239,8'd69} : s = 308;
	{8'd239,8'd70} : s = 309;
	{8'd239,8'd71} : s = 310;
	{8'd239,8'd72} : s = 311;
	{8'd239,8'd73} : s = 312;
	{8'd239,8'd74} : s = 313;
	{8'd239,8'd75} : s = 314;
	{8'd239,8'd76} : s = 315;
	{8'd239,8'd77} : s = 316;
	{8'd239,8'd78} : s = 317;
	{8'd239,8'd79} : s = 318;
	{8'd239,8'd80} : s = 319;
	{8'd239,8'd81} : s = 320;
	{8'd239,8'd82} : s = 321;
	{8'd239,8'd83} : s = 322;
	{8'd239,8'd84} : s = 323;
	{8'd239,8'd85} : s = 324;
	{8'd239,8'd86} : s = 325;
	{8'd239,8'd87} : s = 326;
	{8'd239,8'd88} : s = 327;
	{8'd239,8'd89} : s = 328;
	{8'd239,8'd90} : s = 329;
	{8'd239,8'd91} : s = 330;
	{8'd239,8'd92} : s = 331;
	{8'd239,8'd93} : s = 332;
	{8'd239,8'd94} : s = 333;
	{8'd239,8'd95} : s = 334;
	{8'd239,8'd96} : s = 335;
	{8'd239,8'd97} : s = 336;
	{8'd239,8'd98} : s = 337;
	{8'd239,8'd99} : s = 338;
	{8'd239,8'd100} : s = 339;
	{8'd239,8'd101} : s = 340;
	{8'd239,8'd102} : s = 341;
	{8'd239,8'd103} : s = 342;
	{8'd239,8'd104} : s = 343;
	{8'd239,8'd105} : s = 344;
	{8'd239,8'd106} : s = 345;
	{8'd239,8'd107} : s = 346;
	{8'd239,8'd108} : s = 347;
	{8'd239,8'd109} : s = 348;
	{8'd239,8'd110} : s = 349;
	{8'd239,8'd111} : s = 350;
	{8'd239,8'd112} : s = 351;
	{8'd239,8'd113} : s = 352;
	{8'd239,8'd114} : s = 353;
	{8'd239,8'd115} : s = 354;
	{8'd239,8'd116} : s = 355;
	{8'd239,8'd117} : s = 356;
	{8'd239,8'd118} : s = 357;
	{8'd239,8'd119} : s = 358;
	{8'd239,8'd120} : s = 359;
	{8'd239,8'd121} : s = 360;
	{8'd239,8'd122} : s = 361;
	{8'd239,8'd123} : s = 362;
	{8'd239,8'd124} : s = 363;
	{8'd239,8'd125} : s = 364;
	{8'd239,8'd126} : s = 365;
	{8'd239,8'd127} : s = 366;
	{8'd239,8'd128} : s = 367;
	{8'd239,8'd129} : s = 368;
	{8'd239,8'd130} : s = 369;
	{8'd239,8'd131} : s = 370;
	{8'd239,8'd132} : s = 371;
	{8'd239,8'd133} : s = 372;
	{8'd239,8'd134} : s = 373;
	{8'd239,8'd135} : s = 374;
	{8'd239,8'd136} : s = 375;
	{8'd239,8'd137} : s = 376;
	{8'd239,8'd138} : s = 377;
	{8'd239,8'd139} : s = 378;
	{8'd239,8'd140} : s = 379;
	{8'd239,8'd141} : s = 380;
	{8'd239,8'd142} : s = 381;
	{8'd239,8'd143} : s = 382;
	{8'd239,8'd144} : s = 383;
	{8'd239,8'd145} : s = 384;
	{8'd239,8'd146} : s = 385;
	{8'd239,8'd147} : s = 386;
	{8'd239,8'd148} : s = 387;
	{8'd239,8'd149} : s = 388;
	{8'd239,8'd150} : s = 389;
	{8'd239,8'd151} : s = 390;
	{8'd239,8'd152} : s = 391;
	{8'd239,8'd153} : s = 392;
	{8'd239,8'd154} : s = 393;
	{8'd239,8'd155} : s = 394;
	{8'd239,8'd156} : s = 395;
	{8'd239,8'd157} : s = 396;
	{8'd239,8'd158} : s = 397;
	{8'd239,8'd159} : s = 398;
	{8'd239,8'd160} : s = 399;
	{8'd239,8'd161} : s = 400;
	{8'd239,8'd162} : s = 401;
	{8'd239,8'd163} : s = 402;
	{8'd239,8'd164} : s = 403;
	{8'd239,8'd165} : s = 404;
	{8'd239,8'd166} : s = 405;
	{8'd239,8'd167} : s = 406;
	{8'd239,8'd168} : s = 407;
	{8'd239,8'd169} : s = 408;
	{8'd239,8'd170} : s = 409;
	{8'd239,8'd171} : s = 410;
	{8'd239,8'd172} : s = 411;
	{8'd239,8'd173} : s = 412;
	{8'd239,8'd174} : s = 413;
	{8'd239,8'd175} : s = 414;
	{8'd239,8'd176} : s = 415;
	{8'd239,8'd177} : s = 416;
	{8'd239,8'd178} : s = 417;
	{8'd239,8'd179} : s = 418;
	{8'd239,8'd180} : s = 419;
	{8'd239,8'd181} : s = 420;
	{8'd239,8'd182} : s = 421;
	{8'd239,8'd183} : s = 422;
	{8'd239,8'd184} : s = 423;
	{8'd239,8'd185} : s = 424;
	{8'd239,8'd186} : s = 425;
	{8'd239,8'd187} : s = 426;
	{8'd239,8'd188} : s = 427;
	{8'd239,8'd189} : s = 428;
	{8'd239,8'd190} : s = 429;
	{8'd239,8'd191} : s = 430;
	{8'd239,8'd192} : s = 431;
	{8'd239,8'd193} : s = 432;
	{8'd239,8'd194} : s = 433;
	{8'd239,8'd195} : s = 434;
	{8'd239,8'd196} : s = 435;
	{8'd239,8'd197} : s = 436;
	{8'd239,8'd198} : s = 437;
	{8'd239,8'd199} : s = 438;
	{8'd239,8'd200} : s = 439;
	{8'd239,8'd201} : s = 440;
	{8'd239,8'd202} : s = 441;
	{8'd239,8'd203} : s = 442;
	{8'd239,8'd204} : s = 443;
	{8'd239,8'd205} : s = 444;
	{8'd239,8'd206} : s = 445;
	{8'd239,8'd207} : s = 446;
	{8'd239,8'd208} : s = 447;
	{8'd239,8'd209} : s = 448;
	{8'd239,8'd210} : s = 449;
	{8'd239,8'd211} : s = 450;
	{8'd239,8'd212} : s = 451;
	{8'd239,8'd213} : s = 452;
	{8'd239,8'd214} : s = 453;
	{8'd239,8'd215} : s = 454;
	{8'd239,8'd216} : s = 455;
	{8'd239,8'd217} : s = 456;
	{8'd239,8'd218} : s = 457;
	{8'd239,8'd219} : s = 458;
	{8'd239,8'd220} : s = 459;
	{8'd239,8'd221} : s = 460;
	{8'd239,8'd222} : s = 461;
	{8'd239,8'd223} : s = 462;
	{8'd239,8'd224} : s = 463;
	{8'd239,8'd225} : s = 464;
	{8'd239,8'd226} : s = 465;
	{8'd239,8'd227} : s = 466;
	{8'd239,8'd228} : s = 467;
	{8'd239,8'd229} : s = 468;
	{8'd239,8'd230} : s = 469;
	{8'd239,8'd231} : s = 470;
	{8'd239,8'd232} : s = 471;
	{8'd239,8'd233} : s = 472;
	{8'd239,8'd234} : s = 473;
	{8'd239,8'd235} : s = 474;
	{8'd239,8'd236} : s = 475;
	{8'd239,8'd237} : s = 476;
	{8'd239,8'd238} : s = 477;
	{8'd239,8'd239} : s = 478;
	{8'd239,8'd240} : s = 479;
	{8'd239,8'd241} : s = 480;
	{8'd239,8'd242} : s = 481;
	{8'd239,8'd243} : s = 482;
	{8'd239,8'd244} : s = 483;
	{8'd239,8'd245} : s = 484;
	{8'd239,8'd246} : s = 485;
	{8'd239,8'd247} : s = 486;
	{8'd239,8'd248} : s = 487;
	{8'd239,8'd249} : s = 488;
	{8'd239,8'd250} : s = 489;
	{8'd239,8'd251} : s = 490;
	{8'd239,8'd252} : s = 491;
	{8'd239,8'd253} : s = 492;
	{8'd239,8'd254} : s = 493;
	{8'd239,8'd255} : s = 494;
	{8'd240,8'd0} : s = 240;
	{8'd240,8'd1} : s = 241;
	{8'd240,8'd2} : s = 242;
	{8'd240,8'd3} : s = 243;
	{8'd240,8'd4} : s = 244;
	{8'd240,8'd5} : s = 245;
	{8'd240,8'd6} : s = 246;
	{8'd240,8'd7} : s = 247;
	{8'd240,8'd8} : s = 248;
	{8'd240,8'd9} : s = 249;
	{8'd240,8'd10} : s = 250;
	{8'd240,8'd11} : s = 251;
	{8'd240,8'd12} : s = 252;
	{8'd240,8'd13} : s = 253;
	{8'd240,8'd14} : s = 254;
	{8'd240,8'd15} : s = 255;
	{8'd240,8'd16} : s = 256;
	{8'd240,8'd17} : s = 257;
	{8'd240,8'd18} : s = 258;
	{8'd240,8'd19} : s = 259;
	{8'd240,8'd20} : s = 260;
	{8'd240,8'd21} : s = 261;
	{8'd240,8'd22} : s = 262;
	{8'd240,8'd23} : s = 263;
	{8'd240,8'd24} : s = 264;
	{8'd240,8'd25} : s = 265;
	{8'd240,8'd26} : s = 266;
	{8'd240,8'd27} : s = 267;
	{8'd240,8'd28} : s = 268;
	{8'd240,8'd29} : s = 269;
	{8'd240,8'd30} : s = 270;
	{8'd240,8'd31} : s = 271;
	{8'd240,8'd32} : s = 272;
	{8'd240,8'd33} : s = 273;
	{8'd240,8'd34} : s = 274;
	{8'd240,8'd35} : s = 275;
	{8'd240,8'd36} : s = 276;
	{8'd240,8'd37} : s = 277;
	{8'd240,8'd38} : s = 278;
	{8'd240,8'd39} : s = 279;
	{8'd240,8'd40} : s = 280;
	{8'd240,8'd41} : s = 281;
	{8'd240,8'd42} : s = 282;
	{8'd240,8'd43} : s = 283;
	{8'd240,8'd44} : s = 284;
	{8'd240,8'd45} : s = 285;
	{8'd240,8'd46} : s = 286;
	{8'd240,8'd47} : s = 287;
	{8'd240,8'd48} : s = 288;
	{8'd240,8'd49} : s = 289;
	{8'd240,8'd50} : s = 290;
	{8'd240,8'd51} : s = 291;
	{8'd240,8'd52} : s = 292;
	{8'd240,8'd53} : s = 293;
	{8'd240,8'd54} : s = 294;
	{8'd240,8'd55} : s = 295;
	{8'd240,8'd56} : s = 296;
	{8'd240,8'd57} : s = 297;
	{8'd240,8'd58} : s = 298;
	{8'd240,8'd59} : s = 299;
	{8'd240,8'd60} : s = 300;
	{8'd240,8'd61} : s = 301;
	{8'd240,8'd62} : s = 302;
	{8'd240,8'd63} : s = 303;
	{8'd240,8'd64} : s = 304;
	{8'd240,8'd65} : s = 305;
	{8'd240,8'd66} : s = 306;
	{8'd240,8'd67} : s = 307;
	{8'd240,8'd68} : s = 308;
	{8'd240,8'd69} : s = 309;
	{8'd240,8'd70} : s = 310;
	{8'd240,8'd71} : s = 311;
	{8'd240,8'd72} : s = 312;
	{8'd240,8'd73} : s = 313;
	{8'd240,8'd74} : s = 314;
	{8'd240,8'd75} : s = 315;
	{8'd240,8'd76} : s = 316;
	{8'd240,8'd77} : s = 317;
	{8'd240,8'd78} : s = 318;
	{8'd240,8'd79} : s = 319;
	{8'd240,8'd80} : s = 320;
	{8'd240,8'd81} : s = 321;
	{8'd240,8'd82} : s = 322;
	{8'd240,8'd83} : s = 323;
	{8'd240,8'd84} : s = 324;
	{8'd240,8'd85} : s = 325;
	{8'd240,8'd86} : s = 326;
	{8'd240,8'd87} : s = 327;
	{8'd240,8'd88} : s = 328;
	{8'd240,8'd89} : s = 329;
	{8'd240,8'd90} : s = 330;
	{8'd240,8'd91} : s = 331;
	{8'd240,8'd92} : s = 332;
	{8'd240,8'd93} : s = 333;
	{8'd240,8'd94} : s = 334;
	{8'd240,8'd95} : s = 335;
	{8'd240,8'd96} : s = 336;
	{8'd240,8'd97} : s = 337;
	{8'd240,8'd98} : s = 338;
	{8'd240,8'd99} : s = 339;
	{8'd240,8'd100} : s = 340;
	{8'd240,8'd101} : s = 341;
	{8'd240,8'd102} : s = 342;
	{8'd240,8'd103} : s = 343;
	{8'd240,8'd104} : s = 344;
	{8'd240,8'd105} : s = 345;
	{8'd240,8'd106} : s = 346;
	{8'd240,8'd107} : s = 347;
	{8'd240,8'd108} : s = 348;
	{8'd240,8'd109} : s = 349;
	{8'd240,8'd110} : s = 350;
	{8'd240,8'd111} : s = 351;
	{8'd240,8'd112} : s = 352;
	{8'd240,8'd113} : s = 353;
	{8'd240,8'd114} : s = 354;
	{8'd240,8'd115} : s = 355;
	{8'd240,8'd116} : s = 356;
	{8'd240,8'd117} : s = 357;
	{8'd240,8'd118} : s = 358;
	{8'd240,8'd119} : s = 359;
	{8'd240,8'd120} : s = 360;
	{8'd240,8'd121} : s = 361;
	{8'd240,8'd122} : s = 362;
	{8'd240,8'd123} : s = 363;
	{8'd240,8'd124} : s = 364;
	{8'd240,8'd125} : s = 365;
	{8'd240,8'd126} : s = 366;
	{8'd240,8'd127} : s = 367;
	{8'd240,8'd128} : s = 368;
	{8'd240,8'd129} : s = 369;
	{8'd240,8'd130} : s = 370;
	{8'd240,8'd131} : s = 371;
	{8'd240,8'd132} : s = 372;
	{8'd240,8'd133} : s = 373;
	{8'd240,8'd134} : s = 374;
	{8'd240,8'd135} : s = 375;
	{8'd240,8'd136} : s = 376;
	{8'd240,8'd137} : s = 377;
	{8'd240,8'd138} : s = 378;
	{8'd240,8'd139} : s = 379;
	{8'd240,8'd140} : s = 380;
	{8'd240,8'd141} : s = 381;
	{8'd240,8'd142} : s = 382;
	{8'd240,8'd143} : s = 383;
	{8'd240,8'd144} : s = 384;
	{8'd240,8'd145} : s = 385;
	{8'd240,8'd146} : s = 386;
	{8'd240,8'd147} : s = 387;
	{8'd240,8'd148} : s = 388;
	{8'd240,8'd149} : s = 389;
	{8'd240,8'd150} : s = 390;
	{8'd240,8'd151} : s = 391;
	{8'd240,8'd152} : s = 392;
	{8'd240,8'd153} : s = 393;
	{8'd240,8'd154} : s = 394;
	{8'd240,8'd155} : s = 395;
	{8'd240,8'd156} : s = 396;
	{8'd240,8'd157} : s = 397;
	{8'd240,8'd158} : s = 398;
	{8'd240,8'd159} : s = 399;
	{8'd240,8'd160} : s = 400;
	{8'd240,8'd161} : s = 401;
	{8'd240,8'd162} : s = 402;
	{8'd240,8'd163} : s = 403;
	{8'd240,8'd164} : s = 404;
	{8'd240,8'd165} : s = 405;
	{8'd240,8'd166} : s = 406;
	{8'd240,8'd167} : s = 407;
	{8'd240,8'd168} : s = 408;
	{8'd240,8'd169} : s = 409;
	{8'd240,8'd170} : s = 410;
	{8'd240,8'd171} : s = 411;
	{8'd240,8'd172} : s = 412;
	{8'd240,8'd173} : s = 413;
	{8'd240,8'd174} : s = 414;
	{8'd240,8'd175} : s = 415;
	{8'd240,8'd176} : s = 416;
	{8'd240,8'd177} : s = 417;
	{8'd240,8'd178} : s = 418;
	{8'd240,8'd179} : s = 419;
	{8'd240,8'd180} : s = 420;
	{8'd240,8'd181} : s = 421;
	{8'd240,8'd182} : s = 422;
	{8'd240,8'd183} : s = 423;
	{8'd240,8'd184} : s = 424;
	{8'd240,8'd185} : s = 425;
	{8'd240,8'd186} : s = 426;
	{8'd240,8'd187} : s = 427;
	{8'd240,8'd188} : s = 428;
	{8'd240,8'd189} : s = 429;
	{8'd240,8'd190} : s = 430;
	{8'd240,8'd191} : s = 431;
	{8'd240,8'd192} : s = 432;
	{8'd240,8'd193} : s = 433;
	{8'd240,8'd194} : s = 434;
	{8'd240,8'd195} : s = 435;
	{8'd240,8'd196} : s = 436;
	{8'd240,8'd197} : s = 437;
	{8'd240,8'd198} : s = 438;
	{8'd240,8'd199} : s = 439;
	{8'd240,8'd200} : s = 440;
	{8'd240,8'd201} : s = 441;
	{8'd240,8'd202} : s = 442;
	{8'd240,8'd203} : s = 443;
	{8'd240,8'd204} : s = 444;
	{8'd240,8'd205} : s = 445;
	{8'd240,8'd206} : s = 446;
	{8'd240,8'd207} : s = 447;
	{8'd240,8'd208} : s = 448;
	{8'd240,8'd209} : s = 449;
	{8'd240,8'd210} : s = 450;
	{8'd240,8'd211} : s = 451;
	{8'd240,8'd212} : s = 452;
	{8'd240,8'd213} : s = 453;
	{8'd240,8'd214} : s = 454;
	{8'd240,8'd215} : s = 455;
	{8'd240,8'd216} : s = 456;
	{8'd240,8'd217} : s = 457;
	{8'd240,8'd218} : s = 458;
	{8'd240,8'd219} : s = 459;
	{8'd240,8'd220} : s = 460;
	{8'd240,8'd221} : s = 461;
	{8'd240,8'd222} : s = 462;
	{8'd240,8'd223} : s = 463;
	{8'd240,8'd224} : s = 464;
	{8'd240,8'd225} : s = 465;
	{8'd240,8'd226} : s = 466;
	{8'd240,8'd227} : s = 467;
	{8'd240,8'd228} : s = 468;
	{8'd240,8'd229} : s = 469;
	{8'd240,8'd230} : s = 470;
	{8'd240,8'd231} : s = 471;
	{8'd240,8'd232} : s = 472;
	{8'd240,8'd233} : s = 473;
	{8'd240,8'd234} : s = 474;
	{8'd240,8'd235} : s = 475;
	{8'd240,8'd236} : s = 476;
	{8'd240,8'd237} : s = 477;
	{8'd240,8'd238} : s = 478;
	{8'd240,8'd239} : s = 479;
	{8'd240,8'd240} : s = 480;
	{8'd240,8'd241} : s = 481;
	{8'd240,8'd242} : s = 482;
	{8'd240,8'd243} : s = 483;
	{8'd240,8'd244} : s = 484;
	{8'd240,8'd245} : s = 485;
	{8'd240,8'd246} : s = 486;
	{8'd240,8'd247} : s = 487;
	{8'd240,8'd248} : s = 488;
	{8'd240,8'd249} : s = 489;
	{8'd240,8'd250} : s = 490;
	{8'd240,8'd251} : s = 491;
	{8'd240,8'd252} : s = 492;
	{8'd240,8'd253} : s = 493;
	{8'd240,8'd254} : s = 494;
	{8'd240,8'd255} : s = 495;
	{8'd241,8'd0} : s = 241;
	{8'd241,8'd1} : s = 242;
	{8'd241,8'd2} : s = 243;
	{8'd241,8'd3} : s = 244;
	{8'd241,8'd4} : s = 245;
	{8'd241,8'd5} : s = 246;
	{8'd241,8'd6} : s = 247;
	{8'd241,8'd7} : s = 248;
	{8'd241,8'd8} : s = 249;
	{8'd241,8'd9} : s = 250;
	{8'd241,8'd10} : s = 251;
	{8'd241,8'd11} : s = 252;
	{8'd241,8'd12} : s = 253;
	{8'd241,8'd13} : s = 254;
	{8'd241,8'd14} : s = 255;
	{8'd241,8'd15} : s = 256;
	{8'd241,8'd16} : s = 257;
	{8'd241,8'd17} : s = 258;
	{8'd241,8'd18} : s = 259;
	{8'd241,8'd19} : s = 260;
	{8'd241,8'd20} : s = 261;
	{8'd241,8'd21} : s = 262;
	{8'd241,8'd22} : s = 263;
	{8'd241,8'd23} : s = 264;
	{8'd241,8'd24} : s = 265;
	{8'd241,8'd25} : s = 266;
	{8'd241,8'd26} : s = 267;
	{8'd241,8'd27} : s = 268;
	{8'd241,8'd28} : s = 269;
	{8'd241,8'd29} : s = 270;
	{8'd241,8'd30} : s = 271;
	{8'd241,8'd31} : s = 272;
	{8'd241,8'd32} : s = 273;
	{8'd241,8'd33} : s = 274;
	{8'd241,8'd34} : s = 275;
	{8'd241,8'd35} : s = 276;
	{8'd241,8'd36} : s = 277;
	{8'd241,8'd37} : s = 278;
	{8'd241,8'd38} : s = 279;
	{8'd241,8'd39} : s = 280;
	{8'd241,8'd40} : s = 281;
	{8'd241,8'd41} : s = 282;
	{8'd241,8'd42} : s = 283;
	{8'd241,8'd43} : s = 284;
	{8'd241,8'd44} : s = 285;
	{8'd241,8'd45} : s = 286;
	{8'd241,8'd46} : s = 287;
	{8'd241,8'd47} : s = 288;
	{8'd241,8'd48} : s = 289;
	{8'd241,8'd49} : s = 290;
	{8'd241,8'd50} : s = 291;
	{8'd241,8'd51} : s = 292;
	{8'd241,8'd52} : s = 293;
	{8'd241,8'd53} : s = 294;
	{8'd241,8'd54} : s = 295;
	{8'd241,8'd55} : s = 296;
	{8'd241,8'd56} : s = 297;
	{8'd241,8'd57} : s = 298;
	{8'd241,8'd58} : s = 299;
	{8'd241,8'd59} : s = 300;
	{8'd241,8'd60} : s = 301;
	{8'd241,8'd61} : s = 302;
	{8'd241,8'd62} : s = 303;
	{8'd241,8'd63} : s = 304;
	{8'd241,8'd64} : s = 305;
	{8'd241,8'd65} : s = 306;
	{8'd241,8'd66} : s = 307;
	{8'd241,8'd67} : s = 308;
	{8'd241,8'd68} : s = 309;
	{8'd241,8'd69} : s = 310;
	{8'd241,8'd70} : s = 311;
	{8'd241,8'd71} : s = 312;
	{8'd241,8'd72} : s = 313;
	{8'd241,8'd73} : s = 314;
	{8'd241,8'd74} : s = 315;
	{8'd241,8'd75} : s = 316;
	{8'd241,8'd76} : s = 317;
	{8'd241,8'd77} : s = 318;
	{8'd241,8'd78} : s = 319;
	{8'd241,8'd79} : s = 320;
	{8'd241,8'd80} : s = 321;
	{8'd241,8'd81} : s = 322;
	{8'd241,8'd82} : s = 323;
	{8'd241,8'd83} : s = 324;
	{8'd241,8'd84} : s = 325;
	{8'd241,8'd85} : s = 326;
	{8'd241,8'd86} : s = 327;
	{8'd241,8'd87} : s = 328;
	{8'd241,8'd88} : s = 329;
	{8'd241,8'd89} : s = 330;
	{8'd241,8'd90} : s = 331;
	{8'd241,8'd91} : s = 332;
	{8'd241,8'd92} : s = 333;
	{8'd241,8'd93} : s = 334;
	{8'd241,8'd94} : s = 335;
	{8'd241,8'd95} : s = 336;
	{8'd241,8'd96} : s = 337;
	{8'd241,8'd97} : s = 338;
	{8'd241,8'd98} : s = 339;
	{8'd241,8'd99} : s = 340;
	{8'd241,8'd100} : s = 341;
	{8'd241,8'd101} : s = 342;
	{8'd241,8'd102} : s = 343;
	{8'd241,8'd103} : s = 344;
	{8'd241,8'd104} : s = 345;
	{8'd241,8'd105} : s = 346;
	{8'd241,8'd106} : s = 347;
	{8'd241,8'd107} : s = 348;
	{8'd241,8'd108} : s = 349;
	{8'd241,8'd109} : s = 350;
	{8'd241,8'd110} : s = 351;
	{8'd241,8'd111} : s = 352;
	{8'd241,8'd112} : s = 353;
	{8'd241,8'd113} : s = 354;
	{8'd241,8'd114} : s = 355;
	{8'd241,8'd115} : s = 356;
	{8'd241,8'd116} : s = 357;
	{8'd241,8'd117} : s = 358;
	{8'd241,8'd118} : s = 359;
	{8'd241,8'd119} : s = 360;
	{8'd241,8'd120} : s = 361;
	{8'd241,8'd121} : s = 362;
	{8'd241,8'd122} : s = 363;
	{8'd241,8'd123} : s = 364;
	{8'd241,8'd124} : s = 365;
	{8'd241,8'd125} : s = 366;
	{8'd241,8'd126} : s = 367;
	{8'd241,8'd127} : s = 368;
	{8'd241,8'd128} : s = 369;
	{8'd241,8'd129} : s = 370;
	{8'd241,8'd130} : s = 371;
	{8'd241,8'd131} : s = 372;
	{8'd241,8'd132} : s = 373;
	{8'd241,8'd133} : s = 374;
	{8'd241,8'd134} : s = 375;
	{8'd241,8'd135} : s = 376;
	{8'd241,8'd136} : s = 377;
	{8'd241,8'd137} : s = 378;
	{8'd241,8'd138} : s = 379;
	{8'd241,8'd139} : s = 380;
	{8'd241,8'd140} : s = 381;
	{8'd241,8'd141} : s = 382;
	{8'd241,8'd142} : s = 383;
	{8'd241,8'd143} : s = 384;
	{8'd241,8'd144} : s = 385;
	{8'd241,8'd145} : s = 386;
	{8'd241,8'd146} : s = 387;
	{8'd241,8'd147} : s = 388;
	{8'd241,8'd148} : s = 389;
	{8'd241,8'd149} : s = 390;
	{8'd241,8'd150} : s = 391;
	{8'd241,8'd151} : s = 392;
	{8'd241,8'd152} : s = 393;
	{8'd241,8'd153} : s = 394;
	{8'd241,8'd154} : s = 395;
	{8'd241,8'd155} : s = 396;
	{8'd241,8'd156} : s = 397;
	{8'd241,8'd157} : s = 398;
	{8'd241,8'd158} : s = 399;
	{8'd241,8'd159} : s = 400;
	{8'd241,8'd160} : s = 401;
	{8'd241,8'd161} : s = 402;
	{8'd241,8'd162} : s = 403;
	{8'd241,8'd163} : s = 404;
	{8'd241,8'd164} : s = 405;
	{8'd241,8'd165} : s = 406;
	{8'd241,8'd166} : s = 407;
	{8'd241,8'd167} : s = 408;
	{8'd241,8'd168} : s = 409;
	{8'd241,8'd169} : s = 410;
	{8'd241,8'd170} : s = 411;
	{8'd241,8'd171} : s = 412;
	{8'd241,8'd172} : s = 413;
	{8'd241,8'd173} : s = 414;
	{8'd241,8'd174} : s = 415;
	{8'd241,8'd175} : s = 416;
	{8'd241,8'd176} : s = 417;
	{8'd241,8'd177} : s = 418;
	{8'd241,8'd178} : s = 419;
	{8'd241,8'd179} : s = 420;
	{8'd241,8'd180} : s = 421;
	{8'd241,8'd181} : s = 422;
	{8'd241,8'd182} : s = 423;
	{8'd241,8'd183} : s = 424;
	{8'd241,8'd184} : s = 425;
	{8'd241,8'd185} : s = 426;
	{8'd241,8'd186} : s = 427;
	{8'd241,8'd187} : s = 428;
	{8'd241,8'd188} : s = 429;
	{8'd241,8'd189} : s = 430;
	{8'd241,8'd190} : s = 431;
	{8'd241,8'd191} : s = 432;
	{8'd241,8'd192} : s = 433;
	{8'd241,8'd193} : s = 434;
	{8'd241,8'd194} : s = 435;
	{8'd241,8'd195} : s = 436;
	{8'd241,8'd196} : s = 437;
	{8'd241,8'd197} : s = 438;
	{8'd241,8'd198} : s = 439;
	{8'd241,8'd199} : s = 440;
	{8'd241,8'd200} : s = 441;
	{8'd241,8'd201} : s = 442;
	{8'd241,8'd202} : s = 443;
	{8'd241,8'd203} : s = 444;
	{8'd241,8'd204} : s = 445;
	{8'd241,8'd205} : s = 446;
	{8'd241,8'd206} : s = 447;
	{8'd241,8'd207} : s = 448;
	{8'd241,8'd208} : s = 449;
	{8'd241,8'd209} : s = 450;
	{8'd241,8'd210} : s = 451;
	{8'd241,8'd211} : s = 452;
	{8'd241,8'd212} : s = 453;
	{8'd241,8'd213} : s = 454;
	{8'd241,8'd214} : s = 455;
	{8'd241,8'd215} : s = 456;
	{8'd241,8'd216} : s = 457;
	{8'd241,8'd217} : s = 458;
	{8'd241,8'd218} : s = 459;
	{8'd241,8'd219} : s = 460;
	{8'd241,8'd220} : s = 461;
	{8'd241,8'd221} : s = 462;
	{8'd241,8'd222} : s = 463;
	{8'd241,8'd223} : s = 464;
	{8'd241,8'd224} : s = 465;
	{8'd241,8'd225} : s = 466;
	{8'd241,8'd226} : s = 467;
	{8'd241,8'd227} : s = 468;
	{8'd241,8'd228} : s = 469;
	{8'd241,8'd229} : s = 470;
	{8'd241,8'd230} : s = 471;
	{8'd241,8'd231} : s = 472;
	{8'd241,8'd232} : s = 473;
	{8'd241,8'd233} : s = 474;
	{8'd241,8'd234} : s = 475;
	{8'd241,8'd235} : s = 476;
	{8'd241,8'd236} : s = 477;
	{8'd241,8'd237} : s = 478;
	{8'd241,8'd238} : s = 479;
	{8'd241,8'd239} : s = 480;
	{8'd241,8'd240} : s = 481;
	{8'd241,8'd241} : s = 482;
	{8'd241,8'd242} : s = 483;
	{8'd241,8'd243} : s = 484;
	{8'd241,8'd244} : s = 485;
	{8'd241,8'd245} : s = 486;
	{8'd241,8'd246} : s = 487;
	{8'd241,8'd247} : s = 488;
	{8'd241,8'd248} : s = 489;
	{8'd241,8'd249} : s = 490;
	{8'd241,8'd250} : s = 491;
	{8'd241,8'd251} : s = 492;
	{8'd241,8'd252} : s = 493;
	{8'd241,8'd253} : s = 494;
	{8'd241,8'd254} : s = 495;
	{8'd241,8'd255} : s = 496;
	{8'd242,8'd0} : s = 242;
	{8'd242,8'd1} : s = 243;
	{8'd242,8'd2} : s = 244;
	{8'd242,8'd3} : s = 245;
	{8'd242,8'd4} : s = 246;
	{8'd242,8'd5} : s = 247;
	{8'd242,8'd6} : s = 248;
	{8'd242,8'd7} : s = 249;
	{8'd242,8'd8} : s = 250;
	{8'd242,8'd9} : s = 251;
	{8'd242,8'd10} : s = 252;
	{8'd242,8'd11} : s = 253;
	{8'd242,8'd12} : s = 254;
	{8'd242,8'd13} : s = 255;
	{8'd242,8'd14} : s = 256;
	{8'd242,8'd15} : s = 257;
	{8'd242,8'd16} : s = 258;
	{8'd242,8'd17} : s = 259;
	{8'd242,8'd18} : s = 260;
	{8'd242,8'd19} : s = 261;
	{8'd242,8'd20} : s = 262;
	{8'd242,8'd21} : s = 263;
	{8'd242,8'd22} : s = 264;
	{8'd242,8'd23} : s = 265;
	{8'd242,8'd24} : s = 266;
	{8'd242,8'd25} : s = 267;
	{8'd242,8'd26} : s = 268;
	{8'd242,8'd27} : s = 269;
	{8'd242,8'd28} : s = 270;
	{8'd242,8'd29} : s = 271;
	{8'd242,8'd30} : s = 272;
	{8'd242,8'd31} : s = 273;
	{8'd242,8'd32} : s = 274;
	{8'd242,8'd33} : s = 275;
	{8'd242,8'd34} : s = 276;
	{8'd242,8'd35} : s = 277;
	{8'd242,8'd36} : s = 278;
	{8'd242,8'd37} : s = 279;
	{8'd242,8'd38} : s = 280;
	{8'd242,8'd39} : s = 281;
	{8'd242,8'd40} : s = 282;
	{8'd242,8'd41} : s = 283;
	{8'd242,8'd42} : s = 284;
	{8'd242,8'd43} : s = 285;
	{8'd242,8'd44} : s = 286;
	{8'd242,8'd45} : s = 287;
	{8'd242,8'd46} : s = 288;
	{8'd242,8'd47} : s = 289;
	{8'd242,8'd48} : s = 290;
	{8'd242,8'd49} : s = 291;
	{8'd242,8'd50} : s = 292;
	{8'd242,8'd51} : s = 293;
	{8'd242,8'd52} : s = 294;
	{8'd242,8'd53} : s = 295;
	{8'd242,8'd54} : s = 296;
	{8'd242,8'd55} : s = 297;
	{8'd242,8'd56} : s = 298;
	{8'd242,8'd57} : s = 299;
	{8'd242,8'd58} : s = 300;
	{8'd242,8'd59} : s = 301;
	{8'd242,8'd60} : s = 302;
	{8'd242,8'd61} : s = 303;
	{8'd242,8'd62} : s = 304;
	{8'd242,8'd63} : s = 305;
	{8'd242,8'd64} : s = 306;
	{8'd242,8'd65} : s = 307;
	{8'd242,8'd66} : s = 308;
	{8'd242,8'd67} : s = 309;
	{8'd242,8'd68} : s = 310;
	{8'd242,8'd69} : s = 311;
	{8'd242,8'd70} : s = 312;
	{8'd242,8'd71} : s = 313;
	{8'd242,8'd72} : s = 314;
	{8'd242,8'd73} : s = 315;
	{8'd242,8'd74} : s = 316;
	{8'd242,8'd75} : s = 317;
	{8'd242,8'd76} : s = 318;
	{8'd242,8'd77} : s = 319;
	{8'd242,8'd78} : s = 320;
	{8'd242,8'd79} : s = 321;
	{8'd242,8'd80} : s = 322;
	{8'd242,8'd81} : s = 323;
	{8'd242,8'd82} : s = 324;
	{8'd242,8'd83} : s = 325;
	{8'd242,8'd84} : s = 326;
	{8'd242,8'd85} : s = 327;
	{8'd242,8'd86} : s = 328;
	{8'd242,8'd87} : s = 329;
	{8'd242,8'd88} : s = 330;
	{8'd242,8'd89} : s = 331;
	{8'd242,8'd90} : s = 332;
	{8'd242,8'd91} : s = 333;
	{8'd242,8'd92} : s = 334;
	{8'd242,8'd93} : s = 335;
	{8'd242,8'd94} : s = 336;
	{8'd242,8'd95} : s = 337;
	{8'd242,8'd96} : s = 338;
	{8'd242,8'd97} : s = 339;
	{8'd242,8'd98} : s = 340;
	{8'd242,8'd99} : s = 341;
	{8'd242,8'd100} : s = 342;
	{8'd242,8'd101} : s = 343;
	{8'd242,8'd102} : s = 344;
	{8'd242,8'd103} : s = 345;
	{8'd242,8'd104} : s = 346;
	{8'd242,8'd105} : s = 347;
	{8'd242,8'd106} : s = 348;
	{8'd242,8'd107} : s = 349;
	{8'd242,8'd108} : s = 350;
	{8'd242,8'd109} : s = 351;
	{8'd242,8'd110} : s = 352;
	{8'd242,8'd111} : s = 353;
	{8'd242,8'd112} : s = 354;
	{8'd242,8'd113} : s = 355;
	{8'd242,8'd114} : s = 356;
	{8'd242,8'd115} : s = 357;
	{8'd242,8'd116} : s = 358;
	{8'd242,8'd117} : s = 359;
	{8'd242,8'd118} : s = 360;
	{8'd242,8'd119} : s = 361;
	{8'd242,8'd120} : s = 362;
	{8'd242,8'd121} : s = 363;
	{8'd242,8'd122} : s = 364;
	{8'd242,8'd123} : s = 365;
	{8'd242,8'd124} : s = 366;
	{8'd242,8'd125} : s = 367;
	{8'd242,8'd126} : s = 368;
	{8'd242,8'd127} : s = 369;
	{8'd242,8'd128} : s = 370;
	{8'd242,8'd129} : s = 371;
	{8'd242,8'd130} : s = 372;
	{8'd242,8'd131} : s = 373;
	{8'd242,8'd132} : s = 374;
	{8'd242,8'd133} : s = 375;
	{8'd242,8'd134} : s = 376;
	{8'd242,8'd135} : s = 377;
	{8'd242,8'd136} : s = 378;
	{8'd242,8'd137} : s = 379;
	{8'd242,8'd138} : s = 380;
	{8'd242,8'd139} : s = 381;
	{8'd242,8'd140} : s = 382;
	{8'd242,8'd141} : s = 383;
	{8'd242,8'd142} : s = 384;
	{8'd242,8'd143} : s = 385;
	{8'd242,8'd144} : s = 386;
	{8'd242,8'd145} : s = 387;
	{8'd242,8'd146} : s = 388;
	{8'd242,8'd147} : s = 389;
	{8'd242,8'd148} : s = 390;
	{8'd242,8'd149} : s = 391;
	{8'd242,8'd150} : s = 392;
	{8'd242,8'd151} : s = 393;
	{8'd242,8'd152} : s = 394;
	{8'd242,8'd153} : s = 395;
	{8'd242,8'd154} : s = 396;
	{8'd242,8'd155} : s = 397;
	{8'd242,8'd156} : s = 398;
	{8'd242,8'd157} : s = 399;
	{8'd242,8'd158} : s = 400;
	{8'd242,8'd159} : s = 401;
	{8'd242,8'd160} : s = 402;
	{8'd242,8'd161} : s = 403;
	{8'd242,8'd162} : s = 404;
	{8'd242,8'd163} : s = 405;
	{8'd242,8'd164} : s = 406;
	{8'd242,8'd165} : s = 407;
	{8'd242,8'd166} : s = 408;
	{8'd242,8'd167} : s = 409;
	{8'd242,8'd168} : s = 410;
	{8'd242,8'd169} : s = 411;
	{8'd242,8'd170} : s = 412;
	{8'd242,8'd171} : s = 413;
	{8'd242,8'd172} : s = 414;
	{8'd242,8'd173} : s = 415;
	{8'd242,8'd174} : s = 416;
	{8'd242,8'd175} : s = 417;
	{8'd242,8'd176} : s = 418;
	{8'd242,8'd177} : s = 419;
	{8'd242,8'd178} : s = 420;
	{8'd242,8'd179} : s = 421;
	{8'd242,8'd180} : s = 422;
	{8'd242,8'd181} : s = 423;
	{8'd242,8'd182} : s = 424;
	{8'd242,8'd183} : s = 425;
	{8'd242,8'd184} : s = 426;
	{8'd242,8'd185} : s = 427;
	{8'd242,8'd186} : s = 428;
	{8'd242,8'd187} : s = 429;
	{8'd242,8'd188} : s = 430;
	{8'd242,8'd189} : s = 431;
	{8'd242,8'd190} : s = 432;
	{8'd242,8'd191} : s = 433;
	{8'd242,8'd192} : s = 434;
	{8'd242,8'd193} : s = 435;
	{8'd242,8'd194} : s = 436;
	{8'd242,8'd195} : s = 437;
	{8'd242,8'd196} : s = 438;
	{8'd242,8'd197} : s = 439;
	{8'd242,8'd198} : s = 440;
	{8'd242,8'd199} : s = 441;
	{8'd242,8'd200} : s = 442;
	{8'd242,8'd201} : s = 443;
	{8'd242,8'd202} : s = 444;
	{8'd242,8'd203} : s = 445;
	{8'd242,8'd204} : s = 446;
	{8'd242,8'd205} : s = 447;
	{8'd242,8'd206} : s = 448;
	{8'd242,8'd207} : s = 449;
	{8'd242,8'd208} : s = 450;
	{8'd242,8'd209} : s = 451;
	{8'd242,8'd210} : s = 452;
	{8'd242,8'd211} : s = 453;
	{8'd242,8'd212} : s = 454;
	{8'd242,8'd213} : s = 455;
	{8'd242,8'd214} : s = 456;
	{8'd242,8'd215} : s = 457;
	{8'd242,8'd216} : s = 458;
	{8'd242,8'd217} : s = 459;
	{8'd242,8'd218} : s = 460;
	{8'd242,8'd219} : s = 461;
	{8'd242,8'd220} : s = 462;
	{8'd242,8'd221} : s = 463;
	{8'd242,8'd222} : s = 464;
	{8'd242,8'd223} : s = 465;
	{8'd242,8'd224} : s = 466;
	{8'd242,8'd225} : s = 467;
	{8'd242,8'd226} : s = 468;
	{8'd242,8'd227} : s = 469;
	{8'd242,8'd228} : s = 470;
	{8'd242,8'd229} : s = 471;
	{8'd242,8'd230} : s = 472;
	{8'd242,8'd231} : s = 473;
	{8'd242,8'd232} : s = 474;
	{8'd242,8'd233} : s = 475;
	{8'd242,8'd234} : s = 476;
	{8'd242,8'd235} : s = 477;
	{8'd242,8'd236} : s = 478;
	{8'd242,8'd237} : s = 479;
	{8'd242,8'd238} : s = 480;
	{8'd242,8'd239} : s = 481;
	{8'd242,8'd240} : s = 482;
	{8'd242,8'd241} : s = 483;
	{8'd242,8'd242} : s = 484;
	{8'd242,8'd243} : s = 485;
	{8'd242,8'd244} : s = 486;
	{8'd242,8'd245} : s = 487;
	{8'd242,8'd246} : s = 488;
	{8'd242,8'd247} : s = 489;
	{8'd242,8'd248} : s = 490;
	{8'd242,8'd249} : s = 491;
	{8'd242,8'd250} : s = 492;
	{8'd242,8'd251} : s = 493;
	{8'd242,8'd252} : s = 494;
	{8'd242,8'd253} : s = 495;
	{8'd242,8'd254} : s = 496;
	{8'd242,8'd255} : s = 497;
	{8'd243,8'd0} : s = 243;
	{8'd243,8'd1} : s = 244;
	{8'd243,8'd2} : s = 245;
	{8'd243,8'd3} : s = 246;
	{8'd243,8'd4} : s = 247;
	{8'd243,8'd5} : s = 248;
	{8'd243,8'd6} : s = 249;
	{8'd243,8'd7} : s = 250;
	{8'd243,8'd8} : s = 251;
	{8'd243,8'd9} : s = 252;
	{8'd243,8'd10} : s = 253;
	{8'd243,8'd11} : s = 254;
	{8'd243,8'd12} : s = 255;
	{8'd243,8'd13} : s = 256;
	{8'd243,8'd14} : s = 257;
	{8'd243,8'd15} : s = 258;
	{8'd243,8'd16} : s = 259;
	{8'd243,8'd17} : s = 260;
	{8'd243,8'd18} : s = 261;
	{8'd243,8'd19} : s = 262;
	{8'd243,8'd20} : s = 263;
	{8'd243,8'd21} : s = 264;
	{8'd243,8'd22} : s = 265;
	{8'd243,8'd23} : s = 266;
	{8'd243,8'd24} : s = 267;
	{8'd243,8'd25} : s = 268;
	{8'd243,8'd26} : s = 269;
	{8'd243,8'd27} : s = 270;
	{8'd243,8'd28} : s = 271;
	{8'd243,8'd29} : s = 272;
	{8'd243,8'd30} : s = 273;
	{8'd243,8'd31} : s = 274;
	{8'd243,8'd32} : s = 275;
	{8'd243,8'd33} : s = 276;
	{8'd243,8'd34} : s = 277;
	{8'd243,8'd35} : s = 278;
	{8'd243,8'd36} : s = 279;
	{8'd243,8'd37} : s = 280;
	{8'd243,8'd38} : s = 281;
	{8'd243,8'd39} : s = 282;
	{8'd243,8'd40} : s = 283;
	{8'd243,8'd41} : s = 284;
	{8'd243,8'd42} : s = 285;
	{8'd243,8'd43} : s = 286;
	{8'd243,8'd44} : s = 287;
	{8'd243,8'd45} : s = 288;
	{8'd243,8'd46} : s = 289;
	{8'd243,8'd47} : s = 290;
	{8'd243,8'd48} : s = 291;
	{8'd243,8'd49} : s = 292;
	{8'd243,8'd50} : s = 293;
	{8'd243,8'd51} : s = 294;
	{8'd243,8'd52} : s = 295;
	{8'd243,8'd53} : s = 296;
	{8'd243,8'd54} : s = 297;
	{8'd243,8'd55} : s = 298;
	{8'd243,8'd56} : s = 299;
	{8'd243,8'd57} : s = 300;
	{8'd243,8'd58} : s = 301;
	{8'd243,8'd59} : s = 302;
	{8'd243,8'd60} : s = 303;
	{8'd243,8'd61} : s = 304;
	{8'd243,8'd62} : s = 305;
	{8'd243,8'd63} : s = 306;
	{8'd243,8'd64} : s = 307;
	{8'd243,8'd65} : s = 308;
	{8'd243,8'd66} : s = 309;
	{8'd243,8'd67} : s = 310;
	{8'd243,8'd68} : s = 311;
	{8'd243,8'd69} : s = 312;
	{8'd243,8'd70} : s = 313;
	{8'd243,8'd71} : s = 314;
	{8'd243,8'd72} : s = 315;
	{8'd243,8'd73} : s = 316;
	{8'd243,8'd74} : s = 317;
	{8'd243,8'd75} : s = 318;
	{8'd243,8'd76} : s = 319;
	{8'd243,8'd77} : s = 320;
	{8'd243,8'd78} : s = 321;
	{8'd243,8'd79} : s = 322;
	{8'd243,8'd80} : s = 323;
	{8'd243,8'd81} : s = 324;
	{8'd243,8'd82} : s = 325;
	{8'd243,8'd83} : s = 326;
	{8'd243,8'd84} : s = 327;
	{8'd243,8'd85} : s = 328;
	{8'd243,8'd86} : s = 329;
	{8'd243,8'd87} : s = 330;
	{8'd243,8'd88} : s = 331;
	{8'd243,8'd89} : s = 332;
	{8'd243,8'd90} : s = 333;
	{8'd243,8'd91} : s = 334;
	{8'd243,8'd92} : s = 335;
	{8'd243,8'd93} : s = 336;
	{8'd243,8'd94} : s = 337;
	{8'd243,8'd95} : s = 338;
	{8'd243,8'd96} : s = 339;
	{8'd243,8'd97} : s = 340;
	{8'd243,8'd98} : s = 341;
	{8'd243,8'd99} : s = 342;
	{8'd243,8'd100} : s = 343;
	{8'd243,8'd101} : s = 344;
	{8'd243,8'd102} : s = 345;
	{8'd243,8'd103} : s = 346;
	{8'd243,8'd104} : s = 347;
	{8'd243,8'd105} : s = 348;
	{8'd243,8'd106} : s = 349;
	{8'd243,8'd107} : s = 350;
	{8'd243,8'd108} : s = 351;
	{8'd243,8'd109} : s = 352;
	{8'd243,8'd110} : s = 353;
	{8'd243,8'd111} : s = 354;
	{8'd243,8'd112} : s = 355;
	{8'd243,8'd113} : s = 356;
	{8'd243,8'd114} : s = 357;
	{8'd243,8'd115} : s = 358;
	{8'd243,8'd116} : s = 359;
	{8'd243,8'd117} : s = 360;
	{8'd243,8'd118} : s = 361;
	{8'd243,8'd119} : s = 362;
	{8'd243,8'd120} : s = 363;
	{8'd243,8'd121} : s = 364;
	{8'd243,8'd122} : s = 365;
	{8'd243,8'd123} : s = 366;
	{8'd243,8'd124} : s = 367;
	{8'd243,8'd125} : s = 368;
	{8'd243,8'd126} : s = 369;
	{8'd243,8'd127} : s = 370;
	{8'd243,8'd128} : s = 371;
	{8'd243,8'd129} : s = 372;
	{8'd243,8'd130} : s = 373;
	{8'd243,8'd131} : s = 374;
	{8'd243,8'd132} : s = 375;
	{8'd243,8'd133} : s = 376;
	{8'd243,8'd134} : s = 377;
	{8'd243,8'd135} : s = 378;
	{8'd243,8'd136} : s = 379;
	{8'd243,8'd137} : s = 380;
	{8'd243,8'd138} : s = 381;
	{8'd243,8'd139} : s = 382;
	{8'd243,8'd140} : s = 383;
	{8'd243,8'd141} : s = 384;
	{8'd243,8'd142} : s = 385;
	{8'd243,8'd143} : s = 386;
	{8'd243,8'd144} : s = 387;
	{8'd243,8'd145} : s = 388;
	{8'd243,8'd146} : s = 389;
	{8'd243,8'd147} : s = 390;
	{8'd243,8'd148} : s = 391;
	{8'd243,8'd149} : s = 392;
	{8'd243,8'd150} : s = 393;
	{8'd243,8'd151} : s = 394;
	{8'd243,8'd152} : s = 395;
	{8'd243,8'd153} : s = 396;
	{8'd243,8'd154} : s = 397;
	{8'd243,8'd155} : s = 398;
	{8'd243,8'd156} : s = 399;
	{8'd243,8'd157} : s = 400;
	{8'd243,8'd158} : s = 401;
	{8'd243,8'd159} : s = 402;
	{8'd243,8'd160} : s = 403;
	{8'd243,8'd161} : s = 404;
	{8'd243,8'd162} : s = 405;
	{8'd243,8'd163} : s = 406;
	{8'd243,8'd164} : s = 407;
	{8'd243,8'd165} : s = 408;
	{8'd243,8'd166} : s = 409;
	{8'd243,8'd167} : s = 410;
	{8'd243,8'd168} : s = 411;
	{8'd243,8'd169} : s = 412;
	{8'd243,8'd170} : s = 413;
	{8'd243,8'd171} : s = 414;
	{8'd243,8'd172} : s = 415;
	{8'd243,8'd173} : s = 416;
	{8'd243,8'd174} : s = 417;
	{8'd243,8'd175} : s = 418;
	{8'd243,8'd176} : s = 419;
	{8'd243,8'd177} : s = 420;
	{8'd243,8'd178} : s = 421;
	{8'd243,8'd179} : s = 422;
	{8'd243,8'd180} : s = 423;
	{8'd243,8'd181} : s = 424;
	{8'd243,8'd182} : s = 425;
	{8'd243,8'd183} : s = 426;
	{8'd243,8'd184} : s = 427;
	{8'd243,8'd185} : s = 428;
	{8'd243,8'd186} : s = 429;
	{8'd243,8'd187} : s = 430;
	{8'd243,8'd188} : s = 431;
	{8'd243,8'd189} : s = 432;
	{8'd243,8'd190} : s = 433;
	{8'd243,8'd191} : s = 434;
	{8'd243,8'd192} : s = 435;
	{8'd243,8'd193} : s = 436;
	{8'd243,8'd194} : s = 437;
	{8'd243,8'd195} : s = 438;
	{8'd243,8'd196} : s = 439;
	{8'd243,8'd197} : s = 440;
	{8'd243,8'd198} : s = 441;
	{8'd243,8'd199} : s = 442;
	{8'd243,8'd200} : s = 443;
	{8'd243,8'd201} : s = 444;
	{8'd243,8'd202} : s = 445;
	{8'd243,8'd203} : s = 446;
	{8'd243,8'd204} : s = 447;
	{8'd243,8'd205} : s = 448;
	{8'd243,8'd206} : s = 449;
	{8'd243,8'd207} : s = 450;
	{8'd243,8'd208} : s = 451;
	{8'd243,8'd209} : s = 452;
	{8'd243,8'd210} : s = 453;
	{8'd243,8'd211} : s = 454;
	{8'd243,8'd212} : s = 455;
	{8'd243,8'd213} : s = 456;
	{8'd243,8'd214} : s = 457;
	{8'd243,8'd215} : s = 458;
	{8'd243,8'd216} : s = 459;
	{8'd243,8'd217} : s = 460;
	{8'd243,8'd218} : s = 461;
	{8'd243,8'd219} : s = 462;
	{8'd243,8'd220} : s = 463;
	{8'd243,8'd221} : s = 464;
	{8'd243,8'd222} : s = 465;
	{8'd243,8'd223} : s = 466;
	{8'd243,8'd224} : s = 467;
	{8'd243,8'd225} : s = 468;
	{8'd243,8'd226} : s = 469;
	{8'd243,8'd227} : s = 470;
	{8'd243,8'd228} : s = 471;
	{8'd243,8'd229} : s = 472;
	{8'd243,8'd230} : s = 473;
	{8'd243,8'd231} : s = 474;
	{8'd243,8'd232} : s = 475;
	{8'd243,8'd233} : s = 476;
	{8'd243,8'd234} : s = 477;
	{8'd243,8'd235} : s = 478;
	{8'd243,8'd236} : s = 479;
	{8'd243,8'd237} : s = 480;
	{8'd243,8'd238} : s = 481;
	{8'd243,8'd239} : s = 482;
	{8'd243,8'd240} : s = 483;
	{8'd243,8'd241} : s = 484;
	{8'd243,8'd242} : s = 485;
	{8'd243,8'd243} : s = 486;
	{8'd243,8'd244} : s = 487;
	{8'd243,8'd245} : s = 488;
	{8'd243,8'd246} : s = 489;
	{8'd243,8'd247} : s = 490;
	{8'd243,8'd248} : s = 491;
	{8'd243,8'd249} : s = 492;
	{8'd243,8'd250} : s = 493;
	{8'd243,8'd251} : s = 494;
	{8'd243,8'd252} : s = 495;
	{8'd243,8'd253} : s = 496;
	{8'd243,8'd254} : s = 497;
	{8'd243,8'd255} : s = 498;
	{8'd244,8'd0} : s = 244;
	{8'd244,8'd1} : s = 245;
	{8'd244,8'd2} : s = 246;
	{8'd244,8'd3} : s = 247;
	{8'd244,8'd4} : s = 248;
	{8'd244,8'd5} : s = 249;
	{8'd244,8'd6} : s = 250;
	{8'd244,8'd7} : s = 251;
	{8'd244,8'd8} : s = 252;
	{8'd244,8'd9} : s = 253;
	{8'd244,8'd10} : s = 254;
	{8'd244,8'd11} : s = 255;
	{8'd244,8'd12} : s = 256;
	{8'd244,8'd13} : s = 257;
	{8'd244,8'd14} : s = 258;
	{8'd244,8'd15} : s = 259;
	{8'd244,8'd16} : s = 260;
	{8'd244,8'd17} : s = 261;
	{8'd244,8'd18} : s = 262;
	{8'd244,8'd19} : s = 263;
	{8'd244,8'd20} : s = 264;
	{8'd244,8'd21} : s = 265;
	{8'd244,8'd22} : s = 266;
	{8'd244,8'd23} : s = 267;
	{8'd244,8'd24} : s = 268;
	{8'd244,8'd25} : s = 269;
	{8'd244,8'd26} : s = 270;
	{8'd244,8'd27} : s = 271;
	{8'd244,8'd28} : s = 272;
	{8'd244,8'd29} : s = 273;
	{8'd244,8'd30} : s = 274;
	{8'd244,8'd31} : s = 275;
	{8'd244,8'd32} : s = 276;
	{8'd244,8'd33} : s = 277;
	{8'd244,8'd34} : s = 278;
	{8'd244,8'd35} : s = 279;
	{8'd244,8'd36} : s = 280;
	{8'd244,8'd37} : s = 281;
	{8'd244,8'd38} : s = 282;
	{8'd244,8'd39} : s = 283;
	{8'd244,8'd40} : s = 284;
	{8'd244,8'd41} : s = 285;
	{8'd244,8'd42} : s = 286;
	{8'd244,8'd43} : s = 287;
	{8'd244,8'd44} : s = 288;
	{8'd244,8'd45} : s = 289;
	{8'd244,8'd46} : s = 290;
	{8'd244,8'd47} : s = 291;
	{8'd244,8'd48} : s = 292;
	{8'd244,8'd49} : s = 293;
	{8'd244,8'd50} : s = 294;
	{8'd244,8'd51} : s = 295;
	{8'd244,8'd52} : s = 296;
	{8'd244,8'd53} : s = 297;
	{8'd244,8'd54} : s = 298;
	{8'd244,8'd55} : s = 299;
	{8'd244,8'd56} : s = 300;
	{8'd244,8'd57} : s = 301;
	{8'd244,8'd58} : s = 302;
	{8'd244,8'd59} : s = 303;
	{8'd244,8'd60} : s = 304;
	{8'd244,8'd61} : s = 305;
	{8'd244,8'd62} : s = 306;
	{8'd244,8'd63} : s = 307;
	{8'd244,8'd64} : s = 308;
	{8'd244,8'd65} : s = 309;
	{8'd244,8'd66} : s = 310;
	{8'd244,8'd67} : s = 311;
	{8'd244,8'd68} : s = 312;
	{8'd244,8'd69} : s = 313;
	{8'd244,8'd70} : s = 314;
	{8'd244,8'd71} : s = 315;
	{8'd244,8'd72} : s = 316;
	{8'd244,8'd73} : s = 317;
	{8'd244,8'd74} : s = 318;
	{8'd244,8'd75} : s = 319;
	{8'd244,8'd76} : s = 320;
	{8'd244,8'd77} : s = 321;
	{8'd244,8'd78} : s = 322;
	{8'd244,8'd79} : s = 323;
	{8'd244,8'd80} : s = 324;
	{8'd244,8'd81} : s = 325;
	{8'd244,8'd82} : s = 326;
	{8'd244,8'd83} : s = 327;
	{8'd244,8'd84} : s = 328;
	{8'd244,8'd85} : s = 329;
	{8'd244,8'd86} : s = 330;
	{8'd244,8'd87} : s = 331;
	{8'd244,8'd88} : s = 332;
	{8'd244,8'd89} : s = 333;
	{8'd244,8'd90} : s = 334;
	{8'd244,8'd91} : s = 335;
	{8'd244,8'd92} : s = 336;
	{8'd244,8'd93} : s = 337;
	{8'd244,8'd94} : s = 338;
	{8'd244,8'd95} : s = 339;
	{8'd244,8'd96} : s = 340;
	{8'd244,8'd97} : s = 341;
	{8'd244,8'd98} : s = 342;
	{8'd244,8'd99} : s = 343;
	{8'd244,8'd100} : s = 344;
	{8'd244,8'd101} : s = 345;
	{8'd244,8'd102} : s = 346;
	{8'd244,8'd103} : s = 347;
	{8'd244,8'd104} : s = 348;
	{8'd244,8'd105} : s = 349;
	{8'd244,8'd106} : s = 350;
	{8'd244,8'd107} : s = 351;
	{8'd244,8'd108} : s = 352;
	{8'd244,8'd109} : s = 353;
	{8'd244,8'd110} : s = 354;
	{8'd244,8'd111} : s = 355;
	{8'd244,8'd112} : s = 356;
	{8'd244,8'd113} : s = 357;
	{8'd244,8'd114} : s = 358;
	{8'd244,8'd115} : s = 359;
	{8'd244,8'd116} : s = 360;
	{8'd244,8'd117} : s = 361;
	{8'd244,8'd118} : s = 362;
	{8'd244,8'd119} : s = 363;
	{8'd244,8'd120} : s = 364;
	{8'd244,8'd121} : s = 365;
	{8'd244,8'd122} : s = 366;
	{8'd244,8'd123} : s = 367;
	{8'd244,8'd124} : s = 368;
	{8'd244,8'd125} : s = 369;
	{8'd244,8'd126} : s = 370;
	{8'd244,8'd127} : s = 371;
	{8'd244,8'd128} : s = 372;
	{8'd244,8'd129} : s = 373;
	{8'd244,8'd130} : s = 374;
	{8'd244,8'd131} : s = 375;
	{8'd244,8'd132} : s = 376;
	{8'd244,8'd133} : s = 377;
	{8'd244,8'd134} : s = 378;
	{8'd244,8'd135} : s = 379;
	{8'd244,8'd136} : s = 380;
	{8'd244,8'd137} : s = 381;
	{8'd244,8'd138} : s = 382;
	{8'd244,8'd139} : s = 383;
	{8'd244,8'd140} : s = 384;
	{8'd244,8'd141} : s = 385;
	{8'd244,8'd142} : s = 386;
	{8'd244,8'd143} : s = 387;
	{8'd244,8'd144} : s = 388;
	{8'd244,8'd145} : s = 389;
	{8'd244,8'd146} : s = 390;
	{8'd244,8'd147} : s = 391;
	{8'd244,8'd148} : s = 392;
	{8'd244,8'd149} : s = 393;
	{8'd244,8'd150} : s = 394;
	{8'd244,8'd151} : s = 395;
	{8'd244,8'd152} : s = 396;
	{8'd244,8'd153} : s = 397;
	{8'd244,8'd154} : s = 398;
	{8'd244,8'd155} : s = 399;
	{8'd244,8'd156} : s = 400;
	{8'd244,8'd157} : s = 401;
	{8'd244,8'd158} : s = 402;
	{8'd244,8'd159} : s = 403;
	{8'd244,8'd160} : s = 404;
	{8'd244,8'd161} : s = 405;
	{8'd244,8'd162} : s = 406;
	{8'd244,8'd163} : s = 407;
	{8'd244,8'd164} : s = 408;
	{8'd244,8'd165} : s = 409;
	{8'd244,8'd166} : s = 410;
	{8'd244,8'd167} : s = 411;
	{8'd244,8'd168} : s = 412;
	{8'd244,8'd169} : s = 413;
	{8'd244,8'd170} : s = 414;
	{8'd244,8'd171} : s = 415;
	{8'd244,8'd172} : s = 416;
	{8'd244,8'd173} : s = 417;
	{8'd244,8'd174} : s = 418;
	{8'd244,8'd175} : s = 419;
	{8'd244,8'd176} : s = 420;
	{8'd244,8'd177} : s = 421;
	{8'd244,8'd178} : s = 422;
	{8'd244,8'd179} : s = 423;
	{8'd244,8'd180} : s = 424;
	{8'd244,8'd181} : s = 425;
	{8'd244,8'd182} : s = 426;
	{8'd244,8'd183} : s = 427;
	{8'd244,8'd184} : s = 428;
	{8'd244,8'd185} : s = 429;
	{8'd244,8'd186} : s = 430;
	{8'd244,8'd187} : s = 431;
	{8'd244,8'd188} : s = 432;
	{8'd244,8'd189} : s = 433;
	{8'd244,8'd190} : s = 434;
	{8'd244,8'd191} : s = 435;
	{8'd244,8'd192} : s = 436;
	{8'd244,8'd193} : s = 437;
	{8'd244,8'd194} : s = 438;
	{8'd244,8'd195} : s = 439;
	{8'd244,8'd196} : s = 440;
	{8'd244,8'd197} : s = 441;
	{8'd244,8'd198} : s = 442;
	{8'd244,8'd199} : s = 443;
	{8'd244,8'd200} : s = 444;
	{8'd244,8'd201} : s = 445;
	{8'd244,8'd202} : s = 446;
	{8'd244,8'd203} : s = 447;
	{8'd244,8'd204} : s = 448;
	{8'd244,8'd205} : s = 449;
	{8'd244,8'd206} : s = 450;
	{8'd244,8'd207} : s = 451;
	{8'd244,8'd208} : s = 452;
	{8'd244,8'd209} : s = 453;
	{8'd244,8'd210} : s = 454;
	{8'd244,8'd211} : s = 455;
	{8'd244,8'd212} : s = 456;
	{8'd244,8'd213} : s = 457;
	{8'd244,8'd214} : s = 458;
	{8'd244,8'd215} : s = 459;
	{8'd244,8'd216} : s = 460;
	{8'd244,8'd217} : s = 461;
	{8'd244,8'd218} : s = 462;
	{8'd244,8'd219} : s = 463;
	{8'd244,8'd220} : s = 464;
	{8'd244,8'd221} : s = 465;
	{8'd244,8'd222} : s = 466;
	{8'd244,8'd223} : s = 467;
	{8'd244,8'd224} : s = 468;
	{8'd244,8'd225} : s = 469;
	{8'd244,8'd226} : s = 470;
	{8'd244,8'd227} : s = 471;
	{8'd244,8'd228} : s = 472;
	{8'd244,8'd229} : s = 473;
	{8'd244,8'd230} : s = 474;
	{8'd244,8'd231} : s = 475;
	{8'd244,8'd232} : s = 476;
	{8'd244,8'd233} : s = 477;
	{8'd244,8'd234} : s = 478;
	{8'd244,8'd235} : s = 479;
	{8'd244,8'd236} : s = 480;
	{8'd244,8'd237} : s = 481;
	{8'd244,8'd238} : s = 482;
	{8'd244,8'd239} : s = 483;
	{8'd244,8'd240} : s = 484;
	{8'd244,8'd241} : s = 485;
	{8'd244,8'd242} : s = 486;
	{8'd244,8'd243} : s = 487;
	{8'd244,8'd244} : s = 488;
	{8'd244,8'd245} : s = 489;
	{8'd244,8'd246} : s = 490;
	{8'd244,8'd247} : s = 491;
	{8'd244,8'd248} : s = 492;
	{8'd244,8'd249} : s = 493;
	{8'd244,8'd250} : s = 494;
	{8'd244,8'd251} : s = 495;
	{8'd244,8'd252} : s = 496;
	{8'd244,8'd253} : s = 497;
	{8'd244,8'd254} : s = 498;
	{8'd244,8'd255} : s = 499;
	{8'd245,8'd0} : s = 245;
	{8'd245,8'd1} : s = 246;
	{8'd245,8'd2} : s = 247;
	{8'd245,8'd3} : s = 248;
	{8'd245,8'd4} : s = 249;
	{8'd245,8'd5} : s = 250;
	{8'd245,8'd6} : s = 251;
	{8'd245,8'd7} : s = 252;
	{8'd245,8'd8} : s = 253;
	{8'd245,8'd9} : s = 254;
	{8'd245,8'd10} : s = 255;
	{8'd245,8'd11} : s = 256;
	{8'd245,8'd12} : s = 257;
	{8'd245,8'd13} : s = 258;
	{8'd245,8'd14} : s = 259;
	{8'd245,8'd15} : s = 260;
	{8'd245,8'd16} : s = 261;
	{8'd245,8'd17} : s = 262;
	{8'd245,8'd18} : s = 263;
	{8'd245,8'd19} : s = 264;
	{8'd245,8'd20} : s = 265;
	{8'd245,8'd21} : s = 266;
	{8'd245,8'd22} : s = 267;
	{8'd245,8'd23} : s = 268;
	{8'd245,8'd24} : s = 269;
	{8'd245,8'd25} : s = 270;
	{8'd245,8'd26} : s = 271;
	{8'd245,8'd27} : s = 272;
	{8'd245,8'd28} : s = 273;
	{8'd245,8'd29} : s = 274;
	{8'd245,8'd30} : s = 275;
	{8'd245,8'd31} : s = 276;
	{8'd245,8'd32} : s = 277;
	{8'd245,8'd33} : s = 278;
	{8'd245,8'd34} : s = 279;
	{8'd245,8'd35} : s = 280;
	{8'd245,8'd36} : s = 281;
	{8'd245,8'd37} : s = 282;
	{8'd245,8'd38} : s = 283;
	{8'd245,8'd39} : s = 284;
	{8'd245,8'd40} : s = 285;
	{8'd245,8'd41} : s = 286;
	{8'd245,8'd42} : s = 287;
	{8'd245,8'd43} : s = 288;
	{8'd245,8'd44} : s = 289;
	{8'd245,8'd45} : s = 290;
	{8'd245,8'd46} : s = 291;
	{8'd245,8'd47} : s = 292;
	{8'd245,8'd48} : s = 293;
	{8'd245,8'd49} : s = 294;
	{8'd245,8'd50} : s = 295;
	{8'd245,8'd51} : s = 296;
	{8'd245,8'd52} : s = 297;
	{8'd245,8'd53} : s = 298;
	{8'd245,8'd54} : s = 299;
	{8'd245,8'd55} : s = 300;
	{8'd245,8'd56} : s = 301;
	{8'd245,8'd57} : s = 302;
	{8'd245,8'd58} : s = 303;
	{8'd245,8'd59} : s = 304;
	{8'd245,8'd60} : s = 305;
	{8'd245,8'd61} : s = 306;
	{8'd245,8'd62} : s = 307;
	{8'd245,8'd63} : s = 308;
	{8'd245,8'd64} : s = 309;
	{8'd245,8'd65} : s = 310;
	{8'd245,8'd66} : s = 311;
	{8'd245,8'd67} : s = 312;
	{8'd245,8'd68} : s = 313;
	{8'd245,8'd69} : s = 314;
	{8'd245,8'd70} : s = 315;
	{8'd245,8'd71} : s = 316;
	{8'd245,8'd72} : s = 317;
	{8'd245,8'd73} : s = 318;
	{8'd245,8'd74} : s = 319;
	{8'd245,8'd75} : s = 320;
	{8'd245,8'd76} : s = 321;
	{8'd245,8'd77} : s = 322;
	{8'd245,8'd78} : s = 323;
	{8'd245,8'd79} : s = 324;
	{8'd245,8'd80} : s = 325;
	{8'd245,8'd81} : s = 326;
	{8'd245,8'd82} : s = 327;
	{8'd245,8'd83} : s = 328;
	{8'd245,8'd84} : s = 329;
	{8'd245,8'd85} : s = 330;
	{8'd245,8'd86} : s = 331;
	{8'd245,8'd87} : s = 332;
	{8'd245,8'd88} : s = 333;
	{8'd245,8'd89} : s = 334;
	{8'd245,8'd90} : s = 335;
	{8'd245,8'd91} : s = 336;
	{8'd245,8'd92} : s = 337;
	{8'd245,8'd93} : s = 338;
	{8'd245,8'd94} : s = 339;
	{8'd245,8'd95} : s = 340;
	{8'd245,8'd96} : s = 341;
	{8'd245,8'd97} : s = 342;
	{8'd245,8'd98} : s = 343;
	{8'd245,8'd99} : s = 344;
	{8'd245,8'd100} : s = 345;
	{8'd245,8'd101} : s = 346;
	{8'd245,8'd102} : s = 347;
	{8'd245,8'd103} : s = 348;
	{8'd245,8'd104} : s = 349;
	{8'd245,8'd105} : s = 350;
	{8'd245,8'd106} : s = 351;
	{8'd245,8'd107} : s = 352;
	{8'd245,8'd108} : s = 353;
	{8'd245,8'd109} : s = 354;
	{8'd245,8'd110} : s = 355;
	{8'd245,8'd111} : s = 356;
	{8'd245,8'd112} : s = 357;
	{8'd245,8'd113} : s = 358;
	{8'd245,8'd114} : s = 359;
	{8'd245,8'd115} : s = 360;
	{8'd245,8'd116} : s = 361;
	{8'd245,8'd117} : s = 362;
	{8'd245,8'd118} : s = 363;
	{8'd245,8'd119} : s = 364;
	{8'd245,8'd120} : s = 365;
	{8'd245,8'd121} : s = 366;
	{8'd245,8'd122} : s = 367;
	{8'd245,8'd123} : s = 368;
	{8'd245,8'd124} : s = 369;
	{8'd245,8'd125} : s = 370;
	{8'd245,8'd126} : s = 371;
	{8'd245,8'd127} : s = 372;
	{8'd245,8'd128} : s = 373;
	{8'd245,8'd129} : s = 374;
	{8'd245,8'd130} : s = 375;
	{8'd245,8'd131} : s = 376;
	{8'd245,8'd132} : s = 377;
	{8'd245,8'd133} : s = 378;
	{8'd245,8'd134} : s = 379;
	{8'd245,8'd135} : s = 380;
	{8'd245,8'd136} : s = 381;
	{8'd245,8'd137} : s = 382;
	{8'd245,8'd138} : s = 383;
	{8'd245,8'd139} : s = 384;
	{8'd245,8'd140} : s = 385;
	{8'd245,8'd141} : s = 386;
	{8'd245,8'd142} : s = 387;
	{8'd245,8'd143} : s = 388;
	{8'd245,8'd144} : s = 389;
	{8'd245,8'd145} : s = 390;
	{8'd245,8'd146} : s = 391;
	{8'd245,8'd147} : s = 392;
	{8'd245,8'd148} : s = 393;
	{8'd245,8'd149} : s = 394;
	{8'd245,8'd150} : s = 395;
	{8'd245,8'd151} : s = 396;
	{8'd245,8'd152} : s = 397;
	{8'd245,8'd153} : s = 398;
	{8'd245,8'd154} : s = 399;
	{8'd245,8'd155} : s = 400;
	{8'd245,8'd156} : s = 401;
	{8'd245,8'd157} : s = 402;
	{8'd245,8'd158} : s = 403;
	{8'd245,8'd159} : s = 404;
	{8'd245,8'd160} : s = 405;
	{8'd245,8'd161} : s = 406;
	{8'd245,8'd162} : s = 407;
	{8'd245,8'd163} : s = 408;
	{8'd245,8'd164} : s = 409;
	{8'd245,8'd165} : s = 410;
	{8'd245,8'd166} : s = 411;
	{8'd245,8'd167} : s = 412;
	{8'd245,8'd168} : s = 413;
	{8'd245,8'd169} : s = 414;
	{8'd245,8'd170} : s = 415;
	{8'd245,8'd171} : s = 416;
	{8'd245,8'd172} : s = 417;
	{8'd245,8'd173} : s = 418;
	{8'd245,8'd174} : s = 419;
	{8'd245,8'd175} : s = 420;
	{8'd245,8'd176} : s = 421;
	{8'd245,8'd177} : s = 422;
	{8'd245,8'd178} : s = 423;
	{8'd245,8'd179} : s = 424;
	{8'd245,8'd180} : s = 425;
	{8'd245,8'd181} : s = 426;
	{8'd245,8'd182} : s = 427;
	{8'd245,8'd183} : s = 428;
	{8'd245,8'd184} : s = 429;
	{8'd245,8'd185} : s = 430;
	{8'd245,8'd186} : s = 431;
	{8'd245,8'd187} : s = 432;
	{8'd245,8'd188} : s = 433;
	{8'd245,8'd189} : s = 434;
	{8'd245,8'd190} : s = 435;
	{8'd245,8'd191} : s = 436;
	{8'd245,8'd192} : s = 437;
	{8'd245,8'd193} : s = 438;
	{8'd245,8'd194} : s = 439;
	{8'd245,8'd195} : s = 440;
	{8'd245,8'd196} : s = 441;
	{8'd245,8'd197} : s = 442;
	{8'd245,8'd198} : s = 443;
	{8'd245,8'd199} : s = 444;
	{8'd245,8'd200} : s = 445;
	{8'd245,8'd201} : s = 446;
	{8'd245,8'd202} : s = 447;
	{8'd245,8'd203} : s = 448;
	{8'd245,8'd204} : s = 449;
	{8'd245,8'd205} : s = 450;
	{8'd245,8'd206} : s = 451;
	{8'd245,8'd207} : s = 452;
	{8'd245,8'd208} : s = 453;
	{8'd245,8'd209} : s = 454;
	{8'd245,8'd210} : s = 455;
	{8'd245,8'd211} : s = 456;
	{8'd245,8'd212} : s = 457;
	{8'd245,8'd213} : s = 458;
	{8'd245,8'd214} : s = 459;
	{8'd245,8'd215} : s = 460;
	{8'd245,8'd216} : s = 461;
	{8'd245,8'd217} : s = 462;
	{8'd245,8'd218} : s = 463;
	{8'd245,8'd219} : s = 464;
	{8'd245,8'd220} : s = 465;
	{8'd245,8'd221} : s = 466;
	{8'd245,8'd222} : s = 467;
	{8'd245,8'd223} : s = 468;
	{8'd245,8'd224} : s = 469;
	{8'd245,8'd225} : s = 470;
	{8'd245,8'd226} : s = 471;
	{8'd245,8'd227} : s = 472;
	{8'd245,8'd228} : s = 473;
	{8'd245,8'd229} : s = 474;
	{8'd245,8'd230} : s = 475;
	{8'd245,8'd231} : s = 476;
	{8'd245,8'd232} : s = 477;
	{8'd245,8'd233} : s = 478;
	{8'd245,8'd234} : s = 479;
	{8'd245,8'd235} : s = 480;
	{8'd245,8'd236} : s = 481;
	{8'd245,8'd237} : s = 482;
	{8'd245,8'd238} : s = 483;
	{8'd245,8'd239} : s = 484;
	{8'd245,8'd240} : s = 485;
	{8'd245,8'd241} : s = 486;
	{8'd245,8'd242} : s = 487;
	{8'd245,8'd243} : s = 488;
	{8'd245,8'd244} : s = 489;
	{8'd245,8'd245} : s = 490;
	{8'd245,8'd246} : s = 491;
	{8'd245,8'd247} : s = 492;
	{8'd245,8'd248} : s = 493;
	{8'd245,8'd249} : s = 494;
	{8'd245,8'd250} : s = 495;
	{8'd245,8'd251} : s = 496;
	{8'd245,8'd252} : s = 497;
	{8'd245,8'd253} : s = 498;
	{8'd245,8'd254} : s = 499;
	{8'd245,8'd255} : s = 500;
	{8'd246,8'd0} : s = 246;
	{8'd246,8'd1} : s = 247;
	{8'd246,8'd2} : s = 248;
	{8'd246,8'd3} : s = 249;
	{8'd246,8'd4} : s = 250;
	{8'd246,8'd5} : s = 251;
	{8'd246,8'd6} : s = 252;
	{8'd246,8'd7} : s = 253;
	{8'd246,8'd8} : s = 254;
	{8'd246,8'd9} : s = 255;
	{8'd246,8'd10} : s = 256;
	{8'd246,8'd11} : s = 257;
	{8'd246,8'd12} : s = 258;
	{8'd246,8'd13} : s = 259;
	{8'd246,8'd14} : s = 260;
	{8'd246,8'd15} : s = 261;
	{8'd246,8'd16} : s = 262;
	{8'd246,8'd17} : s = 263;
	{8'd246,8'd18} : s = 264;
	{8'd246,8'd19} : s = 265;
	{8'd246,8'd20} : s = 266;
	{8'd246,8'd21} : s = 267;
	{8'd246,8'd22} : s = 268;
	{8'd246,8'd23} : s = 269;
	{8'd246,8'd24} : s = 270;
	{8'd246,8'd25} : s = 271;
	{8'd246,8'd26} : s = 272;
	{8'd246,8'd27} : s = 273;
	{8'd246,8'd28} : s = 274;
	{8'd246,8'd29} : s = 275;
	{8'd246,8'd30} : s = 276;
	{8'd246,8'd31} : s = 277;
	{8'd246,8'd32} : s = 278;
	{8'd246,8'd33} : s = 279;
	{8'd246,8'd34} : s = 280;
	{8'd246,8'd35} : s = 281;
	{8'd246,8'd36} : s = 282;
	{8'd246,8'd37} : s = 283;
	{8'd246,8'd38} : s = 284;
	{8'd246,8'd39} : s = 285;
	{8'd246,8'd40} : s = 286;
	{8'd246,8'd41} : s = 287;
	{8'd246,8'd42} : s = 288;
	{8'd246,8'd43} : s = 289;
	{8'd246,8'd44} : s = 290;
	{8'd246,8'd45} : s = 291;
	{8'd246,8'd46} : s = 292;
	{8'd246,8'd47} : s = 293;
	{8'd246,8'd48} : s = 294;
	{8'd246,8'd49} : s = 295;
	{8'd246,8'd50} : s = 296;
	{8'd246,8'd51} : s = 297;
	{8'd246,8'd52} : s = 298;
	{8'd246,8'd53} : s = 299;
	{8'd246,8'd54} : s = 300;
	{8'd246,8'd55} : s = 301;
	{8'd246,8'd56} : s = 302;
	{8'd246,8'd57} : s = 303;
	{8'd246,8'd58} : s = 304;
	{8'd246,8'd59} : s = 305;
	{8'd246,8'd60} : s = 306;
	{8'd246,8'd61} : s = 307;
	{8'd246,8'd62} : s = 308;
	{8'd246,8'd63} : s = 309;
	{8'd246,8'd64} : s = 310;
	{8'd246,8'd65} : s = 311;
	{8'd246,8'd66} : s = 312;
	{8'd246,8'd67} : s = 313;
	{8'd246,8'd68} : s = 314;
	{8'd246,8'd69} : s = 315;
	{8'd246,8'd70} : s = 316;
	{8'd246,8'd71} : s = 317;
	{8'd246,8'd72} : s = 318;
	{8'd246,8'd73} : s = 319;
	{8'd246,8'd74} : s = 320;
	{8'd246,8'd75} : s = 321;
	{8'd246,8'd76} : s = 322;
	{8'd246,8'd77} : s = 323;
	{8'd246,8'd78} : s = 324;
	{8'd246,8'd79} : s = 325;
	{8'd246,8'd80} : s = 326;
	{8'd246,8'd81} : s = 327;
	{8'd246,8'd82} : s = 328;
	{8'd246,8'd83} : s = 329;
	{8'd246,8'd84} : s = 330;
	{8'd246,8'd85} : s = 331;
	{8'd246,8'd86} : s = 332;
	{8'd246,8'd87} : s = 333;
	{8'd246,8'd88} : s = 334;
	{8'd246,8'd89} : s = 335;
	{8'd246,8'd90} : s = 336;
	{8'd246,8'd91} : s = 337;
	{8'd246,8'd92} : s = 338;
	{8'd246,8'd93} : s = 339;
	{8'd246,8'd94} : s = 340;
	{8'd246,8'd95} : s = 341;
	{8'd246,8'd96} : s = 342;
	{8'd246,8'd97} : s = 343;
	{8'd246,8'd98} : s = 344;
	{8'd246,8'd99} : s = 345;
	{8'd246,8'd100} : s = 346;
	{8'd246,8'd101} : s = 347;
	{8'd246,8'd102} : s = 348;
	{8'd246,8'd103} : s = 349;
	{8'd246,8'd104} : s = 350;
	{8'd246,8'd105} : s = 351;
	{8'd246,8'd106} : s = 352;
	{8'd246,8'd107} : s = 353;
	{8'd246,8'd108} : s = 354;
	{8'd246,8'd109} : s = 355;
	{8'd246,8'd110} : s = 356;
	{8'd246,8'd111} : s = 357;
	{8'd246,8'd112} : s = 358;
	{8'd246,8'd113} : s = 359;
	{8'd246,8'd114} : s = 360;
	{8'd246,8'd115} : s = 361;
	{8'd246,8'd116} : s = 362;
	{8'd246,8'd117} : s = 363;
	{8'd246,8'd118} : s = 364;
	{8'd246,8'd119} : s = 365;
	{8'd246,8'd120} : s = 366;
	{8'd246,8'd121} : s = 367;
	{8'd246,8'd122} : s = 368;
	{8'd246,8'd123} : s = 369;
	{8'd246,8'd124} : s = 370;
	{8'd246,8'd125} : s = 371;
	{8'd246,8'd126} : s = 372;
	{8'd246,8'd127} : s = 373;
	{8'd246,8'd128} : s = 374;
	{8'd246,8'd129} : s = 375;
	{8'd246,8'd130} : s = 376;
	{8'd246,8'd131} : s = 377;
	{8'd246,8'd132} : s = 378;
	{8'd246,8'd133} : s = 379;
	{8'd246,8'd134} : s = 380;
	{8'd246,8'd135} : s = 381;
	{8'd246,8'd136} : s = 382;
	{8'd246,8'd137} : s = 383;
	{8'd246,8'd138} : s = 384;
	{8'd246,8'd139} : s = 385;
	{8'd246,8'd140} : s = 386;
	{8'd246,8'd141} : s = 387;
	{8'd246,8'd142} : s = 388;
	{8'd246,8'd143} : s = 389;
	{8'd246,8'd144} : s = 390;
	{8'd246,8'd145} : s = 391;
	{8'd246,8'd146} : s = 392;
	{8'd246,8'd147} : s = 393;
	{8'd246,8'd148} : s = 394;
	{8'd246,8'd149} : s = 395;
	{8'd246,8'd150} : s = 396;
	{8'd246,8'd151} : s = 397;
	{8'd246,8'd152} : s = 398;
	{8'd246,8'd153} : s = 399;
	{8'd246,8'd154} : s = 400;
	{8'd246,8'd155} : s = 401;
	{8'd246,8'd156} : s = 402;
	{8'd246,8'd157} : s = 403;
	{8'd246,8'd158} : s = 404;
	{8'd246,8'd159} : s = 405;
	{8'd246,8'd160} : s = 406;
	{8'd246,8'd161} : s = 407;
	{8'd246,8'd162} : s = 408;
	{8'd246,8'd163} : s = 409;
	{8'd246,8'd164} : s = 410;
	{8'd246,8'd165} : s = 411;
	{8'd246,8'd166} : s = 412;
	{8'd246,8'd167} : s = 413;
	{8'd246,8'd168} : s = 414;
	{8'd246,8'd169} : s = 415;
	{8'd246,8'd170} : s = 416;
	{8'd246,8'd171} : s = 417;
	{8'd246,8'd172} : s = 418;
	{8'd246,8'd173} : s = 419;
	{8'd246,8'd174} : s = 420;
	{8'd246,8'd175} : s = 421;
	{8'd246,8'd176} : s = 422;
	{8'd246,8'd177} : s = 423;
	{8'd246,8'd178} : s = 424;
	{8'd246,8'd179} : s = 425;
	{8'd246,8'd180} : s = 426;
	{8'd246,8'd181} : s = 427;
	{8'd246,8'd182} : s = 428;
	{8'd246,8'd183} : s = 429;
	{8'd246,8'd184} : s = 430;
	{8'd246,8'd185} : s = 431;
	{8'd246,8'd186} : s = 432;
	{8'd246,8'd187} : s = 433;
	{8'd246,8'd188} : s = 434;
	{8'd246,8'd189} : s = 435;
	{8'd246,8'd190} : s = 436;
	{8'd246,8'd191} : s = 437;
	{8'd246,8'd192} : s = 438;
	{8'd246,8'd193} : s = 439;
	{8'd246,8'd194} : s = 440;
	{8'd246,8'd195} : s = 441;
	{8'd246,8'd196} : s = 442;
	{8'd246,8'd197} : s = 443;
	{8'd246,8'd198} : s = 444;
	{8'd246,8'd199} : s = 445;
	{8'd246,8'd200} : s = 446;
	{8'd246,8'd201} : s = 447;
	{8'd246,8'd202} : s = 448;
	{8'd246,8'd203} : s = 449;
	{8'd246,8'd204} : s = 450;
	{8'd246,8'd205} : s = 451;
	{8'd246,8'd206} : s = 452;
	{8'd246,8'd207} : s = 453;
	{8'd246,8'd208} : s = 454;
	{8'd246,8'd209} : s = 455;
	{8'd246,8'd210} : s = 456;
	{8'd246,8'd211} : s = 457;
	{8'd246,8'd212} : s = 458;
	{8'd246,8'd213} : s = 459;
	{8'd246,8'd214} : s = 460;
	{8'd246,8'd215} : s = 461;
	{8'd246,8'd216} : s = 462;
	{8'd246,8'd217} : s = 463;
	{8'd246,8'd218} : s = 464;
	{8'd246,8'd219} : s = 465;
	{8'd246,8'd220} : s = 466;
	{8'd246,8'd221} : s = 467;
	{8'd246,8'd222} : s = 468;
	{8'd246,8'd223} : s = 469;
	{8'd246,8'd224} : s = 470;
	{8'd246,8'd225} : s = 471;
	{8'd246,8'd226} : s = 472;
	{8'd246,8'd227} : s = 473;
	{8'd246,8'd228} : s = 474;
	{8'd246,8'd229} : s = 475;
	{8'd246,8'd230} : s = 476;
	{8'd246,8'd231} : s = 477;
	{8'd246,8'd232} : s = 478;
	{8'd246,8'd233} : s = 479;
	{8'd246,8'd234} : s = 480;
	{8'd246,8'd235} : s = 481;
	{8'd246,8'd236} : s = 482;
	{8'd246,8'd237} : s = 483;
	{8'd246,8'd238} : s = 484;
	{8'd246,8'd239} : s = 485;
	{8'd246,8'd240} : s = 486;
	{8'd246,8'd241} : s = 487;
	{8'd246,8'd242} : s = 488;
	{8'd246,8'd243} : s = 489;
	{8'd246,8'd244} : s = 490;
	{8'd246,8'd245} : s = 491;
	{8'd246,8'd246} : s = 492;
	{8'd246,8'd247} : s = 493;
	{8'd246,8'd248} : s = 494;
	{8'd246,8'd249} : s = 495;
	{8'd246,8'd250} : s = 496;
	{8'd246,8'd251} : s = 497;
	{8'd246,8'd252} : s = 498;
	{8'd246,8'd253} : s = 499;
	{8'd246,8'd254} : s = 500;
	{8'd246,8'd255} : s = 501;
	{8'd247,8'd0} : s = 247;
	{8'd247,8'd1} : s = 248;
	{8'd247,8'd2} : s = 249;
	{8'd247,8'd3} : s = 250;
	{8'd247,8'd4} : s = 251;
	{8'd247,8'd5} : s = 252;
	{8'd247,8'd6} : s = 253;
	{8'd247,8'd7} : s = 254;
	{8'd247,8'd8} : s = 255;
	{8'd247,8'd9} : s = 256;
	{8'd247,8'd10} : s = 257;
	{8'd247,8'd11} : s = 258;
	{8'd247,8'd12} : s = 259;
	{8'd247,8'd13} : s = 260;
	{8'd247,8'd14} : s = 261;
	{8'd247,8'd15} : s = 262;
	{8'd247,8'd16} : s = 263;
	{8'd247,8'd17} : s = 264;
	{8'd247,8'd18} : s = 265;
	{8'd247,8'd19} : s = 266;
	{8'd247,8'd20} : s = 267;
	{8'd247,8'd21} : s = 268;
	{8'd247,8'd22} : s = 269;
	{8'd247,8'd23} : s = 270;
	{8'd247,8'd24} : s = 271;
	{8'd247,8'd25} : s = 272;
	{8'd247,8'd26} : s = 273;
	{8'd247,8'd27} : s = 274;
	{8'd247,8'd28} : s = 275;
	{8'd247,8'd29} : s = 276;
	{8'd247,8'd30} : s = 277;
	{8'd247,8'd31} : s = 278;
	{8'd247,8'd32} : s = 279;
	{8'd247,8'd33} : s = 280;
	{8'd247,8'd34} : s = 281;
	{8'd247,8'd35} : s = 282;
	{8'd247,8'd36} : s = 283;
	{8'd247,8'd37} : s = 284;
	{8'd247,8'd38} : s = 285;
	{8'd247,8'd39} : s = 286;
	{8'd247,8'd40} : s = 287;
	{8'd247,8'd41} : s = 288;
	{8'd247,8'd42} : s = 289;
	{8'd247,8'd43} : s = 290;
	{8'd247,8'd44} : s = 291;
	{8'd247,8'd45} : s = 292;
	{8'd247,8'd46} : s = 293;
	{8'd247,8'd47} : s = 294;
	{8'd247,8'd48} : s = 295;
	{8'd247,8'd49} : s = 296;
	{8'd247,8'd50} : s = 297;
	{8'd247,8'd51} : s = 298;
	{8'd247,8'd52} : s = 299;
	{8'd247,8'd53} : s = 300;
	{8'd247,8'd54} : s = 301;
	{8'd247,8'd55} : s = 302;
	{8'd247,8'd56} : s = 303;
	{8'd247,8'd57} : s = 304;
	{8'd247,8'd58} : s = 305;
	{8'd247,8'd59} : s = 306;
	{8'd247,8'd60} : s = 307;
	{8'd247,8'd61} : s = 308;
	{8'd247,8'd62} : s = 309;
	{8'd247,8'd63} : s = 310;
	{8'd247,8'd64} : s = 311;
	{8'd247,8'd65} : s = 312;
	{8'd247,8'd66} : s = 313;
	{8'd247,8'd67} : s = 314;
	{8'd247,8'd68} : s = 315;
	{8'd247,8'd69} : s = 316;
	{8'd247,8'd70} : s = 317;
	{8'd247,8'd71} : s = 318;
	{8'd247,8'd72} : s = 319;
	{8'd247,8'd73} : s = 320;
	{8'd247,8'd74} : s = 321;
	{8'd247,8'd75} : s = 322;
	{8'd247,8'd76} : s = 323;
	{8'd247,8'd77} : s = 324;
	{8'd247,8'd78} : s = 325;
	{8'd247,8'd79} : s = 326;
	{8'd247,8'd80} : s = 327;
	{8'd247,8'd81} : s = 328;
	{8'd247,8'd82} : s = 329;
	{8'd247,8'd83} : s = 330;
	{8'd247,8'd84} : s = 331;
	{8'd247,8'd85} : s = 332;
	{8'd247,8'd86} : s = 333;
	{8'd247,8'd87} : s = 334;
	{8'd247,8'd88} : s = 335;
	{8'd247,8'd89} : s = 336;
	{8'd247,8'd90} : s = 337;
	{8'd247,8'd91} : s = 338;
	{8'd247,8'd92} : s = 339;
	{8'd247,8'd93} : s = 340;
	{8'd247,8'd94} : s = 341;
	{8'd247,8'd95} : s = 342;
	{8'd247,8'd96} : s = 343;
	{8'd247,8'd97} : s = 344;
	{8'd247,8'd98} : s = 345;
	{8'd247,8'd99} : s = 346;
	{8'd247,8'd100} : s = 347;
	{8'd247,8'd101} : s = 348;
	{8'd247,8'd102} : s = 349;
	{8'd247,8'd103} : s = 350;
	{8'd247,8'd104} : s = 351;
	{8'd247,8'd105} : s = 352;
	{8'd247,8'd106} : s = 353;
	{8'd247,8'd107} : s = 354;
	{8'd247,8'd108} : s = 355;
	{8'd247,8'd109} : s = 356;
	{8'd247,8'd110} : s = 357;
	{8'd247,8'd111} : s = 358;
	{8'd247,8'd112} : s = 359;
	{8'd247,8'd113} : s = 360;
	{8'd247,8'd114} : s = 361;
	{8'd247,8'd115} : s = 362;
	{8'd247,8'd116} : s = 363;
	{8'd247,8'd117} : s = 364;
	{8'd247,8'd118} : s = 365;
	{8'd247,8'd119} : s = 366;
	{8'd247,8'd120} : s = 367;
	{8'd247,8'd121} : s = 368;
	{8'd247,8'd122} : s = 369;
	{8'd247,8'd123} : s = 370;
	{8'd247,8'd124} : s = 371;
	{8'd247,8'd125} : s = 372;
	{8'd247,8'd126} : s = 373;
	{8'd247,8'd127} : s = 374;
	{8'd247,8'd128} : s = 375;
	{8'd247,8'd129} : s = 376;
	{8'd247,8'd130} : s = 377;
	{8'd247,8'd131} : s = 378;
	{8'd247,8'd132} : s = 379;
	{8'd247,8'd133} : s = 380;
	{8'd247,8'd134} : s = 381;
	{8'd247,8'd135} : s = 382;
	{8'd247,8'd136} : s = 383;
	{8'd247,8'd137} : s = 384;
	{8'd247,8'd138} : s = 385;
	{8'd247,8'd139} : s = 386;
	{8'd247,8'd140} : s = 387;
	{8'd247,8'd141} : s = 388;
	{8'd247,8'd142} : s = 389;
	{8'd247,8'd143} : s = 390;
	{8'd247,8'd144} : s = 391;
	{8'd247,8'd145} : s = 392;
	{8'd247,8'd146} : s = 393;
	{8'd247,8'd147} : s = 394;
	{8'd247,8'd148} : s = 395;
	{8'd247,8'd149} : s = 396;
	{8'd247,8'd150} : s = 397;
	{8'd247,8'd151} : s = 398;
	{8'd247,8'd152} : s = 399;
	{8'd247,8'd153} : s = 400;
	{8'd247,8'd154} : s = 401;
	{8'd247,8'd155} : s = 402;
	{8'd247,8'd156} : s = 403;
	{8'd247,8'd157} : s = 404;
	{8'd247,8'd158} : s = 405;
	{8'd247,8'd159} : s = 406;
	{8'd247,8'd160} : s = 407;
	{8'd247,8'd161} : s = 408;
	{8'd247,8'd162} : s = 409;
	{8'd247,8'd163} : s = 410;
	{8'd247,8'd164} : s = 411;
	{8'd247,8'd165} : s = 412;
	{8'd247,8'd166} : s = 413;
	{8'd247,8'd167} : s = 414;
	{8'd247,8'd168} : s = 415;
	{8'd247,8'd169} : s = 416;
	{8'd247,8'd170} : s = 417;
	{8'd247,8'd171} : s = 418;
	{8'd247,8'd172} : s = 419;
	{8'd247,8'd173} : s = 420;
	{8'd247,8'd174} : s = 421;
	{8'd247,8'd175} : s = 422;
	{8'd247,8'd176} : s = 423;
	{8'd247,8'd177} : s = 424;
	{8'd247,8'd178} : s = 425;
	{8'd247,8'd179} : s = 426;
	{8'd247,8'd180} : s = 427;
	{8'd247,8'd181} : s = 428;
	{8'd247,8'd182} : s = 429;
	{8'd247,8'd183} : s = 430;
	{8'd247,8'd184} : s = 431;
	{8'd247,8'd185} : s = 432;
	{8'd247,8'd186} : s = 433;
	{8'd247,8'd187} : s = 434;
	{8'd247,8'd188} : s = 435;
	{8'd247,8'd189} : s = 436;
	{8'd247,8'd190} : s = 437;
	{8'd247,8'd191} : s = 438;
	{8'd247,8'd192} : s = 439;
	{8'd247,8'd193} : s = 440;
	{8'd247,8'd194} : s = 441;
	{8'd247,8'd195} : s = 442;
	{8'd247,8'd196} : s = 443;
	{8'd247,8'd197} : s = 444;
	{8'd247,8'd198} : s = 445;
	{8'd247,8'd199} : s = 446;
	{8'd247,8'd200} : s = 447;
	{8'd247,8'd201} : s = 448;
	{8'd247,8'd202} : s = 449;
	{8'd247,8'd203} : s = 450;
	{8'd247,8'd204} : s = 451;
	{8'd247,8'd205} : s = 452;
	{8'd247,8'd206} : s = 453;
	{8'd247,8'd207} : s = 454;
	{8'd247,8'd208} : s = 455;
	{8'd247,8'd209} : s = 456;
	{8'd247,8'd210} : s = 457;
	{8'd247,8'd211} : s = 458;
	{8'd247,8'd212} : s = 459;
	{8'd247,8'd213} : s = 460;
	{8'd247,8'd214} : s = 461;
	{8'd247,8'd215} : s = 462;
	{8'd247,8'd216} : s = 463;
	{8'd247,8'd217} : s = 464;
	{8'd247,8'd218} : s = 465;
	{8'd247,8'd219} : s = 466;
	{8'd247,8'd220} : s = 467;
	{8'd247,8'd221} : s = 468;
	{8'd247,8'd222} : s = 469;
	{8'd247,8'd223} : s = 470;
	{8'd247,8'd224} : s = 471;
	{8'd247,8'd225} : s = 472;
	{8'd247,8'd226} : s = 473;
	{8'd247,8'd227} : s = 474;
	{8'd247,8'd228} : s = 475;
	{8'd247,8'd229} : s = 476;
	{8'd247,8'd230} : s = 477;
	{8'd247,8'd231} : s = 478;
	{8'd247,8'd232} : s = 479;
	{8'd247,8'd233} : s = 480;
	{8'd247,8'd234} : s = 481;
	{8'd247,8'd235} : s = 482;
	{8'd247,8'd236} : s = 483;
	{8'd247,8'd237} : s = 484;
	{8'd247,8'd238} : s = 485;
	{8'd247,8'd239} : s = 486;
	{8'd247,8'd240} : s = 487;
	{8'd247,8'd241} : s = 488;
	{8'd247,8'd242} : s = 489;
	{8'd247,8'd243} : s = 490;
	{8'd247,8'd244} : s = 491;
	{8'd247,8'd245} : s = 492;
	{8'd247,8'd246} : s = 493;
	{8'd247,8'd247} : s = 494;
	{8'd247,8'd248} : s = 495;
	{8'd247,8'd249} : s = 496;
	{8'd247,8'd250} : s = 497;
	{8'd247,8'd251} : s = 498;
	{8'd247,8'd252} : s = 499;
	{8'd247,8'd253} : s = 500;
	{8'd247,8'd254} : s = 501;
	{8'd247,8'd255} : s = 502;
	{8'd248,8'd0} : s = 248;
	{8'd248,8'd1} : s = 249;
	{8'd248,8'd2} : s = 250;
	{8'd248,8'd3} : s = 251;
	{8'd248,8'd4} : s = 252;
	{8'd248,8'd5} : s = 253;
	{8'd248,8'd6} : s = 254;
	{8'd248,8'd7} : s = 255;
	{8'd248,8'd8} : s = 256;
	{8'd248,8'd9} : s = 257;
	{8'd248,8'd10} : s = 258;
	{8'd248,8'd11} : s = 259;
	{8'd248,8'd12} : s = 260;
	{8'd248,8'd13} : s = 261;
	{8'd248,8'd14} : s = 262;
	{8'd248,8'd15} : s = 263;
	{8'd248,8'd16} : s = 264;
	{8'd248,8'd17} : s = 265;
	{8'd248,8'd18} : s = 266;
	{8'd248,8'd19} : s = 267;
	{8'd248,8'd20} : s = 268;
	{8'd248,8'd21} : s = 269;
	{8'd248,8'd22} : s = 270;
	{8'd248,8'd23} : s = 271;
	{8'd248,8'd24} : s = 272;
	{8'd248,8'd25} : s = 273;
	{8'd248,8'd26} : s = 274;
	{8'd248,8'd27} : s = 275;
	{8'd248,8'd28} : s = 276;
	{8'd248,8'd29} : s = 277;
	{8'd248,8'd30} : s = 278;
	{8'd248,8'd31} : s = 279;
	{8'd248,8'd32} : s = 280;
	{8'd248,8'd33} : s = 281;
	{8'd248,8'd34} : s = 282;
	{8'd248,8'd35} : s = 283;
	{8'd248,8'd36} : s = 284;
	{8'd248,8'd37} : s = 285;
	{8'd248,8'd38} : s = 286;
	{8'd248,8'd39} : s = 287;
	{8'd248,8'd40} : s = 288;
	{8'd248,8'd41} : s = 289;
	{8'd248,8'd42} : s = 290;
	{8'd248,8'd43} : s = 291;
	{8'd248,8'd44} : s = 292;
	{8'd248,8'd45} : s = 293;
	{8'd248,8'd46} : s = 294;
	{8'd248,8'd47} : s = 295;
	{8'd248,8'd48} : s = 296;
	{8'd248,8'd49} : s = 297;
	{8'd248,8'd50} : s = 298;
	{8'd248,8'd51} : s = 299;
	{8'd248,8'd52} : s = 300;
	{8'd248,8'd53} : s = 301;
	{8'd248,8'd54} : s = 302;
	{8'd248,8'd55} : s = 303;
	{8'd248,8'd56} : s = 304;
	{8'd248,8'd57} : s = 305;
	{8'd248,8'd58} : s = 306;
	{8'd248,8'd59} : s = 307;
	{8'd248,8'd60} : s = 308;
	{8'd248,8'd61} : s = 309;
	{8'd248,8'd62} : s = 310;
	{8'd248,8'd63} : s = 311;
	{8'd248,8'd64} : s = 312;
	{8'd248,8'd65} : s = 313;
	{8'd248,8'd66} : s = 314;
	{8'd248,8'd67} : s = 315;
	{8'd248,8'd68} : s = 316;
	{8'd248,8'd69} : s = 317;
	{8'd248,8'd70} : s = 318;
	{8'd248,8'd71} : s = 319;
	{8'd248,8'd72} : s = 320;
	{8'd248,8'd73} : s = 321;
	{8'd248,8'd74} : s = 322;
	{8'd248,8'd75} : s = 323;
	{8'd248,8'd76} : s = 324;
	{8'd248,8'd77} : s = 325;
	{8'd248,8'd78} : s = 326;
	{8'd248,8'd79} : s = 327;
	{8'd248,8'd80} : s = 328;
	{8'd248,8'd81} : s = 329;
	{8'd248,8'd82} : s = 330;
	{8'd248,8'd83} : s = 331;
	{8'd248,8'd84} : s = 332;
	{8'd248,8'd85} : s = 333;
	{8'd248,8'd86} : s = 334;
	{8'd248,8'd87} : s = 335;
	{8'd248,8'd88} : s = 336;
	{8'd248,8'd89} : s = 337;
	{8'd248,8'd90} : s = 338;
	{8'd248,8'd91} : s = 339;
	{8'd248,8'd92} : s = 340;
	{8'd248,8'd93} : s = 341;
	{8'd248,8'd94} : s = 342;
	{8'd248,8'd95} : s = 343;
	{8'd248,8'd96} : s = 344;
	{8'd248,8'd97} : s = 345;
	{8'd248,8'd98} : s = 346;
	{8'd248,8'd99} : s = 347;
	{8'd248,8'd100} : s = 348;
	{8'd248,8'd101} : s = 349;
	{8'd248,8'd102} : s = 350;
	{8'd248,8'd103} : s = 351;
	{8'd248,8'd104} : s = 352;
	{8'd248,8'd105} : s = 353;
	{8'd248,8'd106} : s = 354;
	{8'd248,8'd107} : s = 355;
	{8'd248,8'd108} : s = 356;
	{8'd248,8'd109} : s = 357;
	{8'd248,8'd110} : s = 358;
	{8'd248,8'd111} : s = 359;
	{8'd248,8'd112} : s = 360;
	{8'd248,8'd113} : s = 361;
	{8'd248,8'd114} : s = 362;
	{8'd248,8'd115} : s = 363;
	{8'd248,8'd116} : s = 364;
	{8'd248,8'd117} : s = 365;
	{8'd248,8'd118} : s = 366;
	{8'd248,8'd119} : s = 367;
	{8'd248,8'd120} : s = 368;
	{8'd248,8'd121} : s = 369;
	{8'd248,8'd122} : s = 370;
	{8'd248,8'd123} : s = 371;
	{8'd248,8'd124} : s = 372;
	{8'd248,8'd125} : s = 373;
	{8'd248,8'd126} : s = 374;
	{8'd248,8'd127} : s = 375;
	{8'd248,8'd128} : s = 376;
	{8'd248,8'd129} : s = 377;
	{8'd248,8'd130} : s = 378;
	{8'd248,8'd131} : s = 379;
	{8'd248,8'd132} : s = 380;
	{8'd248,8'd133} : s = 381;
	{8'd248,8'd134} : s = 382;
	{8'd248,8'd135} : s = 383;
	{8'd248,8'd136} : s = 384;
	{8'd248,8'd137} : s = 385;
	{8'd248,8'd138} : s = 386;
	{8'd248,8'd139} : s = 387;
	{8'd248,8'd140} : s = 388;
	{8'd248,8'd141} : s = 389;
	{8'd248,8'd142} : s = 390;
	{8'd248,8'd143} : s = 391;
	{8'd248,8'd144} : s = 392;
	{8'd248,8'd145} : s = 393;
	{8'd248,8'd146} : s = 394;
	{8'd248,8'd147} : s = 395;
	{8'd248,8'd148} : s = 396;
	{8'd248,8'd149} : s = 397;
	{8'd248,8'd150} : s = 398;
	{8'd248,8'd151} : s = 399;
	{8'd248,8'd152} : s = 400;
	{8'd248,8'd153} : s = 401;
	{8'd248,8'd154} : s = 402;
	{8'd248,8'd155} : s = 403;
	{8'd248,8'd156} : s = 404;
	{8'd248,8'd157} : s = 405;
	{8'd248,8'd158} : s = 406;
	{8'd248,8'd159} : s = 407;
	{8'd248,8'd160} : s = 408;
	{8'd248,8'd161} : s = 409;
	{8'd248,8'd162} : s = 410;
	{8'd248,8'd163} : s = 411;
	{8'd248,8'd164} : s = 412;
	{8'd248,8'd165} : s = 413;
	{8'd248,8'd166} : s = 414;
	{8'd248,8'd167} : s = 415;
	{8'd248,8'd168} : s = 416;
	{8'd248,8'd169} : s = 417;
	{8'd248,8'd170} : s = 418;
	{8'd248,8'd171} : s = 419;
	{8'd248,8'd172} : s = 420;
	{8'd248,8'd173} : s = 421;
	{8'd248,8'd174} : s = 422;
	{8'd248,8'd175} : s = 423;
	{8'd248,8'd176} : s = 424;
	{8'd248,8'd177} : s = 425;
	{8'd248,8'd178} : s = 426;
	{8'd248,8'd179} : s = 427;
	{8'd248,8'd180} : s = 428;
	{8'd248,8'd181} : s = 429;
	{8'd248,8'd182} : s = 430;
	{8'd248,8'd183} : s = 431;
	{8'd248,8'd184} : s = 432;
	{8'd248,8'd185} : s = 433;
	{8'd248,8'd186} : s = 434;
	{8'd248,8'd187} : s = 435;
	{8'd248,8'd188} : s = 436;
	{8'd248,8'd189} : s = 437;
	{8'd248,8'd190} : s = 438;
	{8'd248,8'd191} : s = 439;
	{8'd248,8'd192} : s = 440;
	{8'd248,8'd193} : s = 441;
	{8'd248,8'd194} : s = 442;
	{8'd248,8'd195} : s = 443;
	{8'd248,8'd196} : s = 444;
	{8'd248,8'd197} : s = 445;
	{8'd248,8'd198} : s = 446;
	{8'd248,8'd199} : s = 447;
	{8'd248,8'd200} : s = 448;
	{8'd248,8'd201} : s = 449;
	{8'd248,8'd202} : s = 450;
	{8'd248,8'd203} : s = 451;
	{8'd248,8'd204} : s = 452;
	{8'd248,8'd205} : s = 453;
	{8'd248,8'd206} : s = 454;
	{8'd248,8'd207} : s = 455;
	{8'd248,8'd208} : s = 456;
	{8'd248,8'd209} : s = 457;
	{8'd248,8'd210} : s = 458;
	{8'd248,8'd211} : s = 459;
	{8'd248,8'd212} : s = 460;
	{8'd248,8'd213} : s = 461;
	{8'd248,8'd214} : s = 462;
	{8'd248,8'd215} : s = 463;
	{8'd248,8'd216} : s = 464;
	{8'd248,8'd217} : s = 465;
	{8'd248,8'd218} : s = 466;
	{8'd248,8'd219} : s = 467;
	{8'd248,8'd220} : s = 468;
	{8'd248,8'd221} : s = 469;
	{8'd248,8'd222} : s = 470;
	{8'd248,8'd223} : s = 471;
	{8'd248,8'd224} : s = 472;
	{8'd248,8'd225} : s = 473;
	{8'd248,8'd226} : s = 474;
	{8'd248,8'd227} : s = 475;
	{8'd248,8'd228} : s = 476;
	{8'd248,8'd229} : s = 477;
	{8'd248,8'd230} : s = 478;
	{8'd248,8'd231} : s = 479;
	{8'd248,8'd232} : s = 480;
	{8'd248,8'd233} : s = 481;
	{8'd248,8'd234} : s = 482;
	{8'd248,8'd235} : s = 483;
	{8'd248,8'd236} : s = 484;
	{8'd248,8'd237} : s = 485;
	{8'd248,8'd238} : s = 486;
	{8'd248,8'd239} : s = 487;
	{8'd248,8'd240} : s = 488;
	{8'd248,8'd241} : s = 489;
	{8'd248,8'd242} : s = 490;
	{8'd248,8'd243} : s = 491;
	{8'd248,8'd244} : s = 492;
	{8'd248,8'd245} : s = 493;
	{8'd248,8'd246} : s = 494;
	{8'd248,8'd247} : s = 495;
	{8'd248,8'd248} : s = 496;
	{8'd248,8'd249} : s = 497;
	{8'd248,8'd250} : s = 498;
	{8'd248,8'd251} : s = 499;
	{8'd248,8'd252} : s = 500;
	{8'd248,8'd253} : s = 501;
	{8'd248,8'd254} : s = 502;
	{8'd248,8'd255} : s = 503;
	{8'd249,8'd0} : s = 249;
	{8'd249,8'd1} : s = 250;
	{8'd249,8'd2} : s = 251;
	{8'd249,8'd3} : s = 252;
	{8'd249,8'd4} : s = 253;
	{8'd249,8'd5} : s = 254;
	{8'd249,8'd6} : s = 255;
	{8'd249,8'd7} : s = 256;
	{8'd249,8'd8} : s = 257;
	{8'd249,8'd9} : s = 258;
	{8'd249,8'd10} : s = 259;
	{8'd249,8'd11} : s = 260;
	{8'd249,8'd12} : s = 261;
	{8'd249,8'd13} : s = 262;
	{8'd249,8'd14} : s = 263;
	{8'd249,8'd15} : s = 264;
	{8'd249,8'd16} : s = 265;
	{8'd249,8'd17} : s = 266;
	{8'd249,8'd18} : s = 267;
	{8'd249,8'd19} : s = 268;
	{8'd249,8'd20} : s = 269;
	{8'd249,8'd21} : s = 270;
	{8'd249,8'd22} : s = 271;
	{8'd249,8'd23} : s = 272;
	{8'd249,8'd24} : s = 273;
	{8'd249,8'd25} : s = 274;
	{8'd249,8'd26} : s = 275;
	{8'd249,8'd27} : s = 276;
	{8'd249,8'd28} : s = 277;
	{8'd249,8'd29} : s = 278;
	{8'd249,8'd30} : s = 279;
	{8'd249,8'd31} : s = 280;
	{8'd249,8'd32} : s = 281;
	{8'd249,8'd33} : s = 282;
	{8'd249,8'd34} : s = 283;
	{8'd249,8'd35} : s = 284;
	{8'd249,8'd36} : s = 285;
	{8'd249,8'd37} : s = 286;
	{8'd249,8'd38} : s = 287;
	{8'd249,8'd39} : s = 288;
	{8'd249,8'd40} : s = 289;
	{8'd249,8'd41} : s = 290;
	{8'd249,8'd42} : s = 291;
	{8'd249,8'd43} : s = 292;
	{8'd249,8'd44} : s = 293;
	{8'd249,8'd45} : s = 294;
	{8'd249,8'd46} : s = 295;
	{8'd249,8'd47} : s = 296;
	{8'd249,8'd48} : s = 297;
	{8'd249,8'd49} : s = 298;
	{8'd249,8'd50} : s = 299;
	{8'd249,8'd51} : s = 300;
	{8'd249,8'd52} : s = 301;
	{8'd249,8'd53} : s = 302;
	{8'd249,8'd54} : s = 303;
	{8'd249,8'd55} : s = 304;
	{8'd249,8'd56} : s = 305;
	{8'd249,8'd57} : s = 306;
	{8'd249,8'd58} : s = 307;
	{8'd249,8'd59} : s = 308;
	{8'd249,8'd60} : s = 309;
	{8'd249,8'd61} : s = 310;
	{8'd249,8'd62} : s = 311;
	{8'd249,8'd63} : s = 312;
	{8'd249,8'd64} : s = 313;
	{8'd249,8'd65} : s = 314;
	{8'd249,8'd66} : s = 315;
	{8'd249,8'd67} : s = 316;
	{8'd249,8'd68} : s = 317;
	{8'd249,8'd69} : s = 318;
	{8'd249,8'd70} : s = 319;
	{8'd249,8'd71} : s = 320;
	{8'd249,8'd72} : s = 321;
	{8'd249,8'd73} : s = 322;
	{8'd249,8'd74} : s = 323;
	{8'd249,8'd75} : s = 324;
	{8'd249,8'd76} : s = 325;
	{8'd249,8'd77} : s = 326;
	{8'd249,8'd78} : s = 327;
	{8'd249,8'd79} : s = 328;
	{8'd249,8'd80} : s = 329;
	{8'd249,8'd81} : s = 330;
	{8'd249,8'd82} : s = 331;
	{8'd249,8'd83} : s = 332;
	{8'd249,8'd84} : s = 333;
	{8'd249,8'd85} : s = 334;
	{8'd249,8'd86} : s = 335;
	{8'd249,8'd87} : s = 336;
	{8'd249,8'd88} : s = 337;
	{8'd249,8'd89} : s = 338;
	{8'd249,8'd90} : s = 339;
	{8'd249,8'd91} : s = 340;
	{8'd249,8'd92} : s = 341;
	{8'd249,8'd93} : s = 342;
	{8'd249,8'd94} : s = 343;
	{8'd249,8'd95} : s = 344;
	{8'd249,8'd96} : s = 345;
	{8'd249,8'd97} : s = 346;
	{8'd249,8'd98} : s = 347;
	{8'd249,8'd99} : s = 348;
	{8'd249,8'd100} : s = 349;
	{8'd249,8'd101} : s = 350;
	{8'd249,8'd102} : s = 351;
	{8'd249,8'd103} : s = 352;
	{8'd249,8'd104} : s = 353;
	{8'd249,8'd105} : s = 354;
	{8'd249,8'd106} : s = 355;
	{8'd249,8'd107} : s = 356;
	{8'd249,8'd108} : s = 357;
	{8'd249,8'd109} : s = 358;
	{8'd249,8'd110} : s = 359;
	{8'd249,8'd111} : s = 360;
	{8'd249,8'd112} : s = 361;
	{8'd249,8'd113} : s = 362;
	{8'd249,8'd114} : s = 363;
	{8'd249,8'd115} : s = 364;
	{8'd249,8'd116} : s = 365;
	{8'd249,8'd117} : s = 366;
	{8'd249,8'd118} : s = 367;
	{8'd249,8'd119} : s = 368;
	{8'd249,8'd120} : s = 369;
	{8'd249,8'd121} : s = 370;
	{8'd249,8'd122} : s = 371;
	{8'd249,8'd123} : s = 372;
	{8'd249,8'd124} : s = 373;
	{8'd249,8'd125} : s = 374;
	{8'd249,8'd126} : s = 375;
	{8'd249,8'd127} : s = 376;
	{8'd249,8'd128} : s = 377;
	{8'd249,8'd129} : s = 378;
	{8'd249,8'd130} : s = 379;
	{8'd249,8'd131} : s = 380;
	{8'd249,8'd132} : s = 381;
	{8'd249,8'd133} : s = 382;
	{8'd249,8'd134} : s = 383;
	{8'd249,8'd135} : s = 384;
	{8'd249,8'd136} : s = 385;
	{8'd249,8'd137} : s = 386;
	{8'd249,8'd138} : s = 387;
	{8'd249,8'd139} : s = 388;
	{8'd249,8'd140} : s = 389;
	{8'd249,8'd141} : s = 390;
	{8'd249,8'd142} : s = 391;
	{8'd249,8'd143} : s = 392;
	{8'd249,8'd144} : s = 393;
	{8'd249,8'd145} : s = 394;
	{8'd249,8'd146} : s = 395;
	{8'd249,8'd147} : s = 396;
	{8'd249,8'd148} : s = 397;
	{8'd249,8'd149} : s = 398;
	{8'd249,8'd150} : s = 399;
	{8'd249,8'd151} : s = 400;
	{8'd249,8'd152} : s = 401;
	{8'd249,8'd153} : s = 402;
	{8'd249,8'd154} : s = 403;
	{8'd249,8'd155} : s = 404;
	{8'd249,8'd156} : s = 405;
	{8'd249,8'd157} : s = 406;
	{8'd249,8'd158} : s = 407;
	{8'd249,8'd159} : s = 408;
	{8'd249,8'd160} : s = 409;
	{8'd249,8'd161} : s = 410;
	{8'd249,8'd162} : s = 411;
	{8'd249,8'd163} : s = 412;
	{8'd249,8'd164} : s = 413;
	{8'd249,8'd165} : s = 414;
	{8'd249,8'd166} : s = 415;
	{8'd249,8'd167} : s = 416;
	{8'd249,8'd168} : s = 417;
	{8'd249,8'd169} : s = 418;
	{8'd249,8'd170} : s = 419;
	{8'd249,8'd171} : s = 420;
	{8'd249,8'd172} : s = 421;
	{8'd249,8'd173} : s = 422;
	{8'd249,8'd174} : s = 423;
	{8'd249,8'd175} : s = 424;
	{8'd249,8'd176} : s = 425;
	{8'd249,8'd177} : s = 426;
	{8'd249,8'd178} : s = 427;
	{8'd249,8'd179} : s = 428;
	{8'd249,8'd180} : s = 429;
	{8'd249,8'd181} : s = 430;
	{8'd249,8'd182} : s = 431;
	{8'd249,8'd183} : s = 432;
	{8'd249,8'd184} : s = 433;
	{8'd249,8'd185} : s = 434;
	{8'd249,8'd186} : s = 435;
	{8'd249,8'd187} : s = 436;
	{8'd249,8'd188} : s = 437;
	{8'd249,8'd189} : s = 438;
	{8'd249,8'd190} : s = 439;
	{8'd249,8'd191} : s = 440;
	{8'd249,8'd192} : s = 441;
	{8'd249,8'd193} : s = 442;
	{8'd249,8'd194} : s = 443;
	{8'd249,8'd195} : s = 444;
	{8'd249,8'd196} : s = 445;
	{8'd249,8'd197} : s = 446;
	{8'd249,8'd198} : s = 447;
	{8'd249,8'd199} : s = 448;
	{8'd249,8'd200} : s = 449;
	{8'd249,8'd201} : s = 450;
	{8'd249,8'd202} : s = 451;
	{8'd249,8'd203} : s = 452;
	{8'd249,8'd204} : s = 453;
	{8'd249,8'd205} : s = 454;
	{8'd249,8'd206} : s = 455;
	{8'd249,8'd207} : s = 456;
	{8'd249,8'd208} : s = 457;
	{8'd249,8'd209} : s = 458;
	{8'd249,8'd210} : s = 459;
	{8'd249,8'd211} : s = 460;
	{8'd249,8'd212} : s = 461;
	{8'd249,8'd213} : s = 462;
	{8'd249,8'd214} : s = 463;
	{8'd249,8'd215} : s = 464;
	{8'd249,8'd216} : s = 465;
	{8'd249,8'd217} : s = 466;
	{8'd249,8'd218} : s = 467;
	{8'd249,8'd219} : s = 468;
	{8'd249,8'd220} : s = 469;
	{8'd249,8'd221} : s = 470;
	{8'd249,8'd222} : s = 471;
	{8'd249,8'd223} : s = 472;
	{8'd249,8'd224} : s = 473;
	{8'd249,8'd225} : s = 474;
	{8'd249,8'd226} : s = 475;
	{8'd249,8'd227} : s = 476;
	{8'd249,8'd228} : s = 477;
	{8'd249,8'd229} : s = 478;
	{8'd249,8'd230} : s = 479;
	{8'd249,8'd231} : s = 480;
	{8'd249,8'd232} : s = 481;
	{8'd249,8'd233} : s = 482;
	{8'd249,8'd234} : s = 483;
	{8'd249,8'd235} : s = 484;
	{8'd249,8'd236} : s = 485;
	{8'd249,8'd237} : s = 486;
	{8'd249,8'd238} : s = 487;
	{8'd249,8'd239} : s = 488;
	{8'd249,8'd240} : s = 489;
	{8'd249,8'd241} : s = 490;
	{8'd249,8'd242} : s = 491;
	{8'd249,8'd243} : s = 492;
	{8'd249,8'd244} : s = 493;
	{8'd249,8'd245} : s = 494;
	{8'd249,8'd246} : s = 495;
	{8'd249,8'd247} : s = 496;
	{8'd249,8'd248} : s = 497;
	{8'd249,8'd249} : s = 498;
	{8'd249,8'd250} : s = 499;
	{8'd249,8'd251} : s = 500;
	{8'd249,8'd252} : s = 501;
	{8'd249,8'd253} : s = 502;
	{8'd249,8'd254} : s = 503;
	{8'd249,8'd255} : s = 504;
	{8'd250,8'd0} : s = 250;
	{8'd250,8'd1} : s = 251;
	{8'd250,8'd2} : s = 252;
	{8'd250,8'd3} : s = 253;
	{8'd250,8'd4} : s = 254;
	{8'd250,8'd5} : s = 255;
	{8'd250,8'd6} : s = 256;
	{8'd250,8'd7} : s = 257;
	{8'd250,8'd8} : s = 258;
	{8'd250,8'd9} : s = 259;
	{8'd250,8'd10} : s = 260;
	{8'd250,8'd11} : s = 261;
	{8'd250,8'd12} : s = 262;
	{8'd250,8'd13} : s = 263;
	{8'd250,8'd14} : s = 264;
	{8'd250,8'd15} : s = 265;
	{8'd250,8'd16} : s = 266;
	{8'd250,8'd17} : s = 267;
	{8'd250,8'd18} : s = 268;
	{8'd250,8'd19} : s = 269;
	{8'd250,8'd20} : s = 270;
	{8'd250,8'd21} : s = 271;
	{8'd250,8'd22} : s = 272;
	{8'd250,8'd23} : s = 273;
	{8'd250,8'd24} : s = 274;
	{8'd250,8'd25} : s = 275;
	{8'd250,8'd26} : s = 276;
	{8'd250,8'd27} : s = 277;
	{8'd250,8'd28} : s = 278;
	{8'd250,8'd29} : s = 279;
	{8'd250,8'd30} : s = 280;
	{8'd250,8'd31} : s = 281;
	{8'd250,8'd32} : s = 282;
	{8'd250,8'd33} : s = 283;
	{8'd250,8'd34} : s = 284;
	{8'd250,8'd35} : s = 285;
	{8'd250,8'd36} : s = 286;
	{8'd250,8'd37} : s = 287;
	{8'd250,8'd38} : s = 288;
	{8'd250,8'd39} : s = 289;
	{8'd250,8'd40} : s = 290;
	{8'd250,8'd41} : s = 291;
	{8'd250,8'd42} : s = 292;
	{8'd250,8'd43} : s = 293;
	{8'd250,8'd44} : s = 294;
	{8'd250,8'd45} : s = 295;
	{8'd250,8'd46} : s = 296;
	{8'd250,8'd47} : s = 297;
	{8'd250,8'd48} : s = 298;
	{8'd250,8'd49} : s = 299;
	{8'd250,8'd50} : s = 300;
	{8'd250,8'd51} : s = 301;
	{8'd250,8'd52} : s = 302;
	{8'd250,8'd53} : s = 303;
	{8'd250,8'd54} : s = 304;
	{8'd250,8'd55} : s = 305;
	{8'd250,8'd56} : s = 306;
	{8'd250,8'd57} : s = 307;
	{8'd250,8'd58} : s = 308;
	{8'd250,8'd59} : s = 309;
	{8'd250,8'd60} : s = 310;
	{8'd250,8'd61} : s = 311;
	{8'd250,8'd62} : s = 312;
	{8'd250,8'd63} : s = 313;
	{8'd250,8'd64} : s = 314;
	{8'd250,8'd65} : s = 315;
	{8'd250,8'd66} : s = 316;
	{8'd250,8'd67} : s = 317;
	{8'd250,8'd68} : s = 318;
	{8'd250,8'd69} : s = 319;
	{8'd250,8'd70} : s = 320;
	{8'd250,8'd71} : s = 321;
	{8'd250,8'd72} : s = 322;
	{8'd250,8'd73} : s = 323;
	{8'd250,8'd74} : s = 324;
	{8'd250,8'd75} : s = 325;
	{8'd250,8'd76} : s = 326;
	{8'd250,8'd77} : s = 327;
	{8'd250,8'd78} : s = 328;
	{8'd250,8'd79} : s = 329;
	{8'd250,8'd80} : s = 330;
	{8'd250,8'd81} : s = 331;
	{8'd250,8'd82} : s = 332;
	{8'd250,8'd83} : s = 333;
	{8'd250,8'd84} : s = 334;
	{8'd250,8'd85} : s = 335;
	{8'd250,8'd86} : s = 336;
	{8'd250,8'd87} : s = 337;
	{8'd250,8'd88} : s = 338;
	{8'd250,8'd89} : s = 339;
	{8'd250,8'd90} : s = 340;
	{8'd250,8'd91} : s = 341;
	{8'd250,8'd92} : s = 342;
	{8'd250,8'd93} : s = 343;
	{8'd250,8'd94} : s = 344;
	{8'd250,8'd95} : s = 345;
	{8'd250,8'd96} : s = 346;
	{8'd250,8'd97} : s = 347;
	{8'd250,8'd98} : s = 348;
	{8'd250,8'd99} : s = 349;
	{8'd250,8'd100} : s = 350;
	{8'd250,8'd101} : s = 351;
	{8'd250,8'd102} : s = 352;
	{8'd250,8'd103} : s = 353;
	{8'd250,8'd104} : s = 354;
	{8'd250,8'd105} : s = 355;
	{8'd250,8'd106} : s = 356;
	{8'd250,8'd107} : s = 357;
	{8'd250,8'd108} : s = 358;
	{8'd250,8'd109} : s = 359;
	{8'd250,8'd110} : s = 360;
	{8'd250,8'd111} : s = 361;
	{8'd250,8'd112} : s = 362;
	{8'd250,8'd113} : s = 363;
	{8'd250,8'd114} : s = 364;
	{8'd250,8'd115} : s = 365;
	{8'd250,8'd116} : s = 366;
	{8'd250,8'd117} : s = 367;
	{8'd250,8'd118} : s = 368;
	{8'd250,8'd119} : s = 369;
	{8'd250,8'd120} : s = 370;
	{8'd250,8'd121} : s = 371;
	{8'd250,8'd122} : s = 372;
	{8'd250,8'd123} : s = 373;
	{8'd250,8'd124} : s = 374;
	{8'd250,8'd125} : s = 375;
	{8'd250,8'd126} : s = 376;
	{8'd250,8'd127} : s = 377;
	{8'd250,8'd128} : s = 378;
	{8'd250,8'd129} : s = 379;
	{8'd250,8'd130} : s = 380;
	{8'd250,8'd131} : s = 381;
	{8'd250,8'd132} : s = 382;
	{8'd250,8'd133} : s = 383;
	{8'd250,8'd134} : s = 384;
	{8'd250,8'd135} : s = 385;
	{8'd250,8'd136} : s = 386;
	{8'd250,8'd137} : s = 387;
	{8'd250,8'd138} : s = 388;
	{8'd250,8'd139} : s = 389;
	{8'd250,8'd140} : s = 390;
	{8'd250,8'd141} : s = 391;
	{8'd250,8'd142} : s = 392;
	{8'd250,8'd143} : s = 393;
	{8'd250,8'd144} : s = 394;
	{8'd250,8'd145} : s = 395;
	{8'd250,8'd146} : s = 396;
	{8'd250,8'd147} : s = 397;
	{8'd250,8'd148} : s = 398;
	{8'd250,8'd149} : s = 399;
	{8'd250,8'd150} : s = 400;
	{8'd250,8'd151} : s = 401;
	{8'd250,8'd152} : s = 402;
	{8'd250,8'd153} : s = 403;
	{8'd250,8'd154} : s = 404;
	{8'd250,8'd155} : s = 405;
	{8'd250,8'd156} : s = 406;
	{8'd250,8'd157} : s = 407;
	{8'd250,8'd158} : s = 408;
	{8'd250,8'd159} : s = 409;
	{8'd250,8'd160} : s = 410;
	{8'd250,8'd161} : s = 411;
	{8'd250,8'd162} : s = 412;
	{8'd250,8'd163} : s = 413;
	{8'd250,8'd164} : s = 414;
	{8'd250,8'd165} : s = 415;
	{8'd250,8'd166} : s = 416;
	{8'd250,8'd167} : s = 417;
	{8'd250,8'd168} : s = 418;
	{8'd250,8'd169} : s = 419;
	{8'd250,8'd170} : s = 420;
	{8'd250,8'd171} : s = 421;
	{8'd250,8'd172} : s = 422;
	{8'd250,8'd173} : s = 423;
	{8'd250,8'd174} : s = 424;
	{8'd250,8'd175} : s = 425;
	{8'd250,8'd176} : s = 426;
	{8'd250,8'd177} : s = 427;
	{8'd250,8'd178} : s = 428;
	{8'd250,8'd179} : s = 429;
	{8'd250,8'd180} : s = 430;
	{8'd250,8'd181} : s = 431;
	{8'd250,8'd182} : s = 432;
	{8'd250,8'd183} : s = 433;
	{8'd250,8'd184} : s = 434;
	{8'd250,8'd185} : s = 435;
	{8'd250,8'd186} : s = 436;
	{8'd250,8'd187} : s = 437;
	{8'd250,8'd188} : s = 438;
	{8'd250,8'd189} : s = 439;
	{8'd250,8'd190} : s = 440;
	{8'd250,8'd191} : s = 441;
	{8'd250,8'd192} : s = 442;
	{8'd250,8'd193} : s = 443;
	{8'd250,8'd194} : s = 444;
	{8'd250,8'd195} : s = 445;
	{8'd250,8'd196} : s = 446;
	{8'd250,8'd197} : s = 447;
	{8'd250,8'd198} : s = 448;
	{8'd250,8'd199} : s = 449;
	{8'd250,8'd200} : s = 450;
	{8'd250,8'd201} : s = 451;
	{8'd250,8'd202} : s = 452;
	{8'd250,8'd203} : s = 453;
	{8'd250,8'd204} : s = 454;
	{8'd250,8'd205} : s = 455;
	{8'd250,8'd206} : s = 456;
	{8'd250,8'd207} : s = 457;
	{8'd250,8'd208} : s = 458;
	{8'd250,8'd209} : s = 459;
	{8'd250,8'd210} : s = 460;
	{8'd250,8'd211} : s = 461;
	{8'd250,8'd212} : s = 462;
	{8'd250,8'd213} : s = 463;
	{8'd250,8'd214} : s = 464;
	{8'd250,8'd215} : s = 465;
	{8'd250,8'd216} : s = 466;
	{8'd250,8'd217} : s = 467;
	{8'd250,8'd218} : s = 468;
	{8'd250,8'd219} : s = 469;
	{8'd250,8'd220} : s = 470;
	{8'd250,8'd221} : s = 471;
	{8'd250,8'd222} : s = 472;
	{8'd250,8'd223} : s = 473;
	{8'd250,8'd224} : s = 474;
	{8'd250,8'd225} : s = 475;
	{8'd250,8'd226} : s = 476;
	{8'd250,8'd227} : s = 477;
	{8'd250,8'd228} : s = 478;
	{8'd250,8'd229} : s = 479;
	{8'd250,8'd230} : s = 480;
	{8'd250,8'd231} : s = 481;
	{8'd250,8'd232} : s = 482;
	{8'd250,8'd233} : s = 483;
	{8'd250,8'd234} : s = 484;
	{8'd250,8'd235} : s = 485;
	{8'd250,8'd236} : s = 486;
	{8'd250,8'd237} : s = 487;
	{8'd250,8'd238} : s = 488;
	{8'd250,8'd239} : s = 489;
	{8'd250,8'd240} : s = 490;
	{8'd250,8'd241} : s = 491;
	{8'd250,8'd242} : s = 492;
	{8'd250,8'd243} : s = 493;
	{8'd250,8'd244} : s = 494;
	{8'd250,8'd245} : s = 495;
	{8'd250,8'd246} : s = 496;
	{8'd250,8'd247} : s = 497;
	{8'd250,8'd248} : s = 498;
	{8'd250,8'd249} : s = 499;
	{8'd250,8'd250} : s = 500;
	{8'd250,8'd251} : s = 501;
	{8'd250,8'd252} : s = 502;
	{8'd250,8'd253} : s = 503;
	{8'd250,8'd254} : s = 504;
	{8'd250,8'd255} : s = 505;
	{8'd251,8'd0} : s = 251;
	{8'd251,8'd1} : s = 252;
	{8'd251,8'd2} : s = 253;
	{8'd251,8'd3} : s = 254;
	{8'd251,8'd4} : s = 255;
	{8'd251,8'd5} : s = 256;
	{8'd251,8'd6} : s = 257;
	{8'd251,8'd7} : s = 258;
	{8'd251,8'd8} : s = 259;
	{8'd251,8'd9} : s = 260;
	{8'd251,8'd10} : s = 261;
	{8'd251,8'd11} : s = 262;
	{8'd251,8'd12} : s = 263;
	{8'd251,8'd13} : s = 264;
	{8'd251,8'd14} : s = 265;
	{8'd251,8'd15} : s = 266;
	{8'd251,8'd16} : s = 267;
	{8'd251,8'd17} : s = 268;
	{8'd251,8'd18} : s = 269;
	{8'd251,8'd19} : s = 270;
	{8'd251,8'd20} : s = 271;
	{8'd251,8'd21} : s = 272;
	{8'd251,8'd22} : s = 273;
	{8'd251,8'd23} : s = 274;
	{8'd251,8'd24} : s = 275;
	{8'd251,8'd25} : s = 276;
	{8'd251,8'd26} : s = 277;
	{8'd251,8'd27} : s = 278;
	{8'd251,8'd28} : s = 279;
	{8'd251,8'd29} : s = 280;
	{8'd251,8'd30} : s = 281;
	{8'd251,8'd31} : s = 282;
	{8'd251,8'd32} : s = 283;
	{8'd251,8'd33} : s = 284;
	{8'd251,8'd34} : s = 285;
	{8'd251,8'd35} : s = 286;
	{8'd251,8'd36} : s = 287;
	{8'd251,8'd37} : s = 288;
	{8'd251,8'd38} : s = 289;
	{8'd251,8'd39} : s = 290;
	{8'd251,8'd40} : s = 291;
	{8'd251,8'd41} : s = 292;
	{8'd251,8'd42} : s = 293;
	{8'd251,8'd43} : s = 294;
	{8'd251,8'd44} : s = 295;
	{8'd251,8'd45} : s = 296;
	{8'd251,8'd46} : s = 297;
	{8'd251,8'd47} : s = 298;
	{8'd251,8'd48} : s = 299;
	{8'd251,8'd49} : s = 300;
	{8'd251,8'd50} : s = 301;
	{8'd251,8'd51} : s = 302;
	{8'd251,8'd52} : s = 303;
	{8'd251,8'd53} : s = 304;
	{8'd251,8'd54} : s = 305;
	{8'd251,8'd55} : s = 306;
	{8'd251,8'd56} : s = 307;
	{8'd251,8'd57} : s = 308;
	{8'd251,8'd58} : s = 309;
	{8'd251,8'd59} : s = 310;
	{8'd251,8'd60} : s = 311;
	{8'd251,8'd61} : s = 312;
	{8'd251,8'd62} : s = 313;
	{8'd251,8'd63} : s = 314;
	{8'd251,8'd64} : s = 315;
	{8'd251,8'd65} : s = 316;
	{8'd251,8'd66} : s = 317;
	{8'd251,8'd67} : s = 318;
	{8'd251,8'd68} : s = 319;
	{8'd251,8'd69} : s = 320;
	{8'd251,8'd70} : s = 321;
	{8'd251,8'd71} : s = 322;
	{8'd251,8'd72} : s = 323;
	{8'd251,8'd73} : s = 324;
	{8'd251,8'd74} : s = 325;
	{8'd251,8'd75} : s = 326;
	{8'd251,8'd76} : s = 327;
	{8'd251,8'd77} : s = 328;
	{8'd251,8'd78} : s = 329;
	{8'd251,8'd79} : s = 330;
	{8'd251,8'd80} : s = 331;
	{8'd251,8'd81} : s = 332;
	{8'd251,8'd82} : s = 333;
	{8'd251,8'd83} : s = 334;
	{8'd251,8'd84} : s = 335;
	{8'd251,8'd85} : s = 336;
	{8'd251,8'd86} : s = 337;
	{8'd251,8'd87} : s = 338;
	{8'd251,8'd88} : s = 339;
	{8'd251,8'd89} : s = 340;
	{8'd251,8'd90} : s = 341;
	{8'd251,8'd91} : s = 342;
	{8'd251,8'd92} : s = 343;
	{8'd251,8'd93} : s = 344;
	{8'd251,8'd94} : s = 345;
	{8'd251,8'd95} : s = 346;
	{8'd251,8'd96} : s = 347;
	{8'd251,8'd97} : s = 348;
	{8'd251,8'd98} : s = 349;
	{8'd251,8'd99} : s = 350;
	{8'd251,8'd100} : s = 351;
	{8'd251,8'd101} : s = 352;
	{8'd251,8'd102} : s = 353;
	{8'd251,8'd103} : s = 354;
	{8'd251,8'd104} : s = 355;
	{8'd251,8'd105} : s = 356;
	{8'd251,8'd106} : s = 357;
	{8'd251,8'd107} : s = 358;
	{8'd251,8'd108} : s = 359;
	{8'd251,8'd109} : s = 360;
	{8'd251,8'd110} : s = 361;
	{8'd251,8'd111} : s = 362;
	{8'd251,8'd112} : s = 363;
	{8'd251,8'd113} : s = 364;
	{8'd251,8'd114} : s = 365;
	{8'd251,8'd115} : s = 366;
	{8'd251,8'd116} : s = 367;
	{8'd251,8'd117} : s = 368;
	{8'd251,8'd118} : s = 369;
	{8'd251,8'd119} : s = 370;
	{8'd251,8'd120} : s = 371;
	{8'd251,8'd121} : s = 372;
	{8'd251,8'd122} : s = 373;
	{8'd251,8'd123} : s = 374;
	{8'd251,8'd124} : s = 375;
	{8'd251,8'd125} : s = 376;
	{8'd251,8'd126} : s = 377;
	{8'd251,8'd127} : s = 378;
	{8'd251,8'd128} : s = 379;
	{8'd251,8'd129} : s = 380;
	{8'd251,8'd130} : s = 381;
	{8'd251,8'd131} : s = 382;
	{8'd251,8'd132} : s = 383;
	{8'd251,8'd133} : s = 384;
	{8'd251,8'd134} : s = 385;
	{8'd251,8'd135} : s = 386;
	{8'd251,8'd136} : s = 387;
	{8'd251,8'd137} : s = 388;
	{8'd251,8'd138} : s = 389;
	{8'd251,8'd139} : s = 390;
	{8'd251,8'd140} : s = 391;
	{8'd251,8'd141} : s = 392;
	{8'd251,8'd142} : s = 393;
	{8'd251,8'd143} : s = 394;
	{8'd251,8'd144} : s = 395;
	{8'd251,8'd145} : s = 396;
	{8'd251,8'd146} : s = 397;
	{8'd251,8'd147} : s = 398;
	{8'd251,8'd148} : s = 399;
	{8'd251,8'd149} : s = 400;
	{8'd251,8'd150} : s = 401;
	{8'd251,8'd151} : s = 402;
	{8'd251,8'd152} : s = 403;
	{8'd251,8'd153} : s = 404;
	{8'd251,8'd154} : s = 405;
	{8'd251,8'd155} : s = 406;
	{8'd251,8'd156} : s = 407;
	{8'd251,8'd157} : s = 408;
	{8'd251,8'd158} : s = 409;
	{8'd251,8'd159} : s = 410;
	{8'd251,8'd160} : s = 411;
	{8'd251,8'd161} : s = 412;
	{8'd251,8'd162} : s = 413;
	{8'd251,8'd163} : s = 414;
	{8'd251,8'd164} : s = 415;
	{8'd251,8'd165} : s = 416;
	{8'd251,8'd166} : s = 417;
	{8'd251,8'd167} : s = 418;
	{8'd251,8'd168} : s = 419;
	{8'd251,8'd169} : s = 420;
	{8'd251,8'd170} : s = 421;
	{8'd251,8'd171} : s = 422;
	{8'd251,8'd172} : s = 423;
	{8'd251,8'd173} : s = 424;
	{8'd251,8'd174} : s = 425;
	{8'd251,8'd175} : s = 426;
	{8'd251,8'd176} : s = 427;
	{8'd251,8'd177} : s = 428;
	{8'd251,8'd178} : s = 429;
	{8'd251,8'd179} : s = 430;
	{8'd251,8'd180} : s = 431;
	{8'd251,8'd181} : s = 432;
	{8'd251,8'd182} : s = 433;
	{8'd251,8'd183} : s = 434;
	{8'd251,8'd184} : s = 435;
	{8'd251,8'd185} : s = 436;
	{8'd251,8'd186} : s = 437;
	{8'd251,8'd187} : s = 438;
	{8'd251,8'd188} : s = 439;
	{8'd251,8'd189} : s = 440;
	{8'd251,8'd190} : s = 441;
	{8'd251,8'd191} : s = 442;
	{8'd251,8'd192} : s = 443;
	{8'd251,8'd193} : s = 444;
	{8'd251,8'd194} : s = 445;
	{8'd251,8'd195} : s = 446;
	{8'd251,8'd196} : s = 447;
	{8'd251,8'd197} : s = 448;
	{8'd251,8'd198} : s = 449;
	{8'd251,8'd199} : s = 450;
	{8'd251,8'd200} : s = 451;
	{8'd251,8'd201} : s = 452;
	{8'd251,8'd202} : s = 453;
	{8'd251,8'd203} : s = 454;
	{8'd251,8'd204} : s = 455;
	{8'd251,8'd205} : s = 456;
	{8'd251,8'd206} : s = 457;
	{8'd251,8'd207} : s = 458;
	{8'd251,8'd208} : s = 459;
	{8'd251,8'd209} : s = 460;
	{8'd251,8'd210} : s = 461;
	{8'd251,8'd211} : s = 462;
	{8'd251,8'd212} : s = 463;
	{8'd251,8'd213} : s = 464;
	{8'd251,8'd214} : s = 465;
	{8'd251,8'd215} : s = 466;
	{8'd251,8'd216} : s = 467;
	{8'd251,8'd217} : s = 468;
	{8'd251,8'd218} : s = 469;
	{8'd251,8'd219} : s = 470;
	{8'd251,8'd220} : s = 471;
	{8'd251,8'd221} : s = 472;
	{8'd251,8'd222} : s = 473;
	{8'd251,8'd223} : s = 474;
	{8'd251,8'd224} : s = 475;
	{8'd251,8'd225} : s = 476;
	{8'd251,8'd226} : s = 477;
	{8'd251,8'd227} : s = 478;
	{8'd251,8'd228} : s = 479;
	{8'd251,8'd229} : s = 480;
	{8'd251,8'd230} : s = 481;
	{8'd251,8'd231} : s = 482;
	{8'd251,8'd232} : s = 483;
	{8'd251,8'd233} : s = 484;
	{8'd251,8'd234} : s = 485;
	{8'd251,8'd235} : s = 486;
	{8'd251,8'd236} : s = 487;
	{8'd251,8'd237} : s = 488;
	{8'd251,8'd238} : s = 489;
	{8'd251,8'd239} : s = 490;
	{8'd251,8'd240} : s = 491;
	{8'd251,8'd241} : s = 492;
	{8'd251,8'd242} : s = 493;
	{8'd251,8'd243} : s = 494;
	{8'd251,8'd244} : s = 495;
	{8'd251,8'd245} : s = 496;
	{8'd251,8'd246} : s = 497;
	{8'd251,8'd247} : s = 498;
	{8'd251,8'd248} : s = 499;
	{8'd251,8'd249} : s = 500;
	{8'd251,8'd250} : s = 501;
	{8'd251,8'd251} : s = 502;
	{8'd251,8'd252} : s = 503;
	{8'd251,8'd253} : s = 504;
	{8'd251,8'd254} : s = 505;
	{8'd251,8'd255} : s = 506;
	{8'd252,8'd0} : s = 252;
	{8'd252,8'd1} : s = 253;
	{8'd252,8'd2} : s = 254;
	{8'd252,8'd3} : s = 255;
	{8'd252,8'd4} : s = 256;
	{8'd252,8'd5} : s = 257;
	{8'd252,8'd6} : s = 258;
	{8'd252,8'd7} : s = 259;
	{8'd252,8'd8} : s = 260;
	{8'd252,8'd9} : s = 261;
	{8'd252,8'd10} : s = 262;
	{8'd252,8'd11} : s = 263;
	{8'd252,8'd12} : s = 264;
	{8'd252,8'd13} : s = 265;
	{8'd252,8'd14} : s = 266;
	{8'd252,8'd15} : s = 267;
	{8'd252,8'd16} : s = 268;
	{8'd252,8'd17} : s = 269;
	{8'd252,8'd18} : s = 270;
	{8'd252,8'd19} : s = 271;
	{8'd252,8'd20} : s = 272;
	{8'd252,8'd21} : s = 273;
	{8'd252,8'd22} : s = 274;
	{8'd252,8'd23} : s = 275;
	{8'd252,8'd24} : s = 276;
	{8'd252,8'd25} : s = 277;
	{8'd252,8'd26} : s = 278;
	{8'd252,8'd27} : s = 279;
	{8'd252,8'd28} : s = 280;
	{8'd252,8'd29} : s = 281;
	{8'd252,8'd30} : s = 282;
	{8'd252,8'd31} : s = 283;
	{8'd252,8'd32} : s = 284;
	{8'd252,8'd33} : s = 285;
	{8'd252,8'd34} : s = 286;
	{8'd252,8'd35} : s = 287;
	{8'd252,8'd36} : s = 288;
	{8'd252,8'd37} : s = 289;
	{8'd252,8'd38} : s = 290;
	{8'd252,8'd39} : s = 291;
	{8'd252,8'd40} : s = 292;
	{8'd252,8'd41} : s = 293;
	{8'd252,8'd42} : s = 294;
	{8'd252,8'd43} : s = 295;
	{8'd252,8'd44} : s = 296;
	{8'd252,8'd45} : s = 297;
	{8'd252,8'd46} : s = 298;
	{8'd252,8'd47} : s = 299;
	{8'd252,8'd48} : s = 300;
	{8'd252,8'd49} : s = 301;
	{8'd252,8'd50} : s = 302;
	{8'd252,8'd51} : s = 303;
	{8'd252,8'd52} : s = 304;
	{8'd252,8'd53} : s = 305;
	{8'd252,8'd54} : s = 306;
	{8'd252,8'd55} : s = 307;
	{8'd252,8'd56} : s = 308;
	{8'd252,8'd57} : s = 309;
	{8'd252,8'd58} : s = 310;
	{8'd252,8'd59} : s = 311;
	{8'd252,8'd60} : s = 312;
	{8'd252,8'd61} : s = 313;
	{8'd252,8'd62} : s = 314;
	{8'd252,8'd63} : s = 315;
	{8'd252,8'd64} : s = 316;
	{8'd252,8'd65} : s = 317;
	{8'd252,8'd66} : s = 318;
	{8'd252,8'd67} : s = 319;
	{8'd252,8'd68} : s = 320;
	{8'd252,8'd69} : s = 321;
	{8'd252,8'd70} : s = 322;
	{8'd252,8'd71} : s = 323;
	{8'd252,8'd72} : s = 324;
	{8'd252,8'd73} : s = 325;
	{8'd252,8'd74} : s = 326;
	{8'd252,8'd75} : s = 327;
	{8'd252,8'd76} : s = 328;
	{8'd252,8'd77} : s = 329;
	{8'd252,8'd78} : s = 330;
	{8'd252,8'd79} : s = 331;
	{8'd252,8'd80} : s = 332;
	{8'd252,8'd81} : s = 333;
	{8'd252,8'd82} : s = 334;
	{8'd252,8'd83} : s = 335;
	{8'd252,8'd84} : s = 336;
	{8'd252,8'd85} : s = 337;
	{8'd252,8'd86} : s = 338;
	{8'd252,8'd87} : s = 339;
	{8'd252,8'd88} : s = 340;
	{8'd252,8'd89} : s = 341;
	{8'd252,8'd90} : s = 342;
	{8'd252,8'd91} : s = 343;
	{8'd252,8'd92} : s = 344;
	{8'd252,8'd93} : s = 345;
	{8'd252,8'd94} : s = 346;
	{8'd252,8'd95} : s = 347;
	{8'd252,8'd96} : s = 348;
	{8'd252,8'd97} : s = 349;
	{8'd252,8'd98} : s = 350;
	{8'd252,8'd99} : s = 351;
	{8'd252,8'd100} : s = 352;
	{8'd252,8'd101} : s = 353;
	{8'd252,8'd102} : s = 354;
	{8'd252,8'd103} : s = 355;
	{8'd252,8'd104} : s = 356;
	{8'd252,8'd105} : s = 357;
	{8'd252,8'd106} : s = 358;
	{8'd252,8'd107} : s = 359;
	{8'd252,8'd108} : s = 360;
	{8'd252,8'd109} : s = 361;
	{8'd252,8'd110} : s = 362;
	{8'd252,8'd111} : s = 363;
	{8'd252,8'd112} : s = 364;
	{8'd252,8'd113} : s = 365;
	{8'd252,8'd114} : s = 366;
	{8'd252,8'd115} : s = 367;
	{8'd252,8'd116} : s = 368;
	{8'd252,8'd117} : s = 369;
	{8'd252,8'd118} : s = 370;
	{8'd252,8'd119} : s = 371;
	{8'd252,8'd120} : s = 372;
	{8'd252,8'd121} : s = 373;
	{8'd252,8'd122} : s = 374;
	{8'd252,8'd123} : s = 375;
	{8'd252,8'd124} : s = 376;
	{8'd252,8'd125} : s = 377;
	{8'd252,8'd126} : s = 378;
	{8'd252,8'd127} : s = 379;
	{8'd252,8'd128} : s = 380;
	{8'd252,8'd129} : s = 381;
	{8'd252,8'd130} : s = 382;
	{8'd252,8'd131} : s = 383;
	{8'd252,8'd132} : s = 384;
	{8'd252,8'd133} : s = 385;
	{8'd252,8'd134} : s = 386;
	{8'd252,8'd135} : s = 387;
	{8'd252,8'd136} : s = 388;
	{8'd252,8'd137} : s = 389;
	{8'd252,8'd138} : s = 390;
	{8'd252,8'd139} : s = 391;
	{8'd252,8'd140} : s = 392;
	{8'd252,8'd141} : s = 393;
	{8'd252,8'd142} : s = 394;
	{8'd252,8'd143} : s = 395;
	{8'd252,8'd144} : s = 396;
	{8'd252,8'd145} : s = 397;
	{8'd252,8'd146} : s = 398;
	{8'd252,8'd147} : s = 399;
	{8'd252,8'd148} : s = 400;
	{8'd252,8'd149} : s = 401;
	{8'd252,8'd150} : s = 402;
	{8'd252,8'd151} : s = 403;
	{8'd252,8'd152} : s = 404;
	{8'd252,8'd153} : s = 405;
	{8'd252,8'd154} : s = 406;
	{8'd252,8'd155} : s = 407;
	{8'd252,8'd156} : s = 408;
	{8'd252,8'd157} : s = 409;
	{8'd252,8'd158} : s = 410;
	{8'd252,8'd159} : s = 411;
	{8'd252,8'd160} : s = 412;
	{8'd252,8'd161} : s = 413;
	{8'd252,8'd162} : s = 414;
	{8'd252,8'd163} : s = 415;
	{8'd252,8'd164} : s = 416;
	{8'd252,8'd165} : s = 417;
	{8'd252,8'd166} : s = 418;
	{8'd252,8'd167} : s = 419;
	{8'd252,8'd168} : s = 420;
	{8'd252,8'd169} : s = 421;
	{8'd252,8'd170} : s = 422;
	{8'd252,8'd171} : s = 423;
	{8'd252,8'd172} : s = 424;
	{8'd252,8'd173} : s = 425;
	{8'd252,8'd174} : s = 426;
	{8'd252,8'd175} : s = 427;
	{8'd252,8'd176} : s = 428;
	{8'd252,8'd177} : s = 429;
	{8'd252,8'd178} : s = 430;
	{8'd252,8'd179} : s = 431;
	{8'd252,8'd180} : s = 432;
	{8'd252,8'd181} : s = 433;
	{8'd252,8'd182} : s = 434;
	{8'd252,8'd183} : s = 435;
	{8'd252,8'd184} : s = 436;
	{8'd252,8'd185} : s = 437;
	{8'd252,8'd186} : s = 438;
	{8'd252,8'd187} : s = 439;
	{8'd252,8'd188} : s = 440;
	{8'd252,8'd189} : s = 441;
	{8'd252,8'd190} : s = 442;
	{8'd252,8'd191} : s = 443;
	{8'd252,8'd192} : s = 444;
	{8'd252,8'd193} : s = 445;
	{8'd252,8'd194} : s = 446;
	{8'd252,8'd195} : s = 447;
	{8'd252,8'd196} : s = 448;
	{8'd252,8'd197} : s = 449;
	{8'd252,8'd198} : s = 450;
	{8'd252,8'd199} : s = 451;
	{8'd252,8'd200} : s = 452;
	{8'd252,8'd201} : s = 453;
	{8'd252,8'd202} : s = 454;
	{8'd252,8'd203} : s = 455;
	{8'd252,8'd204} : s = 456;
	{8'd252,8'd205} : s = 457;
	{8'd252,8'd206} : s = 458;
	{8'd252,8'd207} : s = 459;
	{8'd252,8'd208} : s = 460;
	{8'd252,8'd209} : s = 461;
	{8'd252,8'd210} : s = 462;
	{8'd252,8'd211} : s = 463;
	{8'd252,8'd212} : s = 464;
	{8'd252,8'd213} : s = 465;
	{8'd252,8'd214} : s = 466;
	{8'd252,8'd215} : s = 467;
	{8'd252,8'd216} : s = 468;
	{8'd252,8'd217} : s = 469;
	{8'd252,8'd218} : s = 470;
	{8'd252,8'd219} : s = 471;
	{8'd252,8'd220} : s = 472;
	{8'd252,8'd221} : s = 473;
	{8'd252,8'd222} : s = 474;
	{8'd252,8'd223} : s = 475;
	{8'd252,8'd224} : s = 476;
	{8'd252,8'd225} : s = 477;
	{8'd252,8'd226} : s = 478;
	{8'd252,8'd227} : s = 479;
	{8'd252,8'd228} : s = 480;
	{8'd252,8'd229} : s = 481;
	{8'd252,8'd230} : s = 482;
	{8'd252,8'd231} : s = 483;
	{8'd252,8'd232} : s = 484;
	{8'd252,8'd233} : s = 485;
	{8'd252,8'd234} : s = 486;
	{8'd252,8'd235} : s = 487;
	{8'd252,8'd236} : s = 488;
	{8'd252,8'd237} : s = 489;
	{8'd252,8'd238} : s = 490;
	{8'd252,8'd239} : s = 491;
	{8'd252,8'd240} : s = 492;
	{8'd252,8'd241} : s = 493;
	{8'd252,8'd242} : s = 494;
	{8'd252,8'd243} : s = 495;
	{8'd252,8'd244} : s = 496;
	{8'd252,8'd245} : s = 497;
	{8'd252,8'd246} : s = 498;
	{8'd252,8'd247} : s = 499;
	{8'd252,8'd248} : s = 500;
	{8'd252,8'd249} : s = 501;
	{8'd252,8'd250} : s = 502;
	{8'd252,8'd251} : s = 503;
	{8'd252,8'd252} : s = 504;
	{8'd252,8'd253} : s = 505;
	{8'd252,8'd254} : s = 506;
	{8'd252,8'd255} : s = 507;
	{8'd253,8'd0} : s = 253;
	{8'd253,8'd1} : s = 254;
	{8'd253,8'd2} : s = 255;
	{8'd253,8'd3} : s = 256;
	{8'd253,8'd4} : s = 257;
	{8'd253,8'd5} : s = 258;
	{8'd253,8'd6} : s = 259;
	{8'd253,8'd7} : s = 260;
	{8'd253,8'd8} : s = 261;
	{8'd253,8'd9} : s = 262;
	{8'd253,8'd10} : s = 263;
	{8'd253,8'd11} : s = 264;
	{8'd253,8'd12} : s = 265;
	{8'd253,8'd13} : s = 266;
	{8'd253,8'd14} : s = 267;
	{8'd253,8'd15} : s = 268;
	{8'd253,8'd16} : s = 269;
	{8'd253,8'd17} : s = 270;
	{8'd253,8'd18} : s = 271;
	{8'd253,8'd19} : s = 272;
	{8'd253,8'd20} : s = 273;
	{8'd253,8'd21} : s = 274;
	{8'd253,8'd22} : s = 275;
	{8'd253,8'd23} : s = 276;
	{8'd253,8'd24} : s = 277;
	{8'd253,8'd25} : s = 278;
	{8'd253,8'd26} : s = 279;
	{8'd253,8'd27} : s = 280;
	{8'd253,8'd28} : s = 281;
	{8'd253,8'd29} : s = 282;
	{8'd253,8'd30} : s = 283;
	{8'd253,8'd31} : s = 284;
	{8'd253,8'd32} : s = 285;
	{8'd253,8'd33} : s = 286;
	{8'd253,8'd34} : s = 287;
	{8'd253,8'd35} : s = 288;
	{8'd253,8'd36} : s = 289;
	{8'd253,8'd37} : s = 290;
	{8'd253,8'd38} : s = 291;
	{8'd253,8'd39} : s = 292;
	{8'd253,8'd40} : s = 293;
	{8'd253,8'd41} : s = 294;
	{8'd253,8'd42} : s = 295;
	{8'd253,8'd43} : s = 296;
	{8'd253,8'd44} : s = 297;
	{8'd253,8'd45} : s = 298;
	{8'd253,8'd46} : s = 299;
	{8'd253,8'd47} : s = 300;
	{8'd253,8'd48} : s = 301;
	{8'd253,8'd49} : s = 302;
	{8'd253,8'd50} : s = 303;
	{8'd253,8'd51} : s = 304;
	{8'd253,8'd52} : s = 305;
	{8'd253,8'd53} : s = 306;
	{8'd253,8'd54} : s = 307;
	{8'd253,8'd55} : s = 308;
	{8'd253,8'd56} : s = 309;
	{8'd253,8'd57} : s = 310;
	{8'd253,8'd58} : s = 311;
	{8'd253,8'd59} : s = 312;
	{8'd253,8'd60} : s = 313;
	{8'd253,8'd61} : s = 314;
	{8'd253,8'd62} : s = 315;
	{8'd253,8'd63} : s = 316;
	{8'd253,8'd64} : s = 317;
	{8'd253,8'd65} : s = 318;
	{8'd253,8'd66} : s = 319;
	{8'd253,8'd67} : s = 320;
	{8'd253,8'd68} : s = 321;
	{8'd253,8'd69} : s = 322;
	{8'd253,8'd70} : s = 323;
	{8'd253,8'd71} : s = 324;
	{8'd253,8'd72} : s = 325;
	{8'd253,8'd73} : s = 326;
	{8'd253,8'd74} : s = 327;
	{8'd253,8'd75} : s = 328;
	{8'd253,8'd76} : s = 329;
	{8'd253,8'd77} : s = 330;
	{8'd253,8'd78} : s = 331;
	{8'd253,8'd79} : s = 332;
	{8'd253,8'd80} : s = 333;
	{8'd253,8'd81} : s = 334;
	{8'd253,8'd82} : s = 335;
	{8'd253,8'd83} : s = 336;
	{8'd253,8'd84} : s = 337;
	{8'd253,8'd85} : s = 338;
	{8'd253,8'd86} : s = 339;
	{8'd253,8'd87} : s = 340;
	{8'd253,8'd88} : s = 341;
	{8'd253,8'd89} : s = 342;
	{8'd253,8'd90} : s = 343;
	{8'd253,8'd91} : s = 344;
	{8'd253,8'd92} : s = 345;
	{8'd253,8'd93} : s = 346;
	{8'd253,8'd94} : s = 347;
	{8'd253,8'd95} : s = 348;
	{8'd253,8'd96} : s = 349;
	{8'd253,8'd97} : s = 350;
	{8'd253,8'd98} : s = 351;
	{8'd253,8'd99} : s = 352;
	{8'd253,8'd100} : s = 353;
	{8'd253,8'd101} : s = 354;
	{8'd253,8'd102} : s = 355;
	{8'd253,8'd103} : s = 356;
	{8'd253,8'd104} : s = 357;
	{8'd253,8'd105} : s = 358;
	{8'd253,8'd106} : s = 359;
	{8'd253,8'd107} : s = 360;
	{8'd253,8'd108} : s = 361;
	{8'd253,8'd109} : s = 362;
	{8'd253,8'd110} : s = 363;
	{8'd253,8'd111} : s = 364;
	{8'd253,8'd112} : s = 365;
	{8'd253,8'd113} : s = 366;
	{8'd253,8'd114} : s = 367;
	{8'd253,8'd115} : s = 368;
	{8'd253,8'd116} : s = 369;
	{8'd253,8'd117} : s = 370;
	{8'd253,8'd118} : s = 371;
	{8'd253,8'd119} : s = 372;
	{8'd253,8'd120} : s = 373;
	{8'd253,8'd121} : s = 374;
	{8'd253,8'd122} : s = 375;
	{8'd253,8'd123} : s = 376;
	{8'd253,8'd124} : s = 377;
	{8'd253,8'd125} : s = 378;
	{8'd253,8'd126} : s = 379;
	{8'd253,8'd127} : s = 380;
	{8'd253,8'd128} : s = 381;
	{8'd253,8'd129} : s = 382;
	{8'd253,8'd130} : s = 383;
	{8'd253,8'd131} : s = 384;
	{8'd253,8'd132} : s = 385;
	{8'd253,8'd133} : s = 386;
	{8'd253,8'd134} : s = 387;
	{8'd253,8'd135} : s = 388;
	{8'd253,8'd136} : s = 389;
	{8'd253,8'd137} : s = 390;
	{8'd253,8'd138} : s = 391;
	{8'd253,8'd139} : s = 392;
	{8'd253,8'd140} : s = 393;
	{8'd253,8'd141} : s = 394;
	{8'd253,8'd142} : s = 395;
	{8'd253,8'd143} : s = 396;
	{8'd253,8'd144} : s = 397;
	{8'd253,8'd145} : s = 398;
	{8'd253,8'd146} : s = 399;
	{8'd253,8'd147} : s = 400;
	{8'd253,8'd148} : s = 401;
	{8'd253,8'd149} : s = 402;
	{8'd253,8'd150} : s = 403;
	{8'd253,8'd151} : s = 404;
	{8'd253,8'd152} : s = 405;
	{8'd253,8'd153} : s = 406;
	{8'd253,8'd154} : s = 407;
	{8'd253,8'd155} : s = 408;
	{8'd253,8'd156} : s = 409;
	{8'd253,8'd157} : s = 410;
	{8'd253,8'd158} : s = 411;
	{8'd253,8'd159} : s = 412;
	{8'd253,8'd160} : s = 413;
	{8'd253,8'd161} : s = 414;
	{8'd253,8'd162} : s = 415;
	{8'd253,8'd163} : s = 416;
	{8'd253,8'd164} : s = 417;
	{8'd253,8'd165} : s = 418;
	{8'd253,8'd166} : s = 419;
	{8'd253,8'd167} : s = 420;
	{8'd253,8'd168} : s = 421;
	{8'd253,8'd169} : s = 422;
	{8'd253,8'd170} : s = 423;
	{8'd253,8'd171} : s = 424;
	{8'd253,8'd172} : s = 425;
	{8'd253,8'd173} : s = 426;
	{8'd253,8'd174} : s = 427;
	{8'd253,8'd175} : s = 428;
	{8'd253,8'd176} : s = 429;
	{8'd253,8'd177} : s = 430;
	{8'd253,8'd178} : s = 431;
	{8'd253,8'd179} : s = 432;
	{8'd253,8'd180} : s = 433;
	{8'd253,8'd181} : s = 434;
	{8'd253,8'd182} : s = 435;
	{8'd253,8'd183} : s = 436;
	{8'd253,8'd184} : s = 437;
	{8'd253,8'd185} : s = 438;
	{8'd253,8'd186} : s = 439;
	{8'd253,8'd187} : s = 440;
	{8'd253,8'd188} : s = 441;
	{8'd253,8'd189} : s = 442;
	{8'd253,8'd190} : s = 443;
	{8'd253,8'd191} : s = 444;
	{8'd253,8'd192} : s = 445;
	{8'd253,8'd193} : s = 446;
	{8'd253,8'd194} : s = 447;
	{8'd253,8'd195} : s = 448;
	{8'd253,8'd196} : s = 449;
	{8'd253,8'd197} : s = 450;
	{8'd253,8'd198} : s = 451;
	{8'd253,8'd199} : s = 452;
	{8'd253,8'd200} : s = 453;
	{8'd253,8'd201} : s = 454;
	{8'd253,8'd202} : s = 455;
	{8'd253,8'd203} : s = 456;
	{8'd253,8'd204} : s = 457;
	{8'd253,8'd205} : s = 458;
	{8'd253,8'd206} : s = 459;
	{8'd253,8'd207} : s = 460;
	{8'd253,8'd208} : s = 461;
	{8'd253,8'd209} : s = 462;
	{8'd253,8'd210} : s = 463;
	{8'd253,8'd211} : s = 464;
	{8'd253,8'd212} : s = 465;
	{8'd253,8'd213} : s = 466;
	{8'd253,8'd214} : s = 467;
	{8'd253,8'd215} : s = 468;
	{8'd253,8'd216} : s = 469;
	{8'd253,8'd217} : s = 470;
	{8'd253,8'd218} : s = 471;
	{8'd253,8'd219} : s = 472;
	{8'd253,8'd220} : s = 473;
	{8'd253,8'd221} : s = 474;
	{8'd253,8'd222} : s = 475;
	{8'd253,8'd223} : s = 476;
	{8'd253,8'd224} : s = 477;
	{8'd253,8'd225} : s = 478;
	{8'd253,8'd226} : s = 479;
	{8'd253,8'd227} : s = 480;
	{8'd253,8'd228} : s = 481;
	{8'd253,8'd229} : s = 482;
	{8'd253,8'd230} : s = 483;
	{8'd253,8'd231} : s = 484;
	{8'd253,8'd232} : s = 485;
	{8'd253,8'd233} : s = 486;
	{8'd253,8'd234} : s = 487;
	{8'd253,8'd235} : s = 488;
	{8'd253,8'd236} : s = 489;
	{8'd253,8'd237} : s = 490;
	{8'd253,8'd238} : s = 491;
	{8'd253,8'd239} : s = 492;
	{8'd253,8'd240} : s = 493;
	{8'd253,8'd241} : s = 494;
	{8'd253,8'd242} : s = 495;
	{8'd253,8'd243} : s = 496;
	{8'd253,8'd244} : s = 497;
	{8'd253,8'd245} : s = 498;
	{8'd253,8'd246} : s = 499;
	{8'd253,8'd247} : s = 500;
	{8'd253,8'd248} : s = 501;
	{8'd253,8'd249} : s = 502;
	{8'd253,8'd250} : s = 503;
	{8'd253,8'd251} : s = 504;
	{8'd253,8'd252} : s = 505;
	{8'd253,8'd253} : s = 506;
	{8'd253,8'd254} : s = 507;
	{8'd253,8'd255} : s = 508;
	{8'd254,8'd0} : s = 254;
	{8'd254,8'd1} : s = 255;
	{8'd254,8'd2} : s = 256;
	{8'd254,8'd3} : s = 257;
	{8'd254,8'd4} : s = 258;
	{8'd254,8'd5} : s = 259;
	{8'd254,8'd6} : s = 260;
	{8'd254,8'd7} : s = 261;
	{8'd254,8'd8} : s = 262;
	{8'd254,8'd9} : s = 263;
	{8'd254,8'd10} : s = 264;
	{8'd254,8'd11} : s = 265;
	{8'd254,8'd12} : s = 266;
	{8'd254,8'd13} : s = 267;
	{8'd254,8'd14} : s = 268;
	{8'd254,8'd15} : s = 269;
	{8'd254,8'd16} : s = 270;
	{8'd254,8'd17} : s = 271;
	{8'd254,8'd18} : s = 272;
	{8'd254,8'd19} : s = 273;
	{8'd254,8'd20} : s = 274;
	{8'd254,8'd21} : s = 275;
	{8'd254,8'd22} : s = 276;
	{8'd254,8'd23} : s = 277;
	{8'd254,8'd24} : s = 278;
	{8'd254,8'd25} : s = 279;
	{8'd254,8'd26} : s = 280;
	{8'd254,8'd27} : s = 281;
	{8'd254,8'd28} : s = 282;
	{8'd254,8'd29} : s = 283;
	{8'd254,8'd30} : s = 284;
	{8'd254,8'd31} : s = 285;
	{8'd254,8'd32} : s = 286;
	{8'd254,8'd33} : s = 287;
	{8'd254,8'd34} : s = 288;
	{8'd254,8'd35} : s = 289;
	{8'd254,8'd36} : s = 290;
	{8'd254,8'd37} : s = 291;
	{8'd254,8'd38} : s = 292;
	{8'd254,8'd39} : s = 293;
	{8'd254,8'd40} : s = 294;
	{8'd254,8'd41} : s = 295;
	{8'd254,8'd42} : s = 296;
	{8'd254,8'd43} : s = 297;
	{8'd254,8'd44} : s = 298;
	{8'd254,8'd45} : s = 299;
	{8'd254,8'd46} : s = 300;
	{8'd254,8'd47} : s = 301;
	{8'd254,8'd48} : s = 302;
	{8'd254,8'd49} : s = 303;
	{8'd254,8'd50} : s = 304;
	{8'd254,8'd51} : s = 305;
	{8'd254,8'd52} : s = 306;
	{8'd254,8'd53} : s = 307;
	{8'd254,8'd54} : s = 308;
	{8'd254,8'd55} : s = 309;
	{8'd254,8'd56} : s = 310;
	{8'd254,8'd57} : s = 311;
	{8'd254,8'd58} : s = 312;
	{8'd254,8'd59} : s = 313;
	{8'd254,8'd60} : s = 314;
	{8'd254,8'd61} : s = 315;
	{8'd254,8'd62} : s = 316;
	{8'd254,8'd63} : s = 317;
	{8'd254,8'd64} : s = 318;
	{8'd254,8'd65} : s = 319;
	{8'd254,8'd66} : s = 320;
	{8'd254,8'd67} : s = 321;
	{8'd254,8'd68} : s = 322;
	{8'd254,8'd69} : s = 323;
	{8'd254,8'd70} : s = 324;
	{8'd254,8'd71} : s = 325;
	{8'd254,8'd72} : s = 326;
	{8'd254,8'd73} : s = 327;
	{8'd254,8'd74} : s = 328;
	{8'd254,8'd75} : s = 329;
	{8'd254,8'd76} : s = 330;
	{8'd254,8'd77} : s = 331;
	{8'd254,8'd78} : s = 332;
	{8'd254,8'd79} : s = 333;
	{8'd254,8'd80} : s = 334;
	{8'd254,8'd81} : s = 335;
	{8'd254,8'd82} : s = 336;
	{8'd254,8'd83} : s = 337;
	{8'd254,8'd84} : s = 338;
	{8'd254,8'd85} : s = 339;
	{8'd254,8'd86} : s = 340;
	{8'd254,8'd87} : s = 341;
	{8'd254,8'd88} : s = 342;
	{8'd254,8'd89} : s = 343;
	{8'd254,8'd90} : s = 344;
	{8'd254,8'd91} : s = 345;
	{8'd254,8'd92} : s = 346;
	{8'd254,8'd93} : s = 347;
	{8'd254,8'd94} : s = 348;
	{8'd254,8'd95} : s = 349;
	{8'd254,8'd96} : s = 350;
	{8'd254,8'd97} : s = 351;
	{8'd254,8'd98} : s = 352;
	{8'd254,8'd99} : s = 353;
	{8'd254,8'd100} : s = 354;
	{8'd254,8'd101} : s = 355;
	{8'd254,8'd102} : s = 356;
	{8'd254,8'd103} : s = 357;
	{8'd254,8'd104} : s = 358;
	{8'd254,8'd105} : s = 359;
	{8'd254,8'd106} : s = 360;
	{8'd254,8'd107} : s = 361;
	{8'd254,8'd108} : s = 362;
	{8'd254,8'd109} : s = 363;
	{8'd254,8'd110} : s = 364;
	{8'd254,8'd111} : s = 365;
	{8'd254,8'd112} : s = 366;
	{8'd254,8'd113} : s = 367;
	{8'd254,8'd114} : s = 368;
	{8'd254,8'd115} : s = 369;
	{8'd254,8'd116} : s = 370;
	{8'd254,8'd117} : s = 371;
	{8'd254,8'd118} : s = 372;
	{8'd254,8'd119} : s = 373;
	{8'd254,8'd120} : s = 374;
	{8'd254,8'd121} : s = 375;
	{8'd254,8'd122} : s = 376;
	{8'd254,8'd123} : s = 377;
	{8'd254,8'd124} : s = 378;
	{8'd254,8'd125} : s = 379;
	{8'd254,8'd126} : s = 380;
	{8'd254,8'd127} : s = 381;
	{8'd254,8'd128} : s = 382;
	{8'd254,8'd129} : s = 383;
	{8'd254,8'd130} : s = 384;
	{8'd254,8'd131} : s = 385;
	{8'd254,8'd132} : s = 386;
	{8'd254,8'd133} : s = 387;
	{8'd254,8'd134} : s = 388;
	{8'd254,8'd135} : s = 389;
	{8'd254,8'd136} : s = 390;
	{8'd254,8'd137} : s = 391;
	{8'd254,8'd138} : s = 392;
	{8'd254,8'd139} : s = 393;
	{8'd254,8'd140} : s = 394;
	{8'd254,8'd141} : s = 395;
	{8'd254,8'd142} : s = 396;
	{8'd254,8'd143} : s = 397;
	{8'd254,8'd144} : s = 398;
	{8'd254,8'd145} : s = 399;
	{8'd254,8'd146} : s = 400;
	{8'd254,8'd147} : s = 401;
	{8'd254,8'd148} : s = 402;
	{8'd254,8'd149} : s = 403;
	{8'd254,8'd150} : s = 404;
	{8'd254,8'd151} : s = 405;
	{8'd254,8'd152} : s = 406;
	{8'd254,8'd153} : s = 407;
	{8'd254,8'd154} : s = 408;
	{8'd254,8'd155} : s = 409;
	{8'd254,8'd156} : s = 410;
	{8'd254,8'd157} : s = 411;
	{8'd254,8'd158} : s = 412;
	{8'd254,8'd159} : s = 413;
	{8'd254,8'd160} : s = 414;
	{8'd254,8'd161} : s = 415;
	{8'd254,8'd162} : s = 416;
	{8'd254,8'd163} : s = 417;
	{8'd254,8'd164} : s = 418;
	{8'd254,8'd165} : s = 419;
	{8'd254,8'd166} : s = 420;
	{8'd254,8'd167} : s = 421;
	{8'd254,8'd168} : s = 422;
	{8'd254,8'd169} : s = 423;
	{8'd254,8'd170} : s = 424;
	{8'd254,8'd171} : s = 425;
	{8'd254,8'd172} : s = 426;
	{8'd254,8'd173} : s = 427;
	{8'd254,8'd174} : s = 428;
	{8'd254,8'd175} : s = 429;
	{8'd254,8'd176} : s = 430;
	{8'd254,8'd177} : s = 431;
	{8'd254,8'd178} : s = 432;
	{8'd254,8'd179} : s = 433;
	{8'd254,8'd180} : s = 434;
	{8'd254,8'd181} : s = 435;
	{8'd254,8'd182} : s = 436;
	{8'd254,8'd183} : s = 437;
	{8'd254,8'd184} : s = 438;
	{8'd254,8'd185} : s = 439;
	{8'd254,8'd186} : s = 440;
	{8'd254,8'd187} : s = 441;
	{8'd254,8'd188} : s = 442;
	{8'd254,8'd189} : s = 443;
	{8'd254,8'd190} : s = 444;
	{8'd254,8'd191} : s = 445;
	{8'd254,8'd192} : s = 446;
	{8'd254,8'd193} : s = 447;
	{8'd254,8'd194} : s = 448;
	{8'd254,8'd195} : s = 449;
	{8'd254,8'd196} : s = 450;
	{8'd254,8'd197} : s = 451;
	{8'd254,8'd198} : s = 452;
	{8'd254,8'd199} : s = 453;
	{8'd254,8'd200} : s = 454;
	{8'd254,8'd201} : s = 455;
	{8'd254,8'd202} : s = 456;
	{8'd254,8'd203} : s = 457;
	{8'd254,8'd204} : s = 458;
	{8'd254,8'd205} : s = 459;
	{8'd254,8'd206} : s = 460;
	{8'd254,8'd207} : s = 461;
	{8'd254,8'd208} : s = 462;
	{8'd254,8'd209} : s = 463;
	{8'd254,8'd210} : s = 464;
	{8'd254,8'd211} : s = 465;
	{8'd254,8'd212} : s = 466;
	{8'd254,8'd213} : s = 467;
	{8'd254,8'd214} : s = 468;
	{8'd254,8'd215} : s = 469;
	{8'd254,8'd216} : s = 470;
	{8'd254,8'd217} : s = 471;
	{8'd254,8'd218} : s = 472;
	{8'd254,8'd219} : s = 473;
	{8'd254,8'd220} : s = 474;
	{8'd254,8'd221} : s = 475;
	{8'd254,8'd222} : s = 476;
	{8'd254,8'd223} : s = 477;
	{8'd254,8'd224} : s = 478;
	{8'd254,8'd225} : s = 479;
	{8'd254,8'd226} : s = 480;
	{8'd254,8'd227} : s = 481;
	{8'd254,8'd228} : s = 482;
	{8'd254,8'd229} : s = 483;
	{8'd254,8'd230} : s = 484;
	{8'd254,8'd231} : s = 485;
	{8'd254,8'd232} : s = 486;
	{8'd254,8'd233} : s = 487;
	{8'd254,8'd234} : s = 488;
	{8'd254,8'd235} : s = 489;
	{8'd254,8'd236} : s = 490;
	{8'd254,8'd237} : s = 491;
	{8'd254,8'd238} : s = 492;
	{8'd254,8'd239} : s = 493;
	{8'd254,8'd240} : s = 494;
	{8'd254,8'd241} : s = 495;
	{8'd254,8'd242} : s = 496;
	{8'd254,8'd243} : s = 497;
	{8'd254,8'd244} : s = 498;
	{8'd254,8'd245} : s = 499;
	{8'd254,8'd246} : s = 500;
	{8'd254,8'd247} : s = 501;
	{8'd254,8'd248} : s = 502;
	{8'd254,8'd249} : s = 503;
	{8'd254,8'd250} : s = 504;
	{8'd254,8'd251} : s = 505;
	{8'd254,8'd252} : s = 506;
	{8'd254,8'd253} : s = 507;
	{8'd254,8'd254} : s = 508;
	{8'd254,8'd255} : s = 509;
	{8'd255,8'd0} : s = 255;
	{8'd255,8'd1} : s = 256;
	{8'd255,8'd2} : s = 257;
	{8'd255,8'd3} : s = 258;
	{8'd255,8'd4} : s = 259;
	{8'd255,8'd5} : s = 260;
	{8'd255,8'd6} : s = 261;
	{8'd255,8'd7} : s = 262;
	{8'd255,8'd8} : s = 263;
	{8'd255,8'd9} : s = 264;
	{8'd255,8'd10} : s = 265;
	{8'd255,8'd11} : s = 266;
	{8'd255,8'd12} : s = 267;
	{8'd255,8'd13} : s = 268;
	{8'd255,8'd14} : s = 269;
	{8'd255,8'd15} : s = 270;
	{8'd255,8'd16} : s = 271;
	{8'd255,8'd17} : s = 272;
	{8'd255,8'd18} : s = 273;
	{8'd255,8'd19} : s = 274;
	{8'd255,8'd20} : s = 275;
	{8'd255,8'd21} : s = 276;
	{8'd255,8'd22} : s = 277;
	{8'd255,8'd23} : s = 278;
	{8'd255,8'd24} : s = 279;
	{8'd255,8'd25} : s = 280;
	{8'd255,8'd26} : s = 281;
	{8'd255,8'd27} : s = 282;
	{8'd255,8'd28} : s = 283;
	{8'd255,8'd29} : s = 284;
	{8'd255,8'd30} : s = 285;
	{8'd255,8'd31} : s = 286;
	{8'd255,8'd32} : s = 287;
	{8'd255,8'd33} : s = 288;
	{8'd255,8'd34} : s = 289;
	{8'd255,8'd35} : s = 290;
	{8'd255,8'd36} : s = 291;
	{8'd255,8'd37} : s = 292;
	{8'd255,8'd38} : s = 293;
	{8'd255,8'd39} : s = 294;
	{8'd255,8'd40} : s = 295;
	{8'd255,8'd41} : s = 296;
	{8'd255,8'd42} : s = 297;
	{8'd255,8'd43} : s = 298;
	{8'd255,8'd44} : s = 299;
	{8'd255,8'd45} : s = 300;
	{8'd255,8'd46} : s = 301;
	{8'd255,8'd47} : s = 302;
	{8'd255,8'd48} : s = 303;
	{8'd255,8'd49} : s = 304;
	{8'd255,8'd50} : s = 305;
	{8'd255,8'd51} : s = 306;
	{8'd255,8'd52} : s = 307;
	{8'd255,8'd53} : s = 308;
	{8'd255,8'd54} : s = 309;
	{8'd255,8'd55} : s = 310;
	{8'd255,8'd56} : s = 311;
	{8'd255,8'd57} : s = 312;
	{8'd255,8'd58} : s = 313;
	{8'd255,8'd59} : s = 314;
	{8'd255,8'd60} : s = 315;
	{8'd255,8'd61} : s = 316;
	{8'd255,8'd62} : s = 317;
	{8'd255,8'd63} : s = 318;
	{8'd255,8'd64} : s = 319;
	{8'd255,8'd65} : s = 320;
	{8'd255,8'd66} : s = 321;
	{8'd255,8'd67} : s = 322;
	{8'd255,8'd68} : s = 323;
	{8'd255,8'd69} : s = 324;
	{8'd255,8'd70} : s = 325;
	{8'd255,8'd71} : s = 326;
	{8'd255,8'd72} : s = 327;
	{8'd255,8'd73} : s = 328;
	{8'd255,8'd74} : s = 329;
	{8'd255,8'd75} : s = 330;
	{8'd255,8'd76} : s = 331;
	{8'd255,8'd77} : s = 332;
	{8'd255,8'd78} : s = 333;
	{8'd255,8'd79} : s = 334;
	{8'd255,8'd80} : s = 335;
	{8'd255,8'd81} : s = 336;
	{8'd255,8'd82} : s = 337;
	{8'd255,8'd83} : s = 338;
	{8'd255,8'd84} : s = 339;
	{8'd255,8'd85} : s = 340;
	{8'd255,8'd86} : s = 341;
	{8'd255,8'd87} : s = 342;
	{8'd255,8'd88} : s = 343;
	{8'd255,8'd89} : s = 344;
	{8'd255,8'd90} : s = 345;
	{8'd255,8'd91} : s = 346;
	{8'd255,8'd92} : s = 347;
	{8'd255,8'd93} : s = 348;
	{8'd255,8'd94} : s = 349;
	{8'd255,8'd95} : s = 350;
	{8'd255,8'd96} : s = 351;
	{8'd255,8'd97} : s = 352;
	{8'd255,8'd98} : s = 353;
	{8'd255,8'd99} : s = 354;
	{8'd255,8'd100} : s = 355;
	{8'd255,8'd101} : s = 356;
	{8'd255,8'd102} : s = 357;
	{8'd255,8'd103} : s = 358;
	{8'd255,8'd104} : s = 359;
	{8'd255,8'd105} : s = 360;
	{8'd255,8'd106} : s = 361;
	{8'd255,8'd107} : s = 362;
	{8'd255,8'd108} : s = 363;
	{8'd255,8'd109} : s = 364;
	{8'd255,8'd110} : s = 365;
	{8'd255,8'd111} : s = 366;
	{8'd255,8'd112} : s = 367;
	{8'd255,8'd113} : s = 368;
	{8'd255,8'd114} : s = 369;
	{8'd255,8'd115} : s = 370;
	{8'd255,8'd116} : s = 371;
	{8'd255,8'd117} : s = 372;
	{8'd255,8'd118} : s = 373;
	{8'd255,8'd119} : s = 374;
	{8'd255,8'd120} : s = 375;
	{8'd255,8'd121} : s = 376;
	{8'd255,8'd122} : s = 377;
	{8'd255,8'd123} : s = 378;
	{8'd255,8'd124} : s = 379;
	{8'd255,8'd125} : s = 380;
	{8'd255,8'd126} : s = 381;
	{8'd255,8'd127} : s = 382;
	{8'd255,8'd128} : s = 383;
	{8'd255,8'd129} : s = 384;
	{8'd255,8'd130} : s = 385;
	{8'd255,8'd131} : s = 386;
	{8'd255,8'd132} : s = 387;
	{8'd255,8'd133} : s = 388;
	{8'd255,8'd134} : s = 389;
	{8'd255,8'd135} : s = 390;
	{8'd255,8'd136} : s = 391;
	{8'd255,8'd137} : s = 392;
	{8'd255,8'd138} : s = 393;
	{8'd255,8'd139} : s = 394;
	{8'd255,8'd140} : s = 395;
	{8'd255,8'd141} : s = 396;
	{8'd255,8'd142} : s = 397;
	{8'd255,8'd143} : s = 398;
	{8'd255,8'd144} : s = 399;
	{8'd255,8'd145} : s = 400;
	{8'd255,8'd146} : s = 401;
	{8'd255,8'd147} : s = 402;
	{8'd255,8'd148} : s = 403;
	{8'd255,8'd149} : s = 404;
	{8'd255,8'd150} : s = 405;
	{8'd255,8'd151} : s = 406;
	{8'd255,8'd152} : s = 407;
	{8'd255,8'd153} : s = 408;
	{8'd255,8'd154} : s = 409;
	{8'd255,8'd155} : s = 410;
	{8'd255,8'd156} : s = 411;
	{8'd255,8'd157} : s = 412;
	{8'd255,8'd158} : s = 413;
	{8'd255,8'd159} : s = 414;
	{8'd255,8'd160} : s = 415;
	{8'd255,8'd161} : s = 416;
	{8'd255,8'd162} : s = 417;
	{8'd255,8'd163} : s = 418;
	{8'd255,8'd164} : s = 419;
	{8'd255,8'd165} : s = 420;
	{8'd255,8'd166} : s = 421;
	{8'd255,8'd167} : s = 422;
	{8'd255,8'd168} : s = 423;
	{8'd255,8'd169} : s = 424;
	{8'd255,8'd170} : s = 425;
	{8'd255,8'd171} : s = 426;
	{8'd255,8'd172} : s = 427;
	{8'd255,8'd173} : s = 428;
	{8'd255,8'd174} : s = 429;
	{8'd255,8'd175} : s = 430;
	{8'd255,8'd176} : s = 431;
	{8'd255,8'd177} : s = 432;
	{8'd255,8'd178} : s = 433;
	{8'd255,8'd179} : s = 434;
	{8'd255,8'd180} : s = 435;
	{8'd255,8'd181} : s = 436;
	{8'd255,8'd182} : s = 437;
	{8'd255,8'd183} : s = 438;
	{8'd255,8'd184} : s = 439;
	{8'd255,8'd185} : s = 440;
	{8'd255,8'd186} : s = 441;
	{8'd255,8'd187} : s = 442;
	{8'd255,8'd188} : s = 443;
	{8'd255,8'd189} : s = 444;
	{8'd255,8'd190} : s = 445;
	{8'd255,8'd191} : s = 446;
	{8'd255,8'd192} : s = 447;
	{8'd255,8'd193} : s = 448;
	{8'd255,8'd194} : s = 449;
	{8'd255,8'd195} : s = 450;
	{8'd255,8'd196} : s = 451;
	{8'd255,8'd197} : s = 452;
	{8'd255,8'd198} : s = 453;
	{8'd255,8'd199} : s = 454;
	{8'd255,8'd200} : s = 455;
	{8'd255,8'd201} : s = 456;
	{8'd255,8'd202} : s = 457;
	{8'd255,8'd203} : s = 458;
	{8'd255,8'd204} : s = 459;
	{8'd255,8'd205} : s = 460;
	{8'd255,8'd206} : s = 461;
	{8'd255,8'd207} : s = 462;
	{8'd255,8'd208} : s = 463;
	{8'd255,8'd209} : s = 464;
	{8'd255,8'd210} : s = 465;
	{8'd255,8'd211} : s = 466;
	{8'd255,8'd212} : s = 467;
	{8'd255,8'd213} : s = 468;
	{8'd255,8'd214} : s = 469;
	{8'd255,8'd215} : s = 470;
	{8'd255,8'd216} : s = 471;
	{8'd255,8'd217} : s = 472;
	{8'd255,8'd218} : s = 473;
	{8'd255,8'd219} : s = 474;
	{8'd255,8'd220} : s = 475;
	{8'd255,8'd221} : s = 476;
	{8'd255,8'd222} : s = 477;
	{8'd255,8'd223} : s = 478;
	{8'd255,8'd224} : s = 479;
	{8'd255,8'd225} : s = 480;
	{8'd255,8'd226} : s = 481;
	{8'd255,8'd227} : s = 482;
	{8'd255,8'd228} : s = 483;
	{8'd255,8'd229} : s = 484;
	{8'd255,8'd230} : s = 485;
	{8'd255,8'd231} : s = 486;
	{8'd255,8'd232} : s = 487;
	{8'd255,8'd233} : s = 488;
	{8'd255,8'd234} : s = 489;
	{8'd255,8'd235} : s = 490;
	{8'd255,8'd236} : s = 491;
	{8'd255,8'd237} : s = 492;
	{8'd255,8'd238} : s = 493;
	{8'd255,8'd239} : s = 494;
	{8'd255,8'd240} : s = 495;
	{8'd255,8'd241} : s = 496;
	{8'd255,8'd242} : s = 497;
	{8'd255,8'd243} : s = 498;
	{8'd255,8'd244} : s = 499;
	{8'd255,8'd245} : s = 500;
	{8'd255,8'd246} : s = 501;
	{8'd255,8'd247} : s = 502;
	{8'd255,8'd248} : s = 503;
	{8'd255,8'd249} : s = 504;
	{8'd255,8'd250} : s = 505;
	{8'd255,8'd251} : s = 506;
	{8'd255,8'd252} : s = 507;
	{8'd255,8'd253} : s = 508;
	{8'd255,8'd254} : s = 509;
	{8'd255,8'd255} : s = 510;
    endcase
end
endmodule
