module gen_nonlinear_part(a,b,n);
input  [11:0] a, b; //adder inputs
output [8176:0] n; // non-linear outputs

wire [8177:0] g;

assign g[0] = 0;
//Assigning outputs for input bit 0
assign g[1] = a[0] & b[0];
assign g[2] = a[0] & g[0];
assign g[3] = b[0] & g[0];
//Assigning outputs for input bit 1
assign g[4] = a[1] & b[1];
assign g[5] = a[1] & g[1];
assign g[8] = b[1] & g[1];
assign g[6] = a[1] & g[2];
assign g[9] = b[1] & g[2];
assign g[7] = a[1] & g[3];
assign g[10] = b[1] & g[3];
//Assigning outputs for input bit 2
assign g[11] = a[2] & b[2];
assign g[12] = a[2] & g[4];
assign g[19] = b[2] & g[4];
assign g[13] = a[2] & g[5];
assign g[20] = b[2] & g[5];
assign g[14] = a[2] & g[6];
assign g[21] = b[2] & g[6];
assign g[15] = a[2] & g[7];
assign g[22] = b[2] & g[7];
assign g[16] = a[2] & g[8];
assign g[23] = b[2] & g[8];
assign g[17] = a[2] & g[9];
assign g[24] = b[2] & g[9];
assign g[18] = a[2] & g[10];
assign g[25] = b[2] & g[10];
//Assigning outputs for input bit 3
assign g[26] = a[3] & b[3];
assign g[27] = a[3] & g[11];
assign g[42] = b[3] & g[11];
assign g[28] = a[3] & g[12];
assign g[43] = b[3] & g[12];
assign g[29] = a[3] & g[13];
assign g[44] = b[3] & g[13];
assign g[30] = a[3] & g[14];
assign g[45] = b[3] & g[14];
assign g[31] = a[3] & g[15];
assign g[46] = b[3] & g[15];
assign g[32] = a[3] & g[16];
assign g[47] = b[3] & g[16];
assign g[33] = a[3] & g[17];
assign g[48] = b[3] & g[17];
assign g[34] = a[3] & g[18];
assign g[49] = b[3] & g[18];
assign g[35] = a[3] & g[19];
assign g[50] = b[3] & g[19];
assign g[36] = a[3] & g[20];
assign g[51] = b[3] & g[20];
assign g[37] = a[3] & g[21];
assign g[52] = b[3] & g[21];
assign g[38] = a[3] & g[22];
assign g[53] = b[3] & g[22];
assign g[39] = a[3] & g[23];
assign g[54] = b[3] & g[23];
assign g[40] = a[3] & g[24];
assign g[55] = b[3] & g[24];
assign g[41] = a[3] & g[25];
assign g[56] = b[3] & g[25];
//Assigning outputs for input bit 4
assign g[57] = a[4] & b[4];
assign g[58] = a[4] & g[26];
assign g[89] = b[4] & g[26];
assign g[59] = a[4] & g[27];
assign g[90] = b[4] & g[27];
assign g[60] = a[4] & g[28];
assign g[91] = b[4] & g[28];
assign g[61] = a[4] & g[29];
assign g[92] = b[4] & g[29];
assign g[62] = a[4] & g[30];
assign g[93] = b[4] & g[30];
assign g[63] = a[4] & g[31];
assign g[94] = b[4] & g[31];
assign g[64] = a[4] & g[32];
assign g[95] = b[4] & g[32];
assign g[65] = a[4] & g[33];
assign g[96] = b[4] & g[33];
assign g[66] = a[4] & g[34];
assign g[97] = b[4] & g[34];
assign g[67] = a[4] & g[35];
assign g[98] = b[4] & g[35];
assign g[68] = a[4] & g[36];
assign g[99] = b[4] & g[36];
assign g[69] = a[4] & g[37];
assign g[100] = b[4] & g[37];
assign g[70] = a[4] & g[38];
assign g[101] = b[4] & g[38];
assign g[71] = a[4] & g[39];
assign g[102] = b[4] & g[39];
assign g[72] = a[4] & g[40];
assign g[103] = b[4] & g[40];
assign g[73] = a[4] & g[41];
assign g[104] = b[4] & g[41];
assign g[74] = a[4] & g[42];
assign g[105] = b[4] & g[42];
assign g[75] = a[4] & g[43];
assign g[106] = b[4] & g[43];
assign g[76] = a[4] & g[44];
assign g[107] = b[4] & g[44];
assign g[77] = a[4] & g[45];
assign g[108] = b[4] & g[45];
assign g[78] = a[4] & g[46];
assign g[109] = b[4] & g[46];
assign g[79] = a[4] & g[47];
assign g[110] = b[4] & g[47];
assign g[80] = a[4] & g[48];
assign g[111] = b[4] & g[48];
assign g[81] = a[4] & g[49];
assign g[112] = b[4] & g[49];
assign g[82] = a[4] & g[50];
assign g[113] = b[4] & g[50];
assign g[83] = a[4] & g[51];
assign g[114] = b[4] & g[51];
assign g[84] = a[4] & g[52];
assign g[115] = b[4] & g[52];
assign g[85] = a[4] & g[53];
assign g[116] = b[4] & g[53];
assign g[86] = a[4] & g[54];
assign g[117] = b[4] & g[54];
assign g[87] = a[4] & g[55];
assign g[118] = b[4] & g[55];
assign g[88] = a[4] & g[56];
assign g[119] = b[4] & g[56];
//Assigning outputs for input bit 5
assign g[120] = a[5] & b[5];
assign g[121] = a[5] & g[57];
assign g[184] = b[5] & g[57];
assign g[122] = a[5] & g[58];
assign g[185] = b[5] & g[58];
assign g[123] = a[5] & g[59];
assign g[186] = b[5] & g[59];
assign g[124] = a[5] & g[60];
assign g[187] = b[5] & g[60];
assign g[125] = a[5] & g[61];
assign g[188] = b[5] & g[61];
assign g[126] = a[5] & g[62];
assign g[189] = b[5] & g[62];
assign g[127] = a[5] & g[63];
assign g[190] = b[5] & g[63];
assign g[128] = a[5] & g[64];
assign g[191] = b[5] & g[64];
assign g[129] = a[5] & g[65];
assign g[192] = b[5] & g[65];
assign g[130] = a[5] & g[66];
assign g[193] = b[5] & g[66];
assign g[131] = a[5] & g[67];
assign g[194] = b[5] & g[67];
assign g[132] = a[5] & g[68];
assign g[195] = b[5] & g[68];
assign g[133] = a[5] & g[69];
assign g[196] = b[5] & g[69];
assign g[134] = a[5] & g[70];
assign g[197] = b[5] & g[70];
assign g[135] = a[5] & g[71];
assign g[198] = b[5] & g[71];
assign g[136] = a[5] & g[72];
assign g[199] = b[5] & g[72];
assign g[137] = a[5] & g[73];
assign g[200] = b[5] & g[73];
assign g[138] = a[5] & g[74];
assign g[201] = b[5] & g[74];
assign g[139] = a[5] & g[75];
assign g[202] = b[5] & g[75];
assign g[140] = a[5] & g[76];
assign g[203] = b[5] & g[76];
assign g[141] = a[5] & g[77];
assign g[204] = b[5] & g[77];
assign g[142] = a[5] & g[78];
assign g[205] = b[5] & g[78];
assign g[143] = a[5] & g[79];
assign g[206] = b[5] & g[79];
assign g[144] = a[5] & g[80];
assign g[207] = b[5] & g[80];
assign g[145] = a[5] & g[81];
assign g[208] = b[5] & g[81];
assign g[146] = a[5] & g[82];
assign g[209] = b[5] & g[82];
assign g[147] = a[5] & g[83];
assign g[210] = b[5] & g[83];
assign g[148] = a[5] & g[84];
assign g[211] = b[5] & g[84];
assign g[149] = a[5] & g[85];
assign g[212] = b[5] & g[85];
assign g[150] = a[5] & g[86];
assign g[213] = b[5] & g[86];
assign g[151] = a[5] & g[87];
assign g[214] = b[5] & g[87];
assign g[152] = a[5] & g[88];
assign g[215] = b[5] & g[88];
assign g[153] = a[5] & g[89];
assign g[216] = b[5] & g[89];
assign g[154] = a[5] & g[90];
assign g[217] = b[5] & g[90];
assign g[155] = a[5] & g[91];
assign g[218] = b[5] & g[91];
assign g[156] = a[5] & g[92];
assign g[219] = b[5] & g[92];
assign g[157] = a[5] & g[93];
assign g[220] = b[5] & g[93];
assign g[158] = a[5] & g[94];
assign g[221] = b[5] & g[94];
assign g[159] = a[5] & g[95];
assign g[222] = b[5] & g[95];
assign g[160] = a[5] & g[96];
assign g[223] = b[5] & g[96];
assign g[161] = a[5] & g[97];
assign g[224] = b[5] & g[97];
assign g[162] = a[5] & g[98];
assign g[225] = b[5] & g[98];
assign g[163] = a[5] & g[99];
assign g[226] = b[5] & g[99];
assign g[164] = a[5] & g[100];
assign g[227] = b[5] & g[100];
assign g[165] = a[5] & g[101];
assign g[228] = b[5] & g[101];
assign g[166] = a[5] & g[102];
assign g[229] = b[5] & g[102];
assign g[167] = a[5] & g[103];
assign g[230] = b[5] & g[103];
assign g[168] = a[5] & g[104];
assign g[231] = b[5] & g[104];
assign g[169] = a[5] & g[105];
assign g[232] = b[5] & g[105];
assign g[170] = a[5] & g[106];
assign g[233] = b[5] & g[106];
assign g[171] = a[5] & g[107];
assign g[234] = b[5] & g[107];
assign g[172] = a[5] & g[108];
assign g[235] = b[5] & g[108];
assign g[173] = a[5] & g[109];
assign g[236] = b[5] & g[109];
assign g[174] = a[5] & g[110];
assign g[237] = b[5] & g[110];
assign g[175] = a[5] & g[111];
assign g[238] = b[5] & g[111];
assign g[176] = a[5] & g[112];
assign g[239] = b[5] & g[112];
assign g[177] = a[5] & g[113];
assign g[240] = b[5] & g[113];
assign g[178] = a[5] & g[114];
assign g[241] = b[5] & g[114];
assign g[179] = a[5] & g[115];
assign g[242] = b[5] & g[115];
assign g[180] = a[5] & g[116];
assign g[243] = b[5] & g[116];
assign g[181] = a[5] & g[117];
assign g[244] = b[5] & g[117];
assign g[182] = a[5] & g[118];
assign g[245] = b[5] & g[118];
assign g[183] = a[5] & g[119];
assign g[246] = b[5] & g[119];
//Assigning outputs for input bit 6
assign g[247] = a[6] & b[6];
assign g[248] = a[6] & g[120];
assign g[375] = b[6] & g[120];
assign g[249] = a[6] & g[121];
assign g[376] = b[6] & g[121];
assign g[250] = a[6] & g[122];
assign g[377] = b[6] & g[122];
assign g[251] = a[6] & g[123];
assign g[378] = b[6] & g[123];
assign g[252] = a[6] & g[124];
assign g[379] = b[6] & g[124];
assign g[253] = a[6] & g[125];
assign g[380] = b[6] & g[125];
assign g[254] = a[6] & g[126];
assign g[381] = b[6] & g[126];
assign g[255] = a[6] & g[127];
assign g[382] = b[6] & g[127];
assign g[256] = a[6] & g[128];
assign g[383] = b[6] & g[128];
assign g[257] = a[6] & g[129];
assign g[384] = b[6] & g[129];
assign g[258] = a[6] & g[130];
assign g[385] = b[6] & g[130];
assign g[259] = a[6] & g[131];
assign g[386] = b[6] & g[131];
assign g[260] = a[6] & g[132];
assign g[387] = b[6] & g[132];
assign g[261] = a[6] & g[133];
assign g[388] = b[6] & g[133];
assign g[262] = a[6] & g[134];
assign g[389] = b[6] & g[134];
assign g[263] = a[6] & g[135];
assign g[390] = b[6] & g[135];
assign g[264] = a[6] & g[136];
assign g[391] = b[6] & g[136];
assign g[265] = a[6] & g[137];
assign g[392] = b[6] & g[137];
assign g[266] = a[6] & g[138];
assign g[393] = b[6] & g[138];
assign g[267] = a[6] & g[139];
assign g[394] = b[6] & g[139];
assign g[268] = a[6] & g[140];
assign g[395] = b[6] & g[140];
assign g[269] = a[6] & g[141];
assign g[396] = b[6] & g[141];
assign g[270] = a[6] & g[142];
assign g[397] = b[6] & g[142];
assign g[271] = a[6] & g[143];
assign g[398] = b[6] & g[143];
assign g[272] = a[6] & g[144];
assign g[399] = b[6] & g[144];
assign g[273] = a[6] & g[145];
assign g[400] = b[6] & g[145];
assign g[274] = a[6] & g[146];
assign g[401] = b[6] & g[146];
assign g[275] = a[6] & g[147];
assign g[402] = b[6] & g[147];
assign g[276] = a[6] & g[148];
assign g[403] = b[6] & g[148];
assign g[277] = a[6] & g[149];
assign g[404] = b[6] & g[149];
assign g[278] = a[6] & g[150];
assign g[405] = b[6] & g[150];
assign g[279] = a[6] & g[151];
assign g[406] = b[6] & g[151];
assign g[280] = a[6] & g[152];
assign g[407] = b[6] & g[152];
assign g[281] = a[6] & g[153];
assign g[408] = b[6] & g[153];
assign g[282] = a[6] & g[154];
assign g[409] = b[6] & g[154];
assign g[283] = a[6] & g[155];
assign g[410] = b[6] & g[155];
assign g[284] = a[6] & g[156];
assign g[411] = b[6] & g[156];
assign g[285] = a[6] & g[157];
assign g[412] = b[6] & g[157];
assign g[286] = a[6] & g[158];
assign g[413] = b[6] & g[158];
assign g[287] = a[6] & g[159];
assign g[414] = b[6] & g[159];
assign g[288] = a[6] & g[160];
assign g[415] = b[6] & g[160];
assign g[289] = a[6] & g[161];
assign g[416] = b[6] & g[161];
assign g[290] = a[6] & g[162];
assign g[417] = b[6] & g[162];
assign g[291] = a[6] & g[163];
assign g[418] = b[6] & g[163];
assign g[292] = a[6] & g[164];
assign g[419] = b[6] & g[164];
assign g[293] = a[6] & g[165];
assign g[420] = b[6] & g[165];
assign g[294] = a[6] & g[166];
assign g[421] = b[6] & g[166];
assign g[295] = a[6] & g[167];
assign g[422] = b[6] & g[167];
assign g[296] = a[6] & g[168];
assign g[423] = b[6] & g[168];
assign g[297] = a[6] & g[169];
assign g[424] = b[6] & g[169];
assign g[298] = a[6] & g[170];
assign g[425] = b[6] & g[170];
assign g[299] = a[6] & g[171];
assign g[426] = b[6] & g[171];
assign g[300] = a[6] & g[172];
assign g[427] = b[6] & g[172];
assign g[301] = a[6] & g[173];
assign g[428] = b[6] & g[173];
assign g[302] = a[6] & g[174];
assign g[429] = b[6] & g[174];
assign g[303] = a[6] & g[175];
assign g[430] = b[6] & g[175];
assign g[304] = a[6] & g[176];
assign g[431] = b[6] & g[176];
assign g[305] = a[6] & g[177];
assign g[432] = b[6] & g[177];
assign g[306] = a[6] & g[178];
assign g[433] = b[6] & g[178];
assign g[307] = a[6] & g[179];
assign g[434] = b[6] & g[179];
assign g[308] = a[6] & g[180];
assign g[435] = b[6] & g[180];
assign g[309] = a[6] & g[181];
assign g[436] = b[6] & g[181];
assign g[310] = a[6] & g[182];
assign g[437] = b[6] & g[182];
assign g[311] = a[6] & g[183];
assign g[438] = b[6] & g[183];
assign g[312] = a[6] & g[184];
assign g[439] = b[6] & g[184];
assign g[313] = a[6] & g[185];
assign g[440] = b[6] & g[185];
assign g[314] = a[6] & g[186];
assign g[441] = b[6] & g[186];
assign g[315] = a[6] & g[187];
assign g[442] = b[6] & g[187];
assign g[316] = a[6] & g[188];
assign g[443] = b[6] & g[188];
assign g[317] = a[6] & g[189];
assign g[444] = b[6] & g[189];
assign g[318] = a[6] & g[190];
assign g[445] = b[6] & g[190];
assign g[319] = a[6] & g[191];
assign g[446] = b[6] & g[191];
assign g[320] = a[6] & g[192];
assign g[447] = b[6] & g[192];
assign g[321] = a[6] & g[193];
assign g[448] = b[6] & g[193];
assign g[322] = a[6] & g[194];
assign g[449] = b[6] & g[194];
assign g[323] = a[6] & g[195];
assign g[450] = b[6] & g[195];
assign g[324] = a[6] & g[196];
assign g[451] = b[6] & g[196];
assign g[325] = a[6] & g[197];
assign g[452] = b[6] & g[197];
assign g[326] = a[6] & g[198];
assign g[453] = b[6] & g[198];
assign g[327] = a[6] & g[199];
assign g[454] = b[6] & g[199];
assign g[328] = a[6] & g[200];
assign g[455] = b[6] & g[200];
assign g[329] = a[6] & g[201];
assign g[456] = b[6] & g[201];
assign g[330] = a[6] & g[202];
assign g[457] = b[6] & g[202];
assign g[331] = a[6] & g[203];
assign g[458] = b[6] & g[203];
assign g[332] = a[6] & g[204];
assign g[459] = b[6] & g[204];
assign g[333] = a[6] & g[205];
assign g[460] = b[6] & g[205];
assign g[334] = a[6] & g[206];
assign g[461] = b[6] & g[206];
assign g[335] = a[6] & g[207];
assign g[462] = b[6] & g[207];
assign g[336] = a[6] & g[208];
assign g[463] = b[6] & g[208];
assign g[337] = a[6] & g[209];
assign g[464] = b[6] & g[209];
assign g[338] = a[6] & g[210];
assign g[465] = b[6] & g[210];
assign g[339] = a[6] & g[211];
assign g[466] = b[6] & g[211];
assign g[340] = a[6] & g[212];
assign g[467] = b[6] & g[212];
assign g[341] = a[6] & g[213];
assign g[468] = b[6] & g[213];
assign g[342] = a[6] & g[214];
assign g[469] = b[6] & g[214];
assign g[343] = a[6] & g[215];
assign g[470] = b[6] & g[215];
assign g[344] = a[6] & g[216];
assign g[471] = b[6] & g[216];
assign g[345] = a[6] & g[217];
assign g[472] = b[6] & g[217];
assign g[346] = a[6] & g[218];
assign g[473] = b[6] & g[218];
assign g[347] = a[6] & g[219];
assign g[474] = b[6] & g[219];
assign g[348] = a[6] & g[220];
assign g[475] = b[6] & g[220];
assign g[349] = a[6] & g[221];
assign g[476] = b[6] & g[221];
assign g[350] = a[6] & g[222];
assign g[477] = b[6] & g[222];
assign g[351] = a[6] & g[223];
assign g[478] = b[6] & g[223];
assign g[352] = a[6] & g[224];
assign g[479] = b[6] & g[224];
assign g[353] = a[6] & g[225];
assign g[480] = b[6] & g[225];
assign g[354] = a[6] & g[226];
assign g[481] = b[6] & g[226];
assign g[355] = a[6] & g[227];
assign g[482] = b[6] & g[227];
assign g[356] = a[6] & g[228];
assign g[483] = b[6] & g[228];
assign g[357] = a[6] & g[229];
assign g[484] = b[6] & g[229];
assign g[358] = a[6] & g[230];
assign g[485] = b[6] & g[230];
assign g[359] = a[6] & g[231];
assign g[486] = b[6] & g[231];
assign g[360] = a[6] & g[232];
assign g[487] = b[6] & g[232];
assign g[361] = a[6] & g[233];
assign g[488] = b[6] & g[233];
assign g[362] = a[6] & g[234];
assign g[489] = b[6] & g[234];
assign g[363] = a[6] & g[235];
assign g[490] = b[6] & g[235];
assign g[364] = a[6] & g[236];
assign g[491] = b[6] & g[236];
assign g[365] = a[6] & g[237];
assign g[492] = b[6] & g[237];
assign g[366] = a[6] & g[238];
assign g[493] = b[6] & g[238];
assign g[367] = a[6] & g[239];
assign g[494] = b[6] & g[239];
assign g[368] = a[6] & g[240];
assign g[495] = b[6] & g[240];
assign g[369] = a[6] & g[241];
assign g[496] = b[6] & g[241];
assign g[370] = a[6] & g[242];
assign g[497] = b[6] & g[242];
assign g[371] = a[6] & g[243];
assign g[498] = b[6] & g[243];
assign g[372] = a[6] & g[244];
assign g[499] = b[6] & g[244];
assign g[373] = a[6] & g[245];
assign g[500] = b[6] & g[245];
assign g[374] = a[6] & g[246];
assign g[501] = b[6] & g[246];
//Assigning outputs for input bit 7
assign g[502] = a[7] & b[7];
assign g[503] = a[7] & g[247];
assign g[758] = b[7] & g[247];
assign g[504] = a[7] & g[248];
assign g[759] = b[7] & g[248];
assign g[505] = a[7] & g[249];
assign g[760] = b[7] & g[249];
assign g[506] = a[7] & g[250];
assign g[761] = b[7] & g[250];
assign g[507] = a[7] & g[251];
assign g[762] = b[7] & g[251];
assign g[508] = a[7] & g[252];
assign g[763] = b[7] & g[252];
assign g[509] = a[7] & g[253];
assign g[764] = b[7] & g[253];
assign g[510] = a[7] & g[254];
assign g[765] = b[7] & g[254];
assign g[511] = a[7] & g[255];
assign g[766] = b[7] & g[255];
assign g[512] = a[7] & g[256];
assign g[767] = b[7] & g[256];
assign g[513] = a[7] & g[257];
assign g[768] = b[7] & g[257];
assign g[514] = a[7] & g[258];
assign g[769] = b[7] & g[258];
assign g[515] = a[7] & g[259];
assign g[770] = b[7] & g[259];
assign g[516] = a[7] & g[260];
assign g[771] = b[7] & g[260];
assign g[517] = a[7] & g[261];
assign g[772] = b[7] & g[261];
assign g[518] = a[7] & g[262];
assign g[773] = b[7] & g[262];
assign g[519] = a[7] & g[263];
assign g[774] = b[7] & g[263];
assign g[520] = a[7] & g[264];
assign g[775] = b[7] & g[264];
assign g[521] = a[7] & g[265];
assign g[776] = b[7] & g[265];
assign g[522] = a[7] & g[266];
assign g[777] = b[7] & g[266];
assign g[523] = a[7] & g[267];
assign g[778] = b[7] & g[267];
assign g[524] = a[7] & g[268];
assign g[779] = b[7] & g[268];
assign g[525] = a[7] & g[269];
assign g[780] = b[7] & g[269];
assign g[526] = a[7] & g[270];
assign g[781] = b[7] & g[270];
assign g[527] = a[7] & g[271];
assign g[782] = b[7] & g[271];
assign g[528] = a[7] & g[272];
assign g[783] = b[7] & g[272];
assign g[529] = a[7] & g[273];
assign g[784] = b[7] & g[273];
assign g[530] = a[7] & g[274];
assign g[785] = b[7] & g[274];
assign g[531] = a[7] & g[275];
assign g[786] = b[7] & g[275];
assign g[532] = a[7] & g[276];
assign g[787] = b[7] & g[276];
assign g[533] = a[7] & g[277];
assign g[788] = b[7] & g[277];
assign g[534] = a[7] & g[278];
assign g[789] = b[7] & g[278];
assign g[535] = a[7] & g[279];
assign g[790] = b[7] & g[279];
assign g[536] = a[7] & g[280];
assign g[791] = b[7] & g[280];
assign g[537] = a[7] & g[281];
assign g[792] = b[7] & g[281];
assign g[538] = a[7] & g[282];
assign g[793] = b[7] & g[282];
assign g[539] = a[7] & g[283];
assign g[794] = b[7] & g[283];
assign g[540] = a[7] & g[284];
assign g[795] = b[7] & g[284];
assign g[541] = a[7] & g[285];
assign g[796] = b[7] & g[285];
assign g[542] = a[7] & g[286];
assign g[797] = b[7] & g[286];
assign g[543] = a[7] & g[287];
assign g[798] = b[7] & g[287];
assign g[544] = a[7] & g[288];
assign g[799] = b[7] & g[288];
assign g[545] = a[7] & g[289];
assign g[800] = b[7] & g[289];
assign g[546] = a[7] & g[290];
assign g[801] = b[7] & g[290];
assign g[547] = a[7] & g[291];
assign g[802] = b[7] & g[291];
assign g[548] = a[7] & g[292];
assign g[803] = b[7] & g[292];
assign g[549] = a[7] & g[293];
assign g[804] = b[7] & g[293];
assign g[550] = a[7] & g[294];
assign g[805] = b[7] & g[294];
assign g[551] = a[7] & g[295];
assign g[806] = b[7] & g[295];
assign g[552] = a[7] & g[296];
assign g[807] = b[7] & g[296];
assign g[553] = a[7] & g[297];
assign g[808] = b[7] & g[297];
assign g[554] = a[7] & g[298];
assign g[809] = b[7] & g[298];
assign g[555] = a[7] & g[299];
assign g[810] = b[7] & g[299];
assign g[556] = a[7] & g[300];
assign g[811] = b[7] & g[300];
assign g[557] = a[7] & g[301];
assign g[812] = b[7] & g[301];
assign g[558] = a[7] & g[302];
assign g[813] = b[7] & g[302];
assign g[559] = a[7] & g[303];
assign g[814] = b[7] & g[303];
assign g[560] = a[7] & g[304];
assign g[815] = b[7] & g[304];
assign g[561] = a[7] & g[305];
assign g[816] = b[7] & g[305];
assign g[562] = a[7] & g[306];
assign g[817] = b[7] & g[306];
assign g[563] = a[7] & g[307];
assign g[818] = b[7] & g[307];
assign g[564] = a[7] & g[308];
assign g[819] = b[7] & g[308];
assign g[565] = a[7] & g[309];
assign g[820] = b[7] & g[309];
assign g[566] = a[7] & g[310];
assign g[821] = b[7] & g[310];
assign g[567] = a[7] & g[311];
assign g[822] = b[7] & g[311];
assign g[568] = a[7] & g[312];
assign g[823] = b[7] & g[312];
assign g[569] = a[7] & g[313];
assign g[824] = b[7] & g[313];
assign g[570] = a[7] & g[314];
assign g[825] = b[7] & g[314];
assign g[571] = a[7] & g[315];
assign g[826] = b[7] & g[315];
assign g[572] = a[7] & g[316];
assign g[827] = b[7] & g[316];
assign g[573] = a[7] & g[317];
assign g[828] = b[7] & g[317];
assign g[574] = a[7] & g[318];
assign g[829] = b[7] & g[318];
assign g[575] = a[7] & g[319];
assign g[830] = b[7] & g[319];
assign g[576] = a[7] & g[320];
assign g[831] = b[7] & g[320];
assign g[577] = a[7] & g[321];
assign g[832] = b[7] & g[321];
assign g[578] = a[7] & g[322];
assign g[833] = b[7] & g[322];
assign g[579] = a[7] & g[323];
assign g[834] = b[7] & g[323];
assign g[580] = a[7] & g[324];
assign g[835] = b[7] & g[324];
assign g[581] = a[7] & g[325];
assign g[836] = b[7] & g[325];
assign g[582] = a[7] & g[326];
assign g[837] = b[7] & g[326];
assign g[583] = a[7] & g[327];
assign g[838] = b[7] & g[327];
assign g[584] = a[7] & g[328];
assign g[839] = b[7] & g[328];
assign g[585] = a[7] & g[329];
assign g[840] = b[7] & g[329];
assign g[586] = a[7] & g[330];
assign g[841] = b[7] & g[330];
assign g[587] = a[7] & g[331];
assign g[842] = b[7] & g[331];
assign g[588] = a[7] & g[332];
assign g[843] = b[7] & g[332];
assign g[589] = a[7] & g[333];
assign g[844] = b[7] & g[333];
assign g[590] = a[7] & g[334];
assign g[845] = b[7] & g[334];
assign g[591] = a[7] & g[335];
assign g[846] = b[7] & g[335];
assign g[592] = a[7] & g[336];
assign g[847] = b[7] & g[336];
assign g[593] = a[7] & g[337];
assign g[848] = b[7] & g[337];
assign g[594] = a[7] & g[338];
assign g[849] = b[7] & g[338];
assign g[595] = a[7] & g[339];
assign g[850] = b[7] & g[339];
assign g[596] = a[7] & g[340];
assign g[851] = b[7] & g[340];
assign g[597] = a[7] & g[341];
assign g[852] = b[7] & g[341];
assign g[598] = a[7] & g[342];
assign g[853] = b[7] & g[342];
assign g[599] = a[7] & g[343];
assign g[854] = b[7] & g[343];
assign g[600] = a[7] & g[344];
assign g[855] = b[7] & g[344];
assign g[601] = a[7] & g[345];
assign g[856] = b[7] & g[345];
assign g[602] = a[7] & g[346];
assign g[857] = b[7] & g[346];
assign g[603] = a[7] & g[347];
assign g[858] = b[7] & g[347];
assign g[604] = a[7] & g[348];
assign g[859] = b[7] & g[348];
assign g[605] = a[7] & g[349];
assign g[860] = b[7] & g[349];
assign g[606] = a[7] & g[350];
assign g[861] = b[7] & g[350];
assign g[607] = a[7] & g[351];
assign g[862] = b[7] & g[351];
assign g[608] = a[7] & g[352];
assign g[863] = b[7] & g[352];
assign g[609] = a[7] & g[353];
assign g[864] = b[7] & g[353];
assign g[610] = a[7] & g[354];
assign g[865] = b[7] & g[354];
assign g[611] = a[7] & g[355];
assign g[866] = b[7] & g[355];
assign g[612] = a[7] & g[356];
assign g[867] = b[7] & g[356];
assign g[613] = a[7] & g[357];
assign g[868] = b[7] & g[357];
assign g[614] = a[7] & g[358];
assign g[869] = b[7] & g[358];
assign g[615] = a[7] & g[359];
assign g[870] = b[7] & g[359];
assign g[616] = a[7] & g[360];
assign g[871] = b[7] & g[360];
assign g[617] = a[7] & g[361];
assign g[872] = b[7] & g[361];
assign g[618] = a[7] & g[362];
assign g[873] = b[7] & g[362];
assign g[619] = a[7] & g[363];
assign g[874] = b[7] & g[363];
assign g[620] = a[7] & g[364];
assign g[875] = b[7] & g[364];
assign g[621] = a[7] & g[365];
assign g[876] = b[7] & g[365];
assign g[622] = a[7] & g[366];
assign g[877] = b[7] & g[366];
assign g[623] = a[7] & g[367];
assign g[878] = b[7] & g[367];
assign g[624] = a[7] & g[368];
assign g[879] = b[7] & g[368];
assign g[625] = a[7] & g[369];
assign g[880] = b[7] & g[369];
assign g[626] = a[7] & g[370];
assign g[881] = b[7] & g[370];
assign g[627] = a[7] & g[371];
assign g[882] = b[7] & g[371];
assign g[628] = a[7] & g[372];
assign g[883] = b[7] & g[372];
assign g[629] = a[7] & g[373];
assign g[884] = b[7] & g[373];
assign g[630] = a[7] & g[374];
assign g[885] = b[7] & g[374];
assign g[631] = a[7] & g[375];
assign g[886] = b[7] & g[375];
assign g[632] = a[7] & g[376];
assign g[887] = b[7] & g[376];
assign g[633] = a[7] & g[377];
assign g[888] = b[7] & g[377];
assign g[634] = a[7] & g[378];
assign g[889] = b[7] & g[378];
assign g[635] = a[7] & g[379];
assign g[890] = b[7] & g[379];
assign g[636] = a[7] & g[380];
assign g[891] = b[7] & g[380];
assign g[637] = a[7] & g[381];
assign g[892] = b[7] & g[381];
assign g[638] = a[7] & g[382];
assign g[893] = b[7] & g[382];
assign g[639] = a[7] & g[383];
assign g[894] = b[7] & g[383];
assign g[640] = a[7] & g[384];
assign g[895] = b[7] & g[384];
assign g[641] = a[7] & g[385];
assign g[896] = b[7] & g[385];
assign g[642] = a[7] & g[386];
assign g[897] = b[7] & g[386];
assign g[643] = a[7] & g[387];
assign g[898] = b[7] & g[387];
assign g[644] = a[7] & g[388];
assign g[899] = b[7] & g[388];
assign g[645] = a[7] & g[389];
assign g[900] = b[7] & g[389];
assign g[646] = a[7] & g[390];
assign g[901] = b[7] & g[390];
assign g[647] = a[7] & g[391];
assign g[902] = b[7] & g[391];
assign g[648] = a[7] & g[392];
assign g[903] = b[7] & g[392];
assign g[649] = a[7] & g[393];
assign g[904] = b[7] & g[393];
assign g[650] = a[7] & g[394];
assign g[905] = b[7] & g[394];
assign g[651] = a[7] & g[395];
assign g[906] = b[7] & g[395];
assign g[652] = a[7] & g[396];
assign g[907] = b[7] & g[396];
assign g[653] = a[7] & g[397];
assign g[908] = b[7] & g[397];
assign g[654] = a[7] & g[398];
assign g[909] = b[7] & g[398];
assign g[655] = a[7] & g[399];
assign g[910] = b[7] & g[399];
assign g[656] = a[7] & g[400];
assign g[911] = b[7] & g[400];
assign g[657] = a[7] & g[401];
assign g[912] = b[7] & g[401];
assign g[658] = a[7] & g[402];
assign g[913] = b[7] & g[402];
assign g[659] = a[7] & g[403];
assign g[914] = b[7] & g[403];
assign g[660] = a[7] & g[404];
assign g[915] = b[7] & g[404];
assign g[661] = a[7] & g[405];
assign g[916] = b[7] & g[405];
assign g[662] = a[7] & g[406];
assign g[917] = b[7] & g[406];
assign g[663] = a[7] & g[407];
assign g[918] = b[7] & g[407];
assign g[664] = a[7] & g[408];
assign g[919] = b[7] & g[408];
assign g[665] = a[7] & g[409];
assign g[920] = b[7] & g[409];
assign g[666] = a[7] & g[410];
assign g[921] = b[7] & g[410];
assign g[667] = a[7] & g[411];
assign g[922] = b[7] & g[411];
assign g[668] = a[7] & g[412];
assign g[923] = b[7] & g[412];
assign g[669] = a[7] & g[413];
assign g[924] = b[7] & g[413];
assign g[670] = a[7] & g[414];
assign g[925] = b[7] & g[414];
assign g[671] = a[7] & g[415];
assign g[926] = b[7] & g[415];
assign g[672] = a[7] & g[416];
assign g[927] = b[7] & g[416];
assign g[673] = a[7] & g[417];
assign g[928] = b[7] & g[417];
assign g[674] = a[7] & g[418];
assign g[929] = b[7] & g[418];
assign g[675] = a[7] & g[419];
assign g[930] = b[7] & g[419];
assign g[676] = a[7] & g[420];
assign g[931] = b[7] & g[420];
assign g[677] = a[7] & g[421];
assign g[932] = b[7] & g[421];
assign g[678] = a[7] & g[422];
assign g[933] = b[7] & g[422];
assign g[679] = a[7] & g[423];
assign g[934] = b[7] & g[423];
assign g[680] = a[7] & g[424];
assign g[935] = b[7] & g[424];
assign g[681] = a[7] & g[425];
assign g[936] = b[7] & g[425];
assign g[682] = a[7] & g[426];
assign g[937] = b[7] & g[426];
assign g[683] = a[7] & g[427];
assign g[938] = b[7] & g[427];
assign g[684] = a[7] & g[428];
assign g[939] = b[7] & g[428];
assign g[685] = a[7] & g[429];
assign g[940] = b[7] & g[429];
assign g[686] = a[7] & g[430];
assign g[941] = b[7] & g[430];
assign g[687] = a[7] & g[431];
assign g[942] = b[7] & g[431];
assign g[688] = a[7] & g[432];
assign g[943] = b[7] & g[432];
assign g[689] = a[7] & g[433];
assign g[944] = b[7] & g[433];
assign g[690] = a[7] & g[434];
assign g[945] = b[7] & g[434];
assign g[691] = a[7] & g[435];
assign g[946] = b[7] & g[435];
assign g[692] = a[7] & g[436];
assign g[947] = b[7] & g[436];
assign g[693] = a[7] & g[437];
assign g[948] = b[7] & g[437];
assign g[694] = a[7] & g[438];
assign g[949] = b[7] & g[438];
assign g[695] = a[7] & g[439];
assign g[950] = b[7] & g[439];
assign g[696] = a[7] & g[440];
assign g[951] = b[7] & g[440];
assign g[697] = a[7] & g[441];
assign g[952] = b[7] & g[441];
assign g[698] = a[7] & g[442];
assign g[953] = b[7] & g[442];
assign g[699] = a[7] & g[443];
assign g[954] = b[7] & g[443];
assign g[700] = a[7] & g[444];
assign g[955] = b[7] & g[444];
assign g[701] = a[7] & g[445];
assign g[956] = b[7] & g[445];
assign g[702] = a[7] & g[446];
assign g[957] = b[7] & g[446];
assign g[703] = a[7] & g[447];
assign g[958] = b[7] & g[447];
assign g[704] = a[7] & g[448];
assign g[959] = b[7] & g[448];
assign g[705] = a[7] & g[449];
assign g[960] = b[7] & g[449];
assign g[706] = a[7] & g[450];
assign g[961] = b[7] & g[450];
assign g[707] = a[7] & g[451];
assign g[962] = b[7] & g[451];
assign g[708] = a[7] & g[452];
assign g[963] = b[7] & g[452];
assign g[709] = a[7] & g[453];
assign g[964] = b[7] & g[453];
assign g[710] = a[7] & g[454];
assign g[965] = b[7] & g[454];
assign g[711] = a[7] & g[455];
assign g[966] = b[7] & g[455];
assign g[712] = a[7] & g[456];
assign g[967] = b[7] & g[456];
assign g[713] = a[7] & g[457];
assign g[968] = b[7] & g[457];
assign g[714] = a[7] & g[458];
assign g[969] = b[7] & g[458];
assign g[715] = a[7] & g[459];
assign g[970] = b[7] & g[459];
assign g[716] = a[7] & g[460];
assign g[971] = b[7] & g[460];
assign g[717] = a[7] & g[461];
assign g[972] = b[7] & g[461];
assign g[718] = a[7] & g[462];
assign g[973] = b[7] & g[462];
assign g[719] = a[7] & g[463];
assign g[974] = b[7] & g[463];
assign g[720] = a[7] & g[464];
assign g[975] = b[7] & g[464];
assign g[721] = a[7] & g[465];
assign g[976] = b[7] & g[465];
assign g[722] = a[7] & g[466];
assign g[977] = b[7] & g[466];
assign g[723] = a[7] & g[467];
assign g[978] = b[7] & g[467];
assign g[724] = a[7] & g[468];
assign g[979] = b[7] & g[468];
assign g[725] = a[7] & g[469];
assign g[980] = b[7] & g[469];
assign g[726] = a[7] & g[470];
assign g[981] = b[7] & g[470];
assign g[727] = a[7] & g[471];
assign g[982] = b[7] & g[471];
assign g[728] = a[7] & g[472];
assign g[983] = b[7] & g[472];
assign g[729] = a[7] & g[473];
assign g[984] = b[7] & g[473];
assign g[730] = a[7] & g[474];
assign g[985] = b[7] & g[474];
assign g[731] = a[7] & g[475];
assign g[986] = b[7] & g[475];
assign g[732] = a[7] & g[476];
assign g[987] = b[7] & g[476];
assign g[733] = a[7] & g[477];
assign g[988] = b[7] & g[477];
assign g[734] = a[7] & g[478];
assign g[989] = b[7] & g[478];
assign g[735] = a[7] & g[479];
assign g[990] = b[7] & g[479];
assign g[736] = a[7] & g[480];
assign g[991] = b[7] & g[480];
assign g[737] = a[7] & g[481];
assign g[992] = b[7] & g[481];
assign g[738] = a[7] & g[482];
assign g[993] = b[7] & g[482];
assign g[739] = a[7] & g[483];
assign g[994] = b[7] & g[483];
assign g[740] = a[7] & g[484];
assign g[995] = b[7] & g[484];
assign g[741] = a[7] & g[485];
assign g[996] = b[7] & g[485];
assign g[742] = a[7] & g[486];
assign g[997] = b[7] & g[486];
assign g[743] = a[7] & g[487];
assign g[998] = b[7] & g[487];
assign g[744] = a[7] & g[488];
assign g[999] = b[7] & g[488];
assign g[745] = a[7] & g[489];
assign g[1000] = b[7] & g[489];
assign g[746] = a[7] & g[490];
assign g[1001] = b[7] & g[490];
assign g[747] = a[7] & g[491];
assign g[1002] = b[7] & g[491];
assign g[748] = a[7] & g[492];
assign g[1003] = b[7] & g[492];
assign g[749] = a[7] & g[493];
assign g[1004] = b[7] & g[493];
assign g[750] = a[7] & g[494];
assign g[1005] = b[7] & g[494];
assign g[751] = a[7] & g[495];
assign g[1006] = b[7] & g[495];
assign g[752] = a[7] & g[496];
assign g[1007] = b[7] & g[496];
assign g[753] = a[7] & g[497];
assign g[1008] = b[7] & g[497];
assign g[754] = a[7] & g[498];
assign g[1009] = b[7] & g[498];
assign g[755] = a[7] & g[499];
assign g[1010] = b[7] & g[499];
assign g[756] = a[7] & g[500];
assign g[1011] = b[7] & g[500];
assign g[757] = a[7] & g[501];
assign g[1012] = b[7] & g[501];
//Assigning outputs for input bit 8
assign g[1013] = a[8] & b[8];
assign g[1014] = a[8] & g[502];
assign g[1525] = b[8] & g[502];
assign g[1015] = a[8] & g[503];
assign g[1526] = b[8] & g[503];
assign g[1016] = a[8] & g[504];
assign g[1527] = b[8] & g[504];
assign g[1017] = a[8] & g[505];
assign g[1528] = b[8] & g[505];
assign g[1018] = a[8] & g[506];
assign g[1529] = b[8] & g[506];
assign g[1019] = a[8] & g[507];
assign g[1530] = b[8] & g[507];
assign g[1020] = a[8] & g[508];
assign g[1531] = b[8] & g[508];
assign g[1021] = a[8] & g[509];
assign g[1532] = b[8] & g[509];
assign g[1022] = a[8] & g[510];
assign g[1533] = b[8] & g[510];
assign g[1023] = a[8] & g[511];
assign g[1534] = b[8] & g[511];
assign g[1024] = a[8] & g[512];
assign g[1535] = b[8] & g[512];
assign g[1025] = a[8] & g[513];
assign g[1536] = b[8] & g[513];
assign g[1026] = a[8] & g[514];
assign g[1537] = b[8] & g[514];
assign g[1027] = a[8] & g[515];
assign g[1538] = b[8] & g[515];
assign g[1028] = a[8] & g[516];
assign g[1539] = b[8] & g[516];
assign g[1029] = a[8] & g[517];
assign g[1540] = b[8] & g[517];
assign g[1030] = a[8] & g[518];
assign g[1541] = b[8] & g[518];
assign g[1031] = a[8] & g[519];
assign g[1542] = b[8] & g[519];
assign g[1032] = a[8] & g[520];
assign g[1543] = b[8] & g[520];
assign g[1033] = a[8] & g[521];
assign g[1544] = b[8] & g[521];
assign g[1034] = a[8] & g[522];
assign g[1545] = b[8] & g[522];
assign g[1035] = a[8] & g[523];
assign g[1546] = b[8] & g[523];
assign g[1036] = a[8] & g[524];
assign g[1547] = b[8] & g[524];
assign g[1037] = a[8] & g[525];
assign g[1548] = b[8] & g[525];
assign g[1038] = a[8] & g[526];
assign g[1549] = b[8] & g[526];
assign g[1039] = a[8] & g[527];
assign g[1550] = b[8] & g[527];
assign g[1040] = a[8] & g[528];
assign g[1551] = b[8] & g[528];
assign g[1041] = a[8] & g[529];
assign g[1552] = b[8] & g[529];
assign g[1042] = a[8] & g[530];
assign g[1553] = b[8] & g[530];
assign g[1043] = a[8] & g[531];
assign g[1554] = b[8] & g[531];
assign g[1044] = a[8] & g[532];
assign g[1555] = b[8] & g[532];
assign g[1045] = a[8] & g[533];
assign g[1556] = b[8] & g[533];
assign g[1046] = a[8] & g[534];
assign g[1557] = b[8] & g[534];
assign g[1047] = a[8] & g[535];
assign g[1558] = b[8] & g[535];
assign g[1048] = a[8] & g[536];
assign g[1559] = b[8] & g[536];
assign g[1049] = a[8] & g[537];
assign g[1560] = b[8] & g[537];
assign g[1050] = a[8] & g[538];
assign g[1561] = b[8] & g[538];
assign g[1051] = a[8] & g[539];
assign g[1562] = b[8] & g[539];
assign g[1052] = a[8] & g[540];
assign g[1563] = b[8] & g[540];
assign g[1053] = a[8] & g[541];
assign g[1564] = b[8] & g[541];
assign g[1054] = a[8] & g[542];
assign g[1565] = b[8] & g[542];
assign g[1055] = a[8] & g[543];
assign g[1566] = b[8] & g[543];
assign g[1056] = a[8] & g[544];
assign g[1567] = b[8] & g[544];
assign g[1057] = a[8] & g[545];
assign g[1568] = b[8] & g[545];
assign g[1058] = a[8] & g[546];
assign g[1569] = b[8] & g[546];
assign g[1059] = a[8] & g[547];
assign g[1570] = b[8] & g[547];
assign g[1060] = a[8] & g[548];
assign g[1571] = b[8] & g[548];
assign g[1061] = a[8] & g[549];
assign g[1572] = b[8] & g[549];
assign g[1062] = a[8] & g[550];
assign g[1573] = b[8] & g[550];
assign g[1063] = a[8] & g[551];
assign g[1574] = b[8] & g[551];
assign g[1064] = a[8] & g[552];
assign g[1575] = b[8] & g[552];
assign g[1065] = a[8] & g[553];
assign g[1576] = b[8] & g[553];
assign g[1066] = a[8] & g[554];
assign g[1577] = b[8] & g[554];
assign g[1067] = a[8] & g[555];
assign g[1578] = b[8] & g[555];
assign g[1068] = a[8] & g[556];
assign g[1579] = b[8] & g[556];
assign g[1069] = a[8] & g[557];
assign g[1580] = b[8] & g[557];
assign g[1070] = a[8] & g[558];
assign g[1581] = b[8] & g[558];
assign g[1071] = a[8] & g[559];
assign g[1582] = b[8] & g[559];
assign g[1072] = a[8] & g[560];
assign g[1583] = b[8] & g[560];
assign g[1073] = a[8] & g[561];
assign g[1584] = b[8] & g[561];
assign g[1074] = a[8] & g[562];
assign g[1585] = b[8] & g[562];
assign g[1075] = a[8] & g[563];
assign g[1586] = b[8] & g[563];
assign g[1076] = a[8] & g[564];
assign g[1587] = b[8] & g[564];
assign g[1077] = a[8] & g[565];
assign g[1588] = b[8] & g[565];
assign g[1078] = a[8] & g[566];
assign g[1589] = b[8] & g[566];
assign g[1079] = a[8] & g[567];
assign g[1590] = b[8] & g[567];
assign g[1080] = a[8] & g[568];
assign g[1591] = b[8] & g[568];
assign g[1081] = a[8] & g[569];
assign g[1592] = b[8] & g[569];
assign g[1082] = a[8] & g[570];
assign g[1593] = b[8] & g[570];
assign g[1083] = a[8] & g[571];
assign g[1594] = b[8] & g[571];
assign g[1084] = a[8] & g[572];
assign g[1595] = b[8] & g[572];
assign g[1085] = a[8] & g[573];
assign g[1596] = b[8] & g[573];
assign g[1086] = a[8] & g[574];
assign g[1597] = b[8] & g[574];
assign g[1087] = a[8] & g[575];
assign g[1598] = b[8] & g[575];
assign g[1088] = a[8] & g[576];
assign g[1599] = b[8] & g[576];
assign g[1089] = a[8] & g[577];
assign g[1600] = b[8] & g[577];
assign g[1090] = a[8] & g[578];
assign g[1601] = b[8] & g[578];
assign g[1091] = a[8] & g[579];
assign g[1602] = b[8] & g[579];
assign g[1092] = a[8] & g[580];
assign g[1603] = b[8] & g[580];
assign g[1093] = a[8] & g[581];
assign g[1604] = b[8] & g[581];
assign g[1094] = a[8] & g[582];
assign g[1605] = b[8] & g[582];
assign g[1095] = a[8] & g[583];
assign g[1606] = b[8] & g[583];
assign g[1096] = a[8] & g[584];
assign g[1607] = b[8] & g[584];
assign g[1097] = a[8] & g[585];
assign g[1608] = b[8] & g[585];
assign g[1098] = a[8] & g[586];
assign g[1609] = b[8] & g[586];
assign g[1099] = a[8] & g[587];
assign g[1610] = b[8] & g[587];
assign g[1100] = a[8] & g[588];
assign g[1611] = b[8] & g[588];
assign g[1101] = a[8] & g[589];
assign g[1612] = b[8] & g[589];
assign g[1102] = a[8] & g[590];
assign g[1613] = b[8] & g[590];
assign g[1103] = a[8] & g[591];
assign g[1614] = b[8] & g[591];
assign g[1104] = a[8] & g[592];
assign g[1615] = b[8] & g[592];
assign g[1105] = a[8] & g[593];
assign g[1616] = b[8] & g[593];
assign g[1106] = a[8] & g[594];
assign g[1617] = b[8] & g[594];
assign g[1107] = a[8] & g[595];
assign g[1618] = b[8] & g[595];
assign g[1108] = a[8] & g[596];
assign g[1619] = b[8] & g[596];
assign g[1109] = a[8] & g[597];
assign g[1620] = b[8] & g[597];
assign g[1110] = a[8] & g[598];
assign g[1621] = b[8] & g[598];
assign g[1111] = a[8] & g[599];
assign g[1622] = b[8] & g[599];
assign g[1112] = a[8] & g[600];
assign g[1623] = b[8] & g[600];
assign g[1113] = a[8] & g[601];
assign g[1624] = b[8] & g[601];
assign g[1114] = a[8] & g[602];
assign g[1625] = b[8] & g[602];
assign g[1115] = a[8] & g[603];
assign g[1626] = b[8] & g[603];
assign g[1116] = a[8] & g[604];
assign g[1627] = b[8] & g[604];
assign g[1117] = a[8] & g[605];
assign g[1628] = b[8] & g[605];
assign g[1118] = a[8] & g[606];
assign g[1629] = b[8] & g[606];
assign g[1119] = a[8] & g[607];
assign g[1630] = b[8] & g[607];
assign g[1120] = a[8] & g[608];
assign g[1631] = b[8] & g[608];
assign g[1121] = a[8] & g[609];
assign g[1632] = b[8] & g[609];
assign g[1122] = a[8] & g[610];
assign g[1633] = b[8] & g[610];
assign g[1123] = a[8] & g[611];
assign g[1634] = b[8] & g[611];
assign g[1124] = a[8] & g[612];
assign g[1635] = b[8] & g[612];
assign g[1125] = a[8] & g[613];
assign g[1636] = b[8] & g[613];
assign g[1126] = a[8] & g[614];
assign g[1637] = b[8] & g[614];
assign g[1127] = a[8] & g[615];
assign g[1638] = b[8] & g[615];
assign g[1128] = a[8] & g[616];
assign g[1639] = b[8] & g[616];
assign g[1129] = a[8] & g[617];
assign g[1640] = b[8] & g[617];
assign g[1130] = a[8] & g[618];
assign g[1641] = b[8] & g[618];
assign g[1131] = a[8] & g[619];
assign g[1642] = b[8] & g[619];
assign g[1132] = a[8] & g[620];
assign g[1643] = b[8] & g[620];
assign g[1133] = a[8] & g[621];
assign g[1644] = b[8] & g[621];
assign g[1134] = a[8] & g[622];
assign g[1645] = b[8] & g[622];
assign g[1135] = a[8] & g[623];
assign g[1646] = b[8] & g[623];
assign g[1136] = a[8] & g[624];
assign g[1647] = b[8] & g[624];
assign g[1137] = a[8] & g[625];
assign g[1648] = b[8] & g[625];
assign g[1138] = a[8] & g[626];
assign g[1649] = b[8] & g[626];
assign g[1139] = a[8] & g[627];
assign g[1650] = b[8] & g[627];
assign g[1140] = a[8] & g[628];
assign g[1651] = b[8] & g[628];
assign g[1141] = a[8] & g[629];
assign g[1652] = b[8] & g[629];
assign g[1142] = a[8] & g[630];
assign g[1653] = b[8] & g[630];
assign g[1143] = a[8] & g[631];
assign g[1654] = b[8] & g[631];
assign g[1144] = a[8] & g[632];
assign g[1655] = b[8] & g[632];
assign g[1145] = a[8] & g[633];
assign g[1656] = b[8] & g[633];
assign g[1146] = a[8] & g[634];
assign g[1657] = b[8] & g[634];
assign g[1147] = a[8] & g[635];
assign g[1658] = b[8] & g[635];
assign g[1148] = a[8] & g[636];
assign g[1659] = b[8] & g[636];
assign g[1149] = a[8] & g[637];
assign g[1660] = b[8] & g[637];
assign g[1150] = a[8] & g[638];
assign g[1661] = b[8] & g[638];
assign g[1151] = a[8] & g[639];
assign g[1662] = b[8] & g[639];
assign g[1152] = a[8] & g[640];
assign g[1663] = b[8] & g[640];
assign g[1153] = a[8] & g[641];
assign g[1664] = b[8] & g[641];
assign g[1154] = a[8] & g[642];
assign g[1665] = b[8] & g[642];
assign g[1155] = a[8] & g[643];
assign g[1666] = b[8] & g[643];
assign g[1156] = a[8] & g[644];
assign g[1667] = b[8] & g[644];
assign g[1157] = a[8] & g[645];
assign g[1668] = b[8] & g[645];
assign g[1158] = a[8] & g[646];
assign g[1669] = b[8] & g[646];
assign g[1159] = a[8] & g[647];
assign g[1670] = b[8] & g[647];
assign g[1160] = a[8] & g[648];
assign g[1671] = b[8] & g[648];
assign g[1161] = a[8] & g[649];
assign g[1672] = b[8] & g[649];
assign g[1162] = a[8] & g[650];
assign g[1673] = b[8] & g[650];
assign g[1163] = a[8] & g[651];
assign g[1674] = b[8] & g[651];
assign g[1164] = a[8] & g[652];
assign g[1675] = b[8] & g[652];
assign g[1165] = a[8] & g[653];
assign g[1676] = b[8] & g[653];
assign g[1166] = a[8] & g[654];
assign g[1677] = b[8] & g[654];
assign g[1167] = a[8] & g[655];
assign g[1678] = b[8] & g[655];
assign g[1168] = a[8] & g[656];
assign g[1679] = b[8] & g[656];
assign g[1169] = a[8] & g[657];
assign g[1680] = b[8] & g[657];
assign g[1170] = a[8] & g[658];
assign g[1681] = b[8] & g[658];
assign g[1171] = a[8] & g[659];
assign g[1682] = b[8] & g[659];
assign g[1172] = a[8] & g[660];
assign g[1683] = b[8] & g[660];
assign g[1173] = a[8] & g[661];
assign g[1684] = b[8] & g[661];
assign g[1174] = a[8] & g[662];
assign g[1685] = b[8] & g[662];
assign g[1175] = a[8] & g[663];
assign g[1686] = b[8] & g[663];
assign g[1176] = a[8] & g[664];
assign g[1687] = b[8] & g[664];
assign g[1177] = a[8] & g[665];
assign g[1688] = b[8] & g[665];
assign g[1178] = a[8] & g[666];
assign g[1689] = b[8] & g[666];
assign g[1179] = a[8] & g[667];
assign g[1690] = b[8] & g[667];
assign g[1180] = a[8] & g[668];
assign g[1691] = b[8] & g[668];
assign g[1181] = a[8] & g[669];
assign g[1692] = b[8] & g[669];
assign g[1182] = a[8] & g[670];
assign g[1693] = b[8] & g[670];
assign g[1183] = a[8] & g[671];
assign g[1694] = b[8] & g[671];
assign g[1184] = a[8] & g[672];
assign g[1695] = b[8] & g[672];
assign g[1185] = a[8] & g[673];
assign g[1696] = b[8] & g[673];
assign g[1186] = a[8] & g[674];
assign g[1697] = b[8] & g[674];
assign g[1187] = a[8] & g[675];
assign g[1698] = b[8] & g[675];
assign g[1188] = a[8] & g[676];
assign g[1699] = b[8] & g[676];
assign g[1189] = a[8] & g[677];
assign g[1700] = b[8] & g[677];
assign g[1190] = a[8] & g[678];
assign g[1701] = b[8] & g[678];
assign g[1191] = a[8] & g[679];
assign g[1702] = b[8] & g[679];
assign g[1192] = a[8] & g[680];
assign g[1703] = b[8] & g[680];
assign g[1193] = a[8] & g[681];
assign g[1704] = b[8] & g[681];
assign g[1194] = a[8] & g[682];
assign g[1705] = b[8] & g[682];
assign g[1195] = a[8] & g[683];
assign g[1706] = b[8] & g[683];
assign g[1196] = a[8] & g[684];
assign g[1707] = b[8] & g[684];
assign g[1197] = a[8] & g[685];
assign g[1708] = b[8] & g[685];
assign g[1198] = a[8] & g[686];
assign g[1709] = b[8] & g[686];
assign g[1199] = a[8] & g[687];
assign g[1710] = b[8] & g[687];
assign g[1200] = a[8] & g[688];
assign g[1711] = b[8] & g[688];
assign g[1201] = a[8] & g[689];
assign g[1712] = b[8] & g[689];
assign g[1202] = a[8] & g[690];
assign g[1713] = b[8] & g[690];
assign g[1203] = a[8] & g[691];
assign g[1714] = b[8] & g[691];
assign g[1204] = a[8] & g[692];
assign g[1715] = b[8] & g[692];
assign g[1205] = a[8] & g[693];
assign g[1716] = b[8] & g[693];
assign g[1206] = a[8] & g[694];
assign g[1717] = b[8] & g[694];
assign g[1207] = a[8] & g[695];
assign g[1718] = b[8] & g[695];
assign g[1208] = a[8] & g[696];
assign g[1719] = b[8] & g[696];
assign g[1209] = a[8] & g[697];
assign g[1720] = b[8] & g[697];
assign g[1210] = a[8] & g[698];
assign g[1721] = b[8] & g[698];
assign g[1211] = a[8] & g[699];
assign g[1722] = b[8] & g[699];
assign g[1212] = a[8] & g[700];
assign g[1723] = b[8] & g[700];
assign g[1213] = a[8] & g[701];
assign g[1724] = b[8] & g[701];
assign g[1214] = a[8] & g[702];
assign g[1725] = b[8] & g[702];
assign g[1215] = a[8] & g[703];
assign g[1726] = b[8] & g[703];
assign g[1216] = a[8] & g[704];
assign g[1727] = b[8] & g[704];
assign g[1217] = a[8] & g[705];
assign g[1728] = b[8] & g[705];
assign g[1218] = a[8] & g[706];
assign g[1729] = b[8] & g[706];
assign g[1219] = a[8] & g[707];
assign g[1730] = b[8] & g[707];
assign g[1220] = a[8] & g[708];
assign g[1731] = b[8] & g[708];
assign g[1221] = a[8] & g[709];
assign g[1732] = b[8] & g[709];
assign g[1222] = a[8] & g[710];
assign g[1733] = b[8] & g[710];
assign g[1223] = a[8] & g[711];
assign g[1734] = b[8] & g[711];
assign g[1224] = a[8] & g[712];
assign g[1735] = b[8] & g[712];
assign g[1225] = a[8] & g[713];
assign g[1736] = b[8] & g[713];
assign g[1226] = a[8] & g[714];
assign g[1737] = b[8] & g[714];
assign g[1227] = a[8] & g[715];
assign g[1738] = b[8] & g[715];
assign g[1228] = a[8] & g[716];
assign g[1739] = b[8] & g[716];
assign g[1229] = a[8] & g[717];
assign g[1740] = b[8] & g[717];
assign g[1230] = a[8] & g[718];
assign g[1741] = b[8] & g[718];
assign g[1231] = a[8] & g[719];
assign g[1742] = b[8] & g[719];
assign g[1232] = a[8] & g[720];
assign g[1743] = b[8] & g[720];
assign g[1233] = a[8] & g[721];
assign g[1744] = b[8] & g[721];
assign g[1234] = a[8] & g[722];
assign g[1745] = b[8] & g[722];
assign g[1235] = a[8] & g[723];
assign g[1746] = b[8] & g[723];
assign g[1236] = a[8] & g[724];
assign g[1747] = b[8] & g[724];
assign g[1237] = a[8] & g[725];
assign g[1748] = b[8] & g[725];
assign g[1238] = a[8] & g[726];
assign g[1749] = b[8] & g[726];
assign g[1239] = a[8] & g[727];
assign g[1750] = b[8] & g[727];
assign g[1240] = a[8] & g[728];
assign g[1751] = b[8] & g[728];
assign g[1241] = a[8] & g[729];
assign g[1752] = b[8] & g[729];
assign g[1242] = a[8] & g[730];
assign g[1753] = b[8] & g[730];
assign g[1243] = a[8] & g[731];
assign g[1754] = b[8] & g[731];
assign g[1244] = a[8] & g[732];
assign g[1755] = b[8] & g[732];
assign g[1245] = a[8] & g[733];
assign g[1756] = b[8] & g[733];
assign g[1246] = a[8] & g[734];
assign g[1757] = b[8] & g[734];
assign g[1247] = a[8] & g[735];
assign g[1758] = b[8] & g[735];
assign g[1248] = a[8] & g[736];
assign g[1759] = b[8] & g[736];
assign g[1249] = a[8] & g[737];
assign g[1760] = b[8] & g[737];
assign g[1250] = a[8] & g[738];
assign g[1761] = b[8] & g[738];
assign g[1251] = a[8] & g[739];
assign g[1762] = b[8] & g[739];
assign g[1252] = a[8] & g[740];
assign g[1763] = b[8] & g[740];
assign g[1253] = a[8] & g[741];
assign g[1764] = b[8] & g[741];
assign g[1254] = a[8] & g[742];
assign g[1765] = b[8] & g[742];
assign g[1255] = a[8] & g[743];
assign g[1766] = b[8] & g[743];
assign g[1256] = a[8] & g[744];
assign g[1767] = b[8] & g[744];
assign g[1257] = a[8] & g[745];
assign g[1768] = b[8] & g[745];
assign g[1258] = a[8] & g[746];
assign g[1769] = b[8] & g[746];
assign g[1259] = a[8] & g[747];
assign g[1770] = b[8] & g[747];
assign g[1260] = a[8] & g[748];
assign g[1771] = b[8] & g[748];
assign g[1261] = a[8] & g[749];
assign g[1772] = b[8] & g[749];
assign g[1262] = a[8] & g[750];
assign g[1773] = b[8] & g[750];
assign g[1263] = a[8] & g[751];
assign g[1774] = b[8] & g[751];
assign g[1264] = a[8] & g[752];
assign g[1775] = b[8] & g[752];
assign g[1265] = a[8] & g[753];
assign g[1776] = b[8] & g[753];
assign g[1266] = a[8] & g[754];
assign g[1777] = b[8] & g[754];
assign g[1267] = a[8] & g[755];
assign g[1778] = b[8] & g[755];
assign g[1268] = a[8] & g[756];
assign g[1779] = b[8] & g[756];
assign g[1269] = a[8] & g[757];
assign g[1780] = b[8] & g[757];
assign g[1270] = a[8] & g[758];
assign g[1781] = b[8] & g[758];
assign g[1271] = a[8] & g[759];
assign g[1782] = b[8] & g[759];
assign g[1272] = a[8] & g[760];
assign g[1783] = b[8] & g[760];
assign g[1273] = a[8] & g[761];
assign g[1784] = b[8] & g[761];
assign g[1274] = a[8] & g[762];
assign g[1785] = b[8] & g[762];
assign g[1275] = a[8] & g[763];
assign g[1786] = b[8] & g[763];
assign g[1276] = a[8] & g[764];
assign g[1787] = b[8] & g[764];
assign g[1277] = a[8] & g[765];
assign g[1788] = b[8] & g[765];
assign g[1278] = a[8] & g[766];
assign g[1789] = b[8] & g[766];
assign g[1279] = a[8] & g[767];
assign g[1790] = b[8] & g[767];
assign g[1280] = a[8] & g[768];
assign g[1791] = b[8] & g[768];
assign g[1281] = a[8] & g[769];
assign g[1792] = b[8] & g[769];
assign g[1282] = a[8] & g[770];
assign g[1793] = b[8] & g[770];
assign g[1283] = a[8] & g[771];
assign g[1794] = b[8] & g[771];
assign g[1284] = a[8] & g[772];
assign g[1795] = b[8] & g[772];
assign g[1285] = a[8] & g[773];
assign g[1796] = b[8] & g[773];
assign g[1286] = a[8] & g[774];
assign g[1797] = b[8] & g[774];
assign g[1287] = a[8] & g[775];
assign g[1798] = b[8] & g[775];
assign g[1288] = a[8] & g[776];
assign g[1799] = b[8] & g[776];
assign g[1289] = a[8] & g[777];
assign g[1800] = b[8] & g[777];
assign g[1290] = a[8] & g[778];
assign g[1801] = b[8] & g[778];
assign g[1291] = a[8] & g[779];
assign g[1802] = b[8] & g[779];
assign g[1292] = a[8] & g[780];
assign g[1803] = b[8] & g[780];
assign g[1293] = a[8] & g[781];
assign g[1804] = b[8] & g[781];
assign g[1294] = a[8] & g[782];
assign g[1805] = b[8] & g[782];
assign g[1295] = a[8] & g[783];
assign g[1806] = b[8] & g[783];
assign g[1296] = a[8] & g[784];
assign g[1807] = b[8] & g[784];
assign g[1297] = a[8] & g[785];
assign g[1808] = b[8] & g[785];
assign g[1298] = a[8] & g[786];
assign g[1809] = b[8] & g[786];
assign g[1299] = a[8] & g[787];
assign g[1810] = b[8] & g[787];
assign g[1300] = a[8] & g[788];
assign g[1811] = b[8] & g[788];
assign g[1301] = a[8] & g[789];
assign g[1812] = b[8] & g[789];
assign g[1302] = a[8] & g[790];
assign g[1813] = b[8] & g[790];
assign g[1303] = a[8] & g[791];
assign g[1814] = b[8] & g[791];
assign g[1304] = a[8] & g[792];
assign g[1815] = b[8] & g[792];
assign g[1305] = a[8] & g[793];
assign g[1816] = b[8] & g[793];
assign g[1306] = a[8] & g[794];
assign g[1817] = b[8] & g[794];
assign g[1307] = a[8] & g[795];
assign g[1818] = b[8] & g[795];
assign g[1308] = a[8] & g[796];
assign g[1819] = b[8] & g[796];
assign g[1309] = a[8] & g[797];
assign g[1820] = b[8] & g[797];
assign g[1310] = a[8] & g[798];
assign g[1821] = b[8] & g[798];
assign g[1311] = a[8] & g[799];
assign g[1822] = b[8] & g[799];
assign g[1312] = a[8] & g[800];
assign g[1823] = b[8] & g[800];
assign g[1313] = a[8] & g[801];
assign g[1824] = b[8] & g[801];
assign g[1314] = a[8] & g[802];
assign g[1825] = b[8] & g[802];
assign g[1315] = a[8] & g[803];
assign g[1826] = b[8] & g[803];
assign g[1316] = a[8] & g[804];
assign g[1827] = b[8] & g[804];
assign g[1317] = a[8] & g[805];
assign g[1828] = b[8] & g[805];
assign g[1318] = a[8] & g[806];
assign g[1829] = b[8] & g[806];
assign g[1319] = a[8] & g[807];
assign g[1830] = b[8] & g[807];
assign g[1320] = a[8] & g[808];
assign g[1831] = b[8] & g[808];
assign g[1321] = a[8] & g[809];
assign g[1832] = b[8] & g[809];
assign g[1322] = a[8] & g[810];
assign g[1833] = b[8] & g[810];
assign g[1323] = a[8] & g[811];
assign g[1834] = b[8] & g[811];
assign g[1324] = a[8] & g[812];
assign g[1835] = b[8] & g[812];
assign g[1325] = a[8] & g[813];
assign g[1836] = b[8] & g[813];
assign g[1326] = a[8] & g[814];
assign g[1837] = b[8] & g[814];
assign g[1327] = a[8] & g[815];
assign g[1838] = b[8] & g[815];
assign g[1328] = a[8] & g[816];
assign g[1839] = b[8] & g[816];
assign g[1329] = a[8] & g[817];
assign g[1840] = b[8] & g[817];
assign g[1330] = a[8] & g[818];
assign g[1841] = b[8] & g[818];
assign g[1331] = a[8] & g[819];
assign g[1842] = b[8] & g[819];
assign g[1332] = a[8] & g[820];
assign g[1843] = b[8] & g[820];
assign g[1333] = a[8] & g[821];
assign g[1844] = b[8] & g[821];
assign g[1334] = a[8] & g[822];
assign g[1845] = b[8] & g[822];
assign g[1335] = a[8] & g[823];
assign g[1846] = b[8] & g[823];
assign g[1336] = a[8] & g[824];
assign g[1847] = b[8] & g[824];
assign g[1337] = a[8] & g[825];
assign g[1848] = b[8] & g[825];
assign g[1338] = a[8] & g[826];
assign g[1849] = b[8] & g[826];
assign g[1339] = a[8] & g[827];
assign g[1850] = b[8] & g[827];
assign g[1340] = a[8] & g[828];
assign g[1851] = b[8] & g[828];
assign g[1341] = a[8] & g[829];
assign g[1852] = b[8] & g[829];
assign g[1342] = a[8] & g[830];
assign g[1853] = b[8] & g[830];
assign g[1343] = a[8] & g[831];
assign g[1854] = b[8] & g[831];
assign g[1344] = a[8] & g[832];
assign g[1855] = b[8] & g[832];
assign g[1345] = a[8] & g[833];
assign g[1856] = b[8] & g[833];
assign g[1346] = a[8] & g[834];
assign g[1857] = b[8] & g[834];
assign g[1347] = a[8] & g[835];
assign g[1858] = b[8] & g[835];
assign g[1348] = a[8] & g[836];
assign g[1859] = b[8] & g[836];
assign g[1349] = a[8] & g[837];
assign g[1860] = b[8] & g[837];
assign g[1350] = a[8] & g[838];
assign g[1861] = b[8] & g[838];
assign g[1351] = a[8] & g[839];
assign g[1862] = b[8] & g[839];
assign g[1352] = a[8] & g[840];
assign g[1863] = b[8] & g[840];
assign g[1353] = a[8] & g[841];
assign g[1864] = b[8] & g[841];
assign g[1354] = a[8] & g[842];
assign g[1865] = b[8] & g[842];
assign g[1355] = a[8] & g[843];
assign g[1866] = b[8] & g[843];
assign g[1356] = a[8] & g[844];
assign g[1867] = b[8] & g[844];
assign g[1357] = a[8] & g[845];
assign g[1868] = b[8] & g[845];
assign g[1358] = a[8] & g[846];
assign g[1869] = b[8] & g[846];
assign g[1359] = a[8] & g[847];
assign g[1870] = b[8] & g[847];
assign g[1360] = a[8] & g[848];
assign g[1871] = b[8] & g[848];
assign g[1361] = a[8] & g[849];
assign g[1872] = b[8] & g[849];
assign g[1362] = a[8] & g[850];
assign g[1873] = b[8] & g[850];
assign g[1363] = a[8] & g[851];
assign g[1874] = b[8] & g[851];
assign g[1364] = a[8] & g[852];
assign g[1875] = b[8] & g[852];
assign g[1365] = a[8] & g[853];
assign g[1876] = b[8] & g[853];
assign g[1366] = a[8] & g[854];
assign g[1877] = b[8] & g[854];
assign g[1367] = a[8] & g[855];
assign g[1878] = b[8] & g[855];
assign g[1368] = a[8] & g[856];
assign g[1879] = b[8] & g[856];
assign g[1369] = a[8] & g[857];
assign g[1880] = b[8] & g[857];
assign g[1370] = a[8] & g[858];
assign g[1881] = b[8] & g[858];
assign g[1371] = a[8] & g[859];
assign g[1882] = b[8] & g[859];
assign g[1372] = a[8] & g[860];
assign g[1883] = b[8] & g[860];
assign g[1373] = a[8] & g[861];
assign g[1884] = b[8] & g[861];
assign g[1374] = a[8] & g[862];
assign g[1885] = b[8] & g[862];
assign g[1375] = a[8] & g[863];
assign g[1886] = b[8] & g[863];
assign g[1376] = a[8] & g[864];
assign g[1887] = b[8] & g[864];
assign g[1377] = a[8] & g[865];
assign g[1888] = b[8] & g[865];
assign g[1378] = a[8] & g[866];
assign g[1889] = b[8] & g[866];
assign g[1379] = a[8] & g[867];
assign g[1890] = b[8] & g[867];
assign g[1380] = a[8] & g[868];
assign g[1891] = b[8] & g[868];
assign g[1381] = a[8] & g[869];
assign g[1892] = b[8] & g[869];
assign g[1382] = a[8] & g[870];
assign g[1893] = b[8] & g[870];
assign g[1383] = a[8] & g[871];
assign g[1894] = b[8] & g[871];
assign g[1384] = a[8] & g[872];
assign g[1895] = b[8] & g[872];
assign g[1385] = a[8] & g[873];
assign g[1896] = b[8] & g[873];
assign g[1386] = a[8] & g[874];
assign g[1897] = b[8] & g[874];
assign g[1387] = a[8] & g[875];
assign g[1898] = b[8] & g[875];
assign g[1388] = a[8] & g[876];
assign g[1899] = b[8] & g[876];
assign g[1389] = a[8] & g[877];
assign g[1900] = b[8] & g[877];
assign g[1390] = a[8] & g[878];
assign g[1901] = b[8] & g[878];
assign g[1391] = a[8] & g[879];
assign g[1902] = b[8] & g[879];
assign g[1392] = a[8] & g[880];
assign g[1903] = b[8] & g[880];
assign g[1393] = a[8] & g[881];
assign g[1904] = b[8] & g[881];
assign g[1394] = a[8] & g[882];
assign g[1905] = b[8] & g[882];
assign g[1395] = a[8] & g[883];
assign g[1906] = b[8] & g[883];
assign g[1396] = a[8] & g[884];
assign g[1907] = b[8] & g[884];
assign g[1397] = a[8] & g[885];
assign g[1908] = b[8] & g[885];
assign g[1398] = a[8] & g[886];
assign g[1909] = b[8] & g[886];
assign g[1399] = a[8] & g[887];
assign g[1910] = b[8] & g[887];
assign g[1400] = a[8] & g[888];
assign g[1911] = b[8] & g[888];
assign g[1401] = a[8] & g[889];
assign g[1912] = b[8] & g[889];
assign g[1402] = a[8] & g[890];
assign g[1913] = b[8] & g[890];
assign g[1403] = a[8] & g[891];
assign g[1914] = b[8] & g[891];
assign g[1404] = a[8] & g[892];
assign g[1915] = b[8] & g[892];
assign g[1405] = a[8] & g[893];
assign g[1916] = b[8] & g[893];
assign g[1406] = a[8] & g[894];
assign g[1917] = b[8] & g[894];
assign g[1407] = a[8] & g[895];
assign g[1918] = b[8] & g[895];
assign g[1408] = a[8] & g[896];
assign g[1919] = b[8] & g[896];
assign g[1409] = a[8] & g[897];
assign g[1920] = b[8] & g[897];
assign g[1410] = a[8] & g[898];
assign g[1921] = b[8] & g[898];
assign g[1411] = a[8] & g[899];
assign g[1922] = b[8] & g[899];
assign g[1412] = a[8] & g[900];
assign g[1923] = b[8] & g[900];
assign g[1413] = a[8] & g[901];
assign g[1924] = b[8] & g[901];
assign g[1414] = a[8] & g[902];
assign g[1925] = b[8] & g[902];
assign g[1415] = a[8] & g[903];
assign g[1926] = b[8] & g[903];
assign g[1416] = a[8] & g[904];
assign g[1927] = b[8] & g[904];
assign g[1417] = a[8] & g[905];
assign g[1928] = b[8] & g[905];
assign g[1418] = a[8] & g[906];
assign g[1929] = b[8] & g[906];
assign g[1419] = a[8] & g[907];
assign g[1930] = b[8] & g[907];
assign g[1420] = a[8] & g[908];
assign g[1931] = b[8] & g[908];
assign g[1421] = a[8] & g[909];
assign g[1932] = b[8] & g[909];
assign g[1422] = a[8] & g[910];
assign g[1933] = b[8] & g[910];
assign g[1423] = a[8] & g[911];
assign g[1934] = b[8] & g[911];
assign g[1424] = a[8] & g[912];
assign g[1935] = b[8] & g[912];
assign g[1425] = a[8] & g[913];
assign g[1936] = b[8] & g[913];
assign g[1426] = a[8] & g[914];
assign g[1937] = b[8] & g[914];
assign g[1427] = a[8] & g[915];
assign g[1938] = b[8] & g[915];
assign g[1428] = a[8] & g[916];
assign g[1939] = b[8] & g[916];
assign g[1429] = a[8] & g[917];
assign g[1940] = b[8] & g[917];
assign g[1430] = a[8] & g[918];
assign g[1941] = b[8] & g[918];
assign g[1431] = a[8] & g[919];
assign g[1942] = b[8] & g[919];
assign g[1432] = a[8] & g[920];
assign g[1943] = b[8] & g[920];
assign g[1433] = a[8] & g[921];
assign g[1944] = b[8] & g[921];
assign g[1434] = a[8] & g[922];
assign g[1945] = b[8] & g[922];
assign g[1435] = a[8] & g[923];
assign g[1946] = b[8] & g[923];
assign g[1436] = a[8] & g[924];
assign g[1947] = b[8] & g[924];
assign g[1437] = a[8] & g[925];
assign g[1948] = b[8] & g[925];
assign g[1438] = a[8] & g[926];
assign g[1949] = b[8] & g[926];
assign g[1439] = a[8] & g[927];
assign g[1950] = b[8] & g[927];
assign g[1440] = a[8] & g[928];
assign g[1951] = b[8] & g[928];
assign g[1441] = a[8] & g[929];
assign g[1952] = b[8] & g[929];
assign g[1442] = a[8] & g[930];
assign g[1953] = b[8] & g[930];
assign g[1443] = a[8] & g[931];
assign g[1954] = b[8] & g[931];
assign g[1444] = a[8] & g[932];
assign g[1955] = b[8] & g[932];
assign g[1445] = a[8] & g[933];
assign g[1956] = b[8] & g[933];
assign g[1446] = a[8] & g[934];
assign g[1957] = b[8] & g[934];
assign g[1447] = a[8] & g[935];
assign g[1958] = b[8] & g[935];
assign g[1448] = a[8] & g[936];
assign g[1959] = b[8] & g[936];
assign g[1449] = a[8] & g[937];
assign g[1960] = b[8] & g[937];
assign g[1450] = a[8] & g[938];
assign g[1961] = b[8] & g[938];
assign g[1451] = a[8] & g[939];
assign g[1962] = b[8] & g[939];
assign g[1452] = a[8] & g[940];
assign g[1963] = b[8] & g[940];
assign g[1453] = a[8] & g[941];
assign g[1964] = b[8] & g[941];
assign g[1454] = a[8] & g[942];
assign g[1965] = b[8] & g[942];
assign g[1455] = a[8] & g[943];
assign g[1966] = b[8] & g[943];
assign g[1456] = a[8] & g[944];
assign g[1967] = b[8] & g[944];
assign g[1457] = a[8] & g[945];
assign g[1968] = b[8] & g[945];
assign g[1458] = a[8] & g[946];
assign g[1969] = b[8] & g[946];
assign g[1459] = a[8] & g[947];
assign g[1970] = b[8] & g[947];
assign g[1460] = a[8] & g[948];
assign g[1971] = b[8] & g[948];
assign g[1461] = a[8] & g[949];
assign g[1972] = b[8] & g[949];
assign g[1462] = a[8] & g[950];
assign g[1973] = b[8] & g[950];
assign g[1463] = a[8] & g[951];
assign g[1974] = b[8] & g[951];
assign g[1464] = a[8] & g[952];
assign g[1975] = b[8] & g[952];
assign g[1465] = a[8] & g[953];
assign g[1976] = b[8] & g[953];
assign g[1466] = a[8] & g[954];
assign g[1977] = b[8] & g[954];
assign g[1467] = a[8] & g[955];
assign g[1978] = b[8] & g[955];
assign g[1468] = a[8] & g[956];
assign g[1979] = b[8] & g[956];
assign g[1469] = a[8] & g[957];
assign g[1980] = b[8] & g[957];
assign g[1470] = a[8] & g[958];
assign g[1981] = b[8] & g[958];
assign g[1471] = a[8] & g[959];
assign g[1982] = b[8] & g[959];
assign g[1472] = a[8] & g[960];
assign g[1983] = b[8] & g[960];
assign g[1473] = a[8] & g[961];
assign g[1984] = b[8] & g[961];
assign g[1474] = a[8] & g[962];
assign g[1985] = b[8] & g[962];
assign g[1475] = a[8] & g[963];
assign g[1986] = b[8] & g[963];
assign g[1476] = a[8] & g[964];
assign g[1987] = b[8] & g[964];
assign g[1477] = a[8] & g[965];
assign g[1988] = b[8] & g[965];
assign g[1478] = a[8] & g[966];
assign g[1989] = b[8] & g[966];
assign g[1479] = a[8] & g[967];
assign g[1990] = b[8] & g[967];
assign g[1480] = a[8] & g[968];
assign g[1991] = b[8] & g[968];
assign g[1481] = a[8] & g[969];
assign g[1992] = b[8] & g[969];
assign g[1482] = a[8] & g[970];
assign g[1993] = b[8] & g[970];
assign g[1483] = a[8] & g[971];
assign g[1994] = b[8] & g[971];
assign g[1484] = a[8] & g[972];
assign g[1995] = b[8] & g[972];
assign g[1485] = a[8] & g[973];
assign g[1996] = b[8] & g[973];
assign g[1486] = a[8] & g[974];
assign g[1997] = b[8] & g[974];
assign g[1487] = a[8] & g[975];
assign g[1998] = b[8] & g[975];
assign g[1488] = a[8] & g[976];
assign g[1999] = b[8] & g[976];
assign g[1489] = a[8] & g[977];
assign g[2000] = b[8] & g[977];
assign g[1490] = a[8] & g[978];
assign g[2001] = b[8] & g[978];
assign g[1491] = a[8] & g[979];
assign g[2002] = b[8] & g[979];
assign g[1492] = a[8] & g[980];
assign g[2003] = b[8] & g[980];
assign g[1493] = a[8] & g[981];
assign g[2004] = b[8] & g[981];
assign g[1494] = a[8] & g[982];
assign g[2005] = b[8] & g[982];
assign g[1495] = a[8] & g[983];
assign g[2006] = b[8] & g[983];
assign g[1496] = a[8] & g[984];
assign g[2007] = b[8] & g[984];
assign g[1497] = a[8] & g[985];
assign g[2008] = b[8] & g[985];
assign g[1498] = a[8] & g[986];
assign g[2009] = b[8] & g[986];
assign g[1499] = a[8] & g[987];
assign g[2010] = b[8] & g[987];
assign g[1500] = a[8] & g[988];
assign g[2011] = b[8] & g[988];
assign g[1501] = a[8] & g[989];
assign g[2012] = b[8] & g[989];
assign g[1502] = a[8] & g[990];
assign g[2013] = b[8] & g[990];
assign g[1503] = a[8] & g[991];
assign g[2014] = b[8] & g[991];
assign g[1504] = a[8] & g[992];
assign g[2015] = b[8] & g[992];
assign g[1505] = a[8] & g[993];
assign g[2016] = b[8] & g[993];
assign g[1506] = a[8] & g[994];
assign g[2017] = b[8] & g[994];
assign g[1507] = a[8] & g[995];
assign g[2018] = b[8] & g[995];
assign g[1508] = a[8] & g[996];
assign g[2019] = b[8] & g[996];
assign g[1509] = a[8] & g[997];
assign g[2020] = b[8] & g[997];
assign g[1510] = a[8] & g[998];
assign g[2021] = b[8] & g[998];
assign g[1511] = a[8] & g[999];
assign g[2022] = b[8] & g[999];
assign g[1512] = a[8] & g[1000];
assign g[2023] = b[8] & g[1000];
assign g[1513] = a[8] & g[1001];
assign g[2024] = b[8] & g[1001];
assign g[1514] = a[8] & g[1002];
assign g[2025] = b[8] & g[1002];
assign g[1515] = a[8] & g[1003];
assign g[2026] = b[8] & g[1003];
assign g[1516] = a[8] & g[1004];
assign g[2027] = b[8] & g[1004];
assign g[1517] = a[8] & g[1005];
assign g[2028] = b[8] & g[1005];
assign g[1518] = a[8] & g[1006];
assign g[2029] = b[8] & g[1006];
assign g[1519] = a[8] & g[1007];
assign g[2030] = b[8] & g[1007];
assign g[1520] = a[8] & g[1008];
assign g[2031] = b[8] & g[1008];
assign g[1521] = a[8] & g[1009];
assign g[2032] = b[8] & g[1009];
assign g[1522] = a[8] & g[1010];
assign g[2033] = b[8] & g[1010];
assign g[1523] = a[8] & g[1011];
assign g[2034] = b[8] & g[1011];
assign g[1524] = a[8] & g[1012];
assign g[2035] = b[8] & g[1012];
//Assigning outputs for input bit 9
assign g[2036] = a[9] & b[9];
assign g[2037] = a[9] & g[1013];
assign g[3060] = b[9] & g[1013];
assign g[2038] = a[9] & g[1014];
assign g[3061] = b[9] & g[1014];
assign g[2039] = a[9] & g[1015];
assign g[3062] = b[9] & g[1015];
assign g[2040] = a[9] & g[1016];
assign g[3063] = b[9] & g[1016];
assign g[2041] = a[9] & g[1017];
assign g[3064] = b[9] & g[1017];
assign g[2042] = a[9] & g[1018];
assign g[3065] = b[9] & g[1018];
assign g[2043] = a[9] & g[1019];
assign g[3066] = b[9] & g[1019];
assign g[2044] = a[9] & g[1020];
assign g[3067] = b[9] & g[1020];
assign g[2045] = a[9] & g[1021];
assign g[3068] = b[9] & g[1021];
assign g[2046] = a[9] & g[1022];
assign g[3069] = b[9] & g[1022];
assign g[2047] = a[9] & g[1023];
assign g[3070] = b[9] & g[1023];
assign g[2048] = a[9] & g[1024];
assign g[3071] = b[9] & g[1024];
assign g[2049] = a[9] & g[1025];
assign g[3072] = b[9] & g[1025];
assign g[2050] = a[9] & g[1026];
assign g[3073] = b[9] & g[1026];
assign g[2051] = a[9] & g[1027];
assign g[3074] = b[9] & g[1027];
assign g[2052] = a[9] & g[1028];
assign g[3075] = b[9] & g[1028];
assign g[2053] = a[9] & g[1029];
assign g[3076] = b[9] & g[1029];
assign g[2054] = a[9] & g[1030];
assign g[3077] = b[9] & g[1030];
assign g[2055] = a[9] & g[1031];
assign g[3078] = b[9] & g[1031];
assign g[2056] = a[9] & g[1032];
assign g[3079] = b[9] & g[1032];
assign g[2057] = a[9] & g[1033];
assign g[3080] = b[9] & g[1033];
assign g[2058] = a[9] & g[1034];
assign g[3081] = b[9] & g[1034];
assign g[2059] = a[9] & g[1035];
assign g[3082] = b[9] & g[1035];
assign g[2060] = a[9] & g[1036];
assign g[3083] = b[9] & g[1036];
assign g[2061] = a[9] & g[1037];
assign g[3084] = b[9] & g[1037];
assign g[2062] = a[9] & g[1038];
assign g[3085] = b[9] & g[1038];
assign g[2063] = a[9] & g[1039];
assign g[3086] = b[9] & g[1039];
assign g[2064] = a[9] & g[1040];
assign g[3087] = b[9] & g[1040];
assign g[2065] = a[9] & g[1041];
assign g[3088] = b[9] & g[1041];
assign g[2066] = a[9] & g[1042];
assign g[3089] = b[9] & g[1042];
assign g[2067] = a[9] & g[1043];
assign g[3090] = b[9] & g[1043];
assign g[2068] = a[9] & g[1044];
assign g[3091] = b[9] & g[1044];
assign g[2069] = a[9] & g[1045];
assign g[3092] = b[9] & g[1045];
assign g[2070] = a[9] & g[1046];
assign g[3093] = b[9] & g[1046];
assign g[2071] = a[9] & g[1047];
assign g[3094] = b[9] & g[1047];
assign g[2072] = a[9] & g[1048];
assign g[3095] = b[9] & g[1048];
assign g[2073] = a[9] & g[1049];
assign g[3096] = b[9] & g[1049];
assign g[2074] = a[9] & g[1050];
assign g[3097] = b[9] & g[1050];
assign g[2075] = a[9] & g[1051];
assign g[3098] = b[9] & g[1051];
assign g[2076] = a[9] & g[1052];
assign g[3099] = b[9] & g[1052];
assign g[2077] = a[9] & g[1053];
assign g[3100] = b[9] & g[1053];
assign g[2078] = a[9] & g[1054];
assign g[3101] = b[9] & g[1054];
assign g[2079] = a[9] & g[1055];
assign g[3102] = b[9] & g[1055];
assign g[2080] = a[9] & g[1056];
assign g[3103] = b[9] & g[1056];
assign g[2081] = a[9] & g[1057];
assign g[3104] = b[9] & g[1057];
assign g[2082] = a[9] & g[1058];
assign g[3105] = b[9] & g[1058];
assign g[2083] = a[9] & g[1059];
assign g[3106] = b[9] & g[1059];
assign g[2084] = a[9] & g[1060];
assign g[3107] = b[9] & g[1060];
assign g[2085] = a[9] & g[1061];
assign g[3108] = b[9] & g[1061];
assign g[2086] = a[9] & g[1062];
assign g[3109] = b[9] & g[1062];
assign g[2087] = a[9] & g[1063];
assign g[3110] = b[9] & g[1063];
assign g[2088] = a[9] & g[1064];
assign g[3111] = b[9] & g[1064];
assign g[2089] = a[9] & g[1065];
assign g[3112] = b[9] & g[1065];
assign g[2090] = a[9] & g[1066];
assign g[3113] = b[9] & g[1066];
assign g[2091] = a[9] & g[1067];
assign g[3114] = b[9] & g[1067];
assign g[2092] = a[9] & g[1068];
assign g[3115] = b[9] & g[1068];
assign g[2093] = a[9] & g[1069];
assign g[3116] = b[9] & g[1069];
assign g[2094] = a[9] & g[1070];
assign g[3117] = b[9] & g[1070];
assign g[2095] = a[9] & g[1071];
assign g[3118] = b[9] & g[1071];
assign g[2096] = a[9] & g[1072];
assign g[3119] = b[9] & g[1072];
assign g[2097] = a[9] & g[1073];
assign g[3120] = b[9] & g[1073];
assign g[2098] = a[9] & g[1074];
assign g[3121] = b[9] & g[1074];
assign g[2099] = a[9] & g[1075];
assign g[3122] = b[9] & g[1075];
assign g[2100] = a[9] & g[1076];
assign g[3123] = b[9] & g[1076];
assign g[2101] = a[9] & g[1077];
assign g[3124] = b[9] & g[1077];
assign g[2102] = a[9] & g[1078];
assign g[3125] = b[9] & g[1078];
assign g[2103] = a[9] & g[1079];
assign g[3126] = b[9] & g[1079];
assign g[2104] = a[9] & g[1080];
assign g[3127] = b[9] & g[1080];
assign g[2105] = a[9] & g[1081];
assign g[3128] = b[9] & g[1081];
assign g[2106] = a[9] & g[1082];
assign g[3129] = b[9] & g[1082];
assign g[2107] = a[9] & g[1083];
assign g[3130] = b[9] & g[1083];
assign g[2108] = a[9] & g[1084];
assign g[3131] = b[9] & g[1084];
assign g[2109] = a[9] & g[1085];
assign g[3132] = b[9] & g[1085];
assign g[2110] = a[9] & g[1086];
assign g[3133] = b[9] & g[1086];
assign g[2111] = a[9] & g[1087];
assign g[3134] = b[9] & g[1087];
assign g[2112] = a[9] & g[1088];
assign g[3135] = b[9] & g[1088];
assign g[2113] = a[9] & g[1089];
assign g[3136] = b[9] & g[1089];
assign g[2114] = a[9] & g[1090];
assign g[3137] = b[9] & g[1090];
assign g[2115] = a[9] & g[1091];
assign g[3138] = b[9] & g[1091];
assign g[2116] = a[9] & g[1092];
assign g[3139] = b[9] & g[1092];
assign g[2117] = a[9] & g[1093];
assign g[3140] = b[9] & g[1093];
assign g[2118] = a[9] & g[1094];
assign g[3141] = b[9] & g[1094];
assign g[2119] = a[9] & g[1095];
assign g[3142] = b[9] & g[1095];
assign g[2120] = a[9] & g[1096];
assign g[3143] = b[9] & g[1096];
assign g[2121] = a[9] & g[1097];
assign g[3144] = b[9] & g[1097];
assign g[2122] = a[9] & g[1098];
assign g[3145] = b[9] & g[1098];
assign g[2123] = a[9] & g[1099];
assign g[3146] = b[9] & g[1099];
assign g[2124] = a[9] & g[1100];
assign g[3147] = b[9] & g[1100];
assign g[2125] = a[9] & g[1101];
assign g[3148] = b[9] & g[1101];
assign g[2126] = a[9] & g[1102];
assign g[3149] = b[9] & g[1102];
assign g[2127] = a[9] & g[1103];
assign g[3150] = b[9] & g[1103];
assign g[2128] = a[9] & g[1104];
assign g[3151] = b[9] & g[1104];
assign g[2129] = a[9] & g[1105];
assign g[3152] = b[9] & g[1105];
assign g[2130] = a[9] & g[1106];
assign g[3153] = b[9] & g[1106];
assign g[2131] = a[9] & g[1107];
assign g[3154] = b[9] & g[1107];
assign g[2132] = a[9] & g[1108];
assign g[3155] = b[9] & g[1108];
assign g[2133] = a[9] & g[1109];
assign g[3156] = b[9] & g[1109];
assign g[2134] = a[9] & g[1110];
assign g[3157] = b[9] & g[1110];
assign g[2135] = a[9] & g[1111];
assign g[3158] = b[9] & g[1111];
assign g[2136] = a[9] & g[1112];
assign g[3159] = b[9] & g[1112];
assign g[2137] = a[9] & g[1113];
assign g[3160] = b[9] & g[1113];
assign g[2138] = a[9] & g[1114];
assign g[3161] = b[9] & g[1114];
assign g[2139] = a[9] & g[1115];
assign g[3162] = b[9] & g[1115];
assign g[2140] = a[9] & g[1116];
assign g[3163] = b[9] & g[1116];
assign g[2141] = a[9] & g[1117];
assign g[3164] = b[9] & g[1117];
assign g[2142] = a[9] & g[1118];
assign g[3165] = b[9] & g[1118];
assign g[2143] = a[9] & g[1119];
assign g[3166] = b[9] & g[1119];
assign g[2144] = a[9] & g[1120];
assign g[3167] = b[9] & g[1120];
assign g[2145] = a[9] & g[1121];
assign g[3168] = b[9] & g[1121];
assign g[2146] = a[9] & g[1122];
assign g[3169] = b[9] & g[1122];
assign g[2147] = a[9] & g[1123];
assign g[3170] = b[9] & g[1123];
assign g[2148] = a[9] & g[1124];
assign g[3171] = b[9] & g[1124];
assign g[2149] = a[9] & g[1125];
assign g[3172] = b[9] & g[1125];
assign g[2150] = a[9] & g[1126];
assign g[3173] = b[9] & g[1126];
assign g[2151] = a[9] & g[1127];
assign g[3174] = b[9] & g[1127];
assign g[2152] = a[9] & g[1128];
assign g[3175] = b[9] & g[1128];
assign g[2153] = a[9] & g[1129];
assign g[3176] = b[9] & g[1129];
assign g[2154] = a[9] & g[1130];
assign g[3177] = b[9] & g[1130];
assign g[2155] = a[9] & g[1131];
assign g[3178] = b[9] & g[1131];
assign g[2156] = a[9] & g[1132];
assign g[3179] = b[9] & g[1132];
assign g[2157] = a[9] & g[1133];
assign g[3180] = b[9] & g[1133];
assign g[2158] = a[9] & g[1134];
assign g[3181] = b[9] & g[1134];
assign g[2159] = a[9] & g[1135];
assign g[3182] = b[9] & g[1135];
assign g[2160] = a[9] & g[1136];
assign g[3183] = b[9] & g[1136];
assign g[2161] = a[9] & g[1137];
assign g[3184] = b[9] & g[1137];
assign g[2162] = a[9] & g[1138];
assign g[3185] = b[9] & g[1138];
assign g[2163] = a[9] & g[1139];
assign g[3186] = b[9] & g[1139];
assign g[2164] = a[9] & g[1140];
assign g[3187] = b[9] & g[1140];
assign g[2165] = a[9] & g[1141];
assign g[3188] = b[9] & g[1141];
assign g[2166] = a[9] & g[1142];
assign g[3189] = b[9] & g[1142];
assign g[2167] = a[9] & g[1143];
assign g[3190] = b[9] & g[1143];
assign g[2168] = a[9] & g[1144];
assign g[3191] = b[9] & g[1144];
assign g[2169] = a[9] & g[1145];
assign g[3192] = b[9] & g[1145];
assign g[2170] = a[9] & g[1146];
assign g[3193] = b[9] & g[1146];
assign g[2171] = a[9] & g[1147];
assign g[3194] = b[9] & g[1147];
assign g[2172] = a[9] & g[1148];
assign g[3195] = b[9] & g[1148];
assign g[2173] = a[9] & g[1149];
assign g[3196] = b[9] & g[1149];
assign g[2174] = a[9] & g[1150];
assign g[3197] = b[9] & g[1150];
assign g[2175] = a[9] & g[1151];
assign g[3198] = b[9] & g[1151];
assign g[2176] = a[9] & g[1152];
assign g[3199] = b[9] & g[1152];
assign g[2177] = a[9] & g[1153];
assign g[3200] = b[9] & g[1153];
assign g[2178] = a[9] & g[1154];
assign g[3201] = b[9] & g[1154];
assign g[2179] = a[9] & g[1155];
assign g[3202] = b[9] & g[1155];
assign g[2180] = a[9] & g[1156];
assign g[3203] = b[9] & g[1156];
assign g[2181] = a[9] & g[1157];
assign g[3204] = b[9] & g[1157];
assign g[2182] = a[9] & g[1158];
assign g[3205] = b[9] & g[1158];
assign g[2183] = a[9] & g[1159];
assign g[3206] = b[9] & g[1159];
assign g[2184] = a[9] & g[1160];
assign g[3207] = b[9] & g[1160];
assign g[2185] = a[9] & g[1161];
assign g[3208] = b[9] & g[1161];
assign g[2186] = a[9] & g[1162];
assign g[3209] = b[9] & g[1162];
assign g[2187] = a[9] & g[1163];
assign g[3210] = b[9] & g[1163];
assign g[2188] = a[9] & g[1164];
assign g[3211] = b[9] & g[1164];
assign g[2189] = a[9] & g[1165];
assign g[3212] = b[9] & g[1165];
assign g[2190] = a[9] & g[1166];
assign g[3213] = b[9] & g[1166];
assign g[2191] = a[9] & g[1167];
assign g[3214] = b[9] & g[1167];
assign g[2192] = a[9] & g[1168];
assign g[3215] = b[9] & g[1168];
assign g[2193] = a[9] & g[1169];
assign g[3216] = b[9] & g[1169];
assign g[2194] = a[9] & g[1170];
assign g[3217] = b[9] & g[1170];
assign g[2195] = a[9] & g[1171];
assign g[3218] = b[9] & g[1171];
assign g[2196] = a[9] & g[1172];
assign g[3219] = b[9] & g[1172];
assign g[2197] = a[9] & g[1173];
assign g[3220] = b[9] & g[1173];
assign g[2198] = a[9] & g[1174];
assign g[3221] = b[9] & g[1174];
assign g[2199] = a[9] & g[1175];
assign g[3222] = b[9] & g[1175];
assign g[2200] = a[9] & g[1176];
assign g[3223] = b[9] & g[1176];
assign g[2201] = a[9] & g[1177];
assign g[3224] = b[9] & g[1177];
assign g[2202] = a[9] & g[1178];
assign g[3225] = b[9] & g[1178];
assign g[2203] = a[9] & g[1179];
assign g[3226] = b[9] & g[1179];
assign g[2204] = a[9] & g[1180];
assign g[3227] = b[9] & g[1180];
assign g[2205] = a[9] & g[1181];
assign g[3228] = b[9] & g[1181];
assign g[2206] = a[9] & g[1182];
assign g[3229] = b[9] & g[1182];
assign g[2207] = a[9] & g[1183];
assign g[3230] = b[9] & g[1183];
assign g[2208] = a[9] & g[1184];
assign g[3231] = b[9] & g[1184];
assign g[2209] = a[9] & g[1185];
assign g[3232] = b[9] & g[1185];
assign g[2210] = a[9] & g[1186];
assign g[3233] = b[9] & g[1186];
assign g[2211] = a[9] & g[1187];
assign g[3234] = b[9] & g[1187];
assign g[2212] = a[9] & g[1188];
assign g[3235] = b[9] & g[1188];
assign g[2213] = a[9] & g[1189];
assign g[3236] = b[9] & g[1189];
assign g[2214] = a[9] & g[1190];
assign g[3237] = b[9] & g[1190];
assign g[2215] = a[9] & g[1191];
assign g[3238] = b[9] & g[1191];
assign g[2216] = a[9] & g[1192];
assign g[3239] = b[9] & g[1192];
assign g[2217] = a[9] & g[1193];
assign g[3240] = b[9] & g[1193];
assign g[2218] = a[9] & g[1194];
assign g[3241] = b[9] & g[1194];
assign g[2219] = a[9] & g[1195];
assign g[3242] = b[9] & g[1195];
assign g[2220] = a[9] & g[1196];
assign g[3243] = b[9] & g[1196];
assign g[2221] = a[9] & g[1197];
assign g[3244] = b[9] & g[1197];
assign g[2222] = a[9] & g[1198];
assign g[3245] = b[9] & g[1198];
assign g[2223] = a[9] & g[1199];
assign g[3246] = b[9] & g[1199];
assign g[2224] = a[9] & g[1200];
assign g[3247] = b[9] & g[1200];
assign g[2225] = a[9] & g[1201];
assign g[3248] = b[9] & g[1201];
assign g[2226] = a[9] & g[1202];
assign g[3249] = b[9] & g[1202];
assign g[2227] = a[9] & g[1203];
assign g[3250] = b[9] & g[1203];
assign g[2228] = a[9] & g[1204];
assign g[3251] = b[9] & g[1204];
assign g[2229] = a[9] & g[1205];
assign g[3252] = b[9] & g[1205];
assign g[2230] = a[9] & g[1206];
assign g[3253] = b[9] & g[1206];
assign g[2231] = a[9] & g[1207];
assign g[3254] = b[9] & g[1207];
assign g[2232] = a[9] & g[1208];
assign g[3255] = b[9] & g[1208];
assign g[2233] = a[9] & g[1209];
assign g[3256] = b[9] & g[1209];
assign g[2234] = a[9] & g[1210];
assign g[3257] = b[9] & g[1210];
assign g[2235] = a[9] & g[1211];
assign g[3258] = b[9] & g[1211];
assign g[2236] = a[9] & g[1212];
assign g[3259] = b[9] & g[1212];
assign g[2237] = a[9] & g[1213];
assign g[3260] = b[9] & g[1213];
assign g[2238] = a[9] & g[1214];
assign g[3261] = b[9] & g[1214];
assign g[2239] = a[9] & g[1215];
assign g[3262] = b[9] & g[1215];
assign g[2240] = a[9] & g[1216];
assign g[3263] = b[9] & g[1216];
assign g[2241] = a[9] & g[1217];
assign g[3264] = b[9] & g[1217];
assign g[2242] = a[9] & g[1218];
assign g[3265] = b[9] & g[1218];
assign g[2243] = a[9] & g[1219];
assign g[3266] = b[9] & g[1219];
assign g[2244] = a[9] & g[1220];
assign g[3267] = b[9] & g[1220];
assign g[2245] = a[9] & g[1221];
assign g[3268] = b[9] & g[1221];
assign g[2246] = a[9] & g[1222];
assign g[3269] = b[9] & g[1222];
assign g[2247] = a[9] & g[1223];
assign g[3270] = b[9] & g[1223];
assign g[2248] = a[9] & g[1224];
assign g[3271] = b[9] & g[1224];
assign g[2249] = a[9] & g[1225];
assign g[3272] = b[9] & g[1225];
assign g[2250] = a[9] & g[1226];
assign g[3273] = b[9] & g[1226];
assign g[2251] = a[9] & g[1227];
assign g[3274] = b[9] & g[1227];
assign g[2252] = a[9] & g[1228];
assign g[3275] = b[9] & g[1228];
assign g[2253] = a[9] & g[1229];
assign g[3276] = b[9] & g[1229];
assign g[2254] = a[9] & g[1230];
assign g[3277] = b[9] & g[1230];
assign g[2255] = a[9] & g[1231];
assign g[3278] = b[9] & g[1231];
assign g[2256] = a[9] & g[1232];
assign g[3279] = b[9] & g[1232];
assign g[2257] = a[9] & g[1233];
assign g[3280] = b[9] & g[1233];
assign g[2258] = a[9] & g[1234];
assign g[3281] = b[9] & g[1234];
assign g[2259] = a[9] & g[1235];
assign g[3282] = b[9] & g[1235];
assign g[2260] = a[9] & g[1236];
assign g[3283] = b[9] & g[1236];
assign g[2261] = a[9] & g[1237];
assign g[3284] = b[9] & g[1237];
assign g[2262] = a[9] & g[1238];
assign g[3285] = b[9] & g[1238];
assign g[2263] = a[9] & g[1239];
assign g[3286] = b[9] & g[1239];
assign g[2264] = a[9] & g[1240];
assign g[3287] = b[9] & g[1240];
assign g[2265] = a[9] & g[1241];
assign g[3288] = b[9] & g[1241];
assign g[2266] = a[9] & g[1242];
assign g[3289] = b[9] & g[1242];
assign g[2267] = a[9] & g[1243];
assign g[3290] = b[9] & g[1243];
assign g[2268] = a[9] & g[1244];
assign g[3291] = b[9] & g[1244];
assign g[2269] = a[9] & g[1245];
assign g[3292] = b[9] & g[1245];
assign g[2270] = a[9] & g[1246];
assign g[3293] = b[9] & g[1246];
assign g[2271] = a[9] & g[1247];
assign g[3294] = b[9] & g[1247];
assign g[2272] = a[9] & g[1248];
assign g[3295] = b[9] & g[1248];
assign g[2273] = a[9] & g[1249];
assign g[3296] = b[9] & g[1249];
assign g[2274] = a[9] & g[1250];
assign g[3297] = b[9] & g[1250];
assign g[2275] = a[9] & g[1251];
assign g[3298] = b[9] & g[1251];
assign g[2276] = a[9] & g[1252];
assign g[3299] = b[9] & g[1252];
assign g[2277] = a[9] & g[1253];
assign g[3300] = b[9] & g[1253];
assign g[2278] = a[9] & g[1254];
assign g[3301] = b[9] & g[1254];
assign g[2279] = a[9] & g[1255];
assign g[3302] = b[9] & g[1255];
assign g[2280] = a[9] & g[1256];
assign g[3303] = b[9] & g[1256];
assign g[2281] = a[9] & g[1257];
assign g[3304] = b[9] & g[1257];
assign g[2282] = a[9] & g[1258];
assign g[3305] = b[9] & g[1258];
assign g[2283] = a[9] & g[1259];
assign g[3306] = b[9] & g[1259];
assign g[2284] = a[9] & g[1260];
assign g[3307] = b[9] & g[1260];
assign g[2285] = a[9] & g[1261];
assign g[3308] = b[9] & g[1261];
assign g[2286] = a[9] & g[1262];
assign g[3309] = b[9] & g[1262];
assign g[2287] = a[9] & g[1263];
assign g[3310] = b[9] & g[1263];
assign g[2288] = a[9] & g[1264];
assign g[3311] = b[9] & g[1264];
assign g[2289] = a[9] & g[1265];
assign g[3312] = b[9] & g[1265];
assign g[2290] = a[9] & g[1266];
assign g[3313] = b[9] & g[1266];
assign g[2291] = a[9] & g[1267];
assign g[3314] = b[9] & g[1267];
assign g[2292] = a[9] & g[1268];
assign g[3315] = b[9] & g[1268];
assign g[2293] = a[9] & g[1269];
assign g[3316] = b[9] & g[1269];
assign g[2294] = a[9] & g[1270];
assign g[3317] = b[9] & g[1270];
assign g[2295] = a[9] & g[1271];
assign g[3318] = b[9] & g[1271];
assign g[2296] = a[9] & g[1272];
assign g[3319] = b[9] & g[1272];
assign g[2297] = a[9] & g[1273];
assign g[3320] = b[9] & g[1273];
assign g[2298] = a[9] & g[1274];
assign g[3321] = b[9] & g[1274];
assign g[2299] = a[9] & g[1275];
assign g[3322] = b[9] & g[1275];
assign g[2300] = a[9] & g[1276];
assign g[3323] = b[9] & g[1276];
assign g[2301] = a[9] & g[1277];
assign g[3324] = b[9] & g[1277];
assign g[2302] = a[9] & g[1278];
assign g[3325] = b[9] & g[1278];
assign g[2303] = a[9] & g[1279];
assign g[3326] = b[9] & g[1279];
assign g[2304] = a[9] & g[1280];
assign g[3327] = b[9] & g[1280];
assign g[2305] = a[9] & g[1281];
assign g[3328] = b[9] & g[1281];
assign g[2306] = a[9] & g[1282];
assign g[3329] = b[9] & g[1282];
assign g[2307] = a[9] & g[1283];
assign g[3330] = b[9] & g[1283];
assign g[2308] = a[9] & g[1284];
assign g[3331] = b[9] & g[1284];
assign g[2309] = a[9] & g[1285];
assign g[3332] = b[9] & g[1285];
assign g[2310] = a[9] & g[1286];
assign g[3333] = b[9] & g[1286];
assign g[2311] = a[9] & g[1287];
assign g[3334] = b[9] & g[1287];
assign g[2312] = a[9] & g[1288];
assign g[3335] = b[9] & g[1288];
assign g[2313] = a[9] & g[1289];
assign g[3336] = b[9] & g[1289];
assign g[2314] = a[9] & g[1290];
assign g[3337] = b[9] & g[1290];
assign g[2315] = a[9] & g[1291];
assign g[3338] = b[9] & g[1291];
assign g[2316] = a[9] & g[1292];
assign g[3339] = b[9] & g[1292];
assign g[2317] = a[9] & g[1293];
assign g[3340] = b[9] & g[1293];
assign g[2318] = a[9] & g[1294];
assign g[3341] = b[9] & g[1294];
assign g[2319] = a[9] & g[1295];
assign g[3342] = b[9] & g[1295];
assign g[2320] = a[9] & g[1296];
assign g[3343] = b[9] & g[1296];
assign g[2321] = a[9] & g[1297];
assign g[3344] = b[9] & g[1297];
assign g[2322] = a[9] & g[1298];
assign g[3345] = b[9] & g[1298];
assign g[2323] = a[9] & g[1299];
assign g[3346] = b[9] & g[1299];
assign g[2324] = a[9] & g[1300];
assign g[3347] = b[9] & g[1300];
assign g[2325] = a[9] & g[1301];
assign g[3348] = b[9] & g[1301];
assign g[2326] = a[9] & g[1302];
assign g[3349] = b[9] & g[1302];
assign g[2327] = a[9] & g[1303];
assign g[3350] = b[9] & g[1303];
assign g[2328] = a[9] & g[1304];
assign g[3351] = b[9] & g[1304];
assign g[2329] = a[9] & g[1305];
assign g[3352] = b[9] & g[1305];
assign g[2330] = a[9] & g[1306];
assign g[3353] = b[9] & g[1306];
assign g[2331] = a[9] & g[1307];
assign g[3354] = b[9] & g[1307];
assign g[2332] = a[9] & g[1308];
assign g[3355] = b[9] & g[1308];
assign g[2333] = a[9] & g[1309];
assign g[3356] = b[9] & g[1309];
assign g[2334] = a[9] & g[1310];
assign g[3357] = b[9] & g[1310];
assign g[2335] = a[9] & g[1311];
assign g[3358] = b[9] & g[1311];
assign g[2336] = a[9] & g[1312];
assign g[3359] = b[9] & g[1312];
assign g[2337] = a[9] & g[1313];
assign g[3360] = b[9] & g[1313];
assign g[2338] = a[9] & g[1314];
assign g[3361] = b[9] & g[1314];
assign g[2339] = a[9] & g[1315];
assign g[3362] = b[9] & g[1315];
assign g[2340] = a[9] & g[1316];
assign g[3363] = b[9] & g[1316];
assign g[2341] = a[9] & g[1317];
assign g[3364] = b[9] & g[1317];
assign g[2342] = a[9] & g[1318];
assign g[3365] = b[9] & g[1318];
assign g[2343] = a[9] & g[1319];
assign g[3366] = b[9] & g[1319];
assign g[2344] = a[9] & g[1320];
assign g[3367] = b[9] & g[1320];
assign g[2345] = a[9] & g[1321];
assign g[3368] = b[9] & g[1321];
assign g[2346] = a[9] & g[1322];
assign g[3369] = b[9] & g[1322];
assign g[2347] = a[9] & g[1323];
assign g[3370] = b[9] & g[1323];
assign g[2348] = a[9] & g[1324];
assign g[3371] = b[9] & g[1324];
assign g[2349] = a[9] & g[1325];
assign g[3372] = b[9] & g[1325];
assign g[2350] = a[9] & g[1326];
assign g[3373] = b[9] & g[1326];
assign g[2351] = a[9] & g[1327];
assign g[3374] = b[9] & g[1327];
assign g[2352] = a[9] & g[1328];
assign g[3375] = b[9] & g[1328];
assign g[2353] = a[9] & g[1329];
assign g[3376] = b[9] & g[1329];
assign g[2354] = a[9] & g[1330];
assign g[3377] = b[9] & g[1330];
assign g[2355] = a[9] & g[1331];
assign g[3378] = b[9] & g[1331];
assign g[2356] = a[9] & g[1332];
assign g[3379] = b[9] & g[1332];
assign g[2357] = a[9] & g[1333];
assign g[3380] = b[9] & g[1333];
assign g[2358] = a[9] & g[1334];
assign g[3381] = b[9] & g[1334];
assign g[2359] = a[9] & g[1335];
assign g[3382] = b[9] & g[1335];
assign g[2360] = a[9] & g[1336];
assign g[3383] = b[9] & g[1336];
assign g[2361] = a[9] & g[1337];
assign g[3384] = b[9] & g[1337];
assign g[2362] = a[9] & g[1338];
assign g[3385] = b[9] & g[1338];
assign g[2363] = a[9] & g[1339];
assign g[3386] = b[9] & g[1339];
assign g[2364] = a[9] & g[1340];
assign g[3387] = b[9] & g[1340];
assign g[2365] = a[9] & g[1341];
assign g[3388] = b[9] & g[1341];
assign g[2366] = a[9] & g[1342];
assign g[3389] = b[9] & g[1342];
assign g[2367] = a[9] & g[1343];
assign g[3390] = b[9] & g[1343];
assign g[2368] = a[9] & g[1344];
assign g[3391] = b[9] & g[1344];
assign g[2369] = a[9] & g[1345];
assign g[3392] = b[9] & g[1345];
assign g[2370] = a[9] & g[1346];
assign g[3393] = b[9] & g[1346];
assign g[2371] = a[9] & g[1347];
assign g[3394] = b[9] & g[1347];
assign g[2372] = a[9] & g[1348];
assign g[3395] = b[9] & g[1348];
assign g[2373] = a[9] & g[1349];
assign g[3396] = b[9] & g[1349];
assign g[2374] = a[9] & g[1350];
assign g[3397] = b[9] & g[1350];
assign g[2375] = a[9] & g[1351];
assign g[3398] = b[9] & g[1351];
assign g[2376] = a[9] & g[1352];
assign g[3399] = b[9] & g[1352];
assign g[2377] = a[9] & g[1353];
assign g[3400] = b[9] & g[1353];
assign g[2378] = a[9] & g[1354];
assign g[3401] = b[9] & g[1354];
assign g[2379] = a[9] & g[1355];
assign g[3402] = b[9] & g[1355];
assign g[2380] = a[9] & g[1356];
assign g[3403] = b[9] & g[1356];
assign g[2381] = a[9] & g[1357];
assign g[3404] = b[9] & g[1357];
assign g[2382] = a[9] & g[1358];
assign g[3405] = b[9] & g[1358];
assign g[2383] = a[9] & g[1359];
assign g[3406] = b[9] & g[1359];
assign g[2384] = a[9] & g[1360];
assign g[3407] = b[9] & g[1360];
assign g[2385] = a[9] & g[1361];
assign g[3408] = b[9] & g[1361];
assign g[2386] = a[9] & g[1362];
assign g[3409] = b[9] & g[1362];
assign g[2387] = a[9] & g[1363];
assign g[3410] = b[9] & g[1363];
assign g[2388] = a[9] & g[1364];
assign g[3411] = b[9] & g[1364];
assign g[2389] = a[9] & g[1365];
assign g[3412] = b[9] & g[1365];
assign g[2390] = a[9] & g[1366];
assign g[3413] = b[9] & g[1366];
assign g[2391] = a[9] & g[1367];
assign g[3414] = b[9] & g[1367];
assign g[2392] = a[9] & g[1368];
assign g[3415] = b[9] & g[1368];
assign g[2393] = a[9] & g[1369];
assign g[3416] = b[9] & g[1369];
assign g[2394] = a[9] & g[1370];
assign g[3417] = b[9] & g[1370];
assign g[2395] = a[9] & g[1371];
assign g[3418] = b[9] & g[1371];
assign g[2396] = a[9] & g[1372];
assign g[3419] = b[9] & g[1372];
assign g[2397] = a[9] & g[1373];
assign g[3420] = b[9] & g[1373];
assign g[2398] = a[9] & g[1374];
assign g[3421] = b[9] & g[1374];
assign g[2399] = a[9] & g[1375];
assign g[3422] = b[9] & g[1375];
assign g[2400] = a[9] & g[1376];
assign g[3423] = b[9] & g[1376];
assign g[2401] = a[9] & g[1377];
assign g[3424] = b[9] & g[1377];
assign g[2402] = a[9] & g[1378];
assign g[3425] = b[9] & g[1378];
assign g[2403] = a[9] & g[1379];
assign g[3426] = b[9] & g[1379];
assign g[2404] = a[9] & g[1380];
assign g[3427] = b[9] & g[1380];
assign g[2405] = a[9] & g[1381];
assign g[3428] = b[9] & g[1381];
assign g[2406] = a[9] & g[1382];
assign g[3429] = b[9] & g[1382];
assign g[2407] = a[9] & g[1383];
assign g[3430] = b[9] & g[1383];
assign g[2408] = a[9] & g[1384];
assign g[3431] = b[9] & g[1384];
assign g[2409] = a[9] & g[1385];
assign g[3432] = b[9] & g[1385];
assign g[2410] = a[9] & g[1386];
assign g[3433] = b[9] & g[1386];
assign g[2411] = a[9] & g[1387];
assign g[3434] = b[9] & g[1387];
assign g[2412] = a[9] & g[1388];
assign g[3435] = b[9] & g[1388];
assign g[2413] = a[9] & g[1389];
assign g[3436] = b[9] & g[1389];
assign g[2414] = a[9] & g[1390];
assign g[3437] = b[9] & g[1390];
assign g[2415] = a[9] & g[1391];
assign g[3438] = b[9] & g[1391];
assign g[2416] = a[9] & g[1392];
assign g[3439] = b[9] & g[1392];
assign g[2417] = a[9] & g[1393];
assign g[3440] = b[9] & g[1393];
assign g[2418] = a[9] & g[1394];
assign g[3441] = b[9] & g[1394];
assign g[2419] = a[9] & g[1395];
assign g[3442] = b[9] & g[1395];
assign g[2420] = a[9] & g[1396];
assign g[3443] = b[9] & g[1396];
assign g[2421] = a[9] & g[1397];
assign g[3444] = b[9] & g[1397];
assign g[2422] = a[9] & g[1398];
assign g[3445] = b[9] & g[1398];
assign g[2423] = a[9] & g[1399];
assign g[3446] = b[9] & g[1399];
assign g[2424] = a[9] & g[1400];
assign g[3447] = b[9] & g[1400];
assign g[2425] = a[9] & g[1401];
assign g[3448] = b[9] & g[1401];
assign g[2426] = a[9] & g[1402];
assign g[3449] = b[9] & g[1402];
assign g[2427] = a[9] & g[1403];
assign g[3450] = b[9] & g[1403];
assign g[2428] = a[9] & g[1404];
assign g[3451] = b[9] & g[1404];
assign g[2429] = a[9] & g[1405];
assign g[3452] = b[9] & g[1405];
assign g[2430] = a[9] & g[1406];
assign g[3453] = b[9] & g[1406];
assign g[2431] = a[9] & g[1407];
assign g[3454] = b[9] & g[1407];
assign g[2432] = a[9] & g[1408];
assign g[3455] = b[9] & g[1408];
assign g[2433] = a[9] & g[1409];
assign g[3456] = b[9] & g[1409];
assign g[2434] = a[9] & g[1410];
assign g[3457] = b[9] & g[1410];
assign g[2435] = a[9] & g[1411];
assign g[3458] = b[9] & g[1411];
assign g[2436] = a[9] & g[1412];
assign g[3459] = b[9] & g[1412];
assign g[2437] = a[9] & g[1413];
assign g[3460] = b[9] & g[1413];
assign g[2438] = a[9] & g[1414];
assign g[3461] = b[9] & g[1414];
assign g[2439] = a[9] & g[1415];
assign g[3462] = b[9] & g[1415];
assign g[2440] = a[9] & g[1416];
assign g[3463] = b[9] & g[1416];
assign g[2441] = a[9] & g[1417];
assign g[3464] = b[9] & g[1417];
assign g[2442] = a[9] & g[1418];
assign g[3465] = b[9] & g[1418];
assign g[2443] = a[9] & g[1419];
assign g[3466] = b[9] & g[1419];
assign g[2444] = a[9] & g[1420];
assign g[3467] = b[9] & g[1420];
assign g[2445] = a[9] & g[1421];
assign g[3468] = b[9] & g[1421];
assign g[2446] = a[9] & g[1422];
assign g[3469] = b[9] & g[1422];
assign g[2447] = a[9] & g[1423];
assign g[3470] = b[9] & g[1423];
assign g[2448] = a[9] & g[1424];
assign g[3471] = b[9] & g[1424];
assign g[2449] = a[9] & g[1425];
assign g[3472] = b[9] & g[1425];
assign g[2450] = a[9] & g[1426];
assign g[3473] = b[9] & g[1426];
assign g[2451] = a[9] & g[1427];
assign g[3474] = b[9] & g[1427];
assign g[2452] = a[9] & g[1428];
assign g[3475] = b[9] & g[1428];
assign g[2453] = a[9] & g[1429];
assign g[3476] = b[9] & g[1429];
assign g[2454] = a[9] & g[1430];
assign g[3477] = b[9] & g[1430];
assign g[2455] = a[9] & g[1431];
assign g[3478] = b[9] & g[1431];
assign g[2456] = a[9] & g[1432];
assign g[3479] = b[9] & g[1432];
assign g[2457] = a[9] & g[1433];
assign g[3480] = b[9] & g[1433];
assign g[2458] = a[9] & g[1434];
assign g[3481] = b[9] & g[1434];
assign g[2459] = a[9] & g[1435];
assign g[3482] = b[9] & g[1435];
assign g[2460] = a[9] & g[1436];
assign g[3483] = b[9] & g[1436];
assign g[2461] = a[9] & g[1437];
assign g[3484] = b[9] & g[1437];
assign g[2462] = a[9] & g[1438];
assign g[3485] = b[9] & g[1438];
assign g[2463] = a[9] & g[1439];
assign g[3486] = b[9] & g[1439];
assign g[2464] = a[9] & g[1440];
assign g[3487] = b[9] & g[1440];
assign g[2465] = a[9] & g[1441];
assign g[3488] = b[9] & g[1441];
assign g[2466] = a[9] & g[1442];
assign g[3489] = b[9] & g[1442];
assign g[2467] = a[9] & g[1443];
assign g[3490] = b[9] & g[1443];
assign g[2468] = a[9] & g[1444];
assign g[3491] = b[9] & g[1444];
assign g[2469] = a[9] & g[1445];
assign g[3492] = b[9] & g[1445];
assign g[2470] = a[9] & g[1446];
assign g[3493] = b[9] & g[1446];
assign g[2471] = a[9] & g[1447];
assign g[3494] = b[9] & g[1447];
assign g[2472] = a[9] & g[1448];
assign g[3495] = b[9] & g[1448];
assign g[2473] = a[9] & g[1449];
assign g[3496] = b[9] & g[1449];
assign g[2474] = a[9] & g[1450];
assign g[3497] = b[9] & g[1450];
assign g[2475] = a[9] & g[1451];
assign g[3498] = b[9] & g[1451];
assign g[2476] = a[9] & g[1452];
assign g[3499] = b[9] & g[1452];
assign g[2477] = a[9] & g[1453];
assign g[3500] = b[9] & g[1453];
assign g[2478] = a[9] & g[1454];
assign g[3501] = b[9] & g[1454];
assign g[2479] = a[9] & g[1455];
assign g[3502] = b[9] & g[1455];
assign g[2480] = a[9] & g[1456];
assign g[3503] = b[9] & g[1456];
assign g[2481] = a[9] & g[1457];
assign g[3504] = b[9] & g[1457];
assign g[2482] = a[9] & g[1458];
assign g[3505] = b[9] & g[1458];
assign g[2483] = a[9] & g[1459];
assign g[3506] = b[9] & g[1459];
assign g[2484] = a[9] & g[1460];
assign g[3507] = b[9] & g[1460];
assign g[2485] = a[9] & g[1461];
assign g[3508] = b[9] & g[1461];
assign g[2486] = a[9] & g[1462];
assign g[3509] = b[9] & g[1462];
assign g[2487] = a[9] & g[1463];
assign g[3510] = b[9] & g[1463];
assign g[2488] = a[9] & g[1464];
assign g[3511] = b[9] & g[1464];
assign g[2489] = a[9] & g[1465];
assign g[3512] = b[9] & g[1465];
assign g[2490] = a[9] & g[1466];
assign g[3513] = b[9] & g[1466];
assign g[2491] = a[9] & g[1467];
assign g[3514] = b[9] & g[1467];
assign g[2492] = a[9] & g[1468];
assign g[3515] = b[9] & g[1468];
assign g[2493] = a[9] & g[1469];
assign g[3516] = b[9] & g[1469];
assign g[2494] = a[9] & g[1470];
assign g[3517] = b[9] & g[1470];
assign g[2495] = a[9] & g[1471];
assign g[3518] = b[9] & g[1471];
assign g[2496] = a[9] & g[1472];
assign g[3519] = b[9] & g[1472];
assign g[2497] = a[9] & g[1473];
assign g[3520] = b[9] & g[1473];
assign g[2498] = a[9] & g[1474];
assign g[3521] = b[9] & g[1474];
assign g[2499] = a[9] & g[1475];
assign g[3522] = b[9] & g[1475];
assign g[2500] = a[9] & g[1476];
assign g[3523] = b[9] & g[1476];
assign g[2501] = a[9] & g[1477];
assign g[3524] = b[9] & g[1477];
assign g[2502] = a[9] & g[1478];
assign g[3525] = b[9] & g[1478];
assign g[2503] = a[9] & g[1479];
assign g[3526] = b[9] & g[1479];
assign g[2504] = a[9] & g[1480];
assign g[3527] = b[9] & g[1480];
assign g[2505] = a[9] & g[1481];
assign g[3528] = b[9] & g[1481];
assign g[2506] = a[9] & g[1482];
assign g[3529] = b[9] & g[1482];
assign g[2507] = a[9] & g[1483];
assign g[3530] = b[9] & g[1483];
assign g[2508] = a[9] & g[1484];
assign g[3531] = b[9] & g[1484];
assign g[2509] = a[9] & g[1485];
assign g[3532] = b[9] & g[1485];
assign g[2510] = a[9] & g[1486];
assign g[3533] = b[9] & g[1486];
assign g[2511] = a[9] & g[1487];
assign g[3534] = b[9] & g[1487];
assign g[2512] = a[9] & g[1488];
assign g[3535] = b[9] & g[1488];
assign g[2513] = a[9] & g[1489];
assign g[3536] = b[9] & g[1489];
assign g[2514] = a[9] & g[1490];
assign g[3537] = b[9] & g[1490];
assign g[2515] = a[9] & g[1491];
assign g[3538] = b[9] & g[1491];
assign g[2516] = a[9] & g[1492];
assign g[3539] = b[9] & g[1492];
assign g[2517] = a[9] & g[1493];
assign g[3540] = b[9] & g[1493];
assign g[2518] = a[9] & g[1494];
assign g[3541] = b[9] & g[1494];
assign g[2519] = a[9] & g[1495];
assign g[3542] = b[9] & g[1495];
assign g[2520] = a[9] & g[1496];
assign g[3543] = b[9] & g[1496];
assign g[2521] = a[9] & g[1497];
assign g[3544] = b[9] & g[1497];
assign g[2522] = a[9] & g[1498];
assign g[3545] = b[9] & g[1498];
assign g[2523] = a[9] & g[1499];
assign g[3546] = b[9] & g[1499];
assign g[2524] = a[9] & g[1500];
assign g[3547] = b[9] & g[1500];
assign g[2525] = a[9] & g[1501];
assign g[3548] = b[9] & g[1501];
assign g[2526] = a[9] & g[1502];
assign g[3549] = b[9] & g[1502];
assign g[2527] = a[9] & g[1503];
assign g[3550] = b[9] & g[1503];
assign g[2528] = a[9] & g[1504];
assign g[3551] = b[9] & g[1504];
assign g[2529] = a[9] & g[1505];
assign g[3552] = b[9] & g[1505];
assign g[2530] = a[9] & g[1506];
assign g[3553] = b[9] & g[1506];
assign g[2531] = a[9] & g[1507];
assign g[3554] = b[9] & g[1507];
assign g[2532] = a[9] & g[1508];
assign g[3555] = b[9] & g[1508];
assign g[2533] = a[9] & g[1509];
assign g[3556] = b[9] & g[1509];
assign g[2534] = a[9] & g[1510];
assign g[3557] = b[9] & g[1510];
assign g[2535] = a[9] & g[1511];
assign g[3558] = b[9] & g[1511];
assign g[2536] = a[9] & g[1512];
assign g[3559] = b[9] & g[1512];
assign g[2537] = a[9] & g[1513];
assign g[3560] = b[9] & g[1513];
assign g[2538] = a[9] & g[1514];
assign g[3561] = b[9] & g[1514];
assign g[2539] = a[9] & g[1515];
assign g[3562] = b[9] & g[1515];
assign g[2540] = a[9] & g[1516];
assign g[3563] = b[9] & g[1516];
assign g[2541] = a[9] & g[1517];
assign g[3564] = b[9] & g[1517];
assign g[2542] = a[9] & g[1518];
assign g[3565] = b[9] & g[1518];
assign g[2543] = a[9] & g[1519];
assign g[3566] = b[9] & g[1519];
assign g[2544] = a[9] & g[1520];
assign g[3567] = b[9] & g[1520];
assign g[2545] = a[9] & g[1521];
assign g[3568] = b[9] & g[1521];
assign g[2546] = a[9] & g[1522];
assign g[3569] = b[9] & g[1522];
assign g[2547] = a[9] & g[1523];
assign g[3570] = b[9] & g[1523];
assign g[2548] = a[9] & g[1524];
assign g[3571] = b[9] & g[1524];
assign g[2549] = a[9] & g[1525];
assign g[3572] = b[9] & g[1525];
assign g[2550] = a[9] & g[1526];
assign g[3573] = b[9] & g[1526];
assign g[2551] = a[9] & g[1527];
assign g[3574] = b[9] & g[1527];
assign g[2552] = a[9] & g[1528];
assign g[3575] = b[9] & g[1528];
assign g[2553] = a[9] & g[1529];
assign g[3576] = b[9] & g[1529];
assign g[2554] = a[9] & g[1530];
assign g[3577] = b[9] & g[1530];
assign g[2555] = a[9] & g[1531];
assign g[3578] = b[9] & g[1531];
assign g[2556] = a[9] & g[1532];
assign g[3579] = b[9] & g[1532];
assign g[2557] = a[9] & g[1533];
assign g[3580] = b[9] & g[1533];
assign g[2558] = a[9] & g[1534];
assign g[3581] = b[9] & g[1534];
assign g[2559] = a[9] & g[1535];
assign g[3582] = b[9] & g[1535];
assign g[2560] = a[9] & g[1536];
assign g[3583] = b[9] & g[1536];
assign g[2561] = a[9] & g[1537];
assign g[3584] = b[9] & g[1537];
assign g[2562] = a[9] & g[1538];
assign g[3585] = b[9] & g[1538];
assign g[2563] = a[9] & g[1539];
assign g[3586] = b[9] & g[1539];
assign g[2564] = a[9] & g[1540];
assign g[3587] = b[9] & g[1540];
assign g[2565] = a[9] & g[1541];
assign g[3588] = b[9] & g[1541];
assign g[2566] = a[9] & g[1542];
assign g[3589] = b[9] & g[1542];
assign g[2567] = a[9] & g[1543];
assign g[3590] = b[9] & g[1543];
assign g[2568] = a[9] & g[1544];
assign g[3591] = b[9] & g[1544];
assign g[2569] = a[9] & g[1545];
assign g[3592] = b[9] & g[1545];
assign g[2570] = a[9] & g[1546];
assign g[3593] = b[9] & g[1546];
assign g[2571] = a[9] & g[1547];
assign g[3594] = b[9] & g[1547];
assign g[2572] = a[9] & g[1548];
assign g[3595] = b[9] & g[1548];
assign g[2573] = a[9] & g[1549];
assign g[3596] = b[9] & g[1549];
assign g[2574] = a[9] & g[1550];
assign g[3597] = b[9] & g[1550];
assign g[2575] = a[9] & g[1551];
assign g[3598] = b[9] & g[1551];
assign g[2576] = a[9] & g[1552];
assign g[3599] = b[9] & g[1552];
assign g[2577] = a[9] & g[1553];
assign g[3600] = b[9] & g[1553];
assign g[2578] = a[9] & g[1554];
assign g[3601] = b[9] & g[1554];
assign g[2579] = a[9] & g[1555];
assign g[3602] = b[9] & g[1555];
assign g[2580] = a[9] & g[1556];
assign g[3603] = b[9] & g[1556];
assign g[2581] = a[9] & g[1557];
assign g[3604] = b[9] & g[1557];
assign g[2582] = a[9] & g[1558];
assign g[3605] = b[9] & g[1558];
assign g[2583] = a[9] & g[1559];
assign g[3606] = b[9] & g[1559];
assign g[2584] = a[9] & g[1560];
assign g[3607] = b[9] & g[1560];
assign g[2585] = a[9] & g[1561];
assign g[3608] = b[9] & g[1561];
assign g[2586] = a[9] & g[1562];
assign g[3609] = b[9] & g[1562];
assign g[2587] = a[9] & g[1563];
assign g[3610] = b[9] & g[1563];
assign g[2588] = a[9] & g[1564];
assign g[3611] = b[9] & g[1564];
assign g[2589] = a[9] & g[1565];
assign g[3612] = b[9] & g[1565];
assign g[2590] = a[9] & g[1566];
assign g[3613] = b[9] & g[1566];
assign g[2591] = a[9] & g[1567];
assign g[3614] = b[9] & g[1567];
assign g[2592] = a[9] & g[1568];
assign g[3615] = b[9] & g[1568];
assign g[2593] = a[9] & g[1569];
assign g[3616] = b[9] & g[1569];
assign g[2594] = a[9] & g[1570];
assign g[3617] = b[9] & g[1570];
assign g[2595] = a[9] & g[1571];
assign g[3618] = b[9] & g[1571];
assign g[2596] = a[9] & g[1572];
assign g[3619] = b[9] & g[1572];
assign g[2597] = a[9] & g[1573];
assign g[3620] = b[9] & g[1573];
assign g[2598] = a[9] & g[1574];
assign g[3621] = b[9] & g[1574];
assign g[2599] = a[9] & g[1575];
assign g[3622] = b[9] & g[1575];
assign g[2600] = a[9] & g[1576];
assign g[3623] = b[9] & g[1576];
assign g[2601] = a[9] & g[1577];
assign g[3624] = b[9] & g[1577];
assign g[2602] = a[9] & g[1578];
assign g[3625] = b[9] & g[1578];
assign g[2603] = a[9] & g[1579];
assign g[3626] = b[9] & g[1579];
assign g[2604] = a[9] & g[1580];
assign g[3627] = b[9] & g[1580];
assign g[2605] = a[9] & g[1581];
assign g[3628] = b[9] & g[1581];
assign g[2606] = a[9] & g[1582];
assign g[3629] = b[9] & g[1582];
assign g[2607] = a[9] & g[1583];
assign g[3630] = b[9] & g[1583];
assign g[2608] = a[9] & g[1584];
assign g[3631] = b[9] & g[1584];
assign g[2609] = a[9] & g[1585];
assign g[3632] = b[9] & g[1585];
assign g[2610] = a[9] & g[1586];
assign g[3633] = b[9] & g[1586];
assign g[2611] = a[9] & g[1587];
assign g[3634] = b[9] & g[1587];
assign g[2612] = a[9] & g[1588];
assign g[3635] = b[9] & g[1588];
assign g[2613] = a[9] & g[1589];
assign g[3636] = b[9] & g[1589];
assign g[2614] = a[9] & g[1590];
assign g[3637] = b[9] & g[1590];
assign g[2615] = a[9] & g[1591];
assign g[3638] = b[9] & g[1591];
assign g[2616] = a[9] & g[1592];
assign g[3639] = b[9] & g[1592];
assign g[2617] = a[9] & g[1593];
assign g[3640] = b[9] & g[1593];
assign g[2618] = a[9] & g[1594];
assign g[3641] = b[9] & g[1594];
assign g[2619] = a[9] & g[1595];
assign g[3642] = b[9] & g[1595];
assign g[2620] = a[9] & g[1596];
assign g[3643] = b[9] & g[1596];
assign g[2621] = a[9] & g[1597];
assign g[3644] = b[9] & g[1597];
assign g[2622] = a[9] & g[1598];
assign g[3645] = b[9] & g[1598];
assign g[2623] = a[9] & g[1599];
assign g[3646] = b[9] & g[1599];
assign g[2624] = a[9] & g[1600];
assign g[3647] = b[9] & g[1600];
assign g[2625] = a[9] & g[1601];
assign g[3648] = b[9] & g[1601];
assign g[2626] = a[9] & g[1602];
assign g[3649] = b[9] & g[1602];
assign g[2627] = a[9] & g[1603];
assign g[3650] = b[9] & g[1603];
assign g[2628] = a[9] & g[1604];
assign g[3651] = b[9] & g[1604];
assign g[2629] = a[9] & g[1605];
assign g[3652] = b[9] & g[1605];
assign g[2630] = a[9] & g[1606];
assign g[3653] = b[9] & g[1606];
assign g[2631] = a[9] & g[1607];
assign g[3654] = b[9] & g[1607];
assign g[2632] = a[9] & g[1608];
assign g[3655] = b[9] & g[1608];
assign g[2633] = a[9] & g[1609];
assign g[3656] = b[9] & g[1609];
assign g[2634] = a[9] & g[1610];
assign g[3657] = b[9] & g[1610];
assign g[2635] = a[9] & g[1611];
assign g[3658] = b[9] & g[1611];
assign g[2636] = a[9] & g[1612];
assign g[3659] = b[9] & g[1612];
assign g[2637] = a[9] & g[1613];
assign g[3660] = b[9] & g[1613];
assign g[2638] = a[9] & g[1614];
assign g[3661] = b[9] & g[1614];
assign g[2639] = a[9] & g[1615];
assign g[3662] = b[9] & g[1615];
assign g[2640] = a[9] & g[1616];
assign g[3663] = b[9] & g[1616];
assign g[2641] = a[9] & g[1617];
assign g[3664] = b[9] & g[1617];
assign g[2642] = a[9] & g[1618];
assign g[3665] = b[9] & g[1618];
assign g[2643] = a[9] & g[1619];
assign g[3666] = b[9] & g[1619];
assign g[2644] = a[9] & g[1620];
assign g[3667] = b[9] & g[1620];
assign g[2645] = a[9] & g[1621];
assign g[3668] = b[9] & g[1621];
assign g[2646] = a[9] & g[1622];
assign g[3669] = b[9] & g[1622];
assign g[2647] = a[9] & g[1623];
assign g[3670] = b[9] & g[1623];
assign g[2648] = a[9] & g[1624];
assign g[3671] = b[9] & g[1624];
assign g[2649] = a[9] & g[1625];
assign g[3672] = b[9] & g[1625];
assign g[2650] = a[9] & g[1626];
assign g[3673] = b[9] & g[1626];
assign g[2651] = a[9] & g[1627];
assign g[3674] = b[9] & g[1627];
assign g[2652] = a[9] & g[1628];
assign g[3675] = b[9] & g[1628];
assign g[2653] = a[9] & g[1629];
assign g[3676] = b[9] & g[1629];
assign g[2654] = a[9] & g[1630];
assign g[3677] = b[9] & g[1630];
assign g[2655] = a[9] & g[1631];
assign g[3678] = b[9] & g[1631];
assign g[2656] = a[9] & g[1632];
assign g[3679] = b[9] & g[1632];
assign g[2657] = a[9] & g[1633];
assign g[3680] = b[9] & g[1633];
assign g[2658] = a[9] & g[1634];
assign g[3681] = b[9] & g[1634];
assign g[2659] = a[9] & g[1635];
assign g[3682] = b[9] & g[1635];
assign g[2660] = a[9] & g[1636];
assign g[3683] = b[9] & g[1636];
assign g[2661] = a[9] & g[1637];
assign g[3684] = b[9] & g[1637];
assign g[2662] = a[9] & g[1638];
assign g[3685] = b[9] & g[1638];
assign g[2663] = a[9] & g[1639];
assign g[3686] = b[9] & g[1639];
assign g[2664] = a[9] & g[1640];
assign g[3687] = b[9] & g[1640];
assign g[2665] = a[9] & g[1641];
assign g[3688] = b[9] & g[1641];
assign g[2666] = a[9] & g[1642];
assign g[3689] = b[9] & g[1642];
assign g[2667] = a[9] & g[1643];
assign g[3690] = b[9] & g[1643];
assign g[2668] = a[9] & g[1644];
assign g[3691] = b[9] & g[1644];
assign g[2669] = a[9] & g[1645];
assign g[3692] = b[9] & g[1645];
assign g[2670] = a[9] & g[1646];
assign g[3693] = b[9] & g[1646];
assign g[2671] = a[9] & g[1647];
assign g[3694] = b[9] & g[1647];
assign g[2672] = a[9] & g[1648];
assign g[3695] = b[9] & g[1648];
assign g[2673] = a[9] & g[1649];
assign g[3696] = b[9] & g[1649];
assign g[2674] = a[9] & g[1650];
assign g[3697] = b[9] & g[1650];
assign g[2675] = a[9] & g[1651];
assign g[3698] = b[9] & g[1651];
assign g[2676] = a[9] & g[1652];
assign g[3699] = b[9] & g[1652];
assign g[2677] = a[9] & g[1653];
assign g[3700] = b[9] & g[1653];
assign g[2678] = a[9] & g[1654];
assign g[3701] = b[9] & g[1654];
assign g[2679] = a[9] & g[1655];
assign g[3702] = b[9] & g[1655];
assign g[2680] = a[9] & g[1656];
assign g[3703] = b[9] & g[1656];
assign g[2681] = a[9] & g[1657];
assign g[3704] = b[9] & g[1657];
assign g[2682] = a[9] & g[1658];
assign g[3705] = b[9] & g[1658];
assign g[2683] = a[9] & g[1659];
assign g[3706] = b[9] & g[1659];
assign g[2684] = a[9] & g[1660];
assign g[3707] = b[9] & g[1660];
assign g[2685] = a[9] & g[1661];
assign g[3708] = b[9] & g[1661];
assign g[2686] = a[9] & g[1662];
assign g[3709] = b[9] & g[1662];
assign g[2687] = a[9] & g[1663];
assign g[3710] = b[9] & g[1663];
assign g[2688] = a[9] & g[1664];
assign g[3711] = b[9] & g[1664];
assign g[2689] = a[9] & g[1665];
assign g[3712] = b[9] & g[1665];
assign g[2690] = a[9] & g[1666];
assign g[3713] = b[9] & g[1666];
assign g[2691] = a[9] & g[1667];
assign g[3714] = b[9] & g[1667];
assign g[2692] = a[9] & g[1668];
assign g[3715] = b[9] & g[1668];
assign g[2693] = a[9] & g[1669];
assign g[3716] = b[9] & g[1669];
assign g[2694] = a[9] & g[1670];
assign g[3717] = b[9] & g[1670];
assign g[2695] = a[9] & g[1671];
assign g[3718] = b[9] & g[1671];
assign g[2696] = a[9] & g[1672];
assign g[3719] = b[9] & g[1672];
assign g[2697] = a[9] & g[1673];
assign g[3720] = b[9] & g[1673];
assign g[2698] = a[9] & g[1674];
assign g[3721] = b[9] & g[1674];
assign g[2699] = a[9] & g[1675];
assign g[3722] = b[9] & g[1675];
assign g[2700] = a[9] & g[1676];
assign g[3723] = b[9] & g[1676];
assign g[2701] = a[9] & g[1677];
assign g[3724] = b[9] & g[1677];
assign g[2702] = a[9] & g[1678];
assign g[3725] = b[9] & g[1678];
assign g[2703] = a[9] & g[1679];
assign g[3726] = b[9] & g[1679];
assign g[2704] = a[9] & g[1680];
assign g[3727] = b[9] & g[1680];
assign g[2705] = a[9] & g[1681];
assign g[3728] = b[9] & g[1681];
assign g[2706] = a[9] & g[1682];
assign g[3729] = b[9] & g[1682];
assign g[2707] = a[9] & g[1683];
assign g[3730] = b[9] & g[1683];
assign g[2708] = a[9] & g[1684];
assign g[3731] = b[9] & g[1684];
assign g[2709] = a[9] & g[1685];
assign g[3732] = b[9] & g[1685];
assign g[2710] = a[9] & g[1686];
assign g[3733] = b[9] & g[1686];
assign g[2711] = a[9] & g[1687];
assign g[3734] = b[9] & g[1687];
assign g[2712] = a[9] & g[1688];
assign g[3735] = b[9] & g[1688];
assign g[2713] = a[9] & g[1689];
assign g[3736] = b[9] & g[1689];
assign g[2714] = a[9] & g[1690];
assign g[3737] = b[9] & g[1690];
assign g[2715] = a[9] & g[1691];
assign g[3738] = b[9] & g[1691];
assign g[2716] = a[9] & g[1692];
assign g[3739] = b[9] & g[1692];
assign g[2717] = a[9] & g[1693];
assign g[3740] = b[9] & g[1693];
assign g[2718] = a[9] & g[1694];
assign g[3741] = b[9] & g[1694];
assign g[2719] = a[9] & g[1695];
assign g[3742] = b[9] & g[1695];
assign g[2720] = a[9] & g[1696];
assign g[3743] = b[9] & g[1696];
assign g[2721] = a[9] & g[1697];
assign g[3744] = b[9] & g[1697];
assign g[2722] = a[9] & g[1698];
assign g[3745] = b[9] & g[1698];
assign g[2723] = a[9] & g[1699];
assign g[3746] = b[9] & g[1699];
assign g[2724] = a[9] & g[1700];
assign g[3747] = b[9] & g[1700];
assign g[2725] = a[9] & g[1701];
assign g[3748] = b[9] & g[1701];
assign g[2726] = a[9] & g[1702];
assign g[3749] = b[9] & g[1702];
assign g[2727] = a[9] & g[1703];
assign g[3750] = b[9] & g[1703];
assign g[2728] = a[9] & g[1704];
assign g[3751] = b[9] & g[1704];
assign g[2729] = a[9] & g[1705];
assign g[3752] = b[9] & g[1705];
assign g[2730] = a[9] & g[1706];
assign g[3753] = b[9] & g[1706];
assign g[2731] = a[9] & g[1707];
assign g[3754] = b[9] & g[1707];
assign g[2732] = a[9] & g[1708];
assign g[3755] = b[9] & g[1708];
assign g[2733] = a[9] & g[1709];
assign g[3756] = b[9] & g[1709];
assign g[2734] = a[9] & g[1710];
assign g[3757] = b[9] & g[1710];
assign g[2735] = a[9] & g[1711];
assign g[3758] = b[9] & g[1711];
assign g[2736] = a[9] & g[1712];
assign g[3759] = b[9] & g[1712];
assign g[2737] = a[9] & g[1713];
assign g[3760] = b[9] & g[1713];
assign g[2738] = a[9] & g[1714];
assign g[3761] = b[9] & g[1714];
assign g[2739] = a[9] & g[1715];
assign g[3762] = b[9] & g[1715];
assign g[2740] = a[9] & g[1716];
assign g[3763] = b[9] & g[1716];
assign g[2741] = a[9] & g[1717];
assign g[3764] = b[9] & g[1717];
assign g[2742] = a[9] & g[1718];
assign g[3765] = b[9] & g[1718];
assign g[2743] = a[9] & g[1719];
assign g[3766] = b[9] & g[1719];
assign g[2744] = a[9] & g[1720];
assign g[3767] = b[9] & g[1720];
assign g[2745] = a[9] & g[1721];
assign g[3768] = b[9] & g[1721];
assign g[2746] = a[9] & g[1722];
assign g[3769] = b[9] & g[1722];
assign g[2747] = a[9] & g[1723];
assign g[3770] = b[9] & g[1723];
assign g[2748] = a[9] & g[1724];
assign g[3771] = b[9] & g[1724];
assign g[2749] = a[9] & g[1725];
assign g[3772] = b[9] & g[1725];
assign g[2750] = a[9] & g[1726];
assign g[3773] = b[9] & g[1726];
assign g[2751] = a[9] & g[1727];
assign g[3774] = b[9] & g[1727];
assign g[2752] = a[9] & g[1728];
assign g[3775] = b[9] & g[1728];
assign g[2753] = a[9] & g[1729];
assign g[3776] = b[9] & g[1729];
assign g[2754] = a[9] & g[1730];
assign g[3777] = b[9] & g[1730];
assign g[2755] = a[9] & g[1731];
assign g[3778] = b[9] & g[1731];
assign g[2756] = a[9] & g[1732];
assign g[3779] = b[9] & g[1732];
assign g[2757] = a[9] & g[1733];
assign g[3780] = b[9] & g[1733];
assign g[2758] = a[9] & g[1734];
assign g[3781] = b[9] & g[1734];
assign g[2759] = a[9] & g[1735];
assign g[3782] = b[9] & g[1735];
assign g[2760] = a[9] & g[1736];
assign g[3783] = b[9] & g[1736];
assign g[2761] = a[9] & g[1737];
assign g[3784] = b[9] & g[1737];
assign g[2762] = a[9] & g[1738];
assign g[3785] = b[9] & g[1738];
assign g[2763] = a[9] & g[1739];
assign g[3786] = b[9] & g[1739];
assign g[2764] = a[9] & g[1740];
assign g[3787] = b[9] & g[1740];
assign g[2765] = a[9] & g[1741];
assign g[3788] = b[9] & g[1741];
assign g[2766] = a[9] & g[1742];
assign g[3789] = b[9] & g[1742];
assign g[2767] = a[9] & g[1743];
assign g[3790] = b[9] & g[1743];
assign g[2768] = a[9] & g[1744];
assign g[3791] = b[9] & g[1744];
assign g[2769] = a[9] & g[1745];
assign g[3792] = b[9] & g[1745];
assign g[2770] = a[9] & g[1746];
assign g[3793] = b[9] & g[1746];
assign g[2771] = a[9] & g[1747];
assign g[3794] = b[9] & g[1747];
assign g[2772] = a[9] & g[1748];
assign g[3795] = b[9] & g[1748];
assign g[2773] = a[9] & g[1749];
assign g[3796] = b[9] & g[1749];
assign g[2774] = a[9] & g[1750];
assign g[3797] = b[9] & g[1750];
assign g[2775] = a[9] & g[1751];
assign g[3798] = b[9] & g[1751];
assign g[2776] = a[9] & g[1752];
assign g[3799] = b[9] & g[1752];
assign g[2777] = a[9] & g[1753];
assign g[3800] = b[9] & g[1753];
assign g[2778] = a[9] & g[1754];
assign g[3801] = b[9] & g[1754];
assign g[2779] = a[9] & g[1755];
assign g[3802] = b[9] & g[1755];
assign g[2780] = a[9] & g[1756];
assign g[3803] = b[9] & g[1756];
assign g[2781] = a[9] & g[1757];
assign g[3804] = b[9] & g[1757];
assign g[2782] = a[9] & g[1758];
assign g[3805] = b[9] & g[1758];
assign g[2783] = a[9] & g[1759];
assign g[3806] = b[9] & g[1759];
assign g[2784] = a[9] & g[1760];
assign g[3807] = b[9] & g[1760];
assign g[2785] = a[9] & g[1761];
assign g[3808] = b[9] & g[1761];
assign g[2786] = a[9] & g[1762];
assign g[3809] = b[9] & g[1762];
assign g[2787] = a[9] & g[1763];
assign g[3810] = b[9] & g[1763];
assign g[2788] = a[9] & g[1764];
assign g[3811] = b[9] & g[1764];
assign g[2789] = a[9] & g[1765];
assign g[3812] = b[9] & g[1765];
assign g[2790] = a[9] & g[1766];
assign g[3813] = b[9] & g[1766];
assign g[2791] = a[9] & g[1767];
assign g[3814] = b[9] & g[1767];
assign g[2792] = a[9] & g[1768];
assign g[3815] = b[9] & g[1768];
assign g[2793] = a[9] & g[1769];
assign g[3816] = b[9] & g[1769];
assign g[2794] = a[9] & g[1770];
assign g[3817] = b[9] & g[1770];
assign g[2795] = a[9] & g[1771];
assign g[3818] = b[9] & g[1771];
assign g[2796] = a[9] & g[1772];
assign g[3819] = b[9] & g[1772];
assign g[2797] = a[9] & g[1773];
assign g[3820] = b[9] & g[1773];
assign g[2798] = a[9] & g[1774];
assign g[3821] = b[9] & g[1774];
assign g[2799] = a[9] & g[1775];
assign g[3822] = b[9] & g[1775];
assign g[2800] = a[9] & g[1776];
assign g[3823] = b[9] & g[1776];
assign g[2801] = a[9] & g[1777];
assign g[3824] = b[9] & g[1777];
assign g[2802] = a[9] & g[1778];
assign g[3825] = b[9] & g[1778];
assign g[2803] = a[9] & g[1779];
assign g[3826] = b[9] & g[1779];
assign g[2804] = a[9] & g[1780];
assign g[3827] = b[9] & g[1780];
assign g[2805] = a[9] & g[1781];
assign g[3828] = b[9] & g[1781];
assign g[2806] = a[9] & g[1782];
assign g[3829] = b[9] & g[1782];
assign g[2807] = a[9] & g[1783];
assign g[3830] = b[9] & g[1783];
assign g[2808] = a[9] & g[1784];
assign g[3831] = b[9] & g[1784];
assign g[2809] = a[9] & g[1785];
assign g[3832] = b[9] & g[1785];
assign g[2810] = a[9] & g[1786];
assign g[3833] = b[9] & g[1786];
assign g[2811] = a[9] & g[1787];
assign g[3834] = b[9] & g[1787];
assign g[2812] = a[9] & g[1788];
assign g[3835] = b[9] & g[1788];
assign g[2813] = a[9] & g[1789];
assign g[3836] = b[9] & g[1789];
assign g[2814] = a[9] & g[1790];
assign g[3837] = b[9] & g[1790];
assign g[2815] = a[9] & g[1791];
assign g[3838] = b[9] & g[1791];
assign g[2816] = a[9] & g[1792];
assign g[3839] = b[9] & g[1792];
assign g[2817] = a[9] & g[1793];
assign g[3840] = b[9] & g[1793];
assign g[2818] = a[9] & g[1794];
assign g[3841] = b[9] & g[1794];
assign g[2819] = a[9] & g[1795];
assign g[3842] = b[9] & g[1795];
assign g[2820] = a[9] & g[1796];
assign g[3843] = b[9] & g[1796];
assign g[2821] = a[9] & g[1797];
assign g[3844] = b[9] & g[1797];
assign g[2822] = a[9] & g[1798];
assign g[3845] = b[9] & g[1798];
assign g[2823] = a[9] & g[1799];
assign g[3846] = b[9] & g[1799];
assign g[2824] = a[9] & g[1800];
assign g[3847] = b[9] & g[1800];
assign g[2825] = a[9] & g[1801];
assign g[3848] = b[9] & g[1801];
assign g[2826] = a[9] & g[1802];
assign g[3849] = b[9] & g[1802];
assign g[2827] = a[9] & g[1803];
assign g[3850] = b[9] & g[1803];
assign g[2828] = a[9] & g[1804];
assign g[3851] = b[9] & g[1804];
assign g[2829] = a[9] & g[1805];
assign g[3852] = b[9] & g[1805];
assign g[2830] = a[9] & g[1806];
assign g[3853] = b[9] & g[1806];
assign g[2831] = a[9] & g[1807];
assign g[3854] = b[9] & g[1807];
assign g[2832] = a[9] & g[1808];
assign g[3855] = b[9] & g[1808];
assign g[2833] = a[9] & g[1809];
assign g[3856] = b[9] & g[1809];
assign g[2834] = a[9] & g[1810];
assign g[3857] = b[9] & g[1810];
assign g[2835] = a[9] & g[1811];
assign g[3858] = b[9] & g[1811];
assign g[2836] = a[9] & g[1812];
assign g[3859] = b[9] & g[1812];
assign g[2837] = a[9] & g[1813];
assign g[3860] = b[9] & g[1813];
assign g[2838] = a[9] & g[1814];
assign g[3861] = b[9] & g[1814];
assign g[2839] = a[9] & g[1815];
assign g[3862] = b[9] & g[1815];
assign g[2840] = a[9] & g[1816];
assign g[3863] = b[9] & g[1816];
assign g[2841] = a[9] & g[1817];
assign g[3864] = b[9] & g[1817];
assign g[2842] = a[9] & g[1818];
assign g[3865] = b[9] & g[1818];
assign g[2843] = a[9] & g[1819];
assign g[3866] = b[9] & g[1819];
assign g[2844] = a[9] & g[1820];
assign g[3867] = b[9] & g[1820];
assign g[2845] = a[9] & g[1821];
assign g[3868] = b[9] & g[1821];
assign g[2846] = a[9] & g[1822];
assign g[3869] = b[9] & g[1822];
assign g[2847] = a[9] & g[1823];
assign g[3870] = b[9] & g[1823];
assign g[2848] = a[9] & g[1824];
assign g[3871] = b[9] & g[1824];
assign g[2849] = a[9] & g[1825];
assign g[3872] = b[9] & g[1825];
assign g[2850] = a[9] & g[1826];
assign g[3873] = b[9] & g[1826];
assign g[2851] = a[9] & g[1827];
assign g[3874] = b[9] & g[1827];
assign g[2852] = a[9] & g[1828];
assign g[3875] = b[9] & g[1828];
assign g[2853] = a[9] & g[1829];
assign g[3876] = b[9] & g[1829];
assign g[2854] = a[9] & g[1830];
assign g[3877] = b[9] & g[1830];
assign g[2855] = a[9] & g[1831];
assign g[3878] = b[9] & g[1831];
assign g[2856] = a[9] & g[1832];
assign g[3879] = b[9] & g[1832];
assign g[2857] = a[9] & g[1833];
assign g[3880] = b[9] & g[1833];
assign g[2858] = a[9] & g[1834];
assign g[3881] = b[9] & g[1834];
assign g[2859] = a[9] & g[1835];
assign g[3882] = b[9] & g[1835];
assign g[2860] = a[9] & g[1836];
assign g[3883] = b[9] & g[1836];
assign g[2861] = a[9] & g[1837];
assign g[3884] = b[9] & g[1837];
assign g[2862] = a[9] & g[1838];
assign g[3885] = b[9] & g[1838];
assign g[2863] = a[9] & g[1839];
assign g[3886] = b[9] & g[1839];
assign g[2864] = a[9] & g[1840];
assign g[3887] = b[9] & g[1840];
assign g[2865] = a[9] & g[1841];
assign g[3888] = b[9] & g[1841];
assign g[2866] = a[9] & g[1842];
assign g[3889] = b[9] & g[1842];
assign g[2867] = a[9] & g[1843];
assign g[3890] = b[9] & g[1843];
assign g[2868] = a[9] & g[1844];
assign g[3891] = b[9] & g[1844];
assign g[2869] = a[9] & g[1845];
assign g[3892] = b[9] & g[1845];
assign g[2870] = a[9] & g[1846];
assign g[3893] = b[9] & g[1846];
assign g[2871] = a[9] & g[1847];
assign g[3894] = b[9] & g[1847];
assign g[2872] = a[9] & g[1848];
assign g[3895] = b[9] & g[1848];
assign g[2873] = a[9] & g[1849];
assign g[3896] = b[9] & g[1849];
assign g[2874] = a[9] & g[1850];
assign g[3897] = b[9] & g[1850];
assign g[2875] = a[9] & g[1851];
assign g[3898] = b[9] & g[1851];
assign g[2876] = a[9] & g[1852];
assign g[3899] = b[9] & g[1852];
assign g[2877] = a[9] & g[1853];
assign g[3900] = b[9] & g[1853];
assign g[2878] = a[9] & g[1854];
assign g[3901] = b[9] & g[1854];
assign g[2879] = a[9] & g[1855];
assign g[3902] = b[9] & g[1855];
assign g[2880] = a[9] & g[1856];
assign g[3903] = b[9] & g[1856];
assign g[2881] = a[9] & g[1857];
assign g[3904] = b[9] & g[1857];
assign g[2882] = a[9] & g[1858];
assign g[3905] = b[9] & g[1858];
assign g[2883] = a[9] & g[1859];
assign g[3906] = b[9] & g[1859];
assign g[2884] = a[9] & g[1860];
assign g[3907] = b[9] & g[1860];
assign g[2885] = a[9] & g[1861];
assign g[3908] = b[9] & g[1861];
assign g[2886] = a[9] & g[1862];
assign g[3909] = b[9] & g[1862];
assign g[2887] = a[9] & g[1863];
assign g[3910] = b[9] & g[1863];
assign g[2888] = a[9] & g[1864];
assign g[3911] = b[9] & g[1864];
assign g[2889] = a[9] & g[1865];
assign g[3912] = b[9] & g[1865];
assign g[2890] = a[9] & g[1866];
assign g[3913] = b[9] & g[1866];
assign g[2891] = a[9] & g[1867];
assign g[3914] = b[9] & g[1867];
assign g[2892] = a[9] & g[1868];
assign g[3915] = b[9] & g[1868];
assign g[2893] = a[9] & g[1869];
assign g[3916] = b[9] & g[1869];
assign g[2894] = a[9] & g[1870];
assign g[3917] = b[9] & g[1870];
assign g[2895] = a[9] & g[1871];
assign g[3918] = b[9] & g[1871];
assign g[2896] = a[9] & g[1872];
assign g[3919] = b[9] & g[1872];
assign g[2897] = a[9] & g[1873];
assign g[3920] = b[9] & g[1873];
assign g[2898] = a[9] & g[1874];
assign g[3921] = b[9] & g[1874];
assign g[2899] = a[9] & g[1875];
assign g[3922] = b[9] & g[1875];
assign g[2900] = a[9] & g[1876];
assign g[3923] = b[9] & g[1876];
assign g[2901] = a[9] & g[1877];
assign g[3924] = b[9] & g[1877];
assign g[2902] = a[9] & g[1878];
assign g[3925] = b[9] & g[1878];
assign g[2903] = a[9] & g[1879];
assign g[3926] = b[9] & g[1879];
assign g[2904] = a[9] & g[1880];
assign g[3927] = b[9] & g[1880];
assign g[2905] = a[9] & g[1881];
assign g[3928] = b[9] & g[1881];
assign g[2906] = a[9] & g[1882];
assign g[3929] = b[9] & g[1882];
assign g[2907] = a[9] & g[1883];
assign g[3930] = b[9] & g[1883];
assign g[2908] = a[9] & g[1884];
assign g[3931] = b[9] & g[1884];
assign g[2909] = a[9] & g[1885];
assign g[3932] = b[9] & g[1885];
assign g[2910] = a[9] & g[1886];
assign g[3933] = b[9] & g[1886];
assign g[2911] = a[9] & g[1887];
assign g[3934] = b[9] & g[1887];
assign g[2912] = a[9] & g[1888];
assign g[3935] = b[9] & g[1888];
assign g[2913] = a[9] & g[1889];
assign g[3936] = b[9] & g[1889];
assign g[2914] = a[9] & g[1890];
assign g[3937] = b[9] & g[1890];
assign g[2915] = a[9] & g[1891];
assign g[3938] = b[9] & g[1891];
assign g[2916] = a[9] & g[1892];
assign g[3939] = b[9] & g[1892];
assign g[2917] = a[9] & g[1893];
assign g[3940] = b[9] & g[1893];
assign g[2918] = a[9] & g[1894];
assign g[3941] = b[9] & g[1894];
assign g[2919] = a[9] & g[1895];
assign g[3942] = b[9] & g[1895];
assign g[2920] = a[9] & g[1896];
assign g[3943] = b[9] & g[1896];
assign g[2921] = a[9] & g[1897];
assign g[3944] = b[9] & g[1897];
assign g[2922] = a[9] & g[1898];
assign g[3945] = b[9] & g[1898];
assign g[2923] = a[9] & g[1899];
assign g[3946] = b[9] & g[1899];
assign g[2924] = a[9] & g[1900];
assign g[3947] = b[9] & g[1900];
assign g[2925] = a[9] & g[1901];
assign g[3948] = b[9] & g[1901];
assign g[2926] = a[9] & g[1902];
assign g[3949] = b[9] & g[1902];
assign g[2927] = a[9] & g[1903];
assign g[3950] = b[9] & g[1903];
assign g[2928] = a[9] & g[1904];
assign g[3951] = b[9] & g[1904];
assign g[2929] = a[9] & g[1905];
assign g[3952] = b[9] & g[1905];
assign g[2930] = a[9] & g[1906];
assign g[3953] = b[9] & g[1906];
assign g[2931] = a[9] & g[1907];
assign g[3954] = b[9] & g[1907];
assign g[2932] = a[9] & g[1908];
assign g[3955] = b[9] & g[1908];
assign g[2933] = a[9] & g[1909];
assign g[3956] = b[9] & g[1909];
assign g[2934] = a[9] & g[1910];
assign g[3957] = b[9] & g[1910];
assign g[2935] = a[9] & g[1911];
assign g[3958] = b[9] & g[1911];
assign g[2936] = a[9] & g[1912];
assign g[3959] = b[9] & g[1912];
assign g[2937] = a[9] & g[1913];
assign g[3960] = b[9] & g[1913];
assign g[2938] = a[9] & g[1914];
assign g[3961] = b[9] & g[1914];
assign g[2939] = a[9] & g[1915];
assign g[3962] = b[9] & g[1915];
assign g[2940] = a[9] & g[1916];
assign g[3963] = b[9] & g[1916];
assign g[2941] = a[9] & g[1917];
assign g[3964] = b[9] & g[1917];
assign g[2942] = a[9] & g[1918];
assign g[3965] = b[9] & g[1918];
assign g[2943] = a[9] & g[1919];
assign g[3966] = b[9] & g[1919];
assign g[2944] = a[9] & g[1920];
assign g[3967] = b[9] & g[1920];
assign g[2945] = a[9] & g[1921];
assign g[3968] = b[9] & g[1921];
assign g[2946] = a[9] & g[1922];
assign g[3969] = b[9] & g[1922];
assign g[2947] = a[9] & g[1923];
assign g[3970] = b[9] & g[1923];
assign g[2948] = a[9] & g[1924];
assign g[3971] = b[9] & g[1924];
assign g[2949] = a[9] & g[1925];
assign g[3972] = b[9] & g[1925];
assign g[2950] = a[9] & g[1926];
assign g[3973] = b[9] & g[1926];
assign g[2951] = a[9] & g[1927];
assign g[3974] = b[9] & g[1927];
assign g[2952] = a[9] & g[1928];
assign g[3975] = b[9] & g[1928];
assign g[2953] = a[9] & g[1929];
assign g[3976] = b[9] & g[1929];
assign g[2954] = a[9] & g[1930];
assign g[3977] = b[9] & g[1930];
assign g[2955] = a[9] & g[1931];
assign g[3978] = b[9] & g[1931];
assign g[2956] = a[9] & g[1932];
assign g[3979] = b[9] & g[1932];
assign g[2957] = a[9] & g[1933];
assign g[3980] = b[9] & g[1933];
assign g[2958] = a[9] & g[1934];
assign g[3981] = b[9] & g[1934];
assign g[2959] = a[9] & g[1935];
assign g[3982] = b[9] & g[1935];
assign g[2960] = a[9] & g[1936];
assign g[3983] = b[9] & g[1936];
assign g[2961] = a[9] & g[1937];
assign g[3984] = b[9] & g[1937];
assign g[2962] = a[9] & g[1938];
assign g[3985] = b[9] & g[1938];
assign g[2963] = a[9] & g[1939];
assign g[3986] = b[9] & g[1939];
assign g[2964] = a[9] & g[1940];
assign g[3987] = b[9] & g[1940];
assign g[2965] = a[9] & g[1941];
assign g[3988] = b[9] & g[1941];
assign g[2966] = a[9] & g[1942];
assign g[3989] = b[9] & g[1942];
assign g[2967] = a[9] & g[1943];
assign g[3990] = b[9] & g[1943];
assign g[2968] = a[9] & g[1944];
assign g[3991] = b[9] & g[1944];
assign g[2969] = a[9] & g[1945];
assign g[3992] = b[9] & g[1945];
assign g[2970] = a[9] & g[1946];
assign g[3993] = b[9] & g[1946];
assign g[2971] = a[9] & g[1947];
assign g[3994] = b[9] & g[1947];
assign g[2972] = a[9] & g[1948];
assign g[3995] = b[9] & g[1948];
assign g[2973] = a[9] & g[1949];
assign g[3996] = b[9] & g[1949];
assign g[2974] = a[9] & g[1950];
assign g[3997] = b[9] & g[1950];
assign g[2975] = a[9] & g[1951];
assign g[3998] = b[9] & g[1951];
assign g[2976] = a[9] & g[1952];
assign g[3999] = b[9] & g[1952];
assign g[2977] = a[9] & g[1953];
assign g[4000] = b[9] & g[1953];
assign g[2978] = a[9] & g[1954];
assign g[4001] = b[9] & g[1954];
assign g[2979] = a[9] & g[1955];
assign g[4002] = b[9] & g[1955];
assign g[2980] = a[9] & g[1956];
assign g[4003] = b[9] & g[1956];
assign g[2981] = a[9] & g[1957];
assign g[4004] = b[9] & g[1957];
assign g[2982] = a[9] & g[1958];
assign g[4005] = b[9] & g[1958];
assign g[2983] = a[9] & g[1959];
assign g[4006] = b[9] & g[1959];
assign g[2984] = a[9] & g[1960];
assign g[4007] = b[9] & g[1960];
assign g[2985] = a[9] & g[1961];
assign g[4008] = b[9] & g[1961];
assign g[2986] = a[9] & g[1962];
assign g[4009] = b[9] & g[1962];
assign g[2987] = a[9] & g[1963];
assign g[4010] = b[9] & g[1963];
assign g[2988] = a[9] & g[1964];
assign g[4011] = b[9] & g[1964];
assign g[2989] = a[9] & g[1965];
assign g[4012] = b[9] & g[1965];
assign g[2990] = a[9] & g[1966];
assign g[4013] = b[9] & g[1966];
assign g[2991] = a[9] & g[1967];
assign g[4014] = b[9] & g[1967];
assign g[2992] = a[9] & g[1968];
assign g[4015] = b[9] & g[1968];
assign g[2993] = a[9] & g[1969];
assign g[4016] = b[9] & g[1969];
assign g[2994] = a[9] & g[1970];
assign g[4017] = b[9] & g[1970];
assign g[2995] = a[9] & g[1971];
assign g[4018] = b[9] & g[1971];
assign g[2996] = a[9] & g[1972];
assign g[4019] = b[9] & g[1972];
assign g[2997] = a[9] & g[1973];
assign g[4020] = b[9] & g[1973];
assign g[2998] = a[9] & g[1974];
assign g[4021] = b[9] & g[1974];
assign g[2999] = a[9] & g[1975];
assign g[4022] = b[9] & g[1975];
assign g[3000] = a[9] & g[1976];
assign g[4023] = b[9] & g[1976];
assign g[3001] = a[9] & g[1977];
assign g[4024] = b[9] & g[1977];
assign g[3002] = a[9] & g[1978];
assign g[4025] = b[9] & g[1978];
assign g[3003] = a[9] & g[1979];
assign g[4026] = b[9] & g[1979];
assign g[3004] = a[9] & g[1980];
assign g[4027] = b[9] & g[1980];
assign g[3005] = a[9] & g[1981];
assign g[4028] = b[9] & g[1981];
assign g[3006] = a[9] & g[1982];
assign g[4029] = b[9] & g[1982];
assign g[3007] = a[9] & g[1983];
assign g[4030] = b[9] & g[1983];
assign g[3008] = a[9] & g[1984];
assign g[4031] = b[9] & g[1984];
assign g[3009] = a[9] & g[1985];
assign g[4032] = b[9] & g[1985];
assign g[3010] = a[9] & g[1986];
assign g[4033] = b[9] & g[1986];
assign g[3011] = a[9] & g[1987];
assign g[4034] = b[9] & g[1987];
assign g[3012] = a[9] & g[1988];
assign g[4035] = b[9] & g[1988];
assign g[3013] = a[9] & g[1989];
assign g[4036] = b[9] & g[1989];
assign g[3014] = a[9] & g[1990];
assign g[4037] = b[9] & g[1990];
assign g[3015] = a[9] & g[1991];
assign g[4038] = b[9] & g[1991];
assign g[3016] = a[9] & g[1992];
assign g[4039] = b[9] & g[1992];
assign g[3017] = a[9] & g[1993];
assign g[4040] = b[9] & g[1993];
assign g[3018] = a[9] & g[1994];
assign g[4041] = b[9] & g[1994];
assign g[3019] = a[9] & g[1995];
assign g[4042] = b[9] & g[1995];
assign g[3020] = a[9] & g[1996];
assign g[4043] = b[9] & g[1996];
assign g[3021] = a[9] & g[1997];
assign g[4044] = b[9] & g[1997];
assign g[3022] = a[9] & g[1998];
assign g[4045] = b[9] & g[1998];
assign g[3023] = a[9] & g[1999];
assign g[4046] = b[9] & g[1999];
assign g[3024] = a[9] & g[2000];
assign g[4047] = b[9] & g[2000];
assign g[3025] = a[9] & g[2001];
assign g[4048] = b[9] & g[2001];
assign g[3026] = a[9] & g[2002];
assign g[4049] = b[9] & g[2002];
assign g[3027] = a[9] & g[2003];
assign g[4050] = b[9] & g[2003];
assign g[3028] = a[9] & g[2004];
assign g[4051] = b[9] & g[2004];
assign g[3029] = a[9] & g[2005];
assign g[4052] = b[9] & g[2005];
assign g[3030] = a[9] & g[2006];
assign g[4053] = b[9] & g[2006];
assign g[3031] = a[9] & g[2007];
assign g[4054] = b[9] & g[2007];
assign g[3032] = a[9] & g[2008];
assign g[4055] = b[9] & g[2008];
assign g[3033] = a[9] & g[2009];
assign g[4056] = b[9] & g[2009];
assign g[3034] = a[9] & g[2010];
assign g[4057] = b[9] & g[2010];
assign g[3035] = a[9] & g[2011];
assign g[4058] = b[9] & g[2011];
assign g[3036] = a[9] & g[2012];
assign g[4059] = b[9] & g[2012];
assign g[3037] = a[9] & g[2013];
assign g[4060] = b[9] & g[2013];
assign g[3038] = a[9] & g[2014];
assign g[4061] = b[9] & g[2014];
assign g[3039] = a[9] & g[2015];
assign g[4062] = b[9] & g[2015];
assign g[3040] = a[9] & g[2016];
assign g[4063] = b[9] & g[2016];
assign g[3041] = a[9] & g[2017];
assign g[4064] = b[9] & g[2017];
assign g[3042] = a[9] & g[2018];
assign g[4065] = b[9] & g[2018];
assign g[3043] = a[9] & g[2019];
assign g[4066] = b[9] & g[2019];
assign g[3044] = a[9] & g[2020];
assign g[4067] = b[9] & g[2020];
assign g[3045] = a[9] & g[2021];
assign g[4068] = b[9] & g[2021];
assign g[3046] = a[9] & g[2022];
assign g[4069] = b[9] & g[2022];
assign g[3047] = a[9] & g[2023];
assign g[4070] = b[9] & g[2023];
assign g[3048] = a[9] & g[2024];
assign g[4071] = b[9] & g[2024];
assign g[3049] = a[9] & g[2025];
assign g[4072] = b[9] & g[2025];
assign g[3050] = a[9] & g[2026];
assign g[4073] = b[9] & g[2026];
assign g[3051] = a[9] & g[2027];
assign g[4074] = b[9] & g[2027];
assign g[3052] = a[9] & g[2028];
assign g[4075] = b[9] & g[2028];
assign g[3053] = a[9] & g[2029];
assign g[4076] = b[9] & g[2029];
assign g[3054] = a[9] & g[2030];
assign g[4077] = b[9] & g[2030];
assign g[3055] = a[9] & g[2031];
assign g[4078] = b[9] & g[2031];
assign g[3056] = a[9] & g[2032];
assign g[4079] = b[9] & g[2032];
assign g[3057] = a[9] & g[2033];
assign g[4080] = b[9] & g[2033];
assign g[3058] = a[9] & g[2034];
assign g[4081] = b[9] & g[2034];
assign g[3059] = a[9] & g[2035];
assign g[4082] = b[9] & g[2035];
//Assigning outputs for input bit 10
assign g[4083] = a[10] & b[10];
assign g[4084] = a[10] & g[2036];
assign g[6131] = b[10] & g[2036];
assign g[4085] = a[10] & g[2037];
assign g[6132] = b[10] & g[2037];
assign g[4086] = a[10] & g[2038];
assign g[6133] = b[10] & g[2038];
assign g[4087] = a[10] & g[2039];
assign g[6134] = b[10] & g[2039];
assign g[4088] = a[10] & g[2040];
assign g[6135] = b[10] & g[2040];
assign g[4089] = a[10] & g[2041];
assign g[6136] = b[10] & g[2041];
assign g[4090] = a[10] & g[2042];
assign g[6137] = b[10] & g[2042];
assign g[4091] = a[10] & g[2043];
assign g[6138] = b[10] & g[2043];
assign g[4092] = a[10] & g[2044];
assign g[6139] = b[10] & g[2044];
assign g[4093] = a[10] & g[2045];
assign g[6140] = b[10] & g[2045];
assign g[4094] = a[10] & g[2046];
assign g[6141] = b[10] & g[2046];
assign g[4095] = a[10] & g[2047];
assign g[6142] = b[10] & g[2047];
assign g[4096] = a[10] & g[2048];
assign g[6143] = b[10] & g[2048];
assign g[4097] = a[10] & g[2049];
assign g[6144] = b[10] & g[2049];
assign g[4098] = a[10] & g[2050];
assign g[6145] = b[10] & g[2050];
assign g[4099] = a[10] & g[2051];
assign g[6146] = b[10] & g[2051];
assign g[4100] = a[10] & g[2052];
assign g[6147] = b[10] & g[2052];
assign g[4101] = a[10] & g[2053];
assign g[6148] = b[10] & g[2053];
assign g[4102] = a[10] & g[2054];
assign g[6149] = b[10] & g[2054];
assign g[4103] = a[10] & g[2055];
assign g[6150] = b[10] & g[2055];
assign g[4104] = a[10] & g[2056];
assign g[6151] = b[10] & g[2056];
assign g[4105] = a[10] & g[2057];
assign g[6152] = b[10] & g[2057];
assign g[4106] = a[10] & g[2058];
assign g[6153] = b[10] & g[2058];
assign g[4107] = a[10] & g[2059];
assign g[6154] = b[10] & g[2059];
assign g[4108] = a[10] & g[2060];
assign g[6155] = b[10] & g[2060];
assign g[4109] = a[10] & g[2061];
assign g[6156] = b[10] & g[2061];
assign g[4110] = a[10] & g[2062];
assign g[6157] = b[10] & g[2062];
assign g[4111] = a[10] & g[2063];
assign g[6158] = b[10] & g[2063];
assign g[4112] = a[10] & g[2064];
assign g[6159] = b[10] & g[2064];
assign g[4113] = a[10] & g[2065];
assign g[6160] = b[10] & g[2065];
assign g[4114] = a[10] & g[2066];
assign g[6161] = b[10] & g[2066];
assign g[4115] = a[10] & g[2067];
assign g[6162] = b[10] & g[2067];
assign g[4116] = a[10] & g[2068];
assign g[6163] = b[10] & g[2068];
assign g[4117] = a[10] & g[2069];
assign g[6164] = b[10] & g[2069];
assign g[4118] = a[10] & g[2070];
assign g[6165] = b[10] & g[2070];
assign g[4119] = a[10] & g[2071];
assign g[6166] = b[10] & g[2071];
assign g[4120] = a[10] & g[2072];
assign g[6167] = b[10] & g[2072];
assign g[4121] = a[10] & g[2073];
assign g[6168] = b[10] & g[2073];
assign g[4122] = a[10] & g[2074];
assign g[6169] = b[10] & g[2074];
assign g[4123] = a[10] & g[2075];
assign g[6170] = b[10] & g[2075];
assign g[4124] = a[10] & g[2076];
assign g[6171] = b[10] & g[2076];
assign g[4125] = a[10] & g[2077];
assign g[6172] = b[10] & g[2077];
assign g[4126] = a[10] & g[2078];
assign g[6173] = b[10] & g[2078];
assign g[4127] = a[10] & g[2079];
assign g[6174] = b[10] & g[2079];
assign g[4128] = a[10] & g[2080];
assign g[6175] = b[10] & g[2080];
assign g[4129] = a[10] & g[2081];
assign g[6176] = b[10] & g[2081];
assign g[4130] = a[10] & g[2082];
assign g[6177] = b[10] & g[2082];
assign g[4131] = a[10] & g[2083];
assign g[6178] = b[10] & g[2083];
assign g[4132] = a[10] & g[2084];
assign g[6179] = b[10] & g[2084];
assign g[4133] = a[10] & g[2085];
assign g[6180] = b[10] & g[2085];
assign g[4134] = a[10] & g[2086];
assign g[6181] = b[10] & g[2086];
assign g[4135] = a[10] & g[2087];
assign g[6182] = b[10] & g[2087];
assign g[4136] = a[10] & g[2088];
assign g[6183] = b[10] & g[2088];
assign g[4137] = a[10] & g[2089];
assign g[6184] = b[10] & g[2089];
assign g[4138] = a[10] & g[2090];
assign g[6185] = b[10] & g[2090];
assign g[4139] = a[10] & g[2091];
assign g[6186] = b[10] & g[2091];
assign g[4140] = a[10] & g[2092];
assign g[6187] = b[10] & g[2092];
assign g[4141] = a[10] & g[2093];
assign g[6188] = b[10] & g[2093];
assign g[4142] = a[10] & g[2094];
assign g[6189] = b[10] & g[2094];
assign g[4143] = a[10] & g[2095];
assign g[6190] = b[10] & g[2095];
assign g[4144] = a[10] & g[2096];
assign g[6191] = b[10] & g[2096];
assign g[4145] = a[10] & g[2097];
assign g[6192] = b[10] & g[2097];
assign g[4146] = a[10] & g[2098];
assign g[6193] = b[10] & g[2098];
assign g[4147] = a[10] & g[2099];
assign g[6194] = b[10] & g[2099];
assign g[4148] = a[10] & g[2100];
assign g[6195] = b[10] & g[2100];
assign g[4149] = a[10] & g[2101];
assign g[6196] = b[10] & g[2101];
assign g[4150] = a[10] & g[2102];
assign g[6197] = b[10] & g[2102];
assign g[4151] = a[10] & g[2103];
assign g[6198] = b[10] & g[2103];
assign g[4152] = a[10] & g[2104];
assign g[6199] = b[10] & g[2104];
assign g[4153] = a[10] & g[2105];
assign g[6200] = b[10] & g[2105];
assign g[4154] = a[10] & g[2106];
assign g[6201] = b[10] & g[2106];
assign g[4155] = a[10] & g[2107];
assign g[6202] = b[10] & g[2107];
assign g[4156] = a[10] & g[2108];
assign g[6203] = b[10] & g[2108];
assign g[4157] = a[10] & g[2109];
assign g[6204] = b[10] & g[2109];
assign g[4158] = a[10] & g[2110];
assign g[6205] = b[10] & g[2110];
assign g[4159] = a[10] & g[2111];
assign g[6206] = b[10] & g[2111];
assign g[4160] = a[10] & g[2112];
assign g[6207] = b[10] & g[2112];
assign g[4161] = a[10] & g[2113];
assign g[6208] = b[10] & g[2113];
assign g[4162] = a[10] & g[2114];
assign g[6209] = b[10] & g[2114];
assign g[4163] = a[10] & g[2115];
assign g[6210] = b[10] & g[2115];
assign g[4164] = a[10] & g[2116];
assign g[6211] = b[10] & g[2116];
assign g[4165] = a[10] & g[2117];
assign g[6212] = b[10] & g[2117];
assign g[4166] = a[10] & g[2118];
assign g[6213] = b[10] & g[2118];
assign g[4167] = a[10] & g[2119];
assign g[6214] = b[10] & g[2119];
assign g[4168] = a[10] & g[2120];
assign g[6215] = b[10] & g[2120];
assign g[4169] = a[10] & g[2121];
assign g[6216] = b[10] & g[2121];
assign g[4170] = a[10] & g[2122];
assign g[6217] = b[10] & g[2122];
assign g[4171] = a[10] & g[2123];
assign g[6218] = b[10] & g[2123];
assign g[4172] = a[10] & g[2124];
assign g[6219] = b[10] & g[2124];
assign g[4173] = a[10] & g[2125];
assign g[6220] = b[10] & g[2125];
assign g[4174] = a[10] & g[2126];
assign g[6221] = b[10] & g[2126];
assign g[4175] = a[10] & g[2127];
assign g[6222] = b[10] & g[2127];
assign g[4176] = a[10] & g[2128];
assign g[6223] = b[10] & g[2128];
assign g[4177] = a[10] & g[2129];
assign g[6224] = b[10] & g[2129];
assign g[4178] = a[10] & g[2130];
assign g[6225] = b[10] & g[2130];
assign g[4179] = a[10] & g[2131];
assign g[6226] = b[10] & g[2131];
assign g[4180] = a[10] & g[2132];
assign g[6227] = b[10] & g[2132];
assign g[4181] = a[10] & g[2133];
assign g[6228] = b[10] & g[2133];
assign g[4182] = a[10] & g[2134];
assign g[6229] = b[10] & g[2134];
assign g[4183] = a[10] & g[2135];
assign g[6230] = b[10] & g[2135];
assign g[4184] = a[10] & g[2136];
assign g[6231] = b[10] & g[2136];
assign g[4185] = a[10] & g[2137];
assign g[6232] = b[10] & g[2137];
assign g[4186] = a[10] & g[2138];
assign g[6233] = b[10] & g[2138];
assign g[4187] = a[10] & g[2139];
assign g[6234] = b[10] & g[2139];
assign g[4188] = a[10] & g[2140];
assign g[6235] = b[10] & g[2140];
assign g[4189] = a[10] & g[2141];
assign g[6236] = b[10] & g[2141];
assign g[4190] = a[10] & g[2142];
assign g[6237] = b[10] & g[2142];
assign g[4191] = a[10] & g[2143];
assign g[6238] = b[10] & g[2143];
assign g[4192] = a[10] & g[2144];
assign g[6239] = b[10] & g[2144];
assign g[4193] = a[10] & g[2145];
assign g[6240] = b[10] & g[2145];
assign g[4194] = a[10] & g[2146];
assign g[6241] = b[10] & g[2146];
assign g[4195] = a[10] & g[2147];
assign g[6242] = b[10] & g[2147];
assign g[4196] = a[10] & g[2148];
assign g[6243] = b[10] & g[2148];
assign g[4197] = a[10] & g[2149];
assign g[6244] = b[10] & g[2149];
assign g[4198] = a[10] & g[2150];
assign g[6245] = b[10] & g[2150];
assign g[4199] = a[10] & g[2151];
assign g[6246] = b[10] & g[2151];
assign g[4200] = a[10] & g[2152];
assign g[6247] = b[10] & g[2152];
assign g[4201] = a[10] & g[2153];
assign g[6248] = b[10] & g[2153];
assign g[4202] = a[10] & g[2154];
assign g[6249] = b[10] & g[2154];
assign g[4203] = a[10] & g[2155];
assign g[6250] = b[10] & g[2155];
assign g[4204] = a[10] & g[2156];
assign g[6251] = b[10] & g[2156];
assign g[4205] = a[10] & g[2157];
assign g[6252] = b[10] & g[2157];
assign g[4206] = a[10] & g[2158];
assign g[6253] = b[10] & g[2158];
assign g[4207] = a[10] & g[2159];
assign g[6254] = b[10] & g[2159];
assign g[4208] = a[10] & g[2160];
assign g[6255] = b[10] & g[2160];
assign g[4209] = a[10] & g[2161];
assign g[6256] = b[10] & g[2161];
assign g[4210] = a[10] & g[2162];
assign g[6257] = b[10] & g[2162];
assign g[4211] = a[10] & g[2163];
assign g[6258] = b[10] & g[2163];
assign g[4212] = a[10] & g[2164];
assign g[6259] = b[10] & g[2164];
assign g[4213] = a[10] & g[2165];
assign g[6260] = b[10] & g[2165];
assign g[4214] = a[10] & g[2166];
assign g[6261] = b[10] & g[2166];
assign g[4215] = a[10] & g[2167];
assign g[6262] = b[10] & g[2167];
assign g[4216] = a[10] & g[2168];
assign g[6263] = b[10] & g[2168];
assign g[4217] = a[10] & g[2169];
assign g[6264] = b[10] & g[2169];
assign g[4218] = a[10] & g[2170];
assign g[6265] = b[10] & g[2170];
assign g[4219] = a[10] & g[2171];
assign g[6266] = b[10] & g[2171];
assign g[4220] = a[10] & g[2172];
assign g[6267] = b[10] & g[2172];
assign g[4221] = a[10] & g[2173];
assign g[6268] = b[10] & g[2173];
assign g[4222] = a[10] & g[2174];
assign g[6269] = b[10] & g[2174];
assign g[4223] = a[10] & g[2175];
assign g[6270] = b[10] & g[2175];
assign g[4224] = a[10] & g[2176];
assign g[6271] = b[10] & g[2176];
assign g[4225] = a[10] & g[2177];
assign g[6272] = b[10] & g[2177];
assign g[4226] = a[10] & g[2178];
assign g[6273] = b[10] & g[2178];
assign g[4227] = a[10] & g[2179];
assign g[6274] = b[10] & g[2179];
assign g[4228] = a[10] & g[2180];
assign g[6275] = b[10] & g[2180];
assign g[4229] = a[10] & g[2181];
assign g[6276] = b[10] & g[2181];
assign g[4230] = a[10] & g[2182];
assign g[6277] = b[10] & g[2182];
assign g[4231] = a[10] & g[2183];
assign g[6278] = b[10] & g[2183];
assign g[4232] = a[10] & g[2184];
assign g[6279] = b[10] & g[2184];
assign g[4233] = a[10] & g[2185];
assign g[6280] = b[10] & g[2185];
assign g[4234] = a[10] & g[2186];
assign g[6281] = b[10] & g[2186];
assign g[4235] = a[10] & g[2187];
assign g[6282] = b[10] & g[2187];
assign g[4236] = a[10] & g[2188];
assign g[6283] = b[10] & g[2188];
assign g[4237] = a[10] & g[2189];
assign g[6284] = b[10] & g[2189];
assign g[4238] = a[10] & g[2190];
assign g[6285] = b[10] & g[2190];
assign g[4239] = a[10] & g[2191];
assign g[6286] = b[10] & g[2191];
assign g[4240] = a[10] & g[2192];
assign g[6287] = b[10] & g[2192];
assign g[4241] = a[10] & g[2193];
assign g[6288] = b[10] & g[2193];
assign g[4242] = a[10] & g[2194];
assign g[6289] = b[10] & g[2194];
assign g[4243] = a[10] & g[2195];
assign g[6290] = b[10] & g[2195];
assign g[4244] = a[10] & g[2196];
assign g[6291] = b[10] & g[2196];
assign g[4245] = a[10] & g[2197];
assign g[6292] = b[10] & g[2197];
assign g[4246] = a[10] & g[2198];
assign g[6293] = b[10] & g[2198];
assign g[4247] = a[10] & g[2199];
assign g[6294] = b[10] & g[2199];
assign g[4248] = a[10] & g[2200];
assign g[6295] = b[10] & g[2200];
assign g[4249] = a[10] & g[2201];
assign g[6296] = b[10] & g[2201];
assign g[4250] = a[10] & g[2202];
assign g[6297] = b[10] & g[2202];
assign g[4251] = a[10] & g[2203];
assign g[6298] = b[10] & g[2203];
assign g[4252] = a[10] & g[2204];
assign g[6299] = b[10] & g[2204];
assign g[4253] = a[10] & g[2205];
assign g[6300] = b[10] & g[2205];
assign g[4254] = a[10] & g[2206];
assign g[6301] = b[10] & g[2206];
assign g[4255] = a[10] & g[2207];
assign g[6302] = b[10] & g[2207];
assign g[4256] = a[10] & g[2208];
assign g[6303] = b[10] & g[2208];
assign g[4257] = a[10] & g[2209];
assign g[6304] = b[10] & g[2209];
assign g[4258] = a[10] & g[2210];
assign g[6305] = b[10] & g[2210];
assign g[4259] = a[10] & g[2211];
assign g[6306] = b[10] & g[2211];
assign g[4260] = a[10] & g[2212];
assign g[6307] = b[10] & g[2212];
assign g[4261] = a[10] & g[2213];
assign g[6308] = b[10] & g[2213];
assign g[4262] = a[10] & g[2214];
assign g[6309] = b[10] & g[2214];
assign g[4263] = a[10] & g[2215];
assign g[6310] = b[10] & g[2215];
assign g[4264] = a[10] & g[2216];
assign g[6311] = b[10] & g[2216];
assign g[4265] = a[10] & g[2217];
assign g[6312] = b[10] & g[2217];
assign g[4266] = a[10] & g[2218];
assign g[6313] = b[10] & g[2218];
assign g[4267] = a[10] & g[2219];
assign g[6314] = b[10] & g[2219];
assign g[4268] = a[10] & g[2220];
assign g[6315] = b[10] & g[2220];
assign g[4269] = a[10] & g[2221];
assign g[6316] = b[10] & g[2221];
assign g[4270] = a[10] & g[2222];
assign g[6317] = b[10] & g[2222];
assign g[4271] = a[10] & g[2223];
assign g[6318] = b[10] & g[2223];
assign g[4272] = a[10] & g[2224];
assign g[6319] = b[10] & g[2224];
assign g[4273] = a[10] & g[2225];
assign g[6320] = b[10] & g[2225];
assign g[4274] = a[10] & g[2226];
assign g[6321] = b[10] & g[2226];
assign g[4275] = a[10] & g[2227];
assign g[6322] = b[10] & g[2227];
assign g[4276] = a[10] & g[2228];
assign g[6323] = b[10] & g[2228];
assign g[4277] = a[10] & g[2229];
assign g[6324] = b[10] & g[2229];
assign g[4278] = a[10] & g[2230];
assign g[6325] = b[10] & g[2230];
assign g[4279] = a[10] & g[2231];
assign g[6326] = b[10] & g[2231];
assign g[4280] = a[10] & g[2232];
assign g[6327] = b[10] & g[2232];
assign g[4281] = a[10] & g[2233];
assign g[6328] = b[10] & g[2233];
assign g[4282] = a[10] & g[2234];
assign g[6329] = b[10] & g[2234];
assign g[4283] = a[10] & g[2235];
assign g[6330] = b[10] & g[2235];
assign g[4284] = a[10] & g[2236];
assign g[6331] = b[10] & g[2236];
assign g[4285] = a[10] & g[2237];
assign g[6332] = b[10] & g[2237];
assign g[4286] = a[10] & g[2238];
assign g[6333] = b[10] & g[2238];
assign g[4287] = a[10] & g[2239];
assign g[6334] = b[10] & g[2239];
assign g[4288] = a[10] & g[2240];
assign g[6335] = b[10] & g[2240];
assign g[4289] = a[10] & g[2241];
assign g[6336] = b[10] & g[2241];
assign g[4290] = a[10] & g[2242];
assign g[6337] = b[10] & g[2242];
assign g[4291] = a[10] & g[2243];
assign g[6338] = b[10] & g[2243];
assign g[4292] = a[10] & g[2244];
assign g[6339] = b[10] & g[2244];
assign g[4293] = a[10] & g[2245];
assign g[6340] = b[10] & g[2245];
assign g[4294] = a[10] & g[2246];
assign g[6341] = b[10] & g[2246];
assign g[4295] = a[10] & g[2247];
assign g[6342] = b[10] & g[2247];
assign g[4296] = a[10] & g[2248];
assign g[6343] = b[10] & g[2248];
assign g[4297] = a[10] & g[2249];
assign g[6344] = b[10] & g[2249];
assign g[4298] = a[10] & g[2250];
assign g[6345] = b[10] & g[2250];
assign g[4299] = a[10] & g[2251];
assign g[6346] = b[10] & g[2251];
assign g[4300] = a[10] & g[2252];
assign g[6347] = b[10] & g[2252];
assign g[4301] = a[10] & g[2253];
assign g[6348] = b[10] & g[2253];
assign g[4302] = a[10] & g[2254];
assign g[6349] = b[10] & g[2254];
assign g[4303] = a[10] & g[2255];
assign g[6350] = b[10] & g[2255];
assign g[4304] = a[10] & g[2256];
assign g[6351] = b[10] & g[2256];
assign g[4305] = a[10] & g[2257];
assign g[6352] = b[10] & g[2257];
assign g[4306] = a[10] & g[2258];
assign g[6353] = b[10] & g[2258];
assign g[4307] = a[10] & g[2259];
assign g[6354] = b[10] & g[2259];
assign g[4308] = a[10] & g[2260];
assign g[6355] = b[10] & g[2260];
assign g[4309] = a[10] & g[2261];
assign g[6356] = b[10] & g[2261];
assign g[4310] = a[10] & g[2262];
assign g[6357] = b[10] & g[2262];
assign g[4311] = a[10] & g[2263];
assign g[6358] = b[10] & g[2263];
assign g[4312] = a[10] & g[2264];
assign g[6359] = b[10] & g[2264];
assign g[4313] = a[10] & g[2265];
assign g[6360] = b[10] & g[2265];
assign g[4314] = a[10] & g[2266];
assign g[6361] = b[10] & g[2266];
assign g[4315] = a[10] & g[2267];
assign g[6362] = b[10] & g[2267];
assign g[4316] = a[10] & g[2268];
assign g[6363] = b[10] & g[2268];
assign g[4317] = a[10] & g[2269];
assign g[6364] = b[10] & g[2269];
assign g[4318] = a[10] & g[2270];
assign g[6365] = b[10] & g[2270];
assign g[4319] = a[10] & g[2271];
assign g[6366] = b[10] & g[2271];
assign g[4320] = a[10] & g[2272];
assign g[6367] = b[10] & g[2272];
assign g[4321] = a[10] & g[2273];
assign g[6368] = b[10] & g[2273];
assign g[4322] = a[10] & g[2274];
assign g[6369] = b[10] & g[2274];
assign g[4323] = a[10] & g[2275];
assign g[6370] = b[10] & g[2275];
assign g[4324] = a[10] & g[2276];
assign g[6371] = b[10] & g[2276];
assign g[4325] = a[10] & g[2277];
assign g[6372] = b[10] & g[2277];
assign g[4326] = a[10] & g[2278];
assign g[6373] = b[10] & g[2278];
assign g[4327] = a[10] & g[2279];
assign g[6374] = b[10] & g[2279];
assign g[4328] = a[10] & g[2280];
assign g[6375] = b[10] & g[2280];
assign g[4329] = a[10] & g[2281];
assign g[6376] = b[10] & g[2281];
assign g[4330] = a[10] & g[2282];
assign g[6377] = b[10] & g[2282];
assign g[4331] = a[10] & g[2283];
assign g[6378] = b[10] & g[2283];
assign g[4332] = a[10] & g[2284];
assign g[6379] = b[10] & g[2284];
assign g[4333] = a[10] & g[2285];
assign g[6380] = b[10] & g[2285];
assign g[4334] = a[10] & g[2286];
assign g[6381] = b[10] & g[2286];
assign g[4335] = a[10] & g[2287];
assign g[6382] = b[10] & g[2287];
assign g[4336] = a[10] & g[2288];
assign g[6383] = b[10] & g[2288];
assign g[4337] = a[10] & g[2289];
assign g[6384] = b[10] & g[2289];
assign g[4338] = a[10] & g[2290];
assign g[6385] = b[10] & g[2290];
assign g[4339] = a[10] & g[2291];
assign g[6386] = b[10] & g[2291];
assign g[4340] = a[10] & g[2292];
assign g[6387] = b[10] & g[2292];
assign g[4341] = a[10] & g[2293];
assign g[6388] = b[10] & g[2293];
assign g[4342] = a[10] & g[2294];
assign g[6389] = b[10] & g[2294];
assign g[4343] = a[10] & g[2295];
assign g[6390] = b[10] & g[2295];
assign g[4344] = a[10] & g[2296];
assign g[6391] = b[10] & g[2296];
assign g[4345] = a[10] & g[2297];
assign g[6392] = b[10] & g[2297];
assign g[4346] = a[10] & g[2298];
assign g[6393] = b[10] & g[2298];
assign g[4347] = a[10] & g[2299];
assign g[6394] = b[10] & g[2299];
assign g[4348] = a[10] & g[2300];
assign g[6395] = b[10] & g[2300];
assign g[4349] = a[10] & g[2301];
assign g[6396] = b[10] & g[2301];
assign g[4350] = a[10] & g[2302];
assign g[6397] = b[10] & g[2302];
assign g[4351] = a[10] & g[2303];
assign g[6398] = b[10] & g[2303];
assign g[4352] = a[10] & g[2304];
assign g[6399] = b[10] & g[2304];
assign g[4353] = a[10] & g[2305];
assign g[6400] = b[10] & g[2305];
assign g[4354] = a[10] & g[2306];
assign g[6401] = b[10] & g[2306];
assign g[4355] = a[10] & g[2307];
assign g[6402] = b[10] & g[2307];
assign g[4356] = a[10] & g[2308];
assign g[6403] = b[10] & g[2308];
assign g[4357] = a[10] & g[2309];
assign g[6404] = b[10] & g[2309];
assign g[4358] = a[10] & g[2310];
assign g[6405] = b[10] & g[2310];
assign g[4359] = a[10] & g[2311];
assign g[6406] = b[10] & g[2311];
assign g[4360] = a[10] & g[2312];
assign g[6407] = b[10] & g[2312];
assign g[4361] = a[10] & g[2313];
assign g[6408] = b[10] & g[2313];
assign g[4362] = a[10] & g[2314];
assign g[6409] = b[10] & g[2314];
assign g[4363] = a[10] & g[2315];
assign g[6410] = b[10] & g[2315];
assign g[4364] = a[10] & g[2316];
assign g[6411] = b[10] & g[2316];
assign g[4365] = a[10] & g[2317];
assign g[6412] = b[10] & g[2317];
assign g[4366] = a[10] & g[2318];
assign g[6413] = b[10] & g[2318];
assign g[4367] = a[10] & g[2319];
assign g[6414] = b[10] & g[2319];
assign g[4368] = a[10] & g[2320];
assign g[6415] = b[10] & g[2320];
assign g[4369] = a[10] & g[2321];
assign g[6416] = b[10] & g[2321];
assign g[4370] = a[10] & g[2322];
assign g[6417] = b[10] & g[2322];
assign g[4371] = a[10] & g[2323];
assign g[6418] = b[10] & g[2323];
assign g[4372] = a[10] & g[2324];
assign g[6419] = b[10] & g[2324];
assign g[4373] = a[10] & g[2325];
assign g[6420] = b[10] & g[2325];
assign g[4374] = a[10] & g[2326];
assign g[6421] = b[10] & g[2326];
assign g[4375] = a[10] & g[2327];
assign g[6422] = b[10] & g[2327];
assign g[4376] = a[10] & g[2328];
assign g[6423] = b[10] & g[2328];
assign g[4377] = a[10] & g[2329];
assign g[6424] = b[10] & g[2329];
assign g[4378] = a[10] & g[2330];
assign g[6425] = b[10] & g[2330];
assign g[4379] = a[10] & g[2331];
assign g[6426] = b[10] & g[2331];
assign g[4380] = a[10] & g[2332];
assign g[6427] = b[10] & g[2332];
assign g[4381] = a[10] & g[2333];
assign g[6428] = b[10] & g[2333];
assign g[4382] = a[10] & g[2334];
assign g[6429] = b[10] & g[2334];
assign g[4383] = a[10] & g[2335];
assign g[6430] = b[10] & g[2335];
assign g[4384] = a[10] & g[2336];
assign g[6431] = b[10] & g[2336];
assign g[4385] = a[10] & g[2337];
assign g[6432] = b[10] & g[2337];
assign g[4386] = a[10] & g[2338];
assign g[6433] = b[10] & g[2338];
assign g[4387] = a[10] & g[2339];
assign g[6434] = b[10] & g[2339];
assign g[4388] = a[10] & g[2340];
assign g[6435] = b[10] & g[2340];
assign g[4389] = a[10] & g[2341];
assign g[6436] = b[10] & g[2341];
assign g[4390] = a[10] & g[2342];
assign g[6437] = b[10] & g[2342];
assign g[4391] = a[10] & g[2343];
assign g[6438] = b[10] & g[2343];
assign g[4392] = a[10] & g[2344];
assign g[6439] = b[10] & g[2344];
assign g[4393] = a[10] & g[2345];
assign g[6440] = b[10] & g[2345];
assign g[4394] = a[10] & g[2346];
assign g[6441] = b[10] & g[2346];
assign g[4395] = a[10] & g[2347];
assign g[6442] = b[10] & g[2347];
assign g[4396] = a[10] & g[2348];
assign g[6443] = b[10] & g[2348];
assign g[4397] = a[10] & g[2349];
assign g[6444] = b[10] & g[2349];
assign g[4398] = a[10] & g[2350];
assign g[6445] = b[10] & g[2350];
assign g[4399] = a[10] & g[2351];
assign g[6446] = b[10] & g[2351];
assign g[4400] = a[10] & g[2352];
assign g[6447] = b[10] & g[2352];
assign g[4401] = a[10] & g[2353];
assign g[6448] = b[10] & g[2353];
assign g[4402] = a[10] & g[2354];
assign g[6449] = b[10] & g[2354];
assign g[4403] = a[10] & g[2355];
assign g[6450] = b[10] & g[2355];
assign g[4404] = a[10] & g[2356];
assign g[6451] = b[10] & g[2356];
assign g[4405] = a[10] & g[2357];
assign g[6452] = b[10] & g[2357];
assign g[4406] = a[10] & g[2358];
assign g[6453] = b[10] & g[2358];
assign g[4407] = a[10] & g[2359];
assign g[6454] = b[10] & g[2359];
assign g[4408] = a[10] & g[2360];
assign g[6455] = b[10] & g[2360];
assign g[4409] = a[10] & g[2361];
assign g[6456] = b[10] & g[2361];
assign g[4410] = a[10] & g[2362];
assign g[6457] = b[10] & g[2362];
assign g[4411] = a[10] & g[2363];
assign g[6458] = b[10] & g[2363];
assign g[4412] = a[10] & g[2364];
assign g[6459] = b[10] & g[2364];
assign g[4413] = a[10] & g[2365];
assign g[6460] = b[10] & g[2365];
assign g[4414] = a[10] & g[2366];
assign g[6461] = b[10] & g[2366];
assign g[4415] = a[10] & g[2367];
assign g[6462] = b[10] & g[2367];
assign g[4416] = a[10] & g[2368];
assign g[6463] = b[10] & g[2368];
assign g[4417] = a[10] & g[2369];
assign g[6464] = b[10] & g[2369];
assign g[4418] = a[10] & g[2370];
assign g[6465] = b[10] & g[2370];
assign g[4419] = a[10] & g[2371];
assign g[6466] = b[10] & g[2371];
assign g[4420] = a[10] & g[2372];
assign g[6467] = b[10] & g[2372];
assign g[4421] = a[10] & g[2373];
assign g[6468] = b[10] & g[2373];
assign g[4422] = a[10] & g[2374];
assign g[6469] = b[10] & g[2374];
assign g[4423] = a[10] & g[2375];
assign g[6470] = b[10] & g[2375];
assign g[4424] = a[10] & g[2376];
assign g[6471] = b[10] & g[2376];
assign g[4425] = a[10] & g[2377];
assign g[6472] = b[10] & g[2377];
assign g[4426] = a[10] & g[2378];
assign g[6473] = b[10] & g[2378];
assign g[4427] = a[10] & g[2379];
assign g[6474] = b[10] & g[2379];
assign g[4428] = a[10] & g[2380];
assign g[6475] = b[10] & g[2380];
assign g[4429] = a[10] & g[2381];
assign g[6476] = b[10] & g[2381];
assign g[4430] = a[10] & g[2382];
assign g[6477] = b[10] & g[2382];
assign g[4431] = a[10] & g[2383];
assign g[6478] = b[10] & g[2383];
assign g[4432] = a[10] & g[2384];
assign g[6479] = b[10] & g[2384];
assign g[4433] = a[10] & g[2385];
assign g[6480] = b[10] & g[2385];
assign g[4434] = a[10] & g[2386];
assign g[6481] = b[10] & g[2386];
assign g[4435] = a[10] & g[2387];
assign g[6482] = b[10] & g[2387];
assign g[4436] = a[10] & g[2388];
assign g[6483] = b[10] & g[2388];
assign g[4437] = a[10] & g[2389];
assign g[6484] = b[10] & g[2389];
assign g[4438] = a[10] & g[2390];
assign g[6485] = b[10] & g[2390];
assign g[4439] = a[10] & g[2391];
assign g[6486] = b[10] & g[2391];
assign g[4440] = a[10] & g[2392];
assign g[6487] = b[10] & g[2392];
assign g[4441] = a[10] & g[2393];
assign g[6488] = b[10] & g[2393];
assign g[4442] = a[10] & g[2394];
assign g[6489] = b[10] & g[2394];
assign g[4443] = a[10] & g[2395];
assign g[6490] = b[10] & g[2395];
assign g[4444] = a[10] & g[2396];
assign g[6491] = b[10] & g[2396];
assign g[4445] = a[10] & g[2397];
assign g[6492] = b[10] & g[2397];
assign g[4446] = a[10] & g[2398];
assign g[6493] = b[10] & g[2398];
assign g[4447] = a[10] & g[2399];
assign g[6494] = b[10] & g[2399];
assign g[4448] = a[10] & g[2400];
assign g[6495] = b[10] & g[2400];
assign g[4449] = a[10] & g[2401];
assign g[6496] = b[10] & g[2401];
assign g[4450] = a[10] & g[2402];
assign g[6497] = b[10] & g[2402];
assign g[4451] = a[10] & g[2403];
assign g[6498] = b[10] & g[2403];
assign g[4452] = a[10] & g[2404];
assign g[6499] = b[10] & g[2404];
assign g[4453] = a[10] & g[2405];
assign g[6500] = b[10] & g[2405];
assign g[4454] = a[10] & g[2406];
assign g[6501] = b[10] & g[2406];
assign g[4455] = a[10] & g[2407];
assign g[6502] = b[10] & g[2407];
assign g[4456] = a[10] & g[2408];
assign g[6503] = b[10] & g[2408];
assign g[4457] = a[10] & g[2409];
assign g[6504] = b[10] & g[2409];
assign g[4458] = a[10] & g[2410];
assign g[6505] = b[10] & g[2410];
assign g[4459] = a[10] & g[2411];
assign g[6506] = b[10] & g[2411];
assign g[4460] = a[10] & g[2412];
assign g[6507] = b[10] & g[2412];
assign g[4461] = a[10] & g[2413];
assign g[6508] = b[10] & g[2413];
assign g[4462] = a[10] & g[2414];
assign g[6509] = b[10] & g[2414];
assign g[4463] = a[10] & g[2415];
assign g[6510] = b[10] & g[2415];
assign g[4464] = a[10] & g[2416];
assign g[6511] = b[10] & g[2416];
assign g[4465] = a[10] & g[2417];
assign g[6512] = b[10] & g[2417];
assign g[4466] = a[10] & g[2418];
assign g[6513] = b[10] & g[2418];
assign g[4467] = a[10] & g[2419];
assign g[6514] = b[10] & g[2419];
assign g[4468] = a[10] & g[2420];
assign g[6515] = b[10] & g[2420];
assign g[4469] = a[10] & g[2421];
assign g[6516] = b[10] & g[2421];
assign g[4470] = a[10] & g[2422];
assign g[6517] = b[10] & g[2422];
assign g[4471] = a[10] & g[2423];
assign g[6518] = b[10] & g[2423];
assign g[4472] = a[10] & g[2424];
assign g[6519] = b[10] & g[2424];
assign g[4473] = a[10] & g[2425];
assign g[6520] = b[10] & g[2425];
assign g[4474] = a[10] & g[2426];
assign g[6521] = b[10] & g[2426];
assign g[4475] = a[10] & g[2427];
assign g[6522] = b[10] & g[2427];
assign g[4476] = a[10] & g[2428];
assign g[6523] = b[10] & g[2428];
assign g[4477] = a[10] & g[2429];
assign g[6524] = b[10] & g[2429];
assign g[4478] = a[10] & g[2430];
assign g[6525] = b[10] & g[2430];
assign g[4479] = a[10] & g[2431];
assign g[6526] = b[10] & g[2431];
assign g[4480] = a[10] & g[2432];
assign g[6527] = b[10] & g[2432];
assign g[4481] = a[10] & g[2433];
assign g[6528] = b[10] & g[2433];
assign g[4482] = a[10] & g[2434];
assign g[6529] = b[10] & g[2434];
assign g[4483] = a[10] & g[2435];
assign g[6530] = b[10] & g[2435];
assign g[4484] = a[10] & g[2436];
assign g[6531] = b[10] & g[2436];
assign g[4485] = a[10] & g[2437];
assign g[6532] = b[10] & g[2437];
assign g[4486] = a[10] & g[2438];
assign g[6533] = b[10] & g[2438];
assign g[4487] = a[10] & g[2439];
assign g[6534] = b[10] & g[2439];
assign g[4488] = a[10] & g[2440];
assign g[6535] = b[10] & g[2440];
assign g[4489] = a[10] & g[2441];
assign g[6536] = b[10] & g[2441];
assign g[4490] = a[10] & g[2442];
assign g[6537] = b[10] & g[2442];
assign g[4491] = a[10] & g[2443];
assign g[6538] = b[10] & g[2443];
assign g[4492] = a[10] & g[2444];
assign g[6539] = b[10] & g[2444];
assign g[4493] = a[10] & g[2445];
assign g[6540] = b[10] & g[2445];
assign g[4494] = a[10] & g[2446];
assign g[6541] = b[10] & g[2446];
assign g[4495] = a[10] & g[2447];
assign g[6542] = b[10] & g[2447];
assign g[4496] = a[10] & g[2448];
assign g[6543] = b[10] & g[2448];
assign g[4497] = a[10] & g[2449];
assign g[6544] = b[10] & g[2449];
assign g[4498] = a[10] & g[2450];
assign g[6545] = b[10] & g[2450];
assign g[4499] = a[10] & g[2451];
assign g[6546] = b[10] & g[2451];
assign g[4500] = a[10] & g[2452];
assign g[6547] = b[10] & g[2452];
assign g[4501] = a[10] & g[2453];
assign g[6548] = b[10] & g[2453];
assign g[4502] = a[10] & g[2454];
assign g[6549] = b[10] & g[2454];
assign g[4503] = a[10] & g[2455];
assign g[6550] = b[10] & g[2455];
assign g[4504] = a[10] & g[2456];
assign g[6551] = b[10] & g[2456];
assign g[4505] = a[10] & g[2457];
assign g[6552] = b[10] & g[2457];
assign g[4506] = a[10] & g[2458];
assign g[6553] = b[10] & g[2458];
assign g[4507] = a[10] & g[2459];
assign g[6554] = b[10] & g[2459];
assign g[4508] = a[10] & g[2460];
assign g[6555] = b[10] & g[2460];
assign g[4509] = a[10] & g[2461];
assign g[6556] = b[10] & g[2461];
assign g[4510] = a[10] & g[2462];
assign g[6557] = b[10] & g[2462];
assign g[4511] = a[10] & g[2463];
assign g[6558] = b[10] & g[2463];
assign g[4512] = a[10] & g[2464];
assign g[6559] = b[10] & g[2464];
assign g[4513] = a[10] & g[2465];
assign g[6560] = b[10] & g[2465];
assign g[4514] = a[10] & g[2466];
assign g[6561] = b[10] & g[2466];
assign g[4515] = a[10] & g[2467];
assign g[6562] = b[10] & g[2467];
assign g[4516] = a[10] & g[2468];
assign g[6563] = b[10] & g[2468];
assign g[4517] = a[10] & g[2469];
assign g[6564] = b[10] & g[2469];
assign g[4518] = a[10] & g[2470];
assign g[6565] = b[10] & g[2470];
assign g[4519] = a[10] & g[2471];
assign g[6566] = b[10] & g[2471];
assign g[4520] = a[10] & g[2472];
assign g[6567] = b[10] & g[2472];
assign g[4521] = a[10] & g[2473];
assign g[6568] = b[10] & g[2473];
assign g[4522] = a[10] & g[2474];
assign g[6569] = b[10] & g[2474];
assign g[4523] = a[10] & g[2475];
assign g[6570] = b[10] & g[2475];
assign g[4524] = a[10] & g[2476];
assign g[6571] = b[10] & g[2476];
assign g[4525] = a[10] & g[2477];
assign g[6572] = b[10] & g[2477];
assign g[4526] = a[10] & g[2478];
assign g[6573] = b[10] & g[2478];
assign g[4527] = a[10] & g[2479];
assign g[6574] = b[10] & g[2479];
assign g[4528] = a[10] & g[2480];
assign g[6575] = b[10] & g[2480];
assign g[4529] = a[10] & g[2481];
assign g[6576] = b[10] & g[2481];
assign g[4530] = a[10] & g[2482];
assign g[6577] = b[10] & g[2482];
assign g[4531] = a[10] & g[2483];
assign g[6578] = b[10] & g[2483];
assign g[4532] = a[10] & g[2484];
assign g[6579] = b[10] & g[2484];
assign g[4533] = a[10] & g[2485];
assign g[6580] = b[10] & g[2485];
assign g[4534] = a[10] & g[2486];
assign g[6581] = b[10] & g[2486];
assign g[4535] = a[10] & g[2487];
assign g[6582] = b[10] & g[2487];
assign g[4536] = a[10] & g[2488];
assign g[6583] = b[10] & g[2488];
assign g[4537] = a[10] & g[2489];
assign g[6584] = b[10] & g[2489];
assign g[4538] = a[10] & g[2490];
assign g[6585] = b[10] & g[2490];
assign g[4539] = a[10] & g[2491];
assign g[6586] = b[10] & g[2491];
assign g[4540] = a[10] & g[2492];
assign g[6587] = b[10] & g[2492];
assign g[4541] = a[10] & g[2493];
assign g[6588] = b[10] & g[2493];
assign g[4542] = a[10] & g[2494];
assign g[6589] = b[10] & g[2494];
assign g[4543] = a[10] & g[2495];
assign g[6590] = b[10] & g[2495];
assign g[4544] = a[10] & g[2496];
assign g[6591] = b[10] & g[2496];
assign g[4545] = a[10] & g[2497];
assign g[6592] = b[10] & g[2497];
assign g[4546] = a[10] & g[2498];
assign g[6593] = b[10] & g[2498];
assign g[4547] = a[10] & g[2499];
assign g[6594] = b[10] & g[2499];
assign g[4548] = a[10] & g[2500];
assign g[6595] = b[10] & g[2500];
assign g[4549] = a[10] & g[2501];
assign g[6596] = b[10] & g[2501];
assign g[4550] = a[10] & g[2502];
assign g[6597] = b[10] & g[2502];
assign g[4551] = a[10] & g[2503];
assign g[6598] = b[10] & g[2503];
assign g[4552] = a[10] & g[2504];
assign g[6599] = b[10] & g[2504];
assign g[4553] = a[10] & g[2505];
assign g[6600] = b[10] & g[2505];
assign g[4554] = a[10] & g[2506];
assign g[6601] = b[10] & g[2506];
assign g[4555] = a[10] & g[2507];
assign g[6602] = b[10] & g[2507];
assign g[4556] = a[10] & g[2508];
assign g[6603] = b[10] & g[2508];
assign g[4557] = a[10] & g[2509];
assign g[6604] = b[10] & g[2509];
assign g[4558] = a[10] & g[2510];
assign g[6605] = b[10] & g[2510];
assign g[4559] = a[10] & g[2511];
assign g[6606] = b[10] & g[2511];
assign g[4560] = a[10] & g[2512];
assign g[6607] = b[10] & g[2512];
assign g[4561] = a[10] & g[2513];
assign g[6608] = b[10] & g[2513];
assign g[4562] = a[10] & g[2514];
assign g[6609] = b[10] & g[2514];
assign g[4563] = a[10] & g[2515];
assign g[6610] = b[10] & g[2515];
assign g[4564] = a[10] & g[2516];
assign g[6611] = b[10] & g[2516];
assign g[4565] = a[10] & g[2517];
assign g[6612] = b[10] & g[2517];
assign g[4566] = a[10] & g[2518];
assign g[6613] = b[10] & g[2518];
assign g[4567] = a[10] & g[2519];
assign g[6614] = b[10] & g[2519];
assign g[4568] = a[10] & g[2520];
assign g[6615] = b[10] & g[2520];
assign g[4569] = a[10] & g[2521];
assign g[6616] = b[10] & g[2521];
assign g[4570] = a[10] & g[2522];
assign g[6617] = b[10] & g[2522];
assign g[4571] = a[10] & g[2523];
assign g[6618] = b[10] & g[2523];
assign g[4572] = a[10] & g[2524];
assign g[6619] = b[10] & g[2524];
assign g[4573] = a[10] & g[2525];
assign g[6620] = b[10] & g[2525];
assign g[4574] = a[10] & g[2526];
assign g[6621] = b[10] & g[2526];
assign g[4575] = a[10] & g[2527];
assign g[6622] = b[10] & g[2527];
assign g[4576] = a[10] & g[2528];
assign g[6623] = b[10] & g[2528];
assign g[4577] = a[10] & g[2529];
assign g[6624] = b[10] & g[2529];
assign g[4578] = a[10] & g[2530];
assign g[6625] = b[10] & g[2530];
assign g[4579] = a[10] & g[2531];
assign g[6626] = b[10] & g[2531];
assign g[4580] = a[10] & g[2532];
assign g[6627] = b[10] & g[2532];
assign g[4581] = a[10] & g[2533];
assign g[6628] = b[10] & g[2533];
assign g[4582] = a[10] & g[2534];
assign g[6629] = b[10] & g[2534];
assign g[4583] = a[10] & g[2535];
assign g[6630] = b[10] & g[2535];
assign g[4584] = a[10] & g[2536];
assign g[6631] = b[10] & g[2536];
assign g[4585] = a[10] & g[2537];
assign g[6632] = b[10] & g[2537];
assign g[4586] = a[10] & g[2538];
assign g[6633] = b[10] & g[2538];
assign g[4587] = a[10] & g[2539];
assign g[6634] = b[10] & g[2539];
assign g[4588] = a[10] & g[2540];
assign g[6635] = b[10] & g[2540];
assign g[4589] = a[10] & g[2541];
assign g[6636] = b[10] & g[2541];
assign g[4590] = a[10] & g[2542];
assign g[6637] = b[10] & g[2542];
assign g[4591] = a[10] & g[2543];
assign g[6638] = b[10] & g[2543];
assign g[4592] = a[10] & g[2544];
assign g[6639] = b[10] & g[2544];
assign g[4593] = a[10] & g[2545];
assign g[6640] = b[10] & g[2545];
assign g[4594] = a[10] & g[2546];
assign g[6641] = b[10] & g[2546];
assign g[4595] = a[10] & g[2547];
assign g[6642] = b[10] & g[2547];
assign g[4596] = a[10] & g[2548];
assign g[6643] = b[10] & g[2548];
assign g[4597] = a[10] & g[2549];
assign g[6644] = b[10] & g[2549];
assign g[4598] = a[10] & g[2550];
assign g[6645] = b[10] & g[2550];
assign g[4599] = a[10] & g[2551];
assign g[6646] = b[10] & g[2551];
assign g[4600] = a[10] & g[2552];
assign g[6647] = b[10] & g[2552];
assign g[4601] = a[10] & g[2553];
assign g[6648] = b[10] & g[2553];
assign g[4602] = a[10] & g[2554];
assign g[6649] = b[10] & g[2554];
assign g[4603] = a[10] & g[2555];
assign g[6650] = b[10] & g[2555];
assign g[4604] = a[10] & g[2556];
assign g[6651] = b[10] & g[2556];
assign g[4605] = a[10] & g[2557];
assign g[6652] = b[10] & g[2557];
assign g[4606] = a[10] & g[2558];
assign g[6653] = b[10] & g[2558];
assign g[4607] = a[10] & g[2559];
assign g[6654] = b[10] & g[2559];
assign g[4608] = a[10] & g[2560];
assign g[6655] = b[10] & g[2560];
assign g[4609] = a[10] & g[2561];
assign g[6656] = b[10] & g[2561];
assign g[4610] = a[10] & g[2562];
assign g[6657] = b[10] & g[2562];
assign g[4611] = a[10] & g[2563];
assign g[6658] = b[10] & g[2563];
assign g[4612] = a[10] & g[2564];
assign g[6659] = b[10] & g[2564];
assign g[4613] = a[10] & g[2565];
assign g[6660] = b[10] & g[2565];
assign g[4614] = a[10] & g[2566];
assign g[6661] = b[10] & g[2566];
assign g[4615] = a[10] & g[2567];
assign g[6662] = b[10] & g[2567];
assign g[4616] = a[10] & g[2568];
assign g[6663] = b[10] & g[2568];
assign g[4617] = a[10] & g[2569];
assign g[6664] = b[10] & g[2569];
assign g[4618] = a[10] & g[2570];
assign g[6665] = b[10] & g[2570];
assign g[4619] = a[10] & g[2571];
assign g[6666] = b[10] & g[2571];
assign g[4620] = a[10] & g[2572];
assign g[6667] = b[10] & g[2572];
assign g[4621] = a[10] & g[2573];
assign g[6668] = b[10] & g[2573];
assign g[4622] = a[10] & g[2574];
assign g[6669] = b[10] & g[2574];
assign g[4623] = a[10] & g[2575];
assign g[6670] = b[10] & g[2575];
assign g[4624] = a[10] & g[2576];
assign g[6671] = b[10] & g[2576];
assign g[4625] = a[10] & g[2577];
assign g[6672] = b[10] & g[2577];
assign g[4626] = a[10] & g[2578];
assign g[6673] = b[10] & g[2578];
assign g[4627] = a[10] & g[2579];
assign g[6674] = b[10] & g[2579];
assign g[4628] = a[10] & g[2580];
assign g[6675] = b[10] & g[2580];
assign g[4629] = a[10] & g[2581];
assign g[6676] = b[10] & g[2581];
assign g[4630] = a[10] & g[2582];
assign g[6677] = b[10] & g[2582];
assign g[4631] = a[10] & g[2583];
assign g[6678] = b[10] & g[2583];
assign g[4632] = a[10] & g[2584];
assign g[6679] = b[10] & g[2584];
assign g[4633] = a[10] & g[2585];
assign g[6680] = b[10] & g[2585];
assign g[4634] = a[10] & g[2586];
assign g[6681] = b[10] & g[2586];
assign g[4635] = a[10] & g[2587];
assign g[6682] = b[10] & g[2587];
assign g[4636] = a[10] & g[2588];
assign g[6683] = b[10] & g[2588];
assign g[4637] = a[10] & g[2589];
assign g[6684] = b[10] & g[2589];
assign g[4638] = a[10] & g[2590];
assign g[6685] = b[10] & g[2590];
assign g[4639] = a[10] & g[2591];
assign g[6686] = b[10] & g[2591];
assign g[4640] = a[10] & g[2592];
assign g[6687] = b[10] & g[2592];
assign g[4641] = a[10] & g[2593];
assign g[6688] = b[10] & g[2593];
assign g[4642] = a[10] & g[2594];
assign g[6689] = b[10] & g[2594];
assign g[4643] = a[10] & g[2595];
assign g[6690] = b[10] & g[2595];
assign g[4644] = a[10] & g[2596];
assign g[6691] = b[10] & g[2596];
assign g[4645] = a[10] & g[2597];
assign g[6692] = b[10] & g[2597];
assign g[4646] = a[10] & g[2598];
assign g[6693] = b[10] & g[2598];
assign g[4647] = a[10] & g[2599];
assign g[6694] = b[10] & g[2599];
assign g[4648] = a[10] & g[2600];
assign g[6695] = b[10] & g[2600];
assign g[4649] = a[10] & g[2601];
assign g[6696] = b[10] & g[2601];
assign g[4650] = a[10] & g[2602];
assign g[6697] = b[10] & g[2602];
assign g[4651] = a[10] & g[2603];
assign g[6698] = b[10] & g[2603];
assign g[4652] = a[10] & g[2604];
assign g[6699] = b[10] & g[2604];
assign g[4653] = a[10] & g[2605];
assign g[6700] = b[10] & g[2605];
assign g[4654] = a[10] & g[2606];
assign g[6701] = b[10] & g[2606];
assign g[4655] = a[10] & g[2607];
assign g[6702] = b[10] & g[2607];
assign g[4656] = a[10] & g[2608];
assign g[6703] = b[10] & g[2608];
assign g[4657] = a[10] & g[2609];
assign g[6704] = b[10] & g[2609];
assign g[4658] = a[10] & g[2610];
assign g[6705] = b[10] & g[2610];
assign g[4659] = a[10] & g[2611];
assign g[6706] = b[10] & g[2611];
assign g[4660] = a[10] & g[2612];
assign g[6707] = b[10] & g[2612];
assign g[4661] = a[10] & g[2613];
assign g[6708] = b[10] & g[2613];
assign g[4662] = a[10] & g[2614];
assign g[6709] = b[10] & g[2614];
assign g[4663] = a[10] & g[2615];
assign g[6710] = b[10] & g[2615];
assign g[4664] = a[10] & g[2616];
assign g[6711] = b[10] & g[2616];
assign g[4665] = a[10] & g[2617];
assign g[6712] = b[10] & g[2617];
assign g[4666] = a[10] & g[2618];
assign g[6713] = b[10] & g[2618];
assign g[4667] = a[10] & g[2619];
assign g[6714] = b[10] & g[2619];
assign g[4668] = a[10] & g[2620];
assign g[6715] = b[10] & g[2620];
assign g[4669] = a[10] & g[2621];
assign g[6716] = b[10] & g[2621];
assign g[4670] = a[10] & g[2622];
assign g[6717] = b[10] & g[2622];
assign g[4671] = a[10] & g[2623];
assign g[6718] = b[10] & g[2623];
assign g[4672] = a[10] & g[2624];
assign g[6719] = b[10] & g[2624];
assign g[4673] = a[10] & g[2625];
assign g[6720] = b[10] & g[2625];
assign g[4674] = a[10] & g[2626];
assign g[6721] = b[10] & g[2626];
assign g[4675] = a[10] & g[2627];
assign g[6722] = b[10] & g[2627];
assign g[4676] = a[10] & g[2628];
assign g[6723] = b[10] & g[2628];
assign g[4677] = a[10] & g[2629];
assign g[6724] = b[10] & g[2629];
assign g[4678] = a[10] & g[2630];
assign g[6725] = b[10] & g[2630];
assign g[4679] = a[10] & g[2631];
assign g[6726] = b[10] & g[2631];
assign g[4680] = a[10] & g[2632];
assign g[6727] = b[10] & g[2632];
assign g[4681] = a[10] & g[2633];
assign g[6728] = b[10] & g[2633];
assign g[4682] = a[10] & g[2634];
assign g[6729] = b[10] & g[2634];
assign g[4683] = a[10] & g[2635];
assign g[6730] = b[10] & g[2635];
assign g[4684] = a[10] & g[2636];
assign g[6731] = b[10] & g[2636];
assign g[4685] = a[10] & g[2637];
assign g[6732] = b[10] & g[2637];
assign g[4686] = a[10] & g[2638];
assign g[6733] = b[10] & g[2638];
assign g[4687] = a[10] & g[2639];
assign g[6734] = b[10] & g[2639];
assign g[4688] = a[10] & g[2640];
assign g[6735] = b[10] & g[2640];
assign g[4689] = a[10] & g[2641];
assign g[6736] = b[10] & g[2641];
assign g[4690] = a[10] & g[2642];
assign g[6737] = b[10] & g[2642];
assign g[4691] = a[10] & g[2643];
assign g[6738] = b[10] & g[2643];
assign g[4692] = a[10] & g[2644];
assign g[6739] = b[10] & g[2644];
assign g[4693] = a[10] & g[2645];
assign g[6740] = b[10] & g[2645];
assign g[4694] = a[10] & g[2646];
assign g[6741] = b[10] & g[2646];
assign g[4695] = a[10] & g[2647];
assign g[6742] = b[10] & g[2647];
assign g[4696] = a[10] & g[2648];
assign g[6743] = b[10] & g[2648];
assign g[4697] = a[10] & g[2649];
assign g[6744] = b[10] & g[2649];
assign g[4698] = a[10] & g[2650];
assign g[6745] = b[10] & g[2650];
assign g[4699] = a[10] & g[2651];
assign g[6746] = b[10] & g[2651];
assign g[4700] = a[10] & g[2652];
assign g[6747] = b[10] & g[2652];
assign g[4701] = a[10] & g[2653];
assign g[6748] = b[10] & g[2653];
assign g[4702] = a[10] & g[2654];
assign g[6749] = b[10] & g[2654];
assign g[4703] = a[10] & g[2655];
assign g[6750] = b[10] & g[2655];
assign g[4704] = a[10] & g[2656];
assign g[6751] = b[10] & g[2656];
assign g[4705] = a[10] & g[2657];
assign g[6752] = b[10] & g[2657];
assign g[4706] = a[10] & g[2658];
assign g[6753] = b[10] & g[2658];
assign g[4707] = a[10] & g[2659];
assign g[6754] = b[10] & g[2659];
assign g[4708] = a[10] & g[2660];
assign g[6755] = b[10] & g[2660];
assign g[4709] = a[10] & g[2661];
assign g[6756] = b[10] & g[2661];
assign g[4710] = a[10] & g[2662];
assign g[6757] = b[10] & g[2662];
assign g[4711] = a[10] & g[2663];
assign g[6758] = b[10] & g[2663];
assign g[4712] = a[10] & g[2664];
assign g[6759] = b[10] & g[2664];
assign g[4713] = a[10] & g[2665];
assign g[6760] = b[10] & g[2665];
assign g[4714] = a[10] & g[2666];
assign g[6761] = b[10] & g[2666];
assign g[4715] = a[10] & g[2667];
assign g[6762] = b[10] & g[2667];
assign g[4716] = a[10] & g[2668];
assign g[6763] = b[10] & g[2668];
assign g[4717] = a[10] & g[2669];
assign g[6764] = b[10] & g[2669];
assign g[4718] = a[10] & g[2670];
assign g[6765] = b[10] & g[2670];
assign g[4719] = a[10] & g[2671];
assign g[6766] = b[10] & g[2671];
assign g[4720] = a[10] & g[2672];
assign g[6767] = b[10] & g[2672];
assign g[4721] = a[10] & g[2673];
assign g[6768] = b[10] & g[2673];
assign g[4722] = a[10] & g[2674];
assign g[6769] = b[10] & g[2674];
assign g[4723] = a[10] & g[2675];
assign g[6770] = b[10] & g[2675];
assign g[4724] = a[10] & g[2676];
assign g[6771] = b[10] & g[2676];
assign g[4725] = a[10] & g[2677];
assign g[6772] = b[10] & g[2677];
assign g[4726] = a[10] & g[2678];
assign g[6773] = b[10] & g[2678];
assign g[4727] = a[10] & g[2679];
assign g[6774] = b[10] & g[2679];
assign g[4728] = a[10] & g[2680];
assign g[6775] = b[10] & g[2680];
assign g[4729] = a[10] & g[2681];
assign g[6776] = b[10] & g[2681];
assign g[4730] = a[10] & g[2682];
assign g[6777] = b[10] & g[2682];
assign g[4731] = a[10] & g[2683];
assign g[6778] = b[10] & g[2683];
assign g[4732] = a[10] & g[2684];
assign g[6779] = b[10] & g[2684];
assign g[4733] = a[10] & g[2685];
assign g[6780] = b[10] & g[2685];
assign g[4734] = a[10] & g[2686];
assign g[6781] = b[10] & g[2686];
assign g[4735] = a[10] & g[2687];
assign g[6782] = b[10] & g[2687];
assign g[4736] = a[10] & g[2688];
assign g[6783] = b[10] & g[2688];
assign g[4737] = a[10] & g[2689];
assign g[6784] = b[10] & g[2689];
assign g[4738] = a[10] & g[2690];
assign g[6785] = b[10] & g[2690];
assign g[4739] = a[10] & g[2691];
assign g[6786] = b[10] & g[2691];
assign g[4740] = a[10] & g[2692];
assign g[6787] = b[10] & g[2692];
assign g[4741] = a[10] & g[2693];
assign g[6788] = b[10] & g[2693];
assign g[4742] = a[10] & g[2694];
assign g[6789] = b[10] & g[2694];
assign g[4743] = a[10] & g[2695];
assign g[6790] = b[10] & g[2695];
assign g[4744] = a[10] & g[2696];
assign g[6791] = b[10] & g[2696];
assign g[4745] = a[10] & g[2697];
assign g[6792] = b[10] & g[2697];
assign g[4746] = a[10] & g[2698];
assign g[6793] = b[10] & g[2698];
assign g[4747] = a[10] & g[2699];
assign g[6794] = b[10] & g[2699];
assign g[4748] = a[10] & g[2700];
assign g[6795] = b[10] & g[2700];
assign g[4749] = a[10] & g[2701];
assign g[6796] = b[10] & g[2701];
assign g[4750] = a[10] & g[2702];
assign g[6797] = b[10] & g[2702];
assign g[4751] = a[10] & g[2703];
assign g[6798] = b[10] & g[2703];
assign g[4752] = a[10] & g[2704];
assign g[6799] = b[10] & g[2704];
assign g[4753] = a[10] & g[2705];
assign g[6800] = b[10] & g[2705];
assign g[4754] = a[10] & g[2706];
assign g[6801] = b[10] & g[2706];
assign g[4755] = a[10] & g[2707];
assign g[6802] = b[10] & g[2707];
assign g[4756] = a[10] & g[2708];
assign g[6803] = b[10] & g[2708];
assign g[4757] = a[10] & g[2709];
assign g[6804] = b[10] & g[2709];
assign g[4758] = a[10] & g[2710];
assign g[6805] = b[10] & g[2710];
assign g[4759] = a[10] & g[2711];
assign g[6806] = b[10] & g[2711];
assign g[4760] = a[10] & g[2712];
assign g[6807] = b[10] & g[2712];
assign g[4761] = a[10] & g[2713];
assign g[6808] = b[10] & g[2713];
assign g[4762] = a[10] & g[2714];
assign g[6809] = b[10] & g[2714];
assign g[4763] = a[10] & g[2715];
assign g[6810] = b[10] & g[2715];
assign g[4764] = a[10] & g[2716];
assign g[6811] = b[10] & g[2716];
assign g[4765] = a[10] & g[2717];
assign g[6812] = b[10] & g[2717];
assign g[4766] = a[10] & g[2718];
assign g[6813] = b[10] & g[2718];
assign g[4767] = a[10] & g[2719];
assign g[6814] = b[10] & g[2719];
assign g[4768] = a[10] & g[2720];
assign g[6815] = b[10] & g[2720];
assign g[4769] = a[10] & g[2721];
assign g[6816] = b[10] & g[2721];
assign g[4770] = a[10] & g[2722];
assign g[6817] = b[10] & g[2722];
assign g[4771] = a[10] & g[2723];
assign g[6818] = b[10] & g[2723];
assign g[4772] = a[10] & g[2724];
assign g[6819] = b[10] & g[2724];
assign g[4773] = a[10] & g[2725];
assign g[6820] = b[10] & g[2725];
assign g[4774] = a[10] & g[2726];
assign g[6821] = b[10] & g[2726];
assign g[4775] = a[10] & g[2727];
assign g[6822] = b[10] & g[2727];
assign g[4776] = a[10] & g[2728];
assign g[6823] = b[10] & g[2728];
assign g[4777] = a[10] & g[2729];
assign g[6824] = b[10] & g[2729];
assign g[4778] = a[10] & g[2730];
assign g[6825] = b[10] & g[2730];
assign g[4779] = a[10] & g[2731];
assign g[6826] = b[10] & g[2731];
assign g[4780] = a[10] & g[2732];
assign g[6827] = b[10] & g[2732];
assign g[4781] = a[10] & g[2733];
assign g[6828] = b[10] & g[2733];
assign g[4782] = a[10] & g[2734];
assign g[6829] = b[10] & g[2734];
assign g[4783] = a[10] & g[2735];
assign g[6830] = b[10] & g[2735];
assign g[4784] = a[10] & g[2736];
assign g[6831] = b[10] & g[2736];
assign g[4785] = a[10] & g[2737];
assign g[6832] = b[10] & g[2737];
assign g[4786] = a[10] & g[2738];
assign g[6833] = b[10] & g[2738];
assign g[4787] = a[10] & g[2739];
assign g[6834] = b[10] & g[2739];
assign g[4788] = a[10] & g[2740];
assign g[6835] = b[10] & g[2740];
assign g[4789] = a[10] & g[2741];
assign g[6836] = b[10] & g[2741];
assign g[4790] = a[10] & g[2742];
assign g[6837] = b[10] & g[2742];
assign g[4791] = a[10] & g[2743];
assign g[6838] = b[10] & g[2743];
assign g[4792] = a[10] & g[2744];
assign g[6839] = b[10] & g[2744];
assign g[4793] = a[10] & g[2745];
assign g[6840] = b[10] & g[2745];
assign g[4794] = a[10] & g[2746];
assign g[6841] = b[10] & g[2746];
assign g[4795] = a[10] & g[2747];
assign g[6842] = b[10] & g[2747];
assign g[4796] = a[10] & g[2748];
assign g[6843] = b[10] & g[2748];
assign g[4797] = a[10] & g[2749];
assign g[6844] = b[10] & g[2749];
assign g[4798] = a[10] & g[2750];
assign g[6845] = b[10] & g[2750];
assign g[4799] = a[10] & g[2751];
assign g[6846] = b[10] & g[2751];
assign g[4800] = a[10] & g[2752];
assign g[6847] = b[10] & g[2752];
assign g[4801] = a[10] & g[2753];
assign g[6848] = b[10] & g[2753];
assign g[4802] = a[10] & g[2754];
assign g[6849] = b[10] & g[2754];
assign g[4803] = a[10] & g[2755];
assign g[6850] = b[10] & g[2755];
assign g[4804] = a[10] & g[2756];
assign g[6851] = b[10] & g[2756];
assign g[4805] = a[10] & g[2757];
assign g[6852] = b[10] & g[2757];
assign g[4806] = a[10] & g[2758];
assign g[6853] = b[10] & g[2758];
assign g[4807] = a[10] & g[2759];
assign g[6854] = b[10] & g[2759];
assign g[4808] = a[10] & g[2760];
assign g[6855] = b[10] & g[2760];
assign g[4809] = a[10] & g[2761];
assign g[6856] = b[10] & g[2761];
assign g[4810] = a[10] & g[2762];
assign g[6857] = b[10] & g[2762];
assign g[4811] = a[10] & g[2763];
assign g[6858] = b[10] & g[2763];
assign g[4812] = a[10] & g[2764];
assign g[6859] = b[10] & g[2764];
assign g[4813] = a[10] & g[2765];
assign g[6860] = b[10] & g[2765];
assign g[4814] = a[10] & g[2766];
assign g[6861] = b[10] & g[2766];
assign g[4815] = a[10] & g[2767];
assign g[6862] = b[10] & g[2767];
assign g[4816] = a[10] & g[2768];
assign g[6863] = b[10] & g[2768];
assign g[4817] = a[10] & g[2769];
assign g[6864] = b[10] & g[2769];
assign g[4818] = a[10] & g[2770];
assign g[6865] = b[10] & g[2770];
assign g[4819] = a[10] & g[2771];
assign g[6866] = b[10] & g[2771];
assign g[4820] = a[10] & g[2772];
assign g[6867] = b[10] & g[2772];
assign g[4821] = a[10] & g[2773];
assign g[6868] = b[10] & g[2773];
assign g[4822] = a[10] & g[2774];
assign g[6869] = b[10] & g[2774];
assign g[4823] = a[10] & g[2775];
assign g[6870] = b[10] & g[2775];
assign g[4824] = a[10] & g[2776];
assign g[6871] = b[10] & g[2776];
assign g[4825] = a[10] & g[2777];
assign g[6872] = b[10] & g[2777];
assign g[4826] = a[10] & g[2778];
assign g[6873] = b[10] & g[2778];
assign g[4827] = a[10] & g[2779];
assign g[6874] = b[10] & g[2779];
assign g[4828] = a[10] & g[2780];
assign g[6875] = b[10] & g[2780];
assign g[4829] = a[10] & g[2781];
assign g[6876] = b[10] & g[2781];
assign g[4830] = a[10] & g[2782];
assign g[6877] = b[10] & g[2782];
assign g[4831] = a[10] & g[2783];
assign g[6878] = b[10] & g[2783];
assign g[4832] = a[10] & g[2784];
assign g[6879] = b[10] & g[2784];
assign g[4833] = a[10] & g[2785];
assign g[6880] = b[10] & g[2785];
assign g[4834] = a[10] & g[2786];
assign g[6881] = b[10] & g[2786];
assign g[4835] = a[10] & g[2787];
assign g[6882] = b[10] & g[2787];
assign g[4836] = a[10] & g[2788];
assign g[6883] = b[10] & g[2788];
assign g[4837] = a[10] & g[2789];
assign g[6884] = b[10] & g[2789];
assign g[4838] = a[10] & g[2790];
assign g[6885] = b[10] & g[2790];
assign g[4839] = a[10] & g[2791];
assign g[6886] = b[10] & g[2791];
assign g[4840] = a[10] & g[2792];
assign g[6887] = b[10] & g[2792];
assign g[4841] = a[10] & g[2793];
assign g[6888] = b[10] & g[2793];
assign g[4842] = a[10] & g[2794];
assign g[6889] = b[10] & g[2794];
assign g[4843] = a[10] & g[2795];
assign g[6890] = b[10] & g[2795];
assign g[4844] = a[10] & g[2796];
assign g[6891] = b[10] & g[2796];
assign g[4845] = a[10] & g[2797];
assign g[6892] = b[10] & g[2797];
assign g[4846] = a[10] & g[2798];
assign g[6893] = b[10] & g[2798];
assign g[4847] = a[10] & g[2799];
assign g[6894] = b[10] & g[2799];
assign g[4848] = a[10] & g[2800];
assign g[6895] = b[10] & g[2800];
assign g[4849] = a[10] & g[2801];
assign g[6896] = b[10] & g[2801];
assign g[4850] = a[10] & g[2802];
assign g[6897] = b[10] & g[2802];
assign g[4851] = a[10] & g[2803];
assign g[6898] = b[10] & g[2803];
assign g[4852] = a[10] & g[2804];
assign g[6899] = b[10] & g[2804];
assign g[4853] = a[10] & g[2805];
assign g[6900] = b[10] & g[2805];
assign g[4854] = a[10] & g[2806];
assign g[6901] = b[10] & g[2806];
assign g[4855] = a[10] & g[2807];
assign g[6902] = b[10] & g[2807];
assign g[4856] = a[10] & g[2808];
assign g[6903] = b[10] & g[2808];
assign g[4857] = a[10] & g[2809];
assign g[6904] = b[10] & g[2809];
assign g[4858] = a[10] & g[2810];
assign g[6905] = b[10] & g[2810];
assign g[4859] = a[10] & g[2811];
assign g[6906] = b[10] & g[2811];
assign g[4860] = a[10] & g[2812];
assign g[6907] = b[10] & g[2812];
assign g[4861] = a[10] & g[2813];
assign g[6908] = b[10] & g[2813];
assign g[4862] = a[10] & g[2814];
assign g[6909] = b[10] & g[2814];
assign g[4863] = a[10] & g[2815];
assign g[6910] = b[10] & g[2815];
assign g[4864] = a[10] & g[2816];
assign g[6911] = b[10] & g[2816];
assign g[4865] = a[10] & g[2817];
assign g[6912] = b[10] & g[2817];
assign g[4866] = a[10] & g[2818];
assign g[6913] = b[10] & g[2818];
assign g[4867] = a[10] & g[2819];
assign g[6914] = b[10] & g[2819];
assign g[4868] = a[10] & g[2820];
assign g[6915] = b[10] & g[2820];
assign g[4869] = a[10] & g[2821];
assign g[6916] = b[10] & g[2821];
assign g[4870] = a[10] & g[2822];
assign g[6917] = b[10] & g[2822];
assign g[4871] = a[10] & g[2823];
assign g[6918] = b[10] & g[2823];
assign g[4872] = a[10] & g[2824];
assign g[6919] = b[10] & g[2824];
assign g[4873] = a[10] & g[2825];
assign g[6920] = b[10] & g[2825];
assign g[4874] = a[10] & g[2826];
assign g[6921] = b[10] & g[2826];
assign g[4875] = a[10] & g[2827];
assign g[6922] = b[10] & g[2827];
assign g[4876] = a[10] & g[2828];
assign g[6923] = b[10] & g[2828];
assign g[4877] = a[10] & g[2829];
assign g[6924] = b[10] & g[2829];
assign g[4878] = a[10] & g[2830];
assign g[6925] = b[10] & g[2830];
assign g[4879] = a[10] & g[2831];
assign g[6926] = b[10] & g[2831];
assign g[4880] = a[10] & g[2832];
assign g[6927] = b[10] & g[2832];
assign g[4881] = a[10] & g[2833];
assign g[6928] = b[10] & g[2833];
assign g[4882] = a[10] & g[2834];
assign g[6929] = b[10] & g[2834];
assign g[4883] = a[10] & g[2835];
assign g[6930] = b[10] & g[2835];
assign g[4884] = a[10] & g[2836];
assign g[6931] = b[10] & g[2836];
assign g[4885] = a[10] & g[2837];
assign g[6932] = b[10] & g[2837];
assign g[4886] = a[10] & g[2838];
assign g[6933] = b[10] & g[2838];
assign g[4887] = a[10] & g[2839];
assign g[6934] = b[10] & g[2839];
assign g[4888] = a[10] & g[2840];
assign g[6935] = b[10] & g[2840];
assign g[4889] = a[10] & g[2841];
assign g[6936] = b[10] & g[2841];
assign g[4890] = a[10] & g[2842];
assign g[6937] = b[10] & g[2842];
assign g[4891] = a[10] & g[2843];
assign g[6938] = b[10] & g[2843];
assign g[4892] = a[10] & g[2844];
assign g[6939] = b[10] & g[2844];
assign g[4893] = a[10] & g[2845];
assign g[6940] = b[10] & g[2845];
assign g[4894] = a[10] & g[2846];
assign g[6941] = b[10] & g[2846];
assign g[4895] = a[10] & g[2847];
assign g[6942] = b[10] & g[2847];
assign g[4896] = a[10] & g[2848];
assign g[6943] = b[10] & g[2848];
assign g[4897] = a[10] & g[2849];
assign g[6944] = b[10] & g[2849];
assign g[4898] = a[10] & g[2850];
assign g[6945] = b[10] & g[2850];
assign g[4899] = a[10] & g[2851];
assign g[6946] = b[10] & g[2851];
assign g[4900] = a[10] & g[2852];
assign g[6947] = b[10] & g[2852];
assign g[4901] = a[10] & g[2853];
assign g[6948] = b[10] & g[2853];
assign g[4902] = a[10] & g[2854];
assign g[6949] = b[10] & g[2854];
assign g[4903] = a[10] & g[2855];
assign g[6950] = b[10] & g[2855];
assign g[4904] = a[10] & g[2856];
assign g[6951] = b[10] & g[2856];
assign g[4905] = a[10] & g[2857];
assign g[6952] = b[10] & g[2857];
assign g[4906] = a[10] & g[2858];
assign g[6953] = b[10] & g[2858];
assign g[4907] = a[10] & g[2859];
assign g[6954] = b[10] & g[2859];
assign g[4908] = a[10] & g[2860];
assign g[6955] = b[10] & g[2860];
assign g[4909] = a[10] & g[2861];
assign g[6956] = b[10] & g[2861];
assign g[4910] = a[10] & g[2862];
assign g[6957] = b[10] & g[2862];
assign g[4911] = a[10] & g[2863];
assign g[6958] = b[10] & g[2863];
assign g[4912] = a[10] & g[2864];
assign g[6959] = b[10] & g[2864];
assign g[4913] = a[10] & g[2865];
assign g[6960] = b[10] & g[2865];
assign g[4914] = a[10] & g[2866];
assign g[6961] = b[10] & g[2866];
assign g[4915] = a[10] & g[2867];
assign g[6962] = b[10] & g[2867];
assign g[4916] = a[10] & g[2868];
assign g[6963] = b[10] & g[2868];
assign g[4917] = a[10] & g[2869];
assign g[6964] = b[10] & g[2869];
assign g[4918] = a[10] & g[2870];
assign g[6965] = b[10] & g[2870];
assign g[4919] = a[10] & g[2871];
assign g[6966] = b[10] & g[2871];
assign g[4920] = a[10] & g[2872];
assign g[6967] = b[10] & g[2872];
assign g[4921] = a[10] & g[2873];
assign g[6968] = b[10] & g[2873];
assign g[4922] = a[10] & g[2874];
assign g[6969] = b[10] & g[2874];
assign g[4923] = a[10] & g[2875];
assign g[6970] = b[10] & g[2875];
assign g[4924] = a[10] & g[2876];
assign g[6971] = b[10] & g[2876];
assign g[4925] = a[10] & g[2877];
assign g[6972] = b[10] & g[2877];
assign g[4926] = a[10] & g[2878];
assign g[6973] = b[10] & g[2878];
assign g[4927] = a[10] & g[2879];
assign g[6974] = b[10] & g[2879];
assign g[4928] = a[10] & g[2880];
assign g[6975] = b[10] & g[2880];
assign g[4929] = a[10] & g[2881];
assign g[6976] = b[10] & g[2881];
assign g[4930] = a[10] & g[2882];
assign g[6977] = b[10] & g[2882];
assign g[4931] = a[10] & g[2883];
assign g[6978] = b[10] & g[2883];
assign g[4932] = a[10] & g[2884];
assign g[6979] = b[10] & g[2884];
assign g[4933] = a[10] & g[2885];
assign g[6980] = b[10] & g[2885];
assign g[4934] = a[10] & g[2886];
assign g[6981] = b[10] & g[2886];
assign g[4935] = a[10] & g[2887];
assign g[6982] = b[10] & g[2887];
assign g[4936] = a[10] & g[2888];
assign g[6983] = b[10] & g[2888];
assign g[4937] = a[10] & g[2889];
assign g[6984] = b[10] & g[2889];
assign g[4938] = a[10] & g[2890];
assign g[6985] = b[10] & g[2890];
assign g[4939] = a[10] & g[2891];
assign g[6986] = b[10] & g[2891];
assign g[4940] = a[10] & g[2892];
assign g[6987] = b[10] & g[2892];
assign g[4941] = a[10] & g[2893];
assign g[6988] = b[10] & g[2893];
assign g[4942] = a[10] & g[2894];
assign g[6989] = b[10] & g[2894];
assign g[4943] = a[10] & g[2895];
assign g[6990] = b[10] & g[2895];
assign g[4944] = a[10] & g[2896];
assign g[6991] = b[10] & g[2896];
assign g[4945] = a[10] & g[2897];
assign g[6992] = b[10] & g[2897];
assign g[4946] = a[10] & g[2898];
assign g[6993] = b[10] & g[2898];
assign g[4947] = a[10] & g[2899];
assign g[6994] = b[10] & g[2899];
assign g[4948] = a[10] & g[2900];
assign g[6995] = b[10] & g[2900];
assign g[4949] = a[10] & g[2901];
assign g[6996] = b[10] & g[2901];
assign g[4950] = a[10] & g[2902];
assign g[6997] = b[10] & g[2902];
assign g[4951] = a[10] & g[2903];
assign g[6998] = b[10] & g[2903];
assign g[4952] = a[10] & g[2904];
assign g[6999] = b[10] & g[2904];
assign g[4953] = a[10] & g[2905];
assign g[7000] = b[10] & g[2905];
assign g[4954] = a[10] & g[2906];
assign g[7001] = b[10] & g[2906];
assign g[4955] = a[10] & g[2907];
assign g[7002] = b[10] & g[2907];
assign g[4956] = a[10] & g[2908];
assign g[7003] = b[10] & g[2908];
assign g[4957] = a[10] & g[2909];
assign g[7004] = b[10] & g[2909];
assign g[4958] = a[10] & g[2910];
assign g[7005] = b[10] & g[2910];
assign g[4959] = a[10] & g[2911];
assign g[7006] = b[10] & g[2911];
assign g[4960] = a[10] & g[2912];
assign g[7007] = b[10] & g[2912];
assign g[4961] = a[10] & g[2913];
assign g[7008] = b[10] & g[2913];
assign g[4962] = a[10] & g[2914];
assign g[7009] = b[10] & g[2914];
assign g[4963] = a[10] & g[2915];
assign g[7010] = b[10] & g[2915];
assign g[4964] = a[10] & g[2916];
assign g[7011] = b[10] & g[2916];
assign g[4965] = a[10] & g[2917];
assign g[7012] = b[10] & g[2917];
assign g[4966] = a[10] & g[2918];
assign g[7013] = b[10] & g[2918];
assign g[4967] = a[10] & g[2919];
assign g[7014] = b[10] & g[2919];
assign g[4968] = a[10] & g[2920];
assign g[7015] = b[10] & g[2920];
assign g[4969] = a[10] & g[2921];
assign g[7016] = b[10] & g[2921];
assign g[4970] = a[10] & g[2922];
assign g[7017] = b[10] & g[2922];
assign g[4971] = a[10] & g[2923];
assign g[7018] = b[10] & g[2923];
assign g[4972] = a[10] & g[2924];
assign g[7019] = b[10] & g[2924];
assign g[4973] = a[10] & g[2925];
assign g[7020] = b[10] & g[2925];
assign g[4974] = a[10] & g[2926];
assign g[7021] = b[10] & g[2926];
assign g[4975] = a[10] & g[2927];
assign g[7022] = b[10] & g[2927];
assign g[4976] = a[10] & g[2928];
assign g[7023] = b[10] & g[2928];
assign g[4977] = a[10] & g[2929];
assign g[7024] = b[10] & g[2929];
assign g[4978] = a[10] & g[2930];
assign g[7025] = b[10] & g[2930];
assign g[4979] = a[10] & g[2931];
assign g[7026] = b[10] & g[2931];
assign g[4980] = a[10] & g[2932];
assign g[7027] = b[10] & g[2932];
assign g[4981] = a[10] & g[2933];
assign g[7028] = b[10] & g[2933];
assign g[4982] = a[10] & g[2934];
assign g[7029] = b[10] & g[2934];
assign g[4983] = a[10] & g[2935];
assign g[7030] = b[10] & g[2935];
assign g[4984] = a[10] & g[2936];
assign g[7031] = b[10] & g[2936];
assign g[4985] = a[10] & g[2937];
assign g[7032] = b[10] & g[2937];
assign g[4986] = a[10] & g[2938];
assign g[7033] = b[10] & g[2938];
assign g[4987] = a[10] & g[2939];
assign g[7034] = b[10] & g[2939];
assign g[4988] = a[10] & g[2940];
assign g[7035] = b[10] & g[2940];
assign g[4989] = a[10] & g[2941];
assign g[7036] = b[10] & g[2941];
assign g[4990] = a[10] & g[2942];
assign g[7037] = b[10] & g[2942];
assign g[4991] = a[10] & g[2943];
assign g[7038] = b[10] & g[2943];
assign g[4992] = a[10] & g[2944];
assign g[7039] = b[10] & g[2944];
assign g[4993] = a[10] & g[2945];
assign g[7040] = b[10] & g[2945];
assign g[4994] = a[10] & g[2946];
assign g[7041] = b[10] & g[2946];
assign g[4995] = a[10] & g[2947];
assign g[7042] = b[10] & g[2947];
assign g[4996] = a[10] & g[2948];
assign g[7043] = b[10] & g[2948];
assign g[4997] = a[10] & g[2949];
assign g[7044] = b[10] & g[2949];
assign g[4998] = a[10] & g[2950];
assign g[7045] = b[10] & g[2950];
assign g[4999] = a[10] & g[2951];
assign g[7046] = b[10] & g[2951];
assign g[5000] = a[10] & g[2952];
assign g[7047] = b[10] & g[2952];
assign g[5001] = a[10] & g[2953];
assign g[7048] = b[10] & g[2953];
assign g[5002] = a[10] & g[2954];
assign g[7049] = b[10] & g[2954];
assign g[5003] = a[10] & g[2955];
assign g[7050] = b[10] & g[2955];
assign g[5004] = a[10] & g[2956];
assign g[7051] = b[10] & g[2956];
assign g[5005] = a[10] & g[2957];
assign g[7052] = b[10] & g[2957];
assign g[5006] = a[10] & g[2958];
assign g[7053] = b[10] & g[2958];
assign g[5007] = a[10] & g[2959];
assign g[7054] = b[10] & g[2959];
assign g[5008] = a[10] & g[2960];
assign g[7055] = b[10] & g[2960];
assign g[5009] = a[10] & g[2961];
assign g[7056] = b[10] & g[2961];
assign g[5010] = a[10] & g[2962];
assign g[7057] = b[10] & g[2962];
assign g[5011] = a[10] & g[2963];
assign g[7058] = b[10] & g[2963];
assign g[5012] = a[10] & g[2964];
assign g[7059] = b[10] & g[2964];
assign g[5013] = a[10] & g[2965];
assign g[7060] = b[10] & g[2965];
assign g[5014] = a[10] & g[2966];
assign g[7061] = b[10] & g[2966];
assign g[5015] = a[10] & g[2967];
assign g[7062] = b[10] & g[2967];
assign g[5016] = a[10] & g[2968];
assign g[7063] = b[10] & g[2968];
assign g[5017] = a[10] & g[2969];
assign g[7064] = b[10] & g[2969];
assign g[5018] = a[10] & g[2970];
assign g[7065] = b[10] & g[2970];
assign g[5019] = a[10] & g[2971];
assign g[7066] = b[10] & g[2971];
assign g[5020] = a[10] & g[2972];
assign g[7067] = b[10] & g[2972];
assign g[5021] = a[10] & g[2973];
assign g[7068] = b[10] & g[2973];
assign g[5022] = a[10] & g[2974];
assign g[7069] = b[10] & g[2974];
assign g[5023] = a[10] & g[2975];
assign g[7070] = b[10] & g[2975];
assign g[5024] = a[10] & g[2976];
assign g[7071] = b[10] & g[2976];
assign g[5025] = a[10] & g[2977];
assign g[7072] = b[10] & g[2977];
assign g[5026] = a[10] & g[2978];
assign g[7073] = b[10] & g[2978];
assign g[5027] = a[10] & g[2979];
assign g[7074] = b[10] & g[2979];
assign g[5028] = a[10] & g[2980];
assign g[7075] = b[10] & g[2980];
assign g[5029] = a[10] & g[2981];
assign g[7076] = b[10] & g[2981];
assign g[5030] = a[10] & g[2982];
assign g[7077] = b[10] & g[2982];
assign g[5031] = a[10] & g[2983];
assign g[7078] = b[10] & g[2983];
assign g[5032] = a[10] & g[2984];
assign g[7079] = b[10] & g[2984];
assign g[5033] = a[10] & g[2985];
assign g[7080] = b[10] & g[2985];
assign g[5034] = a[10] & g[2986];
assign g[7081] = b[10] & g[2986];
assign g[5035] = a[10] & g[2987];
assign g[7082] = b[10] & g[2987];
assign g[5036] = a[10] & g[2988];
assign g[7083] = b[10] & g[2988];
assign g[5037] = a[10] & g[2989];
assign g[7084] = b[10] & g[2989];
assign g[5038] = a[10] & g[2990];
assign g[7085] = b[10] & g[2990];
assign g[5039] = a[10] & g[2991];
assign g[7086] = b[10] & g[2991];
assign g[5040] = a[10] & g[2992];
assign g[7087] = b[10] & g[2992];
assign g[5041] = a[10] & g[2993];
assign g[7088] = b[10] & g[2993];
assign g[5042] = a[10] & g[2994];
assign g[7089] = b[10] & g[2994];
assign g[5043] = a[10] & g[2995];
assign g[7090] = b[10] & g[2995];
assign g[5044] = a[10] & g[2996];
assign g[7091] = b[10] & g[2996];
assign g[5045] = a[10] & g[2997];
assign g[7092] = b[10] & g[2997];
assign g[5046] = a[10] & g[2998];
assign g[7093] = b[10] & g[2998];
assign g[5047] = a[10] & g[2999];
assign g[7094] = b[10] & g[2999];
assign g[5048] = a[10] & g[3000];
assign g[7095] = b[10] & g[3000];
assign g[5049] = a[10] & g[3001];
assign g[7096] = b[10] & g[3001];
assign g[5050] = a[10] & g[3002];
assign g[7097] = b[10] & g[3002];
assign g[5051] = a[10] & g[3003];
assign g[7098] = b[10] & g[3003];
assign g[5052] = a[10] & g[3004];
assign g[7099] = b[10] & g[3004];
assign g[5053] = a[10] & g[3005];
assign g[7100] = b[10] & g[3005];
assign g[5054] = a[10] & g[3006];
assign g[7101] = b[10] & g[3006];
assign g[5055] = a[10] & g[3007];
assign g[7102] = b[10] & g[3007];
assign g[5056] = a[10] & g[3008];
assign g[7103] = b[10] & g[3008];
assign g[5057] = a[10] & g[3009];
assign g[7104] = b[10] & g[3009];
assign g[5058] = a[10] & g[3010];
assign g[7105] = b[10] & g[3010];
assign g[5059] = a[10] & g[3011];
assign g[7106] = b[10] & g[3011];
assign g[5060] = a[10] & g[3012];
assign g[7107] = b[10] & g[3012];
assign g[5061] = a[10] & g[3013];
assign g[7108] = b[10] & g[3013];
assign g[5062] = a[10] & g[3014];
assign g[7109] = b[10] & g[3014];
assign g[5063] = a[10] & g[3015];
assign g[7110] = b[10] & g[3015];
assign g[5064] = a[10] & g[3016];
assign g[7111] = b[10] & g[3016];
assign g[5065] = a[10] & g[3017];
assign g[7112] = b[10] & g[3017];
assign g[5066] = a[10] & g[3018];
assign g[7113] = b[10] & g[3018];
assign g[5067] = a[10] & g[3019];
assign g[7114] = b[10] & g[3019];
assign g[5068] = a[10] & g[3020];
assign g[7115] = b[10] & g[3020];
assign g[5069] = a[10] & g[3021];
assign g[7116] = b[10] & g[3021];
assign g[5070] = a[10] & g[3022];
assign g[7117] = b[10] & g[3022];
assign g[5071] = a[10] & g[3023];
assign g[7118] = b[10] & g[3023];
assign g[5072] = a[10] & g[3024];
assign g[7119] = b[10] & g[3024];
assign g[5073] = a[10] & g[3025];
assign g[7120] = b[10] & g[3025];
assign g[5074] = a[10] & g[3026];
assign g[7121] = b[10] & g[3026];
assign g[5075] = a[10] & g[3027];
assign g[7122] = b[10] & g[3027];
assign g[5076] = a[10] & g[3028];
assign g[7123] = b[10] & g[3028];
assign g[5077] = a[10] & g[3029];
assign g[7124] = b[10] & g[3029];
assign g[5078] = a[10] & g[3030];
assign g[7125] = b[10] & g[3030];
assign g[5079] = a[10] & g[3031];
assign g[7126] = b[10] & g[3031];
assign g[5080] = a[10] & g[3032];
assign g[7127] = b[10] & g[3032];
assign g[5081] = a[10] & g[3033];
assign g[7128] = b[10] & g[3033];
assign g[5082] = a[10] & g[3034];
assign g[7129] = b[10] & g[3034];
assign g[5083] = a[10] & g[3035];
assign g[7130] = b[10] & g[3035];
assign g[5084] = a[10] & g[3036];
assign g[7131] = b[10] & g[3036];
assign g[5085] = a[10] & g[3037];
assign g[7132] = b[10] & g[3037];
assign g[5086] = a[10] & g[3038];
assign g[7133] = b[10] & g[3038];
assign g[5087] = a[10] & g[3039];
assign g[7134] = b[10] & g[3039];
assign g[5088] = a[10] & g[3040];
assign g[7135] = b[10] & g[3040];
assign g[5089] = a[10] & g[3041];
assign g[7136] = b[10] & g[3041];
assign g[5090] = a[10] & g[3042];
assign g[7137] = b[10] & g[3042];
assign g[5091] = a[10] & g[3043];
assign g[7138] = b[10] & g[3043];
assign g[5092] = a[10] & g[3044];
assign g[7139] = b[10] & g[3044];
assign g[5093] = a[10] & g[3045];
assign g[7140] = b[10] & g[3045];
assign g[5094] = a[10] & g[3046];
assign g[7141] = b[10] & g[3046];
assign g[5095] = a[10] & g[3047];
assign g[7142] = b[10] & g[3047];
assign g[5096] = a[10] & g[3048];
assign g[7143] = b[10] & g[3048];
assign g[5097] = a[10] & g[3049];
assign g[7144] = b[10] & g[3049];
assign g[5098] = a[10] & g[3050];
assign g[7145] = b[10] & g[3050];
assign g[5099] = a[10] & g[3051];
assign g[7146] = b[10] & g[3051];
assign g[5100] = a[10] & g[3052];
assign g[7147] = b[10] & g[3052];
assign g[5101] = a[10] & g[3053];
assign g[7148] = b[10] & g[3053];
assign g[5102] = a[10] & g[3054];
assign g[7149] = b[10] & g[3054];
assign g[5103] = a[10] & g[3055];
assign g[7150] = b[10] & g[3055];
assign g[5104] = a[10] & g[3056];
assign g[7151] = b[10] & g[3056];
assign g[5105] = a[10] & g[3057];
assign g[7152] = b[10] & g[3057];
assign g[5106] = a[10] & g[3058];
assign g[7153] = b[10] & g[3058];
assign g[5107] = a[10] & g[3059];
assign g[7154] = b[10] & g[3059];
assign g[5108] = a[10] & g[3060];
assign g[7155] = b[10] & g[3060];
assign g[5109] = a[10] & g[3061];
assign g[7156] = b[10] & g[3061];
assign g[5110] = a[10] & g[3062];
assign g[7157] = b[10] & g[3062];
assign g[5111] = a[10] & g[3063];
assign g[7158] = b[10] & g[3063];
assign g[5112] = a[10] & g[3064];
assign g[7159] = b[10] & g[3064];
assign g[5113] = a[10] & g[3065];
assign g[7160] = b[10] & g[3065];
assign g[5114] = a[10] & g[3066];
assign g[7161] = b[10] & g[3066];
assign g[5115] = a[10] & g[3067];
assign g[7162] = b[10] & g[3067];
assign g[5116] = a[10] & g[3068];
assign g[7163] = b[10] & g[3068];
assign g[5117] = a[10] & g[3069];
assign g[7164] = b[10] & g[3069];
assign g[5118] = a[10] & g[3070];
assign g[7165] = b[10] & g[3070];
assign g[5119] = a[10] & g[3071];
assign g[7166] = b[10] & g[3071];
assign g[5120] = a[10] & g[3072];
assign g[7167] = b[10] & g[3072];
assign g[5121] = a[10] & g[3073];
assign g[7168] = b[10] & g[3073];
assign g[5122] = a[10] & g[3074];
assign g[7169] = b[10] & g[3074];
assign g[5123] = a[10] & g[3075];
assign g[7170] = b[10] & g[3075];
assign g[5124] = a[10] & g[3076];
assign g[7171] = b[10] & g[3076];
assign g[5125] = a[10] & g[3077];
assign g[7172] = b[10] & g[3077];
assign g[5126] = a[10] & g[3078];
assign g[7173] = b[10] & g[3078];
assign g[5127] = a[10] & g[3079];
assign g[7174] = b[10] & g[3079];
assign g[5128] = a[10] & g[3080];
assign g[7175] = b[10] & g[3080];
assign g[5129] = a[10] & g[3081];
assign g[7176] = b[10] & g[3081];
assign g[5130] = a[10] & g[3082];
assign g[7177] = b[10] & g[3082];
assign g[5131] = a[10] & g[3083];
assign g[7178] = b[10] & g[3083];
assign g[5132] = a[10] & g[3084];
assign g[7179] = b[10] & g[3084];
assign g[5133] = a[10] & g[3085];
assign g[7180] = b[10] & g[3085];
assign g[5134] = a[10] & g[3086];
assign g[7181] = b[10] & g[3086];
assign g[5135] = a[10] & g[3087];
assign g[7182] = b[10] & g[3087];
assign g[5136] = a[10] & g[3088];
assign g[7183] = b[10] & g[3088];
assign g[5137] = a[10] & g[3089];
assign g[7184] = b[10] & g[3089];
assign g[5138] = a[10] & g[3090];
assign g[7185] = b[10] & g[3090];
assign g[5139] = a[10] & g[3091];
assign g[7186] = b[10] & g[3091];
assign g[5140] = a[10] & g[3092];
assign g[7187] = b[10] & g[3092];
assign g[5141] = a[10] & g[3093];
assign g[7188] = b[10] & g[3093];
assign g[5142] = a[10] & g[3094];
assign g[7189] = b[10] & g[3094];
assign g[5143] = a[10] & g[3095];
assign g[7190] = b[10] & g[3095];
assign g[5144] = a[10] & g[3096];
assign g[7191] = b[10] & g[3096];
assign g[5145] = a[10] & g[3097];
assign g[7192] = b[10] & g[3097];
assign g[5146] = a[10] & g[3098];
assign g[7193] = b[10] & g[3098];
assign g[5147] = a[10] & g[3099];
assign g[7194] = b[10] & g[3099];
assign g[5148] = a[10] & g[3100];
assign g[7195] = b[10] & g[3100];
assign g[5149] = a[10] & g[3101];
assign g[7196] = b[10] & g[3101];
assign g[5150] = a[10] & g[3102];
assign g[7197] = b[10] & g[3102];
assign g[5151] = a[10] & g[3103];
assign g[7198] = b[10] & g[3103];
assign g[5152] = a[10] & g[3104];
assign g[7199] = b[10] & g[3104];
assign g[5153] = a[10] & g[3105];
assign g[7200] = b[10] & g[3105];
assign g[5154] = a[10] & g[3106];
assign g[7201] = b[10] & g[3106];
assign g[5155] = a[10] & g[3107];
assign g[7202] = b[10] & g[3107];
assign g[5156] = a[10] & g[3108];
assign g[7203] = b[10] & g[3108];
assign g[5157] = a[10] & g[3109];
assign g[7204] = b[10] & g[3109];
assign g[5158] = a[10] & g[3110];
assign g[7205] = b[10] & g[3110];
assign g[5159] = a[10] & g[3111];
assign g[7206] = b[10] & g[3111];
assign g[5160] = a[10] & g[3112];
assign g[7207] = b[10] & g[3112];
assign g[5161] = a[10] & g[3113];
assign g[7208] = b[10] & g[3113];
assign g[5162] = a[10] & g[3114];
assign g[7209] = b[10] & g[3114];
assign g[5163] = a[10] & g[3115];
assign g[7210] = b[10] & g[3115];
assign g[5164] = a[10] & g[3116];
assign g[7211] = b[10] & g[3116];
assign g[5165] = a[10] & g[3117];
assign g[7212] = b[10] & g[3117];
assign g[5166] = a[10] & g[3118];
assign g[7213] = b[10] & g[3118];
assign g[5167] = a[10] & g[3119];
assign g[7214] = b[10] & g[3119];
assign g[5168] = a[10] & g[3120];
assign g[7215] = b[10] & g[3120];
assign g[5169] = a[10] & g[3121];
assign g[7216] = b[10] & g[3121];
assign g[5170] = a[10] & g[3122];
assign g[7217] = b[10] & g[3122];
assign g[5171] = a[10] & g[3123];
assign g[7218] = b[10] & g[3123];
assign g[5172] = a[10] & g[3124];
assign g[7219] = b[10] & g[3124];
assign g[5173] = a[10] & g[3125];
assign g[7220] = b[10] & g[3125];
assign g[5174] = a[10] & g[3126];
assign g[7221] = b[10] & g[3126];
assign g[5175] = a[10] & g[3127];
assign g[7222] = b[10] & g[3127];
assign g[5176] = a[10] & g[3128];
assign g[7223] = b[10] & g[3128];
assign g[5177] = a[10] & g[3129];
assign g[7224] = b[10] & g[3129];
assign g[5178] = a[10] & g[3130];
assign g[7225] = b[10] & g[3130];
assign g[5179] = a[10] & g[3131];
assign g[7226] = b[10] & g[3131];
assign g[5180] = a[10] & g[3132];
assign g[7227] = b[10] & g[3132];
assign g[5181] = a[10] & g[3133];
assign g[7228] = b[10] & g[3133];
assign g[5182] = a[10] & g[3134];
assign g[7229] = b[10] & g[3134];
assign g[5183] = a[10] & g[3135];
assign g[7230] = b[10] & g[3135];
assign g[5184] = a[10] & g[3136];
assign g[7231] = b[10] & g[3136];
assign g[5185] = a[10] & g[3137];
assign g[7232] = b[10] & g[3137];
assign g[5186] = a[10] & g[3138];
assign g[7233] = b[10] & g[3138];
assign g[5187] = a[10] & g[3139];
assign g[7234] = b[10] & g[3139];
assign g[5188] = a[10] & g[3140];
assign g[7235] = b[10] & g[3140];
assign g[5189] = a[10] & g[3141];
assign g[7236] = b[10] & g[3141];
assign g[5190] = a[10] & g[3142];
assign g[7237] = b[10] & g[3142];
assign g[5191] = a[10] & g[3143];
assign g[7238] = b[10] & g[3143];
assign g[5192] = a[10] & g[3144];
assign g[7239] = b[10] & g[3144];
assign g[5193] = a[10] & g[3145];
assign g[7240] = b[10] & g[3145];
assign g[5194] = a[10] & g[3146];
assign g[7241] = b[10] & g[3146];
assign g[5195] = a[10] & g[3147];
assign g[7242] = b[10] & g[3147];
assign g[5196] = a[10] & g[3148];
assign g[7243] = b[10] & g[3148];
assign g[5197] = a[10] & g[3149];
assign g[7244] = b[10] & g[3149];
assign g[5198] = a[10] & g[3150];
assign g[7245] = b[10] & g[3150];
assign g[5199] = a[10] & g[3151];
assign g[7246] = b[10] & g[3151];
assign g[5200] = a[10] & g[3152];
assign g[7247] = b[10] & g[3152];
assign g[5201] = a[10] & g[3153];
assign g[7248] = b[10] & g[3153];
assign g[5202] = a[10] & g[3154];
assign g[7249] = b[10] & g[3154];
assign g[5203] = a[10] & g[3155];
assign g[7250] = b[10] & g[3155];
assign g[5204] = a[10] & g[3156];
assign g[7251] = b[10] & g[3156];
assign g[5205] = a[10] & g[3157];
assign g[7252] = b[10] & g[3157];
assign g[5206] = a[10] & g[3158];
assign g[7253] = b[10] & g[3158];
assign g[5207] = a[10] & g[3159];
assign g[7254] = b[10] & g[3159];
assign g[5208] = a[10] & g[3160];
assign g[7255] = b[10] & g[3160];
assign g[5209] = a[10] & g[3161];
assign g[7256] = b[10] & g[3161];
assign g[5210] = a[10] & g[3162];
assign g[7257] = b[10] & g[3162];
assign g[5211] = a[10] & g[3163];
assign g[7258] = b[10] & g[3163];
assign g[5212] = a[10] & g[3164];
assign g[7259] = b[10] & g[3164];
assign g[5213] = a[10] & g[3165];
assign g[7260] = b[10] & g[3165];
assign g[5214] = a[10] & g[3166];
assign g[7261] = b[10] & g[3166];
assign g[5215] = a[10] & g[3167];
assign g[7262] = b[10] & g[3167];
assign g[5216] = a[10] & g[3168];
assign g[7263] = b[10] & g[3168];
assign g[5217] = a[10] & g[3169];
assign g[7264] = b[10] & g[3169];
assign g[5218] = a[10] & g[3170];
assign g[7265] = b[10] & g[3170];
assign g[5219] = a[10] & g[3171];
assign g[7266] = b[10] & g[3171];
assign g[5220] = a[10] & g[3172];
assign g[7267] = b[10] & g[3172];
assign g[5221] = a[10] & g[3173];
assign g[7268] = b[10] & g[3173];
assign g[5222] = a[10] & g[3174];
assign g[7269] = b[10] & g[3174];
assign g[5223] = a[10] & g[3175];
assign g[7270] = b[10] & g[3175];
assign g[5224] = a[10] & g[3176];
assign g[7271] = b[10] & g[3176];
assign g[5225] = a[10] & g[3177];
assign g[7272] = b[10] & g[3177];
assign g[5226] = a[10] & g[3178];
assign g[7273] = b[10] & g[3178];
assign g[5227] = a[10] & g[3179];
assign g[7274] = b[10] & g[3179];
assign g[5228] = a[10] & g[3180];
assign g[7275] = b[10] & g[3180];
assign g[5229] = a[10] & g[3181];
assign g[7276] = b[10] & g[3181];
assign g[5230] = a[10] & g[3182];
assign g[7277] = b[10] & g[3182];
assign g[5231] = a[10] & g[3183];
assign g[7278] = b[10] & g[3183];
assign g[5232] = a[10] & g[3184];
assign g[7279] = b[10] & g[3184];
assign g[5233] = a[10] & g[3185];
assign g[7280] = b[10] & g[3185];
assign g[5234] = a[10] & g[3186];
assign g[7281] = b[10] & g[3186];
assign g[5235] = a[10] & g[3187];
assign g[7282] = b[10] & g[3187];
assign g[5236] = a[10] & g[3188];
assign g[7283] = b[10] & g[3188];
assign g[5237] = a[10] & g[3189];
assign g[7284] = b[10] & g[3189];
assign g[5238] = a[10] & g[3190];
assign g[7285] = b[10] & g[3190];
assign g[5239] = a[10] & g[3191];
assign g[7286] = b[10] & g[3191];
assign g[5240] = a[10] & g[3192];
assign g[7287] = b[10] & g[3192];
assign g[5241] = a[10] & g[3193];
assign g[7288] = b[10] & g[3193];
assign g[5242] = a[10] & g[3194];
assign g[7289] = b[10] & g[3194];
assign g[5243] = a[10] & g[3195];
assign g[7290] = b[10] & g[3195];
assign g[5244] = a[10] & g[3196];
assign g[7291] = b[10] & g[3196];
assign g[5245] = a[10] & g[3197];
assign g[7292] = b[10] & g[3197];
assign g[5246] = a[10] & g[3198];
assign g[7293] = b[10] & g[3198];
assign g[5247] = a[10] & g[3199];
assign g[7294] = b[10] & g[3199];
assign g[5248] = a[10] & g[3200];
assign g[7295] = b[10] & g[3200];
assign g[5249] = a[10] & g[3201];
assign g[7296] = b[10] & g[3201];
assign g[5250] = a[10] & g[3202];
assign g[7297] = b[10] & g[3202];
assign g[5251] = a[10] & g[3203];
assign g[7298] = b[10] & g[3203];
assign g[5252] = a[10] & g[3204];
assign g[7299] = b[10] & g[3204];
assign g[5253] = a[10] & g[3205];
assign g[7300] = b[10] & g[3205];
assign g[5254] = a[10] & g[3206];
assign g[7301] = b[10] & g[3206];
assign g[5255] = a[10] & g[3207];
assign g[7302] = b[10] & g[3207];
assign g[5256] = a[10] & g[3208];
assign g[7303] = b[10] & g[3208];
assign g[5257] = a[10] & g[3209];
assign g[7304] = b[10] & g[3209];
assign g[5258] = a[10] & g[3210];
assign g[7305] = b[10] & g[3210];
assign g[5259] = a[10] & g[3211];
assign g[7306] = b[10] & g[3211];
assign g[5260] = a[10] & g[3212];
assign g[7307] = b[10] & g[3212];
assign g[5261] = a[10] & g[3213];
assign g[7308] = b[10] & g[3213];
assign g[5262] = a[10] & g[3214];
assign g[7309] = b[10] & g[3214];
assign g[5263] = a[10] & g[3215];
assign g[7310] = b[10] & g[3215];
assign g[5264] = a[10] & g[3216];
assign g[7311] = b[10] & g[3216];
assign g[5265] = a[10] & g[3217];
assign g[7312] = b[10] & g[3217];
assign g[5266] = a[10] & g[3218];
assign g[7313] = b[10] & g[3218];
assign g[5267] = a[10] & g[3219];
assign g[7314] = b[10] & g[3219];
assign g[5268] = a[10] & g[3220];
assign g[7315] = b[10] & g[3220];
assign g[5269] = a[10] & g[3221];
assign g[7316] = b[10] & g[3221];
assign g[5270] = a[10] & g[3222];
assign g[7317] = b[10] & g[3222];
assign g[5271] = a[10] & g[3223];
assign g[7318] = b[10] & g[3223];
assign g[5272] = a[10] & g[3224];
assign g[7319] = b[10] & g[3224];
assign g[5273] = a[10] & g[3225];
assign g[7320] = b[10] & g[3225];
assign g[5274] = a[10] & g[3226];
assign g[7321] = b[10] & g[3226];
assign g[5275] = a[10] & g[3227];
assign g[7322] = b[10] & g[3227];
assign g[5276] = a[10] & g[3228];
assign g[7323] = b[10] & g[3228];
assign g[5277] = a[10] & g[3229];
assign g[7324] = b[10] & g[3229];
assign g[5278] = a[10] & g[3230];
assign g[7325] = b[10] & g[3230];
assign g[5279] = a[10] & g[3231];
assign g[7326] = b[10] & g[3231];
assign g[5280] = a[10] & g[3232];
assign g[7327] = b[10] & g[3232];
assign g[5281] = a[10] & g[3233];
assign g[7328] = b[10] & g[3233];
assign g[5282] = a[10] & g[3234];
assign g[7329] = b[10] & g[3234];
assign g[5283] = a[10] & g[3235];
assign g[7330] = b[10] & g[3235];
assign g[5284] = a[10] & g[3236];
assign g[7331] = b[10] & g[3236];
assign g[5285] = a[10] & g[3237];
assign g[7332] = b[10] & g[3237];
assign g[5286] = a[10] & g[3238];
assign g[7333] = b[10] & g[3238];
assign g[5287] = a[10] & g[3239];
assign g[7334] = b[10] & g[3239];
assign g[5288] = a[10] & g[3240];
assign g[7335] = b[10] & g[3240];
assign g[5289] = a[10] & g[3241];
assign g[7336] = b[10] & g[3241];
assign g[5290] = a[10] & g[3242];
assign g[7337] = b[10] & g[3242];
assign g[5291] = a[10] & g[3243];
assign g[7338] = b[10] & g[3243];
assign g[5292] = a[10] & g[3244];
assign g[7339] = b[10] & g[3244];
assign g[5293] = a[10] & g[3245];
assign g[7340] = b[10] & g[3245];
assign g[5294] = a[10] & g[3246];
assign g[7341] = b[10] & g[3246];
assign g[5295] = a[10] & g[3247];
assign g[7342] = b[10] & g[3247];
assign g[5296] = a[10] & g[3248];
assign g[7343] = b[10] & g[3248];
assign g[5297] = a[10] & g[3249];
assign g[7344] = b[10] & g[3249];
assign g[5298] = a[10] & g[3250];
assign g[7345] = b[10] & g[3250];
assign g[5299] = a[10] & g[3251];
assign g[7346] = b[10] & g[3251];
assign g[5300] = a[10] & g[3252];
assign g[7347] = b[10] & g[3252];
assign g[5301] = a[10] & g[3253];
assign g[7348] = b[10] & g[3253];
assign g[5302] = a[10] & g[3254];
assign g[7349] = b[10] & g[3254];
assign g[5303] = a[10] & g[3255];
assign g[7350] = b[10] & g[3255];
assign g[5304] = a[10] & g[3256];
assign g[7351] = b[10] & g[3256];
assign g[5305] = a[10] & g[3257];
assign g[7352] = b[10] & g[3257];
assign g[5306] = a[10] & g[3258];
assign g[7353] = b[10] & g[3258];
assign g[5307] = a[10] & g[3259];
assign g[7354] = b[10] & g[3259];
assign g[5308] = a[10] & g[3260];
assign g[7355] = b[10] & g[3260];
assign g[5309] = a[10] & g[3261];
assign g[7356] = b[10] & g[3261];
assign g[5310] = a[10] & g[3262];
assign g[7357] = b[10] & g[3262];
assign g[5311] = a[10] & g[3263];
assign g[7358] = b[10] & g[3263];
assign g[5312] = a[10] & g[3264];
assign g[7359] = b[10] & g[3264];
assign g[5313] = a[10] & g[3265];
assign g[7360] = b[10] & g[3265];
assign g[5314] = a[10] & g[3266];
assign g[7361] = b[10] & g[3266];
assign g[5315] = a[10] & g[3267];
assign g[7362] = b[10] & g[3267];
assign g[5316] = a[10] & g[3268];
assign g[7363] = b[10] & g[3268];
assign g[5317] = a[10] & g[3269];
assign g[7364] = b[10] & g[3269];
assign g[5318] = a[10] & g[3270];
assign g[7365] = b[10] & g[3270];
assign g[5319] = a[10] & g[3271];
assign g[7366] = b[10] & g[3271];
assign g[5320] = a[10] & g[3272];
assign g[7367] = b[10] & g[3272];
assign g[5321] = a[10] & g[3273];
assign g[7368] = b[10] & g[3273];
assign g[5322] = a[10] & g[3274];
assign g[7369] = b[10] & g[3274];
assign g[5323] = a[10] & g[3275];
assign g[7370] = b[10] & g[3275];
assign g[5324] = a[10] & g[3276];
assign g[7371] = b[10] & g[3276];
assign g[5325] = a[10] & g[3277];
assign g[7372] = b[10] & g[3277];
assign g[5326] = a[10] & g[3278];
assign g[7373] = b[10] & g[3278];
assign g[5327] = a[10] & g[3279];
assign g[7374] = b[10] & g[3279];
assign g[5328] = a[10] & g[3280];
assign g[7375] = b[10] & g[3280];
assign g[5329] = a[10] & g[3281];
assign g[7376] = b[10] & g[3281];
assign g[5330] = a[10] & g[3282];
assign g[7377] = b[10] & g[3282];
assign g[5331] = a[10] & g[3283];
assign g[7378] = b[10] & g[3283];
assign g[5332] = a[10] & g[3284];
assign g[7379] = b[10] & g[3284];
assign g[5333] = a[10] & g[3285];
assign g[7380] = b[10] & g[3285];
assign g[5334] = a[10] & g[3286];
assign g[7381] = b[10] & g[3286];
assign g[5335] = a[10] & g[3287];
assign g[7382] = b[10] & g[3287];
assign g[5336] = a[10] & g[3288];
assign g[7383] = b[10] & g[3288];
assign g[5337] = a[10] & g[3289];
assign g[7384] = b[10] & g[3289];
assign g[5338] = a[10] & g[3290];
assign g[7385] = b[10] & g[3290];
assign g[5339] = a[10] & g[3291];
assign g[7386] = b[10] & g[3291];
assign g[5340] = a[10] & g[3292];
assign g[7387] = b[10] & g[3292];
assign g[5341] = a[10] & g[3293];
assign g[7388] = b[10] & g[3293];
assign g[5342] = a[10] & g[3294];
assign g[7389] = b[10] & g[3294];
assign g[5343] = a[10] & g[3295];
assign g[7390] = b[10] & g[3295];
assign g[5344] = a[10] & g[3296];
assign g[7391] = b[10] & g[3296];
assign g[5345] = a[10] & g[3297];
assign g[7392] = b[10] & g[3297];
assign g[5346] = a[10] & g[3298];
assign g[7393] = b[10] & g[3298];
assign g[5347] = a[10] & g[3299];
assign g[7394] = b[10] & g[3299];
assign g[5348] = a[10] & g[3300];
assign g[7395] = b[10] & g[3300];
assign g[5349] = a[10] & g[3301];
assign g[7396] = b[10] & g[3301];
assign g[5350] = a[10] & g[3302];
assign g[7397] = b[10] & g[3302];
assign g[5351] = a[10] & g[3303];
assign g[7398] = b[10] & g[3303];
assign g[5352] = a[10] & g[3304];
assign g[7399] = b[10] & g[3304];
assign g[5353] = a[10] & g[3305];
assign g[7400] = b[10] & g[3305];
assign g[5354] = a[10] & g[3306];
assign g[7401] = b[10] & g[3306];
assign g[5355] = a[10] & g[3307];
assign g[7402] = b[10] & g[3307];
assign g[5356] = a[10] & g[3308];
assign g[7403] = b[10] & g[3308];
assign g[5357] = a[10] & g[3309];
assign g[7404] = b[10] & g[3309];
assign g[5358] = a[10] & g[3310];
assign g[7405] = b[10] & g[3310];
assign g[5359] = a[10] & g[3311];
assign g[7406] = b[10] & g[3311];
assign g[5360] = a[10] & g[3312];
assign g[7407] = b[10] & g[3312];
assign g[5361] = a[10] & g[3313];
assign g[7408] = b[10] & g[3313];
assign g[5362] = a[10] & g[3314];
assign g[7409] = b[10] & g[3314];
assign g[5363] = a[10] & g[3315];
assign g[7410] = b[10] & g[3315];
assign g[5364] = a[10] & g[3316];
assign g[7411] = b[10] & g[3316];
assign g[5365] = a[10] & g[3317];
assign g[7412] = b[10] & g[3317];
assign g[5366] = a[10] & g[3318];
assign g[7413] = b[10] & g[3318];
assign g[5367] = a[10] & g[3319];
assign g[7414] = b[10] & g[3319];
assign g[5368] = a[10] & g[3320];
assign g[7415] = b[10] & g[3320];
assign g[5369] = a[10] & g[3321];
assign g[7416] = b[10] & g[3321];
assign g[5370] = a[10] & g[3322];
assign g[7417] = b[10] & g[3322];
assign g[5371] = a[10] & g[3323];
assign g[7418] = b[10] & g[3323];
assign g[5372] = a[10] & g[3324];
assign g[7419] = b[10] & g[3324];
assign g[5373] = a[10] & g[3325];
assign g[7420] = b[10] & g[3325];
assign g[5374] = a[10] & g[3326];
assign g[7421] = b[10] & g[3326];
assign g[5375] = a[10] & g[3327];
assign g[7422] = b[10] & g[3327];
assign g[5376] = a[10] & g[3328];
assign g[7423] = b[10] & g[3328];
assign g[5377] = a[10] & g[3329];
assign g[7424] = b[10] & g[3329];
assign g[5378] = a[10] & g[3330];
assign g[7425] = b[10] & g[3330];
assign g[5379] = a[10] & g[3331];
assign g[7426] = b[10] & g[3331];
assign g[5380] = a[10] & g[3332];
assign g[7427] = b[10] & g[3332];
assign g[5381] = a[10] & g[3333];
assign g[7428] = b[10] & g[3333];
assign g[5382] = a[10] & g[3334];
assign g[7429] = b[10] & g[3334];
assign g[5383] = a[10] & g[3335];
assign g[7430] = b[10] & g[3335];
assign g[5384] = a[10] & g[3336];
assign g[7431] = b[10] & g[3336];
assign g[5385] = a[10] & g[3337];
assign g[7432] = b[10] & g[3337];
assign g[5386] = a[10] & g[3338];
assign g[7433] = b[10] & g[3338];
assign g[5387] = a[10] & g[3339];
assign g[7434] = b[10] & g[3339];
assign g[5388] = a[10] & g[3340];
assign g[7435] = b[10] & g[3340];
assign g[5389] = a[10] & g[3341];
assign g[7436] = b[10] & g[3341];
assign g[5390] = a[10] & g[3342];
assign g[7437] = b[10] & g[3342];
assign g[5391] = a[10] & g[3343];
assign g[7438] = b[10] & g[3343];
assign g[5392] = a[10] & g[3344];
assign g[7439] = b[10] & g[3344];
assign g[5393] = a[10] & g[3345];
assign g[7440] = b[10] & g[3345];
assign g[5394] = a[10] & g[3346];
assign g[7441] = b[10] & g[3346];
assign g[5395] = a[10] & g[3347];
assign g[7442] = b[10] & g[3347];
assign g[5396] = a[10] & g[3348];
assign g[7443] = b[10] & g[3348];
assign g[5397] = a[10] & g[3349];
assign g[7444] = b[10] & g[3349];
assign g[5398] = a[10] & g[3350];
assign g[7445] = b[10] & g[3350];
assign g[5399] = a[10] & g[3351];
assign g[7446] = b[10] & g[3351];
assign g[5400] = a[10] & g[3352];
assign g[7447] = b[10] & g[3352];
assign g[5401] = a[10] & g[3353];
assign g[7448] = b[10] & g[3353];
assign g[5402] = a[10] & g[3354];
assign g[7449] = b[10] & g[3354];
assign g[5403] = a[10] & g[3355];
assign g[7450] = b[10] & g[3355];
assign g[5404] = a[10] & g[3356];
assign g[7451] = b[10] & g[3356];
assign g[5405] = a[10] & g[3357];
assign g[7452] = b[10] & g[3357];
assign g[5406] = a[10] & g[3358];
assign g[7453] = b[10] & g[3358];
assign g[5407] = a[10] & g[3359];
assign g[7454] = b[10] & g[3359];
assign g[5408] = a[10] & g[3360];
assign g[7455] = b[10] & g[3360];
assign g[5409] = a[10] & g[3361];
assign g[7456] = b[10] & g[3361];
assign g[5410] = a[10] & g[3362];
assign g[7457] = b[10] & g[3362];
assign g[5411] = a[10] & g[3363];
assign g[7458] = b[10] & g[3363];
assign g[5412] = a[10] & g[3364];
assign g[7459] = b[10] & g[3364];
assign g[5413] = a[10] & g[3365];
assign g[7460] = b[10] & g[3365];
assign g[5414] = a[10] & g[3366];
assign g[7461] = b[10] & g[3366];
assign g[5415] = a[10] & g[3367];
assign g[7462] = b[10] & g[3367];
assign g[5416] = a[10] & g[3368];
assign g[7463] = b[10] & g[3368];
assign g[5417] = a[10] & g[3369];
assign g[7464] = b[10] & g[3369];
assign g[5418] = a[10] & g[3370];
assign g[7465] = b[10] & g[3370];
assign g[5419] = a[10] & g[3371];
assign g[7466] = b[10] & g[3371];
assign g[5420] = a[10] & g[3372];
assign g[7467] = b[10] & g[3372];
assign g[5421] = a[10] & g[3373];
assign g[7468] = b[10] & g[3373];
assign g[5422] = a[10] & g[3374];
assign g[7469] = b[10] & g[3374];
assign g[5423] = a[10] & g[3375];
assign g[7470] = b[10] & g[3375];
assign g[5424] = a[10] & g[3376];
assign g[7471] = b[10] & g[3376];
assign g[5425] = a[10] & g[3377];
assign g[7472] = b[10] & g[3377];
assign g[5426] = a[10] & g[3378];
assign g[7473] = b[10] & g[3378];
assign g[5427] = a[10] & g[3379];
assign g[7474] = b[10] & g[3379];
assign g[5428] = a[10] & g[3380];
assign g[7475] = b[10] & g[3380];
assign g[5429] = a[10] & g[3381];
assign g[7476] = b[10] & g[3381];
assign g[5430] = a[10] & g[3382];
assign g[7477] = b[10] & g[3382];
assign g[5431] = a[10] & g[3383];
assign g[7478] = b[10] & g[3383];
assign g[5432] = a[10] & g[3384];
assign g[7479] = b[10] & g[3384];
assign g[5433] = a[10] & g[3385];
assign g[7480] = b[10] & g[3385];
assign g[5434] = a[10] & g[3386];
assign g[7481] = b[10] & g[3386];
assign g[5435] = a[10] & g[3387];
assign g[7482] = b[10] & g[3387];
assign g[5436] = a[10] & g[3388];
assign g[7483] = b[10] & g[3388];
assign g[5437] = a[10] & g[3389];
assign g[7484] = b[10] & g[3389];
assign g[5438] = a[10] & g[3390];
assign g[7485] = b[10] & g[3390];
assign g[5439] = a[10] & g[3391];
assign g[7486] = b[10] & g[3391];
assign g[5440] = a[10] & g[3392];
assign g[7487] = b[10] & g[3392];
assign g[5441] = a[10] & g[3393];
assign g[7488] = b[10] & g[3393];
assign g[5442] = a[10] & g[3394];
assign g[7489] = b[10] & g[3394];
assign g[5443] = a[10] & g[3395];
assign g[7490] = b[10] & g[3395];
assign g[5444] = a[10] & g[3396];
assign g[7491] = b[10] & g[3396];
assign g[5445] = a[10] & g[3397];
assign g[7492] = b[10] & g[3397];
assign g[5446] = a[10] & g[3398];
assign g[7493] = b[10] & g[3398];
assign g[5447] = a[10] & g[3399];
assign g[7494] = b[10] & g[3399];
assign g[5448] = a[10] & g[3400];
assign g[7495] = b[10] & g[3400];
assign g[5449] = a[10] & g[3401];
assign g[7496] = b[10] & g[3401];
assign g[5450] = a[10] & g[3402];
assign g[7497] = b[10] & g[3402];
assign g[5451] = a[10] & g[3403];
assign g[7498] = b[10] & g[3403];
assign g[5452] = a[10] & g[3404];
assign g[7499] = b[10] & g[3404];
assign g[5453] = a[10] & g[3405];
assign g[7500] = b[10] & g[3405];
assign g[5454] = a[10] & g[3406];
assign g[7501] = b[10] & g[3406];
assign g[5455] = a[10] & g[3407];
assign g[7502] = b[10] & g[3407];
assign g[5456] = a[10] & g[3408];
assign g[7503] = b[10] & g[3408];
assign g[5457] = a[10] & g[3409];
assign g[7504] = b[10] & g[3409];
assign g[5458] = a[10] & g[3410];
assign g[7505] = b[10] & g[3410];
assign g[5459] = a[10] & g[3411];
assign g[7506] = b[10] & g[3411];
assign g[5460] = a[10] & g[3412];
assign g[7507] = b[10] & g[3412];
assign g[5461] = a[10] & g[3413];
assign g[7508] = b[10] & g[3413];
assign g[5462] = a[10] & g[3414];
assign g[7509] = b[10] & g[3414];
assign g[5463] = a[10] & g[3415];
assign g[7510] = b[10] & g[3415];
assign g[5464] = a[10] & g[3416];
assign g[7511] = b[10] & g[3416];
assign g[5465] = a[10] & g[3417];
assign g[7512] = b[10] & g[3417];
assign g[5466] = a[10] & g[3418];
assign g[7513] = b[10] & g[3418];
assign g[5467] = a[10] & g[3419];
assign g[7514] = b[10] & g[3419];
assign g[5468] = a[10] & g[3420];
assign g[7515] = b[10] & g[3420];
assign g[5469] = a[10] & g[3421];
assign g[7516] = b[10] & g[3421];
assign g[5470] = a[10] & g[3422];
assign g[7517] = b[10] & g[3422];
assign g[5471] = a[10] & g[3423];
assign g[7518] = b[10] & g[3423];
assign g[5472] = a[10] & g[3424];
assign g[7519] = b[10] & g[3424];
assign g[5473] = a[10] & g[3425];
assign g[7520] = b[10] & g[3425];
assign g[5474] = a[10] & g[3426];
assign g[7521] = b[10] & g[3426];
assign g[5475] = a[10] & g[3427];
assign g[7522] = b[10] & g[3427];
assign g[5476] = a[10] & g[3428];
assign g[7523] = b[10] & g[3428];
assign g[5477] = a[10] & g[3429];
assign g[7524] = b[10] & g[3429];
assign g[5478] = a[10] & g[3430];
assign g[7525] = b[10] & g[3430];
assign g[5479] = a[10] & g[3431];
assign g[7526] = b[10] & g[3431];
assign g[5480] = a[10] & g[3432];
assign g[7527] = b[10] & g[3432];
assign g[5481] = a[10] & g[3433];
assign g[7528] = b[10] & g[3433];
assign g[5482] = a[10] & g[3434];
assign g[7529] = b[10] & g[3434];
assign g[5483] = a[10] & g[3435];
assign g[7530] = b[10] & g[3435];
assign g[5484] = a[10] & g[3436];
assign g[7531] = b[10] & g[3436];
assign g[5485] = a[10] & g[3437];
assign g[7532] = b[10] & g[3437];
assign g[5486] = a[10] & g[3438];
assign g[7533] = b[10] & g[3438];
assign g[5487] = a[10] & g[3439];
assign g[7534] = b[10] & g[3439];
assign g[5488] = a[10] & g[3440];
assign g[7535] = b[10] & g[3440];
assign g[5489] = a[10] & g[3441];
assign g[7536] = b[10] & g[3441];
assign g[5490] = a[10] & g[3442];
assign g[7537] = b[10] & g[3442];
assign g[5491] = a[10] & g[3443];
assign g[7538] = b[10] & g[3443];
assign g[5492] = a[10] & g[3444];
assign g[7539] = b[10] & g[3444];
assign g[5493] = a[10] & g[3445];
assign g[7540] = b[10] & g[3445];
assign g[5494] = a[10] & g[3446];
assign g[7541] = b[10] & g[3446];
assign g[5495] = a[10] & g[3447];
assign g[7542] = b[10] & g[3447];
assign g[5496] = a[10] & g[3448];
assign g[7543] = b[10] & g[3448];
assign g[5497] = a[10] & g[3449];
assign g[7544] = b[10] & g[3449];
assign g[5498] = a[10] & g[3450];
assign g[7545] = b[10] & g[3450];
assign g[5499] = a[10] & g[3451];
assign g[7546] = b[10] & g[3451];
assign g[5500] = a[10] & g[3452];
assign g[7547] = b[10] & g[3452];
assign g[5501] = a[10] & g[3453];
assign g[7548] = b[10] & g[3453];
assign g[5502] = a[10] & g[3454];
assign g[7549] = b[10] & g[3454];
assign g[5503] = a[10] & g[3455];
assign g[7550] = b[10] & g[3455];
assign g[5504] = a[10] & g[3456];
assign g[7551] = b[10] & g[3456];
assign g[5505] = a[10] & g[3457];
assign g[7552] = b[10] & g[3457];
assign g[5506] = a[10] & g[3458];
assign g[7553] = b[10] & g[3458];
assign g[5507] = a[10] & g[3459];
assign g[7554] = b[10] & g[3459];
assign g[5508] = a[10] & g[3460];
assign g[7555] = b[10] & g[3460];
assign g[5509] = a[10] & g[3461];
assign g[7556] = b[10] & g[3461];
assign g[5510] = a[10] & g[3462];
assign g[7557] = b[10] & g[3462];
assign g[5511] = a[10] & g[3463];
assign g[7558] = b[10] & g[3463];
assign g[5512] = a[10] & g[3464];
assign g[7559] = b[10] & g[3464];
assign g[5513] = a[10] & g[3465];
assign g[7560] = b[10] & g[3465];
assign g[5514] = a[10] & g[3466];
assign g[7561] = b[10] & g[3466];
assign g[5515] = a[10] & g[3467];
assign g[7562] = b[10] & g[3467];
assign g[5516] = a[10] & g[3468];
assign g[7563] = b[10] & g[3468];
assign g[5517] = a[10] & g[3469];
assign g[7564] = b[10] & g[3469];
assign g[5518] = a[10] & g[3470];
assign g[7565] = b[10] & g[3470];
assign g[5519] = a[10] & g[3471];
assign g[7566] = b[10] & g[3471];
assign g[5520] = a[10] & g[3472];
assign g[7567] = b[10] & g[3472];
assign g[5521] = a[10] & g[3473];
assign g[7568] = b[10] & g[3473];
assign g[5522] = a[10] & g[3474];
assign g[7569] = b[10] & g[3474];
assign g[5523] = a[10] & g[3475];
assign g[7570] = b[10] & g[3475];
assign g[5524] = a[10] & g[3476];
assign g[7571] = b[10] & g[3476];
assign g[5525] = a[10] & g[3477];
assign g[7572] = b[10] & g[3477];
assign g[5526] = a[10] & g[3478];
assign g[7573] = b[10] & g[3478];
assign g[5527] = a[10] & g[3479];
assign g[7574] = b[10] & g[3479];
assign g[5528] = a[10] & g[3480];
assign g[7575] = b[10] & g[3480];
assign g[5529] = a[10] & g[3481];
assign g[7576] = b[10] & g[3481];
assign g[5530] = a[10] & g[3482];
assign g[7577] = b[10] & g[3482];
assign g[5531] = a[10] & g[3483];
assign g[7578] = b[10] & g[3483];
assign g[5532] = a[10] & g[3484];
assign g[7579] = b[10] & g[3484];
assign g[5533] = a[10] & g[3485];
assign g[7580] = b[10] & g[3485];
assign g[5534] = a[10] & g[3486];
assign g[7581] = b[10] & g[3486];
assign g[5535] = a[10] & g[3487];
assign g[7582] = b[10] & g[3487];
assign g[5536] = a[10] & g[3488];
assign g[7583] = b[10] & g[3488];
assign g[5537] = a[10] & g[3489];
assign g[7584] = b[10] & g[3489];
assign g[5538] = a[10] & g[3490];
assign g[7585] = b[10] & g[3490];
assign g[5539] = a[10] & g[3491];
assign g[7586] = b[10] & g[3491];
assign g[5540] = a[10] & g[3492];
assign g[7587] = b[10] & g[3492];
assign g[5541] = a[10] & g[3493];
assign g[7588] = b[10] & g[3493];
assign g[5542] = a[10] & g[3494];
assign g[7589] = b[10] & g[3494];
assign g[5543] = a[10] & g[3495];
assign g[7590] = b[10] & g[3495];
assign g[5544] = a[10] & g[3496];
assign g[7591] = b[10] & g[3496];
assign g[5545] = a[10] & g[3497];
assign g[7592] = b[10] & g[3497];
assign g[5546] = a[10] & g[3498];
assign g[7593] = b[10] & g[3498];
assign g[5547] = a[10] & g[3499];
assign g[7594] = b[10] & g[3499];
assign g[5548] = a[10] & g[3500];
assign g[7595] = b[10] & g[3500];
assign g[5549] = a[10] & g[3501];
assign g[7596] = b[10] & g[3501];
assign g[5550] = a[10] & g[3502];
assign g[7597] = b[10] & g[3502];
assign g[5551] = a[10] & g[3503];
assign g[7598] = b[10] & g[3503];
assign g[5552] = a[10] & g[3504];
assign g[7599] = b[10] & g[3504];
assign g[5553] = a[10] & g[3505];
assign g[7600] = b[10] & g[3505];
assign g[5554] = a[10] & g[3506];
assign g[7601] = b[10] & g[3506];
assign g[5555] = a[10] & g[3507];
assign g[7602] = b[10] & g[3507];
assign g[5556] = a[10] & g[3508];
assign g[7603] = b[10] & g[3508];
assign g[5557] = a[10] & g[3509];
assign g[7604] = b[10] & g[3509];
assign g[5558] = a[10] & g[3510];
assign g[7605] = b[10] & g[3510];
assign g[5559] = a[10] & g[3511];
assign g[7606] = b[10] & g[3511];
assign g[5560] = a[10] & g[3512];
assign g[7607] = b[10] & g[3512];
assign g[5561] = a[10] & g[3513];
assign g[7608] = b[10] & g[3513];
assign g[5562] = a[10] & g[3514];
assign g[7609] = b[10] & g[3514];
assign g[5563] = a[10] & g[3515];
assign g[7610] = b[10] & g[3515];
assign g[5564] = a[10] & g[3516];
assign g[7611] = b[10] & g[3516];
assign g[5565] = a[10] & g[3517];
assign g[7612] = b[10] & g[3517];
assign g[5566] = a[10] & g[3518];
assign g[7613] = b[10] & g[3518];
assign g[5567] = a[10] & g[3519];
assign g[7614] = b[10] & g[3519];
assign g[5568] = a[10] & g[3520];
assign g[7615] = b[10] & g[3520];
assign g[5569] = a[10] & g[3521];
assign g[7616] = b[10] & g[3521];
assign g[5570] = a[10] & g[3522];
assign g[7617] = b[10] & g[3522];
assign g[5571] = a[10] & g[3523];
assign g[7618] = b[10] & g[3523];
assign g[5572] = a[10] & g[3524];
assign g[7619] = b[10] & g[3524];
assign g[5573] = a[10] & g[3525];
assign g[7620] = b[10] & g[3525];
assign g[5574] = a[10] & g[3526];
assign g[7621] = b[10] & g[3526];
assign g[5575] = a[10] & g[3527];
assign g[7622] = b[10] & g[3527];
assign g[5576] = a[10] & g[3528];
assign g[7623] = b[10] & g[3528];
assign g[5577] = a[10] & g[3529];
assign g[7624] = b[10] & g[3529];
assign g[5578] = a[10] & g[3530];
assign g[7625] = b[10] & g[3530];
assign g[5579] = a[10] & g[3531];
assign g[7626] = b[10] & g[3531];
assign g[5580] = a[10] & g[3532];
assign g[7627] = b[10] & g[3532];
assign g[5581] = a[10] & g[3533];
assign g[7628] = b[10] & g[3533];
assign g[5582] = a[10] & g[3534];
assign g[7629] = b[10] & g[3534];
assign g[5583] = a[10] & g[3535];
assign g[7630] = b[10] & g[3535];
assign g[5584] = a[10] & g[3536];
assign g[7631] = b[10] & g[3536];
assign g[5585] = a[10] & g[3537];
assign g[7632] = b[10] & g[3537];
assign g[5586] = a[10] & g[3538];
assign g[7633] = b[10] & g[3538];
assign g[5587] = a[10] & g[3539];
assign g[7634] = b[10] & g[3539];
assign g[5588] = a[10] & g[3540];
assign g[7635] = b[10] & g[3540];
assign g[5589] = a[10] & g[3541];
assign g[7636] = b[10] & g[3541];
assign g[5590] = a[10] & g[3542];
assign g[7637] = b[10] & g[3542];
assign g[5591] = a[10] & g[3543];
assign g[7638] = b[10] & g[3543];
assign g[5592] = a[10] & g[3544];
assign g[7639] = b[10] & g[3544];
assign g[5593] = a[10] & g[3545];
assign g[7640] = b[10] & g[3545];
assign g[5594] = a[10] & g[3546];
assign g[7641] = b[10] & g[3546];
assign g[5595] = a[10] & g[3547];
assign g[7642] = b[10] & g[3547];
assign g[5596] = a[10] & g[3548];
assign g[7643] = b[10] & g[3548];
assign g[5597] = a[10] & g[3549];
assign g[7644] = b[10] & g[3549];
assign g[5598] = a[10] & g[3550];
assign g[7645] = b[10] & g[3550];
assign g[5599] = a[10] & g[3551];
assign g[7646] = b[10] & g[3551];
assign g[5600] = a[10] & g[3552];
assign g[7647] = b[10] & g[3552];
assign g[5601] = a[10] & g[3553];
assign g[7648] = b[10] & g[3553];
assign g[5602] = a[10] & g[3554];
assign g[7649] = b[10] & g[3554];
assign g[5603] = a[10] & g[3555];
assign g[7650] = b[10] & g[3555];
assign g[5604] = a[10] & g[3556];
assign g[7651] = b[10] & g[3556];
assign g[5605] = a[10] & g[3557];
assign g[7652] = b[10] & g[3557];
assign g[5606] = a[10] & g[3558];
assign g[7653] = b[10] & g[3558];
assign g[5607] = a[10] & g[3559];
assign g[7654] = b[10] & g[3559];
assign g[5608] = a[10] & g[3560];
assign g[7655] = b[10] & g[3560];
assign g[5609] = a[10] & g[3561];
assign g[7656] = b[10] & g[3561];
assign g[5610] = a[10] & g[3562];
assign g[7657] = b[10] & g[3562];
assign g[5611] = a[10] & g[3563];
assign g[7658] = b[10] & g[3563];
assign g[5612] = a[10] & g[3564];
assign g[7659] = b[10] & g[3564];
assign g[5613] = a[10] & g[3565];
assign g[7660] = b[10] & g[3565];
assign g[5614] = a[10] & g[3566];
assign g[7661] = b[10] & g[3566];
assign g[5615] = a[10] & g[3567];
assign g[7662] = b[10] & g[3567];
assign g[5616] = a[10] & g[3568];
assign g[7663] = b[10] & g[3568];
assign g[5617] = a[10] & g[3569];
assign g[7664] = b[10] & g[3569];
assign g[5618] = a[10] & g[3570];
assign g[7665] = b[10] & g[3570];
assign g[5619] = a[10] & g[3571];
assign g[7666] = b[10] & g[3571];
assign g[5620] = a[10] & g[3572];
assign g[7667] = b[10] & g[3572];
assign g[5621] = a[10] & g[3573];
assign g[7668] = b[10] & g[3573];
assign g[5622] = a[10] & g[3574];
assign g[7669] = b[10] & g[3574];
assign g[5623] = a[10] & g[3575];
assign g[7670] = b[10] & g[3575];
assign g[5624] = a[10] & g[3576];
assign g[7671] = b[10] & g[3576];
assign g[5625] = a[10] & g[3577];
assign g[7672] = b[10] & g[3577];
assign g[5626] = a[10] & g[3578];
assign g[7673] = b[10] & g[3578];
assign g[5627] = a[10] & g[3579];
assign g[7674] = b[10] & g[3579];
assign g[5628] = a[10] & g[3580];
assign g[7675] = b[10] & g[3580];
assign g[5629] = a[10] & g[3581];
assign g[7676] = b[10] & g[3581];
assign g[5630] = a[10] & g[3582];
assign g[7677] = b[10] & g[3582];
assign g[5631] = a[10] & g[3583];
assign g[7678] = b[10] & g[3583];
assign g[5632] = a[10] & g[3584];
assign g[7679] = b[10] & g[3584];
assign g[5633] = a[10] & g[3585];
assign g[7680] = b[10] & g[3585];
assign g[5634] = a[10] & g[3586];
assign g[7681] = b[10] & g[3586];
assign g[5635] = a[10] & g[3587];
assign g[7682] = b[10] & g[3587];
assign g[5636] = a[10] & g[3588];
assign g[7683] = b[10] & g[3588];
assign g[5637] = a[10] & g[3589];
assign g[7684] = b[10] & g[3589];
assign g[5638] = a[10] & g[3590];
assign g[7685] = b[10] & g[3590];
assign g[5639] = a[10] & g[3591];
assign g[7686] = b[10] & g[3591];
assign g[5640] = a[10] & g[3592];
assign g[7687] = b[10] & g[3592];
assign g[5641] = a[10] & g[3593];
assign g[7688] = b[10] & g[3593];
assign g[5642] = a[10] & g[3594];
assign g[7689] = b[10] & g[3594];
assign g[5643] = a[10] & g[3595];
assign g[7690] = b[10] & g[3595];
assign g[5644] = a[10] & g[3596];
assign g[7691] = b[10] & g[3596];
assign g[5645] = a[10] & g[3597];
assign g[7692] = b[10] & g[3597];
assign g[5646] = a[10] & g[3598];
assign g[7693] = b[10] & g[3598];
assign g[5647] = a[10] & g[3599];
assign g[7694] = b[10] & g[3599];
assign g[5648] = a[10] & g[3600];
assign g[7695] = b[10] & g[3600];
assign g[5649] = a[10] & g[3601];
assign g[7696] = b[10] & g[3601];
assign g[5650] = a[10] & g[3602];
assign g[7697] = b[10] & g[3602];
assign g[5651] = a[10] & g[3603];
assign g[7698] = b[10] & g[3603];
assign g[5652] = a[10] & g[3604];
assign g[7699] = b[10] & g[3604];
assign g[5653] = a[10] & g[3605];
assign g[7700] = b[10] & g[3605];
assign g[5654] = a[10] & g[3606];
assign g[7701] = b[10] & g[3606];
assign g[5655] = a[10] & g[3607];
assign g[7702] = b[10] & g[3607];
assign g[5656] = a[10] & g[3608];
assign g[7703] = b[10] & g[3608];
assign g[5657] = a[10] & g[3609];
assign g[7704] = b[10] & g[3609];
assign g[5658] = a[10] & g[3610];
assign g[7705] = b[10] & g[3610];
assign g[5659] = a[10] & g[3611];
assign g[7706] = b[10] & g[3611];
assign g[5660] = a[10] & g[3612];
assign g[7707] = b[10] & g[3612];
assign g[5661] = a[10] & g[3613];
assign g[7708] = b[10] & g[3613];
assign g[5662] = a[10] & g[3614];
assign g[7709] = b[10] & g[3614];
assign g[5663] = a[10] & g[3615];
assign g[7710] = b[10] & g[3615];
assign g[5664] = a[10] & g[3616];
assign g[7711] = b[10] & g[3616];
assign g[5665] = a[10] & g[3617];
assign g[7712] = b[10] & g[3617];
assign g[5666] = a[10] & g[3618];
assign g[7713] = b[10] & g[3618];
assign g[5667] = a[10] & g[3619];
assign g[7714] = b[10] & g[3619];
assign g[5668] = a[10] & g[3620];
assign g[7715] = b[10] & g[3620];
assign g[5669] = a[10] & g[3621];
assign g[7716] = b[10] & g[3621];
assign g[5670] = a[10] & g[3622];
assign g[7717] = b[10] & g[3622];
assign g[5671] = a[10] & g[3623];
assign g[7718] = b[10] & g[3623];
assign g[5672] = a[10] & g[3624];
assign g[7719] = b[10] & g[3624];
assign g[5673] = a[10] & g[3625];
assign g[7720] = b[10] & g[3625];
assign g[5674] = a[10] & g[3626];
assign g[7721] = b[10] & g[3626];
assign g[5675] = a[10] & g[3627];
assign g[7722] = b[10] & g[3627];
assign g[5676] = a[10] & g[3628];
assign g[7723] = b[10] & g[3628];
assign g[5677] = a[10] & g[3629];
assign g[7724] = b[10] & g[3629];
assign g[5678] = a[10] & g[3630];
assign g[7725] = b[10] & g[3630];
assign g[5679] = a[10] & g[3631];
assign g[7726] = b[10] & g[3631];
assign g[5680] = a[10] & g[3632];
assign g[7727] = b[10] & g[3632];
assign g[5681] = a[10] & g[3633];
assign g[7728] = b[10] & g[3633];
assign g[5682] = a[10] & g[3634];
assign g[7729] = b[10] & g[3634];
assign g[5683] = a[10] & g[3635];
assign g[7730] = b[10] & g[3635];
assign g[5684] = a[10] & g[3636];
assign g[7731] = b[10] & g[3636];
assign g[5685] = a[10] & g[3637];
assign g[7732] = b[10] & g[3637];
assign g[5686] = a[10] & g[3638];
assign g[7733] = b[10] & g[3638];
assign g[5687] = a[10] & g[3639];
assign g[7734] = b[10] & g[3639];
assign g[5688] = a[10] & g[3640];
assign g[7735] = b[10] & g[3640];
assign g[5689] = a[10] & g[3641];
assign g[7736] = b[10] & g[3641];
assign g[5690] = a[10] & g[3642];
assign g[7737] = b[10] & g[3642];
assign g[5691] = a[10] & g[3643];
assign g[7738] = b[10] & g[3643];
assign g[5692] = a[10] & g[3644];
assign g[7739] = b[10] & g[3644];
assign g[5693] = a[10] & g[3645];
assign g[7740] = b[10] & g[3645];
assign g[5694] = a[10] & g[3646];
assign g[7741] = b[10] & g[3646];
assign g[5695] = a[10] & g[3647];
assign g[7742] = b[10] & g[3647];
assign g[5696] = a[10] & g[3648];
assign g[7743] = b[10] & g[3648];
assign g[5697] = a[10] & g[3649];
assign g[7744] = b[10] & g[3649];
assign g[5698] = a[10] & g[3650];
assign g[7745] = b[10] & g[3650];
assign g[5699] = a[10] & g[3651];
assign g[7746] = b[10] & g[3651];
assign g[5700] = a[10] & g[3652];
assign g[7747] = b[10] & g[3652];
assign g[5701] = a[10] & g[3653];
assign g[7748] = b[10] & g[3653];
assign g[5702] = a[10] & g[3654];
assign g[7749] = b[10] & g[3654];
assign g[5703] = a[10] & g[3655];
assign g[7750] = b[10] & g[3655];
assign g[5704] = a[10] & g[3656];
assign g[7751] = b[10] & g[3656];
assign g[5705] = a[10] & g[3657];
assign g[7752] = b[10] & g[3657];
assign g[5706] = a[10] & g[3658];
assign g[7753] = b[10] & g[3658];
assign g[5707] = a[10] & g[3659];
assign g[7754] = b[10] & g[3659];
assign g[5708] = a[10] & g[3660];
assign g[7755] = b[10] & g[3660];
assign g[5709] = a[10] & g[3661];
assign g[7756] = b[10] & g[3661];
assign g[5710] = a[10] & g[3662];
assign g[7757] = b[10] & g[3662];
assign g[5711] = a[10] & g[3663];
assign g[7758] = b[10] & g[3663];
assign g[5712] = a[10] & g[3664];
assign g[7759] = b[10] & g[3664];
assign g[5713] = a[10] & g[3665];
assign g[7760] = b[10] & g[3665];
assign g[5714] = a[10] & g[3666];
assign g[7761] = b[10] & g[3666];
assign g[5715] = a[10] & g[3667];
assign g[7762] = b[10] & g[3667];
assign g[5716] = a[10] & g[3668];
assign g[7763] = b[10] & g[3668];
assign g[5717] = a[10] & g[3669];
assign g[7764] = b[10] & g[3669];
assign g[5718] = a[10] & g[3670];
assign g[7765] = b[10] & g[3670];
assign g[5719] = a[10] & g[3671];
assign g[7766] = b[10] & g[3671];
assign g[5720] = a[10] & g[3672];
assign g[7767] = b[10] & g[3672];
assign g[5721] = a[10] & g[3673];
assign g[7768] = b[10] & g[3673];
assign g[5722] = a[10] & g[3674];
assign g[7769] = b[10] & g[3674];
assign g[5723] = a[10] & g[3675];
assign g[7770] = b[10] & g[3675];
assign g[5724] = a[10] & g[3676];
assign g[7771] = b[10] & g[3676];
assign g[5725] = a[10] & g[3677];
assign g[7772] = b[10] & g[3677];
assign g[5726] = a[10] & g[3678];
assign g[7773] = b[10] & g[3678];
assign g[5727] = a[10] & g[3679];
assign g[7774] = b[10] & g[3679];
assign g[5728] = a[10] & g[3680];
assign g[7775] = b[10] & g[3680];
assign g[5729] = a[10] & g[3681];
assign g[7776] = b[10] & g[3681];
assign g[5730] = a[10] & g[3682];
assign g[7777] = b[10] & g[3682];
assign g[5731] = a[10] & g[3683];
assign g[7778] = b[10] & g[3683];
assign g[5732] = a[10] & g[3684];
assign g[7779] = b[10] & g[3684];
assign g[5733] = a[10] & g[3685];
assign g[7780] = b[10] & g[3685];
assign g[5734] = a[10] & g[3686];
assign g[7781] = b[10] & g[3686];
assign g[5735] = a[10] & g[3687];
assign g[7782] = b[10] & g[3687];
assign g[5736] = a[10] & g[3688];
assign g[7783] = b[10] & g[3688];
assign g[5737] = a[10] & g[3689];
assign g[7784] = b[10] & g[3689];
assign g[5738] = a[10] & g[3690];
assign g[7785] = b[10] & g[3690];
assign g[5739] = a[10] & g[3691];
assign g[7786] = b[10] & g[3691];
assign g[5740] = a[10] & g[3692];
assign g[7787] = b[10] & g[3692];
assign g[5741] = a[10] & g[3693];
assign g[7788] = b[10] & g[3693];
assign g[5742] = a[10] & g[3694];
assign g[7789] = b[10] & g[3694];
assign g[5743] = a[10] & g[3695];
assign g[7790] = b[10] & g[3695];
assign g[5744] = a[10] & g[3696];
assign g[7791] = b[10] & g[3696];
assign g[5745] = a[10] & g[3697];
assign g[7792] = b[10] & g[3697];
assign g[5746] = a[10] & g[3698];
assign g[7793] = b[10] & g[3698];
assign g[5747] = a[10] & g[3699];
assign g[7794] = b[10] & g[3699];
assign g[5748] = a[10] & g[3700];
assign g[7795] = b[10] & g[3700];
assign g[5749] = a[10] & g[3701];
assign g[7796] = b[10] & g[3701];
assign g[5750] = a[10] & g[3702];
assign g[7797] = b[10] & g[3702];
assign g[5751] = a[10] & g[3703];
assign g[7798] = b[10] & g[3703];
assign g[5752] = a[10] & g[3704];
assign g[7799] = b[10] & g[3704];
assign g[5753] = a[10] & g[3705];
assign g[7800] = b[10] & g[3705];
assign g[5754] = a[10] & g[3706];
assign g[7801] = b[10] & g[3706];
assign g[5755] = a[10] & g[3707];
assign g[7802] = b[10] & g[3707];
assign g[5756] = a[10] & g[3708];
assign g[7803] = b[10] & g[3708];
assign g[5757] = a[10] & g[3709];
assign g[7804] = b[10] & g[3709];
assign g[5758] = a[10] & g[3710];
assign g[7805] = b[10] & g[3710];
assign g[5759] = a[10] & g[3711];
assign g[7806] = b[10] & g[3711];
assign g[5760] = a[10] & g[3712];
assign g[7807] = b[10] & g[3712];
assign g[5761] = a[10] & g[3713];
assign g[7808] = b[10] & g[3713];
assign g[5762] = a[10] & g[3714];
assign g[7809] = b[10] & g[3714];
assign g[5763] = a[10] & g[3715];
assign g[7810] = b[10] & g[3715];
assign g[5764] = a[10] & g[3716];
assign g[7811] = b[10] & g[3716];
assign g[5765] = a[10] & g[3717];
assign g[7812] = b[10] & g[3717];
assign g[5766] = a[10] & g[3718];
assign g[7813] = b[10] & g[3718];
assign g[5767] = a[10] & g[3719];
assign g[7814] = b[10] & g[3719];
assign g[5768] = a[10] & g[3720];
assign g[7815] = b[10] & g[3720];
assign g[5769] = a[10] & g[3721];
assign g[7816] = b[10] & g[3721];
assign g[5770] = a[10] & g[3722];
assign g[7817] = b[10] & g[3722];
assign g[5771] = a[10] & g[3723];
assign g[7818] = b[10] & g[3723];
assign g[5772] = a[10] & g[3724];
assign g[7819] = b[10] & g[3724];
assign g[5773] = a[10] & g[3725];
assign g[7820] = b[10] & g[3725];
assign g[5774] = a[10] & g[3726];
assign g[7821] = b[10] & g[3726];
assign g[5775] = a[10] & g[3727];
assign g[7822] = b[10] & g[3727];
assign g[5776] = a[10] & g[3728];
assign g[7823] = b[10] & g[3728];
assign g[5777] = a[10] & g[3729];
assign g[7824] = b[10] & g[3729];
assign g[5778] = a[10] & g[3730];
assign g[7825] = b[10] & g[3730];
assign g[5779] = a[10] & g[3731];
assign g[7826] = b[10] & g[3731];
assign g[5780] = a[10] & g[3732];
assign g[7827] = b[10] & g[3732];
assign g[5781] = a[10] & g[3733];
assign g[7828] = b[10] & g[3733];
assign g[5782] = a[10] & g[3734];
assign g[7829] = b[10] & g[3734];
assign g[5783] = a[10] & g[3735];
assign g[7830] = b[10] & g[3735];
assign g[5784] = a[10] & g[3736];
assign g[7831] = b[10] & g[3736];
assign g[5785] = a[10] & g[3737];
assign g[7832] = b[10] & g[3737];
assign g[5786] = a[10] & g[3738];
assign g[7833] = b[10] & g[3738];
assign g[5787] = a[10] & g[3739];
assign g[7834] = b[10] & g[3739];
assign g[5788] = a[10] & g[3740];
assign g[7835] = b[10] & g[3740];
assign g[5789] = a[10] & g[3741];
assign g[7836] = b[10] & g[3741];
assign g[5790] = a[10] & g[3742];
assign g[7837] = b[10] & g[3742];
assign g[5791] = a[10] & g[3743];
assign g[7838] = b[10] & g[3743];
assign g[5792] = a[10] & g[3744];
assign g[7839] = b[10] & g[3744];
assign g[5793] = a[10] & g[3745];
assign g[7840] = b[10] & g[3745];
assign g[5794] = a[10] & g[3746];
assign g[7841] = b[10] & g[3746];
assign g[5795] = a[10] & g[3747];
assign g[7842] = b[10] & g[3747];
assign g[5796] = a[10] & g[3748];
assign g[7843] = b[10] & g[3748];
assign g[5797] = a[10] & g[3749];
assign g[7844] = b[10] & g[3749];
assign g[5798] = a[10] & g[3750];
assign g[7845] = b[10] & g[3750];
assign g[5799] = a[10] & g[3751];
assign g[7846] = b[10] & g[3751];
assign g[5800] = a[10] & g[3752];
assign g[7847] = b[10] & g[3752];
assign g[5801] = a[10] & g[3753];
assign g[7848] = b[10] & g[3753];
assign g[5802] = a[10] & g[3754];
assign g[7849] = b[10] & g[3754];
assign g[5803] = a[10] & g[3755];
assign g[7850] = b[10] & g[3755];
assign g[5804] = a[10] & g[3756];
assign g[7851] = b[10] & g[3756];
assign g[5805] = a[10] & g[3757];
assign g[7852] = b[10] & g[3757];
assign g[5806] = a[10] & g[3758];
assign g[7853] = b[10] & g[3758];
assign g[5807] = a[10] & g[3759];
assign g[7854] = b[10] & g[3759];
assign g[5808] = a[10] & g[3760];
assign g[7855] = b[10] & g[3760];
assign g[5809] = a[10] & g[3761];
assign g[7856] = b[10] & g[3761];
assign g[5810] = a[10] & g[3762];
assign g[7857] = b[10] & g[3762];
assign g[5811] = a[10] & g[3763];
assign g[7858] = b[10] & g[3763];
assign g[5812] = a[10] & g[3764];
assign g[7859] = b[10] & g[3764];
assign g[5813] = a[10] & g[3765];
assign g[7860] = b[10] & g[3765];
assign g[5814] = a[10] & g[3766];
assign g[7861] = b[10] & g[3766];
assign g[5815] = a[10] & g[3767];
assign g[7862] = b[10] & g[3767];
assign g[5816] = a[10] & g[3768];
assign g[7863] = b[10] & g[3768];
assign g[5817] = a[10] & g[3769];
assign g[7864] = b[10] & g[3769];
assign g[5818] = a[10] & g[3770];
assign g[7865] = b[10] & g[3770];
assign g[5819] = a[10] & g[3771];
assign g[7866] = b[10] & g[3771];
assign g[5820] = a[10] & g[3772];
assign g[7867] = b[10] & g[3772];
assign g[5821] = a[10] & g[3773];
assign g[7868] = b[10] & g[3773];
assign g[5822] = a[10] & g[3774];
assign g[7869] = b[10] & g[3774];
assign g[5823] = a[10] & g[3775];
assign g[7870] = b[10] & g[3775];
assign g[5824] = a[10] & g[3776];
assign g[7871] = b[10] & g[3776];
assign g[5825] = a[10] & g[3777];
assign g[7872] = b[10] & g[3777];
assign g[5826] = a[10] & g[3778];
assign g[7873] = b[10] & g[3778];
assign g[5827] = a[10] & g[3779];
assign g[7874] = b[10] & g[3779];
assign g[5828] = a[10] & g[3780];
assign g[7875] = b[10] & g[3780];
assign g[5829] = a[10] & g[3781];
assign g[7876] = b[10] & g[3781];
assign g[5830] = a[10] & g[3782];
assign g[7877] = b[10] & g[3782];
assign g[5831] = a[10] & g[3783];
assign g[7878] = b[10] & g[3783];
assign g[5832] = a[10] & g[3784];
assign g[7879] = b[10] & g[3784];
assign g[5833] = a[10] & g[3785];
assign g[7880] = b[10] & g[3785];
assign g[5834] = a[10] & g[3786];
assign g[7881] = b[10] & g[3786];
assign g[5835] = a[10] & g[3787];
assign g[7882] = b[10] & g[3787];
assign g[5836] = a[10] & g[3788];
assign g[7883] = b[10] & g[3788];
assign g[5837] = a[10] & g[3789];
assign g[7884] = b[10] & g[3789];
assign g[5838] = a[10] & g[3790];
assign g[7885] = b[10] & g[3790];
assign g[5839] = a[10] & g[3791];
assign g[7886] = b[10] & g[3791];
assign g[5840] = a[10] & g[3792];
assign g[7887] = b[10] & g[3792];
assign g[5841] = a[10] & g[3793];
assign g[7888] = b[10] & g[3793];
assign g[5842] = a[10] & g[3794];
assign g[7889] = b[10] & g[3794];
assign g[5843] = a[10] & g[3795];
assign g[7890] = b[10] & g[3795];
assign g[5844] = a[10] & g[3796];
assign g[7891] = b[10] & g[3796];
assign g[5845] = a[10] & g[3797];
assign g[7892] = b[10] & g[3797];
assign g[5846] = a[10] & g[3798];
assign g[7893] = b[10] & g[3798];
assign g[5847] = a[10] & g[3799];
assign g[7894] = b[10] & g[3799];
assign g[5848] = a[10] & g[3800];
assign g[7895] = b[10] & g[3800];
assign g[5849] = a[10] & g[3801];
assign g[7896] = b[10] & g[3801];
assign g[5850] = a[10] & g[3802];
assign g[7897] = b[10] & g[3802];
assign g[5851] = a[10] & g[3803];
assign g[7898] = b[10] & g[3803];
assign g[5852] = a[10] & g[3804];
assign g[7899] = b[10] & g[3804];
assign g[5853] = a[10] & g[3805];
assign g[7900] = b[10] & g[3805];
assign g[5854] = a[10] & g[3806];
assign g[7901] = b[10] & g[3806];
assign g[5855] = a[10] & g[3807];
assign g[7902] = b[10] & g[3807];
assign g[5856] = a[10] & g[3808];
assign g[7903] = b[10] & g[3808];
assign g[5857] = a[10] & g[3809];
assign g[7904] = b[10] & g[3809];
assign g[5858] = a[10] & g[3810];
assign g[7905] = b[10] & g[3810];
assign g[5859] = a[10] & g[3811];
assign g[7906] = b[10] & g[3811];
assign g[5860] = a[10] & g[3812];
assign g[7907] = b[10] & g[3812];
assign g[5861] = a[10] & g[3813];
assign g[7908] = b[10] & g[3813];
assign g[5862] = a[10] & g[3814];
assign g[7909] = b[10] & g[3814];
assign g[5863] = a[10] & g[3815];
assign g[7910] = b[10] & g[3815];
assign g[5864] = a[10] & g[3816];
assign g[7911] = b[10] & g[3816];
assign g[5865] = a[10] & g[3817];
assign g[7912] = b[10] & g[3817];
assign g[5866] = a[10] & g[3818];
assign g[7913] = b[10] & g[3818];
assign g[5867] = a[10] & g[3819];
assign g[7914] = b[10] & g[3819];
assign g[5868] = a[10] & g[3820];
assign g[7915] = b[10] & g[3820];
assign g[5869] = a[10] & g[3821];
assign g[7916] = b[10] & g[3821];
assign g[5870] = a[10] & g[3822];
assign g[7917] = b[10] & g[3822];
assign g[5871] = a[10] & g[3823];
assign g[7918] = b[10] & g[3823];
assign g[5872] = a[10] & g[3824];
assign g[7919] = b[10] & g[3824];
assign g[5873] = a[10] & g[3825];
assign g[7920] = b[10] & g[3825];
assign g[5874] = a[10] & g[3826];
assign g[7921] = b[10] & g[3826];
assign g[5875] = a[10] & g[3827];
assign g[7922] = b[10] & g[3827];
assign g[5876] = a[10] & g[3828];
assign g[7923] = b[10] & g[3828];
assign g[5877] = a[10] & g[3829];
assign g[7924] = b[10] & g[3829];
assign g[5878] = a[10] & g[3830];
assign g[7925] = b[10] & g[3830];
assign g[5879] = a[10] & g[3831];
assign g[7926] = b[10] & g[3831];
assign g[5880] = a[10] & g[3832];
assign g[7927] = b[10] & g[3832];
assign g[5881] = a[10] & g[3833];
assign g[7928] = b[10] & g[3833];
assign g[5882] = a[10] & g[3834];
assign g[7929] = b[10] & g[3834];
assign g[5883] = a[10] & g[3835];
assign g[7930] = b[10] & g[3835];
assign g[5884] = a[10] & g[3836];
assign g[7931] = b[10] & g[3836];
assign g[5885] = a[10] & g[3837];
assign g[7932] = b[10] & g[3837];
assign g[5886] = a[10] & g[3838];
assign g[7933] = b[10] & g[3838];
assign g[5887] = a[10] & g[3839];
assign g[7934] = b[10] & g[3839];
assign g[5888] = a[10] & g[3840];
assign g[7935] = b[10] & g[3840];
assign g[5889] = a[10] & g[3841];
assign g[7936] = b[10] & g[3841];
assign g[5890] = a[10] & g[3842];
assign g[7937] = b[10] & g[3842];
assign g[5891] = a[10] & g[3843];
assign g[7938] = b[10] & g[3843];
assign g[5892] = a[10] & g[3844];
assign g[7939] = b[10] & g[3844];
assign g[5893] = a[10] & g[3845];
assign g[7940] = b[10] & g[3845];
assign g[5894] = a[10] & g[3846];
assign g[7941] = b[10] & g[3846];
assign g[5895] = a[10] & g[3847];
assign g[7942] = b[10] & g[3847];
assign g[5896] = a[10] & g[3848];
assign g[7943] = b[10] & g[3848];
assign g[5897] = a[10] & g[3849];
assign g[7944] = b[10] & g[3849];
assign g[5898] = a[10] & g[3850];
assign g[7945] = b[10] & g[3850];
assign g[5899] = a[10] & g[3851];
assign g[7946] = b[10] & g[3851];
assign g[5900] = a[10] & g[3852];
assign g[7947] = b[10] & g[3852];
assign g[5901] = a[10] & g[3853];
assign g[7948] = b[10] & g[3853];
assign g[5902] = a[10] & g[3854];
assign g[7949] = b[10] & g[3854];
assign g[5903] = a[10] & g[3855];
assign g[7950] = b[10] & g[3855];
assign g[5904] = a[10] & g[3856];
assign g[7951] = b[10] & g[3856];
assign g[5905] = a[10] & g[3857];
assign g[7952] = b[10] & g[3857];
assign g[5906] = a[10] & g[3858];
assign g[7953] = b[10] & g[3858];
assign g[5907] = a[10] & g[3859];
assign g[7954] = b[10] & g[3859];
assign g[5908] = a[10] & g[3860];
assign g[7955] = b[10] & g[3860];
assign g[5909] = a[10] & g[3861];
assign g[7956] = b[10] & g[3861];
assign g[5910] = a[10] & g[3862];
assign g[7957] = b[10] & g[3862];
assign g[5911] = a[10] & g[3863];
assign g[7958] = b[10] & g[3863];
assign g[5912] = a[10] & g[3864];
assign g[7959] = b[10] & g[3864];
assign g[5913] = a[10] & g[3865];
assign g[7960] = b[10] & g[3865];
assign g[5914] = a[10] & g[3866];
assign g[7961] = b[10] & g[3866];
assign g[5915] = a[10] & g[3867];
assign g[7962] = b[10] & g[3867];
assign g[5916] = a[10] & g[3868];
assign g[7963] = b[10] & g[3868];
assign g[5917] = a[10] & g[3869];
assign g[7964] = b[10] & g[3869];
assign g[5918] = a[10] & g[3870];
assign g[7965] = b[10] & g[3870];
assign g[5919] = a[10] & g[3871];
assign g[7966] = b[10] & g[3871];
assign g[5920] = a[10] & g[3872];
assign g[7967] = b[10] & g[3872];
assign g[5921] = a[10] & g[3873];
assign g[7968] = b[10] & g[3873];
assign g[5922] = a[10] & g[3874];
assign g[7969] = b[10] & g[3874];
assign g[5923] = a[10] & g[3875];
assign g[7970] = b[10] & g[3875];
assign g[5924] = a[10] & g[3876];
assign g[7971] = b[10] & g[3876];
assign g[5925] = a[10] & g[3877];
assign g[7972] = b[10] & g[3877];
assign g[5926] = a[10] & g[3878];
assign g[7973] = b[10] & g[3878];
assign g[5927] = a[10] & g[3879];
assign g[7974] = b[10] & g[3879];
assign g[5928] = a[10] & g[3880];
assign g[7975] = b[10] & g[3880];
assign g[5929] = a[10] & g[3881];
assign g[7976] = b[10] & g[3881];
assign g[5930] = a[10] & g[3882];
assign g[7977] = b[10] & g[3882];
assign g[5931] = a[10] & g[3883];
assign g[7978] = b[10] & g[3883];
assign g[5932] = a[10] & g[3884];
assign g[7979] = b[10] & g[3884];
assign g[5933] = a[10] & g[3885];
assign g[7980] = b[10] & g[3885];
assign g[5934] = a[10] & g[3886];
assign g[7981] = b[10] & g[3886];
assign g[5935] = a[10] & g[3887];
assign g[7982] = b[10] & g[3887];
assign g[5936] = a[10] & g[3888];
assign g[7983] = b[10] & g[3888];
assign g[5937] = a[10] & g[3889];
assign g[7984] = b[10] & g[3889];
assign g[5938] = a[10] & g[3890];
assign g[7985] = b[10] & g[3890];
assign g[5939] = a[10] & g[3891];
assign g[7986] = b[10] & g[3891];
assign g[5940] = a[10] & g[3892];
assign g[7987] = b[10] & g[3892];
assign g[5941] = a[10] & g[3893];
assign g[7988] = b[10] & g[3893];
assign g[5942] = a[10] & g[3894];
assign g[7989] = b[10] & g[3894];
assign g[5943] = a[10] & g[3895];
assign g[7990] = b[10] & g[3895];
assign g[5944] = a[10] & g[3896];
assign g[7991] = b[10] & g[3896];
assign g[5945] = a[10] & g[3897];
assign g[7992] = b[10] & g[3897];
assign g[5946] = a[10] & g[3898];
assign g[7993] = b[10] & g[3898];
assign g[5947] = a[10] & g[3899];
assign g[7994] = b[10] & g[3899];
assign g[5948] = a[10] & g[3900];
assign g[7995] = b[10] & g[3900];
assign g[5949] = a[10] & g[3901];
assign g[7996] = b[10] & g[3901];
assign g[5950] = a[10] & g[3902];
assign g[7997] = b[10] & g[3902];
assign g[5951] = a[10] & g[3903];
assign g[7998] = b[10] & g[3903];
assign g[5952] = a[10] & g[3904];
assign g[7999] = b[10] & g[3904];
assign g[5953] = a[10] & g[3905];
assign g[8000] = b[10] & g[3905];
assign g[5954] = a[10] & g[3906];
assign g[8001] = b[10] & g[3906];
assign g[5955] = a[10] & g[3907];
assign g[8002] = b[10] & g[3907];
assign g[5956] = a[10] & g[3908];
assign g[8003] = b[10] & g[3908];
assign g[5957] = a[10] & g[3909];
assign g[8004] = b[10] & g[3909];
assign g[5958] = a[10] & g[3910];
assign g[8005] = b[10] & g[3910];
assign g[5959] = a[10] & g[3911];
assign g[8006] = b[10] & g[3911];
assign g[5960] = a[10] & g[3912];
assign g[8007] = b[10] & g[3912];
assign g[5961] = a[10] & g[3913];
assign g[8008] = b[10] & g[3913];
assign g[5962] = a[10] & g[3914];
assign g[8009] = b[10] & g[3914];
assign g[5963] = a[10] & g[3915];
assign g[8010] = b[10] & g[3915];
assign g[5964] = a[10] & g[3916];
assign g[8011] = b[10] & g[3916];
assign g[5965] = a[10] & g[3917];
assign g[8012] = b[10] & g[3917];
assign g[5966] = a[10] & g[3918];
assign g[8013] = b[10] & g[3918];
assign g[5967] = a[10] & g[3919];
assign g[8014] = b[10] & g[3919];
assign g[5968] = a[10] & g[3920];
assign g[8015] = b[10] & g[3920];
assign g[5969] = a[10] & g[3921];
assign g[8016] = b[10] & g[3921];
assign g[5970] = a[10] & g[3922];
assign g[8017] = b[10] & g[3922];
assign g[5971] = a[10] & g[3923];
assign g[8018] = b[10] & g[3923];
assign g[5972] = a[10] & g[3924];
assign g[8019] = b[10] & g[3924];
assign g[5973] = a[10] & g[3925];
assign g[8020] = b[10] & g[3925];
assign g[5974] = a[10] & g[3926];
assign g[8021] = b[10] & g[3926];
assign g[5975] = a[10] & g[3927];
assign g[8022] = b[10] & g[3927];
assign g[5976] = a[10] & g[3928];
assign g[8023] = b[10] & g[3928];
assign g[5977] = a[10] & g[3929];
assign g[8024] = b[10] & g[3929];
assign g[5978] = a[10] & g[3930];
assign g[8025] = b[10] & g[3930];
assign g[5979] = a[10] & g[3931];
assign g[8026] = b[10] & g[3931];
assign g[5980] = a[10] & g[3932];
assign g[8027] = b[10] & g[3932];
assign g[5981] = a[10] & g[3933];
assign g[8028] = b[10] & g[3933];
assign g[5982] = a[10] & g[3934];
assign g[8029] = b[10] & g[3934];
assign g[5983] = a[10] & g[3935];
assign g[8030] = b[10] & g[3935];
assign g[5984] = a[10] & g[3936];
assign g[8031] = b[10] & g[3936];
assign g[5985] = a[10] & g[3937];
assign g[8032] = b[10] & g[3937];
assign g[5986] = a[10] & g[3938];
assign g[8033] = b[10] & g[3938];
assign g[5987] = a[10] & g[3939];
assign g[8034] = b[10] & g[3939];
assign g[5988] = a[10] & g[3940];
assign g[8035] = b[10] & g[3940];
assign g[5989] = a[10] & g[3941];
assign g[8036] = b[10] & g[3941];
assign g[5990] = a[10] & g[3942];
assign g[8037] = b[10] & g[3942];
assign g[5991] = a[10] & g[3943];
assign g[8038] = b[10] & g[3943];
assign g[5992] = a[10] & g[3944];
assign g[8039] = b[10] & g[3944];
assign g[5993] = a[10] & g[3945];
assign g[8040] = b[10] & g[3945];
assign g[5994] = a[10] & g[3946];
assign g[8041] = b[10] & g[3946];
assign g[5995] = a[10] & g[3947];
assign g[8042] = b[10] & g[3947];
assign g[5996] = a[10] & g[3948];
assign g[8043] = b[10] & g[3948];
assign g[5997] = a[10] & g[3949];
assign g[8044] = b[10] & g[3949];
assign g[5998] = a[10] & g[3950];
assign g[8045] = b[10] & g[3950];
assign g[5999] = a[10] & g[3951];
assign g[8046] = b[10] & g[3951];
assign g[6000] = a[10] & g[3952];
assign g[8047] = b[10] & g[3952];
assign g[6001] = a[10] & g[3953];
assign g[8048] = b[10] & g[3953];
assign g[6002] = a[10] & g[3954];
assign g[8049] = b[10] & g[3954];
assign g[6003] = a[10] & g[3955];
assign g[8050] = b[10] & g[3955];
assign g[6004] = a[10] & g[3956];
assign g[8051] = b[10] & g[3956];
assign g[6005] = a[10] & g[3957];
assign g[8052] = b[10] & g[3957];
assign g[6006] = a[10] & g[3958];
assign g[8053] = b[10] & g[3958];
assign g[6007] = a[10] & g[3959];
assign g[8054] = b[10] & g[3959];
assign g[6008] = a[10] & g[3960];
assign g[8055] = b[10] & g[3960];
assign g[6009] = a[10] & g[3961];
assign g[8056] = b[10] & g[3961];
assign g[6010] = a[10] & g[3962];
assign g[8057] = b[10] & g[3962];
assign g[6011] = a[10] & g[3963];
assign g[8058] = b[10] & g[3963];
assign g[6012] = a[10] & g[3964];
assign g[8059] = b[10] & g[3964];
assign g[6013] = a[10] & g[3965];
assign g[8060] = b[10] & g[3965];
assign g[6014] = a[10] & g[3966];
assign g[8061] = b[10] & g[3966];
assign g[6015] = a[10] & g[3967];
assign g[8062] = b[10] & g[3967];
assign g[6016] = a[10] & g[3968];
assign g[8063] = b[10] & g[3968];
assign g[6017] = a[10] & g[3969];
assign g[8064] = b[10] & g[3969];
assign g[6018] = a[10] & g[3970];
assign g[8065] = b[10] & g[3970];
assign g[6019] = a[10] & g[3971];
assign g[8066] = b[10] & g[3971];
assign g[6020] = a[10] & g[3972];
assign g[8067] = b[10] & g[3972];
assign g[6021] = a[10] & g[3973];
assign g[8068] = b[10] & g[3973];
assign g[6022] = a[10] & g[3974];
assign g[8069] = b[10] & g[3974];
assign g[6023] = a[10] & g[3975];
assign g[8070] = b[10] & g[3975];
assign g[6024] = a[10] & g[3976];
assign g[8071] = b[10] & g[3976];
assign g[6025] = a[10] & g[3977];
assign g[8072] = b[10] & g[3977];
assign g[6026] = a[10] & g[3978];
assign g[8073] = b[10] & g[3978];
assign g[6027] = a[10] & g[3979];
assign g[8074] = b[10] & g[3979];
assign g[6028] = a[10] & g[3980];
assign g[8075] = b[10] & g[3980];
assign g[6029] = a[10] & g[3981];
assign g[8076] = b[10] & g[3981];
assign g[6030] = a[10] & g[3982];
assign g[8077] = b[10] & g[3982];
assign g[6031] = a[10] & g[3983];
assign g[8078] = b[10] & g[3983];
assign g[6032] = a[10] & g[3984];
assign g[8079] = b[10] & g[3984];
assign g[6033] = a[10] & g[3985];
assign g[8080] = b[10] & g[3985];
assign g[6034] = a[10] & g[3986];
assign g[8081] = b[10] & g[3986];
assign g[6035] = a[10] & g[3987];
assign g[8082] = b[10] & g[3987];
assign g[6036] = a[10] & g[3988];
assign g[8083] = b[10] & g[3988];
assign g[6037] = a[10] & g[3989];
assign g[8084] = b[10] & g[3989];
assign g[6038] = a[10] & g[3990];
assign g[8085] = b[10] & g[3990];
assign g[6039] = a[10] & g[3991];
assign g[8086] = b[10] & g[3991];
assign g[6040] = a[10] & g[3992];
assign g[8087] = b[10] & g[3992];
assign g[6041] = a[10] & g[3993];
assign g[8088] = b[10] & g[3993];
assign g[6042] = a[10] & g[3994];
assign g[8089] = b[10] & g[3994];
assign g[6043] = a[10] & g[3995];
assign g[8090] = b[10] & g[3995];
assign g[6044] = a[10] & g[3996];
assign g[8091] = b[10] & g[3996];
assign g[6045] = a[10] & g[3997];
assign g[8092] = b[10] & g[3997];
assign g[6046] = a[10] & g[3998];
assign g[8093] = b[10] & g[3998];
assign g[6047] = a[10] & g[3999];
assign g[8094] = b[10] & g[3999];
assign g[6048] = a[10] & g[4000];
assign g[8095] = b[10] & g[4000];
assign g[6049] = a[10] & g[4001];
assign g[8096] = b[10] & g[4001];
assign g[6050] = a[10] & g[4002];
assign g[8097] = b[10] & g[4002];
assign g[6051] = a[10] & g[4003];
assign g[8098] = b[10] & g[4003];
assign g[6052] = a[10] & g[4004];
assign g[8099] = b[10] & g[4004];
assign g[6053] = a[10] & g[4005];
assign g[8100] = b[10] & g[4005];
assign g[6054] = a[10] & g[4006];
assign g[8101] = b[10] & g[4006];
assign g[6055] = a[10] & g[4007];
assign g[8102] = b[10] & g[4007];
assign g[6056] = a[10] & g[4008];
assign g[8103] = b[10] & g[4008];
assign g[6057] = a[10] & g[4009];
assign g[8104] = b[10] & g[4009];
assign g[6058] = a[10] & g[4010];
assign g[8105] = b[10] & g[4010];
assign g[6059] = a[10] & g[4011];
assign g[8106] = b[10] & g[4011];
assign g[6060] = a[10] & g[4012];
assign g[8107] = b[10] & g[4012];
assign g[6061] = a[10] & g[4013];
assign g[8108] = b[10] & g[4013];
assign g[6062] = a[10] & g[4014];
assign g[8109] = b[10] & g[4014];
assign g[6063] = a[10] & g[4015];
assign g[8110] = b[10] & g[4015];
assign g[6064] = a[10] & g[4016];
assign g[8111] = b[10] & g[4016];
assign g[6065] = a[10] & g[4017];
assign g[8112] = b[10] & g[4017];
assign g[6066] = a[10] & g[4018];
assign g[8113] = b[10] & g[4018];
assign g[6067] = a[10] & g[4019];
assign g[8114] = b[10] & g[4019];
assign g[6068] = a[10] & g[4020];
assign g[8115] = b[10] & g[4020];
assign g[6069] = a[10] & g[4021];
assign g[8116] = b[10] & g[4021];
assign g[6070] = a[10] & g[4022];
assign g[8117] = b[10] & g[4022];
assign g[6071] = a[10] & g[4023];
assign g[8118] = b[10] & g[4023];
assign g[6072] = a[10] & g[4024];
assign g[8119] = b[10] & g[4024];
assign g[6073] = a[10] & g[4025];
assign g[8120] = b[10] & g[4025];
assign g[6074] = a[10] & g[4026];
assign g[8121] = b[10] & g[4026];
assign g[6075] = a[10] & g[4027];
assign g[8122] = b[10] & g[4027];
assign g[6076] = a[10] & g[4028];
assign g[8123] = b[10] & g[4028];
assign g[6077] = a[10] & g[4029];
assign g[8124] = b[10] & g[4029];
assign g[6078] = a[10] & g[4030];
assign g[8125] = b[10] & g[4030];
assign g[6079] = a[10] & g[4031];
assign g[8126] = b[10] & g[4031];
assign g[6080] = a[10] & g[4032];
assign g[8127] = b[10] & g[4032];
assign g[6081] = a[10] & g[4033];
assign g[8128] = b[10] & g[4033];
assign g[6082] = a[10] & g[4034];
assign g[8129] = b[10] & g[4034];
assign g[6083] = a[10] & g[4035];
assign g[8130] = b[10] & g[4035];
assign g[6084] = a[10] & g[4036];
assign g[8131] = b[10] & g[4036];
assign g[6085] = a[10] & g[4037];
assign g[8132] = b[10] & g[4037];
assign g[6086] = a[10] & g[4038];
assign g[8133] = b[10] & g[4038];
assign g[6087] = a[10] & g[4039];
assign g[8134] = b[10] & g[4039];
assign g[6088] = a[10] & g[4040];
assign g[8135] = b[10] & g[4040];
assign g[6089] = a[10] & g[4041];
assign g[8136] = b[10] & g[4041];
assign g[6090] = a[10] & g[4042];
assign g[8137] = b[10] & g[4042];
assign g[6091] = a[10] & g[4043];
assign g[8138] = b[10] & g[4043];
assign g[6092] = a[10] & g[4044];
assign g[8139] = b[10] & g[4044];
assign g[6093] = a[10] & g[4045];
assign g[8140] = b[10] & g[4045];
assign g[6094] = a[10] & g[4046];
assign g[8141] = b[10] & g[4046];
assign g[6095] = a[10] & g[4047];
assign g[8142] = b[10] & g[4047];
assign g[6096] = a[10] & g[4048];
assign g[8143] = b[10] & g[4048];
assign g[6097] = a[10] & g[4049];
assign g[8144] = b[10] & g[4049];
assign g[6098] = a[10] & g[4050];
assign g[8145] = b[10] & g[4050];
assign g[6099] = a[10] & g[4051];
assign g[8146] = b[10] & g[4051];
assign g[6100] = a[10] & g[4052];
assign g[8147] = b[10] & g[4052];
assign g[6101] = a[10] & g[4053];
assign g[8148] = b[10] & g[4053];
assign g[6102] = a[10] & g[4054];
assign g[8149] = b[10] & g[4054];
assign g[6103] = a[10] & g[4055];
assign g[8150] = b[10] & g[4055];
assign g[6104] = a[10] & g[4056];
assign g[8151] = b[10] & g[4056];
assign g[6105] = a[10] & g[4057];
assign g[8152] = b[10] & g[4057];
assign g[6106] = a[10] & g[4058];
assign g[8153] = b[10] & g[4058];
assign g[6107] = a[10] & g[4059];
assign g[8154] = b[10] & g[4059];
assign g[6108] = a[10] & g[4060];
assign g[8155] = b[10] & g[4060];
assign g[6109] = a[10] & g[4061];
assign g[8156] = b[10] & g[4061];
assign g[6110] = a[10] & g[4062];
assign g[8157] = b[10] & g[4062];
assign g[6111] = a[10] & g[4063];
assign g[8158] = b[10] & g[4063];
assign g[6112] = a[10] & g[4064];
assign g[8159] = b[10] & g[4064];
assign g[6113] = a[10] & g[4065];
assign g[8160] = b[10] & g[4065];
assign g[6114] = a[10] & g[4066];
assign g[8161] = b[10] & g[4066];
assign g[6115] = a[10] & g[4067];
assign g[8162] = b[10] & g[4067];
assign g[6116] = a[10] & g[4068];
assign g[8163] = b[10] & g[4068];
assign g[6117] = a[10] & g[4069];
assign g[8164] = b[10] & g[4069];
assign g[6118] = a[10] & g[4070];
assign g[8165] = b[10] & g[4070];
assign g[6119] = a[10] & g[4071];
assign g[8166] = b[10] & g[4071];
assign g[6120] = a[10] & g[4072];
assign g[8167] = b[10] & g[4072];
assign g[6121] = a[10] & g[4073];
assign g[8168] = b[10] & g[4073];
assign g[6122] = a[10] & g[4074];
assign g[8169] = b[10] & g[4074];
assign g[6123] = a[10] & g[4075];
assign g[8170] = b[10] & g[4075];
assign g[6124] = a[10] & g[4076];
assign g[8171] = b[10] & g[4076];
assign g[6125] = a[10] & g[4077];
assign g[8172] = b[10] & g[4077];
assign g[6126] = a[10] & g[4078];
assign g[8173] = b[10] & g[4078];
assign g[6127] = a[10] & g[4079];
assign g[8174] = b[10] & g[4079];
assign g[6128] = a[10] & g[4080];
assign g[8175] = b[10] & g[4080];
assign g[6129] = a[10] & g[4081];
assign g[8176] = b[10] & g[4081];
assign g[6130] = a[10] & g[4082];
assign g[8177] = b[10] & g[4082];
assign n = g[8177:1]; //assign outputs
endmodule